

module b17_C_gen_AntiSAT_k_256_6 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214;

  OAI21_X1 U11242 ( .B1(n15097), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15104), .ZN(n12584) );
  OAI21_X2 U11243 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18877), .A(n16532), 
        .ZN(n17904) );
  NAND2_X1 U11244 ( .A1(n14925), .A2(n12140), .ZN(n12162) );
  OR2_X1 U11245 ( .A1(n14245), .A2(n11847), .ZN(n14651) );
  CLKBUF_X3 U11246 ( .A(n11856), .Z(n15908) );
  NAND3_X1 U11247 ( .A1(n14170), .A2(n14171), .A3(n14169), .ZN(n14176) );
  NAND2_X1 U11248 ( .A1(n12403), .A2(n19074), .ZN(n12427) );
  INV_X2 U11249 ( .A(n16891), .ZN(n9865) );
  NOR2_X1 U11250 ( .A1(n12404), .A2(n10211), .ZN(n9971) );
  INV_X1 U11251 ( .A(n17402), .ZN(n18272) );
  CLKBUF_X2 U11252 ( .A(n10625), .Z(n9798) );
  NOR2_X1 U11253 ( .A1(n9814), .A2(n12312), .ZN(n12334) );
  OAI22_X1 U11254 ( .A1(n13381), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11778), 
        .B2(n11834), .ZN(n11107) );
  INV_X2 U11256 ( .A(n17218), .ZN(n17206) );
  INV_X1 U11257 ( .A(n12307), .ZN(n12312) );
  INV_X2 U11258 ( .A(n19277), .ZN(n12592) );
  INV_X1 U11259 ( .A(n17150), .ZN(n15615) );
  AND2_X1 U11260 ( .A1(n12244), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10636) );
  AND2_X1 U11261 ( .A1(n10353), .A2(n16325), .ZN(n10648) );
  AND2_X1 U11262 ( .A1(n12599), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12004) );
  AND2_X1 U11263 ( .A1(n10387), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10670) );
  AND2_X1 U11264 ( .A1(n9802), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10671) );
  INV_X1 U11265 ( .A(n9850), .ZN(n12031) );
  INV_X1 U11266 ( .A(n12220), .ZN(n9815) );
  CLKBUF_X1 U11267 ( .A(n10974), .Z(n11540) );
  INV_X1 U11268 ( .A(n10240), .ZN(n17196) );
  INV_X1 U11270 ( .A(n20183), .ZN(n11036) );
  INV_X2 U11271 ( .A(n18689), .ZN(n18670) );
  NAND2_X1 U11272 ( .A1(n18839), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12686) );
  BUF_X1 U11273 ( .A(n11038), .Z(n13540) );
  AND2_X1 U11275 ( .A1(n10917), .A2(n10920), .ZN(n11092) );
  AND2_X1 U11276 ( .A1(n13737), .A2(n10918), .ZN(n11091) );
  INV_X1 U11277 ( .A(n19283), .ZN(n11930) );
  NAND2_X1 U11278 ( .A1(n15570), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12220) );
  OR2_X1 U11281 ( .A1(n14651), .A2(n11848), .ZN(n10252) );
  OR2_X1 U11282 ( .A1(n11287), .A2(n10175), .ZN(n11297) );
  AND2_X1 U11283 ( .A1(n10433), .A2(n10432), .ZN(n10434) );
  INV_X1 U11284 ( .A(n13020), .ZN(n13047) );
  AND2_X1 U11285 ( .A1(n12243), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10676) );
  AND3_X1 U11286 ( .A1(n9804), .A2(n19110), .A3(n9970), .ZN(n9829) );
  NAND2_X1 U11287 ( .A1(n12319), .A2(n19256), .ZN(n19492) );
  OAI21_X1 U11288 ( .B1(n14601), .B2(n11855), .A(n15908), .ZN(n14581) );
  OR2_X1 U11289 ( .A1(n10928), .A2(n10927), .ZN(n11034) );
  INV_X1 U11290 ( .A(n19292), .ZN(n10334) );
  CLKBUF_X2 U11291 ( .A(n10481), .Z(n10482) );
  CLKBUF_X2 U11292 ( .A(n12775), .Z(n9799) );
  INV_X1 U11293 ( .A(n12780), .ZN(n17214) );
  OR3_X1 U11294 ( .A1(n14671), .A2(n14667), .A3(n14262), .ZN(n14245) );
  NAND2_X1 U11295 ( .A1(n11287), .A2(n11278), .ZN(n13788) );
  NOR2_X1 U11297 ( .A1(n13933), .A2(n13934), .ZN(n15489) );
  INV_X1 U11298 ( .A(n19264), .ZN(n10431) );
  INV_X1 U11299 ( .A(n15140), .ZN(n12662) );
  NAND3_X1 U11300 ( .A1(n12462), .A2(n12469), .A3(n9854), .ZN(n15442) );
  XNOR2_X1 U11301 ( .A(n12656), .B(n12399), .ZN(n15517) );
  OR2_X1 U11302 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12683), .ZN(
        n10240) );
  OR2_X1 U11304 ( .A1(n16917), .A2(n12686), .ZN(n13841) );
  INV_X1 U11305 ( .A(n18267), .ZN(n12989) );
  NAND2_X1 U11306 ( .A1(n14601), .A2(n14630), .ZN(n14622) );
  MUX2_X1 U11307 ( .A(n14557), .B(n14556), .S(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(n11858) );
  INV_X1 U11308 ( .A(n19041), .ZN(n19076) );
  XNOR2_X1 U11309 ( .A(n12162), .B(n12163), .ZN(n14918) );
  NAND2_X1 U11310 ( .A1(n19259), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14818) );
  XNOR2_X1 U11311 ( .A(n12427), .B(n14181), .ZN(n14167) );
  INV_X1 U11312 ( .A(n16925), .ZN(n16912) );
  INV_X1 U11313 ( .A(n17740), .ZN(n17755) );
  INV_X1 U11314 ( .A(n20075), .ZN(n20109) );
  AND3_X2 U11315 ( .A1(n12787), .A2(n12786), .A3(n12785), .ZN(n10256) );
  NAND2_X1 U11317 ( .A1(n10442), .A2(n10434), .ZN(n10479) );
  BUF_X4 U11318 ( .A(n13115), .Z(n14326) );
  NAND2_X2 U11319 ( .A1(n11762), .A2(n13096), .ZN(n13115) );
  NOR3_X2 U11320 ( .A1(n14256), .A2(n21172), .A3(n15834), .ZN(n14447) );
  AND3_X1 U11321 ( .A1(n10588), .A2(n13446), .A3(n19292), .ZN(n10625) );
  AOI21_X2 U11322 ( .B1(n11949), .B2(n11948), .A(n11947), .ZN(n13413) );
  AND2_X2 U11323 ( .A1(n14487), .A2(n10177), .ZN(n14409) );
  NOR2_X4 U11324 ( .A1(n14494), .A2(n15792), .ZN(n14487) );
  NAND2_X2 U11325 ( .A1(n16933), .A2(n12687), .ZN(n16917) );
  NOR2_X2 U11326 ( .A1(n12682), .A2(n18670), .ZN(n12723) );
  INV_X1 U11327 ( .A(n17150), .ZN(n17222) );
  XNOR2_X2 U11328 ( .A(n13342), .B(n11943), .ZN(n13335) );
  NAND2_X2 U11329 ( .A1(n11937), .A2(n11936), .ZN(n13342) );
  NOR2_X2 U11330 ( .A1(n17778), .A2(n17934), .ZN(n12814) );
  CLKBUF_X3 U11331 ( .A(n12775), .Z(n9800) );
  AND2_X1 U11332 ( .A1(n15571), .A2(n10202), .ZN(n9801) );
  AND2_X1 U11333 ( .A1(n15571), .A2(n10202), .ZN(n9802) );
  NOR2_X1 U11334 ( .A1(n15129), .A2(n10195), .ZN(n15088) );
  CLKBUF_X1 U11335 ( .A(n15186), .Z(n15187) );
  OAI21_X1 U11336 ( .B1(n12648), .B2(n10884), .A(n19061), .ZN(n12460) );
  NOR2_X1 U11337 ( .A1(n14929), .A2(n14919), .ZN(n14920) );
  NAND2_X2 U11338 ( .A1(n17680), .A2(n17740), .ZN(n17899) );
  INV_X1 U11339 ( .A(n15055), .ZN(n15338) );
  INV_X2 U11340 ( .A(n17904), .ZN(n17891) );
  NAND2_X1 U11341 ( .A1(n18136), .A2(n17777), .ZN(n17811) );
  AND2_X1 U11342 ( .A1(n12335), .A2(n19256), .ZN(n12378) );
  AND2_X1 U11343 ( .A1(n12334), .A2(n12330), .ZN(n19785) );
  OR2_X1 U11344 ( .A1(n12809), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10113) );
  AND2_X1 U11345 ( .A1(n12334), .A2(n12333), .ZN(n19706) );
  AND2_X1 U11346 ( .A1(n12334), .A2(n12329), .ZN(n19675) );
  AND2_X1 U11347 ( .A1(n12334), .A2(n12313), .ZN(n19753) );
  OR2_X2 U11348 ( .A1(n9804), .A2(n12307), .ZN(n12332) );
  INV_X1 U11349 ( .A(n12312), .ZN(n19256) );
  NAND2_X1 U11350 ( .A1(n11938), .A2(n11939), .ZN(n10458) );
  AND3_X1 U11351 ( .A1(n10463), .A2(n10462), .A3(n10461), .ZN(n11950) );
  CLKBUF_X3 U11352 ( .A(n10479), .Z(n10480) );
  AND2_X1 U11354 ( .A1(n16363), .A2(n12273), .ZN(n10437) );
  NOR2_X2 U11355 ( .A1(n17418), .A2(n12772), .ZN(n12796) );
  NOR2_X1 U11356 ( .A1(n17623), .A2(n17624), .ZN(n17606) );
  AND2_X1 U11357 ( .A1(n12722), .A2(n12721), .ZN(n17418) );
  AOI211_X2 U11358 ( .C1(n17223), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n12883), .B(n12882), .ZN(n17286) );
  NAND2_X1 U11360 ( .A1(n10587), .A2(n11930), .ZN(n10417) );
  OR2_X1 U11361 ( .A1(n11030), .A2(n11038), .ZN(n11045) );
  NAND2_X1 U11362 ( .A1(n19283), .A2(n10407), .ZN(n10408) );
  BUF_X1 U11363 ( .A(n13100), .Z(n11762) );
  AND4_X1 U11364 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n12735) );
  INV_X1 U11365 ( .A(n12723), .ZN(n17150) );
  BUF_X2 U11366 ( .A(n11115), .Z(n11740) );
  CLKBUF_X2 U11367 ( .A(n11092), .Z(n11093) );
  INV_X4 U11368 ( .A(n13841), .ZN(n17219) );
  BUF_X2 U11369 ( .A(n11141), .Z(n11731) );
  INV_X4 U11370 ( .A(n17216), .ZN(n17175) );
  CLKBUF_X2 U11371 ( .A(n12053), .Z(n9808) );
  BUF_X2 U11372 ( .A(n11098), .Z(n11732) );
  OR3_X2 U11373 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n16917), .ZN(n12697) );
  INV_X4 U11374 ( .A(n17191), .ZN(n17229) );
  INV_X4 U11376 ( .A(n10239), .ZN(n9803) );
  OR2_X1 U11377 ( .A1(n12685), .A2(n12686), .ZN(n9849) );
  NOR3_X1 U11378 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n12685), .ZN(n12775) );
  AND2_X2 U11379 ( .A1(n10920), .A2(n10919), .ZN(n10974) );
  XNOR2_X1 U11380 ( .A(n11858), .B(n10114), .ZN(n14718) );
  AND2_X1 U11381 ( .A1(n9963), .A2(n9962), .ZN(n9961) );
  INV_X1 U11382 ( .A(n14372), .ZN(n14590) );
  OR2_X1 U11383 ( .A1(n14597), .A2(n15953), .ZN(n9963) );
  NAND2_X1 U11384 ( .A1(n12561), .A2(n12560), .ZN(n10024) );
  OR2_X1 U11385 ( .A1(n14370), .A2(n10183), .ZN(n9822) );
  XNOR2_X1 U11386 ( .A(n14396), .B(n14384), .ZN(n14597) );
  NAND2_X1 U11387 ( .A1(n14600), .A2(n10106), .ZN(n14583) );
  OAI21_X1 U11388 ( .B1(n9852), .B2(n9986), .A(n9984), .ZN(n15219) );
  OR2_X1 U11389 ( .A1(n15744), .A2(n17814), .ZN(n10095) );
  NOR2_X1 U11390 ( .A1(n15651), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15744) );
  AND2_X1 U11391 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12652), .ZN(
        n12647) );
  NAND2_X1 U11392 ( .A1(n12426), .A2(n12425), .ZN(n14168) );
  NAND2_X1 U11393 ( .A1(n15517), .A2(n15527), .ZN(n12652) );
  XNOR2_X1 U11394 ( .A(n12657), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15505) );
  XOR2_X1 U11395 ( .A(n12668), .B(n12667), .Z(n16092) );
  XNOR2_X1 U11396 ( .A(n12460), .B(n15542), .ZN(n15243) );
  CLKBUF_X1 U11397 ( .A(n11364), .Z(n14131) );
  NAND2_X1 U11398 ( .A1(n9952), .A2(n14181), .ZN(n14171) );
  AND2_X1 U11399 ( .A1(n14920), .A2(n10150), .ZN(n14897) );
  NAND2_X1 U11400 ( .A1(n12410), .A2(n13975), .ZN(n15550) );
  NOR3_X1 U11401 ( .A1(n10252), .A2(n10108), .A3(n10112), .ZN(n10107) );
  NOR2_X1 U11402 ( .A1(n10252), .A2(n10112), .ZN(n10109) );
  OR2_X1 U11403 ( .A1(n14842), .A2(n14927), .ZN(n14929) );
  AND2_X1 U11404 ( .A1(n12085), .A2(n12108), .ZN(n12086) );
  AND2_X1 U11405 ( .A1(n12406), .A2(n12635), .ZN(n12630) );
  OR2_X1 U11406 ( .A1(n15005), .A2(n14833), .ZN(n15264) );
  AND2_X1 U11407 ( .A1(n14025), .A2(n14026), .ZN(n11315) );
  AND2_X1 U11408 ( .A1(n17675), .A2(n13003), .ZN(n17602) );
  NAND2_X1 U11409 ( .A1(n17599), .A2(n17598), .ZN(n17597) );
  NAND2_X1 U11410 ( .A1(n9960), .A2(n13956), .ZN(n9959) );
  AND2_X1 U11411 ( .A1(n9872), .A2(n10013), .ZN(n17599) );
  AND2_X1 U11412 ( .A1(n11856), .A2(n14270), .ZN(n14667) );
  NAND2_X2 U11413 ( .A1(n14120), .A2(n11988), .ZN(n14121) );
  NOR2_X1 U11414 ( .A1(n14987), .A2(n14860), .ZN(n14977) );
  NAND2_X1 U11415 ( .A1(n17767), .A2(n17966), .ZN(n17705) );
  NOR2_X1 U11416 ( .A1(n17683), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17682) );
  NAND2_X1 U11417 ( .A1(n10199), .A2(n12364), .ZN(n12404) );
  NOR2_X2 U11418 ( .A1(n14053), .A2(n14054), .ZN(n14076) );
  AND2_X1 U11419 ( .A1(n15793), .A2(n10144), .ZN(n14425) );
  NOR2_X1 U11420 ( .A1(n15406), .A2(n9884), .ZN(n15062) );
  NOR2_X2 U11421 ( .A1(n18244), .A2(n16532), .ZN(n17897) );
  AND2_X2 U11422 ( .A1(n12335), .A2(n15594), .ZN(n19330) );
  AOI22_X1 U11423 ( .A1(n19675), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12386), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12339) );
  CLKBUF_X1 U11424 ( .A(n14505), .Z(n15893) );
  NAND2_X1 U11425 ( .A1(n9829), .A2(n19256), .ZN(n12368) );
  OR2_X1 U11426 ( .A1(n11971), .A2(n13415), .ZN(n13416) );
  NAND2_X1 U11427 ( .A1(n15594), .A2(n12319), .ZN(n19361) );
  NAND2_X1 U11428 ( .A1(n12316), .A2(n19256), .ZN(n19427) );
  AND2_X1 U11429 ( .A1(n9858), .A2(n15569), .ZN(n12335) );
  NAND2_X1 U11430 ( .A1(n12316), .A2(n15594), .ZN(n19301) );
  NAND2_X1 U11431 ( .A1(n11189), .A2(n11188), .ZN(n13791) );
  AND2_X1 U11432 ( .A1(n10179), .A2(n10178), .ZN(n10177) );
  NOR2_X1 U11433 ( .A1(n14472), .A2(n14226), .ZN(n14330) );
  CLKBUF_X2 U11434 ( .A(n13421), .Z(n9814) );
  NAND2_X1 U11435 ( .A1(n15489), .A2(n15490), .ZN(n15491) );
  BUF_X2 U11436 ( .A(n13421), .Z(n9804) );
  CLKBUF_X1 U11437 ( .A(n14802), .Z(n20493) );
  NAND2_X1 U11438 ( .A1(n11959), .A2(n11958), .ZN(n11960) );
  AOI21_X1 U11439 ( .B1(n15569), .B2(n11964), .A(n11942), .ZN(n13334) );
  NAND2_X1 U11440 ( .A1(n15536), .A2(n10748), .ZN(n13961) );
  AND2_X1 U11441 ( .A1(n11939), .A2(n11935), .ZN(n15564) );
  NAND2_X1 U11442 ( .A1(n11157), .A2(n11156), .ZN(n20231) );
  NAND2_X1 U11443 ( .A1(n12992), .A2(n12982), .ZN(n15641) );
  NAND2_X2 U11444 ( .A1(n11911), .A2(n11910), .ZN(n15707) );
  NAND2_X1 U11445 ( .A1(n10460), .A2(n10459), .ZN(n11953) );
  NAND2_X1 U11446 ( .A1(n10186), .A2(n10428), .ZN(n10455) );
  NAND2_X1 U11447 ( .A1(n10470), .A2(n10469), .ZN(n10476) );
  AND2_X1 U11448 ( .A1(n11110), .A2(n11108), .ZN(n11155) );
  NAND2_X1 U11449 ( .A1(n11066), .A2(n11065), .ZN(n11110) );
  NAND2_X1 U11450 ( .A1(n17861), .A2(n12798), .ZN(n12801) );
  AOI21_X1 U11451 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20169), .A(
        n11905), .ZN(n11906) );
  NOR2_X1 U11452 ( .A1(n16386), .A2(n18662), .ZN(n18137) );
  NAND2_X1 U11453 ( .A1(n12594), .A2(n9855), .ZN(n12487) );
  NOR2_X1 U11454 ( .A1(n13315), .A2(n10669), .ZN(n13976) );
  INV_X2 U11455 ( .A(n17275), .ZN(n17266) );
  AND3_X1 U11456 ( .A1(n10473), .A2(n10472), .A3(n10471), .ZN(n10474) );
  OR2_X1 U11457 ( .A1(n10669), .A2(n10664), .ZN(n13314) );
  NAND2_X2 U11458 ( .A1(n16386), .A2(n16427), .ZN(n17777) );
  AOI21_X1 U11459 ( .B1(n10662), .B2(n9851), .A(n10663), .ZN(n10669) );
  CLKBUF_X1 U11460 ( .A(n13056), .Z(n15587) );
  NAND2_X1 U11461 ( .A1(n17885), .A2(n12790), .ZN(n12792) );
  NAND2_X1 U11462 ( .A1(n12286), .A2(n10436), .ZN(n13056) );
  NAND2_X1 U11463 ( .A1(n13077), .A2(n12273), .ZN(n10450) );
  NAND2_X1 U11464 ( .A1(n17886), .A2(n17887), .ZN(n17885) );
  AND2_X1 U11465 ( .A1(n10406), .A2(n13050), .ZN(n10447) );
  CLKBUF_X1 U11466 ( .A(n11047), .Z(n11048) );
  NAND2_X1 U11467 ( .A1(n10437), .A2(n19264), .ZN(n10505) );
  AND2_X1 U11468 ( .A1(n13285), .A2(n13286), .ZN(n10646) );
  AND2_X1 U11469 ( .A1(n10422), .A2(n10421), .ZN(n13077) );
  NOR2_X1 U11470 ( .A1(n12411), .A2(n12407), .ZN(n12422) );
  NAND2_X1 U11471 ( .A1(n10611), .A2(n10610), .ZN(n13285) );
  NAND2_X1 U11472 ( .A1(n13131), .A2(n14326), .ZN(n14324) );
  XNOR2_X1 U11473 ( .A(n12789), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17887) );
  NAND2_X1 U11474 ( .A1(n13644), .A2(n14326), .ZN(n13168) );
  AND3_X2 U11475 ( .A1(n10420), .A2(n10429), .A3(n10419), .ZN(n16363) );
  NOR2_X1 U11476 ( .A1(n10256), .A2(n18859), .ZN(n17903) );
  AND2_X1 U11477 ( .A1(n9969), .A2(n10334), .ZN(n9967) );
  AND2_X1 U11478 ( .A1(n10149), .A2(n10402), .ZN(n13226) );
  AND3_X1 U11479 ( .A1(n12895), .A2(n12894), .A3(n10248), .ZN(n17402) );
  NAND2_X1 U11480 ( .A1(n10149), .A2(n10420), .ZN(n13088) );
  NAND2_X2 U11481 ( .A1(n11174), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11907) );
  NAND3_X1 U11482 ( .A1(n13397), .A2(n20209), .A3(n11067), .ZN(n13746) );
  INV_X1 U11483 ( .A(n20819), .ZN(n11838) );
  INV_X1 U11484 ( .A(n13035), .ZN(n10436) );
  INV_X1 U11485 ( .A(n14818), .ZN(n12273) );
  CLKBUF_X1 U11486 ( .A(n11930), .Z(n13668) );
  OR2_X1 U11487 ( .A1(n20183), .A2(n13557), .ZN(n20822) );
  OR2_X1 U11488 ( .A1(n12750), .A2(n12749), .ZN(n17423) );
  NAND2_X1 U11489 ( .A1(n20215), .A2(n11031), .ZN(n11049) );
  CLKBUF_X1 U11490 ( .A(n11039), .Z(n20209) );
  INV_X1 U11491 ( .A(n10407), .ZN(n10587) );
  AND2_X2 U11492 ( .A1(n13557), .A2(n13096), .ZN(n13644) );
  NAND2_X1 U11493 ( .A1(n11032), .A2(n11231), .ZN(n11040) );
  OR2_X2 U11494 ( .A1(n16485), .A2(n16441), .ZN(n16488) );
  OR2_X1 U11495 ( .A1(n10971), .A2(n10970), .ZN(n13100) );
  NAND2_X1 U11496 ( .A1(n10386), .A2(n10385), .ZN(n9953) );
  NAND2_X1 U11497 ( .A1(n10347), .A2(n10346), .ZN(n10407) );
  NAND4_X2 U11498 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(
        n13096) );
  INV_X2 U11499 ( .A(U214), .ZN(n16485) );
  NAND2_X1 U11500 ( .A1(n10358), .A2(n16325), .ZN(n10359) );
  AND4_X1 U11501 ( .A1(n10978), .A2(n10977), .A3(n10976), .A4(n10975), .ZN(
        n10983) );
  AND4_X1 U11502 ( .A1(n11021), .A2(n11020), .A3(n11019), .A4(n11018), .ZN(
        n11027) );
  AND4_X1 U11503 ( .A1(n11017), .A2(n11016), .A3(n11015), .A4(n11014), .ZN(
        n11028) );
  AND4_X1 U11504 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n11007) );
  AND4_X1 U11505 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11006) );
  AND3_X1 U11506 ( .A1(n10952), .A2(n10951), .A3(n10950), .ZN(n10957) );
  AND4_X1 U11507 ( .A1(n10932), .A2(n10931), .A3(n10930), .A4(n10929), .ZN(
        n10938) );
  NAND2_X2 U11508 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20000), .ZN(n19933) );
  BUF_X2 U11509 ( .A(n10973), .Z(n11203) );
  AND4_X1 U11510 ( .A1(n11004), .A2(n11003), .A3(n11002), .A4(n11001), .ZN(
        n11005) );
  BUF_X2 U11511 ( .A(n10961), .Z(n11638) );
  INV_X4 U11512 ( .A(n12737), .ZN(n17201) );
  AND2_X1 U11513 ( .A1(n10381), .A2(n10380), .ZN(n10383) );
  AND4_X1 U11514 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10366) );
  AND3_X1 U11515 ( .A1(n10949), .A2(n10948), .A3(n10947), .ZN(n10952) );
  AND4_X1 U11516 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10379) );
  INV_X2 U11517 ( .A(n18756), .ZN(n9805) );
  NAND2_X2 U11518 ( .A1(n18821), .A2(n18754), .ZN(n18805) );
  NAND2_X2 U11519 ( .A1(n20000), .A2(n19877), .ZN(n19937) );
  BUF_X2 U11520 ( .A(n17221), .Z(n17194) );
  AND2_X2 U11521 ( .A1(n9815), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10647) );
  AND2_X2 U11522 ( .A1(n9808), .A2(n16325), .ZN(n10634) );
  INV_X2 U11523 ( .A(n9849), .ZN(n17200) );
  AND2_X2 U11524 ( .A1(n9815), .A2(n16325), .ZN(n12073) );
  INV_X2 U11525 ( .A(n16521), .ZN(U215) );
  BUF_X2 U11526 ( .A(n11091), .Z(n11738) );
  INV_X1 U11527 ( .A(n12220), .ZN(n10374) );
  INV_X2 U11528 ( .A(n20001), .ZN(n20000) );
  CLKBUF_X2 U11529 ( .A(n12053), .Z(n12245) );
  AND2_X2 U11530 ( .A1(n10921), .A2(n10917), .ZN(n11141) );
  AND2_X2 U11531 ( .A1(n10917), .A2(n13393), .ZN(n11122) );
  NOR3_X1 U11532 ( .A1(n18849), .A2(n18839), .A3(n16917), .ZN(n12680) );
  INV_X1 U11533 ( .A(n12235), .ZN(n9807) );
  AND2_X2 U11534 ( .A1(n10387), .A2(n16325), .ZN(n10616) );
  OR2_X2 U11535 ( .A1(n12682), .A2(n12685), .ZN(n10239) );
  AND2_X2 U11536 ( .A1(n13393), .A2(n10922), .ZN(n11127) );
  AND2_X2 U11537 ( .A1(n11865), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10917) );
  AND2_X1 U11538 ( .A1(n10912), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10921) );
  AND2_X2 U11539 ( .A1(n10920), .A2(n10922), .ZN(n11098) );
  AND2_X2 U11540 ( .A1(n10919), .A2(n13393), .ZN(n10992) );
  AND2_X1 U11541 ( .A1(n10910), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13737) );
  NAND4_X1 U11542 ( .A1(n18849), .A2(n18839), .A3(n12687), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17191) );
  AND2_X2 U11543 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10922) );
  NOR2_X2 U11544 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10919) );
  CLKBUF_X1 U11545 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13751) );
  NAND2_X1 U11546 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18697) );
  AND2_X1 U11547 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10598) );
  INV_X4 U11548 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10202) );
  NOR2_X1 U11549 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10298) );
  AND2_X2 U11550 ( .A1(n11914), .A2(n11035), .ZN(n9809) );
  INV_X1 U11551 ( .A(n9809), .ZN(n13369) );
  NOR2_X2 U11552 ( .A1(n9959), .A2(n13899), .ZN(n13954) );
  XNOR2_X2 U11553 ( .A(n11297), .B(n11296), .ZN(n11805) );
  NAND2_X1 U11554 ( .A1(n10442), .A2(n10434), .ZN(n9810) );
  NAND2_X1 U11555 ( .A1(n10442), .A2(n10434), .ZN(n9811) );
  OAI21_X1 U11556 ( .B1(n9814), .B2(n12673), .A(n11969), .ZN(n11971) );
  NAND2_X2 U11557 ( .A1(n11277), .A2(n11253), .ZN(n11774) );
  AND2_X2 U11558 ( .A1(n11975), .A2(n9823), .ZN(n14120) );
  NOR2_X2 U11559 ( .A1(n15788), .A2(n14332), .ZN(n15766) );
  NOR2_X2 U11560 ( .A1(n14933), .A2(n12111), .ZN(n12138) );
  NOR2_X2 U11561 ( .A1(n14932), .A2(n14934), .ZN(n14933) );
  OR2_X1 U11562 ( .A1(n12656), .A2(n12399), .ZN(n12657) );
  AND4_X1 U11563 ( .A1(n10370), .A2(n10369), .A3(n10368), .A4(n10367), .ZN(
        n10371) );
  NAND2_X1 U11564 ( .A1(n11934), .A2(n11933), .ZN(n11939) );
  AND2_X1 U11565 ( .A1(n12244), .A2(n16325), .ZN(n10692) );
  NOR2_X1 U11566 ( .A1(n18670), .A2(n12686), .ZN(n9813) );
  AND2_X4 U11567 ( .A1(n10598), .A2(n15562), .ZN(n10335) );
  NOR3_X2 U11568 ( .A1(n14399), .A2(n10139), .A3(n13180), .ZN(n10141) );
  NOR2_X2 U11569 ( .A1(n13076), .A2(n12278), .ZN(n13038) );
  NAND4_X2 U11570 ( .A1(n10026), .A2(n10430), .A3(n12283), .A4(n10025), .ZN(
        n13076) );
  NOR2_X2 U11571 ( .A1(n15135), .A2(n9866), .ZN(n15097) );
  AND2_X2 U11572 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15571) );
  OAI211_X2 U11573 ( .C1(n12585), .C2(n15109), .A(n12584), .B(n15101), .ZN(
        n15086) );
  OAI211_X1 U11574 ( .C1(n11963), .C2(n11962), .A(n11961), .B(n11960), .ZN(
        n13421) );
  INV_X1 U11575 ( .A(n12307), .ZN(n15594) );
  XNOR2_X1 U11576 ( .A(n11938), .B(n11939), .ZN(n15569) );
  NOR2_X2 U11577 ( .A1(n14941), .A2(n14940), .ZN(n14939) );
  INV_X1 U11578 ( .A(n9815), .ZN(n9816) );
  INV_X2 U11579 ( .A(n15602), .ZN(n9817) );
  INV_X1 U11580 ( .A(n15602), .ZN(n9818) );
  NAND2_X2 U11581 ( .A1(n15571), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15602) );
  NOR2_X1 U11582 ( .A1(n11072), .A2(n9964), .ZN(n11058) );
  NAND2_X1 U11583 ( .A1(n9853), .A2(n9967), .ZN(n10412) );
  NAND4_X1 U11584 ( .A1(n11315), .A2(n13954), .A3(n14085), .A4(n14132), .ZN(
        n11364) );
  OR2_X1 U11585 ( .A1(n18839), .A2(n12683), .ZN(n10257) );
  NAND2_X1 U11586 ( .A1(n18272), .A2(n18252), .ZN(n12998) );
  NAND2_X1 U11587 ( .A1(n16551), .A2(n18244), .ZN(n12995) );
  CLKBUF_X1 U11588 ( .A(n11730), .Z(n11702) );
  OAI21_X1 U11589 ( .B1(n11903), .B2(n11202), .A(n11201), .ZN(n11286) );
  OAI211_X1 U11590 ( .C1(n20819), .C2(n20202), .A(n11044), .B(n13558), .ZN(
        n11072) );
  NAND2_X1 U11591 ( .A1(n11864), .A2(n11863), .ZN(n11874) );
  NAND2_X1 U11592 ( .A1(n12456), .A2(n12455), .ZN(n12644) );
  NAND2_X1 U11593 ( .A1(n14208), .A2(n14234), .ZN(n9956) );
  INV_X1 U11594 ( .A(n13916), .ZN(n9960) );
  CLKBUF_X1 U11595 ( .A(n11265), .Z(n13998) );
  NAND2_X1 U11596 ( .A1(n11034), .A2(n13557), .ZN(n11174) );
  NAND2_X1 U11597 ( .A1(n9837), .A2(n14975), .ZN(n10234) );
  NOR3_X1 U11598 ( .A1(n9821), .A2(n9896), .A3(n15018), .ZN(n10869) );
  INV_X1 U11599 ( .A(n15004), .ZN(n10079) );
  NOR2_X1 U11600 ( .A1(n14947), .A2(n10158), .ZN(n10157) );
  INV_X1 U11601 ( .A(n10159), .ZN(n10158) );
  AND2_X1 U11602 ( .A1(n12527), .A2(n15179), .ZN(n12528) );
  NAND2_X1 U11603 ( .A1(n13446), .A2(n10592), .ZN(n10841) );
  NOR2_X1 U11604 ( .A1(n10587), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U11606 ( .A1(n10087), .A2(n15451), .ZN(n10086) );
  INV_X1 U11607 ( .A(n15477), .ZN(n10087) );
  INV_X1 U11608 ( .A(n15501), .ZN(n12469) );
  INV_X1 U11609 ( .A(n12405), .ZN(n10212) );
  INV_X1 U11610 ( .A(n10841), .ZN(n10825) );
  NAND2_X1 U11611 ( .A1(n11927), .A2(n19979), .ZN(n11968) );
  AND2_X1 U11612 ( .A1(n18906), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U11613 ( .A1(n18849), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12682) );
  NAND2_X1 U11614 ( .A1(n16933), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12685) );
  OR3_X1 U11615 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18839), .A3(
        n18697), .ZN(n12715) );
  NOR2_X1 U11616 ( .A1(n12873), .A2(n12872), .ZN(n13798) );
  NOR2_X1 U11617 ( .A1(n15639), .A2(n18883), .ZN(n17435) );
  NOR2_X1 U11618 ( .A1(n13557), .A2(n13096), .ZN(n11067) );
  NOR2_X1 U11619 ( .A1(n10181), .A2(n13095), .ZN(n10180) );
  NAND2_X1 U11620 ( .A1(n10182), .A2(n14384), .ZN(n10181) );
  INV_X1 U11621 ( .A(n10183), .ZN(n10182) );
  NAND2_X1 U11622 ( .A1(n10886), .A2(n19277), .ZN(n12594) );
  INV_X1 U11623 ( .A(n11946), .ZN(n11947) );
  AND2_X1 U11624 ( .A1(n13019), .A2(n12617), .ZN(n12670) );
  CLKBUF_X2 U11625 ( .A(n10591), .Z(n13072) );
  OR2_X1 U11626 ( .A1(n10195), .A2(n15251), .ZN(n9946) );
  AND2_X1 U11627 ( .A1(n15376), .A2(n13301), .ZN(n16290) );
  NAND2_X1 U11628 ( .A1(n10325), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10332) );
  NAND2_X1 U11629 ( .A1(n12999), .A2(n18247), .ZN(n12980) );
  NAND2_X2 U11630 ( .A1(n18672), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n17218) );
  OR3_X1 U11631 ( .A1(n16529), .A2(n18880), .A3(n15642), .ZN(n15762) );
  NOR2_X1 U11632 ( .A1(n16412), .A2(n16589), .ZN(n16379) );
  AND2_X1 U11633 ( .A1(n16379), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16408) );
  NAND2_X1 U11634 ( .A1(n12988), .A2(n13000), .ZN(n12993) );
  INV_X1 U11635 ( .A(n12802), .ZN(n12800) );
  INV_X1 U11636 ( .A(n18247), .ZN(n12979) );
  NAND2_X1 U11637 ( .A1(n10071), .A2(n10069), .ZN(n18244) );
  NOR2_X1 U11638 ( .A1(n12860), .A2(n10070), .ZN(n10069) );
  INV_X1 U11639 ( .A(n12859), .ZN(n10071) );
  AND2_X1 U11640 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10070) );
  INV_X1 U11641 ( .A(n15960), .ZN(n15946) );
  OR2_X1 U11642 ( .A1(n11185), .A2(n11184), .ZN(n11795) );
  NAND2_X1 U11643 ( .A1(n11268), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10092) );
  INV_X1 U11644 ( .A(n10166), .ZN(n11912) );
  INV_X1 U11645 ( .A(n11795), .ZN(n11787) );
  AND2_X1 U11646 ( .A1(n10207), .A2(n10209), .ZN(n10204) );
  INV_X1 U11647 ( .A(n15336), .ZN(n10209) );
  AND2_X1 U11648 ( .A1(n10203), .A2(n10020), .ZN(n10019) );
  AND2_X1 U11649 ( .A1(n15161), .A2(n10207), .ZN(n10203) );
  OR2_X1 U11650 ( .A1(n10021), .A2(n12528), .ZN(n10020) );
  INV_X1 U11651 ( .A(n12543), .ZN(n10021) );
  NAND2_X1 U11652 ( .A1(n13047), .A2(n9953), .ZN(n12278) );
  AND2_X1 U11653 ( .A1(n10409), .A2(n10431), .ZN(n10361) );
  NAND2_X1 U11654 ( .A1(n10401), .A2(n19292), .ZN(n10418) );
  NAND3_X1 U11655 ( .A1(n12687), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12683) );
  NAND2_X1 U11656 ( .A1(n18272), .A2(n16551), .ZN(n12927) );
  AND4_X1 U11657 ( .A1(n10936), .A2(n10935), .A3(n10934), .A4(n10933), .ZN(
        n10937) );
  AOI21_X1 U11658 ( .B1(n11731), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A(n9905), .ZN(n11541) );
  AND2_X1 U11659 ( .A1(n9885), .A2(n14434), .ZN(n10179) );
  NOR2_X1 U11660 ( .A1(n9898), .A2(n10174), .ZN(n10173) );
  INV_X1 U11661 ( .A(n14277), .ZN(n10174) );
  INV_X1 U11662 ( .A(n11265), .ZN(n11750) );
  INV_X1 U11663 ( .A(n11286), .ZN(n10175) );
  INV_X1 U11664 ( .A(n13902), .ZN(n11294) );
  AND2_X1 U11665 ( .A1(n11041), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11288) );
  NOR2_X1 U11666 ( .A1(n10107), .A2(n9864), .ZN(n10111) );
  INV_X1 U11667 ( .A(n14154), .ZN(n10143) );
  NOR2_X1 U11668 ( .A1(n10102), .A2(n10098), .ZN(n10097) );
  INV_X1 U11669 ( .A(n13941), .ZN(n10098) );
  INV_X1 U11670 ( .A(n15948), .ZN(n10102) );
  INV_X1 U11671 ( .A(n15947), .ZN(n10100) );
  NAND2_X1 U11672 ( .A1(n11043), .A2(n11031), .ZN(n10166) );
  OR2_X1 U11673 ( .A1(n11121), .A2(n11120), .ZN(n11837) );
  INV_X1 U11674 ( .A(n11837), .ZN(n11833) );
  OR2_X1 U11675 ( .A1(n11151), .A2(n11150), .ZN(n11775) );
  NAND2_X1 U11676 ( .A1(n20202), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11834) );
  INV_X1 U11677 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11865) );
  AND4_X1 U11678 ( .A1(n11013), .A2(n11012), .A3(n11011), .A4(n11010), .ZN(
        n11029) );
  AND3_X1 U11679 ( .A1(n10955), .A2(n10954), .A3(n10953), .ZN(n10956) );
  OAI21_X1 U11680 ( .B1(n20825), .B2(n13761), .A(n14811), .ZN(n20168) );
  NAND2_X1 U11681 ( .A1(n11031), .A2(n11036), .ZN(n11872) );
  OR2_X1 U11682 ( .A1(n11174), .A2(n20169), .ZN(n11903) );
  INV_X1 U11683 ( .A(n12549), .ZN(n10133) );
  OR2_X1 U11684 ( .A1(n12567), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12577) );
  NOR2_X1 U11685 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  INV_X1 U11686 ( .A(n9877), .ZN(n10119) );
  AND2_X1 U11687 ( .A1(n12400), .A2(n10125), .ZN(n12480) );
  NOR2_X1 U11688 ( .A1(n10126), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10125) );
  OR2_X1 U11689 ( .A1(n10129), .A2(n10127), .ZN(n10126) );
  INV_X1 U11690 ( .A(n12468), .ZN(n10127) );
  NOR2_X1 U11691 ( .A1(n12421), .A2(n12401), .ZN(n12400) );
  INV_X1 U11692 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10201) );
  INV_X1 U11693 ( .A(n10223), .ZN(n10222) );
  NAND2_X1 U11694 ( .A1(n9916), .A2(n10224), .ZN(n10223) );
  INV_X1 U11695 ( .A(n14951), .ZN(n10224) );
  INV_X1 U11696 ( .A(n10412), .ZN(n10435) );
  OAI211_X1 U11697 ( .C1(n12413), .C2(n10841), .A(n10660), .B(n10624), .ZN(
        n13286) );
  NOR2_X1 U11698 ( .A1(n10045), .A2(n10044), .ZN(n10043) );
  INV_X1 U11699 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10044) );
  AND4_X1 U11700 ( .A1(n10735), .A2(n10734), .A3(n10733), .A4(n10732), .ZN(
        n10746) );
  AND4_X1 U11701 ( .A1(n10743), .A2(n10742), .A3(n10741), .A4(n10740), .ZN(
        n10744) );
  AND4_X1 U11702 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(
        n10745) );
  NAND2_X1 U11703 ( .A1(n16121), .A2(n12571), .ZN(n12581) );
  INV_X1 U11704 ( .A(n15136), .ZN(n10214) );
  OR2_X1 U11705 ( .A1(n15667), .A2(n12399), .ZN(n12548) );
  NOR2_X1 U11706 ( .A1(n15174), .A2(n15402), .ZN(n9987) );
  OR2_X1 U11707 ( .A1(n18985), .A2(n12504), .ZN(n15173) );
  INV_X1 U11708 ( .A(n14162), .ZN(n10155) );
  AND3_X1 U11709 ( .A1(n10764), .A2(n10763), .A3(n10762), .ZN(n13934) );
  NOR2_X1 U11710 ( .A1(n13425), .A2(n10163), .ZN(n10162) );
  INV_X1 U11711 ( .A(n10164), .ZN(n10163) );
  INV_X1 U11712 ( .A(n12644), .ZN(n12645) );
  INV_X1 U11713 ( .A(n12643), .ZN(n12646) );
  NAND2_X1 U11714 ( .A1(n9949), .A2(n12356), .ZN(n10199) );
  NOR2_X1 U11715 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  OAI22_X1 U11716 ( .A1(n12368), .A2(n12347), .B1(n12346), .B2(n19361), .ZN(
        n12351) );
  NAND2_X1 U11717 ( .A1(n12363), .A2(n10661), .ZN(n12364) );
  INV_X1 U11718 ( .A(n12619), .ZN(n12363) );
  NAND2_X1 U11719 ( .A1(n9853), .A2(n9969), .ZN(n10405) );
  NAND2_X1 U11720 ( .A1(n12307), .A2(n11964), .ZN(n10217) );
  INV_X1 U11721 ( .A(n12378), .ZN(n19461) );
  CLKBUF_X1 U11722 ( .A(n12715), .Z(n17227) );
  AOI21_X1 U11723 ( .B1(n17222), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n10000), .ZN(n9999) );
  AOI21_X1 U11724 ( .B1(n18252), .B2(n12987), .A(n12986), .ZN(n13000) );
  AOI211_X1 U11725 ( .C1(n18257), .C2(n18678), .A(n12998), .B(n12915), .ZN(
        n12926) );
  NAND2_X1 U11726 ( .A1(n12723), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12782) );
  OR2_X1 U11727 ( .A1(n15707), .A2(n13392), .ZN(n13364) );
  NOR2_X1 U11728 ( .A1(n14233), .A2(n9955), .ZN(n9954) );
  INV_X1 U11729 ( .A(n14241), .ZN(n9955) );
  AND4_X1 U11730 ( .A1(n10990), .A2(n10989), .A3(n10988), .A4(n10987), .ZN(
        n11008) );
  INV_X1 U11731 ( .A(n11272), .ZN(n11758) );
  OR2_X1 U11732 ( .A1(n11677), .A2(n14587), .ZN(n11722) );
  AOI21_X1 U11733 ( .B1(n11656), .B2(n11655), .A(n11654), .ZN(n14384) );
  AND2_X1 U11734 ( .A1(n14599), .A2(n13998), .ZN(n11654) );
  OR2_X1 U11735 ( .A1(n11631), .A2(n11630), .ZN(n11675) );
  CLKBUF_X1 U11736 ( .A(n14383), .Z(n14396) );
  NAND2_X1 U11737 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11534), .ZN(
        n11585) );
  NOR2_X1 U11738 ( .A1(n11290), .A2(n13903), .ZN(n11298) );
  INV_X1 U11739 ( .A(n13644), .ZN(n15709) );
  OR2_X1 U11740 ( .A1(n10141), .A2(n13296), .ZN(n10138) );
  NOR2_X1 U11741 ( .A1(n14583), .A2(n10104), .ZN(n14563) );
  NAND2_X1 U11742 ( .A1(n15918), .A2(n10105), .ZN(n10104) );
  NOR2_X1 U11743 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10105) );
  NOR2_X1 U11744 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n14622), .ZN(
        n14600) );
  AND2_X1 U11745 ( .A1(n10145), .A2(n14423), .ZN(n10144) );
  NAND2_X1 U11746 ( .A1(n15793), .A2(n10147), .ZN(n15739) );
  NAND2_X1 U11747 ( .A1(n15793), .A2(n14491), .ZN(n15737) );
  NAND2_X1 U11748 ( .A1(n11037), .A2(n11036), .ZN(n13569) );
  AND2_X1 U11749 ( .A1(n14706), .A2(n14702), .ZN(n14712) );
  NAND2_X1 U11750 ( .A1(n13545), .A2(n13544), .ZN(n13562) );
  INV_X1 U11751 ( .A(n20005), .ZN(n20011) );
  NOR2_X1 U11752 ( .A1(n13788), .A2(n13789), .ZN(n20490) );
  OR2_X1 U11753 ( .A1(n13763), .A2(n20257), .ZN(n20616) );
  NOR2_X1 U11754 ( .A1(n20496), .A2(n20334), .ZN(n20646) );
  INV_X2 U11755 ( .A(n13096), .ZN(n20183) );
  AND2_X1 U11756 ( .A1(n13763), .A2(n20257), .ZN(n20637) );
  NOR2_X1 U11757 ( .A1(n11774), .A2(n13790), .ZN(n20638) );
  INV_X1 U11758 ( .A(n20638), .ZN(n20685) );
  NAND2_X1 U11759 ( .A1(n11869), .A2(n11868), .ZN(n13259) );
  NOR2_X1 U11760 ( .A1(n11903), .A2(n11872), .ZN(n11909) );
  NAND2_X1 U11761 ( .A1(n12570), .A2(n12576), .ZN(n12580) );
  NOR2_X1 U11762 ( .A1(n12580), .A2(n12572), .ZN(n12587) );
  NAND2_X1 U11763 ( .A1(n12594), .A2(n12577), .ZN(n12570) );
  NOR3_X1 U11764 ( .A1(n12550), .A2(n12549), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n12566) );
  NAND2_X1 U11765 ( .A1(n12546), .A2(n12594), .ZN(n12499) );
  NAND2_X1 U11766 ( .A1(n12594), .A2(n12503), .ZN(n12517) );
  NOR2_X1 U11767 ( .A1(n10122), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10121) );
  INV_X1 U11768 ( .A(n10123), .ZN(n10122) );
  OR2_X1 U11769 ( .A1(n12501), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12503) );
  NOR2_X1 U11770 ( .A1(n10227), .A2(n10232), .ZN(n10225) );
  NAND2_X1 U11771 ( .A1(n13581), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10227) );
  AND2_X1 U11772 ( .A1(n15019), .A2(n14832), .ZN(n15005) );
  AND2_X1 U11773 ( .A1(n14122), .A2(n14119), .ZN(n11988) );
  AOI21_X1 U11774 ( .B1(n9827), .B2(n15534), .A(n9901), .ZN(n10076) );
  AND2_X1 U11775 ( .A1(n10265), .A2(n10056), .ZN(n10294) );
  AND2_X1 U11776 ( .A1(n9840), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10056) );
  AND3_X1 U11777 ( .A1(n10539), .A2(n10538), .A3(n10537), .ZN(n14947) );
  AND3_X1 U11778 ( .A1(n10536), .A2(n10535), .A3(n10534), .ZN(n14960) );
  AND2_X1 U11779 ( .A1(n9899), .A2(n14908), .ZN(n10150) );
  INV_X1 U11780 ( .A(n14894), .ZN(n10151) );
  NAND2_X1 U11781 ( .A1(n14910), .A2(n14829), .ZN(n14895) );
  AND2_X1 U11782 ( .A1(n14920), .A2(n14908), .ZN(n14910) );
  NAND2_X1 U11783 ( .A1(n15099), .A2(n15098), .ZN(n15123) );
  NAND2_X1 U11784 ( .A1(n10192), .A2(n10190), .ZN(n15140) );
  NOR2_X1 U11785 ( .A1(n10191), .A2(n15152), .ZN(n10190) );
  INV_X1 U11786 ( .A(n10193), .ZN(n10191) );
  OR2_X1 U11787 ( .A1(n12548), .A2(n15348), .ZN(n15336) );
  NAND2_X1 U11788 ( .A1(n15226), .A2(n12528), .ZN(n10018) );
  INV_X1 U11789 ( .A(n9976), .ZN(n9975) );
  OAI21_X1 U11790 ( .B1(n15179), .B2(n9979), .A(n9977), .ZN(n9976) );
  NAND2_X1 U11791 ( .A1(n9983), .A2(n15195), .ZN(n9977) );
  NAND2_X1 U11792 ( .A1(n14965), .A2(n14966), .ZN(n14957) );
  AND2_X1 U11793 ( .A1(n10843), .A2(n10842), .ZN(n14124) );
  OAI211_X1 U11794 ( .C1(n15167), .C2(n15169), .A(n15168), .B(n15398), .ZN(
        n15170) );
  NAND2_X1 U11795 ( .A1(n14873), .A2(n15405), .ZN(n15406) );
  AND2_X1 U11796 ( .A1(n14076), .A2(n9883), .ZN(n14993) );
  NAND2_X1 U11797 ( .A1(n14076), .A2(n14077), .ZN(n14075) );
  AND3_X1 U11798 ( .A1(n10789), .A2(n10788), .A3(n10787), .ZN(n15477) );
  NAND2_X1 U11799 ( .A1(n15242), .A2(n15243), .ZN(n12462) );
  NAND2_X1 U11800 ( .A1(n15564), .A2(n11964), .ZN(n11937) );
  CLKBUF_X1 U11801 ( .A(n13413), .Z(n13414) );
  AND2_X1 U11802 ( .A1(n13416), .A2(n13497), .ZN(n13418) );
  NAND2_X1 U11803 ( .A1(n19521), .A2(n19520), .ZN(n19491) );
  OR2_X1 U11804 ( .A1(n19521), .A2(n19520), .ZN(n19744) );
  OR2_X1 U11805 ( .A1(n19961), .A2(n19974), .ZN(n19709) );
  AOI21_X1 U11806 ( .B1(n17229), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n12732), .ZN(n12733) );
  AND2_X1 U11807 ( .A1(n9835), .A2(n10036), .ZN(n10035) );
  INV_X1 U11808 ( .A(n16380), .ZN(n10036) );
  INV_X1 U11809 ( .A(n18090), .ZN(n17732) );
  NOR2_X1 U11810 ( .A1(n16532), .A2(n18885), .ZN(n16385) );
  AND2_X1 U11811 ( .A1(n12824), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10014) );
  OR2_X1 U11812 ( .A1(n17692), .A2(n17590), .ZN(n12818) );
  INV_X1 U11813 ( .A(n17636), .ZN(n10012) );
  NAND2_X1 U11814 ( .A1(n18690), .A2(n17286), .ZN(n12992) );
  OAI21_X1 U11815 ( .B1(n17876), .B2(n10009), .A(n10006), .ZN(n17861) );
  INV_X1 U11816 ( .A(n12794), .ZN(n10009) );
  AND2_X1 U11817 ( .A1(n10007), .A2(n17863), .ZN(n10006) );
  NAND2_X1 U11818 ( .A1(n17876), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17875) );
  NAND2_X1 U11819 ( .A1(n17903), .A2(n17895), .ZN(n17894) );
  NAND2_X1 U11820 ( .A1(n12949), .A2(n12926), .ZN(n18662) );
  NOR2_X1 U11821 ( .A1(n18697), .A2(n16933), .ZN(n18672) );
  AOI21_X1 U11822 ( .B1(n15646), .B2(n17435), .A(n15645), .ZN(n18703) );
  NAND2_X1 U11823 ( .A1(n14492), .A2(n20221), .ZN(n15876) );
  AND2_X1 U11824 ( .A1(n14551), .A2(n13575), .ZN(n15888) );
  NAND2_X1 U11825 ( .A1(n15955), .A2(n11916), .ZN(n15960) );
  OR2_X2 U11826 ( .A1(n15714), .A2(n20005), .ZN(n15955) );
  CLKBUF_X1 U11827 ( .A(n13381), .Z(n13382) );
  NAND2_X1 U11828 ( .A1(n15707), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14811) );
  INV_X1 U11829 ( .A(n20439), .ZN(n20460) );
  AND2_X1 U11830 ( .A1(n12487), .A2(n10116), .ZN(n12508) );
  AND2_X1 U11831 ( .A1(n12301), .A2(n12592), .ZN(n16165) );
  NAND2_X1 U11832 ( .A1(n13212), .A2(n12671), .ZN(n16275) );
  AND2_X1 U11833 ( .A1(n12670), .A2(n16362), .ZN(n19248) );
  NAND2_X1 U11834 ( .A1(n13086), .A2(n13080), .ZN(n10073) );
  NAND2_X1 U11835 ( .A1(n15089), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9947) );
  NOR2_X1 U11836 ( .A1(n16092), .A2(n16313), .ZN(n10074) );
  XNOR2_X1 U11837 ( .A(n13075), .B(n13074), .ZN(n19119) );
  NAND2_X1 U11838 ( .A1(n15192), .A2(n9978), .ZN(n9972) );
  AND2_X1 U11839 ( .A1(n15179), .A2(n9983), .ZN(n9978) );
  NAND2_X1 U11840 ( .A1(n15194), .A2(n9974), .ZN(n9973) );
  INV_X1 U11841 ( .A(n9979), .ZN(n9974) );
  AND2_X1 U11842 ( .A1(n13089), .A2(n13079), .ZN(n16307) );
  INV_X1 U11843 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19987) );
  AND2_X1 U11844 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11965), .ZN(
        n19530) );
  INV_X1 U11845 ( .A(n16573), .ZN(n10042) );
  AND2_X1 U11846 ( .A1(n16574), .A2(n10041), .ZN(n10040) );
  OR2_X1 U11847 ( .A1(n16918), .A2(n16575), .ZN(n10041) );
  NAND2_X1 U11848 ( .A1(n16408), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10027) );
  INV_X1 U11849 ( .A(n16902), .ZN(n16918) );
  NOR2_X2 U11850 ( .A1(n18832), .A2(n16901), .ZN(n16902) );
  INV_X1 U11851 ( .A(n12885), .ZN(n12895) );
  AND2_X1 U11852 ( .A1(n17362), .A2(n10062), .ZN(n17320) );
  INV_X1 U11853 ( .A(n17350), .ZN(n17357) );
  INV_X1 U11854 ( .A(n17331), .ZN(n17356) );
  NAND2_X1 U11855 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17367), .ZN(n17363) );
  NOR2_X1 U11856 ( .A1(n17363), .A2(n17539), .ZN(n17362) );
  NOR2_X1 U11857 ( .A1(n17398), .A2(n17369), .ZN(n17367) );
  AOI211_X1 U11858 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n12696), .B(n12695), .ZN(n17404) );
  INV_X1 U11859 ( .A(n17428), .ZN(n17422) );
  INV_X1 U11860 ( .A(n12964), .ZN(n17434) );
  AND2_X1 U11861 ( .A1(n17279), .A2(n18272), .ZN(n17428) );
  NAND2_X1 U11862 ( .A1(n15763), .A2(n17279), .ZN(n17433) );
  AND2_X1 U11863 ( .A1(n10068), .A2(n18878), .ZN(n17279) );
  INV_X1 U11864 ( .A(n17421), .ZN(n17431) );
  NOR2_X1 U11865 ( .A1(n17907), .A2(n16386), .ZN(n17816) );
  INV_X1 U11866 ( .A(n17790), .ZN(n17815) );
  AOI21_X1 U11867 ( .B1(n12830), .B2(n12829), .A(n10011), .ZN(n16388) );
  AOI21_X1 U11868 ( .B1(n9824), .B2(n10095), .A(n10094), .ZN(n10011) );
  NAND2_X1 U11869 ( .A1(n16386), .A2(n18220), .ZN(n18113) );
  INV_X1 U11870 ( .A(n18113), .ZN(n18139) );
  OAI221_X2 U11871 ( .B1(n12950), .B2(n18663), .C1(n12950), .C2(n12949), .A(
        n18878), .ZN(n18222) );
  AOI21_X1 U11872 ( .B1(n11739), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n9908), .ZN(n11688) );
  AOI21_X1 U11873 ( .B1(n11739), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n9907), .ZN(n11643) );
  CLKBUF_X1 U11874 ( .A(n11051), .Z(n11052) );
  AND2_X2 U11875 ( .A1(n10911), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10918) );
  AND2_X1 U11876 ( .A1(n19987), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10582) );
  NAND2_X1 U11877 ( .A1(n10208), .A2(n15336), .ZN(n10207) );
  INV_X1 U11878 ( .A(n15335), .ZN(n10208) );
  NAND2_X1 U11879 ( .A1(n10572), .A2(n10571), .ZN(n10578) );
  OAI21_X1 U11880 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n12687), .A(
        n12916), .ZN(n12924) );
  OR2_X1 U11881 ( .A1(n12937), .A2(n12938), .ZN(n12916) );
  AOI21_X1 U11882 ( .B1(n11707), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A(n9910), .ZN(n11615) );
  AOI21_X1 U11883 ( .B1(n11739), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n9906), .ZN(n11599) );
  NAND2_X1 U11884 ( .A1(n11296), .A2(n11286), .ZN(n10176) );
  INV_X1 U11885 ( .A(n11844), .ZN(n10108) );
  OR2_X1 U11886 ( .A1(n11225), .A2(n11224), .ZN(n11820) );
  OR2_X1 U11887 ( .A1(n11213), .A2(n11212), .ZN(n11808) );
  OR2_X1 U11888 ( .A1(n11200), .A2(n11199), .ZN(n11797) );
  NAND2_X1 U11889 ( .A1(n11762), .A2(n11049), .ZN(n11068) );
  NAND2_X1 U11890 ( .A1(n11127), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11022) );
  INV_X1 U11891 ( .A(n11907), .ZN(n11895) );
  OR2_X1 U11892 ( .A1(n11879), .A2(n15708), .ZN(n11897) );
  AND4_X1 U11893 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10747) );
  NAND2_X1 U11894 ( .A1(n12429), .A2(n9856), .ZN(n12643) );
  AND2_X1 U11895 ( .A1(n10188), .A2(n14172), .ZN(n10187) );
  NAND2_X1 U11896 ( .A1(n10334), .A2(n10333), .ZN(n9969) );
  NAND2_X1 U11897 ( .A1(n11930), .A2(n10401), .ZN(n9968) );
  AND3_X2 U11898 ( .A1(n15574), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12053) );
  NAND2_X1 U11899 ( .A1(n10411), .A2(n10410), .ZN(n13024) );
  OAI21_X1 U11900 ( .B1(n12780), .B2(n17232), .A(n10001), .ZN(n10000) );
  NAND2_X1 U11901 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10001) );
  INV_X1 U11902 ( .A(n10113), .ZN(n17706) );
  INV_X1 U11903 ( .A(n17423), .ZN(n12961) );
  NAND2_X1 U11904 ( .A1(n12979), .A2(n12978), .ZN(n12984) );
  INV_X1 U11905 ( .A(n12932), .ZN(n12928) );
  AND2_X1 U11906 ( .A1(n12989), .A2(n13798), .ZN(n12978) );
  NAND2_X1 U11907 ( .A1(n12995), .A2(n12979), .ZN(n12929) );
  NAND2_X1 U11908 ( .A1(n10258), .A2(n10184), .ZN(n10183) );
  INV_X1 U11909 ( .A(n14371), .ZN(n10184) );
  AND2_X1 U11910 ( .A1(n11586), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11587) );
  INV_X1 U11911 ( .A(n11585), .ZN(n11586) );
  AOI21_X1 U11912 ( .B1(n11657), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n9909), .ZN(n11521) );
  OR2_X1 U11913 ( .A1(n13175), .A2(n10140), .ZN(n10139) );
  INV_X1 U11914 ( .A(n14360), .ZN(n10140) );
  NAND2_X1 U11915 ( .A1(n14629), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14601) );
  AND2_X1 U11916 ( .A1(n10147), .A2(n10146), .ZN(n10145) );
  INV_X1 U11917 ( .A(n14435), .ZN(n10146) );
  NOR2_X1 U11918 ( .A1(n10148), .A2(n15736), .ZN(n10147) );
  INV_X1 U11919 ( .A(n14491), .ZN(n10148) );
  NAND2_X1 U11920 ( .A1(n14217), .A2(n10109), .ZN(n10110) );
  INV_X1 U11921 ( .A(n14214), .ZN(n10142) );
  OAI21_X1 U11922 ( .B1(n13788), .B2(n11872), .A(n11789), .ZN(n11791) );
  OR2_X1 U11923 ( .A1(n11133), .A2(n11132), .ZN(n11776) );
  AND2_X1 U11924 ( .A1(n11154), .A2(n11153), .ZN(n11163) );
  OAI21_X1 U11925 ( .B1(n11269), .B2(n10093), .A(n9863), .ZN(n11139) );
  INV_X1 U11926 ( .A(n11268), .ZN(n10093) );
  AOI21_X1 U11927 ( .B1(n11080), .B2(n13751), .A(n11081), .ZN(n11089) );
  NAND2_X1 U11928 ( .A1(n11912), .A2(n9965), .ZN(n13558) );
  INV_X1 U11929 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20259) );
  AOI21_X1 U11930 ( .B1(n11874), .B2(n11873), .A(n11866), .ZN(n11871) );
  NOR2_X1 U11931 ( .A1(n10124), .A2(n10891), .ZN(n10123) );
  NAND2_X1 U11932 ( .A1(n12480), .A2(n12479), .ZN(n12484) );
  NAND2_X1 U11933 ( .A1(n12457), .A2(n12463), .ZN(n10129) );
  NAND2_X1 U11934 ( .A1(n10883), .A2(n10882), .ZN(n12407) );
  NAND2_X1 U11935 ( .A1(n12592), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U11936 ( .A1(n12604), .A2(n19277), .ZN(n10883) );
  OR2_X1 U11937 ( .A1(n12138), .A2(n12139), .ZN(n12140) );
  INV_X1 U11938 ( .A(n14846), .ZN(n10088) );
  NOR2_X1 U11939 ( .A1(n10090), .A2(n15044), .ZN(n10089) );
  INV_X1 U11940 ( .A(n15339), .ZN(n10090) );
  INV_X1 U11941 ( .A(n14982), .ZN(n10235) );
  OR2_X1 U11942 ( .A1(n10725), .A2(n10724), .ZN(n12453) );
  NOR2_X1 U11943 ( .A1(n10712), .A2(n10711), .ZN(n12396) );
  NOR2_X1 U11944 ( .A1(n15117), .A2(n10058), .ZN(n10057) );
  NOR2_X1 U11945 ( .A1(n10160), .A2(n14960), .ZN(n10159) );
  INV_X1 U11946 ( .A(n14966), .ZN(n10160) );
  NOR2_X1 U11947 ( .A1(n15220), .A2(n10048), .ZN(n10047) );
  NOR2_X1 U11948 ( .A1(n16230), .A2(n10051), .ZN(n10050) );
  INV_X1 U11949 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U11950 ( .A1(n16266), .A2(n10052), .ZN(n10055) );
  OR2_X1 U11951 ( .A1(n10622), .A2(n10621), .ZN(n12624) );
  NAND2_X1 U11952 ( .A1(n10196), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10195) );
  NOR2_X1 U11953 ( .A1(n15109), .A2(n15122), .ZN(n10196) );
  INV_X1 U11954 ( .A(n15100), .ZN(n10213) );
  NAND2_X1 U11955 ( .A1(n10017), .A2(n10016), .ZN(n12558) );
  AOI21_X1 U11956 ( .B1(n10019), .B2(n10021), .A(n9867), .ZN(n10016) );
  NOR2_X1 U11957 ( .A1(n15348), .A2(n10194), .ZN(n10193) );
  INV_X1 U11958 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10194) );
  INV_X1 U11959 ( .A(n15063), .ZN(n10081) );
  OR2_X1 U11960 ( .A1(n12539), .A2(n12538), .ZN(n15176) );
  AND2_X1 U11961 ( .A1(n9883), .A2(n14994), .ZN(n10154) );
  NAND2_X1 U11962 ( .A1(n13961), .A2(n13960), .ZN(n13933) );
  AND2_X1 U11963 ( .A1(n13610), .A2(n13620), .ZN(n10164) );
  OR2_X1 U11964 ( .A1(n10642), .A2(n10641), .ZN(n12622) );
  NAND2_X1 U11965 ( .A1(n10409), .A2(n14108), .ZN(n10026) );
  INV_X1 U11966 ( .A(n15602), .ZN(n12235) );
  INV_X1 U11967 ( .A(n10417), .ZN(n10429) );
  INV_X1 U11968 ( .A(n12982), .ZN(n16549) );
  NOR2_X1 U11969 ( .A1(n10240), .A2(n12731), .ZN(n12732) );
  NOR2_X1 U11970 ( .A1(n17850), .A2(n10034), .ZN(n10033) );
  INV_X1 U11971 ( .A(n17849), .ZN(n10032) );
  OR2_X1 U11972 ( .A1(n16531), .A2(n12995), .ZN(n12982) );
  OR2_X1 U11973 ( .A1(n17415), .A2(n12956), .ZN(n12954) );
  INV_X1 U11974 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10008) );
  XNOR2_X1 U11975 ( .A(n17423), .B(n12964), .ZN(n12789) );
  OAI21_X1 U11976 ( .B1(n12941), .B2(n12940), .A(n12939), .ZN(n16529) );
  CLKBUF_X1 U11977 ( .A(n13262), .Z(n15704) );
  NOR2_X1 U11978 ( .A1(n11450), .A2(n14451), .ZN(n11465) );
  NOR2_X1 U11979 ( .A1(n14399), .A2(n13175), .ZN(n14376) );
  AND2_X1 U11980 ( .A1(n13152), .A2(n13151), .ZN(n14498) );
  AOI21_X1 U11981 ( .B1(n13998), .B2(n14555), .A(n11756), .ZN(n13184) );
  OR2_X1 U11982 ( .A1(n11724), .A2(n14352), .ZN(n11920) );
  NAND2_X1 U11983 ( .A1(n11629), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11631) );
  INV_X1 U11984 ( .A(n11628), .ZN(n11629) );
  AND2_X1 U11985 ( .A1(n11634), .A2(n11633), .ZN(n14394) );
  OR2_X1 U11986 ( .A1(n14607), .A2(n11750), .ZN(n11633) );
  NAND2_X1 U11987 ( .A1(n11587), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11628) );
  CLKBUF_X1 U11988 ( .A(n14409), .Z(n14410) );
  AND2_X1 U11989 ( .A1(n14637), .A2(n13998), .ZN(n11555) );
  NOR2_X1 U11990 ( .A1(n11497), .A2(n15800), .ZN(n11498) );
  NAND2_X1 U11991 ( .A1(n11465), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11497) );
  CLKBUF_X1 U11992 ( .A(n14494), .Z(n14495) );
  NOR2_X1 U11993 ( .A1(n10172), .A2(n15809), .ZN(n10171) );
  INV_X1 U11994 ( .A(n10173), .ZN(n10172) );
  OR2_X1 U11995 ( .A1(n11432), .A2(n15825), .ZN(n11450) );
  INV_X1 U11996 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14451) );
  INV_X1 U11997 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15825) );
  AND2_X1 U11998 ( .A1(n11398), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11415) );
  NAND2_X1 U11999 ( .A1(n11368), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11383) );
  NAND2_X1 U12000 ( .A1(n11367), .A2(n11366), .ZN(n14234) );
  INV_X1 U12001 ( .A(n14131), .ZN(n11367) );
  NOR2_X1 U12002 ( .A1(n11349), .A2(n11348), .ZN(n11368) );
  CLKBUF_X1 U12003 ( .A(n14208), .Z(n14209) );
  NAND2_X1 U12004 ( .A1(n11334), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11349) );
  INV_X1 U12005 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11348) );
  NOR2_X1 U12006 ( .A1(n11317), .A2(n11316), .ZN(n11334) );
  NOR2_X1 U12007 ( .A1(n11306), .A2(n15961), .ZN(n11307) );
  CLKBUF_X1 U12008 ( .A(n13954), .Z(n13955) );
  AOI21_X1 U12009 ( .B1(n11805), .B2(n11395), .A(n11301), .ZN(n13916) );
  NOR2_X1 U12010 ( .A1(n13899), .A2(n13916), .ZN(n13915) );
  AOI21_X1 U12011 ( .B1(n11794), .B2(n11395), .A(n11293), .ZN(n13902) );
  CLKBUF_X1 U12012 ( .A(n13899), .Z(n13900) );
  NAND3_X1 U12013 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11290) );
  AOI21_X1 U12014 ( .B1(n11257), .B2(n11447), .A(n10169), .ZN(n10168) );
  INV_X1 U12015 ( .A(n13657), .ZN(n10169) );
  OR2_X1 U12016 ( .A1(n14399), .A2(n10139), .ZN(n14362) );
  AND2_X1 U12017 ( .A1(n14591), .A2(n14594), .ZN(n10106) );
  NAND2_X1 U12018 ( .A1(n14425), .A2(n14412), .ZN(n14414) );
  NAND2_X1 U12019 ( .A1(n11854), .A2(n15918), .ZN(n14630) );
  NOR2_X1 U12020 ( .A1(n14639), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15734) );
  AND2_X1 U12021 ( .A1(n14497), .A2(n13155), .ZN(n15793) );
  OR2_X1 U12022 ( .A1(n15812), .A2(n15811), .ZN(n15814) );
  OR2_X1 U12023 ( .A1(n14793), .A2(n14251), .ZN(n15823) );
  NOR2_X1 U12024 ( .A1(n15823), .A2(n15824), .ZN(n15822) );
  OR2_X1 U12025 ( .A1(n15908), .A2(n16025), .ZN(n15931) );
  OR2_X1 U12026 ( .A1(n15908), .A2(n11849), .ZN(n15927) );
  OR2_X1 U12027 ( .A1(n14791), .A2(n14790), .ZN(n14793) );
  OR2_X1 U12028 ( .A1(n11856), .A2(n11850), .ZN(n14668) );
  OAI21_X1 U12029 ( .B1(n13598), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13676), .ZN(n14760) );
  NAND2_X1 U12030 ( .A1(n14145), .A2(n9881), .ZN(n14213) );
  OR2_X1 U12031 ( .A1(n14217), .A2(n11844), .ZN(n15938) );
  AND2_X1 U12032 ( .A1(n13130), .A2(n13129), .ZN(n14144) );
  AND2_X1 U12033 ( .A1(n16066), .A2(n14045), .ZN(n14145) );
  NAND2_X1 U12034 ( .A1(n14145), .A2(n14144), .ZN(n14155) );
  AOI21_X1 U12035 ( .B1(n15948), .B2(n10101), .A(n10100), .ZN(n10099) );
  INV_X1 U12036 ( .A(n11826), .ZN(n10101) );
  NOR2_X1 U12037 ( .A1(n16064), .A2(n16063), .ZN(n16066) );
  AND2_X1 U12038 ( .A1(n13122), .A2(n13121), .ZN(n13944) );
  NAND2_X1 U12039 ( .A1(n10136), .A2(n10135), .ZN(n16064) );
  INV_X1 U12040 ( .A(n13944), .ZN(n10135) );
  INV_X1 U12041 ( .A(n13945), .ZN(n10136) );
  OR2_X1 U12042 ( .A1(n13895), .A2(n13894), .ZN(n13945) );
  NAND2_X1 U12043 ( .A1(n13772), .A2(n13771), .ZN(n13895) );
  OR2_X1 U12044 ( .A1(n13596), .A2(n13595), .ZN(n13679) );
  NOR2_X1 U12045 ( .A1(n13679), .A2(n13678), .ZN(n13772) );
  OAI21_X1 U12046 ( .B1(n14802), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11160), 
        .ZN(n11161) );
  CLKBUF_X1 U12047 ( .A(n13253), .Z(n13254) );
  OR2_X1 U12048 ( .A1(n11049), .A2(n11050), .ZN(n14806) );
  INV_X1 U12049 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14810) );
  OR3_X1 U12050 ( .A1(n13380), .A2(n13571), .A3(n13379), .ZN(n15680) );
  NAND2_X1 U12051 ( .A1(n13788), .A2(n11774), .ZN(n20300) );
  INV_X1 U12052 ( .A(n20409), .ZN(n20414) );
  NAND2_X1 U12053 ( .A1(n13763), .A2(n20159), .ZN(n20545) );
  NAND2_X1 U12054 ( .A1(n20166), .A2(n20164), .ZN(n20225) );
  INV_X1 U12055 ( .A(n20298), .ZN(n20684) );
  INV_X1 U12056 ( .A(n20540), .ZN(n20688) );
  AOI21_X1 U12057 ( .B1(n20610), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20334), 
        .ZN(n20687) );
  NAND3_X1 U12058 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20169), .A3(n20168), 
        .ZN(n20222) );
  AND2_X1 U12059 ( .A1(n13025), .A2(n12282), .ZN(n16341) );
  NOR2_X1 U12060 ( .A1(n12545), .A2(n10132), .ZN(n10131) );
  NAND2_X1 U12061 ( .A1(n10133), .A2(n9844), .ZN(n10132) );
  OR2_X1 U12062 ( .A1(n12550), .A2(n12549), .ZN(n12555) );
  NAND2_X1 U12063 ( .A1(n12517), .A2(n10123), .ZN(n12526) );
  NAND2_X1 U12064 ( .A1(n10280), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10279) );
  NOR2_X1 U12065 ( .A1(n10117), .A2(n12509), .ZN(n10116) );
  INV_X1 U12066 ( .A(n10118), .ZN(n10117) );
  NAND2_X1 U12067 ( .A1(n12487), .A2(n10118), .ZN(n12511) );
  NAND2_X1 U12068 ( .A1(n13923), .A2(n13924), .ZN(n14053) );
  NAND2_X1 U12069 ( .A1(n12487), .A2(n12494), .ZN(n12514) );
  AND2_X1 U12070 ( .A1(n12473), .A2(n12472), .ZN(n19050) );
  NOR2_X1 U12071 ( .A1(n10126), .A2(n10130), .ZN(n12470) );
  NOR2_X1 U12072 ( .A1(n10130), .A2(n10128), .ZN(n12465) );
  OR2_X1 U12073 ( .A1(n16338), .A2(n13230), .ZN(n13205) );
  AND3_X1 U12074 ( .A1(n10527), .A2(n10526), .A3(n10525), .ZN(n14860) );
  NAND2_X1 U12075 ( .A1(n15338), .A2(n10089), .ZN(n15046) );
  OAI211_X1 U12076 ( .C1(n14956), .C2(n10221), .A(n10219), .B(n10218), .ZN(
        n14941) );
  NAND2_X1 U12077 ( .A1(n10220), .A2(n10223), .ZN(n10219) );
  NAND2_X1 U12078 ( .A1(n12108), .A2(n10222), .ZN(n10221) );
  NAND2_X1 U12079 ( .A1(n15338), .A2(n15339), .ZN(n15341) );
  INV_X1 U12080 ( .A(n15418), .ZN(n10085) );
  AND3_X1 U12081 ( .A1(n10828), .A2(n10827), .A3(n10826), .ZN(n14875) );
  OR2_X1 U12082 ( .A1(n13978), .A2(n9827), .ZN(n14184) );
  NOR2_X1 U12083 ( .A1(n13205), .A2(n10898), .ZN(n13445) );
  INV_X1 U12084 ( .A(n12298), .ZN(n14107) );
  NAND2_X1 U12085 ( .A1(n10265), .A2(n9840), .ZN(n10292) );
  NAND2_X1 U12086 ( .A1(n10265), .A2(n10057), .ZN(n10290) );
  NAND2_X1 U12087 ( .A1(n10265), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10288) );
  NAND2_X1 U12088 ( .A1(n10283), .A2(n9838), .ZN(n10285) );
  NOR2_X1 U12089 ( .A1(n10282), .A2(n18932), .ZN(n10283) );
  NAND2_X1 U12090 ( .A1(n10283), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10284) );
  NAND2_X1 U12091 ( .A1(n14965), .A2(n10159), .ZN(n14958) );
  NAND2_X1 U12092 ( .A1(n10266), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10282) );
  AND2_X1 U12093 ( .A1(n10280), .A2(n10046), .ZN(n10266) );
  AND2_X1 U12094 ( .A1(n9836), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10046) );
  NAND2_X1 U12095 ( .A1(n10280), .A2(n9836), .ZN(n10281) );
  AND2_X1 U12096 ( .A1(n15375), .A2(n16299), .ZN(n10197) );
  NAND2_X1 U12097 ( .A1(n14076), .A2(n10152), .ZN(n14987) );
  AND2_X1 U12098 ( .A1(n10154), .A2(n10153), .ZN(n10152) );
  INV_X1 U12099 ( .A(n14989), .ZN(n10153) );
  NOR2_X1 U12100 ( .A1(n10277), .A2(n18999), .ZN(n10280) );
  AND2_X1 U12101 ( .A1(n10275), .A2(n10049), .ZN(n10278) );
  AND2_X1 U12102 ( .A1(n9826), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10049) );
  NAND2_X1 U12103 ( .A1(n10278), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10277) );
  NAND2_X1 U12104 ( .A1(n10275), .A2(n9826), .ZN(n10276) );
  NAND2_X1 U12105 ( .A1(n10275), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10274) );
  NOR2_X1 U12106 ( .A1(n16241), .A2(n10272), .ZN(n10275) );
  NAND2_X1 U12107 ( .A1(n10054), .A2(n10053), .ZN(n10272) );
  AND2_X1 U12108 ( .A1(n9828), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10053) );
  NAND2_X1 U12109 ( .A1(n10054), .A2(n10055), .ZN(n10270) );
  AND2_X1 U12110 ( .A1(n10054), .A2(n9828), .ZN(n10273) );
  NOR2_X1 U12111 ( .A1(n10268), .A2(n16266), .ZN(n10271) );
  INV_X1 U12112 ( .A(n12639), .ZN(n9952) );
  NAND2_X1 U12113 ( .A1(n12637), .A2(n14038), .ZN(n14170) );
  NAND2_X1 U12114 ( .A1(n12638), .A2(n14179), .ZN(n14169) );
  NAND2_X1 U12115 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10267) );
  NOR2_X1 U12116 ( .A1(n10267), .A2(n16276), .ZN(n10269) );
  NAND2_X1 U12117 ( .A1(n11957), .A2(n11955), .ZN(n11959) );
  AND2_X1 U12118 ( .A1(n10587), .A2(n19979), .ZN(n10588) );
  NOR2_X1 U12119 ( .A1(n10253), .A2(n12590), .ZN(n12591) );
  NAND2_X1 U12120 ( .A1(n13075), .A2(n10871), .ZN(n14309) );
  AND2_X1 U12121 ( .A1(n10214), .A2(n15128), .ZN(n10022) );
  OR2_X1 U12122 ( .A1(n16109), .A2(n12399), .ZN(n15100) );
  XNOR2_X1 U12123 ( .A(n12581), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15128) );
  NAND2_X1 U12124 ( .A1(n12562), .A2(n10024), .ZN(n15135) );
  NOR3_X1 U12125 ( .A1(n12582), .A2(n12399), .A3(n15303), .ZN(n15138) );
  AND2_X1 U12126 ( .A1(n10024), .A2(n10214), .ZN(n10023) );
  AND2_X1 U12127 ( .A1(n14965), .A2(n9887), .ZN(n14944) );
  INV_X1 U12128 ( .A(n14943), .ZN(n10156) );
  NAND2_X1 U12129 ( .A1(n14965), .A2(n10157), .ZN(n14949) );
  NAND2_X1 U12130 ( .A1(n10192), .A2(n10193), .ZN(n15151) );
  NAND2_X1 U12131 ( .A1(n15182), .A2(n15178), .ZN(n9979) );
  AND2_X1 U12132 ( .A1(n14977), .A2(n14976), .ZN(n14965) );
  NAND2_X1 U12133 ( .A1(n10083), .A2(n14202), .ZN(n10082) );
  INV_X1 U12134 ( .A(n14124), .ZN(n10083) );
  AOI21_X1 U12135 ( .B1(n9987), .B2(n15172), .A(n9985), .ZN(n9984) );
  INV_X1 U12136 ( .A(n9987), .ZN(n9986) );
  INV_X1 U12137 ( .A(n15173), .ZN(n9985) );
  NAND2_X1 U12138 ( .A1(n14076), .A2(n10154), .ZN(n14996) );
  NOR2_X1 U12139 ( .A1(n15491), .A2(n9880), .ZN(n15417) );
  NOR2_X1 U12140 ( .A1(n13911), .A2(n13912), .ZN(n13923) );
  NAND2_X1 U12141 ( .A1(n13780), .A2(n13781), .ZN(n13911) );
  OR2_X1 U12142 ( .A1(n12656), .A2(n12658), .ZN(n12659) );
  NAND2_X1 U12143 ( .A1(n13504), .A2(n10161), .ZN(n13686) );
  AND2_X1 U12144 ( .A1(n10162), .A2(n13577), .ZN(n10161) );
  NOR2_X1 U12145 ( .A1(n13686), .A2(n13687), .ZN(n13780) );
  AND3_X1 U12146 ( .A1(n10494), .A2(n10493), .A3(n10492), .ZN(n13425) );
  AND2_X1 U12147 ( .A1(n13504), .A2(n10162), .ZN(n13576) );
  NAND2_X1 U12148 ( .A1(n13504), .A2(n10164), .ZN(n13609) );
  AND2_X1 U12149 ( .A1(n13299), .A2(n16290), .ZN(n13069) );
  NOR2_X1 U12150 ( .A1(n13082), .A2(n14177), .ZN(n15539) );
  CLKBUF_X1 U12151 ( .A(n15240), .Z(n15241) );
  AND2_X1 U12152 ( .A1(n13504), .A2(n13620), .ZN(n13622) );
  AND3_X1 U12153 ( .A1(n10702), .A2(n10701), .A3(n10700), .ZN(n14031) );
  AND2_X1 U12154 ( .A1(n12364), .A2(n12344), .ZN(n10198) );
  XNOR2_X1 U12155 ( .A(n10646), .B(n10628), .ZN(n13275) );
  INV_X1 U12156 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15562) );
  INV_X1 U12157 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15574) );
  NOR2_X1 U12158 ( .A1(n13207), .A2(n10210), .ZN(n13042) );
  INV_X1 U12159 ( .A(n11929), .ZN(n10216) );
  NAND2_X1 U12160 ( .A1(n13021), .A2(n12274), .ZN(n16340) );
  NAND2_X1 U12161 ( .A1(n13417), .A2(n13418), .ZN(n13499) );
  AND2_X1 U12162 ( .A1(n13020), .A2(n9953), .ZN(n10402) );
  NAND2_X1 U12163 ( .A1(n19521), .A2(n19981), .ZN(n19456) );
  NOR2_X2 U12164 ( .A1(n14105), .A2(n14106), .ZN(n19296) );
  INV_X1 U12165 ( .A(n19295), .ZN(n19288) );
  INV_X1 U12166 ( .A(n19296), .ZN(n19290) );
  AND2_X1 U12167 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19795), .ZN(n19291) );
  INV_X1 U12168 ( .A(n19795), .ZN(n19495) );
  OR2_X1 U12169 ( .A1(n19854), .A2(n19851), .ZN(n13230) );
  INV_X1 U12170 ( .A(n16550), .ZN(n17474) );
  NOR3_X1 U12171 ( .A1(n16550), .A2(n16549), .A3(n18698), .ZN(n18660) );
  OAI22_X1 U12172 ( .A1(n16673), .A2(n9865), .B1(n9865), .B2(n10028), .ZN(
        n16651) );
  INV_X1 U12173 ( .A(n17622), .ZN(n10028) );
  NOR2_X1 U12174 ( .A1(n16651), .A2(n17607), .ZN(n16650) );
  NOR2_X1 U12175 ( .A1(n16692), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n16691) );
  NOR2_X1 U12176 ( .A1(n17495), .A2(n10066), .ZN(n10065) );
  AND2_X1 U12177 ( .A1(n10063), .A2(n9917), .ZN(n10062) );
  NOR2_X1 U12178 ( .A1(n17325), .A2(n10064), .ZN(n10063) );
  INV_X1 U12179 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17190) );
  AOI21_X1 U12180 ( .B1(n17175), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n12745), .ZN(n12746) );
  NOR2_X1 U12181 ( .A1(n12913), .A2(n9998), .ZN(n16551) );
  OAI21_X1 U12182 ( .B1(n13802), .B2(n13801), .A(n15643), .ZN(n15760) );
  NOR2_X1 U12183 ( .A1(n17473), .A2(n17436), .ZN(n17454) );
  INV_X1 U12184 ( .A(n17435), .ZN(n17436) );
  NOR2_X1 U12185 ( .A1(n17474), .A2(n17473), .ZN(n17475) );
  INV_X1 U12186 ( .A(n17914), .ZN(n15655) );
  INV_X1 U12187 ( .A(n16379), .ZN(n16381) );
  NAND2_X1 U12188 ( .A1(n17606), .A2(n9835), .ZN(n17543) );
  NOR2_X1 U12189 ( .A1(n17580), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U12190 ( .A1(n17606), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17579) );
  INV_X1 U12191 ( .A(n16694), .ZN(n17620) );
  NOR2_X1 U12192 ( .A1(n17658), .A2(n17660), .ZN(n17645) );
  AND2_X1 U12193 ( .A1(n10032), .A2(n10030), .ZN(n17719) );
  NOR2_X1 U12194 ( .A1(n17734), .A2(n10031), .ZN(n10030) );
  INV_X1 U12195 ( .A(n10033), .ZN(n10031) );
  NOR2_X1 U12196 ( .A1(n17828), .A2(n17806), .ZN(n17807) );
  INV_X1 U12197 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17806) );
  NAND2_X1 U12198 ( .A1(n10032), .A2(n10033), .ZN(n17733) );
  NOR2_X1 U12199 ( .A1(n17849), .A2(n17850), .ZN(n17768) );
  AND2_X1 U12200 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17868) );
  OR2_X1 U12201 ( .A1(n18737), .A2(n17891), .ZN(n17680) );
  INV_X1 U12202 ( .A(n10015), .ZN(n15745) );
  INV_X1 U12203 ( .A(n10013), .ZN(n17651) );
  NOR2_X1 U12204 ( .A1(n12815), .A2(n12814), .ZN(n17692) );
  NOR2_X1 U12205 ( .A1(n17717), .A2(n18037), .ZN(n18036) );
  NAND2_X1 U12206 ( .A1(n17732), .A2(n17966), .ZN(n18042) );
  INV_X1 U12207 ( .A(n15641), .ZN(n18693) );
  NOR2_X1 U12208 ( .A1(n17286), .A2(n12989), .ZN(n12932) );
  NOR2_X1 U12209 ( .A1(n12996), .A2(n12990), .ZN(n12991) );
  NOR2_X1 U12210 ( .A1(n15641), .A2(n15640), .ZN(n18698) );
  INV_X1 U12211 ( .A(n16551), .ZN(n18238) );
  NOR2_X1 U12212 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18237), .ZN(n18532) );
  OAI211_X1 U12213 ( .C1(n17218), .C2(n17186), .A(n12850), .B(n12849), .ZN(
        n18247) );
  AOI211_X1 U12214 ( .C1(n17043), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n12848), .B(n12847), .ZN(n12849) );
  OAI211_X1 U12215 ( .C1(n10239), .C2(n12906), .A(n12905), .B(n12904), .ZN(
        n18252) );
  INV_X1 U12216 ( .A(n13798), .ZN(n18257) );
  INV_X1 U12217 ( .A(n17286), .ZN(n18262) );
  AOI211_X1 U12218 ( .C1(n17043), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n12838), .B(n12837), .ZN(n12839) );
  INV_X1 U12219 ( .A(n18532), .ZN(n18346) );
  NAND2_X1 U12220 ( .A1(n10003), .A2(n10237), .ZN(n18668) );
  NAND2_X1 U12221 ( .A1(n18665), .A2(n13800), .ZN(n10003) );
  OR2_X1 U12222 ( .A1(n15705), .A2(n20005), .ZN(n13295) );
  OR2_X1 U12224 ( .A1(n20735), .A2(n20169), .ZN(n20005) );
  INV_X1 U12225 ( .A(n15851), .ZN(n20048) );
  AND2_X1 U12226 ( .A1(n14005), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14006) );
  AND2_X1 U12227 ( .A1(n14015), .A2(n14014), .ZN(n20096) );
  INV_X1 U12228 ( .A(n20102), .ZN(n20091) );
  NAND2_X1 U12229 ( .A1(n14015), .A2(n14009), .ZN(n20102) );
  INV_X1 U12230 ( .A(n20030), .ZN(n15767) );
  INV_X1 U12231 ( .A(n20084), .ZN(n20103) );
  INV_X1 U12232 ( .A(n15876), .ZN(n20111) );
  INV_X1 U12233 ( .A(n15900), .ZN(n14543) );
  INV_X1 U12234 ( .A(n14549), .ZN(n14279) );
  OR2_X1 U12235 ( .A1(n13571), .A2(n13570), .ZN(n13572) );
  OR2_X1 U12236 ( .A1(n15891), .A2(n13575), .ZN(n14549) );
  AND2_X1 U12237 ( .A1(n13543), .A2(n13348), .ZN(n20118) );
  INV_X1 U12238 ( .A(n13690), .ZN(n20153) );
  XNOR2_X1 U12239 ( .A(n13094), .B(n13184), .ZN(n14561) );
  OAI21_X1 U12240 ( .B1(n14359), .B2(n10258), .A(n9822), .ZN(n14580) );
  AND2_X1 U12241 ( .A1(n11722), .A2(n11678), .ZN(n14585) );
  OAI21_X1 U12242 ( .B1(n10259), .B2(n14410), .A(n14411), .ZN(n14620) );
  INV_X1 U12243 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15800) );
  INV_X1 U12244 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14677) );
  INV_X1 U12245 ( .A(n15955), .ZN(n20013) );
  INV_X1 U12246 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15961) );
  INV_X1 U12247 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13903) );
  AND3_X1 U12248 ( .A1(n20818), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n20688), 
        .ZN(n20166) );
  NAND2_X1 U12249 ( .A1(n10138), .A2(n10137), .ZN(n14328) );
  NAND2_X1 U12250 ( .A1(n10141), .A2(n14327), .ZN(n10137) );
  OR3_X1 U12251 ( .A1(n14733), .A2(n14714), .A3(n14713), .ZN(n14723) );
  NAND2_X1 U12252 ( .A1(n10103), .A2(n11826), .ZN(n15950) );
  NAND2_X1 U12253 ( .A1(n13942), .A2(n13941), .ZN(n10103) );
  AND2_X1 U12254 ( .A1(n13562), .A2(n13550), .ZN(n16068) );
  NAND2_X1 U12255 ( .A1(n13562), .A2(n15699), .ZN(n14757) );
  INV_X1 U12256 ( .A(n14255), .ZN(n14700) );
  NAND2_X1 U12257 ( .A1(n13562), .A2(n15675), .ZN(n14702) );
  INV_X1 U12258 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20610) );
  INV_X1 U12259 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20157) );
  NAND2_X1 U12260 ( .A1(n13762), .A2(n20334), .ZN(n20156) );
  OAI21_X1 U12261 ( .B1(n20350), .B2(n20335), .A(n20646), .ZN(n20353) );
  NOR2_X2 U12262 ( .A1(n20414), .A2(n20616), .ZN(n20403) );
  OAI211_X1 U12263 ( .C1(n20458), .C2(n20579), .A(n20500), .B(n20443), .ZN(
        n20461) );
  OAI211_X1 U12264 ( .C1(n20601), .C2(n20579), .A(n20646), .B(n20578), .ZN(
        n20604) );
  INV_X1 U12265 ( .A(n20636), .ZN(n20602) );
  AOI22_X1 U12266 ( .A1(n20577), .A2(n20574), .B1(n20572), .B2(n20571), .ZN(
        n20608) );
  OAI211_X1 U12267 ( .C1(n20670), .C2(n20647), .A(n20646), .B(n20645), .ZN(
        n20674) );
  NOR2_X1 U12268 ( .A1(n20334), .A2(n20163), .ZN(n20682) );
  NOR2_X1 U12269 ( .A1(n20334), .A2(n20181), .ZN(n20695) );
  NOR2_X1 U12270 ( .A1(n20334), .A2(n20187), .ZN(n20700) );
  NOR2_X1 U12271 ( .A1(n20334), .A2(n20194), .ZN(n20705) );
  NOR2_X1 U12272 ( .A1(n20334), .A2(n20200), .ZN(n20710) );
  NOR2_X1 U12273 ( .A1(n20334), .A2(n20207), .ZN(n20715) );
  NOR2_X1 U12274 ( .A1(n20334), .A2(n20213), .ZN(n20721) );
  NOR2_X2 U12275 ( .A1(n20685), .A2(n20545), .ZN(n20730) );
  NOR2_X1 U12276 ( .A1(n20334), .A2(n20219), .ZN(n20728) );
  INV_X1 U12277 ( .A(n13259), .ZN(n11908) );
  NAND2_X1 U12278 ( .A1(n16083), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20735) );
  INV_X2 U12279 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20813) );
  AND2_X1 U12280 ( .A1(n15725), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20736) );
  OAI21_X1 U12281 ( .B1(n10295), .B2(n15073), .A(n19094), .ZN(n10296) );
  NAND2_X1 U12282 ( .A1(n14827), .A2(n13929), .ZN(n16102) );
  NAND2_X1 U12283 ( .A1(n16102), .A2(n16103), .ZN(n16101) );
  INV_X1 U12284 ( .A(n12587), .ZN(n12574) );
  NAND2_X1 U12285 ( .A1(n14828), .A2(n15110), .ZN(n14827) );
  NAND2_X1 U12286 ( .A1(n16115), .A2(n16116), .ZN(n16114) );
  NAND2_X1 U12287 ( .A1(n16126), .A2(n16127), .ZN(n16125) );
  NAND2_X1 U12288 ( .A1(n16150), .A2(n16151), .ZN(n16149) );
  NAND2_X1 U12289 ( .A1(n18939), .A2(n13929), .ZN(n15670) );
  NAND2_X1 U12290 ( .A1(n15670), .A2(n16174), .ZN(n15669) );
  NAND2_X1 U12291 ( .A1(n18940), .A2(n18941), .ZN(n18939) );
  AND2_X1 U12292 ( .A1(n12517), .A2(n10121), .ZN(n12498) );
  AND2_X1 U12293 ( .A1(n12521), .A2(n12523), .ZN(n14853) );
  INV_X1 U12294 ( .A(n13929), .ZN(n19092) );
  AND2_X1 U12295 ( .A1(n18907), .A2(n10874), .ZN(n19101) );
  INV_X1 U12296 ( .A(n19049), .ZN(n19102) );
  NOR2_X1 U12297 ( .A1(n13929), .A2(n19048), .ZN(n19113) );
  INV_X1 U12298 ( .A(n19081), .ZN(n19109) );
  OR2_X1 U12299 ( .A1(n10799), .A2(n10798), .ZN(n13910) );
  NAND2_X1 U12300 ( .A1(n9834), .A2(n11974), .ZN(n10233) );
  NOR2_X1 U12301 ( .A1(n10230), .A2(n11973), .ZN(n10226) );
  OR2_X1 U12302 ( .A1(n10761), .A2(n10760), .ZN(n13581) );
  INV_X1 U12303 ( .A(n10230), .ZN(n10228) );
  AND2_X1 U12304 ( .A1(n15007), .A2(n15006), .ZN(n16097) );
  NAND2_X1 U12305 ( .A1(n19147), .A2(n10334), .ZN(n15065) );
  NOR2_X1 U12306 ( .A1(n19181), .A2(n19179), .ZN(n19156) );
  OR2_X1 U12307 ( .A1(n16165), .A2(n13670), .ZN(n19149) );
  NOR2_X1 U12308 ( .A1(n13342), .A2(n13341), .ZN(n19520) );
  INV_X1 U12309 ( .A(n19174), .ZN(n19181) );
  INV_X1 U12310 ( .A(n15065), .ZN(n19179) );
  INV_X1 U12311 ( .A(n19147), .ZN(n19178) );
  INV_X1 U12312 ( .A(n19149), .ZN(n19186) );
  INV_X2 U12313 ( .A(n19191), .ZN(n19223) );
  INV_X1 U12314 ( .A(n13529), .ZN(n19232) );
  XNOR2_X1 U12315 ( .A(n10264), .B(n10263), .ZN(n12675) );
  NAND2_X1 U12316 ( .A1(n10294), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10264) );
  NAND2_X1 U12317 ( .A1(n15232), .A2(n10197), .ZN(n16182) );
  INV_X1 U12318 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16241) );
  INV_X1 U12319 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16266) );
  INV_X1 U12320 ( .A(n16268), .ZN(n19253) );
  INV_X1 U12321 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16276) );
  INV_X1 U12322 ( .A(n19237), .ZN(n19246) );
  AND2_X1 U12323 ( .A1(n16275), .A2(n13269), .ZN(n16268) );
  INV_X1 U12324 ( .A(n16275), .ZN(n19245) );
  OR2_X1 U12325 ( .A1(n14897), .A2(n14896), .ZN(n16099) );
  OR2_X1 U12326 ( .A1(n14910), .A2(n14909), .ZN(n16112) );
  CLKBUF_X1 U12327 ( .A(n15140), .Z(n15141) );
  OR3_X1 U12328 ( .A1(n15357), .A2(n13066), .A3(n15152), .ZN(n15311) );
  NAND2_X1 U12329 ( .A1(n15334), .A2(n15335), .ZN(n10206) );
  NOR2_X1 U12330 ( .A1(n15406), .A2(n14124), .ZN(n14201) );
  NAND2_X1 U12331 ( .A1(n9988), .A2(n15171), .ZN(n9990) );
  NAND2_X1 U12332 ( .A1(n9852), .A2(n9989), .ZN(n9988) );
  AND2_X1 U12333 ( .A1(n14164), .A2(n14163), .ZN(n18995) );
  NAND2_X1 U12334 ( .A1(n15167), .A2(n15434), .ZN(n15438) );
  NOR2_X1 U12335 ( .A1(n15491), .A2(n15477), .ZN(n15450) );
  INV_X1 U12336 ( .A(n16307), .ZN(n16277) );
  NAND2_X1 U12337 ( .A1(n12462), .A2(n12461), .ZN(n15521) );
  INV_X1 U12338 ( .A(n19520), .ZN(n19981) );
  INV_X1 U12339 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19978) );
  XNOR2_X1 U12340 ( .A(n13335), .B(n13334), .ZN(n19974) );
  INV_X1 U12341 ( .A(n19521), .ZN(n19951) );
  INV_X1 U12342 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19960) );
  INV_X1 U12343 ( .A(n19974), .ZN(n19971) );
  XNOR2_X1 U12344 ( .A(n13362), .B(n13361), .ZN(n19961) );
  NAND2_X1 U12345 ( .A1(n16340), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15612) );
  NAND2_X1 U12346 ( .A1(n13499), .A2(n13420), .ZN(n19521) );
  NAND2_X1 U12347 ( .A1(n13414), .A2(n13419), .ZN(n13420) );
  INV_X1 U12348 ( .A(n13418), .ZN(n13419) );
  INV_X1 U12349 ( .A(n19393), .ZN(n19384) );
  OR2_X1 U12350 ( .A1(n19463), .A2(n19462), .ZN(n19488) );
  INV_X1 U12351 ( .A(n19482), .ZN(n19487) );
  NOR2_X1 U12352 ( .A1(n19952), .A2(n19456), .ZN(n19506) );
  OAI21_X1 U12353 ( .B1(n19549), .B2(n19528), .A(n19795), .ZN(n19555) );
  NAND2_X1 U12354 ( .A1(n19532), .A2(n19531), .ZN(n19554) );
  NOR2_X1 U12355 ( .A1(n19705), .A2(n19560), .ZN(n19606) );
  NOR2_X2 U12356 ( .A1(n19744), .A2(n19709), .ZN(n19740) );
  NOR2_X1 U12357 ( .A1(n19744), .A2(n19952), .ZN(n19773) );
  OAI21_X1 U12358 ( .B1(n19756), .B2(n19755), .A(n19754), .ZN(n19780) );
  NOR2_X1 U12359 ( .A1(n19705), .A2(n19709), .ZN(n19779) );
  OAI22_X1 U12360 ( .A1(n20220), .A2(n19290), .B1(n19289), .B2(n19288), .ZN(
        n19778) );
  INV_X1 U12361 ( .A(n19622), .ZN(n19788) );
  INV_X1 U12362 ( .A(n19762), .ZN(n19803) );
  INV_X1 U12363 ( .A(n19634), .ZN(n19801) );
  INV_X1 U12364 ( .A(n19724), .ZN(n19809) );
  INV_X1 U12365 ( .A(n19639), .ZN(n19807) );
  INV_X1 U12366 ( .A(n19644), .ZN(n19813) );
  OAI22_X1 U12367 ( .A1(n20210), .A2(n19290), .B1(n19279), .B2(n19288), .ZN(
        n19827) );
  AND2_X1 U12368 ( .A1(n19277), .A2(n19291), .ZN(n19825) );
  INV_X1 U12369 ( .A(n19738), .ZN(n19833) );
  INV_X1 U12370 ( .A(n19773), .ZN(n19846) );
  NOR2_X2 U12371 ( .A1(n19705), .A2(n19952), .ZN(n19842) );
  INV_X1 U12372 ( .A(n19666), .ZN(n19838) );
  INV_X1 U12373 ( .A(n19778), .ZN(n19847) );
  INV_X1 U12374 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19851) );
  AOI21_X1 U12375 ( .B1(n16366), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16367), 
        .ZN(n19850) );
  AND2_X1 U12376 ( .A1(n12980), .A2(n17474), .ZN(n16531) );
  NAND2_X1 U12377 ( .A1(n18878), .A2(n18661), .ZN(n17473) );
  NOR2_X1 U12378 ( .A1(n18660), .A2(n17473), .ZN(n18882) );
  NOR2_X1 U12379 ( .A1(n16673), .A2(n9865), .ZN(n16662) );
  NOR2_X1 U12380 ( .A1(n16662), .A2(n17622), .ZN(n16661) );
  NOR2_X1 U12381 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16802), .ZN(n16801) );
  INV_X1 U12382 ( .A(n16936), .ZN(n16901) );
  OAI211_X1 U12383 ( .C1(n18719), .C2(n18727), .A(n16881), .B(n18898), .ZN(
        n16936) );
  INV_X1 U12384 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17251) );
  INV_X1 U12385 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17253) );
  INV_X1 U12386 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17261) );
  INV_X1 U12387 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17270) );
  AND2_X1 U12388 ( .A1(n17310), .A2(n9848), .ZN(n17296) );
  NAND2_X1 U12389 ( .A1(n17310), .A2(n9847), .ZN(n17300) );
  INV_X1 U12390 ( .A(n17315), .ZN(n17310) );
  NAND2_X1 U12391 ( .A1(n17310), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17309) );
  AND2_X1 U12392 ( .A1(n17362), .A2(n10059), .ZN(n17316) );
  NOR2_X1 U12393 ( .A1(n18272), .A2(n10061), .ZN(n10059) );
  INV_X1 U12394 ( .A(n17341), .ZN(n17337) );
  NOR3_X1 U12395 ( .A1(n18272), .A2(n17358), .A3(n17325), .ZN(n17346) );
  NAND2_X1 U12396 ( .A1(n17362), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17358) );
  NAND2_X1 U12397 ( .A1(n10068), .A2(n9903), .ZN(n17398) );
  AOI211_X2 U12398 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n12708), .B(n12707), .ZN(n17411) );
  NOR2_X1 U12399 ( .A1(n12714), .A2(n12713), .ZN(n12722) );
  NOR2_X1 U12400 ( .A1(n17508), .A2(n17403), .ZN(n17427) );
  INV_X1 U12401 ( .A(n17433), .ZN(n17424) );
  CLKBUF_X1 U12402 ( .A(n17535), .Z(n17527) );
  NOR2_X1 U12403 ( .A1(n18885), .A2(n17527), .ZN(n17528) );
  OAI21_X1 U12404 ( .B1(n18885), .B2(n18886), .A(n17475), .ZN(n17535) );
  NOR2_X1 U12406 ( .A1(n15655), .A2(n15747), .ZN(n16405) );
  NAND2_X1 U12407 ( .A1(n17666), .A2(n9997), .ZN(n17562) );
  AND2_X1 U12408 ( .A1(n16397), .A2(n16396), .ZN(n9997) );
  NAND2_X1 U12409 ( .A1(n17562), .A2(n17923), .ZN(n9996) );
  INV_X1 U12410 ( .A(n17561), .ZN(n9995) );
  AOI21_X1 U12411 ( .B1(n17919), .B2(n17815), .A(n9993), .ZN(n9992) );
  NOR2_X1 U12412 ( .A1(n18221), .A2(n18808), .ZN(n9993) );
  NOR2_X1 U12413 ( .A1(n17968), .A2(n17705), .ZN(n17666) );
  NOR2_X1 U12414 ( .A1(n17694), .A2(n17698), .ZN(n17679) );
  NAND2_X1 U12415 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17848), .ZN(n17740) );
  NAND2_X1 U12416 ( .A1(n9825), .A2(n10002), .ZN(n17767) );
  INV_X1 U12417 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17828) );
  NOR2_X1 U12418 ( .A1(n17891), .A2(n17866), .ZN(n17848) );
  INV_X1 U12419 ( .A(n18608), .ZN(n18347) );
  INV_X1 U12420 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17892) );
  INV_X1 U12421 ( .A(n17899), .ZN(n17889) );
  NOR2_X2 U12422 ( .A1(n18346), .A2(n18393), .ZN(n18608) );
  INV_X1 U12423 ( .A(n17897), .ZN(n17908) );
  INV_X1 U12424 ( .A(n16385), .ZN(n17907) );
  NAND2_X1 U12425 ( .A1(n12823), .A2(n10014), .ZN(n15652) );
  AND2_X1 U12426 ( .A1(n18679), .A2(n18701), .ZN(n18057) );
  NOR2_X1 U12427 ( .A1(n18222), .A2(n17965), .ZN(n18020) );
  INV_X1 U12428 ( .A(n18679), .ZN(n18691) );
  AND2_X1 U12429 ( .A1(n10005), .A2(n10004), .ZN(n18679) );
  INV_X1 U12430 ( .A(n12993), .ZN(n10004) );
  OR2_X1 U12431 ( .A1(n15641), .A2(n12990), .ZN(n10005) );
  NAND2_X1 U12432 ( .A1(n17875), .A2(n12794), .ZN(n17862) );
  INV_X1 U12433 ( .A(n18665), .ZN(n18198) );
  INV_X1 U12434 ( .A(n18222), .ZN(n18206) );
  NOR2_X1 U12435 ( .A1(n18662), .A2(n18222), .ZN(n18220) );
  INV_X1 U12436 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18684) );
  NOR2_X1 U12437 ( .A1(n15648), .A2(n15647), .ZN(n18862) );
  INV_X1 U12438 ( .A(n18862), .ZN(n18860) );
  INV_X1 U12439 ( .A(n18815), .ZN(n18894) );
  AND2_X1 U12440 ( .A1(n13201), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20164)
         );
  AND2_X1 U12442 ( .A1(n13182), .A2(n10242), .ZN(n13183) );
  OAI21_X1 U12443 ( .B1(n14718), .B2(n15955), .A(n9861), .ZN(P1_U2968) );
  OAI21_X1 U12444 ( .B1(n15971), .B2(n15955), .A(n9961), .ZN(P1_U2973) );
  AOI21_X1 U12445 ( .B1(n15942), .B2(n14599), .A(n14598), .ZN(n9962) );
  NAND2_X1 U12446 ( .A1(n9868), .A2(n9973), .ZN(n15360) );
  AOI211_X1 U12447 ( .C1(n19119), .C2(n16307), .A(n10074), .B(n10072), .ZN(
        n13092) );
  OR2_X1 U12448 ( .A1(n13085), .A2(n10073), .ZN(n10072) );
  AOI21_X1 U12449 ( .B1(n15081), .B2(n16294), .A(n14318), .ZN(n14319) );
  NOR2_X1 U12450 ( .A1(n9857), .A2(n9981), .ZN(n9980) );
  INV_X1 U12451 ( .A(n15359), .ZN(n9981) );
  OAI21_X1 U12452 ( .B1(n16577), .B2(n9902), .A(n9830), .ZN(P3_U2640) );
  NAND2_X1 U12453 ( .A1(n16583), .A2(n16973), .ZN(n10039) );
  INV_X1 U12454 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16900) );
  NAND2_X1 U12455 ( .A1(n17362), .A2(n10060), .ZN(n17319) );
  NAND2_X1 U12456 ( .A1(n10068), .A2(n9843), .ZN(n17429) );
  NAND2_X1 U12457 ( .A1(n10010), .A2(n9819), .ZN(P3_U2799) );
  NAND2_X1 U12458 ( .A1(n16388), .A2(n17815), .ZN(n10010) );
  AOI21_X1 U12459 ( .B1(n16387), .B2(n18218), .A(n13016), .ZN(n13017) );
  AND3_X1 U12460 ( .A1(n16389), .A2(n9873), .A3(n9833), .ZN(n9819) );
  NAND2_X1 U12461 ( .A1(n15762), .A2(n15761), .ZN(n10068) );
  AND3_X1 U12462 ( .A1(n11974), .A2(n9834), .A3(n13910), .ZN(n9820) );
  OR2_X1 U12463 ( .A1(n15027), .A2(n15026), .ZN(n9821) );
  NAND2_X1 U12464 ( .A1(n14240), .A2(n14277), .ZN(n14276) );
  NAND2_X1 U12465 ( .A1(n12462), .A2(n9854), .ZN(n15498) );
  INV_X1 U12466 ( .A(n13557), .ZN(n20170) );
  AND2_X1 U12467 ( .A1(n9820), .A2(n13926), .ZN(n9823) );
  AND2_X1 U12468 ( .A1(n14487), .A2(n9885), .ZN(n14433) );
  AND2_X1 U12469 ( .A1(n10015), .A2(n9919), .ZN(n9824) );
  OR3_X1 U12470 ( .A1(n17907), .A2(n16386), .A3(n18089), .ZN(n9825) );
  AND2_X1 U12471 ( .A1(n10050), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9826) );
  OR2_X1 U12472 ( .A1(n10077), .A2(n14031), .ZN(n9827) );
  AND2_X1 U12473 ( .A1(n10055), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9828) );
  AND3_X1 U12474 ( .A1(n10042), .A2(n10040), .A3(n10039), .ZN(n9830) );
  AND3_X1 U12475 ( .A1(n12909), .A2(n12911), .A3(n9999), .ZN(n9831) );
  AND2_X1 U12476 ( .A1(n9881), .A2(n10142), .ZN(n9832) );
  OR2_X1 U12477 ( .A1(n17730), .A2(n16390), .ZN(n9833) );
  NAND3_X2 U12478 ( .A1(n19945), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19795), 
        .ZN(n14106) );
  OR2_X1 U12479 ( .A1(n10786), .A2(n10785), .ZN(n9834) );
  NAND2_X1 U12480 ( .A1(n10236), .A2(n9915), .ZN(n14200) );
  NAND2_X1 U12481 ( .A1(n14970), .A2(n9916), .ZN(n14950) );
  AND2_X1 U12482 ( .A1(n10037), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9835) );
  AND2_X1 U12483 ( .A1(n10047), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9836) );
  NAND2_X1 U12484 ( .A1(n10399), .A2(n10398), .ZN(n13020) );
  AND2_X1 U12485 ( .A1(n9915), .A2(n10235), .ZN(n9837) );
  NOR2_X1 U12486 ( .A1(n15406), .A2(n9904), .ZN(n14856) );
  AND2_X1 U12487 ( .A1(n10043), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9838) );
  AND2_X1 U12488 ( .A1(n9975), .A2(n16318), .ZN(n9839) );
  NAND2_X1 U12489 ( .A1(n11975), .A2(n11974), .ZN(n13685) );
  NOR2_X1 U12490 ( .A1(n13580), .A2(n10233), .ZN(n13783) );
  AND2_X1 U12491 ( .A1(n10057), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9840) );
  AND2_X1 U12492 ( .A1(n10089), .A2(n10088), .ZN(n9841) );
  AND2_X1 U12493 ( .A1(n10014), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9842) );
  AND2_X1 U12494 ( .A1(n18878), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n9843) );
  AND2_X1 U12495 ( .A1(n14930), .A2(n10134), .ZN(n9844) );
  AND2_X1 U12496 ( .A1(n9843), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n9845) );
  AND2_X1 U12497 ( .A1(n10197), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9846) );
  AND2_X1 U12498 ( .A1(n10065), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9847) );
  AND2_X1 U12499 ( .A1(n9847), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9848) );
  INV_X1 U12500 ( .A(n10480), .ZN(n10498) );
  NAND2_X1 U12501 ( .A1(n9818), .A2(n16325), .ZN(n9850) );
  OR2_X1 U12503 ( .A1(n10646), .A2(n10645), .ZN(n9851) );
  NOR2_X1 U12504 ( .A1(n15188), .A2(n15348), .ZN(n15159) );
  NAND2_X1 U12505 ( .A1(n14487), .A2(n10179), .ZN(n14420) );
  NAND2_X1 U12506 ( .A1(n15115), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15107) );
  AND2_X1 U12507 ( .A1(n14487), .A2(n11516), .ZN(n14488) );
  NAND2_X1 U12508 ( .A1(n15232), .A2(n15375), .ZN(n15223) );
  INV_X1 U12509 ( .A(n10192), .ZN(n15188) );
  NOR2_X1 U12510 ( .A1(n16917), .A2(n12682), .ZN(n12709) );
  AND2_X1 U12511 ( .A1(n9956), .A2(n9957), .ZN(n14232) );
  AND2_X1 U12512 ( .A1(n9956), .A2(n9954), .ZN(n14240) );
  NAND3_X1 U12513 ( .A1(n15170), .A2(n15400), .A3(n15228), .ZN(n9852) );
  AND2_X1 U12514 ( .A1(n14240), .A2(n10171), .ZN(n14493) );
  NAND2_X1 U12515 ( .A1(n14240), .A2(n10173), .ZN(n14445) );
  AND2_X1 U12516 ( .A1(n9968), .A2(n10408), .ZN(n9853) );
  OAI211_X1 U12517 ( .C1(n12697), .C2(n17251), .A(n12840), .B(n12839), .ZN(
        n18267) );
  AND2_X1 U12518 ( .A1(n12461), .A2(n12466), .ZN(n9854) );
  OR2_X1 U12519 ( .A1(n12484), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U12520 ( .A1(n10018), .A2(n12543), .ZN(n15334) );
  NAND2_X1 U12521 ( .A1(n12655), .A2(n12654), .ZN(n15504) );
  NAND2_X1 U12522 ( .A1(n10206), .A2(n15336), .ZN(n15160) );
  AND2_X1 U12523 ( .A1(n14383), .A2(n10180), .ZN(n13094) );
  AND2_X1 U12524 ( .A1(n12398), .A2(n12397), .ZN(n9856) );
  XNOR2_X1 U12525 ( .A(n12643), .B(n12644), .ZN(n12648) );
  INV_X1 U12526 ( .A(n12648), .ZN(n10188) );
  NAND2_X1 U12527 ( .A1(n15938), .A2(n14216), .ZN(n14244) );
  AND2_X1 U12528 ( .A1(n15358), .A2(n16294), .ZN(n9857) );
  NOR2_X1 U12529 ( .A1(n10130), .A2(n10129), .ZN(n10886) );
  AND2_X1 U12530 ( .A1(n14409), .A2(n10259), .ZN(n14395) );
  AND2_X1 U12531 ( .A1(n9814), .A2(n19110), .ZN(n9858) );
  NAND2_X1 U12532 ( .A1(n10423), .A2(n10450), .ZN(n10467) );
  AND2_X1 U12533 ( .A1(n12747), .A2(n12746), .ZN(n9859) );
  OR2_X1 U12534 ( .A1(n13262), .A2(n13345), .ZN(n9860) );
  AND2_X1 U12535 ( .A1(n11925), .A2(n11924), .ZN(n9861) );
  OR2_X1 U12536 ( .A1(n12164), .A2(n12163), .ZN(n9862) );
  AND2_X1 U12537 ( .A1(n10092), .A2(n11266), .ZN(n9863) );
  INV_X2 U12538 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16325) );
  OR2_X1 U12539 ( .A1(n14653), .A2(n11852), .ZN(n9864) );
  NAND2_X1 U12541 ( .A1(n12646), .A2(n12645), .ZN(n12656) );
  NAND3_X1 U12542 ( .A1(n10213), .A2(n10214), .A3(n15128), .ZN(n9866) );
  AND2_X1 U12543 ( .A1(n11054), .A2(n11053), .ZN(n13375) );
  NOR2_X1 U12544 ( .A1(n14956), .A2(n10223), .ZN(n12085) );
  NAND2_X1 U12545 ( .A1(n10205), .A2(n12554), .ZN(n9867) );
  AND2_X1 U12546 ( .A1(n9972), .A2(n9975), .ZN(n9868) );
  INV_X1 U12547 ( .A(n10409), .ZN(n10623) );
  AND2_X1 U12548 ( .A1(n12908), .A2(n12912), .ZN(n9869) );
  AND2_X1 U12549 ( .A1(n16378), .A2(n10033), .ZN(n9870) );
  AND2_X1 U12550 ( .A1(n13416), .A2(n10225), .ZN(n9871) );
  NAND2_X1 U12551 ( .A1(n12818), .A2(n12817), .ZN(n9872) );
  NAND2_X1 U12552 ( .A1(n16387), .A2(n17897), .ZN(n9873) );
  NAND2_X2 U12553 ( .A1(n11030), .A2(n13557), .ZN(n13131) );
  BUF_X1 U12554 ( .A(n11683), .Z(n11707) );
  AND2_X1 U12555 ( .A1(n10068), .A2(n9845), .ZN(n9874) );
  INV_X1 U12556 ( .A(n10268), .ZN(n10054) );
  INV_X1 U12557 ( .A(n12399), .ZN(n12571) );
  AND2_X1 U12558 ( .A1(n15338), .A2(n9841), .ZN(n9875) );
  AND2_X1 U12559 ( .A1(n10236), .A2(n9837), .ZN(n9876) );
  OR2_X1 U12560 ( .A1(n15491), .A2(n10086), .ZN(n14091) );
  OR2_X1 U12561 ( .A1(n19277), .A2(n10888), .ZN(n9877) );
  INV_X1 U12562 ( .A(n14216), .ZN(n10112) );
  AND2_X1 U12563 ( .A1(n17310), .A2(n10065), .ZN(n9878) );
  AND2_X1 U12564 ( .A1(n10275), .A2(n10050), .ZN(n9879) );
  OR2_X1 U12565 ( .A1(n10086), .A2(n14092), .ZN(n9880) );
  AND2_X1 U12566 ( .A1(n14144), .A2(n10143), .ZN(n9881) );
  AND2_X1 U12567 ( .A1(n11315), .A2(n13954), .ZN(n14024) );
  INV_X1 U12568 ( .A(n13797), .ZN(n12990) );
  AND3_X1 U12569 ( .A1(n11315), .A2(n13954), .A3(n14085), .ZN(n14084) );
  NOR2_X1 U12570 ( .A1(n14874), .A2(n14875), .ZN(n14873) );
  AND2_X1 U12571 ( .A1(n15793), .A2(n10145), .ZN(n9882) );
  NAND2_X1 U12572 ( .A1(n15553), .A2(n12632), .ZN(n14037) );
  NAND2_X1 U12573 ( .A1(n18897), .A2(n13799), .ZN(n18701) );
  AND2_X1 U12574 ( .A1(n14077), .A2(n10155), .ZN(n9883) );
  INV_X1 U12575 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20169) );
  OR3_X1 U12576 ( .A1(n10082), .A2(n14857), .A3(n10081), .ZN(n9884) );
  AND2_X1 U12577 ( .A1(n15768), .A2(n11516), .ZN(n9885) );
  INV_X1 U12578 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18906) );
  OR2_X1 U12579 ( .A1(n10658), .A2(n10657), .ZN(n12620) );
  INV_X1 U12580 ( .A(n15172), .ZN(n9989) );
  AND2_X1 U12581 ( .A1(n15062), .A2(n15363), .ZN(n15053) );
  INV_X1 U12582 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16251) );
  INV_X1 U12583 ( .A(n10232), .ZN(n10231) );
  INV_X1 U12584 ( .A(n11856), .ZN(n15918) );
  NOR2_X1 U12585 ( .A1(n9880), .A2(n10085), .ZN(n9886) );
  INV_X1 U12586 ( .A(n15182), .ZN(n9983) );
  AND2_X1 U12587 ( .A1(n10157), .A2(n10156), .ZN(n9887) );
  NOR2_X1 U12588 ( .A1(n11931), .A2(n10216), .ZN(n9888) );
  AND2_X1 U12589 ( .A1(n15208), .A2(n16175), .ZN(n9889) );
  AND2_X1 U12590 ( .A1(n10116), .A2(n12506), .ZN(n9890) );
  AND2_X1 U12591 ( .A1(n10121), .A2(n14961), .ZN(n9891) );
  OR2_X1 U12592 ( .A1(n15406), .A2(n10082), .ZN(n9892) );
  AND2_X1 U12593 ( .A1(n9832), .A2(n14238), .ZN(n9893) );
  INV_X1 U12594 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15231) );
  INV_X1 U12595 ( .A(n16313), .ZN(n16296) );
  NAND2_X1 U12596 ( .A1(n13416), .A2(n10231), .ZN(n10230) );
  INV_X2 U12597 ( .A(n12220), .ZN(n12058) );
  INV_X1 U12598 ( .A(n12108), .ZN(n10220) );
  NAND2_X1 U12599 ( .A1(n10229), .A2(n10228), .ZN(n13424) );
  AND2_X1 U12600 ( .A1(n10283), .A2(n10043), .ZN(n9894) );
  INV_X1 U12601 ( .A(n16318), .ZN(n16287) );
  AND2_X1 U12602 ( .A1(n13089), .A2(n19993), .ZN(n16318) );
  AND2_X1 U12603 ( .A1(n10280), .A2(n10047), .ZN(n9895) );
  AND2_X1 U12604 ( .A1(n13505), .A2(n13506), .ZN(n13504) );
  INV_X1 U12605 ( .A(n12516), .ZN(n10124) );
  OR2_X1 U12606 ( .A1(n10080), .A2(n10079), .ZN(n9896) );
  AND2_X1 U12607 ( .A1(n14145), .A2(n9832), .ZN(n9897) );
  INV_X1 U12608 ( .A(n12494), .ZN(n10120) );
  AOI21_X1 U12609 ( .B1(n10478), .B2(n11957), .A(n10477), .ZN(n13505) );
  INV_X1 U12610 ( .A(n12457), .ZN(n10128) );
  OR2_X1 U12611 ( .A1(n14444), .A2(n14547), .ZN(n9898) );
  NOR2_X1 U12612 ( .A1(n10285), .A2(n15143), .ZN(n10265) );
  AND2_X1 U12613 ( .A1(n10229), .A2(n10226), .ZN(n13579) );
  OR2_X1 U12614 ( .A1(n10699), .A2(n10698), .ZN(n12634) );
  INV_X1 U12615 ( .A(n12634), .ZN(n10211) );
  INV_X1 U12616 ( .A(n14121), .ZN(n10236) );
  INV_X1 U12617 ( .A(n14233), .ZN(n9957) );
  AND2_X1 U12618 ( .A1(n11382), .A2(n11381), .ZN(n14233) );
  AND2_X1 U12619 ( .A1(n14829), .A2(n10151), .ZN(n9899) );
  OR2_X1 U12620 ( .A1(n13978), .A2(n14031), .ZN(n10078) );
  AND2_X1 U12621 ( .A1(n9841), .A2(n15033), .ZN(n9900) );
  INV_X1 U12622 ( .A(n15569), .ZN(n9970) );
  NAND2_X1 U12623 ( .A1(n11042), .A2(n11041), .ZN(n13546) );
  AND2_X1 U12624 ( .A1(n10727), .A2(n10726), .ZN(n9901) );
  OR2_X1 U12625 ( .A1(n16919), .A2(n16578), .ZN(n9902) );
  AND2_X1 U12626 ( .A1(n9845), .A2(n17368), .ZN(n9903) );
  OR2_X1 U12627 ( .A1(n10082), .A2(n14857), .ZN(n9904) );
  AND2_X1 U12628 ( .A1(n11127), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n9905) );
  AND2_X1 U12629 ( .A1(n11127), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n9906) );
  AND2_X1 U12630 ( .A1(n11127), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n9907) );
  AND2_X1 U12631 ( .A1(n11127), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n9908) );
  AND2_X1 U12632 ( .A1(n11127), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n9909) );
  AND2_X1 U12633 ( .A1(n11127), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n9910) );
  OR2_X1 U12634 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9911) );
  AND2_X1 U12635 ( .A1(n13569), .A2(n13366), .ZN(n9912) );
  INV_X1 U12636 ( .A(n13115), .ZN(n13296) );
  INV_X1 U12637 ( .A(n14832), .ZN(n10080) );
  INV_X1 U12638 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10034) );
  INV_X1 U12639 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10045) );
  NOR2_X1 U12640 ( .A1(n20494), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n9913) );
  INV_X1 U12641 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10911) );
  AND2_X1 U12642 ( .A1(n17606), .A2(n10037), .ZN(n9914) );
  OR2_X1 U12643 ( .A1(n11999), .A2(n11998), .ZN(n9915) );
  OR2_X1 U12644 ( .A1(n12041), .A2(n12040), .ZN(n9916) );
  AND4_X1 U12645 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n9917)
         );
  INV_X1 U12646 ( .A(n10061), .ZN(n10060) );
  NAND2_X1 U12647 ( .A1(n10062), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n10061) );
  AND2_X1 U12648 ( .A1(n16006), .A2(n14782), .ZN(n9918) );
  INV_X1 U12649 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n10064) );
  INV_X1 U12650 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n10066) );
  INV_X1 U12651 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n10067) );
  INV_X1 U12652 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10048) );
  INV_X1 U12653 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10114) );
  INV_X1 U12654 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U12655 ( .A1(n18844), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9919) );
  INV_X1 U12656 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10052) );
  INV_X1 U12657 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10134) );
  INV_X1 U12658 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10058) );
  INV_X1 U12659 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11973) );
  OAI22_X2 U12660 ( .A1(n20197), .A2(n20224), .B1(n20196), .B2(n20225), .ZN(
        n20706) );
  OAI22_X2 U12661 ( .A1(n20208), .A2(n20225), .B1(n20973), .B2(n20224), .ZN(
        n20664) );
  NAND2_X1 U12662 ( .A1(n20166), .A2(n20165), .ZN(n20224) );
  INV_X1 U12663 ( .A(n20716), .ZN(n9920) );
  INV_X1 U12664 ( .A(n9920), .ZN(n9921) );
  INV_X1 U12665 ( .A(n20651), .ZN(n9922) );
  INV_X1 U12666 ( .A(n9922), .ZN(n9923) );
  INV_X1 U12667 ( .A(n20654), .ZN(n9924) );
  INV_X1 U12668 ( .A(n9924), .ZN(n9925) );
  INV_X1 U12669 ( .A(n20672), .ZN(n9926) );
  INV_X1 U12670 ( .A(n9926), .ZN(n9927) );
  INV_X1 U12671 ( .A(n20711), .ZN(n9928) );
  INV_X1 U12672 ( .A(n9928), .ZN(n9929) );
  INV_X1 U12673 ( .A(n20722), .ZN(n9930) );
  INV_X1 U12674 ( .A(n9930), .ZN(n9931) );
  INV_X1 U12675 ( .A(n20661), .ZN(n9932) );
  INV_X1 U12676 ( .A(n9932), .ZN(n9933) );
  INV_X1 U12677 ( .A(n20667), .ZN(n9934) );
  INV_X1 U12678 ( .A(n9934), .ZN(n9935) );
  INV_X1 U12679 ( .A(n20696), .ZN(n9936) );
  INV_X1 U12680 ( .A(n9936), .ZN(n9937) );
  INV_X1 U12681 ( .A(n20701), .ZN(n9938) );
  INV_X1 U12682 ( .A(n9938), .ZN(n9939) );
  INV_X1 U12683 ( .A(n20729), .ZN(n9940) );
  INV_X1 U12684 ( .A(n9940), .ZN(n9941) );
  INV_X1 U12685 ( .A(n20690), .ZN(n9942) );
  INV_X1 U12686 ( .A(n9942), .ZN(n9943) );
  INV_X1 U12687 ( .A(n20657), .ZN(n9944) );
  INV_X1 U12688 ( .A(n9944), .ZN(n9945) );
  AOI22_X2 U12689 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19295), .ZN(n19812) );
  NOR2_X2 U12690 ( .A1(n14107), .A2(n14106), .ZN(n19295) );
  OAI22_X2 U12691 ( .A1(n20167), .A2(n20225), .B1(n21012), .B2(n20224), .ZN(
        n20648) );
  NOR3_X4 U12692 ( .A1(n13447), .A2(n13446), .A3(n19869), .ZN(n19229) );
  NOR2_X2 U12693 ( .A1(n15129), .A2(n9946), .ZN(n15089) );
  XNOR2_X2 U12694 ( .A(n9947), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13090) );
  AND2_X2 U12695 ( .A1(n15232), .A2(n9846), .ZN(n15213) );
  NAND2_X2 U12696 ( .A1(n9948), .A2(n12659), .ZN(n15232) );
  NAND2_X1 U12697 ( .A1(n15504), .A2(n15505), .ZN(n9948) );
  AND2_X2 U12698 ( .A1(n15186), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10192) );
  NAND3_X1 U12699 ( .A1(n12362), .A2(n12360), .A3(n12354), .ZN(n9950) );
  NAND4_X1 U12700 ( .A1(n12361), .A2(n12353), .A3(n12359), .A4(n12355), .ZN(
        n9951) );
  XNOR2_X2 U12701 ( .A(n12633), .B(n9856), .ZN(n12639) );
  INV_X2 U12702 ( .A(n9953), .ZN(n14108) );
  NAND2_X1 U12703 ( .A1(n10412), .A2(n9953), .ZN(n10413) );
  NAND2_X1 U12704 ( .A1(n11363), .A2(n11362), .ZN(n14208) );
  INV_X1 U12705 ( .A(n11277), .ZN(n11190) );
  NAND2_X2 U12706 ( .A1(n9958), .A2(n11167), .ZN(n11277) );
  INV_X1 U12707 ( .A(n11251), .ZN(n9958) );
  XNOR2_X1 U12708 ( .A(n11107), .B(n11106), .ZN(n11251) );
  AND2_X2 U12709 ( .A1(n14395), .A2(n14394), .ZN(n14383) );
  NAND2_X1 U12710 ( .A1(n20822), .A2(n11046), .ZN(n9964) );
  INV_X1 U12711 ( .A(n13115), .ZN(n9965) );
  OAI21_X2 U12712 ( .B1(n13788), .B2(n11447), .A(n11284), .ZN(n13656) );
  NAND2_X1 U12713 ( .A1(n14167), .A2(n14168), .ZN(n9966) );
  NAND2_X1 U12714 ( .A1(n9966), .A2(n12428), .ZN(n15242) );
  INV_X2 U12715 ( .A(n12368), .ZN(n12438) );
  NAND2_X2 U12716 ( .A1(n9971), .A2(n10212), .ZN(n12633) );
  NAND3_X1 U12717 ( .A1(n9973), .A2(n9839), .A3(n9972), .ZN(n9982) );
  NAND2_X1 U12718 ( .A1(n9982), .A2(n9980), .ZN(P2_U3025) );
  NAND2_X1 U12719 ( .A1(n16178), .A2(n9889), .ZN(n15192) );
  XNOR2_X1 U12720 ( .A(n9990), .B(n15394), .ZN(n16190) );
  INV_X4 U12721 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16933) );
  NAND4_X1 U12722 ( .A1(n9994), .A2(n17564), .A3(n9992), .A4(n9991), .ZN(
        P3_U2803) );
  INV_X1 U12723 ( .A(n17563), .ZN(n9991) );
  NAND2_X1 U12724 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  NAND3_X1 U12725 ( .A1(n12910), .A2(n9869), .A3(n9831), .ZN(n9998) );
  INV_X1 U12726 ( .A(n17767), .ZN(n17802) );
  NAND2_X1 U12727 ( .A1(n17897), .A2(n17732), .ZN(n10002) );
  NAND2_X1 U12729 ( .A1(n12794), .A2(n10008), .ZN(n10007) );
  NAND2_X1 U12730 ( .A1(n17894), .A2(n12788), .ZN(n17886) );
  XNOR2_X1 U12731 ( .A(n12964), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17895) );
  NAND3_X1 U12732 ( .A1(n17597), .A2(n17602), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12819) );
  NAND2_X2 U12733 ( .A1(n10013), .A2(n10012), .ZN(n17675) );
  OR2_X2 U12734 ( .A1(n17682), .A2(n17814), .ZN(n10013) );
  AND2_X2 U12735 ( .A1(n17811), .A2(n18089), .ZN(n17778) );
  AND2_X2 U12736 ( .A1(n10113), .A2(n18089), .ZN(n18136) );
  AND2_X1 U12737 ( .A1(n12823), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17558) );
  NAND2_X1 U12738 ( .A1(n12823), .A2(n9842), .ZN(n10015) );
  INV_X2 U12739 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18849) );
  NAND2_X1 U12740 ( .A1(n15226), .A2(n10019), .ZN(n10017) );
  NAND3_X1 U12741 ( .A1(n12562), .A2(n10022), .A3(n10024), .ZN(n15102) );
  NAND2_X1 U12742 ( .A1(n10024), .A2(n15149), .ZN(n15150) );
  AND2_X1 U12743 ( .A1(n10023), .A2(n12562), .ZN(n15126) );
  OAI21_X1 U12744 ( .B1(n10417), .B2(n19259), .A(n9953), .ZN(n10025) );
  NAND2_X2 U12745 ( .A1(n13224), .A2(n13035), .ZN(n12283) );
  NAND2_X2 U12746 ( .A1(n19259), .A2(n19264), .ZN(n13035) );
  NAND2_X2 U12747 ( .A1(n10431), .A2(n13048), .ZN(n13224) );
  INV_X4 U12748 ( .A(n19259), .ZN(n13048) );
  NAND2_X1 U12749 ( .A1(n15442), .A2(n12488), .ZN(n15167) );
  XNOR2_X2 U12750 ( .A(n10027), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16891) );
  INV_X1 U12751 ( .A(n17734), .ZN(n10029) );
  NAND3_X1 U12752 ( .A1(n10032), .A2(n9870), .A3(n10029), .ZN(n17694) );
  NAND2_X1 U12753 ( .A1(n17606), .A2(n10035), .ZN(n16412) );
  NOR2_X1 U12754 ( .A1(n16586), .A2(n9865), .ZN(n16577) );
  INV_X2 U12755 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18839) );
  NAND2_X1 U12756 ( .A1(n13978), .A2(n15534), .ZN(n10075) );
  NAND2_X1 U12757 ( .A1(n10075), .A2(n10076), .ZN(n15536) );
  INV_X1 U12758 ( .A(n10078), .ZN(n14032) );
  INV_X1 U12759 ( .A(n14185), .ZN(n10077) );
  NOR2_X1 U12760 ( .A1(n9821), .A2(n15018), .ZN(n15019) );
  INV_X1 U12761 ( .A(n10869), .ZN(n15007) );
  AOI22_X1 U12762 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10675) );
  INV_X1 U12763 ( .A(n15491), .ZN(n10084) );
  NAND2_X1 U12764 ( .A1(n10084), .A2(n9886), .ZN(n14874) );
  NAND2_X1 U12765 ( .A1(n15338), .A2(n9900), .ZN(n15027) );
  NOR2_X2 U12766 ( .A1(n11051), .A2(n11045), .ZN(n11914) );
  NAND2_X1 U12767 ( .A1(n11033), .A2(n11231), .ZN(n11051) );
  XNOR2_X2 U12768 ( .A(n11110), .B(n11109), .ZN(n11269) );
  NAND2_X1 U12769 ( .A1(n10091), .A2(n11268), .ZN(n11267) );
  NAND2_X1 U12770 ( .A1(n11269), .A2(n20169), .ZN(n10091) );
  INV_X1 U12771 ( .A(n10095), .ZN(n12828) );
  INV_X1 U12772 ( .A(n12827), .ZN(n10094) );
  NAND2_X1 U12773 ( .A1(n13942), .A2(n10097), .ZN(n10096) );
  NAND2_X1 U12774 ( .A1(n10096), .A2(n10099), .ZN(n14136) );
  NOR2_X2 U12775 ( .A1(n17565), .A2(n12821), .ZN(n12823) );
  NOR2_X2 U12776 ( .A1(n17566), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17565) );
  AND2_X2 U12777 ( .A1(n10918), .A2(n10917), .ZN(n10973) );
  NAND2_X1 U12778 ( .A1(n10110), .A2(n10111), .ZN(n14647) );
  NAND3_X1 U12779 ( .A1(n10111), .A2(n9918), .A3(n10110), .ZN(n14639) );
  NAND2_X2 U12780 ( .A1(n11190), .A2(n13791), .ZN(n11287) );
  NAND2_X1 U12782 ( .A1(n12487), .A2(n9890), .ZN(n12501) );
  NAND2_X1 U12783 ( .A1(n12517), .A2(n9891), .ZN(n12546) );
  NAND2_X1 U12784 ( .A1(n12517), .A2(n12516), .ZN(n12520) );
  INV_X1 U12785 ( .A(n12400), .ZN(n10130) );
  NAND2_X1 U12786 ( .A1(n12499), .A2(n10131), .ZN(n12567) );
  NAND2_X1 U12787 ( .A1(n12499), .A2(n12544), .ZN(n12550) );
  INV_X1 U12788 ( .A(n10141), .ZN(n14325) );
  NAND2_X1 U12789 ( .A1(n14145), .A2(n9893), .ZN(n14791) );
  NOR2_X2 U12790 ( .A1(n10418), .A2(n10408), .ZN(n10149) );
  NAND4_X1 U12791 ( .A1(n13569), .A2(n13546), .A3(n13366), .A4(n9860), .ZN(
        n10165) );
  NAND2_X1 U12792 ( .A1(n13253), .A2(n20183), .ZN(n13366) );
  NAND2_X2 U12793 ( .A1(n10165), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11076) );
  NAND3_X1 U12794 ( .A1(n11043), .A2(n13540), .A3(n11031), .ZN(n10960) );
  NAND2_X1 U12795 ( .A1(n11774), .A2(n11257), .ZN(n10167) );
  NAND2_X1 U12796 ( .A1(n10167), .A2(n10168), .ZN(n13614) );
  NAND2_X1 U12797 ( .A1(n10170), .A2(n11276), .ZN(n13613) );
  INV_X1 U12798 ( .A(n13614), .ZN(n10170) );
  NOR2_X2 U12799 ( .A1(n11287), .A2(n10176), .ZN(n11302) );
  NAND2_X1 U12800 ( .A1(n11302), .A2(n11303), .ZN(n11816) );
  INV_X1 U12801 ( .A(n14421), .ZN(n10178) );
  XNOR2_X1 U12802 ( .A(n11364), .B(n11365), .ZN(n14210) );
  NAND2_X1 U12803 ( .A1(n14383), .A2(n14384), .ZN(n14370) );
  NOR2_X1 U12804 ( .A1(n14371), .A2(n14370), .ZN(n14359) );
  XNOR2_X2 U12805 ( .A(n10455), .B(n10200), .ZN(n11938) );
  AND3_X2 U12806 ( .A1(n10438), .A2(n10185), .A3(n10439), .ZN(n10200) );
  NAND2_X1 U12807 ( .A1(n9810), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10185) );
  NAND2_X1 U12808 ( .A1(n10467), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10186) );
  NAND2_X1 U12809 ( .A1(n14176), .A2(n10187), .ZN(n10189) );
  NAND2_X1 U12810 ( .A1(n14176), .A2(n14172), .ZN(n12649) );
  NAND3_X1 U12811 ( .A1(n12641), .A2(n10189), .A3(n12642), .ZN(n15240) );
  NOR2_X2 U12812 ( .A1(n15129), .A2(n15286), .ZN(n15115) );
  NAND3_X1 U12813 ( .A1(n12406), .A2(n15552), .A3(n12635), .ZN(n15553) );
  NAND3_X1 U12814 ( .A1(n10199), .A2(n12345), .A3(n10198), .ZN(n12635) );
  NAND2_X1 U12815 ( .A1(n12345), .A2(n12344), .ZN(n12405) );
  NAND2_X1 U12816 ( .A1(n10456), .A2(n10200), .ZN(n10457) );
  AND3_X4 U12817 ( .A1(n10202), .A2(n10201), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U12818 ( .A1(n15161), .A2(n10204), .ZN(n10205) );
  AND2_X2 U12819 ( .A1(n10435), .A2(n13054), .ZN(n12286) );
  AND2_X1 U12820 ( .A1(n10435), .A2(n13041), .ZN(n10210) );
  NAND2_X2 U12821 ( .A1(n13226), .A2(n13048), .ZN(n13231) );
  NAND2_X1 U12822 ( .A1(n11946), .A2(n10215), .ZN(n13361) );
  NAND2_X1 U12823 ( .A1(n10217), .A2(n9888), .ZN(n10215) );
  NAND2_X1 U12824 ( .A1(n10217), .A2(n11929), .ZN(n11932) );
  NAND2_X1 U12825 ( .A1(n14956), .A2(n10220), .ZN(n10218) );
  NAND2_X1 U12826 ( .A1(n13413), .A2(n11970), .ZN(n10229) );
  NAND2_X1 U12827 ( .A1(n10229), .A2(n9871), .ZN(n13580) );
  NAND2_X1 U12828 ( .A1(n19264), .A2(n11972), .ZN(n10232) );
  NAND2_X1 U12829 ( .A1(n11975), .A2(n9820), .ZN(n13908) );
  NOR2_X2 U12830 ( .A1(n14121), .A2(n10234), .ZN(n14969) );
  OAI21_X1 U12831 ( .B1(n14512), .B2(n14503), .A(n13183), .ZN(P1_U2843) );
  AOI21_X1 U12832 ( .B1(n13095), .B2(n9822), .A(n13094), .ZN(n14568) );
  AND2_X1 U12833 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10979) );
  AOI22_X1 U12834 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11141), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10949) );
  INV_X1 U12835 ( .A(n14176), .ZN(n12640) );
  NAND2_X1 U12836 ( .A1(n10371), .A2(n16325), .ZN(n10372) );
  NAND2_X1 U12837 ( .A1(n11063), .A2(n11062), .ZN(n11064) );
  NAND2_X1 U12838 ( .A1(n14944), .A2(n14843), .ZN(n14842) );
  OR2_X1 U12839 ( .A1(n11162), .A2(n11164), .ZN(n11165) );
  NAND2_X1 U12840 ( .A1(n12558), .A2(n12559), .ZN(n15149) );
  NAND2_X1 U12841 ( .A1(n11945), .A2(n11944), .ZN(n13362) );
  AOI22_X1 U12842 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U12843 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10324) );
  NAND2_X1 U12844 ( .A1(n10313), .A2(n16325), .ZN(n10320) );
  NAND2_X1 U12845 ( .A1(n10330), .A2(n16325), .ZN(n10331) );
  NAND2_X1 U12846 ( .A1(n13090), .A2(n19248), .ZN(n12679) );
  AND2_X1 U12847 ( .A1(n15226), .A2(n15436), .ZN(n15227) );
  OAI22_X1 U12848 ( .A1(n10467), .A2(n10440), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10481), .ZN(n10444) );
  INV_X1 U12849 ( .A(n13362), .ZN(n11948) );
  OR2_X1 U12850 ( .A1(n18662), .A2(n16376), .ZN(n10237) );
  XOR2_X1 U12851 ( .A(n12804), .B(n12953), .Z(n10238) );
  INV_X1 U12852 ( .A(n18089), .ZN(n17731) );
  INV_X1 U12853 ( .A(n18221), .ZN(n18144) );
  OR2_X1 U12854 ( .A1(n14315), .A2(n14314), .ZN(n10241) );
  OR2_X1 U12855 ( .A1(n20919), .A2(n14492), .ZN(n10242) );
  NOR2_X1 U12856 ( .A1(n14276), .A2(n14547), .ZN(n10243) );
  OR2_X1 U12857 ( .A1(n17193), .A2(n17157), .ZN(n10244) );
  OR2_X1 U12858 ( .A1(n10239), .A2(n17215), .ZN(n10245) );
  OR2_X1 U12859 ( .A1(n12697), .A2(n17247), .ZN(n10246) );
  OR2_X1 U12860 ( .A1(n21024), .A2(n14492), .ZN(n10247) );
  AND3_X1 U12861 ( .A1(n12893), .A2(n12892), .A3(n10246), .ZN(n10248) );
  AND4_X1 U12862 ( .A1(n10302), .A2(n10301), .A3(n10300), .A4(n10299), .ZN(
        n10249) );
  NOR2_X1 U12863 ( .A1(n15159), .A2(n15333), .ZN(n10250) );
  INV_X1 U12864 ( .A(n17777), .ZN(n17814) );
  NOR2_X1 U12865 ( .A1(n14447), .A2(n15767), .ZN(n10251) );
  INV_X1 U12866 ( .A(n11040), .ZN(n11041) );
  OR2_X1 U12867 ( .A1(n11231), .A2(n20813), .ZN(n11272) );
  INV_X1 U12868 ( .A(n14503), .ZN(n20112) );
  INV_X1 U12869 ( .A(n11447), .ZN(n11395) );
  AND3_X1 U12870 ( .A1(n12588), .A2(n12571), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10253) );
  INV_X1 U12871 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11316) );
  AND3_X1 U12872 ( .A1(n10304), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10303), .ZN(n10254) );
  NAND2_X1 U12873 ( .A1(n20169), .A2(n20168), .ZN(n20334) );
  INV_X1 U12874 ( .A(n20815), .ZN(n14003) );
  AND2_X1 U12875 ( .A1(n10382), .A2(n16325), .ZN(n10255) );
  INV_X1 U12876 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15152) );
  INV_X1 U12877 ( .A(n10482), .ZN(n10486) );
  INV_X1 U12878 ( .A(n9804), .ZN(n13982) );
  INV_X1 U12879 ( .A(n13424), .ZN(n13607) );
  AND2_X1 U12880 ( .A1(n11700), .A2(n11699), .ZN(n10258) );
  AND2_X1 U12881 ( .A1(n11611), .A2(n11610), .ZN(n10259) );
  AND3_X1 U12882 ( .A1(n10982), .A2(n10981), .A3(n10980), .ZN(n10260) );
  AND4_X1 U12883 ( .A1(n10946), .A2(n10945), .A3(n10944), .A4(n10943), .ZN(
        n10261) );
  INV_X1 U12884 ( .A(n14806), .ZN(n13531) );
  AND4_X1 U12885 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10262) );
  INV_X1 U12886 ( .A(n13375), .ZN(n11055) );
  NAND2_X1 U12887 ( .A1(n14806), .A2(n11055), .ZN(n11056) );
  AOI21_X1 U12888 ( .B1(n20209), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11895), 
        .ZN(n11884) );
  OR2_X1 U12889 ( .A1(n11881), .A2(n11880), .ZN(n11861) );
  AOI22_X1 U12890 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U12891 ( .A1(n11139), .A2(n11138), .ZN(n11162) );
  AOI22_X1 U12892 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10342) );
  AND2_X1 U12893 ( .A1(n10333), .A2(n19292), .ZN(n10430) );
  NAND2_X1 U12894 ( .A1(n10623), .A2(n10333), .ZN(n10410) );
  AND2_X1 U12895 ( .A1(n10569), .A2(n10568), .ZN(n10579) );
  INV_X1 U12896 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10912) );
  BUF_X1 U12897 ( .A(n11683), .Z(n11637) );
  NAND2_X1 U12898 ( .A1(n11080), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11066) );
  XNOR2_X1 U12899 ( .A(n11162), .B(n11163), .ZN(n11258) );
  OAI21_X1 U12900 ( .B1(n11962), .B2(n10464), .A(n11950), .ZN(n10466) );
  INV_X1 U12901 ( .A(n12633), .ZN(n12429) );
  NOR2_X1 U12902 ( .A1(n17218), .A2(n17267), .ZN(n12745) );
  AND2_X1 U12903 ( .A1(n11871), .A2(n11870), .ZN(n11904) );
  INV_X1 U12904 ( .A(n14489), .ZN(n11516) );
  INV_X1 U12905 ( .A(n13615), .ZN(n11276) );
  INV_X1 U12906 ( .A(n11808), .ZN(n11818) );
  NOR2_X1 U12907 ( .A1(n10578), .A2(n10573), .ZN(n10574) );
  NAND2_X1 U12908 ( .A1(n10345), .A2(n16325), .ZN(n10346) );
  INV_X1 U12909 ( .A(n15522), .ZN(n12466) );
  NAND2_X1 U12910 ( .A1(n10379), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10386) );
  AND2_X1 U12911 ( .A1(n10876), .A2(n10880), .ZN(n12270) );
  INV_X1 U12912 ( .A(n11365), .ZN(n11366) );
  AND2_X1 U12913 ( .A1(n11537), .A2(n11536), .ZN(n15768) );
  NAND2_X1 U12914 ( .A1(n13531), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11720) );
  NAND2_X1 U12915 ( .A1(n20215), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11447) );
  NOR2_X1 U12916 ( .A1(n11104), .A2(n11103), .ZN(n11778) );
  BUF_X1 U12917 ( .A(n11168), .Z(n13755) );
  INV_X1 U12918 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15688) );
  INV_X1 U12919 ( .A(n11834), .ZN(n11159) );
  AOI21_X1 U12920 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19960), .A(
        n10574), .ZN(n10576) );
  INV_X1 U12921 ( .A(n9798), .ZN(n10666) );
  NAND2_X1 U12922 ( .A1(n12587), .A2(n12586), .ZN(n12593) );
  AND2_X1 U12923 ( .A1(n13047), .A2(n14108), .ZN(n10420) );
  AND2_X1 U12924 ( .A1(n13043), .A2(n10447), .ZN(n10454) );
  INV_X1 U12925 ( .A(n12278), .ZN(n13054) );
  NAND2_X1 U12926 ( .A1(n12782), .A2(n10245), .ZN(n12783) );
  NAND2_X1 U12927 ( .A1(n10238), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12805) );
  OR2_X1 U12928 ( .A1(n11920), .A2(n14553), .ZN(n11922) );
  AND2_X1 U12929 ( .A1(n20813), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11757) );
  AND4_X1 U12930 ( .A1(n11025), .A2(n11024), .A3(n11023), .A4(n11022), .ZN(
        n11026) );
  OR2_X1 U12931 ( .A1(n14566), .A2(n11750), .ZN(n11726) );
  NOR2_X1 U12932 ( .A1(n11531), .A2(n15786), .ZN(n11534) );
  NAND2_X1 U12933 ( .A1(n11173), .A2(n11172), .ZN(n20328) );
  OAI21_X1 U12934 ( .B1(n13259), .B2(n11907), .A(n11906), .ZN(n11911) );
  AOI221_X1 U12935 ( .B1(n10576), .B2(n13228), .C1(n10576), .C2(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n10575), .ZN(n12612) );
  NAND2_X1 U12936 ( .A1(n12412), .A2(n12415), .ZN(n12411) );
  AND3_X1 U12937 ( .A1(n10551), .A2(n10550), .A3(n10549), .ZN(n14919) );
  AND3_X1 U12938 ( .A1(n10542), .A2(n10541), .A3(n10540), .ZN(n14943) );
  INV_X2 U12939 ( .A(n10505), .ZN(n12663) );
  AND3_X1 U12940 ( .A1(n10518), .A2(n10517), .A3(n10516), .ZN(n14162) );
  INV_X1 U12941 ( .A(n15085), .ZN(n12590) );
  INV_X1 U12942 ( .A(n12558), .ZN(n12561) );
  NOR2_X1 U12943 ( .A1(n15507), .A2(n15528), .ZN(n15488) );
  NOR2_X1 U12944 ( .A1(n16664), .A2(n16565), .ZN(n17577) );
  NAND2_X1 U12945 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12711) );
  NOR4_X2 U12946 ( .A1(n12998), .A2(n18262), .A3(n12984), .A4(n16551), .ZN(
        n16550) );
  OR2_X1 U12947 ( .A1(n12807), .A2(n12806), .ZN(n12808) );
  NOR2_X1 U12948 ( .A1(n12784), .A2(n12783), .ZN(n12785) );
  AND2_X1 U12949 ( .A1(n12820), .A2(n17814), .ZN(n12821) );
  INV_X1 U12950 ( .A(n16424), .ZN(n16427) );
  OR2_X1 U12951 ( .A1(n12871), .A2(n12870), .ZN(n12872) );
  AND2_X1 U12952 ( .A1(n14373), .A2(n14335), .ZN(n14336) );
  OR2_X1 U12953 ( .A1(n14406), .A2(n14334), .ZN(n14385) );
  NOR2_X1 U12954 ( .A1(n11383), .A2(n14677), .ZN(n11398) );
  XNOR2_X1 U12955 ( .A(n11922), .B(n11921), .ZN(n14005) );
  NOR2_X1 U12956 ( .A1(n14003), .A2(n9812), .ZN(n14015) );
  INV_X1 U12957 ( .A(n20096), .ZN(n20073) );
  NAND2_X1 U12958 ( .A1(n11314), .A2(n11313), .ZN(n13956) );
  INV_X1 U12959 ( .A(n11759), .ZN(n11760) );
  INV_X1 U12960 ( .A(n14487), .ZN(n15791) );
  NAND2_X1 U12961 ( .A1(n11415), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11432) );
  AND2_X1 U12962 ( .A1(n13593), .A2(n13592), .ZN(n14255) );
  AND2_X1 U12963 ( .A1(n14757), .A2(n14701), .ZN(n14706) );
  OR2_X1 U12964 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20540) );
  INV_X1 U12965 ( .A(n20637), .ZN(n20380) );
  NOR2_X1 U12966 ( .A1(n20572), .A2(n20334), .ZN(n20500) );
  OR2_X1 U12967 ( .A1(n13763), .A2(n20159), .ZN(n20326) );
  INV_X2 U12968 ( .A(n11032), .ZN(n20215) );
  INV_X1 U12969 ( .A(n19107), .ZN(n19087) );
  AND3_X1 U12970 ( .A1(n10524), .A2(n10523), .A3(n10522), .ZN(n14989) );
  NOR2_X1 U12971 ( .A1(n14839), .A2(n12399), .ZN(n15104) );
  AND2_X1 U12972 ( .A1(n15304), .A2(n13070), .ZN(n15248) );
  AND2_X1 U12973 ( .A1(n10847), .A2(n10846), .ZN(n14857) );
  AND2_X1 U12974 ( .A1(n12505), .A2(n15173), .ZN(n15394) );
  OR2_X1 U12975 ( .A1(n12533), .A2(n15415), .ZN(n15398) );
  AND3_X1 U12976 ( .A1(n10607), .A2(n10606), .A3(n10605), .ZN(n14092) );
  XNOR2_X1 U12977 ( .A(n11953), .B(n11950), .ZN(n11926) );
  OAI21_X1 U12978 ( .B1(n16369), .B2(n19984), .A(n15612), .ZN(n12669) );
  AND2_X1 U12979 ( .A1(n13219), .A2(n13218), .ZN(n16351) );
  NAND2_X1 U12980 ( .A1(n19961), .A2(n19971), .ZN(n19560) );
  OR2_X1 U12981 ( .A1(n19627), .A2(n19621), .ZN(n19668) );
  NAND2_X1 U12982 ( .A1(n19951), .A2(n19520), .ZN(n19705) );
  INV_X1 U12983 ( .A(n16529), .ZN(n18661) );
  NOR2_X1 U12984 ( .A1(n18898), .A2(n16551), .ZN(n16552) );
  AND2_X1 U12985 ( .A1(n16683), .A2(n16691), .ZN(n16685) );
  NOR2_X1 U12986 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16768), .ZN(n16754) );
  NOR2_X1 U12987 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16844), .ZN(n16818) );
  INV_X1 U12988 ( .A(n16931), .ZN(n16924) );
  NOR2_X1 U12989 ( .A1(n17618), .A2(n17909), .ZN(n17914) );
  NOR2_X1 U12990 ( .A1(n16724), .A2(n16726), .ZN(n17657) );
  NOR2_X1 U12991 ( .A1(n17411), .A2(n12799), .ZN(n12804) );
  INV_X1 U12992 ( .A(n18136), .ZN(n17813) );
  NOR2_X1 U12993 ( .A1(n12954), .A2(n17411), .ZN(n17837) );
  INV_X1 U12994 ( .A(n18682), .ZN(n18673) );
  INV_X1 U12995 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17186) );
  AND2_X1 U12996 ( .A1(n15707), .A2(n20011), .ZN(n13543) );
  NOR2_X1 U12997 ( .A1(n14226), .A2(n14473), .ZN(n15843) );
  OR2_X1 U12998 ( .A1(n20815), .A2(n14000), .ZN(n20029) );
  NAND2_X1 U12999 ( .A1(n11298), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11306) );
  AND2_X1 U13000 ( .A1(n20029), .A2(n14006), .ZN(n20075) );
  OR2_X1 U13001 ( .A1(n14730), .A2(n15876), .ZN(n13182) );
  NAND2_X1 U13002 ( .A1(n15822), .A2(n14448), .ZN(n15812) );
  INV_X1 U13003 ( .A(n14492), .ZN(n14480) );
  AND2_X1 U13004 ( .A1(n14551), .A2(n14302), .ZN(n15887) );
  INV_X1 U13005 ( .A(n14551), .ZN(n15891) );
  NAND2_X1 U13006 ( .A1(n11498), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11531) );
  NAND2_X1 U13007 ( .A1(n11307), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11317) );
  INV_X1 U13008 ( .A(n15954), .ZN(n15942) );
  INV_X1 U13009 ( .A(n14712), .ZN(n14771) );
  NOR2_X1 U13010 ( .A1(n14250), .A2(n14248), .ZN(n13943) );
  INV_X1 U13011 ( .A(n14757), .ZN(n14692) );
  AND2_X1 U13012 ( .A1(n13562), .A2(n13552), .ZN(n16067) );
  NOR2_X1 U13013 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20798) );
  OAI211_X1 U13014 ( .C1(n20327), .C2(n20813), .A(n20500), .B(n20177), .ZN(
        n20227) );
  NOR2_X2 U13015 ( .A1(n20300), .A2(n20326), .ZN(n20253) );
  OAI211_X1 U13016 ( .C1(n20263), .C2(n20262), .A(n20500), .B(n20261), .ZN(
        n20289) );
  NOR2_X2 U13017 ( .A1(n20300), .A2(n20380), .ZN(n20321) );
  NOR2_X2 U13018 ( .A1(n20300), .A2(n20545), .ZN(n20352) );
  OAI211_X1 U13019 ( .C1(n20402), .C2(n20579), .A(n20646), .B(n20387), .ZN(
        n20404) );
  NOR2_X2 U13020 ( .A1(n20414), .A2(n20380), .ZN(n20432) );
  NOR2_X1 U13021 ( .A1(n11774), .A2(n13791), .ZN(n20409) );
  AND2_X1 U13022 ( .A1(n20490), .A2(n20469), .ZN(n20527) );
  OAI21_X1 U13023 ( .B1(n20544), .B2(n20543), .A(n20542), .ZN(n20563) );
  NOR2_X2 U13024 ( .A1(n20546), .A2(n20545), .ZN(n20603) );
  INV_X1 U13025 ( .A(n20326), .ZN(n20567) );
  NOR2_X2 U13026 ( .A1(n20685), .A2(n20616), .ZN(n20673) );
  NAND2_X1 U13027 ( .A1(n14841), .A2(n15153), .ZN(n14840) );
  NAND2_X1 U13028 ( .A1(n16087), .A2(n10900), .ZN(n19107) );
  INV_X1 U13029 ( .A(n19105), .ZN(n19039) );
  OR2_X1 U13030 ( .A1(n18907), .A2(n10904), .ZN(n19049) );
  AND2_X1 U13031 ( .A1(n10895), .A2(n10586), .ZN(n19081) );
  OR2_X1 U13032 ( .A1(n10604), .A2(n10603), .ZN(n13926) );
  INV_X1 U13033 ( .A(n15000), .ZN(n14984) );
  INV_X1 U13034 ( .A(n13452), .ZN(n13521) );
  NOR2_X1 U13035 ( .A1(n15121), .A2(n15103), .ZN(n15106) );
  AND2_X1 U13036 ( .A1(n10902), .A2(n19851), .ZN(n19235) );
  AND2_X1 U13037 ( .A1(n15176), .A2(n15175), .ZN(n15218) );
  AND2_X1 U13038 ( .A1(n13034), .A2(n16359), .ZN(n13089) );
  AND2_X1 U13039 ( .A1(n12669), .A2(n18906), .ZN(n19795) );
  INV_X1 U13040 ( .A(n16351), .ZN(n16330) );
  OAI21_X1 U13041 ( .B1(n14115), .B2(n14114), .A(n14113), .ZN(n19297) );
  NOR2_X2 U13042 ( .A1(n19560), .A2(n19456), .ZN(n19323) );
  NOR2_X1 U13043 ( .A1(n19560), .A2(n19491), .ZN(n19348) );
  INV_X1 U13044 ( .A(n19424), .ZN(n19416) );
  NAND2_X1 U13045 ( .A1(n19961), .A2(n19974), .ZN(n19946) );
  INV_X1 U13046 ( .A(n19448), .ZN(n19451) );
  AND2_X1 U13047 ( .A1(n19467), .A2(n19466), .ZN(n19486) );
  INV_X1 U13048 ( .A(n19558), .ZN(n19546) );
  OR2_X1 U13049 ( .A1(n19961), .A2(n19971), .ZN(n19952) );
  OAI21_X1 U13050 ( .B1(n19595), .B2(n19611), .A(n19795), .ZN(n19613) );
  NOR2_X1 U13051 ( .A1(n19744), .A2(n19946), .ZN(n19670) );
  NOR2_X1 U13052 ( .A1(n19705), .A2(n19946), .ZN(n19678) );
  INV_X1 U13053 ( .A(n19818), .ZN(n19725) );
  INV_X1 U13054 ( .A(n19830), .ZN(n19769) );
  INV_X1 U13055 ( .A(n19718), .ZN(n19797) );
  OAI22_X1 U13056 ( .A1(n20214), .A2(n19290), .B1(n19282), .B2(n19288), .ZN(
        n19735) );
  INV_X1 U13057 ( .A(n13230), .ZN(n16359) );
  INV_X1 U13058 ( .A(n18882), .ZN(n18898) );
  INV_X1 U13059 ( .A(n18701), .ZN(n18667) );
  NAND2_X1 U13060 ( .A1(n18716), .A2(n16552), .ZN(n16925) );
  NOR2_X1 U13061 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16738), .ZN(n16731) );
  NOR2_X1 U13062 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16792), .ZN(n16772) );
  NOR3_X1 U13063 ( .A1(n16878), .A2(n17257), .A3(n17256), .ZN(n17252) );
  NAND4_X1 U13064 ( .A1(n18878), .A2(n18244), .A3(n18238), .A4(n15760), .ZN(
        n17257) );
  INV_X1 U13065 ( .A(n18036), .ZN(n17618) );
  NOR2_X1 U13066 ( .A1(n12976), .A2(n17803), .ZN(n18090) );
  INV_X1 U13067 ( .A(n17404), .ZN(n16386) );
  INV_X1 U13068 ( .A(n18181), .ZN(n18218) );
  NOR2_X1 U13069 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18832), .ZN(
        n18856) );
  INV_X1 U13070 ( .A(n18715), .ZN(n18878) );
  INV_X1 U13071 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18739) );
  NAND2_X1 U13072 ( .A1(n13543), .A2(n11037), .ZN(n13431) );
  INV_X1 U13073 ( .A(n20098), .ZN(n15826) );
  NAND2_X1 U13074 ( .A1(n20029), .A2(n14001), .ZN(n15851) );
  AND2_X1 U13075 ( .A1(n13572), .A2(n20011), .ZN(n14551) );
  INV_X2 U13076 ( .A(n15888), .ZN(n15896) );
  INV_X1 U13077 ( .A(n20118), .ZN(n20143) );
  NAND2_X1 U13078 ( .A1(n15960), .A2(n11919), .ZN(n15954) );
  INV_X1 U13079 ( .A(n16067), .ZN(n16046) );
  OR3_X1 U13080 ( .A1(n14773), .A2(n14772), .A3(n16052), .ZN(n14781) );
  INV_X1 U13081 ( .A(n16068), .ZN(n16052) );
  INV_X1 U13082 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20573) );
  INV_X1 U13083 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16077) );
  AOI22_X1 U13084 ( .A1(n20176), .A2(n20173), .B1(n20496), .B2(n20327), .ZN(
        n20230) );
  OR2_X1 U13085 ( .A1(n20300), .A2(n20616), .ZN(n20287) );
  AOI22_X1 U13086 ( .A1(n20260), .A2(n20262), .B1(n9913), .B2(n20496), .ZN(
        n20292) );
  INV_X1 U13087 ( .A(n20299), .ZN(n20325) );
  NAND2_X1 U13088 ( .A1(n20409), .A2(n20567), .ZN(n20379) );
  AOI22_X1 U13089 ( .A1(n20386), .A2(n20383), .B1(n9913), .B2(n20572), .ZN(
        n20407) );
  NAND2_X1 U13090 ( .A1(n20409), .A2(n20408), .ZN(n20439) );
  NAND2_X1 U13091 ( .A1(n20490), .A2(n20567), .ZN(n20489) );
  AOI22_X1 U13092 ( .A1(n20497), .A2(n20501), .B1(n20496), .B2(n20495), .ZN(
        n20532) );
  NAND2_X1 U13093 ( .A1(n20490), .A2(n20637), .ZN(n20566) );
  INV_X1 U13094 ( .A(n20695), .ZN(n20585) );
  INV_X1 U13095 ( .A(n20721), .ZN(n20600) );
  NAND2_X1 U13096 ( .A1(n20638), .A2(n20567), .ZN(n20636) );
  NAND2_X1 U13097 ( .A1(n20638), .A2(n20637), .ZN(n20734) );
  INV_X1 U13098 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16083) );
  AND2_X1 U13099 ( .A1(n20003), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20830) );
  NOR2_X1 U13100 ( .A1(n13205), .A2(n10585), .ZN(n18907) );
  NOR2_X1 U13101 ( .A1(n10875), .A2(n10907), .ZN(n10908) );
  OR2_X1 U13102 ( .A1(n10897), .A2(n10896), .ZN(n19105) );
  INV_X1 U13103 ( .A(n19101), .ZN(n19085) );
  INV_X1 U13104 ( .A(n16215), .ZN(n15428) );
  NAND2_X1 U13105 ( .A1(n13337), .A2(n16359), .ZN(n14998) );
  AND2_X1 U13106 ( .A1(n12288), .A2(n16359), .ZN(n19147) );
  NAND2_X1 U13107 ( .A1(n10623), .A2(n19147), .ZN(n19174) );
  NAND2_X1 U13108 ( .A1(n13234), .A2(n19863), .ZN(n19226) );
  NAND2_X1 U13109 ( .A1(n13445), .A2(n13446), .ZN(n13529) );
  OR2_X1 U13110 ( .A1(n12618), .A2(n13035), .ZN(n19237) );
  INV_X1 U13111 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16230) );
  INV_X1 U13112 ( .A(n19248), .ZN(n16260) );
  INV_X1 U13113 ( .A(n15564), .ZN(n19110) );
  INV_X1 U13114 ( .A(n16294), .ZN(n16314) );
  INV_X1 U13115 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19968) );
  INV_X1 U13116 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13228) );
  AOI21_X1 U13117 ( .B1(n14104), .B2(n14114), .A(n14103), .ZN(n19300) );
  INV_X1 U13118 ( .A(n19348), .ZN(n19358) );
  OR2_X1 U13119 ( .A1(n19456), .A2(n19946), .ZN(n19393) );
  OR2_X1 U13120 ( .A1(n19491), .A2(n19946), .ZN(n19424) );
  OR2_X1 U13121 ( .A1(n19456), .A2(n19709), .ZN(n19448) );
  OR2_X1 U13122 ( .A1(n19491), .A2(n19709), .ZN(n19482) );
  INV_X1 U13123 ( .A(n19506), .ZN(n19519) );
  OR2_X1 U13124 ( .A1(n19491), .A2(n19952), .ZN(n19558) );
  NAND2_X1 U13125 ( .A1(n19523), .A2(n19522), .ZN(n19589) );
  INV_X1 U13126 ( .A(n19606), .ZN(n19616) );
  INV_X1 U13127 ( .A(n19670), .ZN(n19664) );
  INV_X1 U13128 ( .A(n19678), .ZN(n19704) );
  INV_X1 U13129 ( .A(n19827), .ZN(n19772) );
  INV_X1 U13130 ( .A(n19779), .ZN(n19776) );
  INV_X1 U13131 ( .A(n19735), .ZN(n19836) );
  INV_X1 U13132 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19855) );
  INV_X1 U13133 ( .A(n19944), .ZN(n19857) );
  INV_X1 U13134 ( .A(n16932), .ZN(n16879) );
  INV_X1 U13135 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17850) );
  NOR2_X1 U13136 ( .A1(n16942), .A2(n16993), .ZN(n16997) );
  AND2_X1 U13137 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17059), .ZN(n17074) );
  INV_X1 U13138 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17247) );
  NAND2_X1 U13139 ( .A1(n18678), .A2(n17428), .ZN(n17421) );
  NAND2_X1 U13140 ( .A1(n17454), .A2(n18238), .ZN(n17453) );
  INV_X1 U13141 ( .A(n17454), .ZN(n17472) );
  INV_X1 U13142 ( .A(n17816), .ZN(n17730) );
  NAND2_X1 U13143 ( .A1(n16386), .A2(n16385), .ZN(n17790) );
  INV_X1 U13144 ( .A(n18020), .ZN(n18034) );
  INV_X1 U13145 ( .A(n18220), .ZN(n18214) );
  INV_X1 U13146 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18683) );
  INV_X1 U13147 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18234) );
  INV_X1 U13148 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18829) );
  INV_X1 U13149 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18832) );
  INV_X1 U13150 ( .A(n18828), .ZN(n18738) );
  INV_X1 U13151 ( .A(n18894), .ZN(n18821) );
  NOR2_X1 U13152 ( .A1(n18739), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18815) );
  CLKBUF_X1 U13153 ( .A(n16524), .Z(n20831) );
  OAI21_X1 U13154 ( .B1(n14561), .B2(n14503), .A(n13189), .ZN(P1_U2842) );
  NAND2_X1 U13155 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10269), .ZN(
        n10268) );
  INV_X1 U13156 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18999) );
  INV_X1 U13157 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15220) );
  INV_X1 U13158 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18957) );
  INV_X1 U13159 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18932) );
  INV_X1 U13160 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15143) );
  INV_X1 U13161 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15117) );
  INV_X1 U13162 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10289) );
  INV_X1 U13163 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15090) );
  XNOR2_X1 U13164 ( .A(n10294), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15073) );
  INV_X1 U13165 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12666) );
  INV_X1 U13166 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10263) );
  AOI22_X4 U13167 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12666), .B1(n12675), 
        .B2(n18906), .ZN(n13929) );
  AOI21_X1 U13168 ( .B1(n15143), .B2(n10285), .A(n10265), .ZN(n15146) );
  INV_X1 U13169 ( .A(n15146), .ZN(n16138) );
  OAI21_X1 U13170 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10266), .A(
        n10282), .ZN(n18951) );
  AOI21_X1 U13171 ( .B1(n18957), .B2(n10281), .A(n10266), .ZN(n18963) );
  AOI21_X1 U13172 ( .B1(n15220), .B2(n10279), .A(n9895), .ZN(n18971) );
  AOI21_X1 U13173 ( .B1(n18999), .B2(n10277), .A(n10280), .ZN(n19005) );
  AOI21_X1 U13174 ( .B1(n15231), .B2(n10276), .A(n10278), .ZN(n19012) );
  AOI21_X1 U13175 ( .B1(n16230), .B2(n10274), .A(n9879), .ZN(n19031) );
  AOI21_X1 U13176 ( .B1(n16241), .B2(n10272), .A(n10275), .ZN(n19056) );
  AOI21_X1 U13177 ( .B1(n16251), .B2(n10270), .A(n10273), .ZN(n16253) );
  AOI21_X1 U13178 ( .B1(n16266), .B2(n10268), .A(n10271), .ZN(n19079) );
  AOI21_X1 U13179 ( .B1(n16276), .B2(n10267), .A(n10269), .ZN(n16267) );
  OAI22_X1 U13180 ( .A1(n18906), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19118) );
  INV_X1 U13181 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14883) );
  OAI22_X1 U13182 ( .A1(n18906), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14883), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14881) );
  AND2_X1 U13183 ( .A1(n19118), .A2(n14881), .ZN(n13988) );
  OAI21_X1 U13184 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n10267), .ZN(n19252) );
  NAND2_X1 U13185 ( .A1(n13988), .A2(n19252), .ZN(n13973) );
  NOR2_X1 U13186 ( .A1(n16267), .A2(n13973), .ZN(n19091) );
  OAI21_X1 U13187 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10269), .A(
        n10268), .ZN(n19243) );
  NAND2_X1 U13188 ( .A1(n19091), .A2(n19243), .ZN(n19077) );
  NOR2_X1 U13189 ( .A1(n19079), .A2(n19077), .ZN(n19064) );
  OAI21_X1 U13190 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10271), .A(
        n10270), .ZN(n19066) );
  NAND2_X1 U13191 ( .A1(n19064), .A2(n19066), .ZN(n13958) );
  NOR2_X1 U13192 ( .A1(n16253), .A2(n13958), .ZN(n13930) );
  OAI21_X1 U13193 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10273), .A(
        n10272), .ZN(n16250) );
  NAND2_X1 U13194 ( .A1(n13930), .A2(n16250), .ZN(n19054) );
  NOR2_X1 U13195 ( .A1(n19056), .A2(n19054), .ZN(n19036) );
  OAI21_X1 U13196 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10275), .A(
        n10274), .ZN(n19038) );
  NAND2_X1 U13197 ( .A1(n19036), .A2(n19038), .ZN(n19029) );
  NOR2_X1 U13198 ( .A1(n19031), .A2(n19029), .ZN(n14088) );
  OAI21_X1 U13199 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9879), .A(
        n10276), .ZN(n16223) );
  NAND2_X1 U13200 ( .A1(n14088), .A2(n16223), .ZN(n19011) );
  NOR2_X1 U13201 ( .A1(n19012), .A2(n19011), .ZN(n19010) );
  OAI21_X1 U13202 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10278), .A(
        n10277), .ZN(n16214) );
  NAND2_X1 U13203 ( .A1(n19010), .A2(n16214), .ZN(n19006) );
  NOR2_X1 U13204 ( .A1(n19005), .A2(n19006), .ZN(n18987) );
  OAI21_X1 U13205 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10280), .A(
        n10279), .ZN(n18988) );
  NAND2_X1 U13206 ( .A1(n18987), .A2(n18988), .ZN(n18970) );
  NOR2_X1 U13207 ( .A1(n18971), .A2(n18970), .ZN(n18969) );
  OAI21_X1 U13208 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n9895), .A(
        n10281), .ZN(n16186) );
  NAND2_X1 U13209 ( .A1(n18969), .A2(n16186), .ZN(n18961) );
  OAI21_X1 U13210 ( .B1(n18963), .B2(n18961), .A(n13929), .ZN(n18950) );
  NAND2_X1 U13211 ( .A1(n18951), .A2(n18950), .ZN(n18949) );
  NAND2_X1 U13212 ( .A1(n18949), .A2(n13929), .ZN(n18940) );
  AOI21_X1 U13213 ( .B1(n10282), .B2(n18932), .A(n10283), .ZN(n15183) );
  INV_X1 U13214 ( .A(n15183), .ZN(n18941) );
  OAI21_X1 U13215 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10283), .A(
        n10284), .ZN(n16174) );
  NAND2_X1 U13216 ( .A1(n13929), .A2(n15669), .ZN(n16150) );
  AOI21_X1 U13217 ( .B1(n10045), .B2(n10284), .A(n9894), .ZN(n15163) );
  INV_X1 U13218 ( .A(n15163), .ZN(n16151) );
  NAND2_X1 U13219 ( .A1(n13929), .A2(n16149), .ZN(n14841) );
  OAI21_X1 U13220 ( .B1(n9894), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n10285), .ZN(n15153) );
  NAND2_X1 U13221 ( .A1(n13929), .A2(n14840), .ZN(n16137) );
  NAND2_X1 U13222 ( .A1(n16138), .A2(n16137), .ZN(n16136) );
  NAND2_X1 U13223 ( .A1(n16136), .A2(n13929), .ZN(n16126) );
  OR2_X1 U13224 ( .A1(n10265), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10286) );
  NAND2_X1 U13225 ( .A1(n10288), .A2(n10286), .ZN(n16127) );
  NAND2_X1 U13226 ( .A1(n13929), .A2(n16125), .ZN(n16115) );
  INV_X1 U13227 ( .A(n10290), .ZN(n10287) );
  AOI21_X1 U13228 ( .B1(n15117), .B2(n10288), .A(n10287), .ZN(n15120) );
  INV_X1 U13229 ( .A(n15120), .ZN(n16116) );
  NAND2_X1 U13230 ( .A1(n13929), .A2(n16114), .ZN(n14828) );
  NAND2_X1 U13231 ( .A1(n10290), .A2(n10289), .ZN(n10291) );
  NAND2_X1 U13232 ( .A1(n10292), .A2(n10291), .ZN(n15110) );
  AND2_X1 U13233 ( .A1(n10292), .A2(n15090), .ZN(n10293) );
  NOR2_X1 U13234 ( .A1(n10294), .A2(n10293), .ZN(n15092) );
  INV_X1 U13235 ( .A(n15092), .ZN(n16103) );
  NAND2_X1 U13236 ( .A1(n13929), .A2(n16101), .ZN(n10295) );
  NAND2_X1 U13237 ( .A1(n15073), .A2(n10295), .ZN(n16095) );
  INV_X1 U13238 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19457) );
  NAND4_X1 U13239 ( .A1(n19851), .A2(n18906), .A3(n19457), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19048) );
  INV_X1 U13240 ( .A(n19048), .ZN(n19094) );
  INV_X1 U13241 ( .A(n10296), .ZN(n10297) );
  NAND2_X1 U13242 ( .A1(n16095), .A2(n10297), .ZN(n10909) );
  AND2_X4 U13243 ( .A1(n15571), .A2(n10202), .ZN(n10353) );
  NOR2_X4 U13244 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15570) );
  AOI22_X1 U13245 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10301) );
  AND2_X4 U13246 ( .A1(n15570), .A2(n10202), .ZN(n10387) );
  AND2_X4 U13247 ( .A1(n10298), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12243) );
  AOI22_X1 U13248 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U13249 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10299) );
  NAND2_X1 U13250 ( .A1(n10249), .A2(n16325), .ZN(n10308) );
  AOI22_X1 U13251 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13252 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13253 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13254 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10305) );
  NAND3_X1 U13255 ( .A1(n10254), .A2(n10306), .A3(n10305), .ZN(n10307) );
  NAND2_X2 U13256 ( .A1(n10308), .A2(n10307), .ZN(n10401) );
  AOI22_X1 U13257 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13258 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13259 ( .A1(n12245), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10310) );
  NAND4_X1 U13260 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n10309), .ZN(
        n10313) );
  AOI22_X1 U13261 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13262 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13263 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U13264 ( .A1(n12245), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10314) );
  NAND4_X1 U13265 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10318) );
  NAND2_X1 U13266 ( .A1(n10318), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10319) );
  NAND2_X2 U13267 ( .A1(n10320), .A2(n10319), .ZN(n19283) );
  AOI22_X1 U13268 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13269 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10322) );
  AOI22_X1 U13270 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10321) );
  NAND4_X1 U13271 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10325) );
  AOI22_X1 U13272 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13273 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12245), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13274 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13275 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10326) );
  NAND4_X1 U13276 ( .A1(n10329), .A2(n10328), .A3(n10327), .A4(n10326), .ZN(
        n10330) );
  NAND2_X4 U13277 ( .A1(n10332), .A2(n10331), .ZN(n19292) );
  INV_X1 U13278 ( .A(n10401), .ZN(n10333) );
  AOI22_X1 U13279 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U13280 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13281 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13282 ( .A1(n12245), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10336) );
  NAND4_X1 U13283 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n10340) );
  NAND2_X1 U13284 ( .A1(n10340), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10347) );
  AOI22_X1 U13285 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13286 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13287 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10341) );
  NAND4_X1 U13288 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10345) );
  NAND2_X2 U13289 ( .A1(n11930), .A2(n10407), .ZN(n10409) );
  AOI22_X1 U13290 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13291 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13292 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13293 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10348) );
  NAND4_X1 U13294 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10352) );
  NAND2_X1 U13295 ( .A1(n10352), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10360) );
  AOI22_X1 U13296 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13297 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13298 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13299 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10354) );
  NAND4_X1 U13300 ( .A1(n10357), .A2(n10356), .A3(n10355), .A4(n10354), .ZN(
        n10358) );
  NAND2_X4 U13301 ( .A1(n10360), .A2(n10359), .ZN(n19264) );
  NAND2_X1 U13302 ( .A1(n10412), .A2(n10361), .ZN(n10445) );
  AOI22_X1 U13303 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13304 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13305 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13306 ( .A1(n12053), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10362) );
  NAND2_X1 U13307 ( .A1(n10366), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10373) );
  AOI22_X1 U13308 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13309 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13310 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10368) );
  AOI22_X1 U13311 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10367) );
  AND2_X4 U13312 ( .A1(n10373), .A2(n10372), .ZN(n19259) );
  NAND2_X1 U13313 ( .A1(n10445), .A2(n13048), .ZN(n10406) );
  AOI22_X1 U13314 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9818), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13315 ( .A1(n9801), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13316 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13317 ( .A1(n12245), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U13318 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13319 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13320 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13321 ( .A1(n12245), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10382) );
  NAND3_X1 U13322 ( .A1(n10384), .A2(n10383), .A3(n10255), .ZN(n10385) );
  NAND2_X1 U13323 ( .A1(n10409), .A2(n14108), .ZN(n10400) );
  AOI22_X1 U13324 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13325 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13326 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13327 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10388) );
  NAND4_X1 U13328 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10392) );
  NAND2_X1 U13329 ( .A1(n10392), .A2(n16325), .ZN(n10399) );
  AOI22_X1 U13330 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9817), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13331 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10335), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U13332 ( .A1(n9808), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13333 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10393) );
  NAND4_X1 U13334 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10397) );
  NAND2_X1 U13335 ( .A1(n10397), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10398) );
  NAND2_X1 U13336 ( .A1(n10400), .A2(n13047), .ZN(n10404) );
  INV_X1 U13337 ( .A(n13226), .ZN(n10403) );
  OAI211_X1 U13338 ( .C1(n10405), .C2(n10404), .A(n10403), .B(n13048), .ZN(
        n13050) );
  NAND2_X1 U13339 ( .A1(n10417), .A2(n10408), .ZN(n12276) );
  NAND2_X1 U13340 ( .A1(n12276), .A2(n10401), .ZN(n10411) );
  NAND2_X1 U13341 ( .A1(n13024), .A2(n19292), .ZN(n13044) );
  NAND2_X1 U13342 ( .A1(n13044), .A2(n14108), .ZN(n10414) );
  NAND2_X1 U13343 ( .A1(n10414), .A2(n10413), .ZN(n10446) );
  NAND2_X1 U13344 ( .A1(n10446), .A2(n10436), .ZN(n10415) );
  NAND2_X1 U13345 ( .A1(n10447), .A2(n10415), .ZN(n10416) );
  NAND2_X1 U13346 ( .A1(n10416), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10423) );
  INV_X1 U13347 ( .A(n10418), .ZN(n10419) );
  INV_X1 U13348 ( .A(n16363), .ZN(n10422) );
  NAND3_X1 U13349 ( .A1(n13088), .A2(n13047), .A3(n19264), .ZN(n10421) );
  NAND2_X1 U13350 ( .A1(n18906), .A2(n19855), .ZN(n14822) );
  INV_X1 U13351 ( .A(n13224), .ZN(n13041) );
  AND3_X1 U13352 ( .A1(n10587), .A2(n19283), .A3(n19292), .ZN(n10424) );
  NAND3_X1 U13353 ( .A1(n13054), .A2(n13041), .A3(n10424), .ZN(n13036) );
  NAND2_X1 U13354 ( .A1(n13036), .A2(n13231), .ZN(n10425) );
  NAND2_X1 U13355 ( .A1(n10425), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10432) );
  INV_X1 U13356 ( .A(n10437), .ZN(n10426) );
  OAI211_X1 U13357 ( .C1(n14822), .C2(n19978), .A(n10432), .B(n10426), .ZN(
        n10427) );
  INV_X1 U13358 ( .A(n10427), .ZN(n10428) );
  NAND2_X1 U13359 ( .A1(n13038), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10442) );
  NAND2_X1 U13360 ( .A1(n10437), .A2(n13446), .ZN(n10433) );
  NOR2_X4 U13361 ( .A1(n13056), .A2(n18906), .ZN(n10481) );
  NAND2_X1 U13362 ( .A1(n10481), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10439) );
  INV_X2 U13363 ( .A(n10505), .ZN(n10511) );
  AOI22_X1 U13364 ( .A1(n10511), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10438) );
  AND3_X1 U13365 ( .A1(n13054), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10436), 
        .ZN(n10440) );
  INV_X1 U13366 ( .A(n14822), .ZN(n10468) );
  NAND2_X1 U13367 ( .A1(n10468), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10441) );
  AND2_X1 U13368 ( .A1(n10442), .A2(n10441), .ZN(n10443) );
  NAND2_X1 U13369 ( .A1(n10444), .A2(n10443), .ZN(n11934) );
  NAND2_X1 U13370 ( .A1(n10446), .A2(n10445), .ZN(n13043) );
  INV_X1 U13371 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18924) );
  NAND2_X1 U13372 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10448) );
  AND2_X1 U13373 ( .A1(n14822), .A2(n10448), .ZN(n10449) );
  OAI211_X1 U13374 ( .C1(n10505), .C2(n18924), .A(n10450), .B(n10449), .ZN(
        n10451) );
  AOI21_X1 U13375 ( .B1(n10481), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10451), .ZN(
        n10453) );
  NAND2_X1 U13376 ( .A1(n10479), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10452) );
  OAI211_X1 U13377 ( .C1(n10454), .C2(n18906), .A(n10453), .B(n10452), .ZN(
        n11933) );
  INV_X1 U13378 ( .A(n10455), .ZN(n10456) );
  NAND2_X2 U13379 ( .A1(n10458), .A2(n10457), .ZN(n11962) );
  NAND2_X1 U13380 ( .A1(n10467), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10460) );
  AOI21_X1 U13381 ( .B1(n18906), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10459) );
  INV_X1 U13382 ( .A(n11953), .ZN(n10464) );
  NAND2_X1 U13383 ( .A1(n10479), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10463) );
  NAND2_X1 U13384 ( .A1(n10481), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13385 ( .A1(n10511), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10461) );
  NAND2_X1 U13386 ( .A1(n11962), .A2(n10464), .ZN(n10465) );
  NAND2_X1 U13387 ( .A1(n10466), .A2(n10465), .ZN(n10478) );
  NAND2_X1 U13388 ( .A1(n10467), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13389 ( .A1(n10468), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10469) );
  NAND2_X1 U13390 ( .A1(n9811), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10473) );
  NAND2_X1 U13391 ( .A1(n10481), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13392 ( .A1(n10511), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10471) );
  XNOR2_X2 U13393 ( .A(n10476), .B(n10474), .ZN(n11957) );
  INV_X1 U13394 ( .A(n10474), .ZN(n10475) );
  NOR2_X1 U13395 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  NAND2_X1 U13396 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10485) );
  NAND2_X1 U13397 ( .A1(n10482), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13398 ( .A1(n12663), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10483) );
  NAND3_X1 U13399 ( .A1(n10485), .A2(n10484), .A3(n10483), .ZN(n13506) );
  NAND2_X1 U13400 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10489) );
  NAND2_X1 U13401 ( .A1(n10482), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13402 ( .A1(n12663), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10487) );
  NAND3_X1 U13403 ( .A1(n10489), .A2(n10488), .A3(n10487), .ZN(n13620) );
  INV_X1 U13404 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U13405 ( .A1(n12663), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10491) );
  NAND2_X1 U13406 ( .A1(n10482), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10490) );
  OAI211_X1 U13407 ( .C1(n10498), .C2(n15542), .A(n10491), .B(n10490), .ZN(
        n13610) );
  NAND2_X1 U13408 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10494) );
  NAND2_X1 U13409 ( .A1(n10482), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13410 ( .A1(n12663), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10492) );
  NAND2_X1 U13411 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10497) );
  NAND2_X1 U13412 ( .A1(n10482), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13413 ( .A1(n12663), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10495) );
  NAND3_X1 U13414 ( .A1(n10497), .A2(n10496), .A3(n10495), .ZN(n13577) );
  INV_X1 U13415 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13416 ( .A1(n12663), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10499) );
  OAI21_X1 U13417 ( .B1(n10486), .B2(n10887), .A(n10499), .ZN(n10500) );
  AOI21_X1 U13418 ( .B1(n10480), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10500), .ZN(n13687) );
  NAND2_X1 U13419 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10503) );
  NAND2_X1 U13420 ( .A1(n10482), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13421 ( .A1(n10511), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10501) );
  NAND3_X1 U13422 ( .A1(n10503), .A2(n10502), .A3(n10501), .ZN(n13781) );
  INV_X1 U13423 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10504) );
  OAI22_X1 U13424 ( .A1(n10505), .A2(n10504), .B1(n19855), .B2(n16230), .ZN(
        n10507) );
  INV_X1 U13425 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15456) );
  NOR2_X1 U13426 ( .A1(n10498), .A2(n15456), .ZN(n10506) );
  AOI211_X1 U13427 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n10482), .A(n10507), .B(
        n10506), .ZN(n13912) );
  NAND2_X1 U13428 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10510) );
  NAND2_X1 U13429 ( .A1(n10482), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13430 ( .A1(n10511), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10508) );
  NAND3_X1 U13431 ( .A1(n10510), .A2(n10509), .A3(n10508), .ZN(n13924) );
  INV_X1 U13432 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U13433 ( .A1(n10511), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10512) );
  OAI21_X1 U13434 ( .B1(n10486), .B2(n10888), .A(n10512), .ZN(n10513) );
  AOI21_X1 U13435 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n10480), .A(
        n10513), .ZN(n14054) );
  INV_X1 U13436 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16321) );
  AOI22_X1 U13437 ( .A1(n12663), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10515) );
  NAND2_X1 U13438 ( .A1(n10482), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10514) );
  OAI211_X1 U13439 ( .C1(n10498), .C2(n16321), .A(n10515), .B(n10514), .ZN(
        n14077) );
  NAND2_X1 U13440 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10518) );
  NAND2_X1 U13441 ( .A1(n10482), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13442 ( .A1(n12663), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10516) );
  NAND2_X1 U13443 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10521) );
  NAND2_X1 U13444 ( .A1(n10482), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13445 ( .A1(n12663), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10519) );
  NAND3_X1 U13446 ( .A1(n10521), .A2(n10520), .A3(n10519), .ZN(n14994) );
  NAND2_X1 U13447 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10524) );
  NAND2_X1 U13448 ( .A1(n10482), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13449 ( .A1(n12663), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10522) );
  NAND2_X1 U13450 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10527) );
  NAND2_X1 U13451 ( .A1(n10482), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13452 ( .A1(n12663), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10525) );
  NAND2_X1 U13453 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10530) );
  NAND2_X1 U13454 ( .A1(n10482), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13455 ( .A1(n12663), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10528) );
  NAND3_X1 U13456 ( .A1(n10530), .A2(n10529), .A3(n10528), .ZN(n14976) );
  NAND2_X1 U13457 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10533) );
  NAND2_X1 U13458 ( .A1(n10482), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13459 ( .A1(n12663), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10531) );
  NAND3_X1 U13460 ( .A1(n10533), .A2(n10532), .A3(n10531), .ZN(n14966) );
  NAND2_X1 U13461 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10536) );
  NAND2_X1 U13462 ( .A1(n10482), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13463 ( .A1(n12663), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10534) );
  NAND2_X1 U13464 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10539) );
  NAND2_X1 U13465 ( .A1(n10482), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13466 ( .A1(n12663), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10537) );
  NAND2_X1 U13467 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10542) );
  NAND2_X1 U13468 ( .A1(n10482), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13469 ( .A1(n12663), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10540) );
  NAND2_X1 U13470 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10545) );
  NAND2_X1 U13471 ( .A1(n10482), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10544) );
  AOI22_X1 U13472 ( .A1(n12663), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10543) );
  NAND3_X1 U13473 ( .A1(n10545), .A2(n10544), .A3(n10543), .ZN(n14843) );
  NAND2_X1 U13474 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10548) );
  NAND2_X1 U13475 ( .A1(n10482), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13476 ( .A1(n12663), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10546) );
  AND3_X1 U13477 ( .A1(n10548), .A2(n10547), .A3(n10546), .ZN(n14927) );
  NAND2_X1 U13478 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10551) );
  NAND2_X1 U13479 ( .A1(n10482), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13480 ( .A1(n12663), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10549) );
  NAND2_X1 U13481 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10554) );
  NAND2_X1 U13482 ( .A1(n10482), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U13483 ( .A1(n12663), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10552) );
  NAND3_X1 U13484 ( .A1(n10554), .A2(n10553), .A3(n10552), .ZN(n14908) );
  NAND2_X1 U13485 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10557) );
  NAND2_X1 U13486 ( .A1(n10482), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13487 ( .A1(n12663), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10555) );
  NAND3_X1 U13488 ( .A1(n10557), .A2(n10556), .A3(n10555), .ZN(n14829) );
  NAND2_X1 U13489 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10560) );
  NAND2_X1 U13490 ( .A1(n10482), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13491 ( .A1(n12663), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10558) );
  AND3_X1 U13492 ( .A1(n10560), .A2(n10559), .A3(n10558), .ZN(n14894) );
  NAND2_X1 U13493 ( .A1(n10480), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10563) );
  NAND2_X1 U13494 ( .A1(n10482), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U13495 ( .A1(n12663), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10561) );
  NAND3_X1 U13496 ( .A1(n10563), .A2(n10562), .A3(n10561), .ZN(n10564) );
  NAND2_X1 U13497 ( .A1(n14897), .A2(n10564), .ZN(n12667) );
  INV_X1 U13498 ( .A(n14897), .ZN(n10566) );
  INV_X1 U13499 ( .A(n10564), .ZN(n10565) );
  NAND2_X1 U13500 ( .A1(n10566), .A2(n10565), .ZN(n10567) );
  NAND2_X1 U13501 ( .A1(n12667), .A2(n10567), .ZN(n15079) );
  XNOR2_X1 U13502 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12255) );
  NAND2_X1 U13503 ( .A1(n12255), .A2(n10582), .ZN(n10569) );
  NAND2_X1 U13504 ( .A1(n19978), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10568) );
  NAND2_X1 U13505 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19968), .ZN(
        n10570) );
  NAND2_X1 U13506 ( .A1(n10579), .A2(n10570), .ZN(n10572) );
  NAND2_X1 U13507 ( .A1(n10202), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10571) );
  MUX2_X1 U13508 ( .A(n19960), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10577) );
  INV_X1 U13509 ( .A(n10577), .ZN(n10573) );
  INV_X1 U13510 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16334) );
  NOR2_X1 U13511 ( .A1(n16334), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10575) );
  NAND3_X1 U13512 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10576), .A3(
        n13228), .ZN(n10876) );
  XNOR2_X1 U13513 ( .A(n10578), .B(n10577), .ZN(n10880) );
  INV_X1 U13514 ( .A(n10579), .ZN(n10581) );
  MUX2_X1 U13515 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n19968), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10580) );
  XNOR2_X1 U13516 ( .A(n10581), .B(n10580), .ZN(n12264) );
  NAND2_X1 U13517 ( .A1(n12270), .A2(n12264), .ZN(n12601) );
  INV_X1 U13518 ( .A(n10582), .ZN(n12257) );
  XNOR2_X1 U13519 ( .A(n12255), .B(n12257), .ZN(n12258) );
  INV_X1 U13520 ( .A(n12258), .ZN(n10583) );
  NOR2_X1 U13521 ( .A1(n12601), .A2(n10583), .ZN(n10584) );
  OR2_X1 U13522 ( .A1(n12612), .A2(n10584), .ZN(n16338) );
  NAND2_X1 U13523 ( .A1(n19855), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19854) );
  NAND2_X1 U13524 ( .A1(n16363), .A2(n19259), .ZN(n10898) );
  NAND2_X1 U13525 ( .A1(n13231), .A2(n10898), .ZN(n16337) );
  INV_X1 U13526 ( .A(n16337), .ZN(n10585) );
  AND2_X1 U13527 ( .A1(n18907), .A2(n10436), .ZN(n10895) );
  NAND2_X1 U13528 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n16356) );
  NAND2_X1 U13529 ( .A1(n19457), .A2(n16356), .ZN(n10899) );
  INV_X1 U13530 ( .A(n10899), .ZN(n10586) );
  NOR2_X1 U13531 ( .A1(n19292), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10591) );
  INV_X2 U13532 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19979) );
  AND2_X2 U13533 ( .A1(n19264), .A2(n19979), .ZN(n10665) );
  AOI22_X1 U13534 ( .A1(n13072), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10590) );
  NAND2_X1 U13535 ( .A1(n9798), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U13536 ( .A1(n10590), .A2(n10589), .ZN(n15339) );
  NAND2_X1 U13537 ( .A1(n9798), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13538 ( .A1(n13072), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13539 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13540 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10596) );
  AND2_X2 U13541 ( .A1(n10593), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10751) );
  AND2_X2 U13542 ( .A1(n10593), .A2(n16325), .ZN(n11989) );
  AOI22_X1 U13543 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10751), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13544 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12031), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10594) );
  NAND4_X1 U13545 ( .A1(n10597), .A2(n10596), .A3(n10595), .A4(n10594), .ZN(
        n10604) );
  AOI22_X1 U13546 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10634), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10602) );
  AND2_X1 U13547 ( .A1(n12243), .A2(n16325), .ZN(n10693) );
  AOI22_X1 U13548 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10692), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10601) );
  INV_X1 U13549 ( .A(n10598), .ZN(n15585) );
  NOR2_X1 U13550 ( .A1(n15585), .A2(n16325), .ZN(n12599) );
  AOI22_X1 U13551 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10600) );
  AND2_X2 U13552 ( .A1(n9808), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10635) );
  AOI22_X1 U13553 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10599) );
  NAND4_X1 U13554 ( .A1(n10602), .A2(n10601), .A3(n10600), .A4(n10599), .ZN(
        n10603) );
  NAND2_X1 U13555 ( .A1(n10825), .A2(n13926), .ZN(n10605) );
  NAND2_X1 U13556 ( .A1(n10625), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10611) );
  INV_X1 U13557 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19227) );
  NAND2_X1 U13558 ( .A1(n19264), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10608) );
  OAI211_X1 U13559 ( .C1(n19292), .C2(n19227), .A(n10608), .B(n19979), .ZN(
        n10609) );
  INV_X1 U13560 ( .A(n10609), .ZN(n10610) );
  AOI22_X1 U13561 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13562 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13563 ( .A1(n10751), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10613) );
  AOI22_X1 U13564 ( .A1(n12031), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10612) );
  NAND4_X1 U13565 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10622) );
  AOI22_X1 U13566 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13567 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13568 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13569 ( .A1(n10635), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10617) );
  NAND4_X1 U13570 ( .A1(n10620), .A2(n10619), .A3(n10618), .A4(n10617), .ZN(
        n10621) );
  INV_X1 U13571 ( .A(n12624), .ZN(n12413) );
  NAND2_X1 U13572 ( .A1(n10623), .A2(n10665), .ZN(n10660) );
  MUX2_X1 U13573 ( .A(n19292), .B(n19987), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10624) );
  INV_X1 U13574 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15580) );
  AOI22_X1 U13575 ( .A1(n10591), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10665), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10627) );
  INV_X1 U13576 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19878) );
  NAND2_X1 U13577 ( .A1(n10625), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10626) );
  NAND2_X1 U13578 ( .A1(n10627), .A2(n10626), .ZN(n10645) );
  INV_X1 U13579 ( .A(n10645), .ZN(n10628) );
  NAND2_X1 U13580 ( .A1(n10409), .A2(n19292), .ZN(n10629) );
  MUX2_X1 U13581 ( .A(n10629), .B(n19978), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10644) );
  AOI22_X1 U13582 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10670), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13583 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13584 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10648), .B1(
        n10751), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10631) );
  AOI22_X1 U13585 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11989), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10630) );
  NAND4_X1 U13586 ( .A1(n10633), .A2(n10632), .A3(n10631), .A4(n10630), .ZN(
        n10642) );
  AOI22_X1 U13587 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10693), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10640) );
  AOI22_X1 U13588 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10634), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10639) );
  AOI22_X1 U13589 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13590 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10635), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10637) );
  NAND4_X1 U13591 ( .A1(n10640), .A2(n10639), .A3(n10638), .A4(n10637), .ZN(
        n10641) );
  NAND2_X1 U13592 ( .A1(n10825), .A2(n12622), .ZN(n10643) );
  AND2_X1 U13593 ( .A1(n10644), .A2(n10643), .ZN(n13274) );
  NAND2_X1 U13594 ( .A1(n13275), .A2(n13274), .ZN(n10662) );
  AOI22_X1 U13595 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13596 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13597 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13598 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11989), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10649) );
  NAND4_X1 U13599 ( .A1(n10652), .A2(n10651), .A3(n10650), .A4(n10649), .ZN(
        n10658) );
  AOI22_X1 U13600 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13601 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13602 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13603 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10653) );
  NAND4_X1 U13604 ( .A1(n10656), .A2(n10655), .A3(n10654), .A4(n10653), .ZN(
        n10657) );
  INV_X1 U13605 ( .A(n12620), .ZN(n10661) );
  NAND2_X1 U13606 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10659) );
  OAI211_X1 U13607 ( .C1(n10661), .C2(n10841), .A(n10660), .B(n10659), .ZN(
        n10663) );
  AND3_X1 U13608 ( .A1(n10662), .A2(n9851), .A3(n10663), .ZN(n10664) );
  AOI22_X1 U13609 ( .A1(n13072), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10665), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U13610 ( .A1(n9798), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10667) );
  NAND2_X1 U13611 ( .A1(n10668), .A2(n10667), .ZN(n13313) );
  NOR2_X1 U13612 ( .A1(n13314), .A2(n13313), .ZN(n13315) );
  NAND2_X1 U13613 ( .A1(n9798), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13614 ( .A1(n10665), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10686) );
  AOI22_X1 U13615 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13616 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13617 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11989), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10672) );
  NAND4_X1 U13618 ( .A1(n10675), .A2(n10674), .A3(n10673), .A4(n10672), .ZN(
        n10682) );
  AOI22_X1 U13619 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13620 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13621 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13622 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10677) );
  NAND4_X1 U13623 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10677), .ZN(
        n10681) );
  NOR2_X1 U13624 ( .A1(n10682), .A2(n10681), .ZN(n12343) );
  INV_X1 U13625 ( .A(n12343), .ZN(n10683) );
  NAND2_X1 U13626 ( .A1(n10825), .A2(n10683), .ZN(n10685) );
  NAND2_X1 U13627 ( .A1(n13072), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10684) );
  NAND4_X1 U13628 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n13977) );
  NAND2_X1 U13629 ( .A1(n13976), .A2(n13977), .ZN(n13978) );
  NAND2_X1 U13630 ( .A1(n9798), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13631 ( .A1(n13072), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10665), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13632 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13633 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13634 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13635 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11989), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10688) );
  NAND4_X1 U13636 ( .A1(n10691), .A2(n10690), .A3(n10689), .A4(n10688), .ZN(
        n10699) );
  AOI22_X1 U13637 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13638 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U13639 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13640 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10694) );
  NAND4_X1 U13641 ( .A1(n10697), .A2(n10696), .A3(n10695), .A4(n10694), .ZN(
        n10698) );
  NAND2_X1 U13642 ( .A1(n10825), .A2(n12634), .ZN(n10700) );
  AOI22_X1 U13643 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13644 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10705) );
  AOI22_X1 U13645 ( .A1(n10751), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10704) );
  AOI22_X1 U13646 ( .A1(n12031), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10703) );
  NAND4_X1 U13647 ( .A1(n10706), .A2(n10705), .A3(n10704), .A4(n10703), .ZN(
        n10712) );
  AOI22_X1 U13648 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13649 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U13650 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13651 ( .A1(n10635), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10707) );
  NAND4_X1 U13652 ( .A1(n10710), .A2(n10709), .A3(n10708), .A4(n10707), .ZN(
        n10711) );
  INV_X1 U13653 ( .A(n12396), .ZN(n10713) );
  AOI22_X1 U13654 ( .A1(n9798), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n10825), .B2(
        n10713), .ZN(n10715) );
  AOI22_X1 U13655 ( .A1(n13072), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10665), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10714) );
  NAND2_X1 U13656 ( .A1(n10715), .A2(n10714), .ZN(n14185) );
  AOI22_X1 U13657 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13658 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13659 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10671), .B1(
        n10751), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13660 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11989), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10716) );
  NAND4_X1 U13661 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n10725) );
  AOI22_X1 U13662 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10693), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13663 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10634), .B1(
        n10635), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13664 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13665 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10676), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10720) );
  NAND4_X1 U13666 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n10720), .ZN(
        n10724) );
  NAND2_X1 U13667 ( .A1(n10825), .A2(n12453), .ZN(n15534) );
  AOI22_X1 U13668 ( .A1(n13072), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10665), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10727) );
  NAND2_X1 U13669 ( .A1(n9798), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10726) );
  NAND2_X1 U13670 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10731) );
  NAND2_X1 U13671 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10730) );
  NAND2_X1 U13672 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10729) );
  NAND2_X1 U13673 ( .A1(n10648), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10728) );
  NAND2_X1 U13674 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10735) );
  NAND2_X1 U13675 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10734) );
  NAND2_X1 U13676 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10733) );
  NAND2_X1 U13677 ( .A1(n10692), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10732) );
  NAND2_X1 U13678 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10739) );
  NAND2_X1 U13679 ( .A1(n10693), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10738) );
  NAND2_X1 U13680 ( .A1(n10635), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10737) );
  NAND2_X1 U13681 ( .A1(n12004), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10736) );
  NAND2_X1 U13682 ( .A1(n10751), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10743) );
  NAND2_X1 U13683 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10742) );
  NAND2_X1 U13684 ( .A1(n12031), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10741) );
  NAND2_X1 U13685 ( .A1(n11989), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10740) );
  NAND4_X1 U13686 ( .A1(n10747), .A2(n10746), .A3(n10745), .A4(n10744), .ZN(
        n10884) );
  INV_X1 U13687 ( .A(n10884), .ZN(n12399) );
  NAND2_X1 U13688 ( .A1(n10825), .A2(n12571), .ZN(n10748) );
  AOI22_X1 U13689 ( .A1(n13072), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10665), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U13690 ( .A1(n9798), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10749) );
  NAND2_X1 U13691 ( .A1(n10750), .A2(n10749), .ZN(n13960) );
  NAND2_X1 U13692 ( .A1(n9798), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13693 ( .A1(n13072), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10665), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13694 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13695 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U13696 ( .A1(n12031), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U13697 ( .A1(n10751), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10752) );
  NAND4_X1 U13698 ( .A1(n10755), .A2(n10754), .A3(n10753), .A4(n10752), .ZN(
        n10761) );
  AOI22_X1 U13699 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13700 ( .A1(n10635), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13701 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10757) );
  AOI22_X1 U13702 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10756) );
  NAND4_X1 U13703 ( .A1(n10759), .A2(n10758), .A3(n10757), .A4(n10756), .ZN(
        n10760) );
  NAND2_X1 U13704 ( .A1(n10825), .A2(n13581), .ZN(n10762) );
  AOI22_X1 U13705 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13706 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U13707 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13708 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11989), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10765) );
  NAND4_X1 U13709 ( .A1(n10768), .A2(n10767), .A3(n10766), .A4(n10765), .ZN(
        n10774) );
  AOI22_X1 U13710 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13711 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13712 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13713 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10769) );
  NAND4_X1 U13714 ( .A1(n10772), .A2(n10771), .A3(n10770), .A4(n10769), .ZN(
        n10773) );
  NOR2_X1 U13715 ( .A1(n10774), .A2(n10773), .ZN(n13684) );
  AOI22_X1 U13716 ( .A1(n13072), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10665), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13717 ( .A1(n9798), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10775) );
  OAI211_X1 U13718 ( .C1(n13684), .C2(n10841), .A(n10776), .B(n10775), .ZN(
        n15490) );
  NAND2_X1 U13719 ( .A1(n9798), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13720 ( .A1(n13072), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13721 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10670), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U13722 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U13723 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n11989), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13724 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10777) );
  NAND4_X1 U13725 ( .A1(n10780), .A2(n10779), .A3(n10778), .A4(n10777), .ZN(
        n10786) );
  AOI22_X1 U13726 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10635), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10784) );
  AOI22_X1 U13727 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13728 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U13729 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10693), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10781) );
  NAND4_X1 U13730 ( .A1(n10784), .A2(n10783), .A3(n10782), .A4(n10781), .ZN(
        n10785) );
  NAND2_X1 U13731 ( .A1(n10825), .A2(n9834), .ZN(n10787) );
  AOI22_X1 U13732 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13733 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13734 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13735 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11989), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10790) );
  NAND4_X1 U13736 ( .A1(n10793), .A2(n10792), .A3(n10791), .A4(n10790), .ZN(
        n10799) );
  AOI22_X1 U13737 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U13738 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U13739 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U13740 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10794) );
  NAND4_X1 U13741 ( .A1(n10797), .A2(n10796), .A3(n10795), .A4(n10794), .ZN(
        n10798) );
  INV_X1 U13742 ( .A(n13910), .ZN(n10802) );
  AOI22_X1 U13743 ( .A1(n13072), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10801) );
  NAND2_X1 U13744 ( .A1(n9798), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10800) );
  OAI211_X1 U13745 ( .C1(n10802), .C2(n10841), .A(n10801), .B(n10800), .ZN(
        n15451) );
  AOI22_X1 U13746 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13747 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13748 ( .A1(n10751), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13749 ( .A1(n12031), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10803) );
  NAND4_X1 U13750 ( .A1(n10806), .A2(n10805), .A3(n10804), .A4(n10803), .ZN(
        n10812) );
  AOI22_X1 U13751 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13752 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13753 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13754 ( .A1(n10635), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10807) );
  NAND4_X1 U13755 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n10811) );
  NOR2_X1 U13756 ( .A1(n10812), .A2(n10811), .ZN(n14055) );
  AOI22_X1 U13757 ( .A1(n13072), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U13758 ( .A1(n9798), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10813) );
  OAI211_X1 U13759 ( .C1(n14055), .C2(n10841), .A(n10814), .B(n10813), .ZN(
        n15418) );
  NAND2_X1 U13760 ( .A1(n9798), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13761 ( .A1(n13072), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13762 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13763 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13764 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12031), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U13765 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10815) );
  NAND4_X1 U13766 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        n10824) );
  AOI22_X1 U13767 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10692), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13768 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13769 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13770 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10634), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10819) );
  NAND4_X1 U13771 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10823) );
  NOR2_X1 U13772 ( .A1(n10824), .A2(n10823), .ZN(n11986) );
  INV_X1 U13773 ( .A(n11986), .ZN(n14080) );
  NAND2_X1 U13774 ( .A1(n10825), .A2(n14080), .ZN(n10826) );
  AOI22_X1 U13775 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13776 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13777 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13778 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11989), .B1(
        n12031), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10829) );
  NAND4_X1 U13779 ( .A1(n10832), .A2(n10831), .A3(n10830), .A4(n10829), .ZN(
        n10838) );
  AOI22_X1 U13780 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13781 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13782 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13783 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10833) );
  NAND4_X1 U13784 ( .A1(n10836), .A2(n10835), .A3(n10834), .A4(n10833), .ZN(
        n10837) );
  NOR2_X1 U13785 ( .A1(n10838), .A2(n10837), .ZN(n14160) );
  AOI22_X1 U13786 ( .A1(n13072), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10840) );
  NAND2_X1 U13787 ( .A1(n9798), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10839) );
  OAI211_X1 U13788 ( .C1(n14160), .C2(n10841), .A(n10840), .B(n10839), .ZN(
        n15405) );
  NAND2_X1 U13789 ( .A1(n9798), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10843) );
  AOI22_X1 U13790 ( .A1(n13072), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10842) );
  AOI22_X1 U13791 ( .A1(n13072), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10845) );
  NAND2_X1 U13792 ( .A1(n9798), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10844) );
  NAND2_X1 U13793 ( .A1(n10845), .A2(n10844), .ZN(n14202) );
  NAND2_X1 U13794 ( .A1(n9798), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13795 ( .A1(n13072), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13796 ( .A1(n13072), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10849) );
  NAND2_X1 U13797 ( .A1(n9798), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10848) );
  NAND2_X1 U13798 ( .A1(n10849), .A2(n10848), .ZN(n15063) );
  AOI22_X1 U13799 ( .A1(n13072), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10851) );
  NAND2_X1 U13800 ( .A1(n9798), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10850) );
  NAND2_X1 U13801 ( .A1(n10851), .A2(n10850), .ZN(n15363) );
  AOI22_X1 U13802 ( .A1(n13072), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10853) );
  NAND2_X1 U13803 ( .A1(n9798), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U13804 ( .A1(n10853), .A2(n10852), .ZN(n15054) );
  NAND2_X1 U13805 ( .A1(n15053), .A2(n15054), .ZN(n15055) );
  NAND2_X1 U13806 ( .A1(n9798), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13807 ( .A1(n13072), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10854) );
  AND2_X1 U13808 ( .A1(n10855), .A2(n10854), .ZN(n15044) );
  NAND2_X1 U13809 ( .A1(n9798), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13810 ( .A1(n13072), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10856) );
  AND2_X1 U13811 ( .A1(n10857), .A2(n10856), .ZN(n14846) );
  INV_X1 U13812 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19923) );
  AOI22_X1 U13813 ( .A1(n13072), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10858) );
  OAI21_X1 U13814 ( .B1(n19923), .B2(n10666), .A(n10858), .ZN(n15033) );
  NAND2_X1 U13815 ( .A1(n9798), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10860) );
  AOI22_X1 U13816 ( .A1(n13072), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10859) );
  AND2_X1 U13817 ( .A1(n10860), .A2(n10859), .ZN(n15026) );
  NAND2_X1 U13818 ( .A1(n9798), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13819 ( .A1(n13072), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10861) );
  AND2_X1 U13820 ( .A1(n10862), .A2(n10861), .ZN(n15018) );
  AOI22_X1 U13821 ( .A1(n13072), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10864) );
  NAND2_X1 U13822 ( .A1(n9798), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10863) );
  NAND2_X1 U13823 ( .A1(n10864), .A2(n10863), .ZN(n14832) );
  INV_X1 U13824 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19931) );
  AOI22_X1 U13825 ( .A1(n13072), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10865) );
  OAI21_X1 U13826 ( .B1(n19931), .B2(n10666), .A(n10865), .ZN(n15004) );
  NAND2_X1 U13827 ( .A1(n9798), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13828 ( .A1(n13072), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n10665), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10866) );
  AND2_X1 U13829 ( .A1(n10867), .A2(n10866), .ZN(n10870) );
  INV_X1 U13830 ( .A(n10870), .ZN(n10868) );
  NAND2_X1 U13831 ( .A1(n10869), .A2(n10868), .ZN(n13075) );
  NAND2_X1 U13832 ( .A1(n15007), .A2(n10870), .ZN(n10871) );
  AND2_X1 U13833 ( .A1(n13446), .A2(n19259), .ZN(n16362) );
  INV_X1 U13834 ( .A(n16356), .ZN(n19869) );
  INV_X1 U13835 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18903) );
  INV_X1 U13836 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19877) );
  NOR2_X1 U13837 ( .A1(n18903), .A2(n19877), .ZN(n19870) );
  NOR2_X1 U13838 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19858) );
  NOR3_X1 U13839 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19870), .A3(n19858), 
        .ZN(n19863) );
  INV_X1 U13840 ( .A(n19863), .ZN(n10872) );
  NOR2_X1 U13841 ( .A1(n19869), .A2(n10872), .ZN(n13215) );
  INV_X1 U13842 ( .A(n13215), .ZN(n10873) );
  NOR2_X1 U13843 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n10873), .ZN(n16361) );
  AND2_X1 U13844 ( .A1(n16362), .A2(n16361), .ZN(n10874) );
  OAI22_X1 U13845 ( .A1(n15079), .A2(n19109), .B1(n14309), .B2(n19085), .ZN(
        n10875) );
  MUX2_X1 U13846 ( .A(n10876), .B(n12634), .S(n10436), .Z(n12611) );
  INV_X1 U13847 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10877) );
  MUX2_X1 U13848 ( .A(n12611), .B(n10877), .S(n12592), .Z(n12423) );
  MUX2_X1 U13849 ( .A(n12620), .B(n12264), .S(n13035), .Z(n12605) );
  INV_X1 U13850 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10878) );
  MUX2_X1 U13851 ( .A(n12605), .B(n10878), .S(n12592), .Z(n12412) );
  NOR2_X1 U13852 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n10879) );
  MUX2_X1 U13853 ( .A(n12622), .B(n10879), .S(n12592), .Z(n12415) );
  INV_X1 U13854 ( .A(n10880), .ZN(n10881) );
  MUX2_X1 U13855 ( .A(n12343), .B(n10881), .S(n13035), .Z(n12604) );
  NAND2_X1 U13856 ( .A1(n12423), .A2(n12422), .ZN(n12421) );
  MUX2_X1 U13857 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12396), .S(n19277), .Z(
        n12401) );
  INV_X1 U13858 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19062) );
  MUX2_X1 U13859 ( .A(n12453), .B(n19062), .S(n12592), .Z(n12457) );
  INV_X1 U13860 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10885) );
  MUX2_X1 U13861 ( .A(n10885), .B(n10884), .S(n19277), .Z(n12463) );
  NAND2_X1 U13862 ( .A1(n12592), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12468) );
  INV_X1 U13863 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U13864 ( .A1(n12592), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12494) );
  INV_X1 U13865 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10889) );
  NOR2_X1 U13866 ( .A1(n19277), .A2(n10889), .ZN(n12509) );
  NAND2_X1 U13867 ( .A1(n12592), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12506) );
  NAND2_X1 U13868 ( .A1(n12592), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12516) );
  NOR2_X1 U13869 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n10890) );
  NOR2_X1 U13870 ( .A1(n19277), .A2(n10890), .ZN(n10891) );
  INV_X1 U13871 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14961) );
  NAND2_X1 U13872 ( .A1(n12592), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12544) );
  INV_X1 U13873 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10892) );
  NOR2_X1 U13874 ( .A1(n19277), .A2(n10892), .ZN(n12549) );
  INV_X1 U13875 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14930) );
  NAND2_X1 U13876 ( .A1(n12592), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12576) );
  INV_X1 U13877 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10893) );
  NOR2_X1 U13878 ( .A1(n19277), .A2(n10893), .ZN(n12572) );
  NAND2_X1 U13879 ( .A1(n12592), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U13880 ( .A1(n12592), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10894) );
  XNOR2_X1 U13881 ( .A(n12593), .B(n10894), .ZN(n12588) );
  INV_X1 U13882 ( .A(n10895), .ZN(n10897) );
  NAND2_X1 U13883 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n10899), .ZN(n10896) );
  OR2_X1 U13884 ( .A1(n13529), .A2(n16361), .ZN(n16087) );
  INV_X1 U13885 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16088) );
  NAND3_X1 U13886 ( .A1(n13445), .A2(n10899), .A3(n16088), .ZN(n10900) );
  AOI22_X1 U13887 ( .A1(n12588), .A2(n19039), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n19107), .ZN(n10906) );
  NOR2_X1 U13888 ( .A1(n19979), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19849) );
  INV_X1 U13889 ( .A(n19849), .ZN(n10901) );
  NOR2_X1 U13890 ( .A1(n19854), .A2(n10901), .ZN(n16358) );
  NAND2_X1 U13891 ( .A1(n19855), .A2(n19979), .ZN(n15611) );
  NOR2_X1 U13892 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15611), .ZN(n10902) );
  INV_X2 U13893 ( .A(n19235), .ZN(n19041) );
  NAND2_X1 U13894 ( .A1(n19041), .A2(n19048), .ZN(n10903) );
  OR2_X1 U13895 ( .A1(n16358), .A2(n10903), .ZN(n10904) );
  NAND2_X1 U13896 ( .A1(n19049), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19072) );
  INV_X2 U13897 ( .A(n19072), .ZN(n19114) );
  AOI22_X1 U13898 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n19102), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19114), .ZN(n10905) );
  NAND2_X1 U13899 ( .A1(n10906), .A2(n10905), .ZN(n10907) );
  NAND2_X1 U13900 ( .A1(n10909), .A2(n10908), .ZN(P2_U2825) );
  INV_X1 U13901 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10910) );
  AND2_X2 U13902 ( .A1(n10921), .A2(n10919), .ZN(n10972) );
  AOI22_X1 U13903 ( .A1(n11091), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10916) );
  AND2_X4 U13904 ( .A1(n10918), .A2(n10922), .ZN(n11730) );
  AOI22_X1 U13905 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11141), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10915) );
  AND2_X4 U13906 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13393) );
  AOI22_X1 U13907 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11122), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10914) );
  NOR2_X4 U13908 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10920) );
  AND2_X2 U13909 ( .A1(n13737), .A2(n10920), .ZN(n10991) );
  AOI22_X1 U13910 ( .A1(n10991), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10913) );
  NAND4_X1 U13911 ( .A1(n10916), .A2(n10915), .A3(n10914), .A4(n10913), .ZN(
        n10928) );
  AOI22_X1 U13913 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10926) );
  AND2_X2 U13914 ( .A1(n10918), .A2(n10919), .ZN(n11683) );
  AOI22_X1 U13915 ( .A1(n11683), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10925) );
  AND2_X2 U13916 ( .A1(n13737), .A2(n13393), .ZN(n10961) );
  AOI22_X1 U13917 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10924) );
  AND2_X4 U13918 ( .A1(n10921), .A2(n10922), .ZN(n11701) );
  AOI22_X1 U13919 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11127), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10923) );
  NAND4_X1 U13920 ( .A1(n10926), .A2(n10925), .A3(n10924), .A4(n10923), .ZN(
        n10927) );
  INV_X1 U13921 ( .A(n11034), .ZN(n11043) );
  AOI22_X1 U13922 ( .A1(n11091), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13923 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10973), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13925 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U13926 ( .A1(n10991), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11127), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13927 ( .A1(n11683), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13928 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11141), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U13929 ( .A1(n11092), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13930 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13932 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13933 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11683), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13934 ( .A1(n11091), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U13935 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U13936 ( .A1(n10991), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U13937 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10945) );
  AOI22_X1 U13938 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11141), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U13939 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11127), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10943) );
  NAND2_X1 U13940 ( .A1(n10262), .A2(n10261), .ZN(n11038) );
  INV_X1 U13941 ( .A(n11038), .ZN(n20190) );
  AOI22_X1 U13942 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U13943 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11127), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10947) );
  AOI22_X1 U13944 ( .A1(n10991), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U13945 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11683), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U13946 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U13947 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U13948 ( .A1(n11091), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10953) );
  NAND2_X2 U13949 ( .A1(n10957), .A2(n10956), .ZN(n11032) );
  NAND2_X1 U13950 ( .A1(n11031), .A2(n11032), .ZN(n10958) );
  NAND2_X1 U13951 ( .A1(n20190), .A2(n10958), .ZN(n10959) );
  NAND2_X1 U13952 ( .A1(n10960), .A2(n10959), .ZN(n10986) );
  AOI22_X1 U13953 ( .A1(n11091), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11115), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U13954 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U13955 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11127), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U13956 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10962) );
  NAND4_X1 U13957 ( .A1(n10965), .A2(n10964), .A3(n10963), .A4(n10962), .ZN(
        n10971) );
  AOI22_X1 U13958 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U13959 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11683), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U13960 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U13961 ( .A1(n10991), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11730), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10966) );
  NAND4_X1 U13962 ( .A1(n10969), .A2(n10968), .A3(n10967), .A4(n10966), .ZN(
        n10970) );
  BUF_X4 U13963 ( .A(n11701), .Z(n11733) );
  AOI22_X1 U13964 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U13965 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U13966 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11683), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U13967 ( .A1(n11091), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11092), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U13968 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10975) );
  AOI21_X1 U13969 ( .B1(n11141), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n10979), .ZN(n10982) );
  AOI22_X1 U13970 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11127), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U13971 ( .A1(n10991), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10980) );
  NAND3_X2 U13972 ( .A1(n10984), .A2(n10983), .A3(n10260), .ZN(n11231) );
  NAND2_X1 U13973 ( .A1(n11231), .A2(n11034), .ZN(n11050) );
  NAND2_X1 U13974 ( .A1(n11050), .A2(n11040), .ZN(n10985) );
  NAND3_X1 U13975 ( .A1(n10986), .A2(n11068), .A3(n10985), .ZN(n11047) );
  NAND2_X1 U13976 ( .A1(n11091), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10990) );
  NAND2_X1 U13977 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10989) );
  NAND2_X1 U13978 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10988) );
  NAND2_X1 U13979 ( .A1(n11092), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10987) );
  BUF_X8 U13980 ( .A(n10991), .Z(n11657) );
  NAND2_X1 U13981 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10996) );
  NAND2_X1 U13982 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10995) );
  NAND2_X1 U13983 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10994) );
  NAND2_X1 U13984 ( .A1(n10992), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10993) );
  NAND2_X1 U13985 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11000) );
  NAND2_X1 U13986 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10999) );
  NAND2_X1 U13987 ( .A1(n11683), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10998) );
  NAND2_X1 U13988 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10997) );
  NAND2_X1 U13989 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11004) );
  NAND2_X1 U13990 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11003) );
  NAND2_X1 U13991 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11002) );
  NAND2_X1 U13992 ( .A1(n11437), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11001) );
  NAND4_X4 U13993 ( .A1(n11008), .A2(n11007), .A3(n11006), .A4(n11005), .ZN(
        n13557) );
  NAND2_X1 U13994 ( .A1(n11912), .A2(n20170), .ZN(n11009) );
  NAND2_X1 U13996 ( .A1(n11091), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11013) );
  NAND2_X1 U13997 ( .A1(n11115), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11012) );
  NAND2_X1 U13998 ( .A1(n10972), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11011) );
  NAND2_X1 U13999 ( .A1(n11092), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11010) );
  NAND2_X1 U14000 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U14001 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11016) );
  NAND2_X1 U14002 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11015) );
  NAND2_X1 U14003 ( .A1(n10992), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11014) );
  NAND2_X1 U14004 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11021) );
  NAND2_X1 U14005 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11020) );
  NAND2_X1 U14006 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11019) );
  NAND2_X1 U14007 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11018) );
  NAND2_X1 U14008 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11025) );
  NAND2_X1 U14009 ( .A1(n11122), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11024) );
  NAND2_X1 U14010 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11023) );
  INV_X1 U14011 ( .A(n13100), .ZN(n11030) );
  INV_X1 U14012 ( .A(n11031), .ZN(n11039) );
  NAND2_X1 U14013 ( .A1(n11039), .A2(n11032), .ZN(n11033) );
  NOR2_X1 U14014 ( .A1(n11031), .A2(n11034), .ZN(n11035) );
  NAND2_X1 U14015 ( .A1(n9809), .A2(n13557), .ZN(n13262) );
  INV_X1 U14016 ( .A(n13262), .ZN(n11037) );
  XNOR2_X1 U14017 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n13345) );
  NOR2_X2 U14018 ( .A1(n13540), .A2(n11762), .ZN(n13397) );
  INV_X1 U14019 ( .A(n13746), .ZN(n11042) );
  NAND2_X2 U14020 ( .A1(n20183), .A2(n13557), .ZN(n20819) );
  NAND2_X1 U14021 ( .A1(n13540), .A2(n13557), .ZN(n11044) );
  INV_X1 U14022 ( .A(n11045), .ZN(n11046) );
  NAND2_X1 U14023 ( .A1(n11048), .A2(n9812), .ZN(n11057) );
  AND2_X1 U14024 ( .A1(n11049), .A2(n20202), .ZN(n11054) );
  INV_X1 U14025 ( .A(n11052), .ZN(n11053) );
  NAND3_X1 U14026 ( .A1(n11058), .A2(n11057), .A3(n11056), .ZN(n11059) );
  NAND2_X1 U14027 ( .A1(n11059), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11060) );
  NAND2_X2 U14028 ( .A1(n11076), .A2(n11060), .ZN(n11080) );
  NAND2_X1 U14029 ( .A1(n11080), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11063) );
  NAND2_X1 U14030 ( .A1(n20798), .A2(n20169), .ZN(n11917) );
  NAND2_X1 U14031 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11083) );
  OAI21_X1 U14032 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11083), .ZN(n20494) );
  NAND2_X1 U14033 ( .A1(n20735), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11077) );
  OAI21_X1 U14034 ( .B1(n11917), .B2(n20494), .A(n11077), .ZN(n11061) );
  INV_X1 U14035 ( .A(n11061), .ZN(n11062) );
  XNOR2_X2 U14036 ( .A(n11064), .B(n11076), .ZN(n20294) );
  INV_X1 U14037 ( .A(n20735), .ZN(n15729) );
  MUX2_X1 U14038 ( .A(n15729), .B(n11917), .S(n20610), .Z(n11065) );
  OAI21_X1 U14039 ( .B1(n15708), .B2(n11068), .A(n11048), .ZN(n11075) );
  NAND2_X1 U14040 ( .A1(n13397), .A2(n20215), .ZN(n13555) );
  NAND2_X1 U14041 ( .A1(n11052), .A2(n11838), .ZN(n11070) );
  INV_X1 U14042 ( .A(n20798), .ZN(n14816) );
  NOR2_X1 U14043 ( .A1(n14816), .A2(n20169), .ZN(n11069) );
  NAND4_X1 U14044 ( .A1(n13555), .A2(n11070), .A3(n11069), .A4(n20822), .ZN(
        n11071) );
  NOR2_X1 U14045 ( .A1(n11072), .A2(n11071), .ZN(n11074) );
  NAND3_X1 U14046 ( .A1(n11055), .A2(n14806), .A3(n11036), .ZN(n11073) );
  NAND3_X1 U14047 ( .A1(n11075), .A2(n11074), .A3(n11073), .ZN(n11108) );
  INV_X1 U14049 ( .A(n11076), .ZN(n11079) );
  NAND2_X1 U14050 ( .A1(n11077), .A2(n14810), .ZN(n11078) );
  NAND2_X1 U14051 ( .A1(n11079), .A2(n11078), .ZN(n11088) );
  NAND2_X1 U14052 ( .A1(n11158), .A2(n11088), .ZN(n11086) );
  AND2_X1 U14053 ( .A1(n20735), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11081) );
  INV_X1 U14054 ( .A(n11917), .ZN(n11171) );
  INV_X1 U14055 ( .A(n11083), .ZN(n11082) );
  NAND2_X1 U14056 ( .A1(n11082), .A2(n20573), .ZN(n20533) );
  NAND2_X1 U14057 ( .A1(n11083), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11084) );
  NAND2_X1 U14058 ( .A1(n20533), .A2(n11084), .ZN(n20171) );
  NAND2_X1 U14059 ( .A1(n11171), .A2(n20171), .ZN(n11087) );
  NAND2_X1 U14060 ( .A1(n11089), .A2(n11087), .ZN(n11085) );
  NAND2_X1 U14061 ( .A1(n11086), .A2(n11085), .ZN(n11168) );
  NAND4_X1 U14062 ( .A1(n11158), .A2(n11089), .A3(n11088), .A4(n11087), .ZN(
        n11090) );
  NAND2_X1 U14063 ( .A1(n11168), .A2(n11090), .ZN(n13381) );
  AOI22_X1 U14064 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14065 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U14066 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11095) );
  AOI22_X1 U14067 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11094) );
  NAND4_X1 U14068 ( .A1(n11097), .A2(n11096), .A3(n11095), .A4(n11094), .ZN(
        n11104) );
  AOI22_X1 U14069 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14070 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U14071 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11100) );
  INV_X1 U14072 ( .A(n11122), .ZN(n11179) );
  BUF_X4 U14073 ( .A(n11127), .Z(n11437) );
  AOI22_X1 U14074 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11099) );
  NAND4_X1 U14075 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n11099), .ZN(
        n11103) );
  INV_X1 U14076 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14077 ( .A1(n9812), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11140) );
  OAI22_X1 U14078 ( .A1(n11903), .A2(n11105), .B1(n11140), .B2(n11778), .ZN(
        n11106) );
  INV_X1 U14079 ( .A(n11108), .ZN(n11109) );
  AOI22_X1 U14080 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14081 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11141), .B1(
        n11730), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14082 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11122), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14083 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11111) );
  NAND4_X1 U14084 ( .A1(n11114), .A2(n11113), .A3(n11112), .A4(n11111), .ZN(
        n11121) );
  AOI22_X1 U14085 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14086 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14087 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14088 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11657), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11116) );
  NAND4_X1 U14089 ( .A1(n11119), .A2(n11118), .A3(n11117), .A4(n11116), .ZN(
        n11120) );
  AOI22_X1 U14090 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11126) );
  AOI22_X1 U14091 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U14092 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11124) );
  AOI22_X1 U14093 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11122), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11123) );
  NAND4_X1 U14094 ( .A1(n11126), .A2(n11125), .A3(n11124), .A4(n11123), .ZN(
        n11133) );
  AOI22_X1 U14095 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11131) );
  AOI22_X1 U14096 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11130) );
  AOI22_X1 U14097 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14098 ( .A1(n11741), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11128) );
  NAND4_X1 U14099 ( .A1(n11131), .A2(n11130), .A3(n11129), .A4(n11128), .ZN(
        n11132) );
  XNOR2_X1 U14100 ( .A(n11833), .B(n11776), .ZN(n11134) );
  NAND2_X1 U14101 ( .A1(n11134), .A2(n11159), .ZN(n11268) );
  INV_X1 U14102 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11137) );
  AOI21_X1 U14103 ( .B1(n9812), .B2(n11776), .A(n20169), .ZN(n11136) );
  NAND2_X1 U14104 ( .A1(n20202), .A2(n11837), .ZN(n11135) );
  OAI211_X1 U14105 ( .C1(n11174), .C2(n11137), .A(n11136), .B(n11135), .ZN(
        n11266) );
  NAND2_X1 U14106 ( .A1(n11159), .A2(n11837), .ZN(n11138) );
  INV_X1 U14107 ( .A(n11140), .ZN(n11152) );
  AOI22_X1 U14108 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11145) );
  AOI22_X1 U14109 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11141), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U14110 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11143) );
  AOI22_X1 U14111 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11142) );
  NAND4_X1 U14112 ( .A1(n11145), .A2(n11144), .A3(n11143), .A4(n11142), .ZN(
        n11151) );
  AOI22_X1 U14113 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14114 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14115 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14116 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11146) );
  NAND4_X1 U14117 ( .A1(n11149), .A2(n11148), .A3(n11147), .A4(n11146), .ZN(
        n11150) );
  AOI22_X1 U14118 ( .A1(n11159), .A2(n11833), .B1(n11152), .B2(n11775), .ZN(
        n11154) );
  INV_X1 U14119 ( .A(n11903), .ZN(n11890) );
  NAND2_X1 U14120 ( .A1(n11890), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11153) );
  INV_X1 U14121 ( .A(n20294), .ZN(n11157) );
  INV_X1 U14122 ( .A(n11155), .ZN(n11156) );
  NAND2_X1 U14123 ( .A1(n11158), .A2(n20231), .ZN(n14802) );
  NAND2_X1 U14124 ( .A1(n11159), .A2(n11775), .ZN(n11160) );
  INV_X1 U14125 ( .A(n11161), .ZN(n11765) );
  NAND2_X1 U14126 ( .A1(n11258), .A2(n11765), .ZN(n11166) );
  INV_X1 U14127 ( .A(n11163), .ZN(n11164) );
  NAND2_X1 U14128 ( .A1(n11166), .A2(n11165), .ZN(n11252) );
  INV_X1 U14129 ( .A(n11252), .ZN(n11167) );
  NAND2_X1 U14130 ( .A1(n11080), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11173) );
  NAND3_X1 U14131 ( .A1(n15688), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20412) );
  INV_X1 U14132 ( .A(n20412), .ZN(n11169) );
  NAND2_X1 U14133 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11169), .ZN(
        n20410) );
  NAND2_X1 U14134 ( .A1(n15688), .A2(n20410), .ZN(n11170) );
  NOR3_X1 U14135 ( .A1(n15688), .A2(n20573), .A3(n20259), .ZN(n20689) );
  NAND2_X1 U14136 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20689), .ZN(
        n20677) );
  AND2_X1 U14137 ( .A1(n11170), .A2(n20677), .ZN(n20437) );
  AOI22_X1 U14138 ( .A1(n11171), .A2(n20437), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20735), .ZN(n11172) );
  XNOR2_X2 U14139 ( .A(n13755), .B(n20328), .ZN(n20436) );
  NAND2_X1 U14140 ( .A1(n20436), .A2(n20169), .ZN(n11189) );
  INV_X1 U14141 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U14142 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11178) );
  AOI22_X1 U14143 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11683), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U14144 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U14145 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11175) );
  NAND4_X1 U14146 ( .A1(n11178), .A2(n11177), .A3(n11176), .A4(n11175), .ZN(
        n11185) );
  AOI22_X1 U14147 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11183) );
  AOI22_X1 U14148 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U14149 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11181) );
  INV_X2 U14150 ( .A(n11179), .ZN(n11739) );
  AOI22_X1 U14151 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11180) );
  NAND4_X1 U14152 ( .A1(n11183), .A2(n11182), .A3(n11181), .A4(n11180), .ZN(
        n11184) );
  OAI22_X1 U14153 ( .A1(n11186), .A2(n11903), .B1(n11907), .B2(n11787), .ZN(
        n11187) );
  INV_X1 U14154 ( .A(n11187), .ZN(n11188) );
  INV_X1 U14155 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14156 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14157 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11683), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14158 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U14159 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11191) );
  NAND4_X1 U14160 ( .A1(n11194), .A2(n11193), .A3(n11192), .A4(n11191), .ZN(
        n11200) );
  AOI22_X1 U14161 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14162 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14163 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14164 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11195) );
  NAND4_X1 U14165 ( .A1(n11198), .A2(n11197), .A3(n11196), .A4(n11195), .ZN(
        n11199) );
  INV_X1 U14166 ( .A(n11797), .ZN(n11806) );
  OR2_X1 U14167 ( .A1(n11907), .A2(n11806), .ZN(n11201) );
  INV_X1 U14168 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14169 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14170 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11206) );
  AOI22_X1 U14171 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14172 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11204) );
  NAND4_X1 U14173 ( .A1(n11207), .A2(n11206), .A3(n11205), .A4(n11204), .ZN(
        n11213) );
  AOI22_X1 U14174 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14175 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14176 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14177 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11208) );
  NAND4_X1 U14178 ( .A1(n11211), .A2(n11210), .A3(n11209), .A4(n11208), .ZN(
        n11212) );
  OR2_X1 U14179 ( .A1(n11907), .A2(n11818), .ZN(n11214) );
  OAI21_X1 U14180 ( .B1(n11903), .B2(n11215), .A(n11214), .ZN(n11296) );
  INV_X1 U14181 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14182 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11203), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14183 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14184 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14185 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11216) );
  NAND4_X1 U14186 ( .A1(n11219), .A2(n11218), .A3(n11217), .A4(n11216), .ZN(
        n11225) );
  AOI22_X1 U14187 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14188 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14189 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14190 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11220) );
  NAND4_X1 U14191 ( .A1(n11223), .A2(n11222), .A3(n11221), .A4(n11220), .ZN(
        n11224) );
  INV_X1 U14192 ( .A(n11820), .ZN(n11226) );
  OR2_X1 U14193 ( .A1(n11907), .A2(n11226), .ZN(n11227) );
  OAI21_X1 U14194 ( .B1(n11903), .B2(n11228), .A(n11227), .ZN(n11303) );
  INV_X1 U14195 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11229) );
  OAI22_X1 U14196 ( .A1(n11229), .A2(n11903), .B1(n11907), .B2(n11833), .ZN(
        n11230) );
  XNOR2_X1 U14197 ( .A(n11816), .B(n11230), .ZN(n11828) );
  NAND2_X1 U14198 ( .A1(n11828), .A2(n11395), .ZN(n11236) );
  INV_X1 U14199 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11233) );
  NOR2_X1 U14200 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11265) );
  OAI21_X1 U14201 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11307), .A(
        n11317), .ZN(n20033) );
  AOI22_X1 U14202 ( .A1(n13998), .A2(n20033), .B1(n11757), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11232) );
  OAI21_X1 U14203 ( .B1(n11272), .B2(n11233), .A(n11232), .ZN(n11234) );
  INV_X1 U14204 ( .A(n11234), .ZN(n11235) );
  NAND2_X1 U14205 ( .A1(n11236), .A2(n11235), .ZN(n14025) );
  XOR2_X1 U14206 ( .A(n11316), .B(n11317), .Z(n14197) );
  AOI22_X1 U14207 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14208 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11203), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U14209 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11238) );
  AOI22_X1 U14210 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11237) );
  NAND4_X1 U14211 ( .A1(n11240), .A2(n11239), .A3(n11238), .A4(n11237), .ZN(
        n11246) );
  AOI22_X1 U14212 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14213 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14214 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14215 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11241) );
  NAND4_X1 U14216 ( .A1(n11244), .A2(n11243), .A3(n11242), .A4(n11241), .ZN(
        n11245) );
  OR2_X1 U14217 ( .A1(n11246), .A2(n11245), .ZN(n11248) );
  INV_X1 U14218 ( .A(n11757), .ZN(n11369) );
  NOR2_X1 U14219 ( .A1(n11369), .A2(n11316), .ZN(n11247) );
  AOI21_X1 U14220 ( .B1(n11395), .B2(n11248), .A(n11247), .ZN(n11250) );
  NAND2_X1 U14221 ( .A1(n11758), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11249) );
  OAI211_X1 U14222 ( .C1(n14197), .C2(n11750), .A(n11250), .B(n11249), .ZN(
        n14026) );
  NAND2_X1 U14223 ( .A1(n11251), .A2(n11252), .ZN(n11253) );
  INV_X1 U14224 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n11255) );
  NAND2_X1 U14225 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11279) );
  OAI21_X1 U14226 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n11279), .ZN(n20094) );
  OAI21_X1 U14227 ( .B1(n20094), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20813), 
        .ZN(n11254) );
  OAI21_X1 U14228 ( .B1(n11272), .B2(n11255), .A(n11254), .ZN(n11256) );
  AOI21_X1 U14229 ( .B1(n11288), .B2(n13751), .A(n11256), .ZN(n11257) );
  NAND2_X1 U14230 ( .A1(n11757), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13657) );
  INV_X1 U14231 ( .A(n11258), .ZN(n11260) );
  INV_X1 U14232 ( .A(n11765), .ZN(n11259) );
  XNOR2_X2 U14233 ( .A(n11260), .B(n11259), .ZN(n13763) );
  NAND2_X1 U14234 ( .A1(n13763), .A2(n11395), .ZN(n11264) );
  INV_X1 U14235 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11261) );
  INV_X1 U14236 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13639) );
  OAI22_X1 U14237 ( .A1(n11272), .A2(n11261), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13639), .ZN(n11262) );
  AOI21_X1 U14238 ( .B1(n11288), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11262), .ZN(n11263) );
  NAND2_X1 U14239 ( .A1(n11264), .A2(n11263), .ZN(n13584) );
  MUX2_X1 U14240 ( .A(n11268), .B(n11267), .S(n11266), .Z(n20257) );
  AOI21_X1 U14241 ( .B1(n20257), .B2(n20215), .A(n20813), .ZN(n13406) );
  NAND2_X1 U14242 ( .A1(n11269), .A2(n11395), .ZN(n11275) );
  INV_X1 U14243 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n11271) );
  INV_X1 U14244 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11270) );
  OAI22_X1 U14245 ( .A1(n11272), .A2(n11271), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11270), .ZN(n11273) );
  AOI21_X1 U14246 ( .B1(n11288), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11273), .ZN(n11274) );
  NAND2_X1 U14247 ( .A1(n11275), .A2(n11274), .ZN(n13404) );
  MUX2_X1 U14248 ( .A(n11265), .B(n13406), .S(n13404), .Z(n13585) );
  NAND2_X1 U14249 ( .A1(n13584), .A2(n13585), .ZN(n13615) );
  NAND2_X1 U14250 ( .A1(n13613), .A2(n13657), .ZN(n11285) );
  INV_X1 U14251 ( .A(n13791), .ZN(n13790) );
  NAND2_X1 U14252 ( .A1(n11277), .A2(n13790), .ZN(n11278) );
  INV_X1 U14253 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11282) );
  INV_X1 U14254 ( .A(n11279), .ZN(n11280) );
  OAI21_X1 U14255 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11280), .A(
        n11290), .ZN(n14063) );
  AOI22_X1 U14256 ( .A1(n13998), .A2(n14063), .B1(n11757), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11281) );
  OAI21_X1 U14257 ( .B1(n11272), .B2(n11282), .A(n11281), .ZN(n11283) );
  AOI21_X1 U14258 ( .B1(n11288), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11283), .ZN(n11284) );
  NAND2_X1 U14259 ( .A1(n11285), .A2(n13656), .ZN(n13655) );
  INV_X1 U14260 ( .A(n13655), .ZN(n11295) );
  XNOR2_X1 U14261 ( .A(n11287), .B(n11286), .ZN(n11794) );
  NAND2_X1 U14262 ( .A1(n11288), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11292) );
  AOI21_X1 U14263 ( .B1(n13903), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11289) );
  AOI21_X1 U14264 ( .B1(n11758), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11289), .ZN(
        n11291) );
  AOI21_X1 U14265 ( .B1(n13903), .B2(n11290), .A(n11298), .ZN(n20076) );
  AOI22_X1 U14266 ( .A1(n11292), .A2(n11291), .B1(n13998), .B2(n20076), .ZN(
        n11293) );
  NAND2_X1 U14267 ( .A1(n11295), .A2(n11294), .ZN(n13899) );
  INV_X1 U14268 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11300) );
  OAI21_X1 U14269 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11298), .A(
        n11306), .ZN(n20066) );
  AOI22_X1 U14270 ( .A1(n13998), .A2(n20066), .B1(n11757), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11299) );
  OAI21_X1 U14271 ( .B1(n11272), .B2(n11300), .A(n11299), .ZN(n11301) );
  INV_X1 U14272 ( .A(n11302), .ZN(n11305) );
  INV_X1 U14273 ( .A(n11303), .ZN(n11304) );
  NAND2_X1 U14274 ( .A1(n11305), .A2(n11304), .ZN(n11817) );
  NAND2_X1 U14275 ( .A1(n11817), .A2(n11395), .ZN(n11314) );
  INV_X1 U14276 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11311) );
  INV_X1 U14277 ( .A(n11306), .ZN(n11309) );
  INV_X1 U14278 ( .A(n11307), .ZN(n11308) );
  OAI21_X1 U14279 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11309), .A(
        n11308), .ZN(n20052) );
  AOI22_X1 U14280 ( .A1(n13998), .A2(n20052), .B1(n11757), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11310) );
  OAI21_X1 U14281 ( .B1(n11272), .B2(n11311), .A(n11310), .ZN(n11312) );
  INV_X1 U14282 ( .A(n11312), .ZN(n11313) );
  XNOR2_X1 U14283 ( .A(n11334), .B(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14469) );
  NAND2_X1 U14284 ( .A1(n14469), .A2(n13998), .ZN(n11333) );
  AOI22_X1 U14285 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14286 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14287 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14288 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11318) );
  NAND4_X1 U14289 ( .A1(n11321), .A2(n11320), .A3(n11319), .A4(n11318), .ZN(
        n11327) );
  AOI22_X1 U14290 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14291 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14292 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14293 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11322) );
  NAND4_X1 U14294 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11326) );
  NOR2_X1 U14295 ( .A1(n11327), .A2(n11326), .ZN(n11330) );
  NAND2_X1 U14296 ( .A1(n11758), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11329) );
  NAND2_X1 U14297 ( .A1(n11757), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11328) );
  OAI211_X1 U14298 ( .C1(n11447), .C2(n11330), .A(n11329), .B(n11328), .ZN(
        n11331) );
  INV_X1 U14299 ( .A(n11331), .ZN(n11332) );
  NAND2_X1 U14300 ( .A1(n11333), .A2(n11332), .ZN(n14085) );
  XOR2_X1 U14301 ( .A(n11348), .B(n11349), .Z(n15941) );
  AOI22_X1 U14302 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14303 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14304 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14305 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11335) );
  NAND4_X1 U14306 ( .A1(n11338), .A2(n11337), .A3(n11336), .A4(n11335), .ZN(
        n11344) );
  AOI22_X1 U14307 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11203), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14308 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14309 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14310 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11339) );
  NAND4_X1 U14311 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n11343) );
  OR2_X1 U14312 ( .A1(n11344), .A2(n11343), .ZN(n11345) );
  AOI22_X1 U14313 ( .A1(n11395), .A2(n11345), .B1(n11757), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11347) );
  NAND2_X1 U14314 ( .A1(n11758), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11346) );
  OAI211_X1 U14315 ( .C1(n15941), .C2(n11750), .A(n11347), .B(n11346), .ZN(
        n14132) );
  XNOR2_X1 U14316 ( .A(n11368), .B(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14685) );
  INV_X1 U14317 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20126) );
  INV_X1 U14318 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14228) );
  OAI22_X1 U14319 ( .A1(n11272), .A2(n20126), .B1(n11369), .B2(n14228), .ZN(
        n11350) );
  AOI21_X1 U14320 ( .B1(n14685), .B2(n13998), .A(n11350), .ZN(n11365) );
  INV_X1 U14321 ( .A(n14210), .ZN(n11363) );
  AOI22_X1 U14322 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11730), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14323 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11740), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14324 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14325 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11351) );
  NAND4_X1 U14326 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11360) );
  AOI22_X1 U14327 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14328 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14329 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11356) );
  AOI22_X1 U14330 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11355) );
  NAND4_X1 U14331 ( .A1(n11358), .A2(n11357), .A3(n11356), .A4(n11355), .ZN(
        n11359) );
  OR2_X1 U14332 ( .A1(n11360), .A2(n11359), .ZN(n11361) );
  NAND2_X1 U14333 ( .A1(n11395), .A2(n11361), .ZN(n14211) );
  INV_X1 U14334 ( .A(n14211), .ZN(n11362) );
  XNOR2_X1 U14335 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11383), .ZN(
        n15849) );
  OAI22_X1 U14336 ( .A1(n11750), .A2(n15849), .B1(n11369), .B2(n14677), .ZN(
        n11370) );
  AOI21_X1 U14337 ( .B1(n11758), .B2(P1_EAX_REG_12__SCAN_IN), .A(n11370), .ZN(
        n11382) );
  AOI22_X1 U14338 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11203), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14339 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14340 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14341 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11371) );
  NAND4_X1 U14342 ( .A1(n11374), .A2(n11373), .A3(n11372), .A4(n11371), .ZN(
        n11380) );
  AOI22_X1 U14343 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14344 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14345 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14346 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11375) );
  NAND4_X1 U14347 ( .A1(n11378), .A2(n11377), .A3(n11376), .A4(n11375), .ZN(
        n11379) );
  OAI21_X1 U14348 ( .B1(n11380), .B2(n11379), .A(n11395), .ZN(n11381) );
  XOR2_X1 U14349 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11398), .Z(
        n15838) );
  AOI22_X1 U14350 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14351 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11203), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11386) );
  AOI22_X1 U14352 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14353 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11384) );
  NAND4_X1 U14354 ( .A1(n11387), .A2(n11386), .A3(n11385), .A4(n11384), .ZN(
        n11393) );
  AOI22_X1 U14355 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14356 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14357 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14358 ( .A1(n11732), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11388) );
  NAND4_X1 U14359 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n11392) );
  OR2_X1 U14360 ( .A1(n11393), .A2(n11392), .ZN(n11394) );
  AOI22_X1 U14361 ( .A1(n11395), .A2(n11394), .B1(n11757), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U14362 ( .A1(n11758), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11396) );
  OAI211_X1 U14363 ( .C1(n15838), .C2(n11750), .A(n11397), .B(n11396), .ZN(
        n14241) );
  XNOR2_X1 U14364 ( .A(n11415), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14662) );
  NAND2_X1 U14365 ( .A1(n14662), .A2(n13998), .ZN(n11414) );
  AOI22_X1 U14366 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14367 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14368 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14369 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11399) );
  NAND4_X1 U14370 ( .A1(n11402), .A2(n11401), .A3(n11400), .A4(n11399), .ZN(
        n11408) );
  AOI22_X1 U14371 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14372 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14373 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14374 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11403) );
  NAND4_X1 U14375 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11407) );
  NOR2_X1 U14376 ( .A1(n11408), .A2(n11407), .ZN(n11411) );
  NAND2_X1 U14377 ( .A1(n11758), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11410) );
  NAND2_X1 U14378 ( .A1(n11757), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11409) );
  OAI211_X1 U14379 ( .C1(n11447), .C2(n11411), .A(n11410), .B(n11409), .ZN(
        n11412) );
  INV_X1 U14380 ( .A(n11412), .ZN(n11413) );
  NAND2_X1 U14381 ( .A1(n11414), .A2(n11413), .ZN(n14277) );
  XNOR2_X1 U14382 ( .A(n11450), .B(n14451), .ZN(n14656) );
  AOI22_X1 U14383 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14384 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11730), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14385 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14386 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11416) );
  NAND4_X1 U14387 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n11427) );
  AOI22_X1 U14388 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11425) );
  NAND2_X1 U14389 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11421) );
  NAND2_X1 U14390 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11420) );
  AND3_X1 U14391 ( .A1(n11421), .A2(n11420), .A3(n11750), .ZN(n11424) );
  AOI22_X1 U14392 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14393 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11422) );
  NAND4_X1 U14394 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11426) );
  NAND2_X1 U14395 ( .A1(n11720), .A2(n11750), .ZN(n11552) );
  OAI21_X1 U14396 ( .B1(n11427), .B2(n11426), .A(n11552), .ZN(n11430) );
  NAND2_X1 U14397 ( .A1(n11758), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n11429) );
  NAND2_X1 U14398 ( .A1(n20813), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11428) );
  NAND3_X1 U14399 ( .A1(n11430), .A2(n11429), .A3(n11428), .ZN(n11431) );
  OAI21_X1 U14400 ( .B1(n14656), .B2(n11750), .A(n11431), .ZN(n14444) );
  XOR2_X1 U14401 ( .A(n15825), .B(n11432), .Z(n15934) );
  INV_X1 U14402 ( .A(n15934), .ZN(n11449) );
  AOI22_X1 U14403 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14404 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14405 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14406 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11702), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U14407 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n11443) );
  AOI22_X1 U14408 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n11657), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14409 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14410 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11637), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14411 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11438) );
  NAND4_X1 U14412 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n11442) );
  NOR2_X1 U14413 ( .A1(n11443), .A2(n11442), .ZN(n11446) );
  NAND2_X1 U14414 ( .A1(n11758), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11445) );
  NAND2_X1 U14415 ( .A1(n11757), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11444) );
  OAI211_X1 U14416 ( .C1(n11447), .C2(n11446), .A(n11445), .B(n11444), .ZN(
        n11448) );
  AOI21_X1 U14417 ( .B1(n11449), .B2(n13998), .A(n11448), .ZN(n14547) );
  XOR2_X1 U14418 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11465), .Z(
        n15808) );
  INV_X1 U14419 ( .A(n15808), .ZN(n15922) );
  AOI22_X1 U14420 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11203), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14421 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14422 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14423 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11451) );
  NAND4_X1 U14424 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(
        n11460) );
  AOI22_X1 U14425 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14426 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14427 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14428 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11455) );
  NAND4_X1 U14429 ( .A1(n11458), .A2(n11457), .A3(n11456), .A4(n11455), .ZN(
        n11459) );
  NOR2_X1 U14430 ( .A1(n11460), .A2(n11459), .ZN(n11463) );
  NAND2_X1 U14431 ( .A1(n11758), .A2(P1_EAX_REG_17__SCAN_IN), .ZN(n11462) );
  NAND2_X1 U14432 ( .A1(n11757), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11461) );
  OAI211_X1 U14433 ( .C1(n11720), .C2(n11463), .A(n11462), .B(n11461), .ZN(
        n11464) );
  AOI21_X1 U14434 ( .B1(n15922), .B2(n13998), .A(n11464), .ZN(n15809) );
  XNOR2_X1 U14435 ( .A(n11497), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15805) );
  AOI22_X1 U14436 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U14437 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11467) );
  NAND2_X1 U14438 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11466) );
  AND3_X1 U14439 ( .A1(n11467), .A2(n11466), .A3(n11750), .ZN(n11470) );
  AOI22_X1 U14440 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14441 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11468) );
  NAND4_X1 U14442 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n11477) );
  AOI22_X1 U14443 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14444 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14445 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14446 ( .A1(n11540), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11472) );
  NAND4_X1 U14447 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(
        n11476) );
  OR2_X1 U14448 ( .A1(n11477), .A2(n11476), .ZN(n11480) );
  INV_X1 U14449 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n11478) );
  OAI22_X1 U14450 ( .A1(n11272), .A2(n11478), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15800), .ZN(n11479) );
  AOI21_X1 U14451 ( .B1(n11552), .B2(n11480), .A(n11479), .ZN(n11481) );
  AOI21_X1 U14452 ( .B1(n15805), .B2(n13998), .A(n11481), .ZN(n14496) );
  NAND2_X1 U14453 ( .A1(n14493), .A2(n14496), .ZN(n14494) );
  AOI22_X1 U14454 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14455 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11730), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14456 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14457 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11482) );
  NAND4_X1 U14458 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11491) );
  AOI22_X1 U14459 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14460 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14461 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14462 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14463 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11490) );
  NOR2_X1 U14464 ( .A1(n11491), .A2(n11490), .ZN(n11496) );
  INV_X1 U14465 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n11493) );
  NAND2_X1 U14466 ( .A1(n20813), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11492) );
  OAI211_X1 U14467 ( .C1(n11272), .C2(n11493), .A(n11750), .B(n11492), .ZN(
        n11494) );
  INV_X1 U14468 ( .A(n11494), .ZN(n11495) );
  OAI21_X1 U14469 ( .B1(n11720), .B2(n11496), .A(n11495), .ZN(n11500) );
  OAI21_X1 U14470 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11498), .A(
        n11531), .ZN(n15915) );
  OR2_X1 U14471 ( .A1(n11750), .A2(n15915), .ZN(n11499) );
  NAND2_X1 U14472 ( .A1(n11500), .A2(n11499), .ZN(n15792) );
  AOI22_X1 U14473 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11203), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14474 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14475 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14476 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11501) );
  NAND4_X1 U14477 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11510) );
  AOI22_X1 U14478 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14479 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14480 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14481 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11505) );
  NAND4_X1 U14482 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n11509) );
  NOR2_X1 U14483 ( .A1(n11510), .A2(n11509), .ZN(n11513) );
  INV_X1 U14484 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15786) );
  AOI21_X1 U14485 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15786), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11511) );
  AOI21_X1 U14486 ( .B1(n11758), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11511), .ZN(
        n11512) );
  OAI21_X1 U14487 ( .B1(n11720), .B2(n11513), .A(n11512), .ZN(n11515) );
  XNOR2_X1 U14488 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11531), .ZN(
        n15776) );
  NAND2_X1 U14489 ( .A1(n13998), .A2(n15776), .ZN(n11514) );
  NAND2_X1 U14490 ( .A1(n11515), .A2(n11514), .ZN(n14489) );
  AOI22_X1 U14491 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14492 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14493 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U14494 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11517) );
  NAND4_X1 U14495 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(
        n11526) );
  AOI22_X1 U14496 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11203), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14497 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14498 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11522) );
  NAND4_X1 U14499 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11525) );
  NOR2_X1 U14500 ( .A1(n11526), .A2(n11525), .ZN(n11530) );
  INV_X1 U14501 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21176) );
  INV_X1 U14502 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21140) );
  OAI21_X1 U14503 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21140), .A(
        n20813), .ZN(n11527) );
  OAI21_X1 U14504 ( .B1(n11272), .B2(n21176), .A(n11527), .ZN(n11528) );
  INV_X1 U14505 ( .A(n11528), .ZN(n11529) );
  OAI21_X1 U14506 ( .B1(n11720), .B2(n11530), .A(n11529), .ZN(n11537) );
  INV_X1 U14507 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11533) );
  INV_X1 U14508 ( .A(n11534), .ZN(n11532) );
  NAND2_X1 U14509 ( .A1(n11533), .A2(n11532), .ZN(n11535) );
  AND2_X1 U14510 ( .A1(n11535), .A2(n11585), .ZN(n15901) );
  NAND2_X1 U14511 ( .A1(n15901), .A2(n13998), .ZN(n11536) );
  NAND2_X1 U14512 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11539) );
  NAND2_X1 U14513 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11538) );
  AND3_X1 U14514 ( .A1(n11539), .A2(n11538), .A3(n11750), .ZN(n11544) );
  AOI22_X1 U14515 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14516 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11542) );
  NAND4_X1 U14517 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .ZN(
        n11550) );
  AOI22_X1 U14518 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U14519 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14520 ( .A1(n11203), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14521 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11545) );
  NAND4_X1 U14522 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n11549) );
  OR2_X1 U14523 ( .A1(n11550), .A2(n11549), .ZN(n11551) );
  NAND2_X1 U14524 ( .A1(n11552), .A2(n11551), .ZN(n11557) );
  INV_X1 U14525 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n11553) );
  INV_X1 U14526 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14633) );
  OAI22_X1 U14527 ( .A1(n11272), .A2(n11553), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14633), .ZN(n11554) );
  INV_X1 U14528 ( .A(n11554), .ZN(n11556) );
  XNOR2_X1 U14529 ( .A(n11585), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14637) );
  AOI21_X1 U14530 ( .B1(n11557), .B2(n11556), .A(n11555), .ZN(n14434) );
  AOI22_X1 U14531 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10961), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14532 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14533 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14534 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11559) );
  NAND4_X1 U14535 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11568) );
  AOI22_X1 U14536 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11203), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14537 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14538 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14539 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11563) );
  NAND4_X1 U14540 ( .A1(n11566), .A2(n11565), .A3(n11564), .A4(n11563), .ZN(
        n11567) );
  NOR2_X1 U14541 ( .A1(n11568), .A2(n11567), .ZN(n11593) );
  AOI22_X1 U14542 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11203), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14543 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11731), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14544 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14545 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11570) );
  NAND4_X1 U14546 ( .A1(n11573), .A2(n11572), .A3(n11571), .A4(n11570), .ZN(
        n11579) );
  AOI22_X1 U14547 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14548 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14549 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14550 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11574) );
  NAND4_X1 U14551 ( .A1(n11577), .A2(n11576), .A3(n11575), .A4(n11574), .ZN(
        n11578) );
  NOR2_X1 U14552 ( .A1(n11579), .A2(n11578), .ZN(n11594) );
  XNOR2_X1 U14553 ( .A(n11593), .B(n11594), .ZN(n11584) );
  INV_X1 U14554 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14555 ( .A1(n20813), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11580) );
  OAI211_X1 U14556 ( .C1(n11272), .C2(n11581), .A(n11750), .B(n11580), .ZN(
        n11582) );
  INV_X1 U14557 ( .A(n11582), .ZN(n11583) );
  OAI21_X1 U14558 ( .B1(n11720), .B2(n11584), .A(n11583), .ZN(n11592) );
  INV_X1 U14559 ( .A(n11587), .ZN(n11589) );
  INV_X1 U14560 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11588) );
  NAND2_X1 U14561 ( .A1(n11589), .A2(n11588), .ZN(n11590) );
  AND2_X1 U14562 ( .A1(n11628), .A2(n11590), .ZN(n14422) );
  NAND2_X1 U14563 ( .A1(n14422), .A2(n11265), .ZN(n11591) );
  NAND2_X1 U14564 ( .A1(n11592), .A2(n11591), .ZN(n14421) );
  NOR2_X1 U14565 ( .A1(n11594), .A2(n11593), .ZN(n11613) );
  AOI22_X1 U14566 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14567 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11683), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14568 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14569 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11595) );
  NAND4_X1 U14570 ( .A1(n11598), .A2(n11597), .A3(n11596), .A4(n11595), .ZN(
        n11604) );
  AOI22_X1 U14571 ( .A1(n11702), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14572 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14573 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11600) );
  NAND4_X1 U14574 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11603) );
  OR2_X1 U14575 ( .A1(n11604), .A2(n11603), .ZN(n11612) );
  XNOR2_X1 U14576 ( .A(n11613), .B(n11612), .ZN(n11609) );
  INV_X1 U14577 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n11606) );
  NAND2_X1 U14578 ( .A1(n20813), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11605) );
  OAI211_X1 U14579 ( .C1(n11272), .C2(n11606), .A(n11750), .B(n11605), .ZN(
        n11607) );
  INV_X1 U14580 ( .A(n11607), .ZN(n11608) );
  OAI21_X1 U14581 ( .B1(n11609), .B2(n11720), .A(n11608), .ZN(n11611) );
  XNOR2_X1 U14582 ( .A(n11628), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14613) );
  NAND2_X1 U14583 ( .A1(n14613), .A2(n13998), .ZN(n11610) );
  NAND2_X1 U14584 ( .A1(n11613), .A2(n11612), .ZN(n11635) );
  AOI22_X1 U14585 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14586 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14587 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11614) );
  NAND4_X1 U14588 ( .A1(n11617), .A2(n11616), .A3(n11615), .A4(n11614), .ZN(
        n11623) );
  AOI22_X1 U14589 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11657), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14590 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11730), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14591 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14592 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11618) );
  NAND4_X1 U14593 ( .A1(n11621), .A2(n11620), .A3(n11619), .A4(n11618), .ZN(
        n11622) );
  NOR2_X1 U14594 ( .A1(n11623), .A2(n11622), .ZN(n11636) );
  XNOR2_X1 U14595 ( .A(n11635), .B(n11636), .ZN(n11627) );
  INV_X1 U14596 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21141) );
  OAI21_X1 U14597 ( .B1(n21140), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n20813), .ZN(n11624) );
  OAI21_X1 U14598 ( .B1(n11272), .B2(n21141), .A(n11624), .ZN(n11625) );
  INV_X1 U14599 ( .A(n11625), .ZN(n11626) );
  OAI21_X1 U14600 ( .B1(n11627), .B2(n11720), .A(n11626), .ZN(n11634) );
  INV_X1 U14601 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11630) );
  NAND2_X1 U14602 ( .A1(n11631), .A2(n11630), .ZN(n11632) );
  NAND2_X1 U14603 ( .A1(n11675), .A2(n11632), .ZN(n14607) );
  NOR2_X1 U14604 ( .A1(n11636), .A2(n11635), .ZN(n11669) );
  AOI22_X1 U14605 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14606 ( .A1(n11638), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11637), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14607 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14608 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11540), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11639) );
  NAND4_X1 U14609 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n11648) );
  AOI22_X1 U14610 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14611 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14612 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11644) );
  NAND4_X1 U14613 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11647) );
  OR2_X1 U14614 ( .A1(n11648), .A2(n11647), .ZN(n11668) );
  INV_X1 U14615 ( .A(n11668), .ZN(n11649) );
  XNOR2_X1 U14616 ( .A(n11669), .B(n11649), .ZN(n11650) );
  INV_X1 U14617 ( .A(n11720), .ZN(n11754) );
  NAND2_X1 U14618 ( .A1(n11650), .A2(n11754), .ZN(n11656) );
  INV_X1 U14619 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n11652) );
  NAND2_X1 U14620 ( .A1(n20813), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11651) );
  OAI211_X1 U14621 ( .C1(n11272), .C2(n11652), .A(n11750), .B(n11651), .ZN(
        n11653) );
  INV_X1 U14622 ( .A(n11653), .ZN(n11655) );
  XNOR2_X1 U14623 ( .A(n11675), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14599) );
  AOI22_X1 U14624 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11569), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14625 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14626 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14627 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11658) );
  NAND4_X1 U14628 ( .A1(n11661), .A2(n11660), .A3(n11659), .A4(n11658), .ZN(
        n11667) );
  AOI22_X1 U14629 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14630 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11730), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14631 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14632 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11662) );
  NAND4_X1 U14633 ( .A1(n11665), .A2(n11664), .A3(n11663), .A4(n11662), .ZN(
        n11666) );
  NOR2_X1 U14634 ( .A1(n11667), .A2(n11666), .ZN(n11682) );
  NAND2_X1 U14635 ( .A1(n11669), .A2(n11668), .ZN(n11681) );
  XNOR2_X1 U14636 ( .A(n11682), .B(n11681), .ZN(n11674) );
  INV_X1 U14637 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n11671) );
  NAND2_X1 U14638 ( .A1(n20813), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11670) );
  OAI211_X1 U14639 ( .C1(n11272), .C2(n11671), .A(n11750), .B(n11670), .ZN(
        n11672) );
  INV_X1 U14640 ( .A(n11672), .ZN(n11673) );
  OAI21_X1 U14641 ( .B1(n11674), .B2(n11720), .A(n11673), .ZN(n11680) );
  INV_X1 U14642 ( .A(n11675), .ZN(n11676) );
  NAND2_X1 U14643 ( .A1(n11676), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11677) );
  INV_X1 U14644 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14587) );
  NAND2_X1 U14645 ( .A1(n11677), .A2(n14587), .ZN(n11678) );
  NAND2_X1 U14646 ( .A1(n14585), .A2(n11265), .ZN(n11679) );
  NAND2_X1 U14647 ( .A1(n11680), .A2(n11679), .ZN(n14371) );
  NOR2_X1 U14648 ( .A1(n11682), .A2(n11681), .ZN(n11715) );
  AOI22_X1 U14649 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14650 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11683), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14651 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14652 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11684) );
  NAND4_X1 U14653 ( .A1(n11687), .A2(n11686), .A3(n11685), .A4(n11684), .ZN(
        n11693) );
  AOI22_X1 U14654 ( .A1(n11730), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11731), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14655 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14656 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U14657 ( .A1(n11691), .A2(n11690), .A3(n11689), .A4(n11688), .ZN(
        n11692) );
  OR2_X1 U14658 ( .A1(n11693), .A2(n11692), .ZN(n11714) );
  XNOR2_X1 U14659 ( .A(n11715), .B(n11714), .ZN(n11698) );
  INV_X1 U14660 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n11695) );
  NAND2_X1 U14661 ( .A1(n20813), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11694) );
  OAI211_X1 U14662 ( .C1(n11272), .C2(n11695), .A(n11750), .B(n11694), .ZN(
        n11696) );
  INV_X1 U14663 ( .A(n11696), .ZN(n11697) );
  OAI21_X1 U14664 ( .B1(n11698), .B2(n11720), .A(n11697), .ZN(n11700) );
  XNOR2_X1 U14665 ( .A(n11722), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14575) );
  NAND2_X1 U14666 ( .A1(n14575), .A2(n13998), .ZN(n11699) );
  AOI22_X1 U14667 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14668 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11702), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14669 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14670 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11703) );
  NAND4_X1 U14671 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(
        n11713) );
  AOI22_X1 U14672 ( .A1(n10973), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14673 ( .A1(n11707), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14674 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14675 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10992), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11708) );
  NAND4_X1 U14676 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11712) );
  NOR2_X1 U14677 ( .A1(n11713), .A2(n11712), .ZN(n11729) );
  NAND2_X1 U14678 ( .A1(n11715), .A2(n11714), .ZN(n11728) );
  XNOR2_X1 U14679 ( .A(n11729), .B(n11728), .ZN(n11721) );
  INV_X1 U14680 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n11717) );
  NAND2_X1 U14681 ( .A1(n20813), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11716) );
  OAI211_X1 U14682 ( .C1(n11272), .C2(n11717), .A(n11750), .B(n11716), .ZN(
        n11718) );
  INV_X1 U14683 ( .A(n11718), .ZN(n11719) );
  OAI21_X1 U14684 ( .B1(n11721), .B2(n11720), .A(n11719), .ZN(n11727) );
  INV_X1 U14685 ( .A(n11722), .ZN(n11723) );
  NAND2_X1 U14686 ( .A1(n11723), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11724) );
  INV_X1 U14687 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14352) );
  NAND2_X1 U14688 ( .A1(n11724), .A2(n14352), .ZN(n11725) );
  NAND2_X1 U14689 ( .A1(n11920), .A2(n11725), .ZN(n14566) );
  NAND2_X1 U14690 ( .A1(n11727), .A2(n11726), .ZN(n13095) );
  XNOR2_X1 U14691 ( .A(n11920), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14555) );
  NOR2_X1 U14692 ( .A1(n11729), .A2(n11728), .ZN(n11749) );
  AOI22_X1 U14693 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n11203), .B1(
        n10972), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14694 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n11731), .B1(
        n11730), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14695 ( .A1(n10961), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U14696 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11437), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11734) );
  NAND4_X1 U14697 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n11747) );
  AOI22_X1 U14698 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U14699 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11637), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U14700 ( .A1(n11740), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14701 ( .A1(n11657), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11742) );
  NAND4_X1 U14702 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11746) );
  NOR2_X1 U14703 ( .A1(n11747), .A2(n11746), .ZN(n11748) );
  XNOR2_X1 U14704 ( .A(n11749), .B(n11748), .ZN(n11755) );
  INV_X1 U14705 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U14706 ( .A1(n20813), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11751) );
  OAI211_X1 U14707 ( .C1(n11272), .C2(n11752), .A(n11751), .B(n11750), .ZN(
        n11753) );
  AOI21_X1 U14708 ( .B1(n11755), .B2(n11754), .A(n11753), .ZN(n11756) );
  NAND2_X1 U14709 ( .A1(n13094), .A2(n13184), .ZN(n11761) );
  AOI22_X1 U14710 ( .A1(n11758), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n11757), .ZN(n11759) );
  XNOR2_X2 U14711 ( .A(n11761), .B(n11760), .ZN(n14323) );
  AND2_X1 U14712 ( .A1(n20169), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20818) );
  NAND2_X1 U14713 ( .A1(n14323), .A2(n20166), .ZN(n11925) );
  NAND2_X1 U14714 ( .A1(n9812), .A2(n11762), .ZN(n11779) );
  OAI21_X1 U14715 ( .B1(n20819), .B2(n11776), .A(n11779), .ZN(n11763) );
  INV_X1 U14716 ( .A(n11763), .ZN(n11764) );
  OAI21_X1 U14717 ( .B1(n20257), .B2(n11872), .A(n11764), .ZN(n13409) );
  NAND2_X1 U14718 ( .A1(n13409), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13408) );
  NAND2_X1 U14719 ( .A1(n11765), .A2(n11036), .ZN(n11769) );
  XNOR2_X1 U14720 ( .A(n11776), .B(n11775), .ZN(n11766) );
  OAI211_X1 U14721 ( .C1(n11766), .C2(n20819), .A(n20190), .B(n11031), .ZN(
        n11767) );
  INV_X1 U14722 ( .A(n11767), .ZN(n11768) );
  NAND2_X1 U14723 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  XNOR2_X1 U14724 ( .A(n13408), .B(n11770), .ZN(n13637) );
  NAND2_X1 U14725 ( .A1(n13637), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11773) );
  INV_X1 U14726 ( .A(n11770), .ZN(n11771) );
  OR2_X1 U14727 ( .A1(n13408), .A2(n11771), .ZN(n11772) );
  NAND2_X1 U14728 ( .A1(n11773), .A2(n11772), .ZN(n11784) );
  INV_X1 U14729 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13109) );
  XNOR2_X1 U14730 ( .A(n11784), .B(n13109), .ZN(n13590) );
  OR2_X1 U14731 ( .A1(n11774), .A2(n11872), .ZN(n11783) );
  NAND2_X1 U14732 ( .A1(n11776), .A2(n11775), .ZN(n11777) );
  NAND2_X1 U14733 ( .A1(n11777), .A2(n11778), .ZN(n11796) );
  OAI21_X1 U14734 ( .B1(n11778), .B2(n11777), .A(n11796), .ZN(n11781) );
  INV_X1 U14735 ( .A(n11779), .ZN(n11780) );
  AOI21_X1 U14736 ( .B1(n11781), .B2(n11838), .A(n11780), .ZN(n11782) );
  NAND2_X1 U14737 ( .A1(n11783), .A2(n11782), .ZN(n13589) );
  NAND2_X1 U14738 ( .A1(n13590), .A2(n13589), .ZN(n11786) );
  NAND2_X1 U14739 ( .A1(n11784), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11785) );
  NAND2_X1 U14740 ( .A1(n11786), .A2(n11785), .ZN(n13674) );
  XNOR2_X1 U14741 ( .A(n11796), .B(n11787), .ZN(n11788) );
  NAND2_X1 U14742 ( .A1(n11788), .A2(n11838), .ZN(n11789) );
  INV_X1 U14743 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11790) );
  XNOR2_X1 U14744 ( .A(n11791), .B(n11790), .ZN(n13675) );
  NAND2_X1 U14745 ( .A1(n13674), .A2(n13675), .ZN(n11793) );
  NAND2_X1 U14746 ( .A1(n11791), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11792) );
  NAND2_X1 U14747 ( .A1(n11793), .A2(n11792), .ZN(n13770) );
  INV_X1 U14748 ( .A(n11872), .ZN(n11827) );
  NAND2_X1 U14749 ( .A1(n11794), .A2(n11827), .ZN(n11800) );
  NAND2_X1 U14750 ( .A1(n11796), .A2(n11795), .ZN(n11807) );
  XNOR2_X1 U14751 ( .A(n11807), .B(n11797), .ZN(n11798) );
  NAND2_X1 U14752 ( .A1(n11798), .A2(n11838), .ZN(n11799) );
  NAND2_X1 U14753 ( .A1(n11800), .A2(n11799), .ZN(n11802) );
  INV_X1 U14754 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11801) );
  XNOR2_X1 U14755 ( .A(n11802), .B(n11801), .ZN(n13769) );
  NAND2_X1 U14756 ( .A1(n13770), .A2(n13769), .ZN(n11804) );
  NAND2_X1 U14757 ( .A1(n11802), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11803) );
  NAND2_X1 U14758 ( .A1(n11804), .A2(n11803), .ZN(n13888) );
  NAND2_X1 U14759 ( .A1(n11805), .A2(n11827), .ZN(n11811) );
  OR2_X1 U14760 ( .A1(n11807), .A2(n11806), .ZN(n11819) );
  XNOR2_X1 U14761 ( .A(n11819), .B(n11808), .ZN(n11809) );
  NAND2_X1 U14762 ( .A1(n11809), .A2(n11838), .ZN(n11810) );
  NAND2_X1 U14763 ( .A1(n11811), .A2(n11810), .ZN(n11813) );
  INV_X1 U14764 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11812) );
  XNOR2_X1 U14765 ( .A(n11813), .B(n11812), .ZN(n13887) );
  NAND2_X1 U14766 ( .A1(n13888), .A2(n13887), .ZN(n11815) );
  NAND2_X1 U14767 ( .A1(n11813), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U14768 ( .A1(n11815), .A2(n11814), .ZN(n13942) );
  NAND3_X1 U14769 ( .A1(n11816), .A2(n11827), .A3(n11817), .ZN(n11823) );
  NOR2_X1 U14770 ( .A1(n11819), .A2(n11818), .ZN(n11821) );
  NAND2_X1 U14771 ( .A1(n11821), .A2(n11820), .ZN(n11836) );
  OAI211_X1 U14772 ( .C1(n11821), .C2(n11820), .A(n11836), .B(n11838), .ZN(
        n11822) );
  NAND2_X1 U14773 ( .A1(n11823), .A2(n11822), .ZN(n11825) );
  INV_X1 U14774 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11824) );
  XNOR2_X1 U14775 ( .A(n11825), .B(n11824), .ZN(n13941) );
  NAND2_X1 U14776 ( .A1(n11825), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11826) );
  NAND2_X1 U14777 ( .A1(n11828), .A2(n11827), .ZN(n11831) );
  XNOR2_X1 U14778 ( .A(n11836), .B(n11837), .ZN(n11829) );
  NAND2_X1 U14779 ( .A1(n11829), .A2(n11838), .ZN(n11830) );
  NAND2_X1 U14780 ( .A1(n11831), .A2(n11830), .ZN(n11832) );
  OR2_X1 U14781 ( .A1(n11832), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15948) );
  NAND2_X1 U14782 ( .A1(n11832), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15947) );
  NOR3_X1 U14783 ( .A1(n11834), .A2(n11872), .A3(n11833), .ZN(n11835) );
  NAND2_X2 U14784 ( .A1(n11816), .A2(n11835), .ZN(n11856) );
  INV_X1 U14785 ( .A(n11836), .ZN(n11839) );
  NAND3_X1 U14786 ( .A1(n11839), .A2(n11838), .A3(n11837), .ZN(n11840) );
  NAND2_X1 U14787 ( .A1(n15908), .A2(n11840), .ZN(n14134) );
  OR2_X1 U14788 ( .A1(n14134), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11841) );
  NAND2_X1 U14789 ( .A1(n14136), .A2(n11841), .ZN(n11843) );
  NAND2_X1 U14790 ( .A1(n14134), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11842) );
  NAND2_X1 U14791 ( .A1(n11843), .A2(n11842), .ZN(n14217) );
  INV_X1 U14792 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11845) );
  NOR2_X1 U14793 ( .A1(n15908), .A2(n11845), .ZN(n11844) );
  NAND2_X1 U14794 ( .A1(n15908), .A2(n11845), .ZN(n14216) );
  XNOR2_X1 U14795 ( .A(n11856), .B(n14794), .ZN(n14671) );
  INV_X1 U14796 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14270) );
  NAND2_X1 U14797 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11846) );
  AND2_X1 U14798 ( .A1(n11856), .A2(n11846), .ZN(n14262) );
  INV_X1 U14799 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14775) );
  AND2_X1 U14800 ( .A1(n15908), .A2(n14775), .ZN(n11847) );
  XNOR2_X1 U14801 ( .A(n15908), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14654) );
  INV_X1 U14802 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16025) );
  NAND2_X1 U14803 ( .A1(n15908), .A2(n16025), .ZN(n15930) );
  OAI211_X1 U14804 ( .C1(n15918), .C2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n14654), .B(n15930), .ZN(n11848) );
  NOR2_X1 U14805 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11849) );
  NAND2_X1 U14806 ( .A1(n15927), .A2(n15931), .ZN(n14653) );
  NOR2_X1 U14807 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11851) );
  NOR2_X1 U14808 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14263) );
  AND2_X1 U14809 ( .A1(n14263), .A2(n14270), .ZN(n11850) );
  OAI21_X1 U14810 ( .B1(n11851), .B2(n15908), .A(n14668), .ZN(n11852) );
  INV_X1 U14811 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16006) );
  INV_X1 U14812 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14782) );
  INV_X1 U14813 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11853) );
  NAND2_X1 U14814 ( .A1(n15734), .A2(n11853), .ZN(n11854) );
  XNOR2_X1 U14815 ( .A(n15908), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14646) );
  NAND2_X2 U14816 ( .A1(n14647), .A2(n14646), .ZN(n15909) );
  AND2_X1 U14817 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15732) );
  NAND2_X1 U14818 ( .A1(n15732), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14695) );
  OAI21_X2 U14819 ( .B1(n15909), .B2(n14695), .A(n15908), .ZN(n14629) );
  NOR2_X1 U14820 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14591) );
  INV_X1 U14821 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14594) );
  INV_X1 U14822 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14722) );
  NAND2_X1 U14823 ( .A1(n14563), .A2(n14722), .ZN(n14557) );
  AND3_X1 U14824 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14703) );
  NAND2_X1 U14825 ( .A1(n14703), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11855) );
  AND2_X1 U14826 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14710) );
  NAND2_X1 U14827 ( .A1(n14581), .A2(n14710), .ZN(n14562) );
  INV_X1 U14828 ( .A(n14562), .ZN(n11857) );
  NAND3_X1 U14829 ( .A1(n11857), .A2(n11856), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14556) );
  NAND2_X1 U14830 ( .A1(n20259), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11860) );
  NAND2_X1 U14831 ( .A1(n14810), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11859) );
  NAND2_X1 U14832 ( .A1(n11860), .A2(n11859), .ZN(n11881) );
  NAND2_X1 U14833 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20610), .ZN(
        n11880) );
  NAND2_X1 U14834 ( .A1(n11861), .A2(n11860), .ZN(n11889) );
  OR2_X1 U14835 ( .A1(n13751), .A2(n20573), .ZN(n11862) );
  NAND2_X1 U14836 ( .A1(n11889), .A2(n11862), .ZN(n11864) );
  NAND2_X1 U14837 ( .A1(n20573), .A2(n13751), .ZN(n11863) );
  MUX2_X1 U14838 ( .A(n15688), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11873) );
  NOR2_X1 U14839 ( .A1(n11865), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11866) );
  NAND2_X1 U14840 ( .A1(n20157), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11867) );
  NAND2_X1 U14841 ( .A1(n11871), .A2(n11867), .ZN(n11869) );
  NAND2_X1 U14842 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16077), .ZN(
        n11868) );
  NOR2_X1 U14843 ( .A1(n20157), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11870) );
  XNOR2_X1 U14844 ( .A(n11874), .B(n11873), .ZN(n13255) );
  INV_X1 U14845 ( .A(n11884), .ZN(n11882) );
  INV_X1 U14846 ( .A(n11904), .ZN(n13261) );
  NOR3_X1 U14847 ( .A1(n11882), .A2(n20183), .A3(n13261), .ZN(n11901) );
  OAI21_X1 U14848 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20610), .A(
        n11880), .ZN(n11876) );
  INV_X1 U14849 ( .A(n11876), .ZN(n11875) );
  OAI21_X1 U14850 ( .B1(n10166), .B2(n9812), .A(n11875), .ZN(n11878) );
  AND2_X1 U14851 ( .A1(n20183), .A2(n11031), .ZN(n11879) );
  NOR2_X1 U14852 ( .A1(n11907), .A2(n11876), .ZN(n11877) );
  OAI22_X1 U14853 ( .A1(n11878), .A2(n11897), .B1(n11909), .B2(n11877), .ZN(
        n11887) );
  INV_X1 U14854 ( .A(n11879), .ZN(n11883) );
  XNOR2_X1 U14855 ( .A(n11881), .B(n11880), .ZN(n13256) );
  AOI22_X1 U14856 ( .A1(n11883), .A2(n11882), .B1(n11890), .B2(n13256), .ZN(
        n11886) );
  NAND2_X1 U14857 ( .A1(n11884), .A2(n11036), .ZN(n11885) );
  AOI22_X1 U14858 ( .A1(n11887), .A2(n11886), .B1(n11885), .B2(n13256), .ZN(
        n11894) );
  NOR2_X1 U14859 ( .A1(n11887), .A2(n11886), .ZN(n11893) );
  MUX2_X1 U14860 ( .A(n20573), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n13751), .Z(n11888) );
  XNOR2_X1 U14861 ( .A(n11889), .B(n11888), .ZN(n13257) );
  AOI21_X1 U14862 ( .B1(n11890), .B2(n13257), .A(n11897), .ZN(n11891) );
  OAI21_X1 U14863 ( .B1(n11907), .B2(n13257), .A(n11891), .ZN(n11892) );
  OAI21_X1 U14864 ( .B1(n11894), .B2(n11893), .A(n11892), .ZN(n11899) );
  INV_X1 U14865 ( .A(n13257), .ZN(n11896) );
  NAND3_X1 U14866 ( .A1(n11897), .A2(n11896), .A3(n11895), .ZN(n11898) );
  AOI22_X1 U14867 ( .A1(n11899), .A2(n11898), .B1(n11903), .B2(n13255), .ZN(
        n11900) );
  AOI211_X1 U14868 ( .C1(n11909), .C2(n13255), .A(n11901), .B(n11900), .ZN(
        n11902) );
  AOI21_X1 U14869 ( .B1(n11904), .B2(n11903), .A(n11902), .ZN(n11905) );
  NAND2_X1 U14870 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  AND2_X1 U14871 ( .A1(n14806), .A2(n9812), .ZN(n11915) );
  NAND2_X1 U14872 ( .A1(n11912), .A2(n20215), .ZN(n11913) );
  NAND2_X1 U14873 ( .A1(n11914), .A2(n11913), .ZN(n13383) );
  OR2_X1 U14874 ( .A1(n11915), .A2(n13383), .ZN(n13376) );
  NOR2_X1 U14875 ( .A1(n13376), .A2(n10166), .ZN(n15696) );
  NAND2_X1 U14876 ( .A1(n15707), .A2(n15696), .ZN(n15714) );
  NAND2_X1 U14877 ( .A1(n20540), .A2(n11917), .ZN(n20816) );
  NAND2_X1 U14878 ( .A1(n20816), .A2(n20169), .ZN(n11916) );
  OR2_X2 U14879 ( .A1(n11917), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20055) );
  INV_X1 U14880 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21183) );
  NOR2_X1 U14881 ( .A1(n20055), .A2(n21183), .ZN(n14698) );
  NAND2_X1 U14882 ( .A1(n20169), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15722) );
  NAND2_X1 U14883 ( .A1(n21140), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11918) );
  AND2_X1 U14884 ( .A1(n15722), .A2(n11918), .ZN(n13407) );
  INV_X1 U14885 ( .A(n13407), .ZN(n11919) );
  INV_X1 U14886 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14553) );
  INV_X1 U14887 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11921) );
  NOR2_X1 U14888 ( .A1(n15954), .A2(n14005), .ZN(n11923) );
  AOI211_X1 U14889 ( .C1(n15946), .C2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14698), .B(n11923), .ZN(n11924) );
  XNOR2_X2 U14890 ( .A(n11962), .B(n11926), .ZN(n12307) );
  NAND2_X1 U14891 ( .A1(n19283), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11927) );
  NOR2_X2 U14892 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19945) );
  NAND2_X1 U14893 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19617) );
  NAND2_X1 U14894 ( .A1(n19617), .A2(n19968), .ZN(n11928) );
  NOR2_X1 U14895 ( .A1(n19968), .A2(n19978), .ZN(n19745) );
  NAND2_X1 U14896 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19745), .ZN(
        n14100) );
  AND2_X1 U14897 ( .A1(n11928), .A2(n14100), .ZN(n19395) );
  AOI22_X1 U14898 ( .A1(n11968), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19945), .B2(n19395), .ZN(n11929) );
  NAND3_X1 U14899 ( .A1(n13668), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19264), 
        .ZN(n13500) );
  INV_X1 U14900 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19272) );
  NOR2_X1 U14901 ( .A1(n13500), .A2(n19272), .ZN(n11931) );
  NAND2_X1 U14902 ( .A1(n11932), .A2(n11931), .ZN(n11946) );
  INV_X1 U14903 ( .A(n13361), .ZN(n11949) );
  OR2_X1 U14904 ( .A1(n11934), .A2(n11933), .ZN(n11935) );
  AOI22_X1 U14905 ( .A1(n11968), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19945), .B2(n19987), .ZN(n11936) );
  INV_X1 U14906 ( .A(n13500), .ZN(n12159) );
  NAND2_X1 U14907 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11943) );
  NAND2_X1 U14908 ( .A1(n11968), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U14909 ( .A1(n19987), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11940) );
  NAND2_X1 U14910 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19978), .ZN(
        n19559) );
  NAND2_X1 U14911 ( .A1(n11940), .A2(n19559), .ZN(n19394) );
  NAND2_X1 U14912 ( .A1(n19945), .A2(n19394), .ZN(n19591) );
  NAND2_X1 U14913 ( .A1(n11941), .A2(n19591), .ZN(n11942) );
  NAND2_X1 U14914 ( .A1(n13335), .A2(n13334), .ZN(n11945) );
  INV_X1 U14915 ( .A(n13342), .ZN(n15566) );
  NAND2_X1 U14916 ( .A1(n15566), .A2(n11943), .ZN(n11944) );
  INV_X1 U14917 ( .A(n11950), .ZN(n11952) );
  NOR2_X1 U14918 ( .A1(n11953), .A2(n11952), .ZN(n11956) );
  INV_X1 U14919 ( .A(n11956), .ZN(n11951) );
  NAND2_X1 U14920 ( .A1(n11957), .A2(n11951), .ZN(n11963) );
  NAND2_X1 U14921 ( .A1(n11953), .A2(n11952), .ZN(n11955) );
  INV_X1 U14922 ( .A(n11957), .ZN(n11954) );
  NAND3_X1 U14923 ( .A1(n11962), .A2(n11955), .A3(n11954), .ZN(n11961) );
  OR2_X2 U14924 ( .A1(n11957), .A2(n11956), .ZN(n11958) );
  INV_X1 U14925 ( .A(n11964), .ZN(n12673) );
  NAND2_X1 U14926 ( .A1(n19745), .A2(n19960), .ZN(n19497) );
  INV_X1 U14927 ( .A(n19497), .ZN(n11965) );
  INV_X1 U14928 ( .A(n19530), .ZN(n19527) );
  NAND2_X1 U14929 ( .A1(n14100), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11966) );
  NAND2_X1 U14930 ( .A1(n19527), .A2(n11966), .ZN(n11967) );
  AND2_X1 U14931 ( .A1(n11967), .A2(n19945), .ZN(n19674) );
  AOI21_X1 U14932 ( .B1(n11968), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19674), .ZN(n11969) );
  NAND2_X1 U14933 ( .A1(n11971), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11970) );
  INV_X1 U14934 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14118) );
  NOR2_X1 U14935 ( .A1(n13500), .A2(n14118), .ZN(n13415) );
  AND3_X1 U14936 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__5__SCAN_IN), 
        .ZN(n11972) );
  INV_X1 U14937 ( .A(n13580), .ZN(n11975) );
  INV_X1 U14938 ( .A(n13684), .ZN(n11974) );
  AOI22_X1 U14939 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U14940 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U14941 ( .A1(n10751), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U14942 ( .A1(n12031), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11976) );
  NAND4_X1 U14943 ( .A1(n11979), .A2(n11978), .A3(n11977), .A4(n11976), .ZN(
        n11985) );
  AOI22_X1 U14944 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U14945 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U14946 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U14947 ( .A1(n10635), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11980) );
  NAND4_X1 U14948 ( .A1(n11983), .A2(n11982), .A3(n11981), .A4(n11980), .ZN(
        n11984) );
  OR2_X1 U14949 ( .A1(n11985), .A2(n11984), .ZN(n14122) );
  INV_X1 U14950 ( .A(n14160), .ZN(n11987) );
  NOR2_X1 U14951 ( .A1(n14055), .A2(n11986), .ZN(n14079) );
  AND2_X1 U14952 ( .A1(n11987), .A2(n14079), .ZN(n14119) );
  AOI22_X1 U14953 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U14954 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U14955 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U14956 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12031), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11990) );
  NAND4_X1 U14957 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n11999) );
  AOI22_X1 U14958 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U14959 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U14960 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U14961 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11994) );
  NAND4_X1 U14962 ( .A1(n11997), .A2(n11996), .A3(n11995), .A4(n11994), .ZN(
        n11998) );
  AOI22_X1 U14963 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U14964 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U14965 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U14966 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12031), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12000) );
  NAND4_X1 U14967 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(
        n12010) );
  AOI22_X1 U14968 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U14969 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U14970 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U14971 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12005) );
  NAND4_X1 U14972 ( .A1(n12008), .A2(n12007), .A3(n12006), .A4(n12005), .ZN(
        n12009) );
  NOR2_X1 U14973 ( .A1(n12010), .A2(n12009), .ZN(n14982) );
  AOI22_X1 U14974 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U14975 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U14976 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U14977 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12031), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12011) );
  NAND4_X1 U14978 ( .A1(n12014), .A2(n12013), .A3(n12012), .A4(n12011), .ZN(
        n12020) );
  AOI22_X1 U14979 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U14980 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U14981 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U14982 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12015) );
  NAND4_X1 U14983 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n12019) );
  OR2_X1 U14984 ( .A1(n12020), .A2(n12019), .ZN(n14975) );
  AOI22_X1 U14985 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U14986 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U14987 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U14988 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12031), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12021) );
  NAND4_X1 U14989 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12030) );
  AOI22_X1 U14990 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U14991 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U14992 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U14993 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12025) );
  NAND4_X1 U14994 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12029) );
  OR2_X1 U14995 ( .A1(n12030), .A2(n12029), .ZN(n14968) );
  NAND2_X1 U14996 ( .A1(n14969), .A2(n14968), .ZN(n14956) );
  AOI22_X1 U14997 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12073), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U14998 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U14999 ( .A1(n10751), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15000 ( .A1(n12031), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12032) );
  NAND4_X1 U15001 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12032), .ZN(
        n12041) );
  AOI22_X1 U15002 ( .A1(n10634), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15003 ( .A1(n10636), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10693), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15004 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15005 ( .A1(n10635), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12036) );
  NAND4_X1 U15006 ( .A1(n12039), .A2(n12038), .A3(n12037), .A4(n12036), .ZN(
        n12040) );
  AOI22_X1 U15007 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12073), .B1(
        n10670), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15008 ( .A1(n10647), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15009 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15010 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12031), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12042) );
  NAND4_X1 U15011 ( .A1(n12045), .A2(n12044), .A3(n12043), .A4(n12042), .ZN(
        n12051) );
  AOI22_X1 U15012 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15013 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15014 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U15015 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12046) );
  NAND4_X1 U15016 ( .A1(n12049), .A2(n12048), .A3(n12047), .A4(n12046), .ZN(
        n12050) );
  NOR2_X1 U15017 ( .A1(n12051), .A2(n12050), .ZN(n14951) );
  INV_X1 U15018 ( .A(n10387), .ZN(n12211) );
  INV_X1 U15019 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12052) );
  INV_X1 U15020 ( .A(n12243), .ZN(n12218) );
  INV_X1 U15021 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19470) );
  OAI22_X1 U15022 ( .A1(n12211), .A2(n12052), .B1(n12218), .B2(n19470), .ZN(
        n12057) );
  INV_X1 U15023 ( .A(n12244), .ZN(n12223) );
  INV_X1 U15024 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12055) );
  INV_X1 U15025 ( .A(n12053), .ZN(n12222) );
  INV_X1 U15026 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12054) );
  OAI22_X1 U15027 ( .A1(n12223), .A2(n12055), .B1(n12222), .B2(n12054), .ZN(
        n12056) );
  NOR2_X1 U15028 ( .A1(n12057), .A2(n12056), .ZN(n12061) );
  AOI22_X1 U15029 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15030 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12059) );
  XNOR2_X1 U15031 ( .A(n16325), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12246) );
  INV_X1 U15032 ( .A(n12246), .ZN(n12238) );
  NAND4_X1 U15033 ( .A1(n12061), .A2(n12060), .A3(n12059), .A4(n12238), .ZN(
        n12072) );
  INV_X1 U15034 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12063) );
  INV_X1 U15035 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12062) );
  OAI22_X1 U15036 ( .A1(n12211), .A2(n12063), .B1(n12223), .B2(n12062), .ZN(
        n12067) );
  INV_X1 U15037 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12065) );
  INV_X1 U15038 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12064) );
  OAI22_X1 U15039 ( .A1(n12222), .A2(n12065), .B1(n12218), .B2(n12064), .ZN(
        n12066) );
  NOR2_X1 U15040 ( .A1(n12067), .A2(n12066), .ZN(n12070) );
  AOI22_X1 U15041 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9802), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15042 ( .A1(n12235), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12068) );
  NAND4_X1 U15043 ( .A1(n12070), .A2(n12246), .A3(n12069), .A4(n12068), .ZN(
        n12071) );
  NAND2_X1 U15044 ( .A1(n12072), .A2(n12071), .ZN(n12110) );
  NOR2_X1 U15045 ( .A1(n13446), .A2(n12110), .ZN(n12084) );
  AOI22_X1 U15046 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10670), .B1(
        n10647), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15047 ( .A1(n12073), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10648), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15048 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10751), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15049 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12031), .B1(
        n11989), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12074) );
  NAND4_X1 U15050 ( .A1(n12077), .A2(n12076), .A3(n12075), .A4(n12074), .ZN(
        n12083) );
  AOI22_X1 U15051 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10635), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15052 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10634), .B1(
        n10692), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15053 ( .A1(n10616), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12004), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15054 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10693), .B1(
        n10636), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12078) );
  NAND4_X1 U15055 ( .A1(n12081), .A2(n12080), .A3(n12079), .A4(n12078), .ZN(
        n12082) );
  NOR2_X1 U15056 ( .A1(n12083), .A2(n12082), .ZN(n12104) );
  XNOR2_X1 U15057 ( .A(n12084), .B(n12104), .ZN(n12108) );
  INV_X1 U15058 ( .A(n12110), .ZN(n12105) );
  NAND2_X1 U15059 ( .A1(n13446), .A2(n12105), .ZN(n14940) );
  NOR2_X2 U15060 ( .A1(n14939), .A2(n12086), .ZN(n14932) );
  INV_X1 U15061 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12347) );
  INV_X1 U15062 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12087) );
  OAI22_X1 U15063 ( .A1(n12211), .A2(n12347), .B1(n12218), .B2(n12087), .ZN(
        n12089) );
  INV_X1 U15064 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12348) );
  INV_X1 U15065 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12349) );
  OAI22_X1 U15066 ( .A1(n12223), .A2(n12348), .B1(n12222), .B2(n12349), .ZN(
        n12088) );
  NOR2_X1 U15067 ( .A1(n12089), .A2(n12088), .ZN(n12092) );
  AOI22_X1 U15068 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15069 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12090) );
  NAND4_X1 U15070 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12238), .ZN(
        n12103) );
  INV_X1 U15071 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12094) );
  INV_X1 U15072 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12093) );
  OAI22_X1 U15073 ( .A1(n12211), .A2(n12094), .B1(n12218), .B2(n12093), .ZN(
        n12098) );
  INV_X1 U15074 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12096) );
  INV_X1 U15075 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12095) );
  OAI22_X1 U15076 ( .A1(n12223), .A2(n12096), .B1(n12222), .B2(n12095), .ZN(
        n12097) );
  NOR2_X1 U15077 ( .A1(n12098), .A2(n12097), .ZN(n12101) );
  AOI22_X1 U15078 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15079 ( .A1(n9801), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U15080 ( .A1(n12101), .A2(n12246), .A3(n12100), .A4(n12099), .ZN(
        n12102) );
  NAND2_X1 U15081 ( .A1(n12103), .A2(n12102), .ZN(n12112) );
  INV_X1 U15082 ( .A(n12104), .ZN(n12106) );
  NAND2_X1 U15083 ( .A1(n12106), .A2(n12105), .ZN(n12113) );
  XOR2_X1 U15084 ( .A(n12112), .B(n12113), .Z(n12107) );
  NAND2_X1 U15085 ( .A1(n12107), .A2(n12159), .ZN(n14934) );
  INV_X1 U15086 ( .A(n12112), .ZN(n12109) );
  NAND2_X1 U15087 ( .A1(n13446), .A2(n12109), .ZN(n14936) );
  NOR3_X1 U15088 ( .A1(n10220), .A2(n12110), .A3(n14936), .ZN(n12111) );
  NOR2_X1 U15089 ( .A1(n12113), .A2(n12112), .ZN(n12134) );
  INV_X1 U15090 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12115) );
  INV_X1 U15091 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12114) );
  OAI22_X1 U15092 ( .A1(n12211), .A2(n12115), .B1(n12218), .B2(n12114), .ZN(
        n12119) );
  INV_X1 U15093 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12117) );
  INV_X1 U15094 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12116) );
  OAI22_X1 U15095 ( .A1(n12223), .A2(n12117), .B1(n12222), .B2(n12116), .ZN(
        n12118) );
  NOR2_X1 U15096 ( .A1(n12119), .A2(n12118), .ZN(n12122) );
  AOI22_X1 U15097 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15098 ( .A1(n9801), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15099 ( .A1(n12122), .A2(n12121), .A3(n12120), .A4(n12238), .ZN(
        n12133) );
  INV_X1 U15100 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12124) );
  INV_X1 U15101 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12123) );
  OAI22_X1 U15102 ( .A1(n12211), .A2(n12124), .B1(n12218), .B2(n12123), .ZN(
        n12128) );
  INV_X1 U15103 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12126) );
  INV_X1 U15104 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12125) );
  OAI22_X1 U15105 ( .A1(n12223), .A2(n12126), .B1(n12222), .B2(n12125), .ZN(
        n12127) );
  NOR2_X1 U15106 ( .A1(n12128), .A2(n12127), .ZN(n12131) );
  AOI22_X1 U15107 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15108 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12129) );
  NAND4_X1 U15109 ( .A1(n12131), .A2(n12246), .A3(n12130), .A4(n12129), .ZN(
        n12132) );
  AND2_X1 U15110 ( .A1(n12133), .A2(n12132), .ZN(n12136) );
  NAND2_X1 U15111 ( .A1(n12134), .A2(n12136), .ZN(n12186) );
  OAI211_X1 U15112 ( .C1(n12134), .C2(n12136), .A(n12159), .B(n12186), .ZN(
        n12139) );
  INV_X1 U15113 ( .A(n12139), .ZN(n12135) );
  XNOR2_X1 U15114 ( .A(n12138), .B(n12135), .ZN(n14924) );
  INV_X1 U15115 ( .A(n12136), .ZN(n12137) );
  NOR2_X1 U15116 ( .A1(n19264), .A2(n12137), .ZN(n14926) );
  NAND2_X1 U15117 ( .A1(n14924), .A2(n14926), .ZN(n14925) );
  INV_X1 U15118 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12142) );
  INV_X1 U15119 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12141) );
  OAI22_X1 U15120 ( .A1(n12211), .A2(n12142), .B1(n12218), .B2(n12141), .ZN(
        n12144) );
  INV_X1 U15121 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12317) );
  INV_X1 U15122 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12318) );
  OAI22_X1 U15123 ( .A1(n12223), .A2(n12317), .B1(n12222), .B2(n12318), .ZN(
        n12143) );
  NOR2_X1 U15124 ( .A1(n12144), .A2(n12143), .ZN(n12147) );
  AOI22_X1 U15125 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15126 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12145) );
  NAND4_X1 U15127 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12238), .ZN(
        n12158) );
  INV_X1 U15128 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12149) );
  INV_X1 U15129 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12148) );
  OAI22_X1 U15130 ( .A1(n12211), .A2(n12149), .B1(n12218), .B2(n12148), .ZN(
        n12153) );
  INV_X1 U15131 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12151) );
  INV_X1 U15132 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12150) );
  OAI22_X1 U15133 ( .A1(n12223), .A2(n12151), .B1(n12222), .B2(n12150), .ZN(
        n12152) );
  NOR2_X1 U15134 ( .A1(n12153), .A2(n12152), .ZN(n12156) );
  AOI22_X1 U15135 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15136 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12154) );
  NAND4_X1 U15137 ( .A1(n12156), .A2(n12246), .A3(n12155), .A4(n12154), .ZN(
        n12157) );
  AND2_X1 U15138 ( .A1(n12158), .A2(n12157), .ZN(n12161) );
  XNOR2_X1 U15139 ( .A(n12186), .B(n12161), .ZN(n12160) );
  NAND2_X1 U15140 ( .A1(n12160), .A2(n12159), .ZN(n12163) );
  INV_X1 U15141 ( .A(n12161), .ZN(n12185) );
  NOR2_X1 U15142 ( .A1(n19264), .A2(n12185), .ZN(n14917) );
  NAND2_X1 U15143 ( .A1(n14918), .A2(n14917), .ZN(n14916) );
  INV_X1 U15144 ( .A(n12162), .ZN(n12164) );
  NAND2_X1 U15145 ( .A1(n14916), .A2(n9862), .ZN(n12189) );
  INV_X1 U15146 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12166) );
  INV_X1 U15147 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12165) );
  OAI22_X1 U15148 ( .A1(n12211), .A2(n12166), .B1(n12218), .B2(n12165), .ZN(
        n12170) );
  INV_X1 U15149 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12168) );
  INV_X1 U15150 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12167) );
  OAI22_X1 U15151 ( .A1(n12223), .A2(n12168), .B1(n12222), .B2(n12167), .ZN(
        n12169) );
  NOR2_X1 U15152 ( .A1(n12170), .A2(n12169), .ZN(n12173) );
  AOI22_X1 U15153 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15154 ( .A1(n9801), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12171) );
  NAND4_X1 U15155 ( .A1(n12173), .A2(n12172), .A3(n12171), .A4(n12238), .ZN(
        n12184) );
  INV_X1 U15156 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12175) );
  INV_X1 U15157 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12174) );
  OAI22_X1 U15158 ( .A1(n12211), .A2(n12175), .B1(n12218), .B2(n12174), .ZN(
        n12179) );
  INV_X1 U15159 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12177) );
  INV_X1 U15160 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12176) );
  OAI22_X1 U15161 ( .A1(n12223), .A2(n12177), .B1(n12222), .B2(n12176), .ZN(
        n12178) );
  NOR2_X1 U15162 ( .A1(n12179), .A2(n12178), .ZN(n12182) );
  AOI22_X1 U15163 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15164 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12180) );
  NAND4_X1 U15165 ( .A1(n12182), .A2(n12246), .A3(n12181), .A4(n12180), .ZN(
        n12183) );
  NAND2_X1 U15166 ( .A1(n12184), .A2(n12183), .ZN(n12191) );
  OR2_X1 U15167 ( .A1(n12186), .A2(n12185), .ZN(n12187) );
  NOR2_X1 U15168 ( .A1(n12187), .A2(n12191), .ZN(n12208) );
  AOI211_X1 U15169 ( .C1(n12191), .C2(n12187), .A(n13500), .B(n12208), .ZN(
        n12188) );
  NAND2_X1 U15170 ( .A1(n12189), .A2(n12188), .ZN(n12193) );
  OR2_X1 U15171 ( .A1(n12189), .A2(n12188), .ZN(n12190) );
  NAND2_X1 U15172 ( .A1(n12193), .A2(n12190), .ZN(n14913) );
  INV_X1 U15173 ( .A(n12191), .ZN(n12192) );
  NAND2_X1 U15174 ( .A1(n13446), .A2(n12192), .ZN(n14912) );
  NOR2_X1 U15175 ( .A1(n14913), .A2(n14912), .ZN(n14911) );
  INV_X1 U15176 ( .A(n12193), .ZN(n12207) );
  INV_X1 U15177 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12367) );
  INV_X1 U15178 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12382) );
  OAI22_X1 U15179 ( .A1(n12211), .A2(n12367), .B1(n12218), .B2(n12382), .ZN(
        n12195) );
  INV_X1 U15180 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12371) );
  INV_X1 U15181 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12369) );
  OAI22_X1 U15182 ( .A1(n12223), .A2(n12371), .B1(n12222), .B2(n12369), .ZN(
        n12194) );
  NOR2_X1 U15183 ( .A1(n12195), .A2(n12194), .ZN(n12198) );
  AOI22_X1 U15184 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15185 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12196) );
  NAND4_X1 U15186 ( .A1(n12198), .A2(n12197), .A3(n12196), .A4(n12238), .ZN(
        n12206) );
  INV_X1 U15187 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12199) );
  INV_X1 U15188 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12384) );
  OAI22_X1 U15189 ( .A1(n12211), .A2(n12199), .B1(n12218), .B2(n12384), .ZN(
        n12201) );
  INV_X1 U15190 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12387) );
  INV_X1 U15191 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12385) );
  OAI22_X1 U15192 ( .A1(n12223), .A2(n12387), .B1(n12222), .B2(n12385), .ZN(
        n12200) );
  NOR2_X1 U15193 ( .A1(n12201), .A2(n12200), .ZN(n12204) );
  AOI22_X1 U15194 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15195 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12202) );
  NAND4_X1 U15196 ( .A1(n12204), .A2(n12246), .A3(n12203), .A4(n12202), .ZN(
        n12205) );
  AND2_X1 U15197 ( .A1(n12206), .A2(n12205), .ZN(n14904) );
  OAI21_X1 U15198 ( .B1(n14911), .B2(n12207), .A(n14904), .ZN(n14899) );
  INV_X1 U15199 ( .A(n12208), .ZN(n14903) );
  NAND2_X1 U15200 ( .A1(n19264), .A2(n14904), .ZN(n12209) );
  NOR2_X1 U15201 ( .A1(n14903), .A2(n12209), .ZN(n12232) );
  INV_X1 U15202 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12210) );
  INV_X1 U15203 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12443) );
  OAI22_X1 U15204 ( .A1(n12211), .A2(n12210), .B1(n12222), .B2(n12443), .ZN(
        n12213) );
  INV_X1 U15205 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12444) );
  INV_X1 U15206 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12432) );
  OAI22_X1 U15207 ( .A1(n12223), .A2(n12444), .B1(n12218), .B2(n12432), .ZN(
        n12212) );
  NOR2_X1 U15208 ( .A1(n12213), .A2(n12212), .ZN(n12216) );
  AOI22_X1 U15209 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15210 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12214) );
  NAND4_X1 U15211 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12238), .ZN(
        n12230) );
  INV_X1 U15212 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12219) );
  INV_X1 U15213 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12217) );
  OAI22_X1 U15214 ( .A1(n9816), .A2(n12219), .B1(n12218), .B2(n12217), .ZN(
        n12225) );
  INV_X1 U15215 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12433) );
  INV_X1 U15216 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12221) );
  OAI22_X1 U15217 ( .A1(n12223), .A2(n12433), .B1(n12222), .B2(n12221), .ZN(
        n12224) );
  NOR2_X1 U15218 ( .A1(n12225), .A2(n12224), .ZN(n12228) );
  AOI22_X1 U15219 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15220 ( .A1(n9801), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12226) );
  NAND4_X1 U15221 ( .A1(n12228), .A2(n12246), .A3(n12227), .A4(n12226), .ZN(
        n12229) );
  AND2_X1 U15222 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  NAND2_X1 U15223 ( .A1(n12232), .A2(n12231), .ZN(n12233) );
  OAI21_X1 U15224 ( .B1(n12232), .B2(n12231), .A(n12233), .ZN(n14900) );
  NOR2_X1 U15225 ( .A1(n14899), .A2(n14900), .ZN(n14898) );
  INV_X1 U15226 ( .A(n12233), .ZN(n12234) );
  NOR2_X1 U15227 ( .A1(n14898), .A2(n12234), .ZN(n12254) );
  AOI22_X1 U15228 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15229 ( .A1(n12235), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12236) );
  NAND2_X1 U15230 ( .A1(n12237), .A2(n12236), .ZN(n12252) );
  AOI22_X1 U15231 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15232 ( .A1(n12245), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12239) );
  NAND3_X1 U15233 ( .A1(n12240), .A2(n12239), .A3(n12238), .ZN(n12251) );
  AOI22_X1 U15234 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12235), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15235 ( .A1(n9801), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10593), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12241) );
  NAND2_X1 U15236 ( .A1(n12242), .A2(n12241), .ZN(n12250) );
  AOI22_X1 U15237 ( .A1(n10387), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12243), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15238 ( .A1(n12245), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12244), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12247) );
  NAND3_X1 U15239 ( .A1(n12248), .A2(n12247), .A3(n12246), .ZN(n12249) );
  OAI22_X1 U15240 ( .A1(n12252), .A2(n12251), .B1(n12250), .B2(n12249), .ZN(
        n12253) );
  XNOR2_X1 U15241 ( .A(n12254), .B(n12253), .ZN(n14322) );
  INV_X1 U15242 ( .A(n12255), .ZN(n12607) );
  NAND2_X1 U15243 ( .A1(n15562), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12256) );
  AND2_X1 U15244 ( .A1(n12257), .A2(n12256), .ZN(n12259) );
  INV_X1 U15245 ( .A(n12259), .ZN(n12600) );
  NOR2_X1 U15246 ( .A1(n12607), .A2(n12600), .ZN(n12261) );
  OAI211_X1 U15247 ( .C1(n19264), .C2(n12259), .A(n13048), .B(n12258), .ZN(
        n12260) );
  OAI21_X1 U15248 ( .B1(n13035), .B2(n12261), .A(n12260), .ZN(n12262) );
  NAND2_X1 U15249 ( .A1(n12270), .A2(n12262), .ZN(n12263) );
  OAI21_X1 U15250 ( .B1(n12601), .B2(n13224), .A(n12263), .ZN(n12268) );
  NAND2_X1 U15251 ( .A1(n14818), .A2(n19264), .ZN(n12266) );
  INV_X1 U15252 ( .A(n12264), .ZN(n12265) );
  MUX2_X1 U15253 ( .A(n13035), .B(n12266), .S(n12265), .Z(n12267) );
  NAND2_X1 U15254 ( .A1(n12268), .A2(n12267), .ZN(n12269) );
  OAI21_X1 U15255 ( .B1(n12270), .B2(n13035), .A(n12269), .ZN(n12271) );
  OR2_X1 U15256 ( .A1(n12271), .A2(n12612), .ZN(n12272) );
  MUX2_X1 U15257 ( .A(n12272), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18906), .Z(n13021) );
  NAND2_X1 U15258 ( .A1(n12612), .A2(n12273), .ZN(n12274) );
  NAND2_X1 U15259 ( .A1(n13446), .A2(n10333), .ZN(n12281) );
  NAND2_X1 U15260 ( .A1(n12281), .A2(n13048), .ZN(n12275) );
  NAND3_X1 U15261 ( .A1(n12275), .A2(n13047), .A3(n19292), .ZN(n12280) );
  NAND2_X1 U15262 ( .A1(n12276), .A2(n19292), .ZN(n12277) );
  NAND2_X1 U15263 ( .A1(n12277), .A2(n16362), .ZN(n13045) );
  NAND2_X1 U15264 ( .A1(n13045), .A2(n12278), .ZN(n12279) );
  AOI21_X1 U15265 ( .B1(n13231), .B2(n12280), .A(n12279), .ZN(n13025) );
  NOR2_X1 U15266 ( .A1(n10409), .A2(n12281), .ZN(n12282) );
  AND2_X1 U15267 ( .A1(n12283), .A2(n16356), .ZN(n13209) );
  NAND2_X1 U15268 ( .A1(n16337), .A2(n13209), .ZN(n12284) );
  NOR2_X1 U15269 ( .A1(n16338), .A2(n12284), .ZN(n12285) );
  AOI21_X1 U15270 ( .B1(n16340), .B2(n16341), .A(n12285), .ZN(n13214) );
  NAND2_X1 U15271 ( .A1(n12286), .A2(n13041), .ZN(n12287) );
  NAND2_X1 U15272 ( .A1(n13214), .A2(n12287), .ZN(n12288) );
  NAND2_X1 U15273 ( .A1(n19147), .A2(n19292), .ZN(n13669) );
  NOR4_X1 U15274 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12292) );
  NOR4_X1 U15275 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12291) );
  NOR4_X1 U15276 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12290) );
  NOR4_X1 U15277 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12289) );
  NAND4_X1 U15278 ( .A1(n12292), .A2(n12291), .A3(n12290), .A4(n12289), .ZN(
        n12297) );
  NOR4_X1 U15279 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12295) );
  NOR4_X1 U15280 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12294) );
  NOR4_X1 U15281 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12293) );
  INV_X1 U15282 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19883) );
  NAND4_X1 U15283 ( .A1(n12295), .A2(n12294), .A3(n12293), .A4(n19883), .ZN(
        n12296) );
  OAI21_X1 U15284 ( .B1(n12297), .B2(n12296), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12298) );
  INV_X2 U15285 ( .A(n14107), .ZN(n14105) );
  NOR3_X4 U15286 ( .A1(n13669), .A2(n13668), .A3(n14105), .ZN(n19120) );
  INV_X1 U15287 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12299) );
  OAI22_X1 U15288 ( .A1(n15065), .A2(n14309), .B1(n19147), .B2(n12299), .ZN(
        n12300) );
  AOI21_X1 U15289 ( .B1(n19120), .B2(BUF1_REG_30__SCAN_IN), .A(n12300), .ZN(
        n12305) );
  NOR3_X2 U15290 ( .A1(n13669), .A2(n13668), .A3(n14107), .ZN(n19121) );
  INV_X1 U15291 ( .A(n13669), .ZN(n12301) );
  NAND2_X1 U15292 ( .A1(n14105), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12303) );
  INV_X1 U15293 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16460) );
  OR2_X1 U15294 ( .A1(n14105), .A2(n16460), .ZN(n12302) );
  NAND2_X1 U15295 ( .A1(n12303), .A2(n12302), .ZN(n19228) );
  AOI22_X1 U15296 ( .A1(n19121), .A2(BUF2_REG_30__SCAN_IN), .B1(n16165), .B2(
        n19228), .ZN(n12304) );
  AND2_X1 U15297 ( .A1(n12305), .A2(n12304), .ZN(n12306) );
  OAI21_X1 U15298 ( .B1(n14322), .B2(n19174), .A(n12306), .ZN(P2_U2889) );
  NAND2_X1 U15299 ( .A1(n9829), .A2(n15594), .ZN(n14101) );
  NAND2_X1 U15300 ( .A1(n12438), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12310) );
  INV_X1 U15301 ( .A(n11938), .ZN(n12308) );
  NAND2_X1 U15302 ( .A1(n15564), .A2(n12308), .ZN(n12315) );
  NOR2_X2 U15303 ( .A1(n12332), .A2(n12315), .ZN(n12352) );
  NAND2_X1 U15304 ( .A1(n12352), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12309) );
  OAI211_X1 U15305 ( .C1(n14118), .C2(n14101), .A(n12310), .B(n12309), .ZN(
        n12311) );
  INV_X1 U15306 ( .A(n12311), .ZN(n12327) );
  AND2_X1 U15307 ( .A1(n15564), .A2(n11938), .ZN(n12330) );
  OR2_X1 U15308 ( .A1(n15569), .A2(n15564), .ZN(n12328) );
  NOR2_X2 U15309 ( .A1(n12332), .A2(n12328), .ZN(n12379) );
  AOI22_X1 U15310 ( .A1(n19785), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12326) );
  AND2_X1 U15311 ( .A1(n15569), .A2(n19110), .ZN(n12313) );
  INV_X1 U15312 ( .A(n12313), .ZN(n12314) );
  NOR2_X2 U15313 ( .A1(n12332), .A2(n12314), .ZN(n12377) );
  AOI22_X1 U15314 ( .A1(n19753), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12377), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12325) );
  INV_X1 U15315 ( .A(n12315), .ZN(n12333) );
  AND2_X1 U15316 ( .A1(n9804), .A2(n12333), .ZN(n12316) );
  OAI22_X1 U15317 ( .A1(n12318), .A2(n19301), .B1(n19427), .B2(n12317), .ZN(
        n12323) );
  INV_X1 U15318 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12321) );
  INV_X1 U15319 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12320) );
  OAI22_X1 U15320 ( .A1(n12321), .A2(n19361), .B1(n19492), .B2(n12320), .ZN(
        n12322) );
  NOR2_X1 U15321 ( .A1(n12323), .A2(n12322), .ZN(n12324) );
  NAND4_X1 U15322 ( .A1(n12327), .A2(n12326), .A3(n12325), .A4(n12324), .ZN(
        n12341) );
  INV_X1 U15323 ( .A(n12328), .ZN(n12329) );
  INV_X1 U15324 ( .A(n12330), .ZN(n12331) );
  NOR2_X2 U15325 ( .A1(n12332), .A2(n12331), .ZN(n12386) );
  NAND2_X1 U15326 ( .A1(n19330), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12338) );
  NAND2_X1 U15327 ( .A1(n19706), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12337) );
  NAND2_X1 U15328 ( .A1(n12378), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12336) );
  NAND4_X1 U15329 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12340) );
  NOR2_X1 U15330 ( .A1(n12341), .A2(n12340), .ZN(n12342) );
  NAND2_X1 U15331 ( .A1(n12342), .A2(n19264), .ZN(n12345) );
  NAND2_X1 U15332 ( .A1(n12343), .A2(n13446), .ZN(n12344) );
  INV_X1 U15333 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12346) );
  OAI22_X1 U15334 ( .A1(n12349), .A2(n19301), .B1(n19427), .B2(n12348), .ZN(
        n12350) );
  NOR2_X1 U15335 ( .A1(n12351), .A2(n12350), .ZN(n12356) );
  AOI22_X1 U15336 ( .A1(n19706), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12355) );
  AOI22_X1 U15337 ( .A1(n19753), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12377), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15338 ( .A1(n19785), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12386), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12353) );
  INV_X1 U15339 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12357) );
  OAI21_X1 U15340 ( .B1(n19492), .B2(n12357), .A(n19264), .ZN(n12358) );
  AOI21_X1 U15341 ( .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n19330), .A(
        n12358), .ZN(n12362) );
  AOI22_X1 U15342 ( .A1(n19675), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12361) );
  INV_X1 U15343 ( .A(n14101), .ZN(n14112) );
  NAND2_X1 U15344 ( .A1(n14112), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12360) );
  NAND2_X1 U15345 ( .A1(n12378), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12359) );
  AND2_X1 U15346 ( .A1(n13446), .A2(n12624), .ZN(n13264) );
  AND2_X1 U15347 ( .A1(n13264), .A2(n12622), .ZN(n12619) );
  NAND2_X1 U15348 ( .A1(n14112), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12366) );
  NAND2_X1 U15349 ( .A1(n19785), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12365) );
  OAI211_X1 U15350 ( .C1(n12368), .C2(n12367), .A(n12366), .B(n12365), .ZN(
        n12376) );
  INV_X1 U15351 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12370) );
  OAI22_X1 U15352 ( .A1(n12370), .A2(n19492), .B1(n19301), .B2(n12369), .ZN(
        n12374) );
  INV_X1 U15353 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12372) );
  OAI22_X1 U15354 ( .A1(n12372), .A2(n19361), .B1(n19427), .B2(n12371), .ZN(
        n12373) );
  OR2_X1 U15355 ( .A1(n12374), .A2(n12373), .ZN(n12375) );
  NOR2_X1 U15356 ( .A1(n12376), .A2(n12375), .ZN(n12395) );
  AOI22_X1 U15357 ( .A1(n19675), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12377), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12394) );
  NAND2_X1 U15358 ( .A1(n19330), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12381) );
  NAND2_X1 U15359 ( .A1(n12379), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12380) );
  OAI211_X1 U15360 ( .C1(n19461), .C2(n12382), .A(n12381), .B(n12380), .ZN(
        n12383) );
  INV_X1 U15361 ( .A(n12383), .ZN(n12393) );
  INV_X1 U15362 ( .A(n12352), .ZN(n19561) );
  INV_X1 U15363 ( .A(n19753), .ZN(n19746) );
  OAI22_X1 U15364 ( .A1(n12385), .A2(n19561), .B1(n19746), .B2(n12384), .ZN(
        n12391) );
  INV_X1 U15365 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12389) );
  INV_X1 U15366 ( .A(n12386), .ZN(n12388) );
  INV_X1 U15367 ( .A(n19706), .ZN(n12434) );
  OAI22_X1 U15368 ( .A1(n12389), .A2(n12388), .B1(n12434), .B2(n12387), .ZN(
        n12390) );
  NOR2_X1 U15369 ( .A1(n12391), .A2(n12390), .ZN(n12392) );
  NAND4_X1 U15370 ( .A1(n12395), .A2(n12394), .A3(n12393), .A4(n12392), .ZN(
        n12398) );
  NAND2_X1 U15371 ( .A1(n12396), .A2(n13446), .ZN(n12397) );
  NAND2_X1 U15372 ( .A1(n12639), .A2(n12399), .ZN(n12403) );
  NAND2_X1 U15373 ( .A1(n12421), .A2(n12401), .ZN(n12402) );
  NAND2_X1 U15374 ( .A1(n10130), .A2(n12402), .ZN(n19074) );
  INV_X1 U15375 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14181) );
  NAND2_X1 U15376 ( .A1(n12405), .A2(n12404), .ZN(n12406) );
  NAND2_X1 U15377 ( .A1(n12630), .A2(n12399), .ZN(n12410) );
  INV_X1 U15378 ( .A(n12422), .ZN(n12409) );
  NAND2_X1 U15379 ( .A1(n12411), .A2(n12407), .ZN(n12408) );
  NAND2_X1 U15380 ( .A1(n12409), .A2(n12408), .ZN(n13975) );
  OAI21_X1 U15381 ( .B1(n12415), .B2(n12412), .A(n12411), .ZN(n13993) );
  INV_X1 U15382 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13058) );
  MUX2_X1 U15383 ( .A(n12413), .B(n12600), .S(n13035), .Z(n12608) );
  INV_X1 U15384 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13343) );
  MUX2_X1 U15385 ( .A(n12608), .B(n13343), .S(n12592), .Z(n19104) );
  INV_X1 U15386 ( .A(n19104), .ZN(n12414) );
  NAND2_X1 U15387 ( .A1(n12414), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13278) );
  INV_X1 U15388 ( .A(n12415), .ZN(n12417) );
  INV_X1 U15389 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13338) );
  NAND3_X1 U15390 ( .A1(n12592), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12416) );
  NAND2_X1 U15391 ( .A1(n12417), .A2(n12416), .ZN(n14882) );
  NOR2_X1 U15392 ( .A1(n13278), .A2(n14882), .ZN(n12418) );
  NAND2_X1 U15393 ( .A1(n13278), .A2(n14882), .ZN(n13277) );
  OAI21_X1 U15394 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12418), .A(
        n13277), .ZN(n13303) );
  XNOR2_X1 U15395 ( .A(n13993), .B(n13058), .ZN(n13302) );
  OR2_X1 U15396 ( .A1(n13303), .A2(n13302), .ZN(n13305) );
  OAI21_X1 U15397 ( .B1(n13993), .B2(n13058), .A(n13305), .ZN(n15548) );
  OAI21_X1 U15398 ( .B1(n15550), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n15548), .ZN(n12420) );
  NAND2_X1 U15399 ( .A1(n15550), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12419) );
  NAND2_X1 U15400 ( .A1(n12420), .A2(n12419), .ZN(n14029) );
  OAI21_X1 U15401 ( .B1(n12423), .B2(n12422), .A(n12421), .ZN(n19086) );
  XNOR2_X1 U15402 ( .A(n19086), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14030) );
  NAND2_X1 U15403 ( .A1(n14029), .A2(n14030), .ZN(n12426) );
  INV_X1 U15404 ( .A(n19086), .ZN(n12424) );
  NAND2_X1 U15405 ( .A1(n12424), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12425) );
  NAND2_X1 U15406 ( .A1(n12427), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12428) );
  NAND2_X1 U15407 ( .A1(n19330), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12431) );
  NAND2_X1 U15408 ( .A1(n19753), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12430) );
  OAI211_X1 U15409 ( .C1(n19461), .C2(n12432), .A(n12431), .B(n12430), .ZN(
        n12437) );
  INV_X1 U15410 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12435) );
  INV_X1 U15411 ( .A(n19675), .ZN(n19682) );
  OAI22_X1 U15412 ( .A1(n12435), .A2(n19682), .B1(n12434), .B2(n12433), .ZN(
        n12436) );
  NOR2_X1 U15413 ( .A1(n12437), .A2(n12436), .ZN(n12452) );
  INV_X1 U15414 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19287) );
  NAND2_X1 U15415 ( .A1(n12438), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12440) );
  NAND2_X1 U15416 ( .A1(n12386), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12439) );
  OAI211_X1 U15417 ( .C1(n14101), .C2(n19287), .A(n12440), .B(n12439), .ZN(
        n12448) );
  INV_X1 U15418 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12442) );
  INV_X1 U15419 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12441) );
  OAI22_X1 U15420 ( .A1(n12442), .A2(n19361), .B1(n19492), .B2(n12441), .ZN(
        n12446) );
  OAI22_X1 U15421 ( .A1(n12444), .A2(n19427), .B1(n19301), .B2(n12443), .ZN(
        n12445) );
  OR2_X1 U15422 ( .A1(n12446), .A2(n12445), .ZN(n12447) );
  NOR2_X1 U15423 ( .A1(n12448), .A2(n12447), .ZN(n12451) );
  AOI22_X1 U15424 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12377), .B1(
        n12352), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15425 ( .A1(n19785), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12379), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12449) );
  NAND4_X1 U15426 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        n12456) );
  INV_X1 U15427 ( .A(n12453), .ZN(n12454) );
  NAND2_X1 U15428 ( .A1(n12454), .A2(n13446), .ZN(n12455) );
  INV_X1 U15429 ( .A(n12465), .ZN(n12459) );
  NAND2_X1 U15430 ( .A1(n10130), .A2(n10128), .ZN(n12458) );
  NAND2_X1 U15431 ( .A1(n12459), .A2(n12458), .ZN(n19061) );
  NAND2_X1 U15432 ( .A1(n12460), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12461) );
  INV_X1 U15433 ( .A(n12463), .ZN(n12464) );
  XNOR2_X1 U15434 ( .A(n12465), .B(n12464), .ZN(n13962) );
  AND2_X1 U15435 ( .A1(n13962), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15522) );
  INV_X1 U15436 ( .A(n12470), .ZN(n12467) );
  OAI21_X1 U15437 ( .B1(n10886), .B2(n12468), .A(n12467), .ZN(n13940) );
  OR2_X1 U15438 ( .A1(n13940), .A2(n12399), .ZN(n12482) );
  INV_X1 U15439 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12481) );
  NOR2_X1 U15440 ( .A1(n12482), .A2(n12481), .ZN(n15501) );
  NAND2_X1 U15441 ( .A1(n12592), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12471) );
  MUX2_X1 U15442 ( .A(n12471), .B(n12592), .S(n12470), .Z(n12473) );
  INV_X1 U15443 ( .A(n12480), .ZN(n12472) );
  NAND2_X1 U15444 ( .A1(n19050), .A2(n12571), .ZN(n12475) );
  INV_X1 U15445 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12474) );
  NAND2_X1 U15446 ( .A1(n12475), .A2(n12474), .ZN(n15482) );
  NOR2_X1 U15447 ( .A1(n12480), .A2(n12479), .ZN(n12476) );
  NAND2_X1 U15448 ( .A1(n12592), .A2(n12476), .ZN(n12477) );
  NAND2_X1 U15449 ( .A1(n12594), .A2(n12477), .ZN(n12478) );
  AOI21_X1 U15450 ( .B1(n12480), .B2(n12479), .A(n12478), .ZN(n19040) );
  NAND2_X1 U15451 ( .A1(n19040), .A2(n12571), .ZN(n12492) );
  INV_X1 U15452 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15474) );
  NAND2_X1 U15453 ( .A1(n12492), .A2(n15474), .ZN(n15466) );
  NAND2_X1 U15454 ( .A1(n12482), .A2(n12481), .ZN(n15499) );
  INV_X1 U15455 ( .A(n13962), .ZN(n12483) );
  INV_X1 U15456 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15527) );
  NAND2_X1 U15457 ( .A1(n12483), .A2(n15527), .ZN(n15520) );
  AND2_X1 U15458 ( .A1(n15499), .A2(n15520), .ZN(n15441) );
  NAND2_X1 U15459 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n12484), .ZN(n12485) );
  NOR2_X1 U15460 ( .A1(n19277), .A2(n12485), .ZN(n12486) );
  OR2_X1 U15461 ( .A1(n12487), .A2(n12486), .ZN(n19026) );
  OAI21_X1 U15462 ( .B1(n19026), .B2(n12399), .A(n15456), .ZN(n15446) );
  AND4_X1 U15463 ( .A1(n15482), .A2(n15466), .A3(n15441), .A4(n15446), .ZN(
        n12488) );
  INV_X1 U15464 ( .A(n19026), .ZN(n12490) );
  AND2_X1 U15465 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12489) );
  NAND2_X1 U15466 ( .A1(n12490), .A2(n12489), .ZN(n15445) );
  AND2_X1 U15467 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12491) );
  NAND2_X1 U15468 ( .A1(n19050), .A2(n12491), .ZN(n15481) );
  OR2_X1 U15469 ( .A1(n15474), .A2(n12492), .ZN(n15465) );
  NAND2_X1 U15470 ( .A1(n15481), .A2(n15465), .ZN(n15444) );
  INV_X1 U15471 ( .A(n15444), .ZN(n12493) );
  AND2_X1 U15472 ( .A1(n15445), .A2(n12493), .ZN(n15434) );
  NAND2_X1 U15473 ( .A1(n10120), .A2(n9855), .ZN(n12495) );
  NAND2_X1 U15474 ( .A1(n12514), .A2(n12495), .ZN(n14098) );
  NAND2_X1 U15475 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12496) );
  OR2_X1 U15476 ( .A1(n14098), .A2(n12496), .ZN(n15435) );
  AND2_X1 U15477 ( .A1(n15434), .A2(n15435), .ZN(n15168) );
  NAND2_X1 U15478 ( .A1(n15167), .A2(n15168), .ZN(n15226) );
  NAND2_X1 U15479 ( .A1(n12592), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12497) );
  NOR2_X1 U15480 ( .A1(n12498), .A2(n12497), .ZN(n12500) );
  OR2_X1 U15481 ( .A1(n12500), .A2(n12499), .ZN(n18937) );
  INV_X1 U15482 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15189) );
  OAI21_X1 U15483 ( .B1(n18937), .B2(n12399), .A(n15189), .ZN(n15181) );
  NAND3_X1 U15484 ( .A1(n12501), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n12592), 
        .ZN(n12502) );
  NAND3_X1 U15485 ( .A1(n12503), .A2(n12594), .A3(n12502), .ZN(n18985) );
  INV_X1 U15486 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16192) );
  OAI21_X1 U15487 ( .B1(n18985), .B2(n12399), .A(n16192), .ZN(n12505) );
  NAND2_X1 U15488 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12504) );
  INV_X1 U15489 ( .A(n12506), .ZN(n12507) );
  XNOR2_X1 U15490 ( .A(n12508), .B(n12507), .ZN(n19003) );
  AOI21_X1 U15491 ( .B1(n19003), .B2(n12571), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15402) );
  INV_X1 U15492 ( .A(n12509), .ZN(n12510) );
  XNOR2_X1 U15493 ( .A(n12511), .B(n12510), .ZN(n14870) );
  NAND2_X1 U15494 ( .A1(n14870), .A2(n12571), .ZN(n12512) );
  NAND2_X1 U15495 ( .A1(n12512), .A2(n16321), .ZN(n15400) );
  OR2_X1 U15496 ( .A1(n14098), .A2(n12399), .ZN(n12513) );
  INV_X1 U15497 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15430) );
  NAND2_X1 U15498 ( .A1(n12513), .A2(n15430), .ZN(n15436) );
  XNOR2_X1 U15499 ( .A(n12514), .B(n9877), .ZN(n19013) );
  NAND2_X1 U15500 ( .A1(n19013), .A2(n12571), .ZN(n12533) );
  INV_X1 U15501 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15415) );
  NAND2_X1 U15502 ( .A1(n12533), .A2(n15415), .ZN(n15228) );
  NAND3_X1 U15503 ( .A1(n15400), .A2(n15436), .A3(n15228), .ZN(n12515) );
  NOR2_X1 U15504 ( .A1(n15402), .A2(n12515), .ZN(n12518) );
  XNOR2_X1 U15505 ( .A(n12517), .B(n10124), .ZN(n18972) );
  NAND2_X1 U15506 ( .A1(n18972), .A2(n12571), .ZN(n12539) );
  INV_X1 U15507 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12538) );
  NAND2_X1 U15508 ( .A1(n12539), .A2(n12538), .ZN(n15175) );
  AND4_X1 U15509 ( .A1(n15181), .A2(n15394), .A3(n12518), .A4(n15175), .ZN(
        n12527) );
  NAND2_X1 U15510 ( .A1(n12592), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12519) );
  MUX2_X1 U15511 ( .A(n12592), .B(n12519), .S(n12520), .Z(n12521) );
  OR2_X1 U15512 ( .A1(n12520), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12523) );
  NAND2_X1 U15513 ( .A1(n14853), .A2(n12571), .ZN(n12522) );
  INV_X1 U15514 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16183) );
  NAND2_X1 U15515 ( .A1(n12522), .A2(n16183), .ZN(n16176) );
  NAND3_X1 U15516 ( .A1(n12523), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n12592), 
        .ZN(n12524) );
  AND2_X1 U15517 ( .A1(n12524), .A2(n12526), .ZN(n18956) );
  NAND2_X1 U15518 ( .A1(n18956), .A2(n12571), .ZN(n12531) );
  INV_X1 U15519 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16280) );
  NAND2_X1 U15520 ( .A1(n12531), .A2(n16280), .ZN(n15207) );
  NAND2_X1 U15521 ( .A1(n16176), .A2(n15207), .ZN(n15193) );
  NAND2_X1 U15522 ( .A1(n12592), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12525) );
  XNOR2_X1 U15523 ( .A(n12526), .B(n12525), .ZN(n18945) );
  AOI21_X1 U15524 ( .B1(n18945), .B2(n12571), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15196) );
  NOR2_X1 U15525 ( .A1(n15193), .A2(n15196), .ZN(n15179) );
  INV_X1 U15526 ( .A(n18937), .ZN(n12530) );
  AND2_X1 U15527 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12529) );
  NAND2_X1 U15528 ( .A1(n12530), .A2(n12529), .ZN(n15180) );
  INV_X1 U15529 ( .A(n12531), .ZN(n12532) );
  NAND2_X1 U15530 ( .A1(n12532), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15208) );
  NAND2_X1 U15531 ( .A1(n15173), .A2(n15398), .ZN(n12536) );
  AND2_X1 U15532 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12534) );
  AND2_X1 U15533 ( .A1(n19003), .A2(n12534), .ZN(n15401) );
  AND2_X1 U15534 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12535) );
  AND2_X1 U15535 ( .A1(n14870), .A2(n12535), .ZN(n16206) );
  OR2_X1 U15536 ( .A1(n15401), .A2(n16206), .ZN(n15172) );
  NOR2_X1 U15537 ( .A1(n12536), .A2(n15172), .ZN(n12540) );
  AND2_X1 U15538 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12537) );
  NAND2_X1 U15539 ( .A1(n18945), .A2(n12537), .ZN(n15178) );
  AND4_X1 U15540 ( .A1(n15208), .A2(n12540), .A3(n15178), .A4(n15176), .ZN(
        n12542) );
  AND2_X1 U15541 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12541) );
  NAND2_X1 U15542 ( .A1(n14853), .A2(n12541), .ZN(n16175) );
  AND3_X1 U15543 ( .A1(n15180), .A2(n12542), .A3(n16175), .ZN(n12543) );
  INV_X1 U15544 ( .A(n12544), .ZN(n12545) );
  NAND2_X1 U15545 ( .A1(n12546), .A2(n12545), .ZN(n12547) );
  NAND2_X1 U15546 ( .A1(n12550), .A2(n12547), .ZN(n15667) );
  NAND2_X1 U15547 ( .A1(n12548), .A2(n15348), .ZN(n15335) );
  NAND2_X1 U15548 ( .A1(n12550), .A2(n12549), .ZN(n12551) );
  NAND2_X1 U15549 ( .A1(n12555), .A2(n12551), .ZN(n16143) );
  OR2_X1 U15550 ( .A1(n16143), .A2(n12399), .ZN(n12552) );
  XNOR2_X1 U15551 ( .A(n12552), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15161) );
  NAND2_X1 U15552 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12553) );
  OR2_X1 U15553 ( .A1(n16143), .A2(n12553), .ZN(n12554) );
  NAND3_X1 U15554 ( .A1(n12555), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n12592), 
        .ZN(n12556) );
  NAND2_X1 U15555 ( .A1(n12556), .A2(n12594), .ZN(n12557) );
  OR2_X1 U15556 ( .A1(n12566), .A2(n12557), .ZN(n14852) );
  NOR2_X1 U15557 ( .A1(n14852), .A2(n12399), .ZN(n12559) );
  NAND2_X1 U15558 ( .A1(n15149), .A2(n15152), .ZN(n12562) );
  INV_X1 U15559 ( .A(n12559), .ZN(n12560) );
  NOR2_X1 U15560 ( .A1(n12566), .A2(n14930), .ZN(n12563) );
  NAND2_X1 U15561 ( .A1(n12592), .A2(n12563), .ZN(n12564) );
  NAND2_X1 U15562 ( .A1(n12594), .A2(n12564), .ZN(n12565) );
  AOI21_X1 U15563 ( .B1(n12566), .B2(n14930), .A(n12565), .ZN(n16132) );
  AOI21_X1 U15564 ( .B1(n16132), .B2(n12571), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15136) );
  NAND2_X1 U15565 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n12567), .ZN(n12568) );
  NOR2_X1 U15566 ( .A1(n19277), .A2(n12568), .ZN(n12569) );
  NOR2_X1 U15567 ( .A1(n12570), .A2(n12569), .ZN(n16121) );
  INV_X1 U15568 ( .A(n15102), .ZN(n12575) );
  NAND2_X1 U15569 ( .A1(n12580), .A2(n12572), .ZN(n12573) );
  NAND2_X1 U15570 ( .A1(n12574), .A2(n12573), .ZN(n14839) );
  AOI21_X1 U15571 ( .B1(n12575), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15104), .ZN(n12585) );
  INV_X1 U15572 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15109) );
  INV_X1 U15573 ( .A(n12576), .ZN(n12578) );
  NAND2_X1 U15574 ( .A1(n12578), .A2(n12577), .ZN(n12579) );
  NAND2_X1 U15575 ( .A1(n12580), .A2(n12579), .ZN(n16109) );
  INV_X1 U15576 ( .A(n12581), .ZN(n12583) );
  INV_X1 U15577 ( .A(n16132), .ZN(n12582) );
  INV_X1 U15578 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15303) );
  AOI21_X1 U15579 ( .B1(n12583), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15138), .ZN(n15101) );
  XNOR2_X1 U15580 ( .A(n12587), .B(n12586), .ZN(n12589) );
  INV_X1 U15581 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15251) );
  OAI21_X1 U15582 ( .B1(n12589), .B2(n12399), .A(n15251), .ZN(n15084) );
  NAND2_X1 U15583 ( .A1(n15086), .A2(n15084), .ZN(n14305) );
  AOI21_X1 U15584 ( .B1(n12588), .B2(n12571), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14306) );
  INV_X1 U15585 ( .A(n12589), .ZN(n16096) );
  NAND3_X1 U15586 ( .A1(n16096), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12571), .ZN(n15085) );
  OAI21_X2 U15587 ( .B1(n14305), .B2(n14306), .A(n12591), .ZN(n12598) );
  OAI21_X1 U15588 ( .B1(n12593), .B2(P2_EBX_REG_30__SCAN_IN), .A(n12592), .ZN(
        n12595) );
  NAND2_X1 U15589 ( .A1(n12595), .A2(n12594), .ZN(n16085) );
  NOR2_X1 U15590 ( .A1(n16085), .A2(n12399), .ZN(n12596) );
  XOR2_X1 U15591 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12596), .Z(
        n12597) );
  XNOR2_X1 U15592 ( .A(n12598), .B(n12597), .ZN(n13093) );
  OR2_X1 U15593 ( .A1(n12599), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13222) );
  INV_X1 U15594 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13220) );
  OAI21_X1 U15595 ( .B1(n10635), .B2(n13222), .A(n13220), .ZN(n19983) );
  NOR2_X1 U15596 ( .A1(n12601), .A2(n12600), .ZN(n12602) );
  NOR2_X1 U15597 ( .A1(n16338), .A2(n12602), .ZN(n12603) );
  MUX2_X1 U15598 ( .A(n19983), .B(n12603), .S(n19855), .Z(n15758) );
  NAND2_X1 U15599 ( .A1(n15758), .A2(n19264), .ZN(n12616) );
  INV_X1 U15600 ( .A(n12604), .ZN(n12610) );
  INV_X1 U15601 ( .A(n12605), .ZN(n12606) );
  OAI21_X1 U15602 ( .B1(n12608), .B2(n12607), .A(n12606), .ZN(n12609) );
  AND3_X1 U15603 ( .A1(n12611), .A2(n12610), .A3(n12609), .ZN(n12613) );
  OR2_X1 U15604 ( .A1(n12613), .A2(n12612), .ZN(n19991) );
  INV_X1 U15605 ( .A(n19991), .ZN(n12614) );
  NAND2_X1 U15606 ( .A1(n12614), .A2(n16362), .ZN(n12615) );
  NAND2_X1 U15607 ( .A1(n12616), .A2(n12615), .ZN(n13019) );
  NOR2_X1 U15608 ( .A1(n13088), .A2(n13230), .ZN(n12617) );
  INV_X1 U15609 ( .A(n12670), .ZN(n12618) );
  XOR2_X1 U15610 ( .A(n12620), .B(n12619), .Z(n13308) );
  INV_X1 U15611 ( .A(n13264), .ZN(n12621) );
  NAND2_X1 U15612 ( .A1(n12621), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13266) );
  INV_X1 U15613 ( .A(n12622), .ZN(n12623) );
  XOR2_X1 U15614 ( .A(n12624), .B(n12623), .Z(n12625) );
  NOR2_X1 U15615 ( .A1(n13266), .A2(n12625), .ZN(n12626) );
  XNOR2_X1 U15616 ( .A(n13266), .B(n12625), .ZN(n13273) );
  NOR2_X1 U15617 ( .A1(n15580), .A2(n13273), .ZN(n13272) );
  NOR2_X1 U15618 ( .A1(n12626), .A2(n13272), .ZN(n12627) );
  XOR2_X1 U15619 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12627), .Z(
        n13307) );
  NOR2_X1 U15620 ( .A1(n13308), .A2(n13307), .ZN(n13306) );
  NOR2_X1 U15621 ( .A1(n12627), .A2(n13058), .ZN(n12628) );
  OR2_X1 U15622 ( .A1(n13306), .A2(n12628), .ZN(n12631) );
  INV_X1 U15623 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12629) );
  XNOR2_X1 U15624 ( .A(n12631), .B(n12629), .ZN(n15552) );
  NAND2_X1 U15625 ( .A1(n12631), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12632) );
  NAND2_X1 U15626 ( .A1(n14037), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12637) );
  NAND2_X1 U15627 ( .A1(n12635), .A2(n10211), .ZN(n12636) );
  NAND2_X1 U15628 ( .A1(n12633), .A2(n12636), .ZN(n14038) );
  INV_X1 U15629 ( .A(n14037), .ZN(n12638) );
  NAND2_X1 U15630 ( .A1(n12639), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14172) );
  INV_X1 U15631 ( .A(n14172), .ZN(n14175) );
  NAND2_X1 U15632 ( .A1(n14175), .A2(n12644), .ZN(n12642) );
  NAND2_X1 U15633 ( .A1(n12640), .A2(n12648), .ZN(n12641) );
  NAND2_X1 U15634 ( .A1(n15240), .A2(n12647), .ZN(n12655) );
  NAND2_X1 U15635 ( .A1(n12649), .A2(n10188), .ZN(n15515) );
  INV_X1 U15636 ( .A(n15517), .ZN(n12650) );
  NAND2_X1 U15637 ( .A1(n12650), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12651) );
  NAND2_X1 U15638 ( .A1(n15515), .A2(n12651), .ZN(n12653) );
  NAND2_X1 U15639 ( .A1(n12653), .A2(n12652), .ZN(n12654) );
  NAND2_X1 U15640 ( .A1(n12571), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12658) );
  NAND3_X1 U15641 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16306) );
  NOR2_X1 U15642 ( .A1(n15474), .A2(n15456), .ZN(n15455) );
  NAND2_X1 U15643 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15455), .ZN(
        n15414) );
  NOR2_X1 U15644 ( .A1(n16306), .A2(n15414), .ZN(n15375) );
  AND2_X1 U15645 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12660) );
  AND2_X1 U15646 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n12660), .ZN(
        n16299) );
  INV_X1 U15647 ( .A(n16299), .ZN(n13062) );
  NAND2_X1 U15648 ( .A1(n15213), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15201) );
  INV_X1 U15649 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12661) );
  NOR2_X2 U15650 ( .A1(n15201), .A2(n12661), .ZN(n15186) );
  NAND2_X2 U15651 ( .A1(n12662), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15129) );
  INV_X1 U15652 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15286) );
  AOI22_X1 U15653 ( .A1(n12663), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12665) );
  NAND2_X1 U15654 ( .A1(n10482), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12664) );
  OAI211_X1 U15655 ( .C1(n10498), .C2(n12666), .A(n12665), .B(n12664), .ZN(
        n12668) );
  NOR2_X1 U15656 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16369) );
  NOR2_X1 U15657 ( .A1(n19851), .A2(n19855), .ZN(n19984) );
  INV_X1 U15658 ( .A(n14106), .ZN(n19255) );
  NOR2_X1 U15659 ( .A1(n16092), .A2(n14106), .ZN(n12677) );
  NAND2_X1 U15660 ( .A1(n12670), .A2(n19259), .ZN(n13212) );
  INV_X1 U15661 ( .A(n15611), .ZN(n19947) );
  OR2_X1 U15662 ( .A1(n19945), .A2(n19947), .ZN(n19969) );
  NAND2_X1 U15663 ( .A1(n19969), .A2(n18906), .ZN(n12671) );
  NAND2_X1 U15664 ( .A1(n19457), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12672) );
  NAND2_X1 U15665 ( .A1(n12673), .A2(n12672), .ZN(n13269) );
  NAND2_X1 U15666 ( .A1(n19076), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n13080) );
  NAND2_X1 U15667 ( .A1(n19245), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12674) );
  OAI211_X1 U15668 ( .C1(n19253), .C2(n12675), .A(n13080), .B(n12674), .ZN(
        n12676) );
  NOR2_X1 U15669 ( .A1(n12677), .A2(n12676), .ZN(n12678) );
  OAI211_X1 U15670 ( .C1(n13093), .C2(n19237), .A(n12679), .B(n12678), .ZN(
        P2_U2983) );
  INV_X4 U15671 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12687) );
  INV_X2 U15672 ( .A(n12680), .ZN(n12737) );
  INV_X2 U15673 ( .A(n12737), .ZN(n17153) );
  INV_X1 U15674 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17128) );
  NOR2_X2 U15675 ( .A1(n16933), .A2(n12687), .ZN(n18689) );
  NAND3_X1 U15676 ( .A1(n18849), .A2(n18839), .A3(n18689), .ZN(n17199) );
  AOI22_X1 U15678 ( .A1(n17222), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12681) );
  OAI21_X1 U15679 ( .B1(n10239), .B2(n17128), .A(n12681), .ZN(n12696) );
  INV_X1 U15680 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16959) );
  INV_X2 U15681 ( .A(n12709), .ZN(n12780) );
  AOI22_X1 U15682 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12694) );
  NOR3_X2 U15684 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n16933), .ZN(n12684) );
  NAND2_X4 U15685 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12684), .ZN(
        n17216) );
  INV_X1 U15686 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17124) );
  OAI22_X1 U15687 ( .A1(n17218), .A2(n17247), .B1(n17216), .B2(n17124), .ZN(
        n12692) );
  INV_X2 U15688 ( .A(n9849), .ZN(n15618) );
  AOI22_X1 U15689 ( .A1(n9800), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12690) );
  NOR2_X2 U15690 ( .A1(n18670), .A2(n12686), .ZN(n17221) );
  AOI22_X1 U15691 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12689) );
  INV_X2 U15692 ( .A(n12715), .ZN(n17043) );
  AOI22_X1 U15693 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12688) );
  NAND3_X1 U15694 ( .A1(n12690), .A2(n12689), .A3(n12688), .ZN(n12691) );
  AOI211_X1 U15695 ( .C1(n17235), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n12692), .B(n12691), .ZN(n12693) );
  OAI211_X1 U15696 ( .C1(n17193), .C2(n16959), .A(n12694), .B(n12693), .ZN(
        n12695) );
  INV_X1 U15697 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13806) );
  INV_X2 U15698 ( .A(n12697), .ZN(n17063) );
  AOI22_X1 U15699 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12698) );
  OAI21_X1 U15700 ( .B1(n13841), .B2(n13806), .A(n12698), .ZN(n12708) );
  INV_X1 U15701 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U15702 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12706) );
  INV_X2 U15703 ( .A(n10257), .ZN(n17220) );
  AOI22_X1 U15704 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12699) );
  OAI21_X1 U15705 ( .B1(n17218), .B2(n17253), .A(n12699), .ZN(n12704) );
  INV_X1 U15706 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15707 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12701) );
  INV_X2 U15708 ( .A(n12780), .ZN(n17090) );
  AOI22_X1 U15709 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12700) );
  OAI211_X1 U15710 ( .C1(n17216), .C2(n12702), .A(n12701), .B(n12700), .ZN(
        n12703) );
  AOI211_X1 U15711 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n12704), .B(n12703), .ZN(n12705) );
  OAI211_X1 U15712 ( .C1(n10239), .C2(n17026), .A(n12706), .B(n12705), .ZN(
        n12707) );
  INV_X1 U15713 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U15714 ( .A1(n12723), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12710) );
  OAI21_X1 U15715 ( .B1(n12780), .B2(n17061), .A(n12710), .ZN(n12714) );
  AOI22_X1 U15716 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12712) );
  INV_X1 U15717 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17157) );
  NAND3_X1 U15718 ( .A1(n12712), .A2(n12711), .A3(n10244), .ZN(n12713) );
  INV_X1 U15719 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U15720 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12716) );
  OAI21_X1 U15721 ( .B1(n17216), .B2(n12906), .A(n12716), .ZN(n12720) );
  INV_X1 U15722 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U15723 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15724 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12717) );
  OAI211_X1 U15725 ( .C1(n17218), .C2(n17263), .A(n12718), .B(n12717), .ZN(
        n12719) );
  AOI211_X1 U15726 ( .C1(n17043), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n12720), .B(n12719), .ZN(n12721) );
  AOI22_X1 U15727 ( .A1(n12680), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15728 ( .A1(n12723), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12724) );
  OAI211_X1 U15729 ( .C1(n17218), .C2(n17270), .A(n12725), .B(n12724), .ZN(
        n12726) );
  INV_X1 U15730 ( .A(n12726), .ZN(n12736) );
  AOI22_X1 U15731 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12709), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15732 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15733 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12728) );
  NAND2_X1 U15734 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12727) );
  AOI22_X1 U15735 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12734) );
  INV_X1 U15736 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12731) );
  NAND4_X2 U15737 ( .A1(n12736), .A2(n12735), .A3(n12734), .A4(n12733), .ZN(
        n12964) );
  AOI22_X1 U15738 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15739 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15740 ( .A1(n12723), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12739) );
  NAND2_X1 U15741 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12738) );
  NAND4_X1 U15742 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12750) );
  INV_X1 U15743 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U15744 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U15745 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12709), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12742) );
  OAI211_X1 U15746 ( .C1(n17191), .C2(n17174), .A(n12743), .B(n12742), .ZN(
        n12744) );
  INV_X1 U15747 ( .A(n12744), .ZN(n12748) );
  AOI22_X1 U15748 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12747) );
  INV_X1 U15749 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17267) );
  NAND2_X1 U15750 ( .A1(n12748), .A2(n9859), .ZN(n12749) );
  NAND2_X1 U15751 ( .A1(n12964), .A2(n17423), .ZN(n12772) );
  AOI22_X1 U15752 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12760) );
  INV_X1 U15753 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U15754 ( .A1(n12723), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U15755 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12751) );
  OAI211_X1 U15756 ( .C1(n17191), .C2(n17140), .A(n12752), .B(n12751), .ZN(
        n12758) );
  AOI22_X1 U15757 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15758 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15759 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12754) );
  NAND2_X1 U15760 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12753) );
  NAND4_X1 U15761 ( .A1(n12756), .A2(n12755), .A3(n12754), .A4(n12753), .ZN(
        n12757) );
  AOI211_X1 U15762 ( .C1(n17175), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n12758), .B(n12757), .ZN(n12759) );
  OAI211_X1 U15763 ( .C1(n17218), .C2(n17261), .A(n12760), .B(n12759), .ZN(
        n12795) );
  NAND2_X1 U15764 ( .A1(n12796), .A2(n12795), .ZN(n12799) );
  AOI22_X1 U15765 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12771) );
  INV_X1 U15766 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U15767 ( .A1(n17222), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U15768 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12761) );
  OAI211_X1 U15769 ( .C1(n17216), .C2(n12763), .A(n12762), .B(n12761), .ZN(
        n12769) );
  AOI22_X1 U15770 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U15771 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U15772 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12765) );
  NAND2_X1 U15773 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12764) );
  NAND4_X1 U15774 ( .A1(n12767), .A2(n12766), .A3(n12765), .A4(n12764), .ZN(
        n12768) );
  AOI211_X1 U15775 ( .C1(n17043), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n12769), .B(n12768), .ZN(n12770) );
  OAI211_X1 U15776 ( .C1(n17218), .C2(n17251), .A(n12771), .B(n12770), .ZN(
        n12953) );
  NAND2_X1 U15777 ( .A1(n12804), .A2(n12953), .ZN(n16424) );
  INV_X1 U15778 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17941) );
  INV_X1 U15779 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18033) );
  XOR2_X1 U15780 ( .A(n12772), .B(n17418), .Z(n12793) );
  INV_X1 U15781 ( .A(n12793), .ZN(n12791) );
  NAND2_X1 U15782 ( .A1(n17434), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12788) );
  INV_X1 U15783 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15784 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12773) );
  OAI21_X1 U15785 ( .B1(n17216), .B2(n12774), .A(n12773), .ZN(n12779) );
  INV_X1 U15786 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U15787 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U15788 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12776) );
  OAI211_X1 U15789 ( .C1(n17218), .C2(n17226), .A(n12777), .B(n12776), .ZN(
        n12778) );
  AOI211_X1 U15790 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n12779), .B(n12778), .ZN(n12787) );
  AOI22_X1 U15791 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12786) );
  INV_X1 U15792 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U15793 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12781) );
  OAI21_X1 U15794 ( .B1(n12697), .B2(n17217), .A(n12781), .ZN(n12784) );
  INV_X1 U15795 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17215) );
  INV_X1 U15796 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18859) );
  INV_X1 U15797 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18843) );
  INV_X1 U15798 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18193) );
  OR2_X1 U15799 ( .A1(n18193), .A2(n12789), .ZN(n12790) );
  XNOR2_X1 U15800 ( .A(n12791), .B(n12792), .ZN(n17876) );
  NAND2_X1 U15801 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  INV_X1 U15802 ( .A(n12795), .ZN(n17415) );
  XNOR2_X1 U15803 ( .A(n12796), .B(n17415), .ZN(n12797) );
  XOR2_X1 U15804 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12797), .Z(
        n17863) );
  NAND2_X1 U15805 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12797), .ZN(
        n12798) );
  XOR2_X1 U15806 ( .A(n12799), .B(n17411), .Z(n12802) );
  XNOR2_X1 U15807 ( .A(n12801), .B(n12800), .ZN(n17852) );
  NAND2_X1 U15808 ( .A1(n17852), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17851) );
  NAND2_X1 U15809 ( .A1(n12802), .A2(n12801), .ZN(n12803) );
  NAND2_X1 U15810 ( .A1(n17851), .A2(n12803), .ZN(n17833) );
  INV_X1 U15811 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18158) );
  XNOR2_X1 U15812 ( .A(n18158), .B(n12953), .ZN(n17839) );
  XOR2_X1 U15813 ( .A(n12804), .B(n17839), .Z(n17834) );
  NAND2_X1 U15814 ( .A1(n17833), .A2(n17834), .ZN(n17832) );
  NAND2_X2 U15815 ( .A1(n17832), .A2(n12805), .ZN(n17691) );
  OAI21_X1 U15816 ( .B1(n16386), .B2(n16427), .A(n17777), .ZN(n12807) );
  XNOR2_X1 U15817 ( .A(n17691), .B(n12807), .ZN(n17820) );
  NAND2_X1 U15818 ( .A1(n17820), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17821) );
  INV_X1 U15819 ( .A(n17691), .ZN(n12806) );
  NAND2_X1 U15820 ( .A1(n17821), .A2(n12808), .ZN(n12809) );
  NAND2_X2 U15821 ( .A1(n12809), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18089) );
  INV_X1 U15822 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18037) );
  NAND2_X1 U15823 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17766) );
  INV_X1 U15824 ( .A(n17766), .ZN(n18094) );
  NAND2_X1 U15825 ( .A1(n18094), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18096) );
  INV_X1 U15826 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18080) );
  NOR2_X1 U15827 ( .A1(n18096), .A2(n18080), .ZN(n18052) );
  NAND2_X1 U15828 ( .A1(n18052), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18055) );
  INV_X1 U15829 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18054) );
  NOR2_X1 U15830 ( .A1(n18055), .A2(n18054), .ZN(n18028) );
  INV_X1 U15831 ( .A(n18028), .ZN(n12810) );
  NOR2_X1 U15832 ( .A1(n18037), .A2(n12810), .ZN(n17966) );
  INV_X1 U15833 ( .A(n17966), .ZN(n17934) );
  INV_X1 U15834 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18125) );
  INV_X1 U15835 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18104) );
  NAND2_X1 U15836 ( .A1(n18125), .A2(n18104), .ZN(n17785) );
  NOR4_X1 U15837 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n17785), .ZN(n12811) );
  NOR2_X1 U15838 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17743) );
  NAND3_X1 U15839 ( .A1(n17706), .A2(n12811), .A3(n17743), .ZN(n12812) );
  NAND2_X1 U15840 ( .A1(n12812), .A2(n17777), .ZN(n12813) );
  OAI221_X1 U15841 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17777), 
        .C1(n18033), .C2(n12814), .A(n12813), .ZN(n17683) );
  INV_X1 U15842 ( .A(n12813), .ZN(n12815) );
  INV_X1 U15843 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18017) );
  NOR2_X1 U15844 ( .A1(n18033), .A2(n18017), .ZN(n18009) );
  INV_X1 U15845 ( .A(n18009), .ZN(n13002) );
  NOR2_X1 U15846 ( .A1(n17692), .A2(n13002), .ZN(n17636) );
  INV_X1 U15847 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17674) );
  NAND2_X1 U15848 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17638) );
  INV_X1 U15849 ( .A(n17638), .ZN(n17986) );
  NAND2_X1 U15850 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17986), .ZN(
        n17975) );
  INV_X1 U15851 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17974) );
  NOR2_X1 U15852 ( .A1(n17975), .A2(n17974), .ZN(n16397) );
  INV_X1 U15853 ( .A(n16397), .ZN(n17605) );
  NOR2_X1 U15854 ( .A1(n17674), .A2(n17605), .ZN(n13003) );
  NAND2_X1 U15855 ( .A1(n18009), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17968) );
  INV_X1 U15856 ( .A(n17968), .ZN(n17982) );
  NAND3_X1 U15857 ( .A1(n17982), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n17986), .ZN(n17972) );
  INV_X1 U15858 ( .A(n17972), .ZN(n17619) );
  NAND2_X1 U15859 ( .A1(n17619), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17959) );
  INV_X1 U15860 ( .A(n17959), .ZN(n13004) );
  NAND2_X1 U15861 ( .A1(n13004), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17590) );
  NAND2_X1 U15862 ( .A1(n17777), .A2(n17674), .ZN(n17673) );
  NOR2_X1 U15863 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17673), .ZN(
        n12816) );
  INV_X1 U15864 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17644) );
  NAND2_X1 U15865 ( .A1(n12816), .A2(n17644), .ZN(n17637) );
  NOR2_X1 U15866 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17637), .ZN(
        n17615) );
  INV_X1 U15867 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17952) );
  NAND3_X1 U15868 ( .A1(n17615), .A2(n17974), .A3(n17952), .ZN(n12817) );
  INV_X1 U15869 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17598) );
  INV_X1 U15870 ( .A(n12819), .ZN(n17585) );
  NAND2_X1 U15871 ( .A1(n17777), .A2(n17597), .ZN(n17584) );
  OAI221_X1 U15872 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17777), 
        .C1(n17941), .C2(n17585), .A(n17584), .ZN(n17566) );
  NAND2_X1 U15873 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17916) );
  OR2_X1 U15874 ( .A1(n12819), .A2(n17916), .ZN(n12820) );
  NOR2_X2 U15875 ( .A1(n12823), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17559) );
  INV_X1 U15876 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17540) );
  AND2_X1 U15877 ( .A1(n17777), .A2(n17540), .ZN(n12822) );
  NAND2_X1 U15878 ( .A1(n17559), .A2(n12822), .ZN(n15651) );
  NOR2_X1 U15879 ( .A1(n17777), .A2(n17540), .ZN(n12824) );
  INV_X1 U15880 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16406) );
  OAI22_X1 U15881 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n12828), .B1(
        n15745), .B2(n17777), .ZN(n12830) );
  NOR2_X1 U15882 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17814), .ZN(
        n12825) );
  AOI21_X1 U15883 ( .B1(n17814), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12825), .ZN(n12829) );
  INV_X1 U15884 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18844) );
  NAND2_X1 U15885 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17814), .ZN(
        n12826) );
  INV_X1 U15886 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15748) );
  OAI22_X1 U15887 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17814), .B1(
        n12826), .B2(n15748), .ZN(n12827) );
  AOI22_X1 U15888 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12840) );
  INV_X1 U15889 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U15890 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U15891 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12831) );
  OAI211_X1 U15892 ( .C1(n17191), .C2(n17011), .A(n12832), .B(n12831), .ZN(
        n12838) );
  AOI22_X1 U15893 ( .A1(n17222), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U15894 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U15895 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12834) );
  NAND2_X1 U15896 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12833) );
  NAND4_X1 U15897 ( .A1(n12836), .A2(n12835), .A3(n12834), .A4(n12833), .ZN(
        n12837) );
  AOI22_X1 U15898 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12850) );
  INV_X1 U15899 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13871) );
  AOI22_X1 U15900 ( .A1(n9799), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U15901 ( .A1(n17222), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12841) );
  OAI211_X1 U15902 ( .C1(n17216), .C2(n13871), .A(n12842), .B(n12841), .ZN(
        n12848) );
  AOI22_X1 U15903 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U15904 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U15905 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12844) );
  NAND2_X1 U15906 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12843) );
  NAND4_X1 U15907 ( .A1(n12846), .A2(n12845), .A3(n12844), .A4(n12843), .ZN(
        n12847) );
  AOI22_X1 U15908 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12851) );
  OAI21_X1 U15909 ( .B1(n17199), .B2(n17190), .A(n12851), .ZN(n12860) );
  AOI22_X1 U15910 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12858) );
  INV_X1 U15911 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17192) );
  INV_X1 U15912 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17092) );
  OAI22_X1 U15913 ( .A1(n17218), .A2(n17192), .B1(n17216), .B2(n17092), .ZN(
        n12856) );
  AOI22_X1 U15914 ( .A1(n9799), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U15915 ( .A1(n17222), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U15916 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12852) );
  NAND3_X1 U15917 ( .A1(n12854), .A2(n12853), .A3(n12852), .ZN(n12855) );
  AOI211_X1 U15918 ( .C1(n17235), .C2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n12856), .B(n12855), .ZN(n12857) );
  OAI211_X1 U15919 ( .C1(n12697), .C2(n17270), .A(n12858), .B(n12857), .ZN(
        n12859) );
  NAND2_X1 U15920 ( .A1(n12979), .A2(n18244), .ZN(n12942) );
  NOR2_X1 U15921 ( .A1(n12989), .A2(n12942), .ZN(n12949) );
  INV_X1 U15922 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U15923 ( .A1(n17222), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12868) );
  INV_X1 U15924 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U15925 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12861) );
  OAI21_X1 U15926 ( .B1(n17216), .B2(n12862), .A(n12861), .ZN(n12866) );
  INV_X1 U15927 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U15928 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U15929 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12863) );
  OAI211_X1 U15930 ( .C1(n17218), .C2(n17141), .A(n12864), .B(n12863), .ZN(
        n12865) );
  AOI211_X1 U15931 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n12866), .B(n12865), .ZN(n12867) );
  OAI211_X1 U15932 ( .C1(n17193), .C2(n17149), .A(n12868), .B(n12867), .ZN(
        n12873) );
  AOI22_X1 U15933 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12869) );
  OAI21_X1 U15934 ( .B1(n12697), .B2(n17261), .A(n12869), .ZN(n12871) );
  AND2_X1 U15935 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12870) );
  AOI22_X1 U15936 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12874) );
  OAI21_X1 U15937 ( .B1(n12697), .B2(n17253), .A(n12874), .ZN(n12883) );
  AOI22_X1 U15938 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12881) );
  AOI22_X1 U15939 ( .A1(n17222), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U15940 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12879) );
  INV_X1 U15941 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U15942 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12875) );
  OAI21_X1 U15943 ( .B1(n12737), .B2(n17031), .A(n12875), .ZN(n12877) );
  INV_X1 U15944 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13811) );
  INV_X1 U15945 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13807) );
  OAI22_X1 U15946 ( .A1(n17193), .A2(n13811), .B1(n17216), .B2(n13807), .ZN(
        n12876) );
  AOI211_X1 U15947 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n12877), .B(n12876), .ZN(n12878) );
  NAND4_X1 U15948 ( .A1(n12881), .A2(n12880), .A3(n12879), .A4(n12878), .ZN(
        n12882) );
  NAND2_X1 U15949 ( .A1(n18262), .A2(n12989), .ZN(n18678) );
  INV_X1 U15950 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17133) );
  AOI22_X1 U15951 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9800), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17194), .ZN(n12884) );
  OAI21_X1 U15952 ( .B1(n12737), .B2(n17133), .A(n12884), .ZN(n12885) );
  INV_X1 U15953 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16958) );
  INV_X1 U15954 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12886) );
  OAI22_X1 U15955 ( .A1(n16958), .A2(n17216), .B1(n10240), .B2(n12886), .ZN(
        n12891) );
  AOI22_X1 U15956 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17200), .ZN(n12889) );
  AOI22_X1 U15957 ( .A1(n17222), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17219), .ZN(n12888) );
  AOI22_X1 U15958 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17229), .B1(
        n17206), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12887) );
  NAND3_X1 U15959 ( .A1(n12889), .A2(n12888), .A3(n12887), .ZN(n12890) );
  AOI211_X1 U15960 ( .C1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .C2(n17043), .A(
        n12891), .B(n12890), .ZN(n12894) );
  NAND2_X1 U15961 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12893) );
  AOI22_X1 U15962 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17220), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12892) );
  AOI22_X1 U15963 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U15964 ( .A1(n12723), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12897) );
  AOI22_X1 U15965 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12896) );
  OAI211_X1 U15966 ( .C1(n17227), .C2(n17157), .A(n12897), .B(n12896), .ZN(
        n12903) );
  AOI22_X1 U15967 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U15968 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U15969 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12899) );
  NAND2_X1 U15970 ( .A1(n17229), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12898) );
  NAND4_X1 U15971 ( .A1(n12901), .A2(n12900), .A3(n12899), .A4(n12898), .ZN(
        n12902) );
  AOI211_X1 U15972 ( .C1(n17206), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n12903), .B(n12902), .ZN(n12904) );
  INV_X1 U15973 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U15974 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12907) );
  OAI21_X1 U15975 ( .B1(n12737), .B2(n17113), .A(n12907), .ZN(n12913) );
  INV_X1 U15976 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U15977 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12912) );
  AOI22_X1 U15978 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U15979 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U15980 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U15981 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12909) );
  INV_X1 U15982 ( .A(n12929), .ZN(n12914) );
  NAND2_X1 U15983 ( .A1(n17286), .A2(n18267), .ZN(n13802) );
  NAND2_X1 U15984 ( .A1(n12914), .A2(n13802), .ZN(n12915) );
  AOI21_X1 U15985 ( .B1(n12979), .B2(n12932), .A(n18257), .ZN(n12945) );
  AOI22_X1 U15986 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18684), .B2(n12687), .ZN(
        n12937) );
  INV_X1 U15987 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18235) );
  AOI22_X1 U15988 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18235), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18849), .ZN(n12923) );
  NAND2_X1 U15989 ( .A1(n18683), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12938) );
  NAND2_X1 U15990 ( .A1(n12923), .A2(n12924), .ZN(n12917) );
  OAI21_X1 U15991 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18849), .A(
        n12917), .ZN(n12918) );
  OAI22_X1 U15992 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18234), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12918), .ZN(n12920) );
  NOR2_X1 U15993 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18234), .ZN(
        n12919) );
  NAND2_X1 U15994 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12918), .ZN(
        n12921) );
  AOI22_X1 U15995 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12920), .B1(
        n12919), .B2(n12921), .ZN(n12925) );
  OAI211_X1 U15996 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18683), .A(
        n12925), .B(n12938), .ZN(n12947) );
  AOI21_X1 U15997 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12921), .A(
        n12920), .ZN(n12922) );
  AOI21_X1 U15998 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18234), .A(
        n12922), .ZN(n12939) );
  XOR2_X1 U15999 ( .A(n12924), .B(n12923), .Z(n12946) );
  NAND2_X1 U16000 ( .A1(n12925), .A2(n12946), .ZN(n12940) );
  OAI211_X1 U16001 ( .C1(n12937), .C2(n12947), .A(n12939), .B(n12940), .ZN(
        n18666) );
  NOR4_X2 U16002 ( .A1(n18252), .A2(n18257), .A3(n12927), .A4(n12928), .ZN(
        n12999) );
  INV_X1 U16003 ( .A(n12926), .ZN(n12936) );
  INV_X1 U16004 ( .A(n12927), .ZN(n12935) );
  NAND2_X1 U16005 ( .A1(n18272), .A2(n12928), .ZN(n12930) );
  AOI22_X1 U16006 ( .A1(n12930), .A2(n18257), .B1(n12929), .B2(n12928), .ZN(
        n12934) );
  OAI21_X1 U16007 ( .B1(n18247), .B2(n18238), .A(n18678), .ZN(n12931) );
  OAI21_X1 U16008 ( .B1(n12978), .B2(n12932), .A(n12931), .ZN(n12933) );
  OAI211_X1 U16009 ( .C1(n12935), .C2(n18252), .A(n12934), .B(n12933), .ZN(
        n12986) );
  NAND2_X1 U16010 ( .A1(n18238), .A2(n18885), .ZN(n12994) );
  AOI21_X1 U16011 ( .B1(n18272), .B2(n18678), .A(n12994), .ZN(n12983) );
  AOI211_X1 U16012 ( .C1(n12980), .C2(n12936), .A(n12986), .B(n12983), .ZN(
        n15644) );
  XNOR2_X1 U16013 ( .A(n12938), .B(n12937), .ZN(n12941) );
  AND2_X1 U16014 ( .A1(n18821), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18756) );
  NOR2_X1 U16015 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18740) );
  NOR3_X1 U16016 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18756), .A3(n18740), 
        .ZN(n15638) );
  AOI21_X1 U16017 ( .B1(n18885), .B2(n18247), .A(n15638), .ZN(n12943) );
  NAND2_X1 U16018 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18886) );
  INV_X1 U16019 ( .A(n18886), .ZN(n18880) );
  AOI21_X1 U16020 ( .B1(n12943), .B2(n12942), .A(n18880), .ZN(n16530) );
  NAND2_X1 U16021 ( .A1(n18262), .A2(n12979), .ZN(n12997) );
  NAND3_X1 U16022 ( .A1(n18661), .A2(n16530), .A3(n12997), .ZN(n12944) );
  OAI211_X1 U16023 ( .C1(n12945), .C2(n18666), .A(n15644), .B(n12944), .ZN(
        n12950) );
  INV_X1 U16024 ( .A(n12946), .ZN(n12948) );
  OAI21_X1 U16025 ( .B1(n12948), .B2(n12947), .A(n18661), .ZN(n16376) );
  INV_X1 U16026 ( .A(n16376), .ZN(n18663) );
  NOR2_X1 U16027 ( .A1(n18829), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18729) );
  NAND2_X1 U16028 ( .A1(n18729), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18715) );
  NAND2_X1 U16029 ( .A1(n16388), .A2(n18139), .ZN(n13018) );
  NAND2_X1 U16030 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16418) );
  INV_X1 U16031 ( .A(n16418), .ZN(n15657) );
  NAND2_X1 U16032 ( .A1(n15657), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15747) );
  NAND2_X1 U16033 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17924) );
  OR2_X1 U16034 ( .A1(n17959), .A2(n17924), .ZN(n17933) );
  NOR2_X1 U16035 ( .A1(n17933), .A2(n17916), .ZN(n16435) );
  INV_X1 U16036 ( .A(n16435), .ZN(n17909) );
  INV_X1 U16037 ( .A(n17418), .ZN(n12951) );
  INV_X1 U16038 ( .A(n10256), .ZN(n15764) );
  NAND2_X1 U16039 ( .A1(n12964), .A2(n15764), .ZN(n12960) );
  NAND2_X1 U16040 ( .A1(n12961), .A2(n12960), .ZN(n12958) );
  NAND2_X1 U16041 ( .A1(n12951), .A2(n12958), .ZN(n12956) );
  NAND2_X1 U16042 ( .A1(n12953), .A2(n17837), .ZN(n12952) );
  NOR2_X1 U16043 ( .A1(n12952), .A2(n17404), .ZN(n12975) );
  INV_X1 U16044 ( .A(n12975), .ZN(n12971) );
  XNOR2_X1 U16045 ( .A(n17404), .B(n12952), .ZN(n17823) );
  INV_X1 U16046 ( .A(n12953), .ZN(n17408) );
  INV_X1 U16047 ( .A(n17837), .ZN(n17835) );
  XOR2_X1 U16048 ( .A(n17408), .B(n17835), .Z(n12970) );
  XOR2_X1 U16049 ( .A(n17411), .B(n12954), .Z(n12955) );
  NAND2_X1 U16050 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12955), .ZN(
        n12969) );
  XOR2_X1 U16051 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n12955), .Z(
        n17847) );
  XOR2_X1 U16052 ( .A(n17415), .B(n12956), .Z(n12957) );
  NAND2_X1 U16053 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12957), .ZN(
        n12968) );
  XOR2_X1 U16054 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12957), .Z(
        n17860) );
  XNOR2_X1 U16055 ( .A(n17418), .B(n12958), .ZN(n12959) );
  NAND2_X1 U16056 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12959), .ZN(
        n12967) );
  XOR2_X1 U16057 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n12959), .Z(
        n17874) );
  XOR2_X1 U16058 ( .A(n12961), .B(n12960), .Z(n12965) );
  OR2_X1 U16059 ( .A1(n18193), .A2(n12965), .ZN(n12966) );
  AOI21_X1 U16060 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12964), .A(
        n15764), .ZN(n12963) );
  NOR2_X1 U16061 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12964), .ZN(
        n12962) );
  AOI221_X1 U16062 ( .B1(n15764), .B2(n12964), .C1(n12963), .C2(n18859), .A(
        n12962), .ZN(n17884) );
  XOR2_X1 U16063 ( .A(n18193), .B(n12965), .Z(n17883) );
  NAND2_X1 U16064 ( .A1(n17884), .A2(n17883), .ZN(n17882) );
  NAND2_X1 U16065 ( .A1(n12966), .A2(n17882), .ZN(n17873) );
  NAND2_X1 U16066 ( .A1(n17874), .A2(n17873), .ZN(n17872) );
  NAND2_X1 U16067 ( .A1(n12967), .A2(n17872), .ZN(n17859) );
  NAND2_X1 U16068 ( .A1(n17860), .A2(n17859), .ZN(n17858) );
  NAND2_X1 U16069 ( .A1(n12968), .A2(n17858), .ZN(n17846) );
  NAND2_X1 U16070 ( .A1(n17847), .A2(n17846), .ZN(n17845) );
  NAND2_X1 U16071 ( .A1(n12969), .A2(n17845), .ZN(n17836) );
  AOI222_X1 U16072 ( .A1(n12970), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n12970), .B2(n17836), .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(
        n17836), .ZN(n17824) );
  NAND2_X1 U16073 ( .A1(n17823), .A2(n17824), .ZN(n17822) );
  NAND2_X1 U16074 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17822), .ZN(
        n12974) );
  NOR2_X1 U16075 ( .A1(n12971), .A2(n12974), .ZN(n12976) );
  NOR2_X1 U16076 ( .A1(n17823), .A2(n17824), .ZN(n12973) );
  NOR2_X1 U16077 ( .A1(n12975), .A2(n12974), .ZN(n12972) );
  AOI211_X1 U16078 ( .C1(n12975), .C2(n12974), .A(n12973), .B(n12972), .ZN(
        n17804) );
  INV_X1 U16079 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18132) );
  NOR2_X1 U16080 ( .A1(n17804), .A2(n18132), .ZN(n17803) );
  NOR2_X1 U16081 ( .A1(n17909), .A2(n18042), .ZN(n17913) );
  INV_X1 U16082 ( .A(n17913), .ZN(n16417) );
  NOR2_X1 U16083 ( .A1(n15747), .A2(n16417), .ZN(n16395) );
  NAND2_X1 U16084 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16395), .ZN(
        n12977) );
  XOR2_X1 U16085 ( .A(n18844), .B(n12977), .Z(n16387) );
  NOR2_X1 U16086 ( .A1(n18252), .A2(n18247), .ZN(n13797) );
  AND2_X1 U16087 ( .A1(n12998), .A2(n18244), .ZN(n12981) );
  NAND2_X1 U16088 ( .A1(n12982), .A2(n12981), .ZN(n12988) );
  AOI21_X1 U16089 ( .B1(n12997), .B2(n12984), .A(n12983), .ZN(n12985) );
  INV_X1 U16090 ( .A(n12985), .ZN(n12987) );
  NAND2_X1 U16091 ( .A1(n18257), .A2(n12989), .ZN(n12996) );
  NOR2_X2 U16092 ( .A1(n12993), .A2(n12991), .ZN(n18690) );
  AND2_X1 U16093 ( .A1(n12995), .A2(n12994), .ZN(n18897) );
  NOR3_X1 U16094 ( .A1(n12998), .A2(n12997), .A3(n12996), .ZN(n13799) );
  NAND2_X1 U16095 ( .A1(n13000), .A2(n12999), .ZN(n15640) );
  NAND2_X2 U16096 ( .A1(n18693), .A2(n15640), .ZN(n18682) );
  NAND2_X2 U16097 ( .A1(n18057), .A2(n18673), .ZN(n18131) );
  NOR2_X4 U16098 ( .A1(n18131), .A2(n18244), .ZN(n18665) );
  NAND2_X1 U16099 ( .A1(n18665), .A2(n18206), .ZN(n18181) );
  NOR2_X1 U16100 ( .A1(n18089), .A2(n18055), .ZN(n17718) );
  NAND2_X1 U16101 ( .A1(n17718), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17717) );
  NAND2_X1 U16102 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16405), .ZN(
        n13001) );
  XOR2_X1 U16103 ( .A(n18844), .B(n13001), .Z(n16377) );
  NOR2_X1 U16104 ( .A1(n17924), .A2(n17916), .ZN(n16396) );
  INV_X1 U16105 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18147) );
  NAND4_X1 U16106 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18146) );
  NOR3_X1 U16107 ( .A1(n18132), .A2(n18147), .A3(n18146), .ZN(n18091) );
  AOI21_X1 U16108 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18195) );
  INV_X1 U16109 ( .A(n18195), .ZN(n18127) );
  NAND2_X1 U16110 ( .A1(n18091), .A2(n18127), .ZN(n18114) );
  NOR3_X1 U16111 ( .A1(n13002), .A2(n17934), .A3(n18114), .ZN(n18008) );
  NAND2_X1 U16112 ( .A1(n13003), .A2(n18008), .ZN(n13008) );
  AOI21_X1 U16113 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18691), .A(
        n18682), .ZN(n18190) );
  NAND3_X1 U16114 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18091), .ZN(n18025) );
  NOR2_X1 U16115 ( .A1(n17934), .A2(n18025), .ZN(n18006) );
  NAND2_X1 U16116 ( .A1(n13004), .A2(n18006), .ZN(n17910) );
  OAI22_X1 U16117 ( .A1(n18701), .A2(n13008), .B1(n18190), .B2(n17910), .ZN(
        n13005) );
  NAND2_X1 U16118 ( .A1(n16396), .A2(n13005), .ZN(n15654) );
  NOR4_X1 U16119 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15747), .A3(
        n15748), .A4(n15654), .ZN(n13006) );
  AOI21_X1 U16120 ( .B1(n18137), .B2(n16377), .A(n13006), .ZN(n13007) );
  OR2_X1 U16121 ( .A1(n13007), .A2(n18222), .ZN(n13015) );
  INV_X1 U16122 ( .A(n18131), .ZN(n18133) );
  NOR2_X1 U16123 ( .A1(n18222), .A2(n18133), .ZN(n18156) );
  INV_X1 U16124 ( .A(n18156), .ZN(n18208) );
  INV_X1 U16125 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18842) );
  NAND2_X1 U16126 ( .A1(n18842), .A2(n18832), .ZN(n18896) );
  OR3_X2 U16127 ( .A1(n18896), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18221) );
  INV_X1 U16128 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17923) );
  NAND2_X1 U16129 ( .A1(n16435), .A2(n18006), .ZN(n13010) );
  NOR3_X1 U16130 ( .A1(n18859), .A2(n17923), .A3(n13010), .ZN(n13012) );
  NOR2_X1 U16131 ( .A1(n16396), .A2(n18701), .ZN(n13009) );
  AND2_X1 U16132 ( .A1(n13008), .A2(n18667), .ZN(n17953) );
  AOI211_X1 U16133 ( .C1(n18682), .C2(n13010), .A(n13009), .B(n17953), .ZN(
        n13011) );
  NOR2_X2 U16134 ( .A1(n18144), .A2(n18206), .ZN(n18201) );
  INV_X1 U16135 ( .A(n18201), .ZN(n18207) );
  OAI211_X1 U16136 ( .C1(n18679), .C2(n13012), .A(n13011), .B(n18207), .ZN(
        n15660) );
  AOI22_X1 U16137 ( .A1(n18156), .A2(n15747), .B1(n18221), .B2(n15660), .ZN(
        n15750) );
  OAI21_X1 U16138 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18208), .A(
        n15750), .ZN(n13013) );
  INV_X1 U16139 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18814) );
  NOR2_X1 U16140 ( .A1(n18814), .A2(n18221), .ZN(n16384) );
  AOI21_X1 U16141 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13013), .A(
        n16384), .ZN(n13014) );
  NAND2_X1 U16142 ( .A1(n13015), .A2(n13014), .ZN(n13016) );
  NAND2_X1 U16143 ( .A1(n13018), .A2(n13017), .ZN(P3_U2831) );
  INV_X1 U16144 ( .A(n13088), .ZN(n16345) );
  NAND2_X1 U16145 ( .A1(n13019), .A2(n16345), .ZN(n13033) );
  NAND2_X1 U16146 ( .A1(n16340), .A2(n19264), .ZN(n13233) );
  INV_X1 U16147 ( .A(n13233), .ZN(n13217) );
  NAND3_X1 U16148 ( .A1(n13217), .A2(n13215), .A3(n13020), .ZN(n13032) );
  AOI21_X1 U16149 ( .B1(n13021), .B2(n13048), .A(n10401), .ZN(n13030) );
  MUX2_X1 U16150 ( .A(n16363), .B(n13020), .S(n13446), .Z(n13022) );
  NAND2_X1 U16151 ( .A1(n13022), .A2(n16356), .ZN(n13028) );
  NAND2_X1 U16152 ( .A1(n16363), .A2(n13215), .ZN(n13023) );
  OR2_X1 U16153 ( .A1(n16338), .A2(n13023), .ZN(n13027) );
  AND2_X1 U16154 ( .A1(n13025), .A2(n13024), .ZN(n13026) );
  AND2_X1 U16155 ( .A1(n13027), .A2(n13026), .ZN(n13213) );
  OAI21_X1 U16156 ( .B1(n16338), .B2(n13028), .A(n13213), .ZN(n13029) );
  AOI21_X1 U16157 ( .B1(n13233), .B2(n13030), .A(n13029), .ZN(n13031) );
  NAND3_X1 U16158 ( .A1(n13033), .A2(n13032), .A3(n13031), .ZN(n13034) );
  NOR2_X1 U16159 ( .A1(n13088), .A2(n13035), .ZN(n19993) );
  INV_X1 U16160 ( .A(n13036), .ZN(n13037) );
  OR2_X1 U16161 ( .A1(n16337), .A2(n13037), .ZN(n15603) );
  NAND2_X1 U16162 ( .A1(n15603), .A2(n13446), .ZN(n13039) );
  INV_X1 U16163 ( .A(n13038), .ZN(n15588) );
  NAND2_X1 U16164 ( .A1(n13039), .A2(n15588), .ZN(n13040) );
  NAND2_X1 U16165 ( .A1(n13089), .A2(n13040), .ZN(n16313) );
  NAND2_X1 U16166 ( .A1(n13089), .A2(n16341), .ZN(n15376) );
  INV_X1 U16167 ( .A(n12283), .ZN(n13207) );
  NAND2_X1 U16168 ( .A1(n13043), .A2(n13042), .ZN(n13055) );
  NAND2_X1 U16169 ( .A1(n13044), .A2(n19264), .ZN(n15561) );
  NAND2_X1 U16170 ( .A1(n15561), .A2(n13045), .ZN(n13046) );
  NAND2_X1 U16171 ( .A1(n13046), .A2(n14108), .ZN(n13052) );
  OAI22_X1 U16172 ( .A1(n12283), .A2(n10401), .B1(n13048), .B2(n13047), .ZN(
        n13049) );
  INV_X1 U16173 ( .A(n13049), .ZN(n13051) );
  NAND3_X1 U16174 ( .A1(n13052), .A2(n13051), .A3(n13050), .ZN(n13053) );
  AOI21_X1 U16175 ( .B1(n13055), .B2(n13054), .A(n13053), .ZN(n15593) );
  NAND2_X1 U16176 ( .A1(n15593), .A2(n15587), .ZN(n13057) );
  NAND2_X1 U16177 ( .A1(n13089), .A2(n13057), .ZN(n13301) );
  NOR2_X1 U16178 ( .A1(n13089), .A2(n19235), .ZN(n13276) );
  INV_X1 U16179 ( .A(n13276), .ZN(n13299) );
  NAND2_X1 U16180 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13082) );
  INV_X1 U16181 ( .A(n13082), .ZN(n14178) );
  INV_X1 U16182 ( .A(n15376), .ZN(n13319) );
  INV_X1 U16183 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15560) );
  NOR2_X1 U16184 ( .A1(n15560), .A2(n15580), .ZN(n13300) );
  INV_X1 U16185 ( .A(n13300), .ZN(n13322) );
  NAND3_X1 U16186 ( .A1(n13319), .A2(n13058), .A3(n13322), .ZN(n13309) );
  INV_X1 U16187 ( .A(n13301), .ZN(n15378) );
  NAND2_X1 U16188 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13300), .ZN(
        n13312) );
  NAND2_X1 U16189 ( .A1(n15378), .A2(n13312), .ZN(n13321) );
  NAND4_X1 U16190 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13309), .A3(
        n13299), .A4(n13321), .ZN(n15554) );
  INV_X1 U16191 ( .A(n13069), .ZN(n13067) );
  NAND2_X1 U16192 ( .A1(n15554), .A2(n13067), .ZN(n14182) );
  OAI21_X1 U16193 ( .B1(n13069), .B2(n14178), .A(n14182), .ZN(n15533) );
  NAND2_X1 U16194 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15507) );
  INV_X1 U16195 ( .A(n15507), .ZN(n13059) );
  AND2_X1 U16196 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13059), .ZN(
        n13060) );
  NOR2_X1 U16197 ( .A1(n13069), .A2(n13060), .ZN(n13061) );
  NOR2_X1 U16198 ( .A1(n15533), .A2(n13061), .ZN(n15453) );
  INV_X1 U16199 ( .A(n15375), .ZN(n13063) );
  NOR3_X1 U16200 ( .A1(n13063), .A2(n16183), .A3(n13062), .ZN(n15362) );
  NAND3_X1 U16201 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n15362), .ZN(n15354) );
  NOR2_X1 U16202 ( .A1(n15189), .A2(n15354), .ZN(n13083) );
  OR2_X1 U16203 ( .A1(n16290), .A2(n13083), .ZN(n13064) );
  NAND2_X1 U16204 ( .A1(n15453), .A2(n13064), .ZN(n15357) );
  NAND2_X1 U16205 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15322) );
  INV_X1 U16206 ( .A(n15322), .ZN(n13065) );
  NOR2_X1 U16207 ( .A1(n16290), .A2(n13065), .ZN(n13066) );
  NAND2_X1 U16208 ( .A1(n15311), .A2(n13067), .ZN(n15304) );
  NAND2_X1 U16209 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15288) );
  INV_X1 U16210 ( .A(n15288), .ZN(n13068) );
  OR2_X1 U16211 ( .A1(n13069), .A2(n13068), .ZN(n13070) );
  AND2_X1 U16212 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13084) );
  NAND2_X1 U16213 ( .A1(n15248), .A2(n13084), .ZN(n15250) );
  INV_X1 U16214 ( .A(n16290), .ZN(n15413) );
  INV_X1 U16215 ( .A(n15248), .ZN(n15280) );
  OAI22_X1 U16216 ( .A1(n15250), .A2(n15251), .B1(n15413), .B2(n15280), .ZN(
        n14315) );
  OAI21_X1 U16217 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16290), .A(
        n14315), .ZN(n13071) );
  NAND2_X1 U16218 ( .A1(n13071), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13086) );
  AOI222_X1 U16219 ( .A1(n9798), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n13072), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n10665), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13073) );
  INV_X1 U16220 ( .A(n13073), .ZN(n13074) );
  NOR2_X1 U16221 ( .A1(n13077), .A2(n13076), .ZN(n16339) );
  AND2_X1 U16222 ( .A1(n16337), .A2(n19264), .ZN(n13078) );
  OR2_X1 U16223 ( .A1(n16339), .A2(n13078), .ZN(n13079) );
  NOR2_X1 U16224 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13300), .ZN(
        n13081) );
  AOI211_X1 U16225 ( .C1(n15376), .C2(n13312), .A(n13081), .B(n16290), .ZN(
        n15555) );
  NAND2_X1 U16226 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15555), .ZN(
        n14177) );
  NAND2_X1 U16227 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15539), .ZN(
        n15528) );
  NAND2_X1 U16228 ( .A1(n13083), .A2(n15488), .ZN(n15344) );
  NOR2_X1 U16229 ( .A1(n15322), .A2(n15344), .ZN(n15312) );
  NAND2_X1 U16230 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15312), .ZN(
        n15287) );
  NOR2_X1 U16231 ( .A1(n15288), .A2(n15287), .ZN(n15261) );
  NAND2_X1 U16232 ( .A1(n13084), .A2(n15261), .ZN(n15253) );
  INV_X1 U16233 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14314) );
  NOR4_X1 U16234 ( .A1(n15253), .A2(n15251), .A3(n14314), .A4(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13085) );
  INV_X1 U16235 ( .A(n16362), .ZN(n13087) );
  NOR2_X1 U16236 ( .A1(n13088), .A2(n13087), .ZN(n19992) );
  AND2_X2 U16237 ( .A1(n13089), .A2(n19992), .ZN(n16294) );
  NAND2_X1 U16238 ( .A1(n13090), .A2(n16294), .ZN(n13091) );
  OAI211_X1 U16239 ( .C1(n13093), .C2(n16287), .A(n13092), .B(n13091), .ZN(
        P2_U3015) );
  INV_X1 U16240 ( .A(n14568), .ZN(n14512) );
  AND2_X1 U16241 ( .A1(n11046), .A2(n13644), .ZN(n13097) );
  NAND2_X1 U16242 ( .A1(n13531), .A2(n13097), .ZN(n13392) );
  INV_X1 U16243 ( .A(n11231), .ZN(n20221) );
  NAND3_X1 U16244 ( .A1(n20221), .A2(n20202), .A3(n11032), .ZN(n13568) );
  INV_X1 U16245 ( .A(n13568), .ZN(n13098) );
  NAND4_X1 U16246 ( .A1(n13098), .A2(n20209), .A3(n13397), .A4(n13644), .ZN(
        n13099) );
  AOI21_X4 U16247 ( .B1(n13364), .B2(n13099), .A(n20005), .ZN(n14492) );
  NAND2_X2 U16248 ( .A1(n14492), .A2(n11231), .ZN(n14503) );
  INV_X1 U16249 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13101) );
  NAND2_X1 U16250 ( .A1(n13131), .A2(n13101), .ZN(n13103) );
  INV_X1 U16251 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21056) );
  NAND2_X1 U16252 ( .A1(n13644), .A2(n21056), .ZN(n13102) );
  NAND3_X1 U16253 ( .A1(n13103), .A2(n14326), .A3(n13102), .ZN(n13105) );
  NAND2_X1 U16254 ( .A1(n13296), .A2(n21056), .ZN(n13104) );
  NAND2_X1 U16255 ( .A1(n13105), .A2(n13104), .ZN(n13108) );
  NAND2_X1 U16256 ( .A1(n13131), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13107) );
  INV_X1 U16257 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14016) );
  NAND2_X1 U16258 ( .A1(n14326), .A2(n14016), .ZN(n13106) );
  NAND2_X1 U16259 ( .A1(n13107), .A2(n13106), .ZN(n13553) );
  XNOR2_X1 U16260 ( .A(n13108), .B(n13553), .ZN(n13645) );
  NAND2_X1 U16261 ( .A1(n13645), .A2(n13644), .ZN(n13647) );
  NAND2_X1 U16262 ( .A1(n13647), .A2(n13108), .ZN(n13596) );
  NAND2_X1 U16263 ( .A1(n13131), .A2(n13109), .ZN(n13111) );
  INV_X1 U16264 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13112) );
  NAND2_X1 U16265 ( .A1(n13644), .A2(n13112), .ZN(n13110) );
  NAND3_X1 U16266 ( .A1(n13111), .A2(n14326), .A3(n13110), .ZN(n13114) );
  NAND2_X1 U16267 ( .A1(n13296), .A2(n13112), .ZN(n13113) );
  AND2_X1 U16268 ( .A1(n13114), .A2(n13113), .ZN(n13595) );
  MUX2_X1 U16269 ( .A(n13168), .B(n14326), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13116) );
  OAI21_X1 U16270 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14324), .A(
        n13116), .ZN(n13678) );
  MUX2_X1 U16271 ( .A(n14326), .B(n13131), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13118) );
  NAND2_X1 U16272 ( .A1(n15709), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13117) );
  NAND2_X1 U16273 ( .A1(n13118), .A2(n13117), .ZN(n13771) );
  NAND2_X1 U16274 ( .A1(n14326), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13119) );
  OAI211_X1 U16275 ( .C1(n15709), .C2(P1_EBX_REG_5__SCAN_IN), .A(n13131), .B(
        n13119), .ZN(n13120) );
  OAI21_X1 U16276 ( .B1(n13168), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13120), .ZN(
        n13894) );
  MUX2_X1 U16277 ( .A(n14326), .B(n13131), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13122) );
  NAND2_X1 U16278 ( .A1(n15709), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13121) );
  NAND2_X1 U16279 ( .A1(n14326), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13123) );
  OAI211_X1 U16280 ( .C1(n15709), .C2(P1_EBX_REG_7__SCAN_IN), .A(n13131), .B(
        n13123), .ZN(n13124) );
  OAI21_X1 U16281 ( .B1(n13168), .B2(P1_EBX_REG_7__SCAN_IN), .A(n13124), .ZN(
        n16063) );
  MUX2_X1 U16282 ( .A(n14326), .B(n13131), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13126) );
  NAND2_X1 U16283 ( .A1(n15709), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13125) );
  NAND2_X1 U16284 ( .A1(n13126), .A2(n13125), .ZN(n14045) );
  INV_X1 U16285 ( .A(n13168), .ZN(n13127) );
  INV_X1 U16286 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20921) );
  NAND2_X1 U16287 ( .A1(n13127), .A2(n20921), .ZN(n13130) );
  NAND2_X1 U16288 ( .A1(n14326), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13128) );
  OAI211_X1 U16289 ( .C1(n15709), .C2(P1_EBX_REG_9__SCAN_IN), .A(n13131), .B(
        n13128), .ZN(n13129) );
  INV_X1 U16290 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15939) );
  NAND2_X1 U16291 ( .A1(n13131), .A2(n15939), .ZN(n13133) );
  INV_X1 U16292 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15859) );
  NAND2_X1 U16293 ( .A1(n13644), .A2(n15859), .ZN(n13132) );
  NAND3_X1 U16294 ( .A1(n13133), .A2(n14326), .A3(n13132), .ZN(n13135) );
  NAND2_X1 U16295 ( .A1(n13296), .A2(n15859), .ZN(n13134) );
  AND2_X1 U16296 ( .A1(n13135), .A2(n13134), .ZN(n14154) );
  MUX2_X1 U16297 ( .A(n13168), .B(n14326), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13136) );
  OAI21_X1 U16298 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14324), .A(
        n13136), .ZN(n14214) );
  MUX2_X1 U16299 ( .A(n14326), .B(n13131), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13138) );
  NAND2_X1 U16300 ( .A1(n15709), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13137) );
  NAND2_X1 U16301 ( .A1(n13138), .A2(n13137), .ZN(n14238) );
  MUX2_X1 U16302 ( .A(n13168), .B(n14326), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13139) );
  OAI21_X1 U16303 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14324), .A(
        n13139), .ZN(n14790) );
  NAND2_X1 U16304 ( .A1(n13131), .A2(n14775), .ZN(n13141) );
  INV_X1 U16305 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13142) );
  NAND2_X1 U16306 ( .A1(n13644), .A2(n13142), .ZN(n13140) );
  NAND3_X1 U16307 ( .A1(n13141), .A2(n14326), .A3(n13140), .ZN(n13144) );
  NAND2_X1 U16308 ( .A1(n13296), .A2(n13142), .ZN(n13143) );
  AND2_X1 U16309 ( .A1(n13144), .A2(n13143), .ZN(n14251) );
  MUX2_X1 U16310 ( .A(n13168), .B(n14326), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13145) );
  OAI21_X1 U16311 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14324), .A(
        n13145), .ZN(n15824) );
  MUX2_X1 U16312 ( .A(n14326), .B(n13131), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13147) );
  NAND2_X1 U16313 ( .A1(n15709), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13146) );
  NAND2_X1 U16314 ( .A1(n13147), .A2(n13146), .ZN(n14448) );
  MUX2_X1 U16315 ( .A(n13168), .B(n14326), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13148) );
  OAI21_X1 U16316 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n14324), .A(
        n13148), .ZN(n15811) );
  NAND2_X1 U16317 ( .A1(n13131), .A2(n14782), .ZN(n13150) );
  INV_X1 U16318 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21008) );
  NAND2_X1 U16319 ( .A1(n13644), .A2(n21008), .ZN(n13149) );
  NAND3_X1 U16320 ( .A1(n13150), .A2(n13115), .A3(n13149), .ZN(n13152) );
  NAND2_X1 U16321 ( .A1(n13296), .A2(n21008), .ZN(n13151) );
  NOR2_X2 U16322 ( .A1(n15814), .A2(n14498), .ZN(n14497) );
  MUX2_X1 U16323 ( .A(n13168), .B(n14326), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n13154) );
  OR2_X1 U16324 ( .A1(n14324), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13153) );
  NAND2_X1 U16325 ( .A1(n13154), .A2(n13153), .ZN(n15795) );
  INV_X1 U16326 ( .A(n15795), .ZN(n13155) );
  MUX2_X1 U16327 ( .A(n14326), .B(n13131), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13157) );
  NAND2_X1 U16328 ( .A1(n15709), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13156) );
  NAND2_X1 U16329 ( .A1(n13157), .A2(n13156), .ZN(n14491) );
  MUX2_X1 U16330 ( .A(n13168), .B(n14326), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13158) );
  OAI21_X1 U16331 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14324), .A(
        n13158), .ZN(n15736) );
  MUX2_X1 U16332 ( .A(n14326), .B(n13131), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13160) );
  NAND2_X1 U16333 ( .A1(n15709), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13159) );
  AND2_X1 U16334 ( .A1(n13160), .A2(n13159), .ZN(n14435) );
  MUX2_X1 U16335 ( .A(n13168), .B(n13115), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13162) );
  OR2_X1 U16336 ( .A1(n14324), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13161) );
  AND2_X1 U16337 ( .A1(n13162), .A2(n13161), .ZN(n14423) );
  INV_X1 U16338 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15985) );
  NAND2_X1 U16339 ( .A1(n13131), .A2(n15985), .ZN(n13163) );
  OAI211_X1 U16340 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n15709), .A(n13163), .B(
        n14326), .ZN(n13165) );
  INV_X1 U16341 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21128) );
  NAND2_X1 U16342 ( .A1(n13296), .A2(n21128), .ZN(n13164) );
  NAND2_X1 U16343 ( .A1(n13165), .A2(n13164), .ZN(n14412) );
  NAND2_X1 U16344 ( .A1(n13115), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13166) );
  OAI211_X1 U16345 ( .C1(n15709), .C2(P1_EBX_REG_25__SCAN_IN), .A(n13131), .B(
        n13166), .ZN(n13167) );
  OAI21_X1 U16346 ( .B1(n13168), .B2(P1_EBX_REG_25__SCAN_IN), .A(n13167), .ZN(
        n14398) );
  OR2_X2 U16347 ( .A1(n14414), .A2(n14398), .ZN(n14399) );
  MUX2_X1 U16348 ( .A(n13168), .B(n13115), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13170) );
  OR2_X1 U16349 ( .A1(n14324), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13169) );
  AND2_X1 U16350 ( .A1(n13170), .A2(n13169), .ZN(n14375) );
  NAND2_X1 U16351 ( .A1(n13131), .A2(n14594), .ZN(n13172) );
  INV_X1 U16352 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14483) );
  NAND2_X1 U16353 ( .A1(n13644), .A2(n14483), .ZN(n13171) );
  NAND3_X1 U16354 ( .A1(n13172), .A2(n14326), .A3(n13171), .ZN(n13174) );
  NAND2_X1 U16355 ( .A1(n13296), .A2(n14483), .ZN(n13173) );
  NAND2_X1 U16356 ( .A1(n13174), .A2(n13173), .ZN(n14386) );
  NAND2_X1 U16357 ( .A1(n14375), .A2(n14386), .ZN(n13175) );
  MUX2_X1 U16358 ( .A(n13115), .B(n13131), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13177) );
  NAND2_X1 U16359 ( .A1(n15709), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13176) );
  NAND2_X1 U16360 ( .A1(n13177), .A2(n13176), .ZN(n14360) );
  OR2_X1 U16361 ( .A1(n14324), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13179) );
  INV_X1 U16362 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n20919) );
  NAND2_X1 U16363 ( .A1(n13644), .A2(n20919), .ZN(n13178) );
  NAND2_X1 U16364 ( .A1(n13179), .A2(n13178), .ZN(n13186) );
  MUX2_X1 U16365 ( .A(P1_EBX_REG_29__SCAN_IN), .B(n13186), .S(n13115), .Z(
        n13180) );
  NAND2_X1 U16366 ( .A1(n14362), .A2(n13180), .ZN(n13181) );
  NAND2_X1 U16367 ( .A1(n14325), .A2(n13181), .ZN(n14730) );
  AND2_X1 U16368 ( .A1(n15709), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13185) );
  AOI21_X1 U16369 ( .B1(n14324), .B2(P1_EBX_REG_30__SCAN_IN), .A(n13185), .ZN(
        n14327) );
  OAI22_X1 U16370 ( .A1(n10141), .A2(n14326), .B1(n13186), .B2(n14362), .ZN(
        n13187) );
  XOR2_X1 U16371 ( .A(n14327), .B(n13187), .Z(n14345) );
  INV_X1 U16372 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n21024) );
  OAI21_X1 U16373 ( .B1(n14345), .B2(n15876), .A(n10247), .ZN(n13188) );
  INV_X1 U16374 ( .A(n13188), .ZN(n13189) );
  NOR2_X1 U16375 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13191) );
  NOR4_X1 U16376 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13190) );
  NAND4_X1 U16377 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13191), .A4(n13190), .ZN(n13204) );
  NOR2_X1 U16378 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13204), .ZN(n16513)
         );
  NOR4_X1 U16379 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13195) );
  NOR4_X1 U16380 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13194) );
  NOR4_X1 U16381 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13193) );
  NOR4_X1 U16382 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13192) );
  AND4_X1 U16383 ( .A1(n13195), .A2(n13194), .A3(n13193), .A4(n13192), .ZN(
        n13200) );
  NOR4_X1 U16384 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13198) );
  NOR4_X1 U16385 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13197) );
  NOR4_X1 U16386 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13196) );
  INV_X1 U16387 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20752) );
  AND4_X1 U16388 ( .A1(n13198), .A2(n13197), .A3(n13196), .A4(n20752), .ZN(
        n13199) );
  NAND2_X1 U16389 ( .A1(n13200), .A2(n13199), .ZN(n13201) );
  INV_X1 U16390 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20966) );
  INV_X1 U16391 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21156) );
  NOR4_X1 U16392 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n20966), .A4(n21156), .ZN(n13203) );
  NOR4_X1 U16393 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13202)
         );
  NAND3_X1 U16394 ( .A1(n20164), .A2(n13203), .A3(n13202), .ZN(U214) );
  NOR2_X1 U16395 ( .A1(n14105), .A2(n13204), .ZN(n16441) );
  NAND2_X1 U16396 ( .A1(n16441), .A2(U214), .ZN(U212) );
  NOR2_X1 U16397 ( .A1(n13205), .A2(n13231), .ZN(n19112) );
  INV_X1 U16398 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13206) );
  INV_X1 U16399 ( .A(n13445), .ZN(n13447) );
  NAND2_X1 U16400 ( .A1(n19945), .A2(n19855), .ZN(n18905) );
  OAI211_X1 U16401 ( .C1(n19112), .C2(n13206), .A(n13447), .B(n18905), .ZN(
        P2_U2814) );
  NOR2_X1 U16402 ( .A1(n18907), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13208)
         );
  AOI22_X1 U16403 ( .A1(n13208), .A2(n18905), .B1(n13207), .B2(n18907), .ZN(
        P2_U3612) );
  NOR2_X1 U16404 ( .A1(n13209), .A2(n13215), .ZN(n13210) );
  NAND2_X1 U16405 ( .A1(n16337), .A2(n13210), .ZN(n13211) );
  NOR2_X1 U16406 ( .A1(n16338), .A2(n13211), .ZN(n16346) );
  NOR2_X1 U16407 ( .A1(n16346), .A2(n13230), .ZN(n19990) );
  OAI21_X1 U16408 ( .B1(n13220), .B2(n19990), .A(n13212), .ZN(P2_U2819) );
  INV_X1 U16409 ( .A(n16340), .ZN(n16342) );
  NAND2_X1 U16410 ( .A1(n16342), .A2(n16339), .ZN(n13336) );
  AND3_X1 U16411 ( .A1(n13214), .A2(n13336), .A3(n13213), .ZN(n13219) );
  INV_X1 U16412 ( .A(n13231), .ZN(n13216) );
  NAND3_X1 U16413 ( .A1(n13217), .A2(n13216), .A3(n13215), .ZN(n13218) );
  NAND2_X1 U16414 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19984), .ZN(n16374) );
  OAI22_X1 U16415 ( .A1(n19979), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13220), 
        .B2(n16374), .ZN(n13221) );
  AOI21_X1 U16416 ( .B1(n16330), .B2(n16359), .A(n13221), .ZN(n15613) );
  INV_X1 U16417 ( .A(n15613), .ZN(n13229) );
  INV_X1 U16418 ( .A(n13222), .ZN(n13223) );
  NOR2_X1 U16419 ( .A1(n13224), .A2(n13223), .ZN(n13225) );
  NAND2_X1 U16420 ( .A1(n13226), .A2(n13225), .ZN(n16347) );
  OR3_X1 U16421 ( .A1(n15613), .A2(n15611), .A3(n16347), .ZN(n13227) );
  OAI21_X1 U16422 ( .B1(n13229), .B2(n13228), .A(n13227), .ZN(P2_U3595) );
  INV_X1 U16423 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15034) );
  OR2_X1 U16424 ( .A1(n13231), .A2(n13230), .ZN(n13232) );
  OAI21_X1 U16425 ( .B1(n13233), .B2(n13232), .A(n13529), .ZN(n13234) );
  OR2_X1 U16426 ( .A1(n19226), .A2(n14818), .ZN(n19188) );
  NAND2_X1 U16427 ( .A1(n19984), .A2(n18906), .ZN(n14823) );
  INV_X1 U16428 ( .A(n14823), .ZN(n19220) );
  CLKBUF_X1 U16429 ( .A(n19220), .Z(n19224) );
  NAND2_X1 U16430 ( .A1(n19226), .A2(n14823), .ZN(n19191) );
  AOI22_X1 U16431 ( .A1(n19224), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13235) );
  OAI21_X1 U16432 ( .B1(n15034), .B2(n19188), .A(n13235), .ZN(P2_U2926) );
  INV_X1 U16433 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15047) );
  AOI22_X1 U16434 ( .A1(n19224), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13236) );
  OAI21_X1 U16435 ( .B1(n15047), .B2(n19188), .A(n13236), .ZN(P2_U2928) );
  INV_X1 U16436 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U16437 ( .A1(n19224), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13237) );
  OAI21_X1 U16438 ( .B1(n13238), .B2(n19188), .A(n13237), .ZN(P2_U2929) );
  INV_X1 U16439 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15057) );
  AOI22_X1 U16440 ( .A1(n19224), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13239) );
  OAI21_X1 U16441 ( .B1(n15057), .B2(n19188), .A(n13239), .ZN(P2_U2930) );
  INV_X1 U16442 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14203) );
  AOI22_X1 U16443 ( .A1(n19224), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13240) );
  OAI21_X1 U16444 ( .B1(n14203), .B2(n19188), .A(n13240), .ZN(P2_U2934) );
  INV_X1 U16445 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15064) );
  AOI22_X1 U16446 ( .A1(n19224), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13241) );
  OAI21_X1 U16447 ( .B1(n15064), .B2(n19188), .A(n13241), .ZN(P2_U2932) );
  INV_X1 U16448 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13530) );
  AOI22_X1 U16449 ( .A1(n19224), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13242) );
  OAI21_X1 U16450 ( .B1(n13530), .B2(n19188), .A(n13242), .ZN(P2_U2925) );
  INV_X1 U16451 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U16452 ( .A1(n19224), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13243) );
  OAI21_X1 U16453 ( .B1(n15021), .B2(n19188), .A(n13243), .ZN(P2_U2924) );
  INV_X1 U16454 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U16455 ( .A1(n19224), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13244) );
  OAI21_X1 U16456 ( .B1(n14125), .B2(n19188), .A(n13244), .ZN(P2_U2935) );
  INV_X1 U16457 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13526) );
  AOI22_X1 U16458 ( .A1(n19224), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13245) );
  OAI21_X1 U16459 ( .B1(n13526), .B2(n19188), .A(n13245), .ZN(P2_U2923) );
  INV_X1 U16460 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16461 ( .A1(n19224), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13246) );
  OAI21_X1 U16462 ( .B1(n13247), .B2(n19188), .A(n13246), .ZN(P2_U2931) );
  INV_X1 U16463 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13249) );
  AOI22_X1 U16464 ( .A1(n19224), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13248) );
  OAI21_X1 U16465 ( .B1(n13249), .B2(n19188), .A(n13248), .ZN(P2_U2922) );
  INV_X1 U16466 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13251) );
  AOI22_X1 U16467 ( .A1(n19224), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13250) );
  OAI21_X1 U16468 ( .B1(n13251), .B2(n19188), .A(n13250), .ZN(P2_U2933) );
  INV_X1 U16469 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13514) );
  AOI22_X1 U16470 ( .A1(n19224), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13252) );
  OAI21_X1 U16471 ( .B1(n13514), .B2(n19188), .A(n13252), .ZN(P2_U2927) );
  OR3_X1 U16472 ( .A1(n13257), .A2(n13256), .A3(n13255), .ZN(n13258) );
  NAND2_X1 U16473 ( .A1(n13259), .A2(n13258), .ZN(n13260) );
  NAND2_X1 U16474 ( .A1(n13261), .A2(n13260), .ZN(n15697) );
  NAND2_X1 U16475 ( .A1(n13254), .A2(n15697), .ZN(n15705) );
  INV_X1 U16476 ( .A(n13295), .ZN(n13263) );
  INV_X1 U16477 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21188) );
  NAND2_X1 U16478 ( .A1(n20688), .A2(n16083), .ZN(n20008) );
  OAI211_X1 U16479 ( .C1(n13263), .C2(n21188), .A(n13431), .B(n20008), .ZN(
        P1_U2801) );
  NAND2_X1 U16480 ( .A1(n13264), .A2(n15560), .ZN(n13265) );
  AND2_X1 U16481 ( .A1(n13266), .A2(n13265), .ZN(n13287) );
  NAND2_X1 U16482 ( .A1(n19104), .A2(n15560), .ZN(n13267) );
  NAND2_X1 U16483 ( .A1(n13278), .A2(n13267), .ZN(n13290) );
  NAND2_X1 U16484 ( .A1(n19076), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13288) );
  OAI21_X1 U16485 ( .B1(n19237), .B2(n13290), .A(n13288), .ZN(n13268) );
  AOI21_X1 U16486 ( .B1(n19248), .B2(n13287), .A(n13268), .ZN(n13271) );
  OAI21_X1 U16487 ( .B1(n19245), .B2(n13269), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13270) );
  OAI211_X1 U16488 ( .C1(n14106), .C2(n19110), .A(n13271), .B(n13270), .ZN(
        P2_U3014) );
  OAI211_X1 U16489 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15413), .B(n13322), .ZN(n13283) );
  AOI21_X1 U16490 ( .B1(n15580), .B2(n13273), .A(n13272), .ZN(n13329) );
  AND2_X1 U16491 ( .A1(n19076), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13327) );
  AOI21_X1 U16492 ( .B1(n16294), .B2(n13329), .A(n13327), .ZN(n13282) );
  OAI21_X1 U16493 ( .B1(n13275), .B2(n13274), .A(n10662), .ZN(n19976) );
  AOI22_X1 U16494 ( .A1(n13276), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16307), .B2(n19976), .ZN(n13281) );
  OAI21_X1 U16495 ( .B1(n14882), .B2(n13278), .A(n13277), .ZN(n13279) );
  XOR2_X1 U16496 ( .A(n13279), .B(n15580), .Z(n13328) );
  NAND2_X1 U16497 ( .A1(n16318), .A2(n13328), .ZN(n13280) );
  AND4_X1 U16498 ( .A1(n13283), .A2(n13282), .A3(n13281), .A4(n13280), .ZN(
        n13284) );
  OAI21_X1 U16499 ( .B1(n9970), .B2(n16313), .A(n13284), .ZN(P2_U3045) );
  XNOR2_X1 U16500 ( .A(n13286), .B(n13285), .ZN(n13662) );
  INV_X1 U16501 ( .A(n13662), .ZN(n19183) );
  AOI22_X1 U16502 ( .A1(n16294), .A2(n13287), .B1(n16307), .B2(n19183), .ZN(
        n13289) );
  OAI211_X1 U16503 ( .C1(n16313), .C2(n19110), .A(n13289), .B(n13288), .ZN(
        n13292) );
  OAI22_X1 U16504 ( .A1(n15560), .A2(n13299), .B1(n16287), .B2(n13290), .ZN(
        n13291) );
  AOI211_X1 U16505 ( .C1(n15560), .C2(n15413), .A(n13292), .B(n13291), .ZN(
        n13293) );
  INV_X1 U16506 ( .A(n13293), .ZN(P2_U3046) );
  INV_X1 U16507 ( .A(n20008), .ZN(n13294) );
  NOR2_X1 U16508 ( .A1(n13294), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13298)
         );
  NAND2_X2 U16509 ( .A1(n13431), .A2(n13295), .ZN(n20815) );
  OAI21_X1 U16510 ( .B1(n15708), .B2(n13296), .A(n20815), .ZN(n13297) );
  OAI21_X1 U16511 ( .B1(n13298), .B2(n20815), .A(n13297), .ZN(P1_U3487) );
  OAI21_X1 U16512 ( .B1(n13301), .B2(n13300), .A(n13299), .ZN(n13325) );
  NAND2_X1 U16513 ( .A1(n13303), .A2(n13302), .ZN(n13304) );
  NAND2_X1 U16514 ( .A1(n13305), .A2(n13304), .ZN(n19244) );
  AOI21_X1 U16515 ( .B1(n13308), .B2(n13307), .A(n13306), .ZN(n19249) );
  NAND2_X1 U16516 ( .A1(n19076), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19251) );
  NAND2_X1 U16517 ( .A1(n19251), .A2(n13309), .ZN(n13310) );
  AOI21_X1 U16518 ( .B1(n16294), .B2(n19249), .A(n13310), .ZN(n13311) );
  OAI21_X1 U16519 ( .B1(n16287), .B2(n19244), .A(n13311), .ZN(n13324) );
  INV_X1 U16520 ( .A(n13312), .ZN(n13318) );
  NAND2_X1 U16521 ( .A1(n13314), .A2(n13313), .ZN(n13317) );
  INV_X1 U16522 ( .A(n13315), .ZN(n13316) );
  AND2_X1 U16523 ( .A1(n13317), .A2(n13316), .ZN(n19962) );
  INV_X1 U16524 ( .A(n19962), .ZN(n13667) );
  AOI22_X1 U16525 ( .A1(n13319), .A2(n13318), .B1(n16307), .B2(n13667), .ZN(
        n13320) );
  OAI21_X1 U16526 ( .B1(n13322), .B2(n13321), .A(n13320), .ZN(n13323) );
  AOI211_X1 U16527 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13325), .A(
        n13324), .B(n13323), .ZN(n13326) );
  OAI21_X1 U16528 ( .B1(n15594), .B2(n16313), .A(n13326), .ZN(P2_U3044) );
  AOI21_X1 U16529 ( .B1(n13328), .B2(n19246), .A(n13327), .ZN(n13331) );
  NAND2_X1 U16530 ( .A1(n19248), .A2(n13329), .ZN(n13330) );
  OAI211_X1 U16531 ( .C1(n16275), .C2(n14883), .A(n13331), .B(n13330), .ZN(
        n13332) );
  AOI21_X1 U16532 ( .B1(n16268), .B2(n14883), .A(n13332), .ZN(n13333) );
  OAI21_X1 U16533 ( .B1(n9970), .B2(n14106), .A(n13333), .ZN(P2_U3013) );
  NAND2_X1 U16534 ( .A1(n13336), .A2(n15587), .ZN(n13337) );
  INV_X1 U16535 ( .A(n14998), .ZN(n14962) );
  NAND2_X1 U16536 ( .A1(n14962), .A2(n19292), .ZN(n15000) );
  MUX2_X1 U16537 ( .A(n13338), .B(n9970), .S(n14962), .Z(n13339) );
  OAI21_X1 U16538 ( .B1(n19971), .B2(n15000), .A(n13339), .ZN(P2_U2886) );
  NAND2_X1 U16539 ( .A1(n19264), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13340) );
  AND4_X1 U16540 ( .A1(n13668), .A2(n13340), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19979), .ZN(n13341) );
  MUX2_X1 U16541 ( .A(n19110), .B(n13343), .S(n14980), .Z(n13344) );
  OAI21_X1 U16542 ( .B1(n19981), .B2(n15000), .A(n13344), .ZN(P2_U2887) );
  OR2_X1 U16543 ( .A1(n15704), .A2(n11036), .ZN(n13551) );
  INV_X1 U16544 ( .A(n13551), .ZN(n13347) );
  INV_X1 U16545 ( .A(n13345), .ZN(n13346) );
  INV_X1 U16546 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20003) );
  NAND2_X1 U16547 ( .A1(n13346), .A2(n20003), .ZN(n15756) );
  INV_X1 U16548 ( .A(n15756), .ZN(n20821) );
  NAND2_X1 U16549 ( .A1(n13347), .A2(n20821), .ZN(n15719) );
  AND2_X1 U16550 ( .A1(n13254), .A2(n11036), .ZN(n15675) );
  NAND2_X1 U16551 ( .A1(n15675), .A2(n20821), .ZN(n13370) );
  NAND2_X1 U16552 ( .A1(n15719), .A2(n13370), .ZN(n13348) );
  NAND2_X1 U16553 ( .A1(n20118), .A2(n13557), .ZN(n13631) );
  NOR2_X1 U16554 ( .A1(n16083), .A2(n20813), .ZN(n13761) );
  INV_X1 U16555 ( .A(n13761), .ZN(n16084) );
  OR2_X1 U16556 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16084), .ZN(n20116) );
  INV_X2 U16557 ( .A(n20116), .ZN(n20141) );
  NOR2_X4 U16558 ( .A1(n20118), .A2(n20141), .ZN(n15757) );
  AOI22_X1 U16559 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13349) );
  OAI21_X1 U16560 ( .B1(n11493), .B2(n13631), .A(n13349), .ZN(P1_U2917) );
  AOI22_X1 U16561 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13350) );
  OAI21_X1 U16562 ( .B1(n11581), .B2(n13631), .A(n13350), .ZN(P1_U2913) );
  AOI22_X1 U16563 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13351) );
  OAI21_X1 U16564 ( .B1(n11606), .B2(n13631), .A(n13351), .ZN(P1_U2912) );
  AOI22_X1 U16565 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13352) );
  OAI21_X1 U16566 ( .B1(n11478), .B2(n13631), .A(n13352), .ZN(P1_U2918) );
  AOI22_X1 U16567 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13353) );
  OAI21_X1 U16568 ( .B1(n11717), .B2(n13631), .A(n13353), .ZN(P1_U2907) );
  INV_X1 U16569 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13355) );
  AOI22_X1 U16570 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13354) );
  OAI21_X1 U16571 ( .B1(n13355), .B2(n13631), .A(n13354), .ZN(P1_U2920) );
  AOI22_X1 U16572 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13356) );
  OAI21_X1 U16573 ( .B1(n11695), .B2(n13631), .A(n13356), .ZN(P1_U2908) );
  AOI22_X1 U16574 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13357) );
  OAI21_X1 U16575 ( .B1(n11671), .B2(n13631), .A(n13357), .ZN(P1_U2909) );
  INV_X1 U16576 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13359) );
  AOI22_X1 U16577 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13358) );
  OAI21_X1 U16578 ( .B1(n13359), .B2(n13631), .A(n13358), .ZN(P1_U2919) );
  AOI22_X1 U16579 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13360) );
  OAI21_X1 U16580 ( .B1(n21141), .B2(n13631), .A(n13360), .ZN(P1_U2911) );
  MUX2_X1 U16581 ( .A(n10878), .B(n15594), .S(n14962), .Z(n13363) );
  OAI21_X1 U16582 ( .B1(n19961), .B2(n15000), .A(n13363), .ZN(P2_U2885) );
  INV_X1 U16583 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20579) );
  INV_X1 U16584 ( .A(n13364), .ZN(n13380) );
  NAND2_X1 U16585 ( .A1(n11046), .A2(n15708), .ZN(n13365) );
  NOR2_X1 U16586 ( .A1(n13365), .A2(n14806), .ZN(n15693) );
  NAND2_X1 U16587 ( .A1(n15707), .A2(n15693), .ZN(n13368) );
  NAND2_X1 U16588 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20820) );
  NAND2_X1 U16589 ( .A1(n20820), .A2(n15697), .ZN(n13532) );
  OR2_X1 U16590 ( .A1(n13366), .A2(n13532), .ZN(n13367) );
  NAND2_X1 U16591 ( .A1(n13368), .A2(n13367), .ZN(n13571) );
  NOR2_X1 U16592 ( .A1(n13644), .A2(n20821), .ZN(n13371) );
  OAI21_X1 U16593 ( .B1(n13371), .B2(n13369), .A(n13370), .ZN(n13373) );
  NAND2_X1 U16594 ( .A1(n15707), .A2(n20820), .ZN(n15720) );
  INV_X1 U16595 ( .A(n15720), .ZN(n13372) );
  NAND2_X1 U16596 ( .A1(n13373), .A2(n13372), .ZN(n13378) );
  INV_X1 U16597 ( .A(n13254), .ZN(n13377) );
  OAI21_X1 U16598 ( .B1(n11049), .B2(n20183), .A(n13557), .ZN(n13374) );
  NOR2_X1 U16599 ( .A1(n13375), .A2(n13374), .ZN(n13388) );
  AOI21_X1 U16600 ( .B1(n13377), .B2(n13376), .A(n13388), .ZN(n13536) );
  OAI211_X1 U16601 ( .C1(n20822), .C2(n13540), .A(n13378), .B(n13536), .ZN(
        n13379) );
  NOR2_X1 U16602 ( .A1(n20169), .A2(n16084), .ZN(n13760) );
  AOI22_X1 U16603 ( .A1(n20011), .A2(n15680), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n13760), .ZN(n16079) );
  OAI21_X1 U16604 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20579), .A(n16079), 
        .ZN(n16076) );
  INV_X1 U16605 ( .A(n16076), .ZN(n20801) );
  AND2_X1 U16606 ( .A1(n13383), .A2(n14324), .ZN(n13387) );
  INV_X1 U16607 ( .A(n20822), .ZN(n14004) );
  OAI21_X1 U16608 ( .B1(n10166), .B2(n13397), .A(n14004), .ZN(n13385) );
  OAI21_X1 U16609 ( .B1(n11040), .B2(n13557), .A(n13540), .ZN(n13384) );
  NAND2_X1 U16610 ( .A1(n13385), .A2(n13384), .ZN(n13386) );
  OR3_X1 U16611 ( .A1(n13388), .A2(n13387), .A3(n13386), .ZN(n13390) );
  AND2_X1 U16612 ( .A1(n11048), .A2(n15708), .ZN(n13389) );
  NOR2_X1 U16613 ( .A1(n13390), .A2(n13389), .ZN(n13556) );
  AND3_X1 U16614 ( .A1(n13369), .A2(n13746), .A3(n13558), .ZN(n13391) );
  AND3_X1 U16615 ( .A1(n13556), .A2(n13391), .A3(n13366), .ZN(n14807) );
  INV_X1 U16616 ( .A(n13751), .ZN(n13394) );
  XNOR2_X1 U16617 ( .A(n13394), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13396) );
  INV_X1 U16618 ( .A(n13392), .ZN(n15699) );
  OR2_X1 U16619 ( .A1(n15699), .A2(n15693), .ZN(n13742) );
  XNOR2_X1 U16620 ( .A(n13393), .B(n13394), .ZN(n13400) );
  INV_X1 U16621 ( .A(n13400), .ZN(n13395) );
  AOI22_X1 U16622 ( .A1(n15675), .A2(n13396), .B1(n13742), .B2(n13395), .ZN(
        n13399) );
  AND2_X1 U16623 ( .A1(n13556), .A2(n13397), .ZN(n13747) );
  NAND3_X1 U16624 ( .A1(n13747), .A2(n13400), .A3(n13746), .ZN(n13398) );
  OAI211_X1 U16625 ( .C1(n13382), .C2(n14807), .A(n13399), .B(n13398), .ZN(
        n13750) );
  INV_X1 U16626 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13648) );
  NOR2_X1 U16627 ( .A1(n16083), .A2(n13648), .ZN(n14813) );
  OAI22_X1 U16628 ( .A1(n10114), .A2(n13101), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14814) );
  INV_X1 U16629 ( .A(n14814), .ZN(n13401) );
  INV_X1 U16630 ( .A(n14811), .ZN(n20796) );
  AOI222_X1 U16631 ( .A1(n13750), .A2(n20798), .B1(n14813), .B2(n13401), .C1(
        n20796), .C2(n13400), .ZN(n13403) );
  NAND2_X1 U16632 ( .A1(n20801), .A2(n13751), .ZN(n13402) );
  OAI21_X1 U16633 ( .B1(n20801), .B2(n13403), .A(n13402), .ZN(P1_U3472) );
  INV_X1 U16634 ( .A(n13404), .ZN(n13405) );
  XNOR2_X1 U16635 ( .A(n13406), .B(n13405), .ZN(n14019) );
  INV_X1 U16636 ( .A(n14019), .ZN(n14022) );
  INV_X1 U16637 ( .A(n20166), .ZN(n15953) );
  NAND2_X1 U16638 ( .A1(n13407), .A2(n15960), .ZN(n13411) );
  INV_X1 U16639 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14021) );
  NOR2_X1 U16640 ( .A1(n20055), .A2(n14021), .ZN(n13564) );
  OAI21_X1 U16641 ( .B1(n13409), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13408), .ZN(n13567) );
  NOR2_X1 U16642 ( .A1(n13567), .A2(n15955), .ZN(n13410) );
  AOI211_X1 U16643 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13411), .A(
        n13564), .B(n13410), .ZN(n13412) );
  OAI21_X1 U16644 ( .B1(n14022), .B2(n15953), .A(n13412), .ZN(P1_U2999) );
  INV_X1 U16645 ( .A(n13414), .ZN(n13417) );
  NAND2_X1 U16646 ( .A1(n11971), .A2(n13415), .ZN(n13497) );
  INV_X1 U16647 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13422) );
  MUX2_X1 U16648 ( .A(n9804), .B(n13422), .S(n14980), .Z(n13423) );
  OAI21_X1 U16649 ( .B1(n19521), .B2(n15000), .A(n13423), .ZN(P2_U2884) );
  XNOR2_X1 U16650 ( .A(n13607), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13429) );
  NAND2_X1 U16651 ( .A1(n13425), .A2(n13609), .ZN(n13427) );
  INV_X1 U16652 ( .A(n13576), .ZN(n13426) );
  NAND2_X1 U16653 ( .A1(n13427), .A2(n13426), .ZN(n15529) );
  MUX2_X1 U16654 ( .A(n15529), .B(n10885), .S(n14980), .Z(n13428) );
  OAI21_X1 U16655 ( .B1(n13429), .B2(n15000), .A(n13428), .ZN(P2_U2880) );
  INV_X1 U16656 ( .A(n20820), .ZN(n20814) );
  AND2_X1 U16657 ( .A1(n20819), .A2(n20814), .ZN(n13430) );
  OR2_X2 U16658 ( .A1(n13431), .A2(n13430), .ZN(n20152) );
  OR2_X1 U16659 ( .A1(n20152), .A2(n11036), .ZN(n13690) );
  NAND2_X1 U16660 ( .A1(n20152), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13432) );
  NOR2_X2 U16661 ( .A1(n20152), .A2(n20183), .ZN(n13725) );
  MUX2_X1 U16662 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20164), .Z(
        n14513) );
  NAND2_X1 U16663 ( .A1(n13725), .A2(n14513), .ZN(n20148) );
  OAI211_X1 U16664 ( .C1(n13690), .C2(n11695), .A(n13432), .B(n20148), .ZN(
        P1_U2949) );
  NAND2_X1 U16665 ( .A1(n20152), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13433) );
  MUX2_X1 U16666 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20164), .Z(
        n14506) );
  NAND2_X1 U16667 ( .A1(n13725), .A2(n14506), .ZN(n20154) );
  OAI211_X1 U16668 ( .C1(n13690), .C2(n11752), .A(n13433), .B(n20154), .ZN(
        P1_U2951) );
  NAND2_X1 U16669 ( .A1(n20152), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13434) );
  MUX2_X1 U16670 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20164), .Z(
        n14509) );
  NAND2_X1 U16671 ( .A1(n13725), .A2(n14509), .ZN(n20150) );
  OAI211_X1 U16672 ( .C1(n13690), .C2(n11717), .A(n13434), .B(n20150), .ZN(
        P1_U2950) );
  NAND2_X1 U16673 ( .A1(n20152), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13435) );
  MUX2_X1 U16674 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20164), .Z(
        n14519) );
  NAND2_X1 U16675 ( .A1(n13725), .A2(n14519), .ZN(n20146) );
  OAI211_X1 U16676 ( .C1(n13690), .C2(n11652), .A(n13435), .B(n20146), .ZN(
        P1_U2947) );
  AOI21_X1 U16677 ( .B1(n20798), .B2(n15675), .A(n20801), .ZN(n13438) );
  INV_X1 U16678 ( .A(n11269), .ZN(n14008) );
  OAI22_X1 U16679 ( .A1(n14008), .A2(n14807), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14806), .ZN(n15676) );
  OAI22_X1 U16680 ( .A1(n16083), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14811), .ZN(n13436) );
  AOI21_X1 U16681 ( .B1(n15676), .B2(n20798), .A(n13436), .ZN(n13437) );
  OAI22_X1 U16682 ( .A1(n13438), .A2(n10911), .B1(n13437), .B2(n20801), .ZN(
        P1_U3474) );
  INV_X1 U16683 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14550) );
  INV_X1 U16684 ( .A(n13725), .ZN(n13441) );
  INV_X1 U16685 ( .A(DATAI_15_), .ZN(n13439) );
  NOR2_X1 U16686 ( .A1(n20164), .A2(n13439), .ZN(n13440) );
  AOI21_X1 U16687 ( .B1(n20164), .B2(BUF1_REG_15__SCAN_IN), .A(n13440), .ZN(
        n14548) );
  INV_X1 U16688 ( .A(n20152), .ZN(n13691) );
  INV_X1 U16689 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20117) );
  OAI222_X1 U16690 ( .A1(n13690), .A2(n14550), .B1(n13441), .B2(n14548), .C1(
        n13691), .C2(n20117), .ZN(P1_U2967) );
  NAND2_X1 U16691 ( .A1(n20152), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13442) );
  MUX2_X1 U16692 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20164), .Z(
        n14526) );
  NAND2_X1 U16693 ( .A1(n13725), .A2(n14526), .ZN(n13443) );
  OAI211_X1 U16694 ( .C1(n13690), .C2(n11606), .A(n13442), .B(n13443), .ZN(
        P1_U2945) );
  INV_X1 U16695 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20132) );
  NAND2_X1 U16696 ( .A1(n20152), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13444) );
  OAI211_X1 U16697 ( .C1(n13690), .C2(n20132), .A(n13444), .B(n13443), .ZN(
        P1_U2960) );
  INV_X1 U16698 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13450) );
  INV_X1 U16699 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13449) );
  OAI21_X1 U16700 ( .B1(n13446), .B2(n16356), .A(n13445), .ZN(n19231) );
  INV_X1 U16701 ( .A(n19231), .ZN(n13452) );
  INV_X1 U16702 ( .A(n19229), .ZN(n13448) );
  AOI22_X1 U16703 ( .A1(n14107), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14105), .ZN(n19124) );
  OAI222_X1 U16704 ( .A1(n13529), .A2(n13450), .B1(n13449), .B2(n13452), .C1(
        n13448), .C2(n19124), .ZN(P2_U2982) );
  AOI22_X1 U16705 ( .A1(n14107), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14105), .ZN(n19265) );
  INV_X1 U16706 ( .A(n19265), .ZN(n13451) );
  NAND2_X1 U16707 ( .A1(n19229), .A2(n13451), .ZN(n13482) );
  AOI22_X1 U16708 ( .A1(n19232), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13521), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13453) );
  NAND2_X1 U16709 ( .A1(n13482), .A2(n13453), .ZN(P2_U2968) );
  AOI22_X1 U16710 ( .A1(n14107), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14105), .ZN(n19260) );
  INV_X1 U16711 ( .A(n19260), .ZN(n13454) );
  NAND2_X1 U16712 ( .A1(n19229), .A2(n13454), .ZN(n13486) );
  AOI22_X1 U16713 ( .A1(n19232), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19231), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13455) );
  NAND2_X1 U16714 ( .A1(n13486), .A2(n13455), .ZN(P2_U2952) );
  INV_X1 U16715 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13456) );
  OR2_X1 U16716 ( .A1(n14105), .A2(n13456), .ZN(n13458) );
  NAND2_X1 U16717 ( .A1(n14105), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13457) );
  AND2_X1 U16718 ( .A1(n13458), .A2(n13457), .ZN(n19129) );
  INV_X1 U16719 ( .A(n19129), .ZN(n15008) );
  NAND2_X1 U16720 ( .A1(n19229), .A2(n15008), .ZN(n13467) );
  AOI22_X1 U16721 ( .A1(n19232), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13521), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13459) );
  NAND2_X1 U16722 ( .A1(n13467), .A2(n13459), .ZN(P2_U2965) );
  INV_X1 U16723 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16478) );
  INV_X1 U16724 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18259) );
  AOI22_X1 U16725 ( .A1(n14107), .A2(n16478), .B1(n18259), .B2(n14105), .ZN(
        n19157) );
  NAND2_X1 U16726 ( .A1(n19229), .A2(n19157), .ZN(n13475) );
  AOI22_X1 U16727 ( .A1(n19232), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13521), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13460) );
  NAND2_X1 U16728 ( .A1(n13475), .A2(n13460), .ZN(P2_U2956) );
  INV_X1 U16729 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13461) );
  OR2_X1 U16730 ( .A1(n14105), .A2(n13461), .ZN(n13463) );
  NAND2_X1 U16731 ( .A1(n14105), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13462) );
  AND2_X1 U16732 ( .A1(n13463), .A2(n13462), .ZN(n19134) );
  INV_X1 U16733 ( .A(n19134), .ZN(n13464) );
  NAND2_X1 U16734 ( .A1(n19229), .A2(n13464), .ZN(n13477) );
  AOI22_X1 U16735 ( .A1(n19232), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13521), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13465) );
  NAND2_X1 U16736 ( .A1(n13477), .A2(n13465), .ZN(P2_U2963) );
  AOI22_X1 U16737 ( .A1(n19232), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13521), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13466) );
  NAND2_X1 U16738 ( .A1(n13467), .A2(n13466), .ZN(P2_U2980) );
  AOI22_X1 U16739 ( .A1(n14107), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14105), .ZN(n19171) );
  INV_X1 U16740 ( .A(n19171), .ZN(n13468) );
  NAND2_X1 U16741 ( .A1(n19229), .A2(n13468), .ZN(n13484) );
  AOI22_X1 U16742 ( .A1(n19232), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19231), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U16743 ( .A1(n13484), .A2(n13469), .ZN(P2_U2955) );
  AOI22_X1 U16744 ( .A1(n14107), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14105), .ZN(n19294) );
  INV_X1 U16745 ( .A(n19294), .ZN(n13470) );
  NAND2_X1 U16746 ( .A1(n19229), .A2(n13470), .ZN(n13480) );
  AOI22_X1 U16747 ( .A1(n19232), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n19231), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13471) );
  NAND2_X1 U16748 ( .A1(n13480), .A2(n13471), .ZN(P2_U2974) );
  INV_X1 U16749 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16474) );
  INV_X1 U16750 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18269) );
  AOI22_X1 U16751 ( .A1(n14107), .A2(n16474), .B1(n18269), .B2(n14105), .ZN(
        n19146) );
  NAND2_X1 U16752 ( .A1(n19229), .A2(n19146), .ZN(n13490) );
  AOI22_X1 U16753 ( .A1(n19232), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13521), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13472) );
  NAND2_X1 U16754 ( .A1(n13490), .A2(n13472), .ZN(P2_U2973) );
  AOI22_X1 U16755 ( .A1(n14107), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14105), .ZN(n19278) );
  INV_X1 U16756 ( .A(n19278), .ZN(n19150) );
  NAND2_X1 U16757 ( .A1(n19229), .A2(n19150), .ZN(n13488) );
  AOI22_X1 U16758 ( .A1(n19232), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13521), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13473) );
  NAND2_X1 U16759 ( .A1(n13488), .A2(n13473), .ZN(P2_U2972) );
  AOI22_X1 U16760 ( .A1(n19232), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13521), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U16761 ( .A1(n13475), .A2(n13474), .ZN(P2_U2971) );
  AOI22_X1 U16762 ( .A1(n19232), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n19231), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13476) );
  NAND2_X1 U16763 ( .A1(n13477), .A2(n13476), .ZN(P2_U2978) );
  OAI22_X1 U16764 ( .A1(n14105), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14107), .ZN(n19269) );
  INV_X1 U16765 ( .A(n19269), .ZN(n16164) );
  NAND2_X1 U16766 ( .A1(n19229), .A2(n16164), .ZN(n13492) );
  AOI22_X1 U16767 ( .A1(n19232), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13521), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13478) );
  NAND2_X1 U16768 ( .A1(n13492), .A2(n13478), .ZN(P2_U2969) );
  AOI22_X1 U16769 ( .A1(n19232), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13521), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13479) );
  NAND2_X1 U16770 ( .A1(n13480), .A2(n13479), .ZN(P2_U2959) );
  AOI22_X1 U16771 ( .A1(n19232), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13521), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13481) );
  NAND2_X1 U16772 ( .A1(n13482), .A2(n13481), .ZN(P2_U2953) );
  AOI22_X1 U16773 ( .A1(n19232), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13521), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13483) );
  NAND2_X1 U16774 ( .A1(n13484), .A2(n13483), .ZN(P2_U2970) );
  AOI22_X1 U16775 ( .A1(n19232), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n13521), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13485) );
  NAND2_X1 U16776 ( .A1(n13486), .A2(n13485), .ZN(P2_U2967) );
  AOI22_X1 U16777 ( .A1(n19232), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13521), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13487) );
  NAND2_X1 U16778 ( .A1(n13488), .A2(n13487), .ZN(P2_U2957) );
  AOI22_X1 U16779 ( .A1(n19232), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n13521), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13489) );
  NAND2_X1 U16780 ( .A1(n13490), .A2(n13489), .ZN(P2_U2958) );
  AOI22_X1 U16781 ( .A1(n19232), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n19231), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13491) );
  NAND2_X1 U16782 ( .A1(n13492), .A2(n13491), .ZN(P2_U2954) );
  NAND2_X1 U16783 ( .A1(n14105), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13494) );
  INV_X1 U16784 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16468) );
  OR2_X1 U16785 ( .A1(n14105), .A2(n16468), .ZN(n13493) );
  NAND2_X1 U16786 ( .A1(n13494), .A2(n13493), .ZN(n19139) );
  NAND2_X1 U16787 ( .A1(n19229), .A2(n19139), .ZN(n13510) );
  AOI22_X1 U16788 ( .A1(n19232), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13521), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13495) );
  NAND2_X1 U16789 ( .A1(n13510), .A2(n13495), .ZN(P2_U2961) );
  NAND2_X1 U16790 ( .A1(n19283), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13496) );
  AND2_X1 U16791 ( .A1(n13497), .A2(n13496), .ZN(n13498) );
  NAND2_X1 U16792 ( .A1(n13499), .A2(n13498), .ZN(n13502) );
  INV_X1 U16793 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19276) );
  NOR2_X1 U16794 ( .A1(n13500), .A2(n19276), .ZN(n13501) );
  NAND2_X1 U16795 ( .A1(n13502), .A2(n13501), .ZN(n13619) );
  OR2_X1 U16796 ( .A1(n13502), .A2(n13501), .ZN(n13503) );
  NAND2_X1 U16797 ( .A1(n13619), .A2(n13503), .ZN(n19160) );
  NOR2_X1 U16798 ( .A1(n13505), .A2(n13506), .ZN(n13507) );
  OR2_X1 U16799 ( .A1(n13504), .A2(n13507), .ZN(n19236) );
  MUX2_X1 U16800 ( .A(n10877), .B(n19236), .S(n14962), .Z(n13508) );
  OAI21_X1 U16801 ( .B1(n19160), .B2(n15000), .A(n13508), .ZN(P2_U2883) );
  INV_X1 U16802 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19205) );
  NAND2_X1 U16803 ( .A1(n13521), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13509) );
  OAI211_X1 U16804 ( .C1(n19205), .C2(n13529), .A(n13510), .B(n13509), .ZN(
        P2_U2976) );
  NAND2_X1 U16805 ( .A1(n14105), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13512) );
  INV_X1 U16806 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16470) );
  OR2_X1 U16807 ( .A1(n14105), .A2(n16470), .ZN(n13511) );
  NAND2_X1 U16808 ( .A1(n13512), .A2(n13511), .ZN(n19142) );
  NAND2_X1 U16809 ( .A1(n19229), .A2(n19142), .ZN(n13523) );
  NAND2_X1 U16810 ( .A1(n19231), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13513) );
  OAI211_X1 U16811 ( .C1(n13514), .C2(n13529), .A(n13523), .B(n13513), .ZN(
        P2_U2960) );
  INV_X1 U16812 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19203) );
  NAND2_X1 U16813 ( .A1(n14105), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13516) );
  INV_X1 U16814 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16466) );
  OR2_X1 U16815 ( .A1(n14105), .A2(n16466), .ZN(n13515) );
  NAND2_X1 U16816 ( .A1(n13516), .A2(n13515), .ZN(n19136) );
  NAND2_X1 U16817 ( .A1(n19229), .A2(n19136), .ZN(n13528) );
  NAND2_X1 U16818 ( .A1(n13521), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13517) );
  OAI211_X1 U16819 ( .C1(n19203), .C2(n13529), .A(n13528), .B(n13517), .ZN(
        P2_U2977) );
  INV_X1 U16820 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19199) );
  NAND2_X1 U16821 ( .A1(n14105), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13519) );
  INV_X1 U16822 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16463) );
  OR2_X1 U16823 ( .A1(n14105), .A2(n16463), .ZN(n13518) );
  NAND2_X1 U16824 ( .A1(n13519), .A2(n13518), .ZN(n19131) );
  NAND2_X1 U16825 ( .A1(n19229), .A2(n19131), .ZN(n13525) );
  NAND2_X1 U16826 ( .A1(n13521), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13520) );
  OAI211_X1 U16827 ( .C1(n19199), .C2(n13529), .A(n13525), .B(n13520), .ZN(
        P2_U2979) );
  INV_X1 U16828 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19207) );
  NAND2_X1 U16829 ( .A1(n13521), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13522) );
  OAI211_X1 U16830 ( .C1(n19207), .C2(n13529), .A(n13523), .B(n13522), .ZN(
        P2_U2975) );
  NAND2_X1 U16831 ( .A1(n19231), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13524) );
  OAI211_X1 U16832 ( .C1(n13526), .C2(n13529), .A(n13525), .B(n13524), .ZN(
        P2_U2964) );
  NAND2_X1 U16833 ( .A1(n19231), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13527) );
  OAI211_X1 U16834 ( .C1(n13530), .C2(n13529), .A(n13528), .B(n13527), .ZN(
        P2_U2962) );
  NAND2_X1 U16835 ( .A1(n13531), .A2(n11036), .ZN(n13537) );
  NAND2_X1 U16836 ( .A1(n11036), .A2(n15756), .ZN(n13534) );
  INV_X1 U16837 ( .A(n13532), .ZN(n13533) );
  NAND3_X1 U16838 ( .A1(n13534), .A2(n13540), .A3(n13533), .ZN(n13535) );
  OAI211_X1 U16839 ( .C1(n15707), .C2(n13537), .A(n13536), .B(n13535), .ZN(
        n13538) );
  NAND2_X1 U16840 ( .A1(n13538), .A2(n20011), .ZN(n13545) );
  OAI21_X1 U16841 ( .B1(n13369), .B2(n20814), .A(n13557), .ZN(n13539) );
  OAI21_X1 U16842 ( .B1(n20821), .B2(n20819), .A(n13539), .ZN(n13541) );
  AOI21_X1 U16843 ( .B1(n13541), .B2(n11040), .A(n13540), .ZN(n13542) );
  NAND2_X1 U16844 ( .A1(n13543), .A2(n13542), .ZN(n13544) );
  INV_X1 U16845 ( .A(n13546), .ZN(n13547) );
  AOI21_X1 U16846 ( .B1(n13547), .B2(n11034), .A(n15693), .ZN(n13549) );
  INV_X1 U16847 ( .A(n15696), .ZN(n13548) );
  NAND3_X1 U16848 ( .A1(n9912), .A2(n13549), .A3(n13548), .ZN(n13550) );
  OAI21_X1 U16849 ( .B1(n13546), .B2(n11034), .A(n13551), .ZN(n13552) );
  OR2_X1 U16850 ( .A1(n14324), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13554) );
  NAND2_X1 U16851 ( .A1(n13554), .A2(n13553), .ZN(n14023) );
  INV_X1 U16852 ( .A(n14023), .ZN(n13565) );
  OAI211_X1 U16853 ( .C1(n13558), .C2(n13557), .A(n13556), .B(n13555), .ZN(
        n13559) );
  NAND2_X1 U16854 ( .A1(n13562), .A2(n13559), .ZN(n14701) );
  INV_X1 U16855 ( .A(n14706), .ZN(n13561) );
  INV_X2 U16856 ( .A(n20055), .ZN(n20070) );
  OR2_X1 U16857 ( .A1(n13562), .A2(n20070), .ZN(n13592) );
  INV_X1 U16858 ( .A(n13592), .ZN(n13560) );
  AOI21_X1 U16859 ( .B1(n13561), .B2(n13648), .A(n13560), .ZN(n13643) );
  AOI22_X1 U16860 ( .A1(n13643), .A2(n14702), .B1(n14706), .B2(n13648), .ZN(
        n13563) );
  AOI211_X1 U16861 ( .C1(n16067), .C2(n13565), .A(n13564), .B(n13563), .ZN(
        n13566) );
  OAI21_X1 U16862 ( .B1(n16052), .B2(n13567), .A(n13566), .ZN(P1_U3031) );
  OAI22_X1 U16863 ( .A1(n13569), .A2(n15720), .B1(n13746), .B2(n13568), .ZN(
        n13570) );
  NAND2_X1 U16864 ( .A1(n11049), .A2(n11231), .ZN(n13575) );
  INV_X1 U16865 ( .A(n20164), .ZN(n20165) );
  NAND2_X1 U16866 ( .A1(n20165), .A2(DATAI_0_), .ZN(n13574) );
  NAND2_X1 U16867 ( .A1(n20164), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13573) );
  AND2_X1 U16868 ( .A1(n13574), .A2(n13573), .ZN(n20163) );
  OAI222_X1 U16869 ( .A1(n14549), .A2(n20163), .B1(n15896), .B2(n14022), .C1(
        n11271), .C2(n14551), .ZN(P1_U2904) );
  OR2_X1 U16870 ( .A1(n13577), .A2(n13576), .ZN(n13578) );
  NAND2_X1 U16871 ( .A1(n13578), .A2(n13686), .ZN(n16246) );
  OAI211_X1 U16872 ( .C1(n13579), .C2(n13581), .A(n13580), .B(n14984), .ZN(
        n13583) );
  NAND2_X1 U16873 ( .A1(n14998), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13582) );
  OAI211_X1 U16874 ( .C1(n16246), .C2(n14998), .A(n13583), .B(n13582), .ZN(
        P2_U2879) );
  OR2_X1 U16875 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  AND2_X1 U16876 ( .A1(n13615), .A2(n13586), .ZN(n20107) );
  INV_X1 U16877 ( .A(n20107), .ZN(n14149) );
  NAND2_X1 U16878 ( .A1(n20165), .A2(DATAI_1_), .ZN(n13588) );
  NAND2_X1 U16879 ( .A1(n20164), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13587) );
  AND2_X1 U16880 ( .A1(n13588), .A2(n13587), .ZN(n20181) );
  OAI222_X1 U16881 ( .A1(n15896), .A2(n14149), .B1(n14551), .B2(n11261), .C1(
        n14549), .C2(n20181), .ZN(P1_U2903) );
  XNOR2_X1 U16882 ( .A(n13590), .B(n13589), .ZN(n13636) );
  NAND2_X1 U16883 ( .A1(n14702), .A2(n14701), .ZN(n13676) );
  INV_X1 U16884 ( .A(n13676), .ZN(n14266) );
  NAND2_X1 U16885 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13591) );
  OAI22_X1 U16886 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14266), .B1(
        n13591), .B2(n14757), .ZN(n13594) );
  OR2_X1 U16887 ( .A1(n14701), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13593) );
  OAI21_X1 U16888 ( .B1(n13594), .B2(n14700), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13605) );
  AOI21_X1 U16889 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U16890 ( .A1(n13596), .A2(n13595), .ZN(n13597) );
  AND2_X1 U16891 ( .A1(n13679), .A2(n13597), .ZN(n20085) );
  NAND2_X1 U16892 ( .A1(n16067), .A2(n20085), .ZN(n13602) );
  INV_X1 U16893 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21191) );
  NOR2_X1 U16894 ( .A1(n20055), .A2(n21191), .ZN(n13632) );
  INV_X1 U16895 ( .A(n13632), .ZN(n13601) );
  INV_X1 U16896 ( .A(n14702), .ZN(n13598) );
  NOR2_X1 U16897 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14760), .ZN(
        n13599) );
  NAND2_X1 U16898 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13599), .ZN(
        n13600) );
  NAND3_X1 U16899 ( .A1(n13602), .A2(n13601), .A3(n13600), .ZN(n13603) );
  AOI21_X1 U16900 ( .B1(n14692), .B2(n14250), .A(n13603), .ZN(n13604) );
  OAI211_X1 U16901 ( .C1(n13636), .C2(n16052), .A(n13605), .B(n13604), .ZN(
        P1_U3029) );
  INV_X1 U16902 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13606) );
  NOR2_X1 U16903 ( .A1(n13619), .A2(n13606), .ZN(n13608) );
  OAI211_X1 U16904 ( .C1(n13608), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14984), .B(n13424), .ZN(n13612) );
  OAI21_X1 U16905 ( .B1(n13622), .B2(n13610), .A(n13609), .ZN(n19067) );
  INV_X1 U16906 ( .A(n19067), .ZN(n15538) );
  NAND2_X1 U16907 ( .A1(n15538), .A2(n14962), .ZN(n13611) );
  OAI211_X1 U16908 ( .C1(n14962), .C2(n19062), .A(n13612), .B(n13611), .ZN(
        P2_U2881) );
  NAND2_X1 U16909 ( .A1(n13614), .A2(n13615), .ZN(n13616) );
  AND2_X1 U16910 ( .A1(n13613), .A2(n13616), .ZN(n20083) );
  INV_X1 U16911 ( .A(n20083), .ZN(n14151) );
  NAND2_X1 U16912 ( .A1(n20165), .A2(DATAI_2_), .ZN(n13618) );
  NAND2_X1 U16913 ( .A1(n20164), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13617) );
  AND2_X1 U16914 ( .A1(n13618), .A2(n13617), .ZN(n20187) );
  OAI222_X1 U16915 ( .A1(n15896), .A2(n14151), .B1(n14551), .B2(n11255), .C1(
        n14549), .C2(n20187), .ZN(P1_U2902) );
  XOR2_X1 U16916 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13619), .Z(n13625)
         );
  INV_X1 U16917 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13623) );
  NOR2_X1 U16918 ( .A1(n13504), .A2(n13620), .ZN(n13621) );
  OR2_X1 U16919 ( .A1(n13622), .A2(n13621), .ZN(n16259) );
  MUX2_X1 U16920 ( .A(n13623), .B(n16259), .S(n14962), .Z(n13624) );
  OAI21_X1 U16921 ( .B1(n13625), .B2(n15000), .A(n13624), .ZN(P2_U2882) );
  AOI22_X1 U16922 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20141), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15757), .ZN(n13626) );
  OAI21_X1 U16923 ( .B1(n11752), .B2(n13631), .A(n13626), .ZN(P1_U2906) );
  AOI22_X1 U16924 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13627) );
  OAI21_X1 U16925 ( .B1(n11553), .B2(n13631), .A(n13627), .ZN(P1_U2914) );
  AOI22_X1 U16926 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13628) );
  OAI21_X1 U16927 ( .B1(n21176), .B2(n13631), .A(n13628), .ZN(P1_U2915) );
  INV_X1 U16928 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n21192) );
  AOI22_X1 U16929 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13629) );
  OAI21_X1 U16930 ( .B1(n21192), .B2(n13631), .A(n13629), .ZN(P1_U2916) );
  AOI22_X1 U16931 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13630) );
  OAI21_X1 U16932 ( .B1(n11652), .B2(n13631), .A(n13630), .ZN(P1_U2910) );
  AOI21_X1 U16933 ( .B1(n15946), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13632), .ZN(n13633) );
  OAI21_X1 U16934 ( .B1(n20094), .B2(n15954), .A(n13633), .ZN(n13634) );
  AOI21_X1 U16935 ( .B1(n20083), .B2(n20166), .A(n13634), .ZN(n13635) );
  OAI21_X1 U16936 ( .B1(n13636), .B2(n15955), .A(n13635), .ZN(P1_U2997) );
  XNOR2_X1 U16937 ( .A(n13637), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13654) );
  INV_X1 U16938 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13638) );
  NOR2_X1 U16939 ( .A1(n20055), .A2(n13638), .ZN(n13651) );
  NOR2_X1 U16940 ( .A1(n15960), .A2(n13639), .ZN(n13640) );
  AOI211_X1 U16941 ( .C1(n13639), .C2(n15942), .A(n13651), .B(n13640), .ZN(
        n13642) );
  NAND2_X1 U16942 ( .A1(n20107), .A2(n20166), .ZN(n13641) );
  OAI211_X1 U16943 ( .C1(n13654), .C2(n15955), .A(n13642), .B(n13641), .ZN(
        P1_U2998) );
  NOR2_X1 U16944 ( .A1(n13643), .A2(n13101), .ZN(n13652) );
  OR2_X1 U16945 ( .A1(n13645), .A2(n13644), .ZN(n13646) );
  NAND2_X1 U16946 ( .A1(n13647), .A2(n13646), .ZN(n20095) );
  AND2_X1 U16947 ( .A1(n16067), .A2(n20095), .ZN(n13650) );
  AOI211_X1 U16948 ( .C1(n13648), .C2(n14702), .A(n14712), .B(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13649) );
  NOR4_X1 U16949 ( .A1(n13652), .A2(n13651), .A3(n13650), .A4(n13649), .ZN(
        n13653) );
  OAI21_X1 U16950 ( .B1(n13654), .B2(n16052), .A(n13653), .ZN(P1_U3030) );
  INV_X1 U16951 ( .A(n13656), .ZN(n13658) );
  NAND3_X1 U16952 ( .A1(n13658), .A2(n13657), .A3(n13613), .ZN(n13659) );
  NAND2_X1 U16953 ( .A1(n13655), .A2(n13659), .ZN(n14073) );
  NAND2_X1 U16954 ( .A1(n20165), .A2(DATAI_3_), .ZN(n13661) );
  NAND2_X1 U16955 ( .A1(n20164), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13660) );
  AND2_X1 U16956 ( .A1(n13661), .A2(n13660), .ZN(n20194) );
  OAI222_X1 U16957 ( .A1(n15896), .A2(n14073), .B1(n14551), .B2(n11282), .C1(
        n14549), .C2(n20194), .ZN(P1_U2901) );
  XNOR2_X1 U16958 ( .A(n19961), .B(n19962), .ZN(n13666) );
  INV_X1 U16959 ( .A(n19976), .ZN(n14886) );
  NAND2_X1 U16960 ( .A1(n19971), .A2(n14886), .ZN(n13663) );
  OAI21_X1 U16961 ( .B1(n19971), .B2(n14886), .A(n13663), .ZN(n19173) );
  NOR2_X1 U16962 ( .A1(n19981), .A2(n13662), .ZN(n19180) );
  NOR2_X1 U16963 ( .A1(n19173), .A2(n19180), .ZN(n19172) );
  INV_X1 U16964 ( .A(n13663), .ZN(n13664) );
  NOR2_X1 U16965 ( .A1(n19172), .A2(n13664), .ZN(n13665) );
  NOR2_X1 U16966 ( .A1(n13665), .A2(n13666), .ZN(n19151) );
  AOI21_X1 U16967 ( .B1(n13666), .B2(n13665), .A(n19151), .ZN(n13673) );
  AOI22_X1 U16968 ( .A1(n19179), .A2(n13667), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19178), .ZN(n13672) );
  NOR2_X1 U16969 ( .A1(n13669), .A2(n13668), .ZN(n13670) );
  NAND2_X1 U16970 ( .A1(n19149), .A2(n16164), .ZN(n13671) );
  OAI211_X1 U16971 ( .C1(n13673), .C2(n19174), .A(n13672), .B(n13671), .ZN(
        P2_U2917) );
  XNOR2_X1 U16972 ( .A(n13675), .B(n13674), .ZN(n13734) );
  AOI21_X1 U16973 ( .B1(n14692), .B2(n14250), .A(n14700), .ZN(n13889) );
  NAND2_X1 U16974 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13677) );
  NAND2_X1 U16975 ( .A1(n13676), .A2(n13677), .ZN(n13890) );
  NAND2_X1 U16976 ( .A1(n13889), .A2(n13890), .ZN(n16040) );
  NOR2_X1 U16977 ( .A1(n14760), .A2(n13677), .ZN(n13949) );
  NOR2_X1 U16978 ( .A1(n14692), .A2(n13949), .ZN(n14248) );
  AOI22_X1 U16979 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16040), .B1(
        n13943), .B2(n11790), .ZN(n13683) );
  AND2_X1 U16980 ( .A1(n13679), .A2(n13678), .ZN(n13680) );
  OR2_X1 U16981 ( .A1(n13772), .A2(n13680), .ZN(n14069) );
  INV_X1 U16982 ( .A(n14069), .ZN(n13681) );
  INV_X1 U16983 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20912) );
  NOR2_X1 U16984 ( .A1(n20055), .A2(n20912), .ZN(n13729) );
  AOI21_X1 U16985 ( .B1(n16067), .B2(n13681), .A(n13729), .ZN(n13682) );
  OAI211_X1 U16986 ( .C1(n16052), .C2(n13734), .A(n13683), .B(n13682), .ZN(
        P1_U3028) );
  OAI211_X1 U16987 ( .C1(n11975), .C2(n11974), .A(n14984), .B(n13685), .ZN(
        n13689) );
  AOI21_X1 U16988 ( .B1(n13687), .B2(n13686), .A(n13780), .ZN(n19057) );
  NAND2_X1 U16989 ( .A1(n19057), .A2(n14962), .ZN(n13688) );
  OAI211_X1 U16990 ( .C1(n14962), .C2(n10887), .A(n13689), .B(n13688), .ZN(
        P2_U2878) );
  AOI22_X1 U16991 ( .A1(n20153), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20152), .ZN(n13694) );
  NAND2_X1 U16992 ( .A1(n20165), .A2(DATAI_5_), .ZN(n13693) );
  NAND2_X1 U16993 ( .A1(n20164), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13692) );
  AND2_X1 U16994 ( .A1(n13693), .A2(n13692), .ZN(n20207) );
  INV_X1 U16995 ( .A(n20207), .ZN(n15881) );
  NAND2_X1 U16996 ( .A1(n13725), .A2(n15881), .ZN(n13697) );
  NAND2_X1 U16997 ( .A1(n13694), .A2(n13697), .ZN(P1_U2957) );
  AOI22_X1 U16998 ( .A1(n20153), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20152), .ZN(n13695) );
  INV_X1 U16999 ( .A(n20187), .ZN(n14539) );
  NAND2_X1 U17000 ( .A1(n13725), .A2(n14539), .ZN(n13703) );
  NAND2_X1 U17001 ( .A1(n13695), .A2(n13703), .ZN(P1_U2954) );
  AOI22_X1 U17002 ( .A1(n20153), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20152), .ZN(n13696) );
  INV_X1 U17003 ( .A(n20194), .ZN(n15886) );
  NAND2_X1 U17004 ( .A1(n13725), .A2(n15886), .ZN(n13713) );
  NAND2_X1 U17005 ( .A1(n13696), .A2(n13713), .ZN(P1_U2955) );
  AOI22_X1 U17006 ( .A1(n20153), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20152), .ZN(n13698) );
  NAND2_X1 U17007 ( .A1(n13698), .A2(n13697), .ZN(P1_U2942) );
  AOI22_X1 U17008 ( .A1(n20153), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20152), .ZN(n13699) );
  INV_X1 U17009 ( .A(n20181), .ZN(n15892) );
  NAND2_X1 U17010 ( .A1(n13725), .A2(n15892), .ZN(n13705) );
  NAND2_X1 U17011 ( .A1(n13699), .A2(n13705), .ZN(P1_U2953) );
  AOI22_X1 U17012 ( .A1(n20153), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20152), .ZN(n13702) );
  NAND2_X1 U17013 ( .A1(n20165), .A2(DATAI_6_), .ZN(n13701) );
  NAND2_X1 U17014 ( .A1(n20164), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13700) );
  AND2_X1 U17015 ( .A1(n13701), .A2(n13700), .ZN(n20213) );
  INV_X1 U17016 ( .A(n20213), .ZN(n14533) );
  NAND2_X1 U17017 ( .A1(n13725), .A2(n14533), .ZN(n13707) );
  NAND2_X1 U17018 ( .A1(n13702), .A2(n13707), .ZN(P1_U2958) );
  AOI22_X1 U17019 ( .A1(n20153), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20152), .ZN(n13704) );
  NAND2_X1 U17020 ( .A1(n13704), .A2(n13703), .ZN(P1_U2939) );
  AOI22_X1 U17021 ( .A1(n20153), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20152), .ZN(n13706) );
  NAND2_X1 U17022 ( .A1(n13706), .A2(n13705), .ZN(P1_U2938) );
  AOI22_X1 U17023 ( .A1(n20153), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20152), .ZN(n13708) );
  NAND2_X1 U17024 ( .A1(n13708), .A2(n13707), .ZN(P1_U2943) );
  AOI22_X1 U17025 ( .A1(n20153), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20152), .ZN(n13711) );
  NAND2_X1 U17026 ( .A1(n20165), .A2(DATAI_4_), .ZN(n13710) );
  NAND2_X1 U17027 ( .A1(n20164), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13709) );
  AND2_X1 U17028 ( .A1(n13710), .A2(n13709), .ZN(n20200) );
  INV_X1 U17029 ( .A(n20200), .ZN(n14536) );
  NAND2_X1 U17030 ( .A1(n13725), .A2(n14536), .ZN(n13716) );
  NAND2_X1 U17031 ( .A1(n13711), .A2(n13716), .ZN(P1_U2941) );
  AOI22_X1 U17032 ( .A1(n20153), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20152), .ZN(n13712) );
  INV_X1 U17033 ( .A(n20163), .ZN(n14542) );
  NAND2_X1 U17034 ( .A1(n13725), .A2(n14542), .ZN(n13718) );
  NAND2_X1 U17035 ( .A1(n13712), .A2(n13718), .ZN(P1_U2937) );
  AOI22_X1 U17036 ( .A1(n20153), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20152), .ZN(n13714) );
  NAND2_X1 U17037 ( .A1(n13714), .A2(n13713), .ZN(P1_U2940) );
  AOI22_X1 U17038 ( .A1(n20153), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20152), .ZN(n13715) );
  MUX2_X1 U17039 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20164), .Z(
        n14516) );
  NAND2_X1 U17040 ( .A1(n13725), .A2(n14516), .ZN(n13720) );
  NAND2_X1 U17041 ( .A1(n13715), .A2(n13720), .ZN(P1_U2948) );
  AOI22_X1 U17042 ( .A1(n20153), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20152), .ZN(n13717) );
  NAND2_X1 U17043 ( .A1(n13717), .A2(n13716), .ZN(P1_U2956) );
  AOI22_X1 U17044 ( .A1(n20153), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20152), .ZN(n13719) );
  NAND2_X1 U17045 ( .A1(n13719), .A2(n13718), .ZN(P1_U2952) );
  AOI22_X1 U17046 ( .A1(n20153), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20152), .ZN(n13721) );
  NAND2_X1 U17047 ( .A1(n13721), .A2(n13720), .ZN(P1_U2963) );
  AOI22_X1 U17048 ( .A1(n20153), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20152), .ZN(n13722) );
  MUX2_X1 U17049 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20164), .Z(
        n14522) );
  NAND2_X1 U17050 ( .A1(n13725), .A2(n14522), .ZN(n20144) );
  NAND2_X1 U17051 ( .A1(n13722), .A2(n20144), .ZN(P1_U2946) );
  AOI22_X1 U17052 ( .A1(n20153), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20152), .ZN(n13726) );
  NAND2_X1 U17053 ( .A1(n20165), .A2(DATAI_7_), .ZN(n13724) );
  NAND2_X1 U17054 ( .A1(n20164), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13723) );
  AND2_X1 U17055 ( .A1(n13724), .A2(n13723), .ZN(n20219) );
  INV_X1 U17056 ( .A(n20219), .ZN(n14529) );
  NAND2_X1 U17057 ( .A1(n13725), .A2(n14529), .ZN(n13727) );
  NAND2_X1 U17058 ( .A1(n13726), .A2(n13727), .ZN(P1_U2959) );
  AOI22_X1 U17059 ( .A1(n20153), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20152), .ZN(n13728) );
  NAND2_X1 U17060 ( .A1(n13728), .A2(n13727), .ZN(P1_U2944) );
  INV_X1 U17061 ( .A(n14073), .ZN(n13732) );
  AOI21_X1 U17062 ( .B1(n15946), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13729), .ZN(n13730) );
  OAI21_X1 U17063 ( .B1(n14063), .B2(n15954), .A(n13730), .ZN(n13731) );
  AOI21_X1 U17064 ( .B1(n13732), .B2(n20166), .A(n13731), .ZN(n13733) );
  OAI21_X1 U17065 ( .B1(n13734), .B2(n15955), .A(n13733), .ZN(P1_U2996) );
  INV_X1 U17066 ( .A(n20436), .ZN(n14067) );
  AND2_X1 U17067 ( .A1(n13751), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13736) );
  INV_X1 U17068 ( .A(n13736), .ZN(n13735) );
  MUX2_X1 U17069 ( .A(n13736), .B(n13735), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13743) );
  INV_X1 U17070 ( .A(n13393), .ZN(n13738) );
  NAND2_X1 U17071 ( .A1(n13738), .A2(n13737), .ZN(n13740) );
  OAI21_X1 U17072 ( .B1(n13393), .B2(n13751), .A(n11865), .ZN(n13739) );
  NAND2_X1 U17073 ( .A1(n13740), .A2(n13739), .ZN(n13741) );
  AOI22_X1 U17074 ( .A1(n15675), .A2(n13743), .B1(n13742), .B2(n13741), .ZN(
        n13749) );
  NAND2_X1 U17075 ( .A1(n13393), .A2(n13751), .ZN(n13744) );
  NAND2_X1 U17076 ( .A1(n13744), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13745) );
  NAND2_X1 U17077 ( .A1(n11179), .A2(n13745), .ZN(n20797) );
  NAND3_X1 U17078 ( .A1(n13747), .A2(n13746), .A3(n20797), .ZN(n13748) );
  OAI211_X1 U17079 ( .C1(n14067), .C2(n14807), .A(n13749), .B(n13748), .ZN(
        n20799) );
  MUX2_X1 U17080 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20799), .S(
        n15680), .Z(n15689) );
  NOR2_X1 U17081 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16083), .ZN(n13752) );
  AOI22_X1 U17082 ( .A1(n15689), .A2(n16083), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13752), .ZN(n13754) );
  MUX2_X1 U17083 ( .A(n13751), .B(n13750), .S(n15680), .Z(n15687) );
  AOI22_X1 U17084 ( .A1(n13752), .A2(n13751), .B1(n16083), .B2(n15687), .ZN(
        n13753) );
  NOR2_X1 U17085 ( .A1(n13754), .A2(n13753), .ZN(n15717) );
  INV_X1 U17086 ( .A(n15717), .ZN(n13759) );
  INV_X1 U17087 ( .A(n20328), .ZN(n20570) );
  NOR2_X1 U17088 ( .A1(n13755), .A2(n20570), .ZN(n13756) );
  XOR2_X1 U17089 ( .A(n16077), .B(n13756), .Z(n20068) );
  NOR2_X1 U17090 ( .A1(n20068), .A2(n13366), .ZN(n16075) );
  NAND2_X1 U17091 ( .A1(n15680), .A2(n16083), .ZN(n13758) );
  OAI21_X1 U17092 ( .B1(n16077), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13758), .ZN(
        n13757) );
  OAI21_X1 U17093 ( .B1(n16075), .B2(n13758), .A(n13757), .ZN(n15715) );
  OAI21_X1 U17094 ( .B1(n13759), .B2(n10920), .A(n15715), .ZN(n13777) );
  OAI21_X1 U17095 ( .B1(n13777), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13760), .ZN(
        n13762) );
  NOR2_X1 U17096 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20825) );
  AND2_X1 U17097 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20579), .ZN(n14803) );
  OR2_X1 U17098 ( .A1(n13763), .A2(n20540), .ZN(n13764) );
  NAND2_X1 U17099 ( .A1(n20688), .A2(n21140), .ZN(n20568) );
  AND2_X1 U17100 ( .A1(n13764), .A2(n20568), .ZN(n20298) );
  NAND3_X1 U17101 ( .A1(n13763), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n20688), 
        .ZN(n13765) );
  MUX2_X1 U17102 ( .A(n20298), .B(n13765), .S(n11774), .Z(n13766) );
  OAI21_X1 U17103 ( .B1(n14803), .B2(n13382), .A(n13766), .ZN(n13767) );
  NAND2_X1 U17104 ( .A1(n20156), .A2(n13767), .ZN(n13768) );
  OAI21_X1 U17105 ( .B1(n20156), .B2(n20573), .A(n13768), .ZN(P1_U3476) );
  XNOR2_X1 U17106 ( .A(n13770), .B(n13769), .ZN(n13907) );
  NAND2_X1 U17107 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13893) );
  OAI211_X1 U17108 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13943), .B(n13893), .ZN(n13776) );
  OR2_X1 U17109 ( .A1(n13772), .A2(n13771), .ZN(n13773) );
  NAND2_X1 U17110 ( .A1(n13895), .A2(n13773), .ZN(n20072) );
  INV_X1 U17111 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20962) );
  OAI22_X1 U17112 ( .A1(n16046), .A2(n20072), .B1(n20962), .B2(n20055), .ZN(
        n13774) );
  AOI21_X1 U17113 ( .B1(n16040), .B2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13774), .ZN(n13775) );
  OAI211_X1 U17114 ( .C1(n16052), .C2(n13907), .A(n13776), .B(n13775), .ZN(
        P1_U3027) );
  NOR2_X1 U17115 ( .A1(n13777), .A2(n16084), .ZN(n15727) );
  OAI22_X1 U17116 ( .A1(n20257), .A2(n20540), .B1(n14008), .B2(n14803), .ZN(
        n13778) );
  OAI21_X1 U17117 ( .B1(n15727), .B2(n13778), .A(n20156), .ZN(n13779) );
  OAI21_X1 U17118 ( .B1(n20156), .B2(n20610), .A(n13779), .ZN(P1_U3478) );
  OR2_X1 U17119 ( .A1(n13781), .A2(n13780), .ZN(n13782) );
  NAND2_X1 U17120 ( .A1(n13782), .A2(n13911), .ZN(n19043) );
  INV_X2 U17121 ( .A(n14962), .ZN(n14980) );
  INV_X1 U17122 ( .A(n13685), .ZN(n13785) );
  INV_X1 U17123 ( .A(n13783), .ZN(n13784) );
  OAI211_X1 U17124 ( .C1(n13785), .C2(n9834), .A(n13784), .B(n14984), .ZN(
        n13787) );
  NAND2_X1 U17125 ( .A1(n14998), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13786) );
  OAI211_X1 U17126 ( .C1(n19043), .C2(n14980), .A(n13787), .B(n13786), .ZN(
        P2_U2877) );
  INV_X1 U17127 ( .A(n11774), .ZN(n13789) );
  MUX2_X1 U17128 ( .A(n20638), .B(n20409), .S(n13763), .Z(n13792) );
  NOR3_X1 U17129 ( .A1(n20490), .A2(n13792), .A3(n21140), .ZN(n13793) );
  AOI211_X1 U17130 ( .C1(n21140), .C2(n13788), .A(n20540), .B(n13793), .ZN(
        n13795) );
  NOR2_X1 U17131 ( .A1(n14067), .A2(n14803), .ZN(n13794) );
  OAI21_X1 U17132 ( .B1(n13795), .B2(n13794), .A(n20156), .ZN(n13796) );
  OAI21_X1 U17133 ( .B1(n15688), .B2(n20156), .A(n13796), .ZN(P1_U3475) );
  AND2_X1 U17134 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16981) );
  NAND3_X1 U17135 ( .A1(n17402), .A2(n13798), .A3(n13797), .ZN(n13801) );
  INV_X1 U17136 ( .A(n18666), .ZN(n13800) );
  NAND2_X1 U17137 ( .A1(n13800), .A2(n13799), .ZN(n15643) );
  NOR2_X1 U17138 ( .A1(n18272), .A2(n17257), .ZN(n17274) );
  INV_X1 U17139 ( .A(n17274), .ZN(n17272) );
  NOR2_X2 U17140 ( .A1(n17257), .A2(n17402), .ZN(n17275) );
  INV_X1 U17141 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16942) );
  INV_X1 U17142 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16940) );
  INV_X1 U17143 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17003) );
  INV_X1 U17144 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16683) );
  INV_X1 U17145 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17085) );
  AND3_X1 U17146 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n14281) );
  NAND4_X1 U17147 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(P3_EBX_REG_2__SCAN_IN), .ZN(n17256) );
  NAND4_X1 U17148 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_11__SCAN_IN), .A4(P3_EBX_REG_10__SCAN_IN), .ZN(n15628)
         );
  NAND4_X1 U17149 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(P3_EBX_REG_4__SCAN_IN), .ZN(n13803) );
  NOR3_X1 U17150 ( .A1(n17256), .A2(n15628), .A3(n13803), .ZN(n13804) );
  NAND4_X1 U17151 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(n14281), .A4(n13804), .ZN(n17103) );
  NOR3_X1 U17152 ( .A1(n17085), .A2(n17257), .A3(n17103), .ZN(n17089) );
  AND2_X1 U17153 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17089), .ZN(n17059) );
  NAND2_X1 U17154 ( .A1(n17402), .A2(n17074), .ZN(n17055) );
  NOR2_X1 U17155 ( .A1(n16683), .A2(n17055), .ZN(n17040) );
  NAND2_X1 U17156 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17040), .ZN(n17009) );
  NOR3_X1 U17157 ( .A1(n16940), .A2(n17003), .A3(n17009), .ZN(n17008) );
  NAND2_X1 U17158 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17008), .ZN(n16993) );
  NAND2_X1 U17159 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16997), .ZN(n16991) );
  NAND2_X1 U17160 ( .A1(n17266), .A2(n16991), .ZN(n13805) );
  OAI21_X1 U17161 ( .B1(n16981), .B2(n17272), .A(n13805), .ZN(n16979) );
  OAI22_X1 U17162 ( .A1(n10240), .A2(n13807), .B1(n17191), .B2(n13806), .ZN(
        n13818) );
  AOI22_X1 U17163 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U17164 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17195), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13815) );
  AOI22_X1 U17165 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13808) );
  OAI21_X1 U17166 ( .B1(n12780), .B2(n17031), .A(n13808), .ZN(n13813) );
  AOI22_X1 U17167 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17223), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U17168 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13809) );
  OAI211_X1 U17169 ( .C1(n17216), .C2(n13811), .A(n13810), .B(n13809), .ZN(
        n13812) );
  AOI211_X1 U17170 ( .C1(n17206), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n13813), .B(n13812), .ZN(n13814) );
  NAND3_X1 U17171 ( .A1(n13816), .A2(n13815), .A3(n13814), .ZN(n13817) );
  AOI211_X1 U17172 ( .C1(n17043), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n13818), .B(n13817), .ZN(n13882) );
  AOI22_X1 U17173 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13819) );
  OAI21_X1 U17174 ( .B1(n10239), .B2(n17157), .A(n13819), .ZN(n13829) );
  INV_X1 U17175 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U17176 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13827) );
  AOI22_X1 U17177 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13820) );
  OAI21_X1 U17178 ( .B1(n10240), .B2(n17061), .A(n13820), .ZN(n13825) );
  INV_X1 U17179 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13823) );
  AOI22_X1 U17180 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13822) );
  AOI22_X1 U17181 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13821) );
  OAI211_X1 U17182 ( .C1(n17216), .C2(n13823), .A(n13822), .B(n13821), .ZN(
        n13824) );
  AOI211_X1 U17183 ( .C1(n17206), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n13825), .B(n13824), .ZN(n13826) );
  OAI211_X1 U17184 ( .C1(n17193), .C2(n17066), .A(n13827), .B(n13826), .ZN(
        n13828) );
  AOI211_X1 U17185 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n13829), .B(n13828), .ZN(n16989) );
  INV_X1 U17186 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U17187 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13830) );
  OAI21_X1 U17188 ( .B1(n13841), .B2(n17093), .A(n13830), .ZN(n13839) );
  AOI22_X1 U17189 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13837) );
  INV_X1 U17190 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17198) );
  OAI22_X1 U17191 ( .A1(n17218), .A2(n17190), .B1(n17191), .B2(n17198), .ZN(
        n13835) );
  AOI22_X1 U17192 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U17193 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U17194 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13831) );
  NAND3_X1 U17195 ( .A1(n13833), .A2(n13832), .A3(n13831), .ZN(n13834) );
  AOI211_X1 U17196 ( .C1(n17220), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n13835), .B(n13834), .ZN(n13836) );
  OAI211_X1 U17197 ( .C1(n10240), .C2(n17092), .A(n13837), .B(n13836), .ZN(
        n13838) );
  AOI211_X1 U17198 ( .C1(n9803), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n13839), .B(n13838), .ZN(n16999) );
  INV_X1 U17199 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U17200 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13850) );
  AOI22_X1 U17201 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13840) );
  OAI21_X1 U17202 ( .B1(n12737), .B2(n17226), .A(n13840), .ZN(n13848) );
  OAI22_X1 U17203 ( .A1(n17193), .A2(n17217), .B1(n13841), .B2(n17232), .ZN(
        n13842) );
  AOI21_X1 U17204 ( .B1(n17194), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n13842), .ZN(n13846) );
  AOI22_X1 U17205 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U17206 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17207 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13843) );
  NAND4_X1 U17208 ( .A1(n13846), .A2(n13845), .A3(n13844), .A4(n13843), .ZN(
        n13847) );
  AOI211_X1 U17209 ( .C1(n12723), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n13848), .B(n13847), .ZN(n13849) );
  OAI211_X1 U17210 ( .C1(n10240), .C2(n17109), .A(n13850), .B(n13849), .ZN(
        n17005) );
  AOI22_X1 U17211 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17229), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17043), .ZN(n13860) );
  AOI22_X1 U17212 ( .A1(n9799), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17219), .ZN(n13852) );
  AOI22_X1 U17213 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17214), .ZN(n13851) );
  OAI211_X1 U17214 ( .C1(n17133), .C2(n17216), .A(n13852), .B(n13851), .ZN(
        n13858) );
  AOI22_X1 U17215 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n9803), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13856) );
  AOI22_X1 U17216 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U17217 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17200), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17194), .ZN(n13854) );
  NAND2_X1 U17218 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n13853) );
  NAND4_X1 U17219 ( .A1(n13856), .A2(n13855), .A3(n13854), .A4(n13853), .ZN(
        n13857) );
  AOI211_X1 U17220 ( .C1(n17206), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n13858), .B(n13857), .ZN(n13859) );
  OAI211_X1 U17221 ( .C1(n17193), .C2(n17247), .A(n13860), .B(n13859), .ZN(
        n17006) );
  NAND2_X1 U17222 ( .A1(n17005), .A2(n17006), .ZN(n17004) );
  NOR2_X1 U17223 ( .A1(n16999), .A2(n17004), .ZN(n16998) );
  AOI22_X1 U17224 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13870) );
  AOI22_X1 U17225 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13862) );
  AOI22_X1 U17226 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13861) );
  OAI211_X1 U17227 ( .C1(n17227), .C2(n17174), .A(n13862), .B(n13861), .ZN(
        n13868) );
  AOI22_X1 U17228 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13866) );
  AOI22_X1 U17229 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13865) );
  AOI22_X1 U17230 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13864) );
  NAND2_X1 U17231 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13863) );
  NAND4_X1 U17232 ( .A1(n13866), .A2(n13865), .A3(n13864), .A4(n13863), .ZN(
        n13867) );
  AOI211_X1 U17233 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n13868), .B(n13867), .ZN(n13869) );
  OAI211_X1 U17234 ( .C1(n10240), .C2(n13871), .A(n13870), .B(n13869), .ZN(
        n16995) );
  NAND2_X1 U17235 ( .A1(n16998), .A2(n16995), .ZN(n16994) );
  NOR2_X1 U17236 ( .A1(n16989), .A2(n16994), .ZN(n16988) );
  AOI22_X1 U17237 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13881) );
  AOI22_X1 U17238 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13873) );
  AOI22_X1 U17239 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13872) );
  OAI211_X1 U17240 ( .C1(n17227), .C2(n17140), .A(n13873), .B(n13872), .ZN(
        n13879) );
  AOI22_X1 U17241 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13877) );
  AOI22_X1 U17242 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U17243 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13875) );
  NAND2_X1 U17244 ( .A1(n15618), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13874) );
  NAND4_X1 U17245 ( .A1(n13877), .A2(n13876), .A3(n13875), .A4(n13874), .ZN(
        n13878) );
  AOI211_X1 U17246 ( .C1(n17206), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n13879), .B(n13878), .ZN(n13880) );
  OAI211_X1 U17247 ( .C1(n17216), .C2(n17149), .A(n13881), .B(n13880), .ZN(
        n16985) );
  NAND2_X1 U17248 ( .A1(n16988), .A2(n16985), .ZN(n16984) );
  NOR2_X1 U17249 ( .A1(n13882), .A2(n16984), .ZN(n16978) );
  AOI21_X1 U17250 ( .B1(n13882), .B2(n16984), .A(n16978), .ZN(n17295) );
  AOI22_X1 U17251 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16979), .B1(n17295), 
        .B2(n17275), .ZN(n13886) );
  INV_X1 U17252 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n13884) );
  INV_X1 U17253 ( .A(n16991), .ZN(n13883) );
  NAND3_X1 U17254 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n13884), .A3(n13883), 
        .ZN(n13885) );
  NAND2_X1 U17255 ( .A1(n13886), .A2(n13885), .ZN(P3_U2675) );
  XNOR2_X1 U17256 ( .A(n13888), .B(n13887), .ZN(n13922) );
  INV_X1 U17257 ( .A(n13893), .ZN(n13892) );
  NAND2_X1 U17258 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13892), .ZN(
        n14249) );
  INV_X1 U17259 ( .A(n14249), .ZN(n14253) );
  OAI21_X1 U17260 ( .B1(n14253), .B2(n14757), .A(n13889), .ZN(n14268) );
  INV_X1 U17261 ( .A(n14268), .ZN(n13891) );
  OAI211_X1 U17262 ( .C1(n14266), .C2(n13892), .A(n13891), .B(n13890), .ZN(
        n13947) );
  NOR2_X1 U17263 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13893), .ZN(
        n13948) );
  AOI22_X1 U17264 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13947), .B1(
        n13943), .B2(n13948), .ZN(n13898) );
  NAND2_X1 U17265 ( .A1(n13895), .A2(n13894), .ZN(n13896) );
  AND2_X1 U17266 ( .A1(n13945), .A2(n13896), .ZN(n20054) );
  INV_X1 U17267 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20984) );
  NOR2_X1 U17268 ( .A1(n20055), .A2(n20984), .ZN(n13918) );
  AOI21_X1 U17269 ( .B1(n16067), .B2(n20054), .A(n13918), .ZN(n13897) );
  OAI211_X1 U17270 ( .C1(n16052), .C2(n13922), .A(n13898), .B(n13897), .ZN(
        P1_U3026) );
  INV_X1 U17271 ( .A(n13900), .ZN(n13901) );
  AOI21_X1 U17272 ( .B1(n13902), .B2(n13655), .A(n13901), .ZN(n20077) );
  NAND2_X1 U17273 ( .A1(n20077), .A2(n20166), .ZN(n13906) );
  OAI22_X1 U17274 ( .A1(n15960), .A2(n13903), .B1(n20055), .B2(n20962), .ZN(
        n13904) );
  AOI21_X1 U17275 ( .B1(n15942), .B2(n20076), .A(n13904), .ZN(n13905) );
  OAI211_X1 U17276 ( .C1(n13907), .C2(n15955), .A(n13906), .B(n13905), .ZN(
        P1_U2995) );
  INV_X1 U17277 ( .A(n20077), .ZN(n13971) );
  INV_X1 U17278 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20137) );
  OAI222_X1 U17279 ( .A1(n15896), .A2(n13971), .B1(n14551), .B2(n20137), .C1(
        n14549), .C2(n20200), .ZN(P1_U2900) );
  INV_X1 U17280 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19025) );
  INV_X1 U17281 ( .A(n13908), .ZN(n13909) );
  OAI211_X1 U17282 ( .C1(n13783), .C2(n13910), .A(n13908), .B(n14984), .ZN(
        n13914) );
  AOI21_X1 U17283 ( .B1(n13912), .B2(n13911), .A(n13923), .ZN(n19032) );
  NAND2_X1 U17284 ( .A1(n19032), .A2(n14962), .ZN(n13913) );
  OAI211_X1 U17285 ( .C1(n14962), .C2(n19025), .A(n13914), .B(n13913), .ZN(
        P2_U2876) );
  AND2_X1 U17286 ( .A1(n13900), .A2(n13916), .ZN(n13917) );
  NOR2_X1 U17287 ( .A1(n13915), .A2(n13917), .ZN(n20061) );
  AOI21_X1 U17288 ( .B1(n15946), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13918), .ZN(n13919) );
  OAI21_X1 U17289 ( .B1(n20066), .B2(n15954), .A(n13919), .ZN(n13920) );
  AOI21_X1 U17290 ( .B1(n20061), .B2(n20166), .A(n13920), .ZN(n13921) );
  OAI21_X1 U17291 ( .B1(n13922), .B2(n15955), .A(n13921), .ZN(P1_U2994) );
  OR2_X1 U17292 ( .A1(n13924), .A2(n13923), .ZN(n13925) );
  AND2_X1 U17293 ( .A1(n13925), .A2(n14053), .ZN(n16215) );
  INV_X1 U17294 ( .A(n14120), .ZN(n14056) );
  OAI211_X1 U17295 ( .C1(n13909), .C2(n13926), .A(n14056), .B(n14984), .ZN(
        n13928) );
  NAND2_X1 U17296 ( .A1(n14998), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13927) );
  OAI211_X1 U17297 ( .C1(n15428), .C2(n14998), .A(n13928), .B(n13927), .ZN(
        P2_U2875) );
  INV_X1 U17298 ( .A(n20061), .ZN(n14153) );
  OAI222_X1 U17299 ( .A1(n15896), .A2(n14153), .B1(n14551), .B2(n11300), .C1(
        n14549), .C2(n20207), .ZN(P1_U2899) );
  NOR2_X1 U17300 ( .A1(n19092), .A2(n13930), .ZN(n13931) );
  XNOR2_X1 U17301 ( .A(n13931), .B(n16250), .ZN(n13932) );
  INV_X1 U17302 ( .A(n19048), .ZN(n14868) );
  NAND2_X1 U17303 ( .A1(n13932), .A2(n14868), .ZN(n13939) );
  AOI21_X1 U17304 ( .B1(n13934), .B2(n13933), .A(n15489), .ZN(n15509) );
  INV_X1 U17305 ( .A(n15509), .ZN(n19144) );
  AOI22_X1 U17306 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19114), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19107), .ZN(n13935) );
  OAI211_X1 U17307 ( .C1(n19085), .C2(n19144), .A(n13935), .B(n19041), .ZN(
        n13937) );
  NOR2_X1 U17308 ( .A1(n19109), .A2(n16246), .ZN(n13936) );
  AOI211_X1 U17309 ( .C1(n19102), .C2(P2_REIP_REG_8__SCAN_IN), .A(n13937), .B(
        n13936), .ZN(n13938) );
  OAI211_X1 U17310 ( .C1(n19105), .C2(n13940), .A(n13939), .B(n13938), .ZN(
        P2_U2847) );
  XNOR2_X1 U17311 ( .A(n13942), .B(n13941), .ZN(n15956) );
  NAND2_X1 U17312 ( .A1(n14253), .A2(n13943), .ZN(n16048) );
  INV_X1 U17313 ( .A(n16048), .ZN(n13952) );
  NAND2_X1 U17314 ( .A1(n13945), .A2(n13944), .ZN(n13946) );
  NAND2_X1 U17315 ( .A1(n16064), .A2(n13946), .ZN(n20041) );
  NAND2_X1 U17316 ( .A1(n20070), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n15958) );
  OAI21_X1 U17317 ( .B1(n16046), .B2(n20041), .A(n15958), .ZN(n13951) );
  AOI21_X1 U17318 ( .B1(n13949), .B2(n13948), .A(n13947), .ZN(n14138) );
  NOR2_X1 U17319 ( .A1(n14138), .A2(n11824), .ZN(n13950) );
  AOI211_X1 U17320 ( .C1(n11824), .C2(n13952), .A(n13951), .B(n13950), .ZN(
        n13953) );
  OAI21_X1 U17321 ( .B1(n16052), .B2(n15956), .A(n13953), .ZN(P1_U3025) );
  NOR2_X1 U17322 ( .A1(n13915), .A2(n13956), .ZN(n13957) );
  OR2_X1 U17323 ( .A1(n13955), .A2(n13957), .ZN(n20044) );
  OAI222_X1 U17324 ( .A1(n15896), .A2(n20044), .B1(n14551), .B2(n11311), .C1(
        n14549), .C2(n20213), .ZN(P1_U2898) );
  NAND2_X1 U17325 ( .A1(n13929), .A2(n13958), .ZN(n13959) );
  XNOR2_X1 U17326 ( .A(n16253), .B(n13959), .ZN(n13968) );
  XNOR2_X1 U17327 ( .A(n13961), .B(n13960), .ZN(n19145) );
  INV_X1 U17328 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19889) );
  AOI22_X1 U17329 ( .A1(n19039), .A2(n13962), .B1(n19107), .B2(
        P2_EBX_REG_7__SCAN_IN), .ZN(n13963) );
  OAI211_X1 U17330 ( .C1(n19889), .C2(n19049), .A(n13963), .B(n19041), .ZN(
        n13964) );
  AOI21_X1 U17331 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19114), .A(
        n13964), .ZN(n13966) );
  INV_X1 U17332 ( .A(n15529), .ZN(n16254) );
  NAND2_X1 U17333 ( .A1(n19081), .A2(n16254), .ZN(n13965) );
  OAI211_X1 U17334 ( .C1(n19145), .C2(n19085), .A(n13966), .B(n13965), .ZN(
        n13967) );
  AOI21_X1 U17335 ( .B1(n13968), .B2(n14868), .A(n13967), .ZN(n13969) );
  INV_X1 U17336 ( .A(n13969), .ZN(P2_U2848) );
  INV_X1 U17337 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13970) );
  OAI222_X1 U17338 ( .A1(n13971), .A2(n14503), .B1(n14492), .B2(n13970), .C1(
        n20072), .C2(n15876), .ZN(P1_U2868) );
  INV_X1 U17339 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13972) );
  OAI222_X1 U17340 ( .A1(n14073), .A2(n14503), .B1(n13972), .B2(n14492), .C1(
        n14069), .C2(n15876), .ZN(P1_U2869) );
  NAND2_X1 U17341 ( .A1(n13929), .A2(n13973), .ZN(n13974) );
  XNOR2_X1 U17342 ( .A(n16267), .B(n13974), .ZN(n13986) );
  INV_X1 U17343 ( .A(n19112), .ZN(n19089) );
  INV_X1 U17344 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19882) );
  OAI22_X1 U17345 ( .A1(n19105), .A2(n13975), .B1(n19882), .B2(n19049), .ZN(
        n13981) );
  OR2_X1 U17346 ( .A1(n13977), .A2(n13976), .ZN(n13979) );
  NAND2_X1 U17347 ( .A1(n13979), .A2(n13978), .ZN(n19957) );
  OAI22_X1 U17348 ( .A1(n16276), .A2(n19072), .B1(n19085), .B2(n19957), .ZN(
        n13980) );
  AOI211_X1 U17349 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19107), .A(n13981), .B(
        n13980), .ZN(n13984) );
  NAND2_X1 U17350 ( .A1(n13982), .A2(n19081), .ZN(n13983) );
  OAI211_X1 U17351 ( .C1(n19089), .C2(n19521), .A(n13984), .B(n13983), .ZN(
        n13985) );
  AOI21_X1 U17352 ( .B1(n13986), .B2(n14868), .A(n13985), .ZN(n13987) );
  INV_X1 U17353 ( .A(n13987), .ZN(P2_U2852) );
  NOR2_X1 U17354 ( .A1(n19092), .A2(n13988), .ZN(n14880) );
  XNOR2_X1 U17355 ( .A(n14880), .B(n19252), .ZN(n13989) );
  NAND2_X1 U17356 ( .A1(n13989), .A2(n19094), .ZN(n13996) );
  OAI22_X1 U17357 ( .A1(n19087), .A2(n10878), .B1(n19962), .B2(n19085), .ZN(
        n13991) );
  INV_X1 U17358 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19880) );
  NOR2_X1 U17359 ( .A1(n19049), .A2(n19880), .ZN(n13990) );
  AOI211_X1 U17360 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n19114), .A(
        n13991), .B(n13990), .ZN(n13992) );
  OAI21_X1 U17361 ( .B1(n13993), .B2(n19105), .A(n13992), .ZN(n13994) );
  AOI21_X1 U17362 ( .B1(n19256), .B2(n19081), .A(n13994), .ZN(n13995) );
  OAI211_X1 U17363 ( .C1(n19089), .C2(n19961), .A(n13996), .B(n13995), .ZN(
        P2_U2853) );
  AND2_X1 U17364 ( .A1(n20820), .A2(n21140), .ZN(n14012) );
  INV_X1 U17365 ( .A(n14012), .ZN(n13997) );
  AOI21_X1 U17366 ( .B1(n20183), .B2(n15756), .A(n13997), .ZN(n14009) );
  NAND2_X1 U17367 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20825), .ZN(n15726) );
  NAND2_X1 U17368 ( .A1(n20818), .A2(n13998), .ZN(n13999) );
  OAI211_X1 U17369 ( .C1(n15726), .C2(n20169), .A(n20055), .B(n13999), .ZN(
        n14000) );
  NAND2_X1 U17370 ( .A1(n20102), .A2(n20029), .ZN(n20030) );
  INV_X1 U17371 ( .A(n15708), .ZN(n14002) );
  NOR2_X1 U17372 ( .A1(n14005), .A2(n16083), .ZN(n14001) );
  OAI21_X1 U17373 ( .B1(n14003), .B2(n14002), .A(n15851), .ZN(n20106) );
  NAND2_X1 U17374 ( .A1(n20815), .A2(n14004), .ZN(n20101) );
  AND2_X2 U17375 ( .A1(n20029), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20098) );
  OAI21_X1 U17376 ( .B1(n20098), .B2(n20075), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14007) );
  OAI21_X1 U17377 ( .B1(n20101), .B2(n14008), .A(n14007), .ZN(n14018) );
  AND2_X1 U17378 ( .A1(n11036), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14011) );
  NOR2_X1 U17379 ( .A1(n14009), .A2(n14011), .ZN(n14010) );
  AND2_X2 U17380 ( .A1(n14015), .A2(n14010), .ZN(n20084) );
  INV_X1 U17381 ( .A(n14011), .ZN(n14013) );
  NOR2_X1 U17382 ( .A1(n14013), .A2(n14012), .ZN(n14014) );
  OAI22_X1 U17383 ( .A1(n14016), .A2(n20103), .B1(n20073), .B2(n14023), .ZN(
        n14017) );
  AOI211_X1 U17384 ( .C1(n20106), .C2(n14019), .A(n14018), .B(n14017), .ZN(
        n14020) );
  OAI21_X1 U17385 ( .B1(n15767), .B2(n14021), .A(n14020), .ZN(P1_U2840) );
  OAI222_X1 U17386 ( .A1(n14023), .A2(n15876), .B1(n14016), .B2(n14492), .C1(
        n14503), .C2(n14022), .ZN(P1_U2872) );
  AOI21_X1 U17387 ( .B1(n13955), .B2(n14025), .A(n14026), .ZN(n14027) );
  OR2_X1 U17388 ( .A1(n14024), .A2(n14027), .ZN(n14194) );
  AOI22_X1 U17389 ( .A1(n14279), .A2(n14526), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15891), .ZN(n14028) );
  OAI21_X1 U17390 ( .B1(n14194), .B2(n15896), .A(n14028), .ZN(P1_U2896) );
  XNOR2_X1 U17391 ( .A(n14029), .B(n14030), .ZN(n19238) );
  NAND2_X1 U17392 ( .A1(n14031), .A2(n13978), .ZN(n14033) );
  AND2_X1 U17393 ( .A1(n14033), .A2(n10078), .ZN(n19158) );
  NOR2_X1 U17394 ( .A1(n19236), .A2(n16313), .ZN(n14036) );
  INV_X1 U17395 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14179) );
  NAND2_X1 U17396 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19235), .ZN(n14034) );
  OAI221_X1 U17397 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14177), .C1(
        n14179), .C2(n14182), .A(n14034), .ZN(n14035) );
  AOI211_X1 U17398 ( .C1(n16307), .C2(n19158), .A(n14036), .B(n14035), .ZN(
        n14041) );
  XOR2_X1 U17399 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n14038), .Z(
        n14039) );
  XNOR2_X1 U17400 ( .A(n14037), .B(n14039), .ZN(n19240) );
  NAND2_X1 U17401 ( .A1(n19240), .A2(n16294), .ZN(n14040) );
  OAI211_X1 U17402 ( .C1(n19238), .C2(n16287), .A(n14041), .B(n14040), .ZN(
        P2_U3042) );
  INV_X1 U17403 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20040) );
  NOR3_X1 U17404 ( .A1(n20912), .A2(n13638), .A3(n21191), .ZN(n20067) );
  NAND2_X1 U17405 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20067), .ZN(n20053) );
  INV_X1 U17406 ( .A(n20053), .ZN(n20045) );
  NAND3_X1 U17407 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(n20045), .ZN(n20031) );
  NOR2_X1 U17408 ( .A1(n20040), .A2(n20031), .ZN(n14225) );
  INV_X1 U17409 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n14193) );
  NAND2_X1 U17410 ( .A1(n14225), .A2(n14193), .ZN(n14050) );
  NAND3_X1 U17411 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14225), .A3(n20029), 
        .ZN(n14472) );
  NAND2_X1 U17412 ( .A1(n20030), .A2(n14472), .ZN(n14043) );
  AOI22_X1 U17413 ( .A1(n20084), .A2(P1_EBX_REG_8__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20098), .ZN(n14042) );
  OAI211_X1 U17414 ( .C1(n14193), .C2(n14043), .A(n14042), .B(n20055), .ZN(
        n14044) );
  INV_X1 U17415 ( .A(n14044), .ZN(n14049) );
  NOR2_X1 U17416 ( .A1(n16066), .A2(n14045), .ZN(n14046) );
  OR2_X1 U17417 ( .A1(n14145), .A2(n14046), .ZN(n14139) );
  INV_X1 U17418 ( .A(n14139), .ZN(n14047) );
  AOI22_X1 U17419 ( .A1(n20096), .A2(n14047), .B1(n20075), .B2(n14197), .ZN(
        n14048) );
  OAI211_X1 U17420 ( .C1(n20102), .C2(n14050), .A(n14049), .B(n14048), .ZN(
        n14051) );
  INV_X1 U17421 ( .A(n14051), .ZN(n14052) );
  OAI21_X1 U17422 ( .B1(n15851), .B2(n14194), .A(n14052), .ZN(P1_U2832) );
  AOI21_X1 U17423 ( .B1(n14054), .B2(n14053), .A(n14076), .ZN(n19020) );
  INV_X1 U17424 ( .A(n19020), .ZN(n15236) );
  INV_X1 U17425 ( .A(n14055), .ZN(n14057) );
  OR2_X1 U17426 ( .A1(n14056), .A2(n14055), .ZN(n14078) );
  OAI211_X1 U17427 ( .C1(n14120), .C2(n14057), .A(n14984), .B(n14078), .ZN(
        n14059) );
  NAND2_X1 U17428 ( .A1(n14998), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n14058) );
  OAI211_X1 U17429 ( .C1(n15236), .C2(n14998), .A(n14059), .B(n14058), .ZN(
        P2_U2874) );
  INV_X1 U17430 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14060) );
  OAI222_X1 U17431 ( .A1(n14194), .A2(n14503), .B1(n14492), .B2(n14060), .C1(
        n14139), .C2(n15876), .ZN(P1_U2864) );
  INV_X1 U17432 ( .A(n20106), .ZN(n14074) );
  NAND2_X1 U17433 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n14061) );
  NAND2_X1 U17434 ( .A1(n20091), .A2(n14061), .ZN(n14062) );
  NAND2_X1 U17435 ( .A1(n20029), .A2(n14062), .ZN(n20090) );
  NAND2_X1 U17436 ( .A1(n20084), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n14066) );
  INV_X1 U17437 ( .A(n14063), .ZN(n14064) );
  AOI22_X1 U17438 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20098), .B1(
        n20075), .B2(n14064), .ZN(n14065) );
  OAI211_X1 U17439 ( .C1(n14067), .C2(n20101), .A(n14066), .B(n14065), .ZN(
        n14071) );
  NAND4_X1 U17440 ( .A1(n20091), .A2(n20912), .A3(P1_REIP_REG_2__SCAN_IN), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n14068) );
  OAI21_X1 U17441 ( .B1(n20073), .B2(n14069), .A(n14068), .ZN(n14070) );
  AOI211_X1 U17442 ( .C1(n20090), .C2(P1_REIP_REG_3__SCAN_IN), .A(n14071), .B(
        n14070), .ZN(n14072) );
  OAI21_X1 U17443 ( .B1(n14074), .B2(n14073), .A(n14072), .ZN(P1_U2837) );
  OAI21_X1 U17444 ( .B1(n14077), .B2(n14076), .A(n14075), .ZN(n16312) );
  INV_X1 U17445 ( .A(n14078), .ZN(n14081) );
  NAND2_X1 U17446 ( .A1(n14120), .A2(n14079), .ZN(n14159) );
  OAI211_X1 U17447 ( .C1(n14081), .C2(n14080), .A(n14984), .B(n14159), .ZN(
        n14083) );
  NAND2_X1 U17448 ( .A1(n14998), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14082) );
  OAI211_X1 U17449 ( .C1(n16312), .C2(n14980), .A(n14083), .B(n14082), .ZN(
        P2_U2873) );
  NOR2_X1 U17450 ( .A1(n14024), .A2(n14085), .ZN(n14086) );
  OR2_X1 U17451 ( .A1(n14084), .A2(n14086), .ZN(n14478) );
  AOI22_X1 U17452 ( .A1(n14279), .A2(n14522), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15891), .ZN(n14087) );
  OAI21_X1 U17453 ( .B1(n14478), .B2(n15896), .A(n14087), .ZN(P1_U2895) );
  NOR2_X1 U17454 ( .A1(n19092), .A2(n14088), .ZN(n14089) );
  XNOR2_X1 U17455 ( .A(n14089), .B(n16223), .ZN(n14090) );
  NAND2_X1 U17456 ( .A1(n14090), .A2(n19094), .ZN(n14097) );
  AOI21_X1 U17457 ( .B1(n14092), .B2(n14091), .A(n15417), .ZN(n15433) );
  INV_X1 U17458 ( .A(n15433), .ZN(n19133) );
  AOI22_X1 U17459 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19114), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19107), .ZN(n14093) );
  OAI211_X1 U17460 ( .C1(n19085), .C2(n19133), .A(n14093), .B(n19041), .ZN(
        n14095) );
  NOR2_X1 U17461 ( .A1(n19109), .A2(n15428), .ZN(n14094) );
  AOI211_X1 U17462 ( .C1(n19102), .C2(P2_REIP_REG_12__SCAN_IN), .A(n14095), 
        .B(n14094), .ZN(n14096) );
  OAI211_X1 U17463 ( .C1(n19105), .C2(n14098), .A(n14097), .B(n14096), .ZN(
        P2_U2843) );
  INV_X1 U17464 ( .A(n19945), .ZN(n19953) );
  NOR3_X1 U17465 ( .A1(n19842), .A2(n19323), .A3(n19953), .ZN(n14099) );
  AND2_X1 U17466 ( .A1(n19945), .A2(n19457), .ZN(n19948) );
  NOR2_X1 U17467 ( .A1(n14099), .A2(n19948), .ZN(n14115) );
  INV_X1 U17468 ( .A(n14115), .ZN(n14104) );
  NOR2_X1 U17469 ( .A1(n14100), .A2(n19960), .ZN(n19837) );
  NAND2_X1 U17470 ( .A1(n19960), .A2(n19968), .ZN(n19360) );
  INV_X1 U17471 ( .A(n19360), .ZN(n19327) );
  NAND2_X1 U17472 ( .A1(n19327), .A2(n19978), .ZN(n19304) );
  NOR2_X1 U17473 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19304), .ZN(
        n19293) );
  NOR2_X1 U17474 ( .A1(n19837), .A2(n19293), .ZN(n14114) );
  AOI21_X1 U17475 ( .B1(n14101), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14102) );
  OAI21_X1 U17476 ( .B1(n14102), .B2(n19293), .A(n19795), .ZN(n14103) );
  AOI22_X1 U17477 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19295), .ZN(n19818) );
  AOI22_X1 U17478 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19295), .ZN(n19728) );
  INV_X1 U17479 ( .A(n19323), .ZN(n14110) );
  NAND2_X1 U17480 ( .A1(n14108), .A2(n19291), .ZN(n19644) );
  INV_X1 U17481 ( .A(n19293), .ZN(n14109) );
  OAI22_X1 U17482 ( .A1(n19728), .A2(n14110), .B1(n19644), .B2(n14109), .ZN(
        n14111) );
  AOI21_X1 U17483 ( .B1(n19842), .B2(n19725), .A(n14111), .ZN(n14117) );
  OAI21_X1 U17484 ( .B1(n14112), .B2(n19293), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14113) );
  NOR2_X2 U17485 ( .A1(n19171), .A2(n19495), .ZN(n19814) );
  NAND2_X1 U17486 ( .A1(n19297), .A2(n19814), .ZN(n14116) );
  OAI211_X1 U17487 ( .C1(n19300), .C2(n14118), .A(n14117), .B(n14116), .ZN(
        P2_U3051) );
  AND2_X1 U17488 ( .A1(n14120), .A2(n14119), .ZN(n14158) );
  OAI21_X1 U17489 ( .B1(n14158), .B2(n14122), .A(n14121), .ZN(n15001) );
  INV_X1 U17490 ( .A(n15406), .ZN(n14123) );
  XNOR2_X1 U17491 ( .A(n14124), .B(n14123), .ZN(n15393) );
  INV_X1 U17492 ( .A(n15393), .ZN(n18989) );
  OAI22_X1 U17493 ( .A1(n15065), .A2(n18989), .B1(n19147), .B2(n14125), .ZN(
        n14127) );
  INV_X1 U17494 ( .A(n19121), .ZN(n15068) );
  INV_X1 U17495 ( .A(n16165), .ZN(n15066) );
  OAI22_X1 U17496 ( .A1(n15068), .A2(n18240), .B1(n19260), .B2(n15066), .ZN(
        n14126) );
  AOI211_X1 U17497 ( .C1(n19120), .C2(BUF1_REG_16__SCAN_IN), .A(n14127), .B(
        n14126), .ZN(n14128) );
  OAI21_X1 U17498 ( .B1(n15001), .B2(n19174), .A(n14128), .ZN(P2_U2903) );
  INV_X1 U17499 ( .A(n14025), .ZN(n14129) );
  XNOR2_X1 U17500 ( .A(n13955), .B(n14129), .ZN(n20113) );
  INV_X1 U17501 ( .A(n20113), .ZN(n14130) );
  OAI222_X1 U17502 ( .A1(n14549), .A2(n20219), .B1(n15896), .B2(n14130), .C1(
        n11233), .C2(n14551), .ZN(P1_U2897) );
  OAI21_X1 U17503 ( .B1(n14084), .B2(n14132), .A(n14131), .ZN(n15861) );
  AOI22_X1 U17504 ( .A1(n14279), .A2(n14519), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15891), .ZN(n14133) );
  OAI21_X1 U17505 ( .B1(n15861), .B2(n15896), .A(n14133), .ZN(P1_U2894) );
  XOR2_X1 U17506 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14134), .Z(
        n14135) );
  XNOR2_X1 U17507 ( .A(n14136), .B(n14135), .ZN(n14199) );
  INV_X1 U17508 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14137) );
  INV_X1 U17509 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16073) );
  NOR2_X1 U17510 ( .A1(n11824), .A2(n16048), .ZN(n16070) );
  OAI221_X1 U17511 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n14137), .C2(n16073), .A(
        n16070), .ZN(n14143) );
  OAI21_X1 U17512 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14712), .A(
        n14138), .ZN(n16062) );
  NOR2_X1 U17513 ( .A1(n20055), .A2(n14193), .ZN(n14141) );
  NOR2_X1 U17514 ( .A1(n16046), .A2(n14139), .ZN(n14140) );
  AOI211_X1 U17515 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n16062), .A(
        n14141), .B(n14140), .ZN(n14142) );
  OAI211_X1 U17516 ( .C1(n14199), .C2(n16052), .A(n14143), .B(n14142), .ZN(
        P1_U3023) );
  OAI21_X1 U17517 ( .B1(n14145), .B2(n14144), .A(n14155), .ZN(n14146) );
  INV_X1 U17518 ( .A(n14146), .ZN(n16056) );
  AOI22_X1 U17519 ( .A1(n20111), .A2(n16056), .B1(n14480), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n14147) );
  OAI21_X1 U17520 ( .B1(n14478), .B2(n14503), .A(n14147), .ZN(P1_U2863) );
  AOI22_X1 U17521 ( .A1(n20111), .A2(n20095), .B1(n14480), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n14148) );
  OAI21_X1 U17522 ( .B1(n14149), .B2(n14503), .A(n14148), .ZN(P1_U2871) );
  AOI22_X1 U17523 ( .A1(n20111), .A2(n20085), .B1(n14480), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n14150) );
  OAI21_X1 U17524 ( .B1(n14151), .B2(n14503), .A(n14150), .ZN(P1_U2870) );
  AOI22_X1 U17525 ( .A1(n20111), .A2(n20054), .B1(n14480), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n14152) );
  OAI21_X1 U17526 ( .B1(n14153), .B2(n14503), .A(n14152), .ZN(P1_U2867) );
  NAND2_X1 U17527 ( .A1(n14155), .A2(n14154), .ZN(n14156) );
  AND2_X1 U17528 ( .A1(n14213), .A2(n14156), .ZN(n15858) );
  AOI22_X1 U17529 ( .A1(n20111), .A2(n15858), .B1(n14480), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14157) );
  OAI21_X1 U17530 ( .B1(n15861), .B2(n14503), .A(n14157), .ZN(P1_U2862) );
  INV_X1 U17531 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n19000) );
  AOI211_X1 U17532 ( .C1(n14160), .C2(n14159), .A(n15000), .B(n14158), .ZN(
        n14161) );
  INV_X1 U17533 ( .A(n14161), .ZN(n14166) );
  NAND2_X1 U17534 ( .A1(n14162), .A2(n14075), .ZN(n14164) );
  INV_X1 U17535 ( .A(n14993), .ZN(n14163) );
  NAND2_X1 U17536 ( .A1(n14962), .A2(n18995), .ZN(n14165) );
  OAI211_X1 U17537 ( .C1(n14962), .C2(n19000), .A(n14166), .B(n14165), .ZN(
        P2_U2872) );
  XNOR2_X1 U17538 ( .A(n14167), .B(n14168), .ZN(n16262) );
  AND2_X1 U17539 ( .A1(n14170), .A2(n14169), .ZN(n14174) );
  AND2_X1 U17540 ( .A1(n14172), .A2(n14171), .ZN(n14173) );
  OAI22_X1 U17541 ( .A1(n14176), .A2(n14175), .B1(n14174), .B2(n14173), .ZN(
        n16261) );
  INV_X1 U17542 ( .A(n16261), .ZN(n14191) );
  AOI211_X1 U17543 ( .C1(n14181), .C2(n14179), .A(n14178), .B(n14177), .ZN(
        n14190) );
  INV_X1 U17544 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n14180) );
  OAI22_X1 U17545 ( .A1(n14182), .A2(n14181), .B1(n19041), .B2(n14180), .ZN(
        n14183) );
  INV_X1 U17546 ( .A(n14183), .ZN(n14188) );
  OAI21_X1 U17547 ( .B1(n14032), .B2(n14185), .A(n14184), .ZN(n19155) );
  INV_X1 U17548 ( .A(n19155), .ZN(n14186) );
  NAND2_X1 U17549 ( .A1(n14186), .A2(n16307), .ZN(n14187) );
  OAI211_X1 U17550 ( .C1(n16259), .C2(n16313), .A(n14188), .B(n14187), .ZN(
        n14189) );
  AOI211_X1 U17551 ( .C1(n14191), .C2(n16294), .A(n14190), .B(n14189), .ZN(
        n14192) );
  OAI21_X1 U17552 ( .B1(n16287), .B2(n16262), .A(n14192), .ZN(P2_U3041) );
  INV_X1 U17553 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20907) );
  OAI222_X1 U17554 ( .A1(n20041), .A2(n15876), .B1(n14492), .B2(n20907), .C1(
        n20044), .C2(n14503), .ZN(P1_U2866) );
  OAI22_X1 U17555 ( .A1(n15960), .A2(n11316), .B1(n20055), .B2(n14193), .ZN(
        n14196) );
  NOR2_X1 U17556 ( .A1(n14194), .A2(n15953), .ZN(n14195) );
  AOI211_X1 U17557 ( .C1(n15942), .C2(n14197), .A(n14196), .B(n14195), .ZN(
        n14198) );
  OAI21_X1 U17558 ( .B1(n15955), .B2(n14199), .A(n14198), .ZN(P1_U2991) );
  OAI21_X1 U17559 ( .B1(n10236), .B2(n9915), .A(n14200), .ZN(n14992) );
  XNOR2_X1 U17560 ( .A(n14202), .B(n14201), .ZN(n18978) );
  OAI22_X1 U17561 ( .A1(n15065), .A2(n18978), .B1(n19147), .B2(n14203), .ZN(
        n14206) );
  INV_X1 U17562 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14204) );
  OAI22_X1 U17563 ( .A1(n15068), .A2(n14204), .B1(n19265), .B2(n15066), .ZN(
        n14205) );
  AOI211_X1 U17564 ( .C1(n19120), .C2(BUF1_REG_17__SCAN_IN), .A(n14206), .B(
        n14205), .ZN(n14207) );
  OAI21_X1 U17565 ( .B1(n14992), .B2(n19174), .A(n14207), .ZN(P2_U2902) );
  NAND2_X1 U17566 ( .A1(n14210), .A2(n14211), .ZN(n14212) );
  NAND2_X1 U17567 ( .A1(n14209), .A2(n14212), .ZN(n14689) );
  AOI21_X1 U17568 ( .B1(n14214), .B2(n14213), .A(n9897), .ZN(n16032) );
  AOI22_X1 U17569 ( .A1(n20111), .A2(n16032), .B1(n14480), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n14215) );
  OAI21_X1 U17570 ( .B1(n14689), .B2(n14503), .A(n14215), .ZN(P1_U2861) );
  INV_X1 U17571 ( .A(n14217), .ZN(n14219) );
  AOI21_X1 U17572 ( .B1(n15918), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10112), .ZN(n14218) );
  OAI22_X1 U17573 ( .A1(n10112), .A2(n15938), .B1(n14219), .B2(n14218), .ZN(
        n16058) );
  NAND2_X1 U17574 ( .A1(n16058), .A2(n20013), .ZN(n14222) );
  NOR2_X1 U17575 ( .A1(n20055), .A2(n14474), .ZN(n16055) );
  NOR2_X1 U17576 ( .A1(n15954), .A2(n14469), .ZN(n14220) );
  AOI211_X1 U17577 ( .C1(n15946), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16055), .B(n14220), .ZN(n14221) );
  OAI211_X1 U17578 ( .C1(n15953), .C2(n14478), .A(n14222), .B(n14221), .ZN(
        P1_U2990) );
  INV_X1 U17579 ( .A(n14516), .ZN(n14223) );
  OAI222_X1 U17580 ( .A1(n14689), .A2(n15896), .B1(n20126), .B2(n14551), .C1(
        n14549), .C2(n14223), .ZN(P1_U2893) );
  INV_X1 U17581 ( .A(n14689), .ZN(n14224) );
  NAND2_X1 U17582 ( .A1(n14224), .A2(n20048), .ZN(n14231) );
  NAND2_X1 U17583 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n14226) );
  NOR2_X1 U17584 ( .A1(n15767), .A2(n14330), .ZN(n15862) );
  NAND3_X1 U17585 ( .A1(n20091), .A2(P1_REIP_REG_8__SCAN_IN), .A3(n14225), 
        .ZN(n14473) );
  INV_X1 U17586 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21053) );
  AOI22_X1 U17587 ( .A1(n20096), .A2(n16032), .B1(n20084), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n14227) );
  OAI211_X1 U17588 ( .C1(n15826), .C2(n14228), .A(n14227), .B(n20055), .ZN(
        n14229) );
  AOI221_X1 U17589 ( .B1(n15862), .B2(P1_REIP_REG_11__SCAN_IN), .C1(n15843), 
        .C2(n21053), .A(n14229), .ZN(n14230) );
  OAI211_X1 U17590 ( .C1(n20109), .C2(n14685), .A(n14231), .B(n14230), .ZN(
        P1_U2829) );
  AND2_X1 U17591 ( .A1(n14234), .A2(n14233), .ZN(n14235) );
  AND2_X1 U17592 ( .A1(n14209), .A2(n14235), .ZN(n14236) );
  OR2_X1 U17593 ( .A1(n14232), .A2(n14236), .ZN(n15852) );
  AOI22_X1 U17594 ( .A1(n14279), .A2(n14513), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15891), .ZN(n14237) );
  OAI21_X1 U17595 ( .B1(n15852), .B2(n15896), .A(n14237), .ZN(P1_U2892) );
  INV_X1 U17596 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n20975) );
  OR2_X1 U17597 ( .A1(n9897), .A2(n14238), .ZN(n14239) );
  NAND2_X1 U17598 ( .A1(n14791), .A2(n14239), .ZN(n15844) );
  OAI222_X1 U17599 ( .A1(n15852), .A2(n14503), .B1(n14492), .B2(n20975), .C1(
        n15844), .C2(n15876), .ZN(P1_U2860) );
  NOR2_X1 U17600 ( .A1(n14232), .A2(n14241), .ZN(n14242) );
  OR2_X1 U17601 ( .A1(n14240), .A2(n14242), .ZN(n15877) );
  AOI22_X1 U17602 ( .A1(n14279), .A2(n14509), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15891), .ZN(n14243) );
  OAI21_X1 U17603 ( .B1(n15877), .B2(n15896), .A(n14243), .ZN(P1_U2891) );
  AND2_X1 U17604 ( .A1(n14244), .A2(n14668), .ZN(n14652) );
  OAI22_X1 U17605 ( .A1(n14652), .A2(n14245), .B1(n15908), .B2(n14794), .ZN(
        n14247) );
  XNOR2_X1 U17606 ( .A(n11856), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14246) );
  XNOR2_X1 U17607 ( .A(n14247), .B(n14246), .ZN(n14666) );
  NOR2_X1 U17608 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14248), .ZN(
        n14260) );
  INV_X1 U17609 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14794) );
  NAND3_X1 U17610 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16049) );
  NOR3_X1 U17611 ( .A1(n15939), .A2(n11845), .A3(n16049), .ZN(n16035) );
  NAND2_X1 U17612 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16035), .ZN(
        n14271) );
  NOR2_X1 U17613 ( .A1(n14270), .A2(n14271), .ZN(n14254) );
  NOR2_X1 U17614 ( .A1(n14250), .A2(n14249), .ZN(n16043) );
  NAND2_X1 U17615 ( .A1(n14254), .A2(n16043), .ZN(n14758) );
  NOR2_X1 U17616 ( .A1(n14794), .A2(n14758), .ZN(n14693) );
  NAND2_X1 U17617 ( .A1(n14793), .A2(n14251), .ZN(n14252) );
  AND2_X1 U17618 ( .A1(n15823), .A2(n14252), .ZN(n14464) );
  INV_X1 U17619 ( .A(n14464), .ZN(n14258) );
  NOR2_X1 U17620 ( .A1(n14693), .A2(n14757), .ZN(n14768) );
  AND3_X1 U17621 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n14253), .ZN(n14267) );
  NAND2_X1 U17622 ( .A1(n14267), .A2(n14254), .ZN(n14759) );
  NOR2_X1 U17623 ( .A1(n14794), .A2(n14759), .ZN(n14690) );
  OAI21_X1 U17624 ( .B1(n14266), .B2(n14690), .A(n14255), .ZN(n14767) );
  OR2_X1 U17625 ( .A1(n14768), .A2(n14767), .ZN(n14799) );
  NAND2_X1 U17626 ( .A1(n14799), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14257) );
  INV_X1 U17627 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14256) );
  OR2_X1 U17628 ( .A1(n20055), .A2(n14256), .ZN(n14661) );
  OAI211_X1 U17629 ( .C1(n16046), .C2(n14258), .A(n14257), .B(n14661), .ZN(
        n14259) );
  AOI21_X1 U17630 ( .B1(n14260), .B2(n14693), .A(n14259), .ZN(n14261) );
  OAI21_X1 U17631 ( .B1(n14666), .B2(n16052), .A(n14261), .ZN(P1_U3017) );
  OR2_X1 U17632 ( .A1(n14244), .A2(n14262), .ZN(n14669) );
  OAI21_X1 U17633 ( .B1(n14263), .B2(n15908), .A(n14669), .ZN(n14265) );
  AOI21_X1 U17634 ( .B1(n15918), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14667), .ZN(n14264) );
  XNOR2_X1 U17635 ( .A(n14265), .B(n14264), .ZN(n14681) );
  AOI21_X1 U17636 ( .B1(n14267), .B2(n16035), .A(n14266), .ZN(n14269) );
  AOI211_X1 U17637 ( .C1(n14692), .C2(n14271), .A(n14269), .B(n14268), .ZN(
        n16039) );
  AOI221_X1 U17638 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16039), 
        .C1(n14760), .C2(n16039), .A(n14270), .ZN(n14274) );
  NOR3_X1 U17639 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14271), .A3(
        n16048), .ZN(n14273) );
  NAND2_X1 U17640 ( .A1(n20070), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n14676) );
  OAI21_X1 U17641 ( .B1(n16046), .B2(n15844), .A(n14676), .ZN(n14272) );
  NOR3_X1 U17642 ( .A1(n14274), .A2(n14273), .A3(n14272), .ZN(n14275) );
  OAI21_X1 U17643 ( .B1(n14681), .B2(n16052), .A(n14275), .ZN(P1_U3019) );
  OAI21_X1 U17644 ( .B1(n14240), .B2(n14277), .A(n14276), .ZN(n14458) );
  AOI22_X1 U17645 ( .A1(n14464), .A2(n20111), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14480), .ZN(n14278) );
  OAI21_X1 U17646 ( .B1(n14458), .B2(n14503), .A(n14278), .ZN(P1_U2858) );
  AOI22_X1 U17647 ( .A1(n14279), .A2(n14506), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15891), .ZN(n14280) );
  OAI21_X1 U17648 ( .B1(n14458), .B2(n15896), .A(n14280), .ZN(P1_U2890) );
  INV_X1 U17649 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n14282) );
  INV_X1 U17650 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n14283) );
  INV_X1 U17651 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16878) );
  NAND2_X1 U17652 ( .A1(n14281), .A2(n17252), .ZN(n17239) );
  NOR2_X1 U17653 ( .A1(n14283), .A2(n17239), .ZN(n17242) );
  NAND2_X1 U17654 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17242), .ZN(n17172) );
  NOR3_X1 U17655 ( .A1(n14282), .A2(n15628), .A3(n17172), .ZN(n17136) );
  INV_X1 U17656 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n15627) );
  INV_X1 U17657 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16820) );
  NOR4_X1 U17658 ( .A1(n18272), .A2(n16820), .A3(n14283), .A4(n17239), .ZN(
        n17187) );
  NAND3_X1 U17659 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n17187), .ZN(n17155) );
  NOR2_X1 U17660 ( .A1(n15627), .A2(n17155), .ZN(n14284) );
  AOI21_X1 U17661 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n14284), .A(
        P3_EBX_REG_14__SCAN_IN), .ZN(n14285) );
  NOR2_X1 U17662 ( .A1(n17136), .A2(n14285), .ZN(n14299) );
  INV_X1 U17663 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14287) );
  AOI22_X1 U17664 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14286) );
  OAI21_X1 U17665 ( .B1(n12697), .B2(n14287), .A(n14286), .ZN(n14297) );
  INV_X1 U17666 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14295) );
  AOI22_X1 U17667 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14294) );
  OAI22_X1 U17668 ( .A1(n17218), .A2(n17011), .B1(n17227), .B2(n17251), .ZN(
        n14292) );
  AOI22_X1 U17669 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14290) );
  AOI22_X1 U17670 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14289) );
  AOI22_X1 U17671 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14288) );
  NAND3_X1 U17672 ( .A1(n14290), .A2(n14289), .A3(n14288), .ZN(n14291) );
  AOI211_X1 U17673 ( .C1(n17235), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n14292), .B(n14291), .ZN(n14293) );
  OAI211_X1 U17674 ( .C1(n17150), .C2(n14295), .A(n14294), .B(n14293), .ZN(
        n14296) );
  AOI211_X1 U17675 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n14297), .B(n14296), .ZN(n17373) );
  INV_X1 U17676 ( .A(n17373), .ZN(n14298) );
  MUX2_X1 U17677 ( .A(n14299), .B(n14298), .S(n17275), .Z(P3_U2689) );
  NOR2_X1 U17678 ( .A1(n11040), .A2(n20165), .ZN(n14300) );
  NAND2_X1 U17679 ( .A1(n14551), .A2(n14300), .ZN(n15900) );
  INV_X1 U17680 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20220) );
  AND2_X1 U17681 ( .A1(n14551), .A2(n20221), .ZN(n14301) );
  NAND2_X1 U17682 ( .A1(n14323), .A2(n14301), .ZN(n14304) );
  NOR2_X1 U17683 ( .A1(n11040), .A2(n20164), .ZN(n14302) );
  AOI22_X1 U17684 ( .A1(n15887), .A2(DATAI_31_), .B1(n15891), .B2(
        P1_EAX_REG_31__SCAN_IN), .ZN(n14303) );
  OAI211_X1 U17685 ( .C1(n15900), .C2(n20220), .A(n14304), .B(n14303), .ZN(
        P1_U2873) );
  NAND2_X1 U17686 ( .A1(n14305), .A2(n15085), .ZN(n14308) );
  NOR2_X1 U17687 ( .A1(n14306), .A2(n10253), .ZN(n14307) );
  XNOR2_X1 U17688 ( .A(n14308), .B(n14307), .ZN(n15083) );
  XNOR2_X1 U17689 ( .A(n15089), .B(n14314), .ZN(n15081) );
  INV_X1 U17690 ( .A(n14309), .ZN(n14312) );
  NAND2_X1 U17691 ( .A1(n14314), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14310) );
  NAND2_X1 U17692 ( .A1(n19076), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15074) );
  OAI21_X1 U17693 ( .B1(n15253), .B2(n14310), .A(n15074), .ZN(n14311) );
  AOI21_X1 U17694 ( .B1(n16307), .B2(n14312), .A(n14311), .ZN(n14317) );
  INV_X1 U17695 ( .A(n15079), .ZN(n14313) );
  NAND2_X1 U17696 ( .A1(n14313), .A2(n16296), .ZN(n14316) );
  NAND3_X1 U17697 ( .A1(n14317), .A2(n14316), .A3(n10241), .ZN(n14318) );
  OAI21_X1 U17698 ( .B1(n15083), .B2(n16287), .A(n14319), .ZN(P2_U3016) );
  NOR2_X1 U17699 ( .A1(n15079), .A2(n14980), .ZN(n14320) );
  AOI21_X1 U17700 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14980), .A(n14320), .ZN(
        n14321) );
  OAI21_X1 U17701 ( .B1(n14322), .B2(n15000), .A(n14321), .ZN(P2_U2857) );
  INV_X1 U17702 ( .A(n14323), .ZN(n14344) );
  AOI22_X1 U17703 ( .A1(n14324), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n15709), .ZN(n14329) );
  XOR2_X1 U17704 ( .A(n14329), .B(n14328), .Z(n14699) );
  NAND2_X1 U17705 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14338) );
  INV_X1 U17706 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21172) );
  NAND3_X1 U17707 ( .A1(n14330), .A2(P1_REIP_REG_11__SCAN_IN), .A3(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15834) );
  NAND4_X1 U17708 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14447), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_15__SCAN_IN), .ZN(n15788) );
  NAND2_X1 U17709 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15787) );
  INV_X1 U17710 ( .A(n15787), .ZN(n14331) );
  NAND2_X1 U17711 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14331), .ZN(n14332) );
  AND3_X1 U17712 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(P1_REIP_REG_23__SCAN_IN), .ZN(n14333) );
  NAND2_X1 U17713 ( .A1(n15766), .A2(n14333), .ZN(n14406) );
  NAND2_X1 U17714 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14334) );
  INV_X1 U17715 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21040) );
  NOR2_X2 U17716 ( .A1(n14385), .A2(n21040), .ZN(n14373) );
  AND2_X1 U17717 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14335) );
  NOR2_X1 U17718 ( .A1(n14336), .A2(n15767), .ZN(n14366) );
  AOI21_X1 U17719 ( .B1(n20030), .B2(n14338), .A(n14366), .ZN(n14349) );
  AOI22_X1 U17720 ( .A1(n20084), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20098), .ZN(n14341) );
  INV_X1 U17721 ( .A(n14336), .ZN(n14337) );
  NOR2_X1 U17722 ( .A1(n14337), .A2(n20102), .ZN(n14354) );
  INV_X1 U17723 ( .A(n14338), .ZN(n14339) );
  NAND3_X1 U17724 ( .A1(n14354), .A2(n14339), .A3(n21183), .ZN(n14340) );
  OAI211_X1 U17725 ( .C1(n14349), .C2(n21183), .A(n14341), .B(n14340), .ZN(
        n14342) );
  AOI21_X1 U17726 ( .B1(n14699), .B2(n20096), .A(n14342), .ZN(n14343) );
  OAI21_X1 U17727 ( .B1(n14344), .B2(n15851), .A(n14343), .ZN(P1_U2809) );
  INV_X1 U17728 ( .A(n14345), .ZN(n14721) );
  AOI21_X1 U17729 ( .B1(n14354), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14348) );
  AOI22_X1 U17730 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20098), .B1(
        n20075), .B2(n14555), .ZN(n14347) );
  NAND2_X1 U17731 ( .A1(n20084), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14346) );
  OAI211_X1 U17732 ( .C1(n14349), .C2(n14348), .A(n14347), .B(n14346), .ZN(
        n14350) );
  AOI21_X1 U17733 ( .B1(n14721), .B2(n20096), .A(n14350), .ZN(n14351) );
  OAI21_X1 U17734 ( .B1(n14561), .B2(n15851), .A(n14351), .ZN(P1_U2810) );
  OAI22_X1 U17735 ( .A1(n14352), .A2(n15826), .B1(n20109), .B2(n14566), .ZN(
        n14353) );
  AOI21_X1 U17736 ( .B1(n20084), .B2(P1_EBX_REG_29__SCAN_IN), .A(n14353), .ZN(
        n14356) );
  INV_X1 U17737 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20908) );
  NAND2_X1 U17738 ( .A1(n14354), .A2(n20908), .ZN(n14355) );
  OAI211_X1 U17739 ( .C1(n14730), .C2(n20073), .A(n14356), .B(n14355), .ZN(
        n14357) );
  AOI21_X1 U17740 ( .B1(n14366), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14357), 
        .ZN(n14358) );
  OAI21_X1 U17741 ( .B1(n14512), .B2(n15851), .A(n14358), .ZN(P1_U2811) );
  OR2_X1 U17742 ( .A1(n14376), .A2(n14360), .ZN(n14361) );
  NAND2_X1 U17743 ( .A1(n14362), .A2(n14361), .ZN(n14739) );
  INV_X1 U17744 ( .A(n14739), .ZN(n14365) );
  INV_X1 U17745 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n20924) );
  AOI22_X1 U17746 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20098), .B1(
        n20075), .B2(n14575), .ZN(n14363) );
  OAI21_X1 U17747 ( .B1(n20103), .B2(n20924), .A(n14363), .ZN(n14364) );
  AOI21_X1 U17748 ( .B1(n14365), .B2(n20096), .A(n14364), .ZN(n14369) );
  INV_X1 U17749 ( .A(n14373), .ZN(n14374) );
  INV_X1 U17750 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21046) );
  NOR2_X1 U17751 ( .A1(n14374), .A2(n21046), .ZN(n14367) );
  OAI21_X1 U17752 ( .B1(n14367), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14366), 
        .ZN(n14368) );
  OAI211_X1 U17753 ( .C1(n14580), .C2(n15851), .A(n14369), .B(n14368), .ZN(
        P1_U2812) );
  AOI21_X1 U17754 ( .B1(n14371), .B2(n14370), .A(n14359), .ZN(n14372) );
  NOR2_X1 U17755 ( .A1(n14373), .A2(n15767), .ZN(n14392) );
  NOR3_X1 U17756 ( .A1(n14374), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n20102), 
        .ZN(n14381) );
  INV_X1 U17757 ( .A(n14399), .ZN(n14387) );
  AOI21_X1 U17758 ( .B1(n14387), .B2(n14386), .A(n14375), .ZN(n14377) );
  NOR2_X1 U17759 ( .A1(n14377), .A2(n14376), .ZN(n14481) );
  INV_X1 U17760 ( .A(n14481), .ZN(n14748) );
  AOI22_X1 U17761 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20098), .B1(
        n20075), .B2(n14585), .ZN(n14379) );
  NAND2_X1 U17762 ( .A1(n20084), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n14378) );
  OAI211_X1 U17763 ( .C1(n14748), .C2(n20073), .A(n14379), .B(n14378), .ZN(
        n14380) );
  AOI211_X1 U17764 ( .C1(n14392), .C2(P1_REIP_REG_27__SCAN_IN), .A(n14381), 
        .B(n14380), .ZN(n14382) );
  OAI21_X1 U17765 ( .B1(n14590), .B2(n15851), .A(n14382), .ZN(P1_U2813) );
  NAND2_X1 U17766 ( .A1(n21040), .A2(n14385), .ZN(n14391) );
  XNOR2_X1 U17767 ( .A(n14387), .B(n14386), .ZN(n15962) );
  AOI22_X1 U17768 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20098), .B1(
        n20075), .B2(n14599), .ZN(n14389) );
  NAND2_X1 U17769 ( .A1(n20084), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14388) );
  OAI211_X1 U17770 ( .C1(n15962), .C2(n20073), .A(n14389), .B(n14388), .ZN(
        n14390) );
  AOI21_X1 U17771 ( .B1(n14392), .B2(n14391), .A(n14390), .ZN(n14393) );
  OAI21_X1 U17772 ( .B1(n14597), .B2(n15851), .A(n14393), .ZN(P1_U2814) );
  INV_X1 U17773 ( .A(n14394), .ZN(n14397) );
  INV_X1 U17774 ( .A(n14395), .ZN(n14411) );
  AOI21_X1 U17775 ( .B1(n14397), .B2(n14411), .A(n14396), .ZN(n14609) );
  INV_X1 U17776 ( .A(n14609), .ZN(n14525) );
  INV_X1 U17777 ( .A(n14414), .ZN(n14401) );
  INV_X1 U17778 ( .A(n14398), .ZN(n14400) );
  OAI21_X1 U17779 ( .B1(n14401), .B2(n14400), .A(n14399), .ZN(n14484) );
  INV_X1 U17780 ( .A(n14484), .ZN(n15974) );
  INV_X1 U17781 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21036) );
  NOR4_X1 U17782 ( .A1(n14406), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n21036), 
        .A4(n20102), .ZN(n14405) );
  INV_X1 U17783 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21047) );
  INV_X1 U17784 ( .A(n14607), .ZN(n14402) );
  AOI22_X1 U17785 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20098), .B1(
        n20075), .B2(n14402), .ZN(n14403) );
  OAI21_X1 U17786 ( .B1(n20103), .B2(n21047), .A(n14403), .ZN(n14404) );
  AOI211_X1 U17787 ( .C1(n15974), .C2(n20096), .A(n14405), .B(n14404), .ZN(
        n14408) );
  NOR3_X1 U17788 ( .A1(n14406), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n20102), 
        .ZN(n14418) );
  AND2_X1 U17789 ( .A1(n14406), .A2(n20030), .ZN(n14429) );
  OAI21_X1 U17790 ( .B1(n14418), .B2(n14429), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14407) );
  OAI211_X1 U17791 ( .C1(n14525), .C2(n15851), .A(n14408), .B(n14407), .ZN(
        P1_U2815) );
  OR2_X1 U17792 ( .A1(n14425), .A2(n14412), .ZN(n14413) );
  NAND2_X1 U17793 ( .A1(n14414), .A2(n14413), .ZN(n15981) );
  AOI22_X1 U17794 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20098), .B1(
        n20075), .B2(n14613), .ZN(n14416) );
  NAND2_X1 U17795 ( .A1(n20084), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14415) );
  OAI211_X1 U17796 ( .C1(n15981), .C2(n20073), .A(n14416), .B(n14415), .ZN(
        n14417) );
  AOI211_X1 U17797 ( .C1(n14429), .C2(P1_REIP_REG_24__SCAN_IN), .A(n14418), 
        .B(n14417), .ZN(n14419) );
  OAI21_X1 U17798 ( .B1(n14620), .B2(n15851), .A(n14419), .ZN(P1_U2816) );
  AOI21_X1 U17799 ( .B1(n14421), .B2(n14420), .A(n14410), .ZN(n14627) );
  INV_X1 U17800 ( .A(n14627), .ZN(n14532) );
  INV_X1 U17801 ( .A(n14422), .ZN(n14625) );
  OAI22_X1 U17802 ( .A1(n11588), .A2(n15826), .B1(n20109), .B2(n14625), .ZN(
        n14427) );
  NOR2_X1 U17803 ( .A1(n9882), .A2(n14423), .ZN(n14424) );
  OR2_X1 U17804 ( .A1(n14425), .A2(n14424), .ZN(n15988) );
  NOR2_X1 U17805 ( .A1(n15988), .A2(n20073), .ZN(n14426) );
  AOI211_X1 U17806 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n20084), .A(n14427), .B(
        n14426), .ZN(n14432) );
  NAND2_X1 U17807 ( .A1(n15766), .A2(n20091), .ZN(n15771) );
  NAND2_X1 U17808 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14428) );
  NOR2_X1 U17809 ( .A1(n15771), .A2(n14428), .ZN(n14430) );
  OAI21_X1 U17810 ( .B1(n14430), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14429), 
        .ZN(n14431) );
  OAI211_X1 U17811 ( .C1(n14532), .C2(n15851), .A(n14432), .B(n14431), .ZN(
        P1_U2817) );
  OAI21_X1 U17812 ( .B1(n14433), .B2(n14434), .A(n14420), .ZN(n14634) );
  XOR2_X1 U17813 ( .A(P1_REIP_REG_22__SCAN_IN), .B(P1_REIP_REG_21__SCAN_IN), 
        .Z(n14442) );
  INV_X1 U17814 ( .A(n15771), .ZN(n14441) );
  AND2_X1 U17815 ( .A1(n15739), .A2(n14435), .ZN(n14436) );
  OR2_X1 U17816 ( .A1(n14436), .A2(n9882), .ZN(n15996) );
  AOI22_X1 U17817 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20098), .B1(
        n20075), .B2(n14637), .ZN(n14438) );
  NAND2_X1 U17818 ( .A1(n20084), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n14437) );
  OAI211_X1 U17819 ( .C1(n15996), .C2(n20073), .A(n14438), .B(n14437), .ZN(
        n14440) );
  INV_X1 U17820 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14632) );
  NOR3_X1 U17821 ( .A1(n15766), .A2(n15767), .A3(n14632), .ZN(n14439) );
  AOI211_X1 U17822 ( .C1(n14442), .C2(n14441), .A(n14440), .B(n14439), .ZN(
        n14443) );
  OAI21_X1 U17823 ( .B1(n14634), .B2(n15851), .A(n14443), .ZN(P1_U2818) );
  INV_X1 U17824 ( .A(n14444), .ZN(n14446) );
  OAI21_X1 U17825 ( .B1(n10243), .B2(n14446), .A(n14445), .ZN(n14546) );
  INV_X1 U17826 ( .A(n14546), .ZN(n14658) );
  INV_X1 U17827 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21138) );
  NAND3_X1 U17828 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(n15843), .ZN(n15842) );
  NOR2_X1 U17829 ( .A1(n21172), .A2(n15842), .ZN(n14459) );
  NAND2_X1 U17830 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n14459), .ZN(n15777) );
  NOR3_X1 U17831 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n21138), .A3(n15777), 
        .ZN(n14456) );
  NOR2_X1 U17832 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15777), .ZN(n15830) );
  OAI21_X1 U17833 ( .B1(n10251), .B2(n15830), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14454) );
  OR2_X1 U17834 ( .A1(n15822), .A2(n14448), .ZN(n14449) );
  NAND2_X1 U17835 ( .A1(n15812), .A2(n14449), .ZN(n14502) );
  INV_X1 U17836 ( .A(n14502), .ZN(n14786) );
  AOI22_X1 U17837 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n20084), .B1(n20096), 
        .B2(n14786), .ZN(n14450) );
  OAI211_X1 U17838 ( .C1(n15826), .C2(n14451), .A(n14450), .B(n20055), .ZN(
        n14452) );
  INV_X1 U17839 ( .A(n14452), .ZN(n14453) );
  OAI211_X1 U17840 ( .C1(n20109), .C2(n14656), .A(n14454), .B(n14453), .ZN(
        n14455) );
  AOI211_X1 U17841 ( .C1(n14658), .C2(n20048), .A(n14456), .B(n14455), .ZN(
        n14457) );
  INV_X1 U17842 ( .A(n14457), .ZN(P1_U2824) );
  INV_X1 U17843 ( .A(n14458), .ZN(n14664) );
  NAND2_X1 U17844 ( .A1(n14664), .A2(n20048), .ZN(n14468) );
  OAI21_X1 U17845 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14459), .A(n10251), 
        .ZN(n14467) );
  INV_X1 U17846 ( .A(n14662), .ZN(n14460) );
  NAND2_X1 U17847 ( .A1(n20075), .A2(n14460), .ZN(n14462) );
  NAND2_X1 U17848 ( .A1(n20098), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14461) );
  NAND3_X1 U17849 ( .A1(n14462), .A2(n14461), .A3(n20055), .ZN(n14463) );
  AOI21_X1 U17850 ( .B1(n20084), .B2(P1_EBX_REG_14__SCAN_IN), .A(n14463), .ZN(
        n14466) );
  NAND2_X1 U17851 ( .A1(n20096), .A2(n14464), .ZN(n14465) );
  NAND4_X1 U17852 ( .A1(n14468), .A2(n14467), .A3(n14466), .A4(n14465), .ZN(
        P1_U2826) );
  NOR2_X1 U17853 ( .A1(n20109), .A2(n14469), .ZN(n14470) );
  AOI211_X1 U17854 ( .C1(n20098), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20070), .B(n14470), .ZN(n14471) );
  OAI21_X1 U17855 ( .B1(n20921), .B2(n20103), .A(n14471), .ZN(n14476) );
  INV_X1 U17856 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14474) );
  AOI21_X1 U17857 ( .B1(n20030), .B2(n14472), .A(n14474), .ZN(n15863) );
  AOI21_X1 U17858 ( .B1(n14474), .B2(n14473), .A(n15863), .ZN(n14475) );
  AOI211_X1 U17859 ( .C1(n16056), .C2(n20096), .A(n14476), .B(n14475), .ZN(
        n14477) );
  OAI21_X1 U17860 ( .B1(n15851), .B2(n14478), .A(n14477), .ZN(P1_U2831) );
  INV_X1 U17861 ( .A(n14699), .ZN(n14479) );
  INV_X1 U17862 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n20986) );
  OAI22_X1 U17863 ( .A1(n14479), .A2(n15876), .B1(n14492), .B2(n20986), .ZN(
        P1_U2841) );
  OAI222_X1 U17864 ( .A1(n14739), .A2(n15876), .B1(n20924), .B2(n14492), .C1(
        n14580), .C2(n14503), .ZN(P1_U2844) );
  AOI22_X1 U17865 ( .A1(n14481), .A2(n20111), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n14480), .ZN(n14482) );
  OAI21_X1 U17866 ( .B1(n14590), .B2(n14503), .A(n14482), .ZN(P1_U2845) );
  OAI222_X1 U17867 ( .A1(n14503), .A2(n14597), .B1(n14483), .B2(n14492), .C1(
        n15876), .C2(n15962), .ZN(P1_U2846) );
  OAI222_X1 U17868 ( .A1(n14484), .A2(n15876), .B1(n21047), .B2(n14492), .C1(
        n14525), .C2(n14503), .ZN(P1_U2847) );
  OAI222_X1 U17869 ( .A1(n15981), .A2(n15876), .B1(n21128), .B2(n14492), .C1(
        n14620), .C2(n14503), .ZN(P1_U2848) );
  INV_X1 U17870 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14485) );
  OAI222_X1 U17871 ( .A1(n15988), .A2(n15876), .B1(n14485), .B2(n14492), .C1(
        n14532), .C2(n14503), .ZN(P1_U2849) );
  INV_X1 U17872 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14486) );
  OAI222_X1 U17873 ( .A1(n15996), .A2(n15876), .B1(n14486), .B2(n14492), .C1(
        n14634), .C2(n14503), .ZN(P1_U2850) );
  AOI21_X1 U17874 ( .B1(n14489), .B2(n15791), .A(n14488), .ZN(n14490) );
  INV_X1 U17875 ( .A(n14490), .ZN(n15780) );
  INV_X1 U17876 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n20977) );
  OAI21_X1 U17877 ( .B1(n15793), .B2(n14491), .A(n15737), .ZN(n15779) );
  OAI222_X1 U17878 ( .A1(n15780), .A2(n14503), .B1(n14492), .B2(n20977), .C1(
        n15779), .C2(n15876), .ZN(P1_U2852) );
  OAI21_X1 U17879 ( .B1(n14493), .B2(n14496), .A(n14495), .ZN(n15802) );
  INV_X1 U17880 ( .A(n14497), .ZN(n15794) );
  NAND2_X1 U17881 ( .A1(n15814), .A2(n14498), .ZN(n14499) );
  NAND2_X1 U17882 ( .A1(n15794), .A2(n14499), .ZN(n15801) );
  OAI22_X1 U17883 ( .A1(n15801), .A2(n15876), .B1(n21008), .B2(n14492), .ZN(
        n14500) );
  INV_X1 U17884 ( .A(n14500), .ZN(n14501) );
  OAI21_X1 U17885 ( .B1(n15802), .B2(n14503), .A(n14501), .ZN(P1_U2854) );
  INV_X1 U17886 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21050) );
  OAI222_X1 U17887 ( .A1(n14546), .A2(n14503), .B1(n14492), .B2(n21050), .C1(
        n14502), .C2(n15876), .ZN(P1_U2856) );
  AOI22_X1 U17888 ( .A1(n15887), .A2(DATAI_30_), .B1(n15891), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14508) );
  NOR3_X1 U17889 ( .A1(n15891), .A2(n20221), .A3(n11031), .ZN(n14505) );
  AOI22_X1 U17890 ( .A1(n15893), .A2(n14506), .B1(BUF1_REG_30__SCAN_IN), .B2(
        n14543), .ZN(n14507) );
  OAI211_X1 U17891 ( .C1(n14561), .C2(n15896), .A(n14508), .B(n14507), .ZN(
        P1_U2874) );
  AOI22_X1 U17892 ( .A1(n15887), .A2(DATAI_29_), .B1(n15891), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14511) );
  AOI22_X1 U17893 ( .A1(n15893), .A2(n14509), .B1(BUF1_REG_29__SCAN_IN), .B2(
        n14543), .ZN(n14510) );
  OAI211_X1 U17894 ( .C1(n14512), .C2(n15896), .A(n14511), .B(n14510), .ZN(
        P1_U2875) );
  AOI22_X1 U17895 ( .A1(n15887), .A2(DATAI_28_), .B1(n15891), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14515) );
  AOI22_X1 U17896 ( .A1(n15893), .A2(n14513), .B1(BUF1_REG_28__SCAN_IN), .B2(
        n14543), .ZN(n14514) );
  OAI211_X1 U17897 ( .C1(n14580), .C2(n15896), .A(n14515), .B(n14514), .ZN(
        P1_U2876) );
  AOI22_X1 U17898 ( .A1(n15887), .A2(DATAI_27_), .B1(n15891), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n14518) );
  AOI22_X1 U17899 ( .A1(n15893), .A2(n14516), .B1(BUF1_REG_27__SCAN_IN), .B2(
        n14543), .ZN(n14517) );
  OAI211_X1 U17900 ( .C1(n14590), .C2(n15896), .A(n14518), .B(n14517), .ZN(
        P1_U2877) );
  AOI22_X1 U17901 ( .A1(n15887), .A2(DATAI_26_), .B1(n15891), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n14521) );
  AOI22_X1 U17902 ( .A1(n15893), .A2(n14519), .B1(BUF1_REG_26__SCAN_IN), .B2(
        n14543), .ZN(n14520) );
  OAI211_X1 U17903 ( .C1(n14597), .C2(n15896), .A(n14521), .B(n14520), .ZN(
        P1_U2878) );
  AOI22_X1 U17904 ( .A1(n15887), .A2(DATAI_25_), .B1(n15891), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14524) );
  AOI22_X1 U17905 ( .A1(n15893), .A2(n14522), .B1(n14543), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14523) );
  OAI211_X1 U17906 ( .C1(n14525), .C2(n15896), .A(n14524), .B(n14523), .ZN(
        P1_U2879) );
  AOI22_X1 U17907 ( .A1(n15887), .A2(DATAI_24_), .B1(n15891), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n14528) );
  AOI22_X1 U17908 ( .A1(n15893), .A2(n14526), .B1(n14543), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14527) );
  OAI211_X1 U17909 ( .C1(n14620), .C2(n15896), .A(n14528), .B(n14527), .ZN(
        P1_U2880) );
  AOI22_X1 U17910 ( .A1(n15893), .A2(n14529), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n15891), .ZN(n14531) );
  AOI22_X1 U17911 ( .A1(n14543), .A2(BUF1_REG_23__SCAN_IN), .B1(n15887), .B2(
        DATAI_23_), .ZN(n14530) );
  OAI211_X1 U17912 ( .C1(n14532), .C2(n15896), .A(n14531), .B(n14530), .ZN(
        P1_U2881) );
  AOI22_X1 U17913 ( .A1(n15893), .A2(n14533), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n15891), .ZN(n14535) );
  AOI22_X1 U17914 ( .A1(n14543), .A2(BUF1_REG_22__SCAN_IN), .B1(n15887), .B2(
        DATAI_22_), .ZN(n14534) );
  OAI211_X1 U17915 ( .C1(n14634), .C2(n15896), .A(n14535), .B(n14534), .ZN(
        P1_U2882) );
  AOI22_X1 U17916 ( .A1(n15893), .A2(n14536), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n15891), .ZN(n14538) );
  AOI22_X1 U17917 ( .A1(n14543), .A2(BUF1_REG_20__SCAN_IN), .B1(n15887), .B2(
        DATAI_20_), .ZN(n14537) );
  OAI211_X1 U17918 ( .C1(n15780), .C2(n15896), .A(n14538), .B(n14537), .ZN(
        P1_U2884) );
  AOI22_X1 U17919 ( .A1(n15893), .A2(n14539), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n15891), .ZN(n14541) );
  AOI22_X1 U17920 ( .A1(n14543), .A2(BUF1_REG_18__SCAN_IN), .B1(n15887), .B2(
        DATAI_18_), .ZN(n14540) );
  OAI211_X1 U17921 ( .C1(n15802), .C2(n15896), .A(n14541), .B(n14540), .ZN(
        P1_U2886) );
  AOI22_X1 U17922 ( .A1(n15893), .A2(n14542), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15891), .ZN(n14545) );
  AOI22_X1 U17923 ( .A1(n14543), .A2(BUF1_REG_16__SCAN_IN), .B1(n15887), .B2(
        DATAI_16_), .ZN(n14544) );
  OAI211_X1 U17924 ( .C1(n14546), .C2(n15896), .A(n14545), .B(n14544), .ZN(
        P1_U2888) );
  AOI21_X1 U17925 ( .B1(n14547), .B2(n14276), .A(n10243), .ZN(n15935) );
  INV_X1 U17926 ( .A(n15935), .ZN(n14552) );
  OAI222_X1 U17927 ( .A1(n15896), .A2(n14552), .B1(n14551), .B2(n14550), .C1(
        n14549), .C2(n14548), .ZN(P1_U2889) );
  INV_X1 U17928 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20910) );
  NOR2_X1 U17929 ( .A1(n20055), .A2(n20910), .ZN(n14720) );
  NOR2_X1 U17930 ( .A1(n15960), .A2(n14553), .ZN(n14554) );
  AOI211_X1 U17931 ( .C1(n15942), .C2(n14555), .A(n14720), .B(n14554), .ZN(
        n14560) );
  NAND2_X1 U17932 ( .A1(n14557), .A2(n14556), .ZN(n14558) );
  XOR2_X1 U17933 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n14558), .Z(
        n14719) );
  NAND2_X1 U17934 ( .A1(n14719), .A2(n20013), .ZN(n14559) );
  OAI211_X1 U17935 ( .C1(n14561), .C2(n15953), .A(n14560), .B(n14559), .ZN(
        P1_U2969) );
  MUX2_X1 U17936 ( .A(n11856), .B(n14563), .S(n14562), .Z(n14564) );
  XNOR2_X1 U17937 ( .A(n14564), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14735) );
  OR2_X1 U17938 ( .A1(n20055), .A2(n20908), .ZN(n14729) );
  NAND2_X1 U17939 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14565) );
  OAI211_X1 U17940 ( .C1(n15954), .C2(n14566), .A(n14729), .B(n14565), .ZN(
        n14567) );
  AOI21_X1 U17941 ( .B1(n14568), .B2(n20166), .A(n14567), .ZN(n14569) );
  OAI21_X1 U17942 ( .B1(n15955), .B2(n14735), .A(n14569), .ZN(P1_U2970) );
  OAI21_X1 U17943 ( .B1(n15918), .B2(n14703), .A(n14622), .ZN(n14573) );
  INV_X1 U17944 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14696) );
  INV_X1 U17945 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15994) );
  NAND4_X1 U17946 ( .A1(n14696), .A2(n15985), .A3(n15994), .A4(n14594), .ZN(
        n14570) );
  NAND2_X1 U17947 ( .A1(n14573), .A2(n14570), .ZN(n14572) );
  INV_X1 U17948 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14753) );
  MUX2_X1 U17949 ( .A(n14753), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15908), .Z(n14571) );
  OAI211_X1 U17950 ( .C1(n14573), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14572), .B(n14571), .ZN(n14574) );
  XNOR2_X1 U17951 ( .A(n14574), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14736) );
  INV_X1 U17952 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14577) );
  NAND2_X1 U17953 ( .A1(n15942), .A2(n14575), .ZN(n14576) );
  NAND2_X1 U17954 ( .A1(n20070), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14738) );
  OAI211_X1 U17955 ( .C1(n15960), .C2(n14577), .A(n14576), .B(n14738), .ZN(
        n14578) );
  AOI21_X1 U17956 ( .B1(n14736), .B2(n20013), .A(n14578), .ZN(n14579) );
  OAI21_X1 U17957 ( .B1(n14580), .B2(n15953), .A(n14579), .ZN(P1_U2971) );
  INV_X1 U17958 ( .A(n14581), .ZN(n14582) );
  AOI21_X1 U17959 ( .B1(n14583), .B2(n15918), .A(n14582), .ZN(n14584) );
  XNOR2_X1 U17960 ( .A(n14584), .B(n14753), .ZN(n14746) );
  NAND2_X1 U17961 ( .A1(n15942), .A2(n14585), .ZN(n14586) );
  NAND2_X1 U17962 ( .A1(n20070), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14747) );
  OAI211_X1 U17963 ( .C1(n15960), .C2(n14587), .A(n14586), .B(n14747), .ZN(
        n14588) );
  AOI21_X1 U17964 ( .B1(n14746), .B2(n20013), .A(n14588), .ZN(n14589) );
  OAI21_X1 U17965 ( .B1(n14590), .B2(n15953), .A(n14589), .ZN(P1_U2972) );
  NAND2_X1 U17966 ( .A1(n14622), .A2(n14703), .ZN(n14593) );
  NAND2_X1 U17967 ( .A1(n14600), .A2(n14591), .ZN(n14592) );
  MUX2_X1 U17968 ( .A(n14593), .B(n14592), .S(n15918), .Z(n14595) );
  XNOR2_X1 U17969 ( .A(n14595), .B(n14594), .ZN(n15971) );
  INV_X1 U17970 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U17971 ( .A1(n20070), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15963) );
  OAI21_X1 U17972 ( .B1(n15960), .B2(n14596), .A(n15963), .ZN(n14598) );
  MUX2_X1 U17973 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14600), .S(
        n15918), .Z(n14604) );
  NAND2_X1 U17974 ( .A1(n14601), .A2(n15908), .ZN(n14602) );
  NAND2_X1 U17975 ( .A1(n14602), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14616) );
  NAND2_X1 U17976 ( .A1(n14616), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14603) );
  NAND2_X1 U17977 ( .A1(n14604), .A2(n14603), .ZN(n14605) );
  XNOR2_X1 U17978 ( .A(n14605), .B(n14696), .ZN(n15978) );
  AOI22_X1 U17979 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n20070), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n14606) );
  OAI21_X1 U17980 ( .B1(n14607), .B2(n15954), .A(n14606), .ZN(n14608) );
  AOI21_X1 U17981 ( .B1(n14609), .B2(n20166), .A(n14608), .ZN(n14610) );
  OAI21_X1 U17982 ( .B1(n15955), .B2(n15978), .A(n14610), .ZN(P1_U2974) );
  INV_X1 U17983 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14611) );
  OAI22_X1 U17984 ( .A1(n15960), .A2(n14611), .B1(n20055), .B2(n21036), .ZN(
        n14612) );
  AOI21_X1 U17985 ( .B1(n15942), .B2(n14613), .A(n14612), .ZN(n14619) );
  INV_X1 U17986 ( .A(n14622), .ZN(n14614) );
  NAND2_X1 U17987 ( .A1(n14614), .A2(n14616), .ZN(n14615) );
  MUX2_X1 U17988 ( .A(n14616), .B(n14615), .S(n15918), .Z(n14617) );
  XNOR2_X1 U17989 ( .A(n14617), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15984) );
  NAND2_X1 U17990 ( .A1(n15984), .A2(n20013), .ZN(n14618) );
  OAI211_X1 U17991 ( .C1(n14620), .C2(n15953), .A(n14619), .B(n14618), .ZN(
        P1_U2975) );
  XNOR2_X1 U17992 ( .A(n15908), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14621) );
  XNOR2_X1 U17993 ( .A(n14622), .B(n14621), .ZN(n15989) );
  INV_X1 U17994 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21159) );
  NOR2_X1 U17995 ( .A1(n20055), .A2(n21159), .ZN(n15991) );
  INV_X1 U17996 ( .A(n15991), .ZN(n14624) );
  NAND2_X1 U17997 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14623) );
  OAI211_X1 U17998 ( .C1(n15954), .C2(n14625), .A(n14624), .B(n14623), .ZN(
        n14626) );
  AOI21_X1 U17999 ( .B1(n14627), .B2(n20166), .A(n14626), .ZN(n14628) );
  OAI21_X1 U18000 ( .B1(n15989), .B2(n15955), .A(n14628), .ZN(P1_U2976) );
  NAND2_X1 U18001 ( .A1(n14630), .A2(n14629), .ZN(n14631) );
  XOR2_X1 U18002 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14631), .Z(
        n16004) );
  OAI22_X1 U18003 ( .A1(n15960), .A2(n14633), .B1(n20055), .B2(n14632), .ZN(
        n14636) );
  NOR2_X1 U18004 ( .A1(n14634), .A2(n15953), .ZN(n14635) );
  AOI211_X1 U18005 ( .C1(n15942), .C2(n14637), .A(n14636), .B(n14635), .ZN(
        n14638) );
  OAI21_X1 U18006 ( .B1(n15955), .B2(n16004), .A(n14638), .ZN(P1_U2977) );
  NOR2_X1 U18007 ( .A1(n16006), .A2(n15909), .ZN(n14641) );
  INV_X1 U18008 ( .A(n14639), .ZN(n14640) );
  MUX2_X1 U18009 ( .A(n14641), .B(n14640), .S(n15918), .Z(n14642) );
  XOR2_X1 U18010 ( .A(n14642), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n14764) );
  AOI22_X1 U18011 ( .A1(n20013), .A2(n14764), .B1(n20070), .B2(
        P1_REIP_REG_20__SCAN_IN), .ZN(n14643) );
  OAI21_X1 U18012 ( .B1(n15960), .B2(n15786), .A(n14643), .ZN(n14644) );
  AOI21_X1 U18013 ( .B1(n15942), .B2(n15776), .A(n14644), .ZN(n14645) );
  OAI21_X1 U18014 ( .B1(n15780), .B2(n15953), .A(n14645), .ZN(P1_U2979) );
  NAND2_X1 U18015 ( .A1(n20070), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14776) );
  OAI21_X1 U18016 ( .B1(n15960), .B2(n15800), .A(n14776), .ZN(n14649) );
  NOR2_X1 U18017 ( .A1(n14647), .A2(n14646), .ZN(n14772) );
  INV_X1 U18018 ( .A(n15909), .ZN(n14773) );
  NOR3_X1 U18019 ( .A1(n14772), .A2(n14773), .A3(n15955), .ZN(n14648) );
  AOI211_X1 U18020 ( .C1(n15942), .C2(n15805), .A(n14649), .B(n14648), .ZN(
        n14650) );
  OAI21_X1 U18021 ( .B1(n15802), .B2(n15953), .A(n14650), .ZN(P1_U2981) );
  NOR2_X1 U18022 ( .A1(n14652), .A2(n14651), .ZN(n15929) );
  OAI21_X1 U18023 ( .B1(n15929), .B2(n14653), .A(n15930), .ZN(n15917) );
  INV_X1 U18024 ( .A(n14654), .ZN(n15916) );
  XNOR2_X1 U18025 ( .A(n15917), .B(n15916), .ZN(n14789) );
  AOI22_X1 U18026 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20070), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14655) );
  OAI21_X1 U18027 ( .B1(n14656), .B2(n15954), .A(n14655), .ZN(n14657) );
  AOI21_X1 U18028 ( .B1(n14658), .B2(n20166), .A(n14657), .ZN(n14659) );
  OAI21_X1 U18029 ( .B1(n15955), .B2(n14789), .A(n14659), .ZN(P1_U2983) );
  NAND2_X1 U18030 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14660) );
  OAI211_X1 U18031 ( .C1(n15954), .C2(n14662), .A(n14661), .B(n14660), .ZN(
        n14663) );
  AOI21_X1 U18032 ( .B1(n14664), .B2(n20166), .A(n14663), .ZN(n14665) );
  OAI21_X1 U18033 ( .B1(n14666), .B2(n15955), .A(n14665), .ZN(P1_U2985) );
  AOI21_X1 U18034 ( .B1(n14669), .B2(n14668), .A(n14667), .ZN(n14670) );
  XOR2_X1 U18035 ( .A(n14671), .B(n14670), .Z(n14801) );
  INV_X1 U18036 ( .A(n15877), .ZN(n15839) );
  INV_X1 U18037 ( .A(n15838), .ZN(n14673) );
  OR2_X1 U18038 ( .A1(n20055), .A2(n21172), .ZN(n14796) );
  NAND2_X1 U18039 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14672) );
  OAI211_X1 U18040 ( .C1(n15954), .C2(n14673), .A(n14796), .B(n14672), .ZN(
        n14674) );
  AOI21_X1 U18041 ( .B1(n15839), .B2(n20166), .A(n14674), .ZN(n14675) );
  OAI21_X1 U18042 ( .B1(n14801), .B2(n15955), .A(n14675), .ZN(P1_U2986) );
  OAI21_X1 U18043 ( .B1(n15960), .B2(n14677), .A(n14676), .ZN(n14679) );
  NOR2_X1 U18044 ( .A1(n15852), .A2(n15953), .ZN(n14678) );
  AOI211_X1 U18045 ( .C1(n15942), .C2(n15849), .A(n14679), .B(n14678), .ZN(
        n14680) );
  OAI21_X1 U18046 ( .B1(n14681), .B2(n15955), .A(n14680), .ZN(P1_U2987) );
  NOR2_X1 U18047 ( .A1(n15938), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14683) );
  NOR2_X1 U18048 ( .A1(n14244), .A2(n15939), .ZN(n14682) );
  MUX2_X1 U18049 ( .A(n14683), .B(n14682), .S(n15908), .Z(n14684) );
  XOR2_X1 U18050 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n14684), .Z(
        n16033) );
  NAND2_X1 U18051 ( .A1(n16033), .A2(n20013), .ZN(n14688) );
  NOR2_X1 U18052 ( .A1(n20055), .A2(n21053), .ZN(n16031) );
  NOR2_X1 U18053 ( .A1(n15954), .A2(n14685), .ZN(n14686) );
  AOI211_X1 U18054 ( .C1(n15946), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16031), .B(n14686), .ZN(n14687) );
  OAI211_X1 U18055 ( .C1(n15953), .C2(n14689), .A(n14688), .B(n14687), .ZN(
        P1_U2988) );
  INV_X1 U18056 ( .A(n14690), .ZN(n14691) );
  NOR2_X1 U18057 ( .A1(n14760), .A2(n14691), .ZN(n15980) );
  AOI21_X1 U18058 ( .B1(n14693), .B2(n14692), .A(n15980), .ZN(n14774) );
  INV_X1 U18059 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14694) );
  INV_X1 U18060 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16014) );
  NAND2_X1 U18061 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16015) );
  NOR2_X1 U18062 ( .A1(n16014), .A2(n16015), .ZN(n14778) );
  NAND3_X1 U18063 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n14778), .ZN(n14756) );
  NOR4_X1 U18064 ( .A1(n14774), .A2(n14695), .A3(n14694), .A4(n14756), .ZN(
        n15992) );
  NAND3_X1 U18065 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n15992), .ZN(n15966) );
  NOR2_X1 U18066 ( .A1(n14696), .A2(n15966), .ZN(n15968) );
  NAND2_X1 U18067 ( .A1(n15968), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14737) );
  INV_X1 U18068 ( .A(n14737), .ZN(n14750) );
  NAND2_X1 U18069 ( .A1(n14750), .A2(n14710), .ZN(n14728) );
  INV_X1 U18070 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14713) );
  NOR4_X1 U18071 ( .A1(n14728), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14713), .A4(n14722), .ZN(n14697) );
  AOI211_X1 U18072 ( .C1(n14699), .C2(n16067), .A(n14698), .B(n14697), .ZN(
        n14717) );
  NAND2_X1 U18073 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15998) );
  AOI211_X1 U18074 ( .C1(n14771), .C2(n14756), .A(n14768), .B(n14767), .ZN(
        n16005) );
  NOR2_X1 U18075 ( .A1(n14771), .A2(n14700), .ZN(n16041) );
  AOI21_X1 U18076 ( .B1(n15732), .B2(n16005), .A(n16041), .ZN(n16000) );
  AOI21_X1 U18077 ( .B1(n14771), .B2(n15998), .A(n16000), .ZN(n15995) );
  OAI21_X1 U18078 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14757), .A(
        n15995), .ZN(n15979) );
  OAI22_X1 U18079 ( .A1(n14703), .A2(n14702), .B1(n14701), .B2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14704) );
  INV_X1 U18080 ( .A(n14704), .ZN(n14705) );
  OAI21_X1 U18081 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14706), .A(
        n14705), .ZN(n14707) );
  NOR2_X1 U18082 ( .A1(n15979), .A2(n14707), .ZN(n15973) );
  NAND2_X1 U18083 ( .A1(n15973), .A2(n14712), .ZN(n14715) );
  NAND2_X1 U18084 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15973), .ZN(
        n15967) );
  INV_X1 U18085 ( .A(n15967), .ZN(n14708) );
  NAND2_X1 U18086 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n14708), .ZN(
        n14709) );
  NAND2_X1 U18087 ( .A1(n14715), .A2(n14709), .ZN(n14754) );
  INV_X1 U18088 ( .A(n14710), .ZN(n14741) );
  NAND2_X1 U18089 ( .A1(n14715), .A2(n14741), .ZN(n14711) );
  NAND2_X1 U18090 ( .A1(n14754), .A2(n14711), .ZN(n14733) );
  NOR2_X1 U18091 ( .A1(n14712), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14714) );
  NAND3_X1 U18092 ( .A1(n14723), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14715), .ZN(n14716) );
  OAI211_X1 U18093 ( .C1(n14718), .C2(n16052), .A(n14717), .B(n14716), .ZN(
        P1_U3000) );
  INV_X1 U18094 ( .A(n14719), .ZN(n14727) );
  AOI21_X1 U18095 ( .B1(n14721), .B2(n16067), .A(n14720), .ZN(n14726) );
  NOR2_X1 U18096 ( .A1(n14728), .A2(n14722), .ZN(n14724) );
  OAI21_X1 U18097 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14724), .A(
        n14723), .ZN(n14725) );
  OAI211_X1 U18098 ( .C1(n14727), .C2(n16052), .A(n14726), .B(n14725), .ZN(
        P1_U3001) );
  NOR2_X1 U18099 ( .A1(n14728), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14732) );
  OAI21_X1 U18100 ( .B1(n14730), .B2(n16046), .A(n14729), .ZN(n14731) );
  AOI211_X1 U18101 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14733), .A(
        n14732), .B(n14731), .ZN(n14734) );
  OAI21_X1 U18102 ( .B1(n14735), .B2(n16052), .A(n14734), .ZN(P1_U3002) );
  INV_X1 U18103 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14745) );
  NAND2_X1 U18104 ( .A1(n14736), .A2(n16068), .ZN(n14744) );
  AOI21_X1 U18105 ( .B1(n14745), .B2(n14753), .A(n14737), .ZN(n14742) );
  OAI21_X1 U18106 ( .B1(n14739), .B2(n16046), .A(n14738), .ZN(n14740) );
  AOI21_X1 U18107 ( .B1(n14742), .B2(n14741), .A(n14740), .ZN(n14743) );
  OAI211_X1 U18108 ( .C1(n14754), .C2(n14745), .A(n14744), .B(n14743), .ZN(
        P1_U3003) );
  NAND2_X1 U18109 ( .A1(n14746), .A2(n16068), .ZN(n14752) );
  OAI21_X1 U18110 ( .B1(n14748), .B2(n16046), .A(n14747), .ZN(n14749) );
  AOI21_X1 U18111 ( .B1(n14750), .B2(n14753), .A(n14749), .ZN(n14751) );
  OAI211_X1 U18112 ( .C1(n14754), .C2(n14753), .A(n14752), .B(n14751), .ZN(
        P1_U3004) );
  INV_X1 U18113 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14762) );
  INV_X1 U18114 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15778) );
  OAI22_X1 U18115 ( .A1(n16005), .A2(n14762), .B1(n20055), .B2(n15778), .ZN(
        n14755) );
  INV_X1 U18116 ( .A(n14755), .ZN(n14766) );
  INV_X1 U18117 ( .A(n14756), .ZN(n14761) );
  OAI22_X1 U18118 ( .A1(n14760), .A2(n14759), .B1(n14758), .B2(n14757), .ZN(
        n14795) );
  NAND3_X1 U18119 ( .A1(n14761), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n14795), .ZN(n16012) );
  AOI211_X1 U18120 ( .C1(n14762), .C2(n16006), .A(n15732), .B(n16012), .ZN(
        n14763) );
  AOI21_X1 U18121 ( .B1(n16068), .B2(n14764), .A(n14763), .ZN(n14765) );
  OAI211_X1 U18122 ( .C1(n15779), .C2(n16046), .A(n14766), .B(n14765), .ZN(
        P1_U3011) );
  INV_X1 U18123 ( .A(n14778), .ZN(n14770) );
  AOI211_X1 U18124 ( .C1(n14775), .C2(n14771), .A(n14768), .B(n14767), .ZN(
        n16024) );
  INV_X1 U18125 ( .A(n16024), .ZN(n14769) );
  AOI21_X1 U18126 ( .B1(n14771), .B2(n14770), .A(n14769), .ZN(n16013) );
  NOR2_X1 U18127 ( .A1(n14775), .A2(n14774), .ZN(n14783) );
  INV_X1 U18128 ( .A(n14783), .ZN(n16026) );
  NOR2_X1 U18129 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16026), .ZN(
        n14779) );
  OAI21_X1 U18130 ( .B1(n15801), .B2(n16046), .A(n14776), .ZN(n14777) );
  AOI21_X1 U18131 ( .B1(n14779), .B2(n14778), .A(n14777), .ZN(n14780) );
  OAI211_X1 U18132 ( .C1(n16013), .C2(n14782), .A(n14781), .B(n14780), .ZN(
        P1_U3013) );
  OAI211_X1 U18133 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n14783), .B(n16015), .ZN(
        n14788) );
  INV_X1 U18134 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14784) );
  INV_X1 U18135 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20931) );
  OAI22_X1 U18136 ( .A1(n16024), .A2(n14784), .B1(n20055), .B2(n20931), .ZN(
        n14785) );
  AOI21_X1 U18137 ( .B1(n16067), .B2(n14786), .A(n14785), .ZN(n14787) );
  OAI211_X1 U18138 ( .C1(n14789), .C2(n16052), .A(n14788), .B(n14787), .ZN(
        P1_U3015) );
  NAND2_X1 U18139 ( .A1(n14791), .A2(n14790), .ZN(n14792) );
  NAND2_X1 U18140 ( .A1(n14793), .A2(n14792), .ZN(n15875) );
  NAND2_X1 U18141 ( .A1(n14795), .A2(n14794), .ZN(n14797) );
  OAI211_X1 U18142 ( .C1(n16046), .C2(n15875), .A(n14797), .B(n14796), .ZN(
        n14798) );
  AOI21_X1 U18143 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14799), .A(
        n14798), .ZN(n14800) );
  OAI21_X1 U18144 ( .B1(n14801), .B2(n16052), .A(n14800), .ZN(P1_U3018) );
  NOR2_X1 U18145 ( .A1(n13763), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14804) );
  OAI22_X1 U18146 ( .A1(n20298), .A2(n14804), .B1(n20493), .B2(n14803), .ZN(
        n14805) );
  MUX2_X1 U18147 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14805), .S(
        n20156), .Z(P1_U3477) );
  NOR3_X1 U18148 ( .A1(n14806), .A2(n10920), .A3(n13393), .ZN(n14809) );
  NOR2_X1 U18149 ( .A1(n20493), .A2(n14807), .ZN(n14808) );
  AOI211_X1 U18150 ( .C1(n15675), .C2(n14810), .A(n14809), .B(n14808), .ZN(
        n15679) );
  NOR3_X1 U18151 ( .A1(n10920), .A2(n13393), .A3(n14811), .ZN(n14812) );
  AOI21_X1 U18152 ( .B1(n14814), .B2(n14813), .A(n14812), .ZN(n14815) );
  OAI21_X1 U18153 ( .B1(n15679), .B2(n14816), .A(n14815), .ZN(n14817) );
  MUX2_X1 U18154 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14817), .S(
        n16076), .Z(P1_U3473) );
  OAI22_X1 U18155 ( .A1(n14818), .A2(P2_STATEBS16_REG_SCAN_IN), .B1(n18906), 
        .B2(n19863), .ZN(n14819) );
  INV_X1 U18156 ( .A(n14819), .ZN(n14821) );
  OAI22_X1 U18157 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16369), .B1(n19869), 
        .B2(n19851), .ZN(n14820) );
  OAI21_X1 U18158 ( .B1(n14821), .B2(n12283), .A(n14820), .ZN(n14826) );
  AND2_X1 U18159 ( .A1(n14822), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16364) );
  OAI22_X1 U18160 ( .A1(n19869), .A2(n14823), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n16364), .ZN(n14824) );
  NOR2_X1 U18161 ( .A1(n18907), .A2(n14824), .ZN(n14825) );
  MUX2_X1 U18162 ( .A(n14826), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14825), 
        .Z(P2_U3610) );
  OAI211_X1 U18163 ( .C1(n14828), .C2(n15110), .A(n19094), .B(n14827), .ZN(
        n14838) );
  OR2_X1 U18164 ( .A1(n14910), .A2(n14829), .ZN(n14830) );
  NAND2_X1 U18165 ( .A1(n14895), .A2(n14830), .ZN(n15268) );
  INV_X1 U18166 ( .A(n15268), .ZN(n14836) );
  AOI22_X1 U18167 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19114), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19102), .ZN(n14831) );
  INV_X1 U18168 ( .A(n14831), .ZN(n14835) );
  NOR2_X1 U18169 ( .A1(n15019), .A2(n14832), .ZN(n14833) );
  OAI22_X1 U18170 ( .A1(n19087), .A2(n10893), .B1(n15264), .B2(n19085), .ZN(
        n14834) );
  AOI211_X1 U18171 ( .C1(n14836), .C2(n19081), .A(n14835), .B(n14834), .ZN(
        n14837) );
  OAI211_X1 U18172 ( .C1(n14839), .C2(n19105), .A(n14838), .B(n14837), .ZN(
        P2_U2827) );
  OAI211_X1 U18173 ( .C1(n14841), .C2(n15153), .A(n19094), .B(n14840), .ZN(
        n14851) );
  OR2_X1 U18174 ( .A1(n14944), .A2(n14843), .ZN(n14844) );
  NAND2_X1 U18175 ( .A1(n14842), .A2(n14844), .ZN(n15317) );
  INV_X1 U18176 ( .A(n15317), .ZN(n14849) );
  AOI22_X1 U18177 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19102), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19114), .ZN(n14845) );
  INV_X1 U18178 ( .A(n14845), .ZN(n14848) );
  AOI21_X1 U18179 ( .B1(n14846), .B2(n15046), .A(n9875), .ZN(n15314) );
  INV_X1 U18180 ( .A(n15314), .ZN(n15039) );
  OAI22_X1 U18181 ( .A1(n19087), .A2(n10134), .B1(n15039), .B2(n19085), .ZN(
        n14847) );
  AOI211_X1 U18182 ( .C1(n14849), .C2(n19081), .A(n14848), .B(n14847), .ZN(
        n14850) );
  OAI211_X1 U18183 ( .C1(n19105), .C2(n14852), .A(n14851), .B(n14850), .ZN(
        P2_U2831) );
  INV_X1 U18184 ( .A(n14853), .ZN(n14866) );
  NOR2_X1 U18185 ( .A1(n19092), .A2(n18969), .ZN(n14854) );
  XNOR2_X1 U18186 ( .A(n14854), .B(n16186), .ZN(n14855) );
  NAND2_X1 U18187 ( .A1(n14855), .A2(n19094), .ZN(n14865) );
  AOI21_X1 U18188 ( .B1(n14857), .B2(n9892), .A(n14856), .ZN(n16291) );
  INV_X1 U18189 ( .A(n16291), .ZN(n14859) );
  AOI22_X1 U18190 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19114), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19107), .ZN(n14858) );
  OAI211_X1 U18191 ( .C1(n19085), .C2(n14859), .A(n14858), .B(n19041), .ZN(
        n14863) );
  AND2_X1 U18192 ( .A1(n14987), .A2(n14860), .ZN(n14861) );
  OR2_X1 U18193 ( .A1(n14861), .A2(n14977), .ZN(n16181) );
  NOR2_X1 U18194 ( .A1(n16181), .A2(n19109), .ZN(n14862) );
  AOI211_X1 U18195 ( .C1(n19102), .C2(P2_REIP_REG_18__SCAN_IN), .A(n14863), 
        .B(n14862), .ZN(n14864) );
  OAI211_X1 U18196 ( .C1(n19105), .C2(n14866), .A(n14865), .B(n14864), .ZN(
        P2_U2837) );
  NOR2_X1 U18197 ( .A1(n19092), .A2(n19010), .ZN(n14867) );
  XNOR2_X1 U18198 ( .A(n14867), .B(n16214), .ZN(n14869) );
  NAND2_X1 U18199 ( .A1(n14869), .A2(n14868), .ZN(n14879) );
  INV_X1 U18200 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19902) );
  AOI22_X1 U18201 ( .A1(n14870), .A2(n19039), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19107), .ZN(n14871) );
  OAI211_X1 U18202 ( .C1(n19902), .C2(n19049), .A(n14871), .B(n19041), .ZN(
        n14872) );
  AOI21_X1 U18203 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19114), .A(
        n14872), .ZN(n14878) );
  INV_X1 U18204 ( .A(n16312), .ZN(n14876) );
  AOI21_X1 U18205 ( .B1(n14875), .B2(n14874), .A(n14873), .ZN(n19126) );
  AOI22_X1 U18206 ( .A1(n14876), .A2(n19081), .B1(n19101), .B2(n19126), .ZN(
        n14877) );
  NAND3_X1 U18207 ( .A1(n14879), .A2(n14878), .A3(n14877), .ZN(P2_U2841) );
  OAI21_X1 U18208 ( .B1(n19118), .B2(n14881), .A(n14880), .ZN(n15579) );
  NOR2_X1 U18209 ( .A1(n19105), .A2(n14882), .ZN(n14888) );
  AOI22_X1 U18210 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19114), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19102), .ZN(n14885) );
  NAND2_X1 U18211 ( .A1(n19113), .A2(n14883), .ZN(n14884) );
  OAI211_X1 U18212 ( .C1(n19085), .C2(n14886), .A(n14885), .B(n14884), .ZN(
        n14887) );
  AOI211_X1 U18213 ( .C1(n19107), .C2(P2_EBX_REG_1__SCAN_IN), .A(n14888), .B(
        n14887), .ZN(n14889) );
  OAI21_X1 U18214 ( .B1(n9970), .B2(n19109), .A(n14889), .ZN(n14890) );
  AOI21_X1 U18215 ( .B1(n19974), .B2(n19112), .A(n14890), .ZN(n14891) );
  OAI21_X1 U18216 ( .B1(n15579), .B2(n19048), .A(n14891), .ZN(P2_U2854) );
  INV_X1 U18217 ( .A(n16092), .ZN(n14892) );
  NAND2_X1 U18218 ( .A1(n14892), .A2(n14962), .ZN(n14893) );
  OAI21_X1 U18219 ( .B1(n14962), .B2(n16088), .A(n14893), .ZN(P2_U2856) );
  AND2_X1 U18220 ( .A1(n14895), .A2(n14894), .ZN(n14896) );
  INV_X1 U18221 ( .A(n14898), .ZN(n15003) );
  NAND2_X1 U18222 ( .A1(n14899), .A2(n14900), .ZN(n15002) );
  NAND3_X1 U18223 ( .A1(n15003), .A2(n14984), .A3(n15002), .ZN(n14902) );
  NAND2_X1 U18224 ( .A1(n14998), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14901) );
  OAI211_X1 U18225 ( .C1(n14980), .C2(n16099), .A(n14902), .B(n14901), .ZN(
        P2_U2858) );
  NAND2_X1 U18226 ( .A1(n12193), .A2(n14903), .ZN(n14905) );
  XNOR2_X1 U18227 ( .A(n14905), .B(n14904), .ZN(n15016) );
  NOR2_X1 U18228 ( .A1(n15268), .A2(n14980), .ZN(n14906) );
  AOI21_X1 U18229 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14980), .A(n14906), .ZN(
        n14907) );
  OAI21_X1 U18230 ( .B1(n15016), .B2(n15000), .A(n14907), .ZN(P2_U2859) );
  NOR2_X1 U18231 ( .A1(n14920), .A2(n14908), .ZN(n14909) );
  AOI21_X1 U18232 ( .B1(n14913), .B2(n14912), .A(n14911), .ZN(n15017) );
  NAND2_X1 U18233 ( .A1(n15017), .A2(n14984), .ZN(n14915) );
  NAND2_X1 U18234 ( .A1(n14980), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14914) );
  OAI211_X1 U18235 ( .C1(n14980), .C2(n16112), .A(n14915), .B(n14914), .ZN(
        P2_U2860) );
  OAI21_X1 U18236 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(n15032) );
  AND2_X1 U18237 ( .A1(n14929), .A2(n14919), .ZN(n14921) );
  OR2_X1 U18238 ( .A1(n14921), .A2(n14920), .ZN(n16123) );
  NOR2_X1 U18239 ( .A1(n16123), .A2(n14980), .ZN(n14922) );
  AOI21_X1 U18240 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n14980), .A(n14922), .ZN(
        n14923) );
  OAI21_X1 U18241 ( .B1(n15032), .B2(n15000), .A(n14923), .ZN(P2_U2861) );
  OAI21_X1 U18242 ( .B1(n14924), .B2(n14926), .A(n14925), .ZN(n15038) );
  NAND2_X1 U18243 ( .A1(n14842), .A2(n14927), .ZN(n14928) );
  NAND2_X1 U18244 ( .A1(n14929), .A2(n14928), .ZN(n16134) );
  MUX2_X1 U18245 ( .A(n16134), .B(n14930), .S(n14980), .Z(n14931) );
  OAI21_X1 U18246 ( .B1(n15038), .B2(n15000), .A(n14931), .ZN(P2_U2862) );
  AOI21_X1 U18247 ( .B1(n14932), .B2(n14934), .A(n14933), .ZN(n14935) );
  XOR2_X1 U18248 ( .A(n14936), .B(n14935), .Z(n15043) );
  NOR2_X1 U18249 ( .A1(n15317), .A2(n14980), .ZN(n14937) );
  AOI21_X1 U18250 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14980), .A(n14937), .ZN(
        n14938) );
  OAI21_X1 U18251 ( .B1(n15043), .B2(n15000), .A(n14938), .ZN(P2_U2863) );
  AOI21_X1 U18252 ( .B1(n14941), .B2(n14940), .A(n14939), .ZN(n14942) );
  INV_X1 U18253 ( .A(n14942), .ZN(n15052) );
  AND2_X1 U18254 ( .A1(n14949), .A2(n14943), .ZN(n14945) );
  OR2_X1 U18255 ( .A1(n14945), .A2(n14944), .ZN(n16146) );
  MUX2_X1 U18256 ( .A(n16146), .B(n10892), .S(n14980), .Z(n14946) );
  OAI21_X1 U18257 ( .B1(n15052), .B2(n15000), .A(n14946), .ZN(P2_U2864) );
  NAND2_X1 U18258 ( .A1(n14958), .A2(n14947), .ZN(n14948) );
  AND2_X1 U18259 ( .A1(n14949), .A2(n14948), .ZN(n16170) );
  INV_X1 U18260 ( .A(n16170), .ZN(n14955) );
  AND2_X1 U18261 ( .A1(n14950), .A2(n14951), .ZN(n14952) );
  NOR2_X1 U18262 ( .A1(n12085), .A2(n14952), .ZN(n16156) );
  NAND2_X1 U18263 ( .A1(n16156), .A2(n14984), .ZN(n14954) );
  NAND2_X1 U18264 ( .A1(n14980), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14953) );
  OAI211_X1 U18265 ( .C1(n14955), .C2(n14980), .A(n14954), .B(n14953), .ZN(
        P2_U2865) );
  INV_X1 U18266 ( .A(n14956), .ZN(n14970) );
  OAI21_X1 U18267 ( .B1(n14970), .B2(n9916), .A(n14950), .ZN(n15061) );
  INV_X1 U18268 ( .A(n14958), .ZN(n14959) );
  AOI21_X1 U18269 ( .B1(n14960), .B2(n14957), .A(n14959), .ZN(n18935) );
  NOR2_X1 U18270 ( .A1(n14962), .A2(n14961), .ZN(n14963) );
  AOI21_X1 U18271 ( .B1(n18935), .B2(n14962), .A(n14963), .ZN(n14964) );
  OAI21_X1 U18272 ( .B1(n15061), .B2(n15000), .A(n14964), .ZN(P2_U2866) );
  OR2_X1 U18273 ( .A1(n14965), .A2(n14966), .ZN(n14967) );
  NAND2_X1 U18274 ( .A1(n14957), .A2(n14967), .ZN(n18946) );
  INV_X1 U18275 ( .A(n14968), .ZN(n14971) );
  INV_X1 U18276 ( .A(n14969), .ZN(n14974) );
  AOI21_X1 U18277 ( .B1(n14971), .B2(n14974), .A(n14970), .ZN(n16160) );
  NAND2_X1 U18278 ( .A1(n16160), .A2(n14984), .ZN(n14973) );
  NAND2_X1 U18279 ( .A1(n14980), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14972) );
  OAI211_X1 U18280 ( .C1(n18946), .C2(n14980), .A(n14973), .B(n14972), .ZN(
        P2_U2867) );
  OAI21_X1 U18281 ( .B1(n9876), .B2(n14975), .A(n14974), .ZN(n15072) );
  NOR2_X1 U18282 ( .A1(n14977), .A2(n14976), .ZN(n14978) );
  OR2_X1 U18283 ( .A1(n14965), .A2(n14978), .ZN(n16282) );
  NOR2_X1 U18284 ( .A1(n16282), .A2(n14980), .ZN(n14979) );
  AOI21_X1 U18285 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n14980), .A(n14979), .ZN(
        n14981) );
  OAI21_X1 U18286 ( .B1(n15072), .B2(n15000), .A(n14981), .ZN(P2_U2868) );
  AND2_X1 U18287 ( .A1(n14200), .A2(n14982), .ZN(n14983) );
  NOR2_X1 U18288 ( .A1(n9876), .A2(n14983), .ZN(n16166) );
  NAND2_X1 U18289 ( .A1(n16166), .A2(n14984), .ZN(n14986) );
  NAND2_X1 U18290 ( .A1(n14998), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n14985) );
  OAI211_X1 U18291 ( .C1(n16181), .C2(n14998), .A(n14986), .B(n14985), .ZN(
        P2_U2869) );
  NAND2_X1 U18292 ( .A1(n14998), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14991) );
  INV_X1 U18293 ( .A(n14987), .ZN(n14988) );
  AOI21_X1 U18294 ( .B1(n14989), .B2(n14996), .A(n14988), .ZN(n18980) );
  NAND2_X1 U18295 ( .A1(n18980), .A2(n14962), .ZN(n14990) );
  OAI211_X1 U18296 ( .C1(n14992), .C2(n15000), .A(n14991), .B(n14990), .ZN(
        P2_U2870) );
  OR2_X1 U18297 ( .A1(n14994), .A2(n14993), .ZN(n14995) );
  NAND2_X1 U18298 ( .A1(n14996), .A2(n14995), .ZN(n18990) );
  NOR2_X1 U18299 ( .A1(n14980), .A2(n18990), .ZN(n14997) );
  AOI21_X1 U18300 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n14998), .A(n14997), .ZN(
        n14999) );
  OAI21_X1 U18301 ( .B1(n15001), .B2(n15000), .A(n14999), .ZN(P2_U2871) );
  NAND3_X1 U18302 ( .A1(n15003), .A2(n19181), .A3(n15002), .ZN(n15012) );
  OR2_X1 U18303 ( .A1(n15005), .A2(n15004), .ZN(n15006) );
  AOI22_X1 U18304 ( .A1(n19179), .A2(n16097), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n19178), .ZN(n15011) );
  AOI22_X1 U18305 ( .A1(n19121), .A2(BUF2_REG_29__SCAN_IN), .B1(n16165), .B2(
        n15008), .ZN(n15010) );
  NAND2_X1 U18306 ( .A1(n19120), .A2(BUF1_REG_29__SCAN_IN), .ZN(n15009) );
  NAND4_X1 U18307 ( .A1(n15012), .A2(n15011), .A3(n15010), .A4(n15009), .ZN(
        P2_U2890) );
  OAI22_X1 U18308 ( .A1(n15065), .A2(n15264), .B1(n19147), .B2(n13526), .ZN(
        n15013) );
  AOI21_X1 U18309 ( .B1(n19120), .B2(BUF1_REG_28__SCAN_IN), .A(n15013), .ZN(
        n15015) );
  AOI22_X1 U18310 ( .A1(n19121), .A2(BUF2_REG_28__SCAN_IN), .B1(n16165), .B2(
        n19131), .ZN(n15014) );
  OAI211_X1 U18311 ( .C1(n15016), .C2(n19174), .A(n15015), .B(n15014), .ZN(
        P2_U2891) );
  INV_X1 U18312 ( .A(n15017), .ZN(n15025) );
  AND2_X1 U18313 ( .A1(n9821), .A2(n15018), .ZN(n15020) );
  OR2_X1 U18314 ( .A1(n15020), .A2(n15019), .ZN(n16111) );
  OAI22_X1 U18315 ( .A1(n15065), .A2(n16111), .B1(n19147), .B2(n15021), .ZN(
        n15023) );
  OAI22_X1 U18316 ( .A1(n15068), .A2(n18253), .B1(n19134), .B2(n15066), .ZN(
        n15022) );
  AOI211_X1 U18317 ( .C1(n19120), .C2(BUF1_REG_27__SCAN_IN), .A(n15023), .B(
        n15022), .ZN(n15024) );
  OAI21_X1 U18318 ( .B1(n15025), .B2(n19174), .A(n15024), .ZN(P2_U2892) );
  NAND2_X1 U18319 ( .A1(n15027), .A2(n15026), .ZN(n15028) );
  AND2_X1 U18320 ( .A1(n9821), .A2(n15028), .ZN(n15292) );
  INV_X1 U18321 ( .A(n15292), .ZN(n16122) );
  OAI22_X1 U18322 ( .A1(n15065), .A2(n16122), .B1(n19147), .B2(n13530), .ZN(
        n15029) );
  AOI21_X1 U18323 ( .B1(n19120), .B2(BUF1_REG_26__SCAN_IN), .A(n15029), .ZN(
        n15031) );
  AOI22_X1 U18324 ( .A1(n19121), .A2(BUF2_REG_26__SCAN_IN), .B1(n16165), .B2(
        n19136), .ZN(n15030) );
  OAI211_X1 U18325 ( .C1(n15032), .C2(n19174), .A(n15031), .B(n15030), .ZN(
        P2_U2893) );
  XNOR2_X1 U18326 ( .A(n9875), .B(n15033), .ZN(n16133) );
  OAI22_X1 U18327 ( .A1(n15065), .A2(n16133), .B1(n19147), .B2(n15034), .ZN(
        n15035) );
  AOI21_X1 U18328 ( .B1(n19120), .B2(BUF1_REG_25__SCAN_IN), .A(n15035), .ZN(
        n15037) );
  AOI22_X1 U18329 ( .A1(n19121), .A2(BUF2_REG_25__SCAN_IN), .B1(n16165), .B2(
        n19139), .ZN(n15036) );
  OAI211_X1 U18330 ( .C1(n15038), .C2(n19174), .A(n15037), .B(n15036), .ZN(
        P2_U2894) );
  OAI22_X1 U18331 ( .A1(n15065), .A2(n15039), .B1(n19147), .B2(n13514), .ZN(
        n15040) );
  AOI21_X1 U18332 ( .B1(n19120), .B2(BUF1_REG_24__SCAN_IN), .A(n15040), .ZN(
        n15042) );
  AOI22_X1 U18333 ( .A1(n19121), .A2(BUF2_REG_24__SCAN_IN), .B1(n16165), .B2(
        n19142), .ZN(n15041) );
  OAI211_X1 U18334 ( .C1(n15043), .C2(n19174), .A(n15042), .B(n15041), .ZN(
        P2_U2895) );
  NAND2_X1 U18335 ( .A1(n15341), .A2(n15044), .ZN(n15045) );
  NAND2_X1 U18336 ( .A1(n15046), .A2(n15045), .ZN(n16154) );
  OAI22_X1 U18337 ( .A1(n15065), .A2(n16154), .B1(n19147), .B2(n15047), .ZN(
        n15050) );
  INV_X1 U18338 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15048) );
  OAI22_X1 U18339 ( .A1(n15068), .A2(n15048), .B1(n19294), .B2(n15066), .ZN(
        n15049) );
  AOI211_X1 U18340 ( .C1(n19120), .C2(BUF1_REG_23__SCAN_IN), .A(n15050), .B(
        n15049), .ZN(n15051) );
  OAI21_X1 U18341 ( .B1(n15052), .B2(n19174), .A(n15051), .ZN(P2_U2896) );
  OR2_X1 U18342 ( .A1(n15053), .A2(n15054), .ZN(n15056) );
  NAND2_X1 U18343 ( .A1(n15056), .A2(n15055), .ZN(n18944) );
  OAI22_X1 U18344 ( .A1(n15065), .A2(n18944), .B1(n19147), .B2(n15057), .ZN(
        n15058) );
  AOI21_X1 U18345 ( .B1(n19120), .B2(BUF1_REG_21__SCAN_IN), .A(n15058), .ZN(
        n15060) );
  AOI22_X1 U18346 ( .A1(n19121), .A2(BUF2_REG_21__SCAN_IN), .B1(n16165), .B2(
        n19150), .ZN(n15059) );
  OAI211_X1 U18347 ( .C1(n15061), .C2(n19174), .A(n15060), .B(n15059), .ZN(
        P2_U2898) );
  INV_X1 U18348 ( .A(n15062), .ZN(n15364) );
  OAI21_X1 U18349 ( .B1(n14856), .B2(n15063), .A(n15364), .ZN(n18968) );
  OAI22_X1 U18350 ( .A1(n15065), .A2(n18968), .B1(n19147), .B2(n15064), .ZN(
        n15070) );
  INV_X1 U18351 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15067) );
  OAI22_X1 U18352 ( .A1(n15068), .A2(n15067), .B1(n19171), .B2(n15066), .ZN(
        n15069) );
  AOI211_X1 U18353 ( .C1(n19120), .C2(BUF1_REG_19__SCAN_IN), .A(n15070), .B(
        n15069), .ZN(n15071) );
  OAI21_X1 U18354 ( .B1(n15072), .B2(n19174), .A(n15071), .ZN(P2_U2900) );
  INV_X1 U18355 ( .A(n15073), .ZN(n15077) );
  INV_X1 U18356 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15075) );
  OAI21_X1 U18357 ( .B1(n16275), .B2(n15075), .A(n15074), .ZN(n15076) );
  AOI21_X1 U18358 ( .B1(n16268), .B2(n15077), .A(n15076), .ZN(n15078) );
  OAI21_X1 U18359 ( .B1(n15079), .B2(n14106), .A(n15078), .ZN(n15080) );
  AOI21_X1 U18360 ( .B1(n15081), .B2(n19248), .A(n15080), .ZN(n15082) );
  OAI21_X1 U18361 ( .B1(n15083), .B2(n19237), .A(n15082), .ZN(P2_U2984) );
  NAND2_X1 U18362 ( .A1(n15085), .A2(n15084), .ZN(n15087) );
  XOR2_X1 U18363 ( .A(n15087), .B(n15086), .Z(n15260) );
  INV_X1 U18364 ( .A(n15088), .ZN(n15108) );
  AOI21_X1 U18365 ( .B1(n15251), .B2(n15108), .A(n15089), .ZN(n15258) );
  NAND2_X1 U18366 ( .A1(n19076), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15252) );
  OAI21_X1 U18367 ( .B1(n16275), .B2(n15090), .A(n15252), .ZN(n15091) );
  AOI21_X1 U18368 ( .B1(n16268), .B2(n15092), .A(n15091), .ZN(n15093) );
  OAI21_X1 U18369 ( .B1(n16099), .B2(n14106), .A(n15093), .ZN(n15094) );
  AOI21_X1 U18370 ( .B1(n15258), .B2(n19248), .A(n15094), .ZN(n15095) );
  OAI21_X1 U18371 ( .B1(n15260), .B2(n19237), .A(n15095), .ZN(P2_U2985) );
  NAND2_X1 U18372 ( .A1(n15102), .A2(n15100), .ZN(n15096) );
  AND2_X1 U18373 ( .A1(n15101), .A2(n15096), .ZN(n15099) );
  INV_X1 U18374 ( .A(n15097), .ZN(n15098) );
  INV_X1 U18375 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15122) );
  NOR2_X1 U18376 ( .A1(n15123), .A2(n15122), .ZN(n15121) );
  AOI21_X1 U18377 ( .B1(n15102), .B2(n15101), .A(n15100), .ZN(n15103) );
  XNOR2_X1 U18378 ( .A(n15104), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15105) );
  XNOR2_X1 U18379 ( .A(n15106), .B(n15105), .ZN(n15273) );
  AOI21_X1 U18380 ( .B1(n15109), .B2(n15107), .A(n15088), .ZN(n15271) );
  AND2_X1 U18381 ( .A1(n19076), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15265) );
  NOR2_X1 U18382 ( .A1(n19253), .A2(n15110), .ZN(n15111) );
  AOI211_X1 U18383 ( .C1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n19245), .A(
        n15265), .B(n15111), .ZN(n15112) );
  OAI21_X1 U18384 ( .B1(n15268), .B2(n14106), .A(n15112), .ZN(n15113) );
  AOI21_X1 U18385 ( .B1(n15271), .B2(n19248), .A(n15113), .ZN(n15114) );
  OAI21_X1 U18386 ( .B1(n15273), .B2(n19237), .A(n15114), .ZN(P2_U2986) );
  BUF_X1 U18387 ( .A(n15115), .Z(n15116) );
  OAI21_X1 U18388 ( .B1(n15116), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15107), .ZN(n15285) );
  NAND2_X1 U18389 ( .A1(n19076), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15274) );
  OAI21_X1 U18390 ( .B1(n16275), .B2(n15117), .A(n15274), .ZN(n15119) );
  NOR2_X1 U18391 ( .A1(n16112), .A2(n14106), .ZN(n15118) );
  AOI211_X1 U18392 ( .C1(n16268), .C2(n15120), .A(n15119), .B(n15118), .ZN(
        n15125) );
  INV_X1 U18393 ( .A(n15121), .ZN(n15282) );
  NAND2_X1 U18394 ( .A1(n15123), .A2(n15122), .ZN(n15281) );
  NAND3_X1 U18395 ( .A1(n15282), .A2(n19246), .A3(n15281), .ZN(n15124) );
  OAI211_X1 U18396 ( .C1(n15285), .C2(n16260), .A(n15125), .B(n15124), .ZN(
        P2_U2987) );
  NOR2_X1 U18397 ( .A1(n15126), .A2(n15138), .ZN(n15127) );
  XOR2_X1 U18398 ( .A(n15128), .B(n15127), .Z(n15298) );
  AOI21_X1 U18399 ( .B1(n15286), .B2(n15129), .A(n15116), .ZN(n15296) );
  INV_X1 U18400 ( .A(n16127), .ZN(n15131) );
  NAND2_X1 U18401 ( .A1(n19076), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15290) );
  OAI21_X1 U18402 ( .B1(n16275), .B2(n10058), .A(n15290), .ZN(n15130) );
  AOI21_X1 U18403 ( .B1(n16268), .B2(n15131), .A(n15130), .ZN(n15132) );
  OAI21_X1 U18404 ( .B1(n16123), .B2(n14106), .A(n15132), .ZN(n15133) );
  AOI21_X1 U18405 ( .B1(n15296), .B2(n19248), .A(n15133), .ZN(n15134) );
  OAI21_X1 U18406 ( .B1(n15298), .B2(n19237), .A(n15134), .ZN(P2_U2988) );
  INV_X1 U18407 ( .A(n15126), .ZN(n15139) );
  OAI21_X1 U18408 ( .B1(n15136), .B2(n15138), .A(n15135), .ZN(n15137) );
  OAI21_X1 U18409 ( .B1(n15139), .B2(n15138), .A(n15137), .ZN(n15310) );
  INV_X1 U18410 ( .A(n15129), .ZN(n15142) );
  AOI21_X1 U18411 ( .B1(n15303), .B2(n15141), .A(n15142), .ZN(n15299) );
  NAND2_X1 U18412 ( .A1(n15299), .A2(n19248), .ZN(n15148) );
  NAND2_X1 U18413 ( .A1(n19076), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15302) );
  OAI21_X1 U18414 ( .B1(n16275), .B2(n15143), .A(n15302), .ZN(n15145) );
  NOR2_X1 U18415 ( .A1(n16134), .A2(n14106), .ZN(n15144) );
  AOI211_X1 U18416 ( .C1(n16268), .C2(n15146), .A(n15145), .B(n15144), .ZN(
        n15147) );
  OAI211_X1 U18417 ( .C1(n19237), .C2(n15310), .A(n15148), .B(n15147), .ZN(
        P2_U2989) );
  XNOR2_X1 U18418 ( .A(n15150), .B(n15152), .ZN(n15321) );
  AOI21_X1 U18419 ( .B1(n15152), .B2(n15151), .A(n12662), .ZN(n15319) );
  AND2_X1 U18420 ( .A1(n19076), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15313) );
  AOI21_X1 U18421 ( .B1(n19245), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15313), .ZN(n15156) );
  INV_X1 U18422 ( .A(n15153), .ZN(n15154) );
  NAND2_X1 U18423 ( .A1(n16268), .A2(n15154), .ZN(n15155) );
  OAI211_X1 U18424 ( .C1(n15317), .C2(n14106), .A(n15156), .B(n15155), .ZN(
        n15157) );
  AOI21_X1 U18425 ( .B1(n15319), .B2(n19248), .A(n15157), .ZN(n15158) );
  OAI21_X1 U18426 ( .B1(n19237), .B2(n15321), .A(n15158), .ZN(P2_U2990) );
  OAI21_X1 U18427 ( .B1(n15159), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15151), .ZN(n15332) );
  XOR2_X1 U18428 ( .A(n15160), .B(n15161), .Z(n15330) );
  INV_X1 U18429 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19919) );
  OAI22_X1 U18430 ( .A1(n16275), .A2(n10045), .B1(n19919), .B2(n19041), .ZN(
        n15162) );
  AOI21_X1 U18431 ( .B1(n16268), .B2(n15163), .A(n15162), .ZN(n15164) );
  OAI21_X1 U18432 ( .B1(n16146), .B2(n14106), .A(n15164), .ZN(n15165) );
  AOI21_X1 U18433 ( .B1(n15330), .B2(n19246), .A(n15165), .ZN(n15166) );
  OAI21_X1 U18434 ( .B1(n15332), .B2(n16260), .A(n15166), .ZN(P2_U2991) );
  INV_X1 U18435 ( .A(n15436), .ZN(n15169) );
  INV_X1 U18436 ( .A(n15402), .ZN(n15171) );
  INV_X1 U18437 ( .A(n15394), .ZN(n15174) );
  INV_X1 U18438 ( .A(n15176), .ZN(n15177) );
  AOI21_X1 U18439 ( .B1(n15219), .B2(n15218), .A(n15177), .ZN(n16178) );
  INV_X1 U18440 ( .A(n15178), .ZN(n15195) );
  NAND2_X1 U18441 ( .A1(n15181), .A2(n15180), .ZN(n15182) );
  NAND2_X1 U18442 ( .A1(n15183), .A2(n16268), .ZN(n15184) );
  NAND2_X1 U18443 ( .A1(n19076), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15352) );
  OAI211_X1 U18444 ( .C1(n16275), .C2(n18932), .A(n15184), .B(n15352), .ZN(
        n15185) );
  AOI21_X1 U18445 ( .B1(n19255), .B2(n18935), .A(n15185), .ZN(n15191) );
  INV_X1 U18446 ( .A(n15187), .ZN(n15202) );
  AOI21_X1 U18447 ( .B1(n15189), .B2(n15202), .A(n10192), .ZN(n15358) );
  NAND2_X1 U18448 ( .A1(n15358), .A2(n19248), .ZN(n15190) );
  OAI211_X1 U18449 ( .C1(n15360), .C2(n19237), .A(n15191), .B(n15190), .ZN(
        P2_U2993) );
  INV_X1 U18450 ( .A(n15192), .ZN(n15194) );
  NOR2_X1 U18451 ( .A1(n15194), .A2(n15193), .ZN(n15198) );
  NOR2_X1 U18452 ( .A1(n15196), .A2(n15195), .ZN(n15197) );
  XNOR2_X1 U18453 ( .A(n15198), .B(n15197), .ZN(n15374) );
  INV_X1 U18454 ( .A(n18951), .ZN(n15205) );
  INV_X1 U18455 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15199) );
  NOR2_X1 U18456 ( .A1(n19041), .A2(n15199), .ZN(n15366) );
  AOI21_X1 U18457 ( .B1(n19245), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15366), .ZN(n15200) );
  OAI21_X1 U18458 ( .B1(n14106), .B2(n18946), .A(n15200), .ZN(n15204) );
  INV_X1 U18459 ( .A(n15201), .ZN(n15214) );
  OAI21_X1 U18460 ( .B1(n15214), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15202), .ZN(n15369) );
  NOR2_X1 U18461 ( .A1(n15369), .A2(n16260), .ZN(n15203) );
  AOI211_X1 U18462 ( .C1(n16268), .C2(n15205), .A(n15204), .B(n15203), .ZN(
        n15206) );
  OAI21_X1 U18463 ( .B1(n15374), .B2(n19237), .A(n15206), .ZN(P2_U2994) );
  NAND2_X1 U18464 ( .A1(n16178), .A2(n16175), .ZN(n16180) );
  NAND2_X1 U18465 ( .A1(n16180), .A2(n16176), .ZN(n15210) );
  NAND2_X1 U18466 ( .A1(n15208), .A2(n15207), .ZN(n15209) );
  XNOR2_X1 U18467 ( .A(n15210), .B(n15209), .ZN(n16286) );
  INV_X1 U18468 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19912) );
  OAI22_X1 U18469 ( .A1(n16275), .A2(n18957), .B1(n19912), .B2(n19041), .ZN(
        n15212) );
  NOR2_X1 U18470 ( .A1(n14106), .A2(n16282), .ZN(n15211) );
  AOI211_X1 U18471 ( .C1(n18963), .C2(n16268), .A(n15212), .B(n15211), .ZN(
        n15217) );
  INV_X1 U18472 ( .A(n15213), .ZN(n15215) );
  AOI21_X1 U18473 ( .B1(n16280), .B2(n15215), .A(n15214), .ZN(n16283) );
  NAND2_X1 U18474 ( .A1(n16283), .A2(n19248), .ZN(n15216) );
  OAI211_X1 U18475 ( .C1(n16286), .C2(n19237), .A(n15217), .B(n15216), .ZN(
        P2_U2995) );
  XNOR2_X1 U18476 ( .A(n15219), .B(n15218), .ZN(n15388) );
  INV_X1 U18477 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19908) );
  NOR2_X1 U18478 ( .A1(n19908), .A2(n19041), .ZN(n15222) );
  INV_X1 U18479 ( .A(n18971), .ZN(n18983) );
  OAI22_X1 U18480 ( .A1(n16275), .A2(n15220), .B1(n19253), .B2(n18983), .ZN(
        n15221) );
  AOI211_X1 U18481 ( .C1(n19255), .C2(n18980), .A(n15222), .B(n15221), .ZN(
        n15225) );
  NAND2_X1 U18482 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15382) );
  NOR2_X1 U18483 ( .A1(n15223), .A2(n15382), .ZN(n16191) );
  OAI211_X1 U18484 ( .C1(n16191), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19248), .B(n16182), .ZN(n15224) );
  OAI211_X1 U18485 ( .C1(n15388), .C2(n19237), .A(n15225), .B(n15224), .ZN(
        P2_U2997) );
  NAND2_X1 U18486 ( .A1(n15227), .A2(n15228), .ZN(n15399) );
  INV_X1 U18487 ( .A(n15399), .ZN(n15230) );
  AOI21_X1 U18488 ( .B1(n15228), .B2(n15398), .A(n15227), .ZN(n15229) );
  AOI21_X1 U18489 ( .B1(n15230), .B2(n15398), .A(n15229), .ZN(n15424) );
  INV_X1 U18490 ( .A(n19012), .ZN(n19024) );
  OAI22_X1 U18491 ( .A1(n16275), .A2(n15231), .B1(n19253), .B2(n19024), .ZN(
        n15238) );
  INV_X1 U18492 ( .A(n15414), .ZN(n15233) );
  AND2_X1 U18493 ( .A1(n15232), .A2(n15233), .ZN(n15449) );
  NAND2_X1 U18494 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15449), .ZN(
        n15426) );
  INV_X1 U18495 ( .A(n15449), .ZN(n15234) );
  NAND2_X1 U18496 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16304) );
  NOR2_X1 U18497 ( .A1(n15234), .A2(n16304), .ZN(n16210) );
  AOI21_X1 U18498 ( .B1(n15415), .B2(n15426), .A(n16210), .ZN(n15419) );
  AOI22_X1 U18499 ( .A1(n19248), .A2(n15419), .B1(n19076), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n15235) );
  OAI21_X1 U18500 ( .B1(n14106), .B2(n15236), .A(n15235), .ZN(n15237) );
  AOI211_X1 U18501 ( .C1(n15424), .C2(n19246), .A(n15238), .B(n15237), .ZN(
        n15239) );
  INV_X1 U18502 ( .A(n15239), .ZN(P2_U3001) );
  XNOR2_X1 U18503 ( .A(n15241), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15547) );
  XOR2_X1 U18504 ( .A(n15242), .B(n15243), .Z(n15545) );
  INV_X1 U18505 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19887) );
  OAI22_X1 U18506 ( .A1(n19887), .A2(n19041), .B1(n19253), .B2(n19066), .ZN(
        n15244) );
  AOI21_X1 U18507 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19245), .A(
        n15244), .ZN(n15245) );
  OAI21_X1 U18508 ( .B1(n19067), .B2(n14106), .A(n15245), .ZN(n15246) );
  AOI21_X1 U18509 ( .B1(n15545), .B2(n19246), .A(n15246), .ZN(n15247) );
  OAI21_X1 U18510 ( .B1(n15547), .B2(n16260), .A(n15247), .ZN(P2_U3008) );
  INV_X1 U18511 ( .A(n15261), .ZN(n15275) );
  NAND2_X1 U18512 ( .A1(n15248), .A2(n15275), .ZN(n15249) );
  NAND2_X1 U18513 ( .A1(n15250), .A2(n15249), .ZN(n15263) );
  NOR2_X1 U18514 ( .A1(n15263), .A2(n15251), .ZN(n15257) );
  OAI21_X1 U18515 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15253), .A(
        n15252), .ZN(n15254) );
  AOI21_X1 U18516 ( .B1(n16307), .B2(n16097), .A(n15254), .ZN(n15255) );
  OAI21_X1 U18517 ( .B1(n16099), .B2(n16313), .A(n15255), .ZN(n15256) );
  AOI211_X1 U18518 ( .C1(n15258), .C2(n16294), .A(n15257), .B(n15256), .ZN(
        n15259) );
  OAI21_X1 U18519 ( .B1(n15260), .B2(n16287), .A(n15259), .ZN(P2_U3017) );
  AOI21_X1 U18520 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15261), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15262) );
  NOR2_X1 U18521 ( .A1(n15263), .A2(n15262), .ZN(n15270) );
  INV_X1 U18522 ( .A(n15264), .ZN(n15266) );
  AOI21_X1 U18523 ( .B1(n16307), .B2(n15266), .A(n15265), .ZN(n15267) );
  OAI21_X1 U18524 ( .B1(n15268), .B2(n16313), .A(n15267), .ZN(n15269) );
  AOI211_X1 U18525 ( .C1(n15271), .C2(n16294), .A(n15270), .B(n15269), .ZN(
        n15272) );
  OAI21_X1 U18526 ( .B1(n15273), .B2(n16287), .A(n15272), .ZN(P2_U3018) );
  INV_X1 U18527 ( .A(n16111), .ZN(n15277) );
  OAI21_X1 U18528 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15275), .A(
        n15274), .ZN(n15276) );
  AOI21_X1 U18529 ( .B1(n16307), .B2(n15277), .A(n15276), .ZN(n15278) );
  OAI21_X1 U18530 ( .B1(n16112), .B2(n16313), .A(n15278), .ZN(n15279) );
  AOI21_X1 U18531 ( .B1(n15280), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15279), .ZN(n15284) );
  NAND3_X1 U18532 ( .A1(n15282), .A2(n16318), .A3(n15281), .ZN(n15283) );
  OAI211_X1 U18533 ( .C1(n15285), .C2(n16314), .A(n15284), .B(n15283), .ZN(
        P2_U3019) );
  NOR2_X1 U18534 ( .A1(n15304), .A2(n15286), .ZN(n15295) );
  INV_X1 U18535 ( .A(n15287), .ZN(n15300) );
  OAI211_X1 U18536 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15288), .B(n15300), .ZN(
        n15289) );
  NAND2_X1 U18537 ( .A1(n15290), .A2(n15289), .ZN(n15291) );
  AOI21_X1 U18538 ( .B1(n16307), .B2(n15292), .A(n15291), .ZN(n15293) );
  OAI21_X1 U18539 ( .B1(n16123), .B2(n16313), .A(n15293), .ZN(n15294) );
  AOI211_X1 U18540 ( .C1(n15296), .C2(n16294), .A(n15295), .B(n15294), .ZN(
        n15297) );
  OAI21_X1 U18541 ( .B1(n15298), .B2(n16287), .A(n15297), .ZN(P2_U3020) );
  NAND2_X1 U18542 ( .A1(n15299), .A2(n16294), .ZN(n15309) );
  INV_X1 U18543 ( .A(n16134), .ZN(n15307) );
  NAND2_X1 U18544 ( .A1(n15303), .A2(n15300), .ZN(n15301) );
  OAI211_X1 U18545 ( .C1(n16277), .C2(n16133), .A(n15302), .B(n15301), .ZN(
        n15306) );
  NOR2_X1 U18546 ( .A1(n15304), .A2(n15303), .ZN(n15305) );
  AOI211_X1 U18547 ( .C1(n15307), .C2(n16296), .A(n15306), .B(n15305), .ZN(
        n15308) );
  OAI211_X1 U18548 ( .C1(n15310), .C2(n16287), .A(n15309), .B(n15308), .ZN(
        P2_U3021) );
  OAI21_X1 U18549 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15312), .A(
        n15311), .ZN(n15316) );
  AOI21_X1 U18550 ( .B1(n16307), .B2(n15314), .A(n15313), .ZN(n15315) );
  OAI211_X1 U18551 ( .C1(n16313), .C2(n15317), .A(n15316), .B(n15315), .ZN(
        n15318) );
  AOI21_X1 U18552 ( .B1(n15319), .B2(n16294), .A(n15318), .ZN(n15320) );
  OAI21_X1 U18553 ( .B1(n16287), .B2(n15321), .A(n15320), .ZN(P2_U3022) );
  NAND2_X1 U18554 ( .A1(n15357), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15328) );
  INV_X1 U18555 ( .A(n16154), .ZN(n15326) );
  NOR2_X1 U18556 ( .A1(n19919), .A2(n19041), .ZN(n15325) );
  OAI21_X1 U18557 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15322), .ZN(n15323) );
  NOR2_X1 U18558 ( .A1(n15323), .A2(n15344), .ZN(n15324) );
  AOI211_X1 U18559 ( .C1(n16307), .C2(n15326), .A(n15325), .B(n15324), .ZN(
        n15327) );
  OAI211_X1 U18560 ( .C1(n16146), .C2(n16313), .A(n15328), .B(n15327), .ZN(
        n15329) );
  AOI21_X1 U18561 ( .B1(n15330), .B2(n16318), .A(n15329), .ZN(n15331) );
  OAI21_X1 U18562 ( .B1(n15332), .B2(n16314), .A(n15331), .ZN(P2_U3023) );
  NOR2_X1 U18563 ( .A1(n10192), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15333) );
  INV_X1 U18564 ( .A(n15357), .ZN(n15349) );
  INV_X1 U18565 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15348) );
  NAND2_X1 U18566 ( .A1(n15336), .A2(n15335), .ZN(n15337) );
  XNOR2_X1 U18567 ( .A(n15334), .B(n15337), .ZN(n16171) );
  NAND2_X1 U18568 ( .A1(n16171), .A2(n16318), .ZN(n15347) );
  OR2_X1 U18569 ( .A1(n15339), .A2(n15338), .ZN(n15340) );
  AND2_X1 U18570 ( .A1(n15341), .A2(n15340), .ZN(n16155) );
  NAND2_X1 U18571 ( .A1(n16307), .A2(n16155), .ZN(n15343) );
  NAND2_X1 U18572 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19076), .ZN(n15342) );
  OAI211_X1 U18573 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15344), .A(
        n15343), .B(n15342), .ZN(n15345) );
  AOI21_X1 U18574 ( .B1(n16170), .B2(n16296), .A(n15345), .ZN(n15346) );
  OAI211_X1 U18575 ( .C1(n15349), .C2(n15348), .A(n15347), .B(n15346), .ZN(
        n15350) );
  AOI21_X1 U18576 ( .B1(n10250), .B2(n16294), .A(n15350), .ZN(n15351) );
  INV_X1 U18577 ( .A(n15351), .ZN(P2_U3024) );
  NAND2_X1 U18578 ( .A1(n18935), .A2(n16296), .ZN(n15353) );
  OAI211_X1 U18579 ( .C1(n16277), .C2(n18944), .A(n15353), .B(n15352), .ZN(
        n15356) );
  INV_X1 U18580 ( .A(n15488), .ZN(n15379) );
  NOR3_X1 U18581 ( .A1(n15379), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15354), .ZN(n15355) );
  AOI211_X1 U18582 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15357), .A(
        n15356), .B(n15355), .ZN(n15359) );
  XNOR2_X1 U18583 ( .A(n16280), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15372) );
  INV_X1 U18584 ( .A(n15362), .ZN(n15361) );
  NOR2_X1 U18585 ( .A1(n15379), .A2(n15361), .ZN(n16281) );
  OAI21_X1 U18586 ( .B1(n16290), .B2(n15362), .A(n15453), .ZN(n16279) );
  NAND2_X1 U18587 ( .A1(n16279), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15368) );
  INV_X1 U18588 ( .A(n15363), .ZN(n15365) );
  AOI21_X1 U18589 ( .B1(n15365), .B2(n15364), .A(n15053), .ZN(n18947) );
  AOI21_X1 U18590 ( .B1(n16307), .B2(n18947), .A(n15366), .ZN(n15367) );
  OAI211_X1 U18591 ( .C1(n18946), .C2(n16313), .A(n15368), .B(n15367), .ZN(
        n15371) );
  NOR2_X1 U18592 ( .A1(n15369), .A2(n16314), .ZN(n15370) );
  AOI211_X1 U18593 ( .C1(n15372), .C2(n16281), .A(n15371), .B(n15370), .ZN(
        n15373) );
  OAI21_X1 U18594 ( .B1(n15374), .B2(n16287), .A(n15373), .ZN(P2_U3026) );
  INV_X1 U18595 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16193) );
  OAI21_X1 U18596 ( .B1(n15375), .B2(n16290), .A(n15453), .ZN(n16288) );
  AOI21_X1 U18597 ( .B1(n16314), .B2(n15376), .A(n16191), .ZN(n15377) );
  AOI211_X1 U18598 ( .C1(n15378), .C2(n16193), .A(n16288), .B(n15377), .ZN(
        n15397) );
  OAI211_X1 U18599 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16290), .A(
        n15397), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15386) );
  NOR2_X1 U18600 ( .A1(n12474), .A2(n15379), .ZN(n15475) );
  NAND2_X1 U18601 ( .A1(n15455), .A2(n15475), .ZN(n16310) );
  NOR2_X1 U18602 ( .A1(n16310), .A2(n16306), .ZN(n16298) );
  INV_X1 U18603 ( .A(n16298), .ZN(n15381) );
  NAND2_X1 U18604 ( .A1(n16191), .A2(n16294), .ZN(n15380) );
  OAI211_X1 U18605 ( .C1(n15382), .C2(n15381), .A(n15380), .B(n12538), .ZN(
        n15385) );
  AOI22_X1 U18606 ( .A1(n16296), .A2(n18980), .B1(P2_REIP_REG_17__SCAN_IN), 
        .B2(n19076), .ZN(n15383) );
  OAI21_X1 U18607 ( .B1(n18978), .B2(n16277), .A(n15383), .ZN(n15384) );
  AOI21_X1 U18608 ( .B1(n15386), .B2(n15385), .A(n15384), .ZN(n15387) );
  OAI21_X1 U18609 ( .B1(n15388), .B2(n16287), .A(n15387), .ZN(P2_U3029) );
  NAND2_X1 U18610 ( .A1(n19076), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16187) );
  OAI21_X1 U18611 ( .B1(n16313), .B2(n18990), .A(n16187), .ZN(n15392) );
  INV_X1 U18612 ( .A(n15223), .ZN(n15389) );
  AOI21_X1 U18613 ( .B1(n15389), .B2(n16294), .A(n16298), .ZN(n15390) );
  NOR3_X1 U18614 ( .A1(n15390), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16193), .ZN(n15391) );
  AOI211_X1 U18615 ( .C1(n16307), .C2(n15393), .A(n15392), .B(n15391), .ZN(
        n15396) );
  NAND2_X1 U18616 ( .A1(n16190), .A2(n16318), .ZN(n15395) );
  OAI211_X1 U18617 ( .C1(n15397), .C2(n16192), .A(n15396), .B(n15395), .ZN(
        P2_U3030) );
  NAND2_X1 U18618 ( .A1(n15399), .A2(n15398), .ZN(n16205) );
  NOR2_X1 U18619 ( .A1(n16205), .A2(n16206), .ZN(n16204) );
  INV_X1 U18620 ( .A(n15400), .ZN(n16208) );
  NOR2_X1 U18621 ( .A1(n16204), .A2(n16208), .ZN(n15404) );
  NOR2_X1 U18622 ( .A1(n15402), .A2(n15401), .ZN(n15403) );
  XNOR2_X1 U18623 ( .A(n15404), .B(n15403), .ZN(n16200) );
  XNOR2_X1 U18624 ( .A(n15223), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16198) );
  OR2_X1 U18625 ( .A1(n15405), .A2(n14873), .ZN(n15407) );
  NAND2_X1 U18626 ( .A1(n15407), .A2(n15406), .ZN(n19125) );
  INV_X1 U18627 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19904) );
  NOR2_X1 U18628 ( .A1(n19904), .A2(n19041), .ZN(n15408) );
  AOI221_X1 U18629 ( .B1(n16298), .B2(n16193), .C1(n16288), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n15408), .ZN(n15410) );
  NAND2_X1 U18630 ( .A1(n16296), .A2(n18995), .ZN(n15409) );
  OAI211_X1 U18631 ( .C1(n16277), .C2(n19125), .A(n15410), .B(n15409), .ZN(
        n15411) );
  AOI21_X1 U18632 ( .B1(n16198), .B2(n16294), .A(n15411), .ZN(n15412) );
  OAI21_X1 U18633 ( .B1(n16200), .B2(n16287), .A(n15412), .ZN(P2_U3031) );
  XOR2_X1 U18634 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n15430), .Z(
        n15416) );
  INV_X1 U18635 ( .A(n15453), .ZN(n15487) );
  AOI21_X1 U18636 ( .B1(n15414), .B2(n15413), .A(n15487), .ZN(n16322) );
  OAI22_X1 U18637 ( .A1(n16310), .A2(n15416), .B1(n15415), .B2(n16322), .ZN(
        n15423) );
  XNOR2_X1 U18638 ( .A(n15418), .B(n15417), .ZN(n19130) );
  AOI22_X1 U18639 ( .A1(n16296), .A2(n19020), .B1(n16294), .B2(n15419), .ZN(
        n15421) );
  NAND2_X1 U18640 ( .A1(n19076), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15420) );
  OAI211_X1 U18641 ( .C1(n19130), .C2(n16277), .A(n15421), .B(n15420), .ZN(
        n15422) );
  AOI211_X1 U18642 ( .C1(n15424), .C2(n16318), .A(n15423), .B(n15422), .ZN(
        n15425) );
  INV_X1 U18643 ( .A(n15425), .ZN(P2_U3033) );
  OR2_X1 U18644 ( .A1(n15449), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15427) );
  NAND2_X1 U18645 ( .A1(n15427), .A2(n15426), .ZN(n16219) );
  NOR2_X1 U18646 ( .A1(n16313), .A2(n15428), .ZN(n15432) );
  NAND2_X1 U18647 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19235), .ZN(n15429) );
  OAI221_X1 U18648 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16310), 
        .C1(n15430), .C2(n16322), .A(n15429), .ZN(n15431) );
  AOI211_X1 U18649 ( .C1(n16307), .C2(n15433), .A(n15432), .B(n15431), .ZN(
        n15440) );
  NAND2_X1 U18650 ( .A1(n15436), .A2(n15435), .ZN(n15437) );
  XNOR2_X1 U18651 ( .A(n15438), .B(n15437), .ZN(n16216) );
  NAND2_X1 U18652 ( .A1(n16216), .A2(n16318), .ZN(n15439) );
  OAI211_X1 U18653 ( .C1(n16219), .C2(n16314), .A(n15440), .B(n15439), .ZN(
        P2_U3034) );
  NAND2_X1 U18654 ( .A1(n15442), .A2(n15441), .ZN(n15484) );
  INV_X1 U18655 ( .A(n15482), .ZN(n15443) );
  NOR2_X1 U18656 ( .A1(n15484), .A2(n15443), .ZN(n15464) );
  AOI21_X1 U18657 ( .B1(n15464), .B2(n15466), .A(n15444), .ZN(n15448) );
  NAND2_X1 U18658 ( .A1(n15446), .A2(n15445), .ZN(n15447) );
  XNOR2_X1 U18659 ( .A(n15448), .B(n15447), .ZN(n16225) );
  AND2_X1 U18660 ( .A1(n15232), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15469) );
  NAND2_X1 U18661 ( .A1(n15469), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15470) );
  AOI21_X1 U18662 ( .B1(n15470), .B2(n15456), .A(n15449), .ZN(n16224) );
  OR2_X1 U18663 ( .A1(n15451), .A2(n15450), .ZN(n15452) );
  NAND2_X1 U18664 ( .A1(n15452), .A2(n14091), .ZN(n19135) );
  OAI21_X1 U18665 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16290), .A(
        n15453), .ZN(n15473) );
  INV_X1 U18666 ( .A(n15475), .ZN(n15454) );
  AOI211_X1 U18667 ( .C1(n15474), .C2(n15456), .A(n15455), .B(n15454), .ZN(
        n15458) );
  NOR2_X1 U18668 ( .A1(n10504), .A2(n19041), .ZN(n15457) );
  AOI211_X1 U18669 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15473), .A(
        n15458), .B(n15457), .ZN(n15460) );
  NAND2_X1 U18670 ( .A1(n19032), .A2(n16296), .ZN(n15459) );
  OAI211_X1 U18671 ( .C1(n16277), .C2(n19135), .A(n15460), .B(n15459), .ZN(
        n15461) );
  AOI21_X1 U18672 ( .B1(n16224), .B2(n16294), .A(n15461), .ZN(n15462) );
  OAI21_X1 U18673 ( .B1(n16225), .B2(n16287), .A(n15462), .ZN(P2_U3035) );
  INV_X1 U18674 ( .A(n15481), .ZN(n15463) );
  NOR2_X1 U18675 ( .A1(n15464), .A2(n15463), .ZN(n15468) );
  NAND2_X1 U18676 ( .A1(n15466), .A2(n15465), .ZN(n15467) );
  XNOR2_X1 U18677 ( .A(n15468), .B(n15467), .ZN(n16231) );
  INV_X1 U18678 ( .A(n15469), .ZN(n15485) );
  INV_X1 U18679 ( .A(n15470), .ZN(n15471) );
  AOI21_X1 U18680 ( .B1(n15474), .B2(n15485), .A(n15471), .ZN(n16233) );
  INV_X1 U18681 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19895) );
  NOR2_X1 U18682 ( .A1(n19895), .A2(n19041), .ZN(n15472) );
  AOI221_X1 U18683 ( .B1(n15475), .B2(n15474), .C1(n15473), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15472), .ZN(n15476) );
  INV_X1 U18684 ( .A(n15476), .ZN(n15479) );
  XNOR2_X1 U18685 ( .A(n15477), .B(n15491), .ZN(n19138) );
  OAI22_X1 U18686 ( .A1(n16277), .A2(n19138), .B1(n16313), .B2(n19043), .ZN(
        n15478) );
  AOI211_X1 U18687 ( .C1(n16233), .C2(n16294), .A(n15479), .B(n15478), .ZN(
        n15480) );
  OAI21_X1 U18688 ( .B1(n16231), .B2(n16287), .A(n15480), .ZN(P2_U3036) );
  NAND2_X1 U18689 ( .A1(n15482), .A2(n15481), .ZN(n15483) );
  XNOR2_X1 U18690 ( .A(n15484), .B(n15483), .ZN(n16236) );
  OAI21_X1 U18691 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15232), .A(
        n15485), .ZN(n16237) );
  INV_X1 U18692 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19893) );
  NOR2_X1 U18693 ( .A1(n19893), .A2(n19041), .ZN(n15486) );
  AOI221_X1 U18694 ( .B1(n15488), .B2(n12474), .C1(n15487), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15486), .ZN(n15495) );
  OR2_X1 U18695 ( .A1(n15490), .A2(n15489), .ZN(n15492) );
  NAND2_X1 U18696 ( .A1(n15492), .A2(n15491), .ZN(n19141) );
  INV_X1 U18697 ( .A(n19141), .ZN(n15493) );
  AOI22_X1 U18698 ( .A1(n16296), .A2(n19057), .B1(n16307), .B2(n15493), .ZN(
        n15494) );
  OAI211_X1 U18699 ( .C1(n16237), .C2(n16314), .A(n15495), .B(n15494), .ZN(
        n15496) );
  INV_X1 U18700 ( .A(n15496), .ZN(n15497) );
  OAI21_X1 U18701 ( .B1(n16287), .B2(n16236), .A(n15497), .ZN(P2_U3037) );
  NAND2_X1 U18702 ( .A1(n15498), .A2(n15520), .ZN(n15503) );
  INV_X1 U18703 ( .A(n15499), .ZN(n15500) );
  NOR2_X1 U18704 ( .A1(n15501), .A2(n15500), .ZN(n15502) );
  XNOR2_X1 U18705 ( .A(n15503), .B(n15502), .ZN(n16243) );
  INV_X1 U18706 ( .A(n16243), .ZN(n15514) );
  INV_X1 U18707 ( .A(n15505), .ZN(n15506) );
  XNOR2_X1 U18708 ( .A(n15504), .B(n15506), .ZN(n16242) );
  AOI21_X1 U18709 ( .B1(n15539), .B2(n15542), .A(n15533), .ZN(n15526) );
  OAI21_X1 U18710 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15507), .ZN(n15508) );
  OAI22_X1 U18711 ( .A1(n15526), .A2(n12481), .B1(n15528), .B2(n15508), .ZN(
        n15512) );
  AOI22_X1 U18712 ( .A1(n16307), .A2(n15509), .B1(n19076), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n15510) );
  OAI21_X1 U18713 ( .B1(n16313), .B2(n16246), .A(n15510), .ZN(n15511) );
  AOI211_X1 U18714 ( .C1(n16242), .C2(n16294), .A(n15512), .B(n15511), .ZN(
        n15513) );
  OAI21_X1 U18715 ( .B1(n16287), .B2(n15514), .A(n15513), .ZN(P2_U3038) );
  NAND2_X1 U18716 ( .A1(n15241), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15516) );
  NAND2_X1 U18717 ( .A1(n15516), .A2(n15515), .ZN(n15519) );
  XNOR2_X1 U18718 ( .A(n15517), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15518) );
  XNOR2_X1 U18719 ( .A(n15519), .B(n15518), .ZN(n16258) );
  INV_X1 U18720 ( .A(n15520), .ZN(n15524) );
  OAI21_X1 U18721 ( .B1(n15522), .B2(n15524), .A(n15521), .ZN(n15523) );
  OAI21_X1 U18722 ( .B1(n15498), .B2(n15524), .A(n15523), .ZN(n16255) );
  NAND2_X1 U18723 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19235), .ZN(n15525) );
  OAI221_X1 U18724 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15528), .C1(
        n15527), .C2(n15526), .A(n15525), .ZN(n15531) );
  OAI22_X1 U18725 ( .A1(n19145), .A2(n16277), .B1(n16313), .B2(n15529), .ZN(
        n15530) );
  AOI211_X1 U18726 ( .C1(n16255), .C2(n16318), .A(n15531), .B(n15530), .ZN(
        n15532) );
  OAI21_X1 U18727 ( .B1(n16314), .B2(n16258), .A(n15532), .ZN(P2_U3039) );
  INV_X1 U18728 ( .A(n15533), .ZN(n15543) );
  NAND3_X1 U18729 ( .A1(n14184), .A2(n9901), .A3(n15534), .ZN(n15535) );
  NAND2_X1 U18730 ( .A1(n15536), .A2(n15535), .ZN(n19148) );
  OAI22_X1 U18731 ( .A1(n19148), .A2(n16277), .B1(n19041), .B2(n19887), .ZN(
        n15537) );
  AOI21_X1 U18732 ( .B1(n16296), .B2(n15538), .A(n15537), .ZN(n15541) );
  NAND2_X1 U18733 ( .A1(n15539), .A2(n15542), .ZN(n15540) );
  OAI211_X1 U18734 ( .C1(n15543), .C2(n15542), .A(n15541), .B(n15540), .ZN(
        n15544) );
  AOI21_X1 U18735 ( .B1(n15545), .B2(n16318), .A(n15544), .ZN(n15546) );
  OAI21_X1 U18736 ( .B1(n15547), .B2(n16314), .A(n15546), .ZN(P2_U3040) );
  XNOR2_X1 U18737 ( .A(n15548), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15549) );
  XNOR2_X1 U18738 ( .A(n15550), .B(n15549), .ZN(n16272) );
  NAND2_X1 U18739 ( .A1(n16272), .A2(n16318), .ZN(n15559) );
  OAI22_X1 U18740 ( .A1(n16277), .A2(n19957), .B1(n19882), .B2(n19041), .ZN(
        n15551) );
  AOI21_X1 U18741 ( .B1(n13982), .B2(n16296), .A(n15551), .ZN(n15558) );
  OR2_X1 U18742 ( .A1(n12630), .A2(n15552), .ZN(n16269) );
  NAND3_X1 U18743 ( .A1(n16269), .A2(n16294), .A3(n15553), .ZN(n15557) );
  OAI21_X1 U18744 ( .B1(n15555), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n15554), .ZN(n15556) );
  NAND4_X1 U18745 ( .A1(n15559), .A2(n15558), .A3(n15557), .A4(n15556), .ZN(
        P2_U3043) );
  OAI22_X1 U18746 ( .A1(n13929), .A2(n15560), .B1(n19118), .B2(n19092), .ZN(
        n15577) );
  INV_X1 U18747 ( .A(n15593), .ZN(n15610) );
  NAND2_X1 U18748 ( .A1(n15561), .A2(n13076), .ZN(n15573) );
  MUX2_X1 U18749 ( .A(n15603), .B(n15573), .S(n15562), .Z(n15563) );
  AOI21_X1 U18750 ( .B1(n15564), .B2(n15610), .A(n15563), .ZN(n15565) );
  INV_X1 U18751 ( .A(n15565), .ZN(n16332) );
  INV_X1 U18752 ( .A(n15612), .ZN(n16370) );
  AOI22_X1 U18753 ( .A1(n16332), .A2(n19947), .B1(n15566), .B2(n16370), .ZN(
        n15567) );
  OAI21_X1 U18754 ( .B1(n15577), .B2(n19855), .A(n15567), .ZN(n15568) );
  MUX2_X1 U18755 ( .A(n15568), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15613), .Z(P2_U3601) );
  NAND2_X1 U18756 ( .A1(n15569), .A2(n15610), .ZN(n15576) );
  NOR2_X1 U18757 ( .A1(n15570), .A2(n15571), .ZN(n15572) );
  AOI22_X1 U18758 ( .A1(n15574), .A2(n15603), .B1(n15573), .B2(n15572), .ZN(
        n15575) );
  NAND2_X1 U18759 ( .A1(n15576), .A2(n15575), .ZN(n16326) );
  INV_X1 U18760 ( .A(n15577), .ZN(n15578) );
  NOR2_X1 U18761 ( .A1(n15578), .A2(n19855), .ZN(n15596) );
  OAI21_X1 U18762 ( .B1(n13929), .B2(n15580), .A(n15579), .ZN(n15595) );
  INV_X1 U18763 ( .A(n15595), .ZN(n15581) );
  AOI22_X1 U18764 ( .A1(n16326), .A2(n19947), .B1(n15596), .B2(n15581), .ZN(
        n15582) );
  OAI21_X1 U18765 ( .B1(n19971), .B2(n15612), .A(n15582), .ZN(n15583) );
  MUX2_X1 U18766 ( .A(n15583), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15613), .Z(P2_U3600) );
  OR2_X1 U18767 ( .A1(n16341), .A2(n16339), .ZN(n15605) );
  INV_X1 U18768 ( .A(n15571), .ZN(n15584) );
  NAND2_X1 U18769 ( .A1(n15584), .A2(n10202), .ZN(n15604) );
  NAND2_X1 U18770 ( .A1(n9807), .A2(n15604), .ZN(n15589) );
  NAND2_X1 U18771 ( .A1(n15603), .A2(n15585), .ZN(n15599) );
  INV_X1 U18772 ( .A(n15599), .ZN(n15586) );
  AOI22_X1 U18773 ( .A1(n15605), .A2(n15589), .B1(n15586), .B2(n9911), .ZN(
        n15592) );
  NAND2_X1 U18774 ( .A1(n15588), .A2(n15587), .ZN(n15601) );
  INV_X1 U18775 ( .A(n15589), .ZN(n15590) );
  NAND2_X1 U18776 ( .A1(n15601), .A2(n15590), .ZN(n15591) );
  OAI211_X1 U18777 ( .C1(n15594), .C2(n15593), .A(n15592), .B(n15591), .ZN(
        n16323) );
  AOI22_X1 U18778 ( .A1(n16323), .A2(n19947), .B1(n15596), .B2(n15595), .ZN(
        n15597) );
  OAI21_X1 U18779 ( .B1(n19961), .B2(n15612), .A(n15597), .ZN(n15598) );
  MUX2_X1 U18780 ( .A(n15598), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15613), .Z(P2_U3599) );
  NAND2_X1 U18781 ( .A1(n15599), .A2(n15604), .ZN(n15600) );
  AOI21_X1 U18782 ( .B1(n9807), .B2(n15601), .A(n15600), .ZN(n15607) );
  AOI22_X1 U18783 ( .A1(n15605), .A2(n15604), .B1(n10598), .B2(n15603), .ZN(
        n15606) );
  MUX2_X1 U18784 ( .A(n15607), .B(n15606), .S(n16325), .Z(n15608) );
  NAND2_X1 U18785 ( .A1(n15608), .A2(n9850), .ZN(n15609) );
  AOI21_X1 U18786 ( .B1(n13982), .B2(n15610), .A(n15609), .ZN(n16324) );
  OAI22_X1 U18787 ( .A1(n19521), .A2(n15612), .B1(n15611), .B2(n16324), .ZN(
        n15614) );
  MUX2_X1 U18788 ( .A(n15614), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15613), .Z(P2_U3596) );
  INV_X1 U18789 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U18790 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15626) );
  AOI22_X1 U18791 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15617) );
  AOI22_X1 U18792 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15616) );
  OAI211_X1 U18793 ( .C1(n17216), .C2(n17026), .A(n15617), .B(n15616), .ZN(
        n15624) );
  AOI22_X1 U18794 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15618), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15622) );
  AOI22_X1 U18795 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15621) );
  AOI22_X1 U18796 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15620) );
  NAND2_X1 U18797 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n15619) );
  NAND4_X1 U18798 ( .A1(n15622), .A2(n15621), .A3(n15620), .A4(n15619), .ZN(
        n15623) );
  AOI211_X1 U18799 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n15624), .B(n15623), .ZN(n15625) );
  OAI211_X1 U18800 ( .C1(n17218), .C2(n17028), .A(n15626), .B(n15625), .ZN(
        n17375) );
  INV_X1 U18801 ( .A(n17375), .ZN(n15631) );
  NAND2_X1 U18802 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .ZN(n17169) );
  NOR3_X1 U18803 ( .A1(n15627), .A2(n17169), .A3(n17172), .ZN(n15629) );
  OAI22_X1 U18804 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n15629), .B1(n17172), 
        .B2(n15628), .ZN(n15630) );
  AOI22_X1 U18805 ( .A1(n17275), .A2(n15631), .B1(n15630), .B2(n17266), .ZN(
        P3_U2690) );
  NAND2_X1 U18806 ( .A1(n18683), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18279) );
  NOR2_X1 U18807 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18888) );
  AOI21_X1 U18808 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18888), .ZN(n18734) );
  NOR2_X1 U18809 ( .A1(n18856), .A2(n18734), .ZN(n18237) );
  INV_X1 U18810 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16872) );
  OAI21_X1 U18811 ( .B1(n18697), .B2(n18839), .A(n16872), .ZN(n15649) );
  NOR2_X1 U18812 ( .A1(n17220), .A2(n15649), .ZN(n18226) );
  INV_X1 U18813 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16533) );
  NAND3_X1 U18814 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18831)
         );
  AOI21_X1 U18815 ( .B1(n18226), .B2(n16533), .A(n18831), .ZN(n15632) );
  NOR2_X1 U18816 ( .A1(n18532), .A2(n15632), .ZN(n18227) );
  INV_X1 U18817 ( .A(n18227), .ZN(n18233) );
  NAND2_X1 U18818 ( .A1(n18279), .A2(n18233), .ZN(n15635) );
  INV_X1 U18819 ( .A(n15635), .ZN(n15634) );
  INV_X1 U18820 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18718) );
  NAND3_X1 U18821 ( .A1(n18718), .A2(n18832), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18393) );
  NAND2_X1 U18822 ( .A1(n18718), .A2(n18832), .ZN(n16527) );
  AND2_X1 U18823 ( .A1(n18896), .A2(n16527), .ZN(n18877) );
  INV_X1 U18824 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18884) );
  NOR2_X1 U18825 ( .A1(n18842), .A2(n18884), .ZN(n17866) );
  OAI22_X1 U18826 ( .A1(n18877), .A2(n17866), .B1(n18683), .B2(n18832), .ZN(
        n15637) );
  NAND3_X1 U18827 ( .A1(n18684), .A2(n18233), .A3(n15637), .ZN(n15633) );
  OAI221_X1 U18828 ( .B1(n18684), .B2(n15634), .C1(n18684), .C2(n18393), .A(
        n15633), .ZN(P3_U2864) );
  NAND2_X1 U18829 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18416) );
  NOR2_X1 U18830 ( .A1(n18877), .A2(n17866), .ZN(n15636) );
  AOI221_X1 U18831 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18416), .C1(n15636), 
        .C2(n18416), .A(n15635), .ZN(n18232) );
  INV_X1 U18832 ( .A(n18393), .ZN(n18581) );
  OAI221_X1 U18833 ( .B1(n18581), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18581), .C2(n15637), .A(n18233), .ZN(n18230) );
  AOI22_X1 U18834 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18232), .B1(
        n18230), .B2(n18235), .ZN(P3_U2865) );
  NAND2_X1 U18835 ( .A1(n18829), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18236) );
  INV_X1 U18836 ( .A(n18236), .ZN(n15648) );
  NOR2_X1 U18837 ( .A1(n18880), .A2(n16529), .ZN(n15646) );
  NOR2_X1 U18838 ( .A1(n18244), .A2(n17474), .ZN(n18717) );
  NOR2_X1 U18839 ( .A1(n16549), .A2(n18717), .ZN(n15639) );
  INV_X1 U18840 ( .A(n15638), .ZN(n18883) );
  AOI21_X1 U18841 ( .B1(n18244), .B2(n16550), .A(n18698), .ZN(n15642) );
  NAND3_X1 U18842 ( .A1(n15644), .A2(n15762), .A3(n15643), .ZN(n15645) );
  OAI22_X1 U18843 ( .A1(n18703), .A2(n18715), .B1(n16533), .B2(n18831), .ZN(
        n15647) );
  INV_X1 U18844 ( .A(n18896), .ZN(n18858) );
  AND2_X1 U18845 ( .A1(n15649), .A2(n18698), .ZN(n18669) );
  NAND3_X1 U18846 ( .A1(n18860), .A2(n18858), .A3(n18669), .ZN(n15650) );
  OAI21_X1 U18847 ( .B1(n18860), .B2(n16872), .A(n15650), .ZN(P3_U3284) );
  NAND2_X1 U18848 ( .A1(n15652), .A2(n15651), .ZN(n15653) );
  XOR2_X1 U18849 ( .A(n15653), .B(n16406), .Z(n16422) );
  OAI21_X1 U18850 ( .B1(n16417), .B2(n18198), .A(n15654), .ZN(n15656) );
  NOR2_X1 U18851 ( .A1(n15655), .A2(n16418), .ZN(n16404) );
  AOI22_X1 U18852 ( .A1(n15657), .A2(n15656), .B1(n18137), .B2(n16404), .ZN(
        n15658) );
  NOR2_X1 U18853 ( .A1(n15658), .A2(n18222), .ZN(n15752) );
  INV_X1 U18854 ( .A(n15752), .ZN(n15664) );
  NOR2_X1 U18855 ( .A1(n16405), .A2(n18222), .ZN(n15659) );
  INV_X1 U18856 ( .A(n16395), .ZN(n16419) );
  AOI22_X1 U18857 ( .A1(n15659), .A2(n18137), .B1(n18218), .B2(n16419), .ZN(
        n15749) );
  INV_X1 U18858 ( .A(n15749), .ZN(n15662) );
  NOR2_X1 U18859 ( .A1(n18682), .A2(n18667), .ZN(n18073) );
  INV_X1 U18860 ( .A(n18073), .ZN(n18103) );
  AOI21_X1 U18861 ( .B1(n17923), .B2(n18103), .A(n15660), .ZN(n16431) );
  OAI22_X1 U18862 ( .A1(n18122), .A2(n16431), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18208), .ZN(n15661) );
  NOR2_X1 U18863 ( .A1(n15662), .A2(n15661), .ZN(n15663) );
  MUX2_X1 U18864 ( .A(n15664), .B(n15663), .S(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(n15665) );
  INV_X2 U18865 ( .A(n18221), .ZN(n18122) );
  NAND2_X1 U18866 ( .A1(n18122), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16411) );
  OAI211_X1 U18867 ( .C1(n16422), .C2(n18113), .A(n15665), .B(n16411), .ZN(
        P3_U2833) );
  AOI22_X1 U18868 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19114), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19102), .ZN(n15674) );
  INV_X1 U18869 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15666) );
  OAI22_X1 U18870 ( .A1(n15667), .A2(n19105), .B1(n19087), .B2(n15666), .ZN(
        n15668) );
  INV_X1 U18871 ( .A(n15668), .ZN(n15673) );
  AOI22_X1 U18872 ( .A1(n16170), .A2(n19081), .B1(n16155), .B2(n19101), .ZN(
        n15672) );
  OAI211_X1 U18873 ( .C1(n16174), .C2(n15670), .A(n19094), .B(n15669), .ZN(
        n15671) );
  NAND4_X1 U18874 ( .A1(n15674), .A2(n15673), .A3(n15672), .A4(n15671), .ZN(
        P2_U2833) );
  INV_X1 U18875 ( .A(n15707), .ZN(n15723) );
  INV_X1 U18876 ( .A(n15675), .ZN(n15678) );
  INV_X1 U18877 ( .A(n15676), .ZN(n15677) );
  OAI211_X1 U18878 ( .C1(n10911), .C2(n15678), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15677), .ZN(n15682) );
  INV_X1 U18879 ( .A(n15679), .ZN(n15681) );
  OAI211_X1 U18880 ( .C1(n20259), .C2(n15682), .A(n15681), .B(n15680), .ZN(
        n15684) );
  NAND2_X1 U18881 ( .A1(n20259), .A2(n15682), .ZN(n15683) );
  NAND2_X1 U18882 ( .A1(n15684), .A2(n15683), .ZN(n15685) );
  AND2_X1 U18883 ( .A1(n20573), .A2(n15685), .ZN(n15686) );
  OAI22_X1 U18884 ( .A1(n15687), .A2(n15686), .B1(n20573), .B2(n15685), .ZN(
        n15692) );
  NOR2_X1 U18885 ( .A1(n15689), .A2(n15688), .ZN(n15691) );
  INV_X1 U18886 ( .A(n15689), .ZN(n15690) );
  OAI22_X1 U18887 ( .A1(n15692), .A2(n15691), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15690), .ZN(n15718) );
  INV_X1 U18888 ( .A(n15693), .ZN(n15694) );
  NAND2_X1 U18889 ( .A1(n15704), .A2(n15694), .ZN(n15695) );
  NOR2_X1 U18890 ( .A1(n15696), .A2(n15695), .ZN(n15702) );
  INV_X1 U18891 ( .A(n15697), .ZN(n15698) );
  NAND2_X1 U18892 ( .A1(n13254), .A2(n15698), .ZN(n15701) );
  NAND2_X1 U18893 ( .A1(n15707), .A2(n15699), .ZN(n15700) );
  OAI211_X1 U18894 ( .C1(n15707), .C2(n15702), .A(n15701), .B(n15700), .ZN(
        n15703) );
  INV_X1 U18895 ( .A(n15703), .ZN(n20811) );
  NAND2_X1 U18896 ( .A1(n15705), .A2(n15704), .ZN(n15706) );
  OAI21_X1 U18897 ( .B1(n15707), .B2(n15708), .A(n15706), .ZN(n20006) );
  NOR2_X1 U18898 ( .A1(n15708), .A2(n20821), .ZN(n15710) );
  AOI21_X1 U18899 ( .B1(n15710), .B2(n15709), .A(n20814), .ZN(n15711) );
  OR2_X1 U18900 ( .A1(n20006), .A2(n15711), .ZN(n20012) );
  INV_X1 U18901 ( .A(n20012), .ZN(n15712) );
  OAI21_X1 U18902 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15712), .ZN(n15713) );
  NAND4_X1 U18903 ( .A1(n15715), .A2(n20811), .A3(n15714), .A4(n15713), .ZN(
        n15716) );
  AOI211_X1 U18904 ( .C1(n20157), .C2(n15718), .A(n15717), .B(n15716), .ZN(
        n15724) );
  NOR3_X1 U18905 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n15720), .A3(n15719), 
        .ZN(n15721) );
  AOI221_X1 U18906 ( .B1(n15722), .B2(n20735), .C1(n20820), .C2(n20735), .A(
        n15721), .ZN(n16080) );
  OAI221_X1 U18907 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15724), 
        .A(n16080), .ZN(n15725) );
  OAI21_X1 U18908 ( .B1(n15723), .B2(n15726), .A(n15725), .ZN(n15731) );
  INV_X1 U18909 ( .A(n15724), .ZN(n15728) );
  OAI211_X1 U18910 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20820), .A(n20736), 
        .B(n15726), .ZN(n16082) );
  AOI211_X1 U18911 ( .C1(n15729), .C2(n15728), .A(n15727), .B(n16082), .ZN(
        n15730) );
  AOI21_X1 U18912 ( .B1(n20169), .B2(n15731), .A(n15730), .ZN(P1_U3161) );
  INV_X1 U18913 ( .A(n15732), .ZN(n15740) );
  NOR2_X1 U18914 ( .A1(n15909), .A2(n15740), .ZN(n15733) );
  MUX2_X1 U18915 ( .A(n15734), .B(n15733), .S(n11856), .Z(n15735) );
  XOR2_X1 U18916 ( .A(n11853), .B(n15735), .Z(n15907) );
  AOI22_X1 U18917 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n16000), .B1(
        n20070), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15743) );
  NAND2_X1 U18918 ( .A1(n15737), .A2(n15736), .ZN(n15738) );
  NAND2_X1 U18919 ( .A1(n15739), .A2(n15738), .ZN(n15867) );
  INV_X1 U18920 ( .A(n15867), .ZN(n15741) );
  NOR2_X1 U18921 ( .A1(n16012), .A2(n15740), .ZN(n15999) );
  AOI22_X1 U18922 ( .A1(n15741), .A2(n16067), .B1(n15999), .B2(n11853), .ZN(
        n15742) );
  OAI211_X1 U18923 ( .C1(n15907), .C2(n16052), .A(n15743), .B(n15742), .ZN(
        P1_U3010) );
  NOR2_X1 U18924 ( .A1(n15745), .A2(n15744), .ZN(n15746) );
  XOR2_X1 U18925 ( .A(n15746), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16403) );
  NOR2_X1 U18926 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15747), .ZN(
        n16398) );
  AOI21_X1 U18927 ( .B1(n15750), .B2(n15749), .A(n15748), .ZN(n15751) );
  AOI21_X1 U18928 ( .B1(n15752), .B2(n16398), .A(n15751), .ZN(n15753) );
  NAND2_X1 U18929 ( .A1(n18122), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16391) );
  OAI211_X1 U18930 ( .C1(n16403), .C2(n18113), .A(n15753), .B(n16391), .ZN(
        P3_U2832) );
  INV_X1 U18931 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20748) );
  INV_X1 U18932 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21175) );
  NOR2_X1 U18933 ( .A1(n20003), .A2(n21175), .ZN(n15754) );
  INV_X1 U18934 ( .A(HOLD), .ZN(n20988) );
  NOR2_X1 U18935 ( .A1(n20748), .A2(n20988), .ZN(n20739) );
  INV_X1 U18936 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20749) );
  OAI22_X1 U18937 ( .A1(n15754), .A2(n20739), .B1(n20749), .B2(n20988), .ZN(
        n15755) );
  OAI211_X1 U18938 ( .C1(n20820), .C2(n20748), .A(n15756), .B(n15755), .ZN(
        P1_U3195) );
  AND2_X1 U18939 ( .A1(n15757), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U18940 ( .A(n16374), .ZN(n15759) );
  AOI221_X1 U18941 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16356), .C1(n18906), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(P2_STATE2_REG_2__SCAN_IN), .ZN(
        n19848) );
  NOR3_X1 U18942 ( .A1(n16369), .A2(n15759), .A3(n19848), .ZN(P2_U3178) );
  INV_X1 U18943 ( .A(n15758), .ZN(n19994) );
  AOI221_X1 U18944 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15759), .C1(n19994), .C2(
        n15759), .A(n19795), .ZN(n19988) );
  INV_X1 U18945 ( .A(n19988), .ZN(n19985) );
  NOR2_X1 U18946 ( .A1(n16334), .A2(n19985), .ZN(P2_U3047) );
  NAND3_X1 U18947 ( .A1(n16551), .A2(n18885), .A3(n15760), .ZN(n15761) );
  NAND2_X1 U18948 ( .A1(n17402), .A2(n17279), .ZN(n17326) );
  INV_X1 U18949 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17504) );
  INV_X1 U18950 ( .A(n18678), .ZN(n15763) );
  AOI22_X1 U18951 ( .A1(n17431), .A2(BUF2_REG_0__SCAN_IN), .B1(n17424), .B2(
        n15764), .ZN(n15765) );
  OAI221_X1 U18952 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17326), .C1(n17504), 
        .C2(n17279), .A(n15765), .ZN(P3_U2735) );
  NOR2_X1 U18953 ( .A1(n15767), .A2(n15766), .ZN(n15783) );
  AOI22_X1 U18954 ( .A1(n15901), .A2(n20075), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n15783), .ZN(n15775) );
  AOI22_X1 U18955 ( .A1(n20084), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20098), .ZN(n15774) );
  NOR2_X1 U18956 ( .A1(n14488), .A2(n15768), .ZN(n15769) );
  OR2_X1 U18957 ( .A1(n14433), .A2(n15769), .ZN(n15903) );
  OAI22_X1 U18958 ( .A1(n15903), .A2(n15851), .B1(n20073), .B2(n15867), .ZN(
        n15770) );
  INV_X1 U18959 ( .A(n15770), .ZN(n15773) );
  OR2_X1 U18960 ( .A1(n15771), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15772) );
  NAND4_X1 U18961 ( .A1(n15775), .A2(n15774), .A3(n15773), .A4(n15772), .ZN(
        P1_U2819) );
  AOI22_X1 U18962 ( .A1(n20084), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n20075), 
        .B2(n15776), .ZN(n15785) );
  NOR3_X1 U18963 ( .A1(n20931), .A2(n21138), .A3(n15777), .ZN(n15817) );
  NAND2_X1 U18964 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n15817), .ZN(n15807) );
  OAI21_X1 U18965 ( .B1(n15787), .B2(n15807), .A(n15778), .ZN(n15782) );
  OAI22_X1 U18966 ( .A1(n15780), .A2(n15851), .B1(n20073), .B2(n15779), .ZN(
        n15781) );
  AOI21_X1 U18967 ( .B1(n15783), .B2(n15782), .A(n15781), .ZN(n15784) );
  OAI211_X1 U18968 ( .C1(n15786), .C2(n15826), .A(n15785), .B(n15784), .ZN(
        P1_U2820) );
  OAI21_X1 U18969 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(P1_REIP_REG_19__SCAN_IN), 
        .A(n15787), .ZN(n15798) );
  AND2_X1 U18970 ( .A1(n15788), .A2(n20030), .ZN(n15816) );
  AOI22_X1 U18971 ( .A1(n15816), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_EBX_REG_19__SCAN_IN), .B2(n20084), .ZN(n15789) );
  OAI21_X1 U18972 ( .B1(n15915), .B2(n20109), .A(n15789), .ZN(n15790) );
  AOI211_X1 U18973 ( .C1(n20098), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20070), .B(n15790), .ZN(n15797) );
  AOI21_X1 U18974 ( .B1(n15792), .B2(n14495), .A(n14487), .ZN(n15912) );
  AOI21_X1 U18975 ( .B1(n15795), .B2(n15794), .A(n15793), .ZN(n16008) );
  AOI22_X1 U18976 ( .A1(n15912), .A2(n20048), .B1(n20096), .B2(n16008), .ZN(
        n15796) );
  OAI211_X1 U18977 ( .C1(n15807), .C2(n15798), .A(n15797), .B(n15796), .ZN(
        P1_U2821) );
  AOI22_X1 U18978 ( .A1(n15816), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n20084), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n15799) );
  OAI211_X1 U18979 ( .C1(n15826), .C2(n15800), .A(n15799), .B(n20055), .ZN(
        n15804) );
  OAI22_X1 U18980 ( .A1(n15802), .A2(n15851), .B1(n20073), .B2(n15801), .ZN(
        n15803) );
  AOI211_X1 U18981 ( .C1(n15805), .C2(n20075), .A(n15804), .B(n15803), .ZN(
        n15806) );
  OAI21_X1 U18982 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15807), .A(n15806), 
        .ZN(P1_U2822) );
  AOI22_X1 U18983 ( .A1(n20084), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20098), .ZN(n15821) );
  AOI21_X1 U18984 ( .B1(n20075), .B2(n15808), .A(n20070), .ZN(n15820) );
  AND2_X1 U18985 ( .A1(n14445), .A2(n15809), .ZN(n15810) );
  OR2_X1 U18986 ( .A1(n15810), .A2(n14493), .ZN(n15923) );
  NAND2_X1 U18987 ( .A1(n15812), .A2(n15811), .ZN(n15813) );
  NAND2_X1 U18988 ( .A1(n15814), .A2(n15813), .ZN(n16016) );
  OAI22_X1 U18989 ( .A1(n15923), .A2(n15851), .B1(n20073), .B2(n16016), .ZN(
        n15815) );
  INV_X1 U18990 ( .A(n15815), .ZN(n15819) );
  OAI21_X1 U18991 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15817), .A(n15816), 
        .ZN(n15818) );
  NAND4_X1 U18992 ( .A1(n15821), .A2(n15820), .A3(n15819), .A4(n15818), .ZN(
        P1_U2823) );
  AOI22_X1 U18993 ( .A1(n15935), .A2(n20048), .B1(n20075), .B2(n15934), .ZN(
        n15833) );
  AOI21_X1 U18994 ( .B1(n15824), .B2(n15823), .A(n15822), .ZN(n16028) );
  INV_X1 U18995 ( .A(n16028), .ZN(n15829) );
  OAI21_X1 U18996 ( .B1(n15826), .B2(n15825), .A(n20055), .ZN(n15827) );
  AOI21_X1 U18997 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(n20084), .A(n15827), .ZN(
        n15828) );
  OAI21_X1 U18998 ( .B1(n20073), .B2(n15829), .A(n15828), .ZN(n15831) );
  AOI211_X1 U18999 ( .C1(n10251), .C2(P1_REIP_REG_15__SCAN_IN), .A(n15831), 
        .B(n15830), .ZN(n15832) );
  NAND2_X1 U19000 ( .A1(n15833), .A2(n15832), .ZN(P1_U2825) );
  NAND2_X1 U19001 ( .A1(n20030), .A2(n15834), .ZN(n15856) );
  INV_X1 U19002 ( .A(n15875), .ZN(n15835) );
  AOI22_X1 U19003 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n20084), .B1(n20096), 
        .B2(n15835), .ZN(n15836) );
  OAI21_X1 U19004 ( .B1(n21172), .B2(n15856), .A(n15836), .ZN(n15837) );
  AOI211_X1 U19005 ( .C1(n20098), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20070), .B(n15837), .ZN(n15841) );
  AOI22_X1 U19006 ( .A1(n15839), .A2(n20048), .B1(n20075), .B2(n15838), .ZN(
        n15840) );
  OAI211_X1 U19007 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n15842), .A(n15841), 
        .B(n15840), .ZN(P1_U2827) );
  AOI21_X1 U19008 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15843), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15857) );
  INV_X1 U19009 ( .A(n15844), .ZN(n15845) );
  NAND2_X1 U19010 ( .A1(n20096), .A2(n15845), .ZN(n15848) );
  NAND2_X1 U19011 ( .A1(n20084), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n15847) );
  NAND2_X1 U19012 ( .A1(n20098), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15846) );
  AND4_X1 U19013 ( .A1(n15848), .A2(n15847), .A3(n20055), .A4(n15846), .ZN(
        n15855) );
  INV_X1 U19014 ( .A(n15849), .ZN(n15850) );
  OAI22_X1 U19015 ( .A1(n15852), .A2(n15851), .B1(n15850), .B2(n20109), .ZN(
        n15853) );
  INV_X1 U19016 ( .A(n15853), .ZN(n15854) );
  OAI211_X1 U19017 ( .C1(n15857), .C2(n15856), .A(n15855), .B(n15854), .ZN(
        P1_U2828) );
  INV_X1 U19018 ( .A(n15858), .ZN(n16045) );
  OAI22_X1 U19019 ( .A1(n15859), .A2(n20103), .B1(n20073), .B2(n16045), .ZN(
        n15860) );
  AOI211_X1 U19020 ( .C1(n20098), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20070), .B(n15860), .ZN(n15866) );
  INV_X1 U19021 ( .A(n15861), .ZN(n15943) );
  AOI22_X1 U19022 ( .A1(n15943), .A2(n20048), .B1(n20075), .B2(n15941), .ZN(
        n15865) );
  OAI21_X1 U19023 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n15863), .A(n15862), 
        .ZN(n15864) );
  NAND3_X1 U19024 ( .A1(n15866), .A2(n15865), .A3(n15864), .ZN(P1_U2830) );
  INV_X1 U19025 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n21026) );
  OAI22_X1 U19026 ( .A1(n15903), .A2(n14503), .B1(n15876), .B2(n15867), .ZN(
        n15868) );
  INV_X1 U19027 ( .A(n15868), .ZN(n15869) );
  OAI21_X1 U19028 ( .B1(n14492), .B2(n21026), .A(n15869), .ZN(P1_U2851) );
  INV_X1 U19029 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21186) );
  AOI22_X1 U19030 ( .A1(n15912), .A2(n20112), .B1(n20111), .B2(n16008), .ZN(
        n15870) );
  OAI21_X1 U19031 ( .B1(n14492), .B2(n21186), .A(n15870), .ZN(P1_U2853) );
  INV_X1 U19032 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15873) );
  OAI22_X1 U19033 ( .A1(n15923), .A2(n14503), .B1(n15876), .B2(n16016), .ZN(
        n15871) );
  INV_X1 U19034 ( .A(n15871), .ZN(n15872) );
  OAI21_X1 U19035 ( .B1(n14492), .B2(n15873), .A(n15872), .ZN(P1_U2855) );
  INV_X1 U19036 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n20905) );
  AOI22_X1 U19037 ( .A1(n15935), .A2(n20112), .B1(n20111), .B2(n16028), .ZN(
        n15874) );
  OAI21_X1 U19038 ( .B1(n14492), .B2(n20905), .A(n15874), .ZN(P1_U2857) );
  INV_X1 U19039 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15880) );
  OAI22_X1 U19040 ( .A1(n15877), .A2(n14503), .B1(n15876), .B2(n15875), .ZN(
        n15878) );
  INV_X1 U19041 ( .A(n15878), .ZN(n15879) );
  OAI21_X1 U19042 ( .B1(n14492), .B2(n15880), .A(n15879), .ZN(P1_U2859) );
  INV_X1 U19043 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20210) );
  AOI22_X1 U19044 ( .A1(n15893), .A2(n15881), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n15891), .ZN(n15885) );
  INV_X1 U19045 ( .A(n15887), .ZN(n15895) );
  INV_X1 U19046 ( .A(DATAI_21_), .ZN(n15882) );
  OAI22_X1 U19047 ( .A1(n15903), .A2(n15896), .B1(n15895), .B2(n15882), .ZN(
        n15883) );
  INV_X1 U19048 ( .A(n15883), .ZN(n15884) );
  OAI211_X1 U19049 ( .C1(n15900), .C2(n20210), .A(n15885), .B(n15884), .ZN(
        P1_U2883) );
  INV_X1 U19050 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20196) );
  AOI22_X1 U19051 ( .A1(n15893), .A2(n15886), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15891), .ZN(n15890) );
  AOI22_X1 U19052 ( .A1(n15912), .A2(n15888), .B1(n15887), .B2(DATAI_19_), 
        .ZN(n15889) );
  OAI211_X1 U19053 ( .C1(n15900), .C2(n20196), .A(n15890), .B(n15889), .ZN(
        P1_U2885) );
  INV_X1 U19054 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20184) );
  AOI22_X1 U19055 ( .A1(n15893), .A2(n15892), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n15891), .ZN(n15899) );
  INV_X1 U19056 ( .A(DATAI_17_), .ZN(n15894) );
  OAI22_X1 U19057 ( .A1(n15923), .A2(n15896), .B1(n15895), .B2(n15894), .ZN(
        n15897) );
  INV_X1 U19058 ( .A(n15897), .ZN(n15898) );
  OAI211_X1 U19059 ( .C1(n15900), .C2(n20184), .A(n15899), .B(n15898), .ZN(
        P1_U2887) );
  AOI22_X1 U19060 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20070), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15906) );
  INV_X1 U19061 ( .A(n15901), .ZN(n15902) );
  OAI22_X1 U19062 ( .A1(n15903), .A2(n15953), .B1(n15902), .B2(n15954), .ZN(
        n15904) );
  INV_X1 U19063 ( .A(n15904), .ZN(n15905) );
  OAI211_X1 U19064 ( .C1(n15907), .C2(n15955), .A(n15906), .B(n15905), .ZN(
        P1_U2978) );
  AOI22_X1 U19065 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20070), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15914) );
  NOR2_X1 U19066 ( .A1(n11856), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15910) );
  MUX2_X1 U19067 ( .A(n15908), .B(n15910), .S(n15909), .Z(n15911) );
  XNOR2_X1 U19068 ( .A(n15911), .B(n16006), .ZN(n16009) );
  AOI22_X1 U19069 ( .A1(n15912), .A2(n20166), .B1(n20013), .B2(n16009), .ZN(
        n15913) );
  OAI211_X1 U19070 ( .C1(n15954), .C2(n15915), .A(n15914), .B(n15913), .ZN(
        P1_U2980) );
  NOR2_X1 U19071 ( .A1(n15917), .A2(n15916), .ZN(n15920) );
  NOR2_X1 U19072 ( .A1(n15920), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15919) );
  MUX2_X1 U19073 ( .A(n15920), .B(n15919), .S(n15918), .Z(n15921) );
  XNOR2_X1 U19074 ( .A(n15921), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16022) );
  AOI22_X1 U19075 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20070), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15926) );
  OAI22_X1 U19076 ( .A1(n15923), .A2(n15953), .B1(n15922), .B2(n15954), .ZN(
        n15924) );
  INV_X1 U19077 ( .A(n15924), .ZN(n15925) );
  OAI211_X1 U19078 ( .C1(n15955), .C2(n16022), .A(n15926), .B(n15925), .ZN(
        P1_U2982) );
  INV_X1 U19079 ( .A(n15927), .ZN(n15928) );
  NOR2_X1 U19080 ( .A1(n15929), .A2(n15928), .ZN(n15933) );
  NAND2_X1 U19081 ( .A1(n15931), .A2(n15930), .ZN(n15932) );
  XNOR2_X1 U19082 ( .A(n15933), .B(n15932), .ZN(n16030) );
  AOI22_X1 U19083 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20070), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15937) );
  AOI22_X1 U19084 ( .A1(n15935), .A2(n20166), .B1(n15942), .B2(n15934), .ZN(
        n15936) );
  OAI211_X1 U19085 ( .C1(n16030), .C2(n15955), .A(n15937), .B(n15936), .ZN(
        P1_U2984) );
  MUX2_X1 U19086 ( .A(n15938), .B(n14244), .S(n15908), .Z(n15940) );
  XNOR2_X1 U19087 ( .A(n15940), .B(n15939), .ZN(n16053) );
  AOI22_X1 U19088 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20070), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n15945) );
  AOI22_X1 U19089 ( .A1(n15943), .A2(n20166), .B1(n15942), .B2(n15941), .ZN(
        n15944) );
  OAI211_X1 U19090 ( .C1(n15955), .C2(n16053), .A(n15945), .B(n15944), .ZN(
        P1_U2989) );
  AOI22_X1 U19091 ( .A1(n15946), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20070), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15952) );
  NAND2_X1 U19092 ( .A1(n15948), .A2(n15947), .ZN(n15949) );
  XNOR2_X1 U19093 ( .A(n15950), .B(n15949), .ZN(n16069) );
  AOI22_X1 U19094 ( .A1(n16069), .A2(n20013), .B1(n20166), .B2(n20113), .ZN(
        n15951) );
  OAI211_X1 U19095 ( .C1(n15954), .C2(n20033), .A(n15952), .B(n15951), .ZN(
        P1_U2992) );
  OAI222_X1 U19096 ( .A1(n15956), .A2(n15955), .B1(n15954), .B2(n20052), .C1(
        n15953), .C2(n20044), .ZN(n15957) );
  INV_X1 U19097 ( .A(n15957), .ZN(n15959) );
  OAI211_X1 U19098 ( .C1(n15961), .C2(n15960), .A(n15959), .B(n15958), .ZN(
        P1_U2993) );
  INV_X1 U19099 ( .A(n15962), .ZN(n15965) );
  INV_X1 U19100 ( .A(n15963), .ZN(n15964) );
  AOI21_X1 U19101 ( .B1(n15965), .B2(n16067), .A(n15964), .ZN(n15970) );
  NOR2_X1 U19102 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15966), .ZN(
        n15972) );
  OAI22_X1 U19103 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15968), .B1(
        n15972), .B2(n15967), .ZN(n15969) );
  OAI211_X1 U19104 ( .C1(n15971), .C2(n16052), .A(n15970), .B(n15969), .ZN(
        P1_U3005) );
  AOI21_X1 U19105 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n20070), .A(n15972), 
        .ZN(n15977) );
  INV_X1 U19106 ( .A(n15973), .ZN(n15975) );
  AOI22_X1 U19107 ( .A1(n15975), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n16067), .B2(n15974), .ZN(n15976) );
  OAI211_X1 U19108 ( .C1(n16052), .C2(n15978), .A(n15977), .B(n15976), .ZN(
        P1_U3006) );
  AOI21_X1 U19109 ( .B1(n15980), .B2(n15994), .A(n15979), .ZN(n15982) );
  OAI22_X1 U19110 ( .A1(n15982), .A2(n15985), .B1(n16046), .B2(n15981), .ZN(
        n15983) );
  AOI21_X1 U19111 ( .B1(n16068), .B2(n15984), .A(n15983), .ZN(n15987) );
  NAND3_X1 U19112 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n15992), .A3(
        n15985), .ZN(n15986) );
  OAI211_X1 U19113 ( .C1(n21036), .C2(n20055), .A(n15987), .B(n15986), .ZN(
        P1_U3007) );
  OAI22_X1 U19114 ( .A1(n15989), .A2(n16052), .B1(n16046), .B2(n15988), .ZN(
        n15990) );
  AOI211_X1 U19115 ( .C1(n15992), .C2(n15994), .A(n15991), .B(n15990), .ZN(
        n15993) );
  OAI21_X1 U19116 ( .B1(n15995), .B2(n15994), .A(n15993), .ZN(P1_U3008) );
  OAI22_X1 U19117 ( .A1(n15996), .A2(n16046), .B1(n14632), .B2(n20055), .ZN(
        n15997) );
  INV_X1 U19118 ( .A(n15997), .ZN(n16003) );
  AND2_X1 U19119 ( .A1(n15999), .A2(n15998), .ZN(n16001) );
  AOI222_X1 U19120 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16001), 
        .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16000), .C1(n16001), 
        .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16002) );
  OAI211_X1 U19121 ( .C1(n16004), .C2(n16052), .A(n16003), .B(n16002), .ZN(
        P1_U3009) );
  INV_X1 U19122 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21157) );
  OAI22_X1 U19123 ( .A1(n16006), .A2(n16005), .B1(n20055), .B2(n21157), .ZN(
        n16007) );
  INV_X1 U19124 ( .A(n16007), .ZN(n16011) );
  AOI22_X1 U19125 ( .A1(n16009), .A2(n16068), .B1(n16067), .B2(n16008), .ZN(
        n16010) );
  OAI211_X1 U19126 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16012), .A(
        n16011), .B(n16010), .ZN(P1_U3012) );
  INV_X1 U19127 ( .A(n16013), .ZN(n16019) );
  OAI21_X1 U19128 ( .B1(n16015), .B2(n16026), .A(n16014), .ZN(n16018) );
  INV_X1 U19129 ( .A(n16016), .ZN(n16017) );
  AOI22_X1 U19130 ( .A1(n16019), .A2(n16018), .B1(n16067), .B2(n16017), .ZN(
        n16021) );
  NAND2_X1 U19131 ( .A1(n20070), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16020) );
  OAI211_X1 U19132 ( .C1(n16022), .C2(n16052), .A(n16021), .B(n16020), .ZN(
        P1_U3014) );
  NAND2_X1 U19133 ( .A1(n20070), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16023) );
  OAI221_X1 U19134 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16026), 
        .C1(n16025), .C2(n16024), .A(n16023), .ZN(n16027) );
  AOI21_X1 U19135 ( .B1(n16028), .B2(n16067), .A(n16027), .ZN(n16029) );
  OAI21_X1 U19136 ( .B1(n16030), .B2(n16052), .A(n16029), .ZN(P1_U3016) );
  INV_X1 U19137 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16038) );
  AOI21_X1 U19138 ( .B1(n16067), .B2(n16032), .A(n16031), .ZN(n16037) );
  NOR2_X1 U19139 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16048), .ZN(
        n16034) );
  AOI22_X1 U19140 ( .A1(n16035), .A2(n16034), .B1(n16068), .B2(n16033), .ZN(
        n16036) );
  OAI211_X1 U19141 ( .C1(n16039), .C2(n16038), .A(n16037), .B(n16036), .ZN(
        P1_U3020) );
  NOR2_X1 U19142 ( .A1(n16049), .A2(n16040), .ZN(n16042) );
  AOI21_X1 U19143 ( .B1(n16043), .B2(n16042), .A(n16041), .ZN(n16054) );
  INV_X1 U19144 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n16044) );
  OAI22_X1 U19145 ( .A1(n16046), .A2(n16045), .B1(n16044), .B2(n20055), .ZN(
        n16047) );
  AOI21_X1 U19146 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16054), .A(
        n16047), .ZN(n16051) );
  NOR2_X1 U19147 ( .A1(n16049), .A2(n16048), .ZN(n16057) );
  OAI221_X1 U19148 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n15939), .C2(n11845), .A(
        n16057), .ZN(n16050) );
  OAI211_X1 U19149 ( .C1(n16053), .C2(n16052), .A(n16051), .B(n16050), .ZN(
        P1_U3021) );
  INV_X1 U19150 ( .A(n16054), .ZN(n16061) );
  AOI21_X1 U19151 ( .B1(n16067), .B2(n16056), .A(n16055), .ZN(n16060) );
  AOI22_X1 U19152 ( .A1(n16058), .A2(n16068), .B1(n11845), .B2(n16057), .ZN(
        n16059) );
  OAI211_X1 U19153 ( .C1(n11845), .C2(n16061), .A(n16060), .B(n16059), .ZN(
        P1_U3022) );
  INV_X1 U19154 ( .A(n16062), .ZN(n16074) );
  AND2_X1 U19155 ( .A1(n16064), .A2(n16063), .ZN(n16065) );
  NOR2_X1 U19156 ( .A1(n16066), .A2(n16065), .ZN(n20110) );
  AOI22_X1 U19157 ( .A1(n16067), .A2(n20110), .B1(n20070), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16072) );
  AOI22_X1 U19158 ( .A1(n16070), .A2(n16073), .B1(n16069), .B2(n16068), .ZN(
        n16071) );
  OAI211_X1 U19159 ( .C1(n16074), .C2(n16073), .A(n16072), .B(n16071), .ZN(
        P1_U3024) );
  NAND2_X1 U19160 ( .A1(n16075), .A2(n20798), .ZN(n16078) );
  OAI22_X1 U19161 ( .A1(n16079), .A2(n16078), .B1(n16077), .B2(n16076), .ZN(
        P1_U3468) );
  OAI221_X1 U19162 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20169), .C2(n20820), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20737) );
  AOI21_X1 U19163 ( .B1(n16084), .B2(n20737), .A(n16080), .ZN(n16081) );
  AOI21_X1 U19164 ( .B1(n16083), .B2(n16082), .A(n16081), .ZN(P1_U3162) );
  OAI22_X1 U19165 ( .A1(n20736), .A2(n20579), .B1(n20169), .B2(n16084), .ZN(
        P1_U3466) );
  NAND2_X1 U19166 ( .A1(n19094), .A2(n13929), .ZN(n19117) );
  INV_X1 U19167 ( .A(n16085), .ZN(n16090) );
  AOI22_X1 U19168 ( .A1(n19102), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19114), .ZN(n16086) );
  OAI21_X1 U19169 ( .B1(n16088), .B2(n16087), .A(n16086), .ZN(n16089) );
  AOI21_X1 U19170 ( .B1(n16090), .B2(n19039), .A(n16089), .ZN(n16091) );
  OAI21_X1 U19171 ( .B1(n16092), .B2(n19109), .A(n16091), .ZN(n16093) );
  AOI21_X1 U19172 ( .B1(n19101), .B2(n19119), .A(n16093), .ZN(n16094) );
  OAI21_X1 U19173 ( .B1(n19117), .B2(n16095), .A(n16094), .ZN(P2_U2824) );
  AOI22_X1 U19174 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19114), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19102), .ZN(n16107) );
  AOI22_X1 U19175 ( .A1(n16096), .A2(n19039), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n19107), .ZN(n16106) );
  INV_X1 U19176 ( .A(n16097), .ZN(n16098) );
  OAI22_X1 U19177 ( .A1(n16099), .A2(n19109), .B1(n16098), .B2(n19085), .ZN(
        n16100) );
  INV_X1 U19178 ( .A(n16100), .ZN(n16105) );
  OAI211_X1 U19179 ( .C1(n16103), .C2(n16102), .A(n19094), .B(n16101), .ZN(
        n16104) );
  NAND4_X1 U19180 ( .A1(n16107), .A2(n16106), .A3(n16105), .A4(n16104), .ZN(
        P2_U2826) );
  AOI22_X1 U19181 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n19102), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19114), .ZN(n16120) );
  INV_X1 U19182 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n16108) );
  OAI22_X1 U19183 ( .A1(n16109), .A2(n19105), .B1(n19087), .B2(n16108), .ZN(
        n16110) );
  INV_X1 U19184 ( .A(n16110), .ZN(n16119) );
  OAI22_X1 U19185 ( .A1(n16112), .A2(n19109), .B1(n16111), .B2(n19085), .ZN(
        n16113) );
  INV_X1 U19186 ( .A(n16113), .ZN(n16118) );
  OAI211_X1 U19187 ( .C1(n16116), .C2(n16115), .A(n19094), .B(n16114), .ZN(
        n16117) );
  NAND4_X1 U19188 ( .A1(n16120), .A2(n16119), .A3(n16118), .A4(n16117), .ZN(
        P2_U2828) );
  AOI22_X1 U19189 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19114), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19102), .ZN(n16131) );
  AOI22_X1 U19190 ( .A1(n16121), .A2(n19039), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n19107), .ZN(n16130) );
  OAI22_X1 U19191 ( .A1(n16123), .A2(n19109), .B1(n16122), .B2(n19085), .ZN(
        n16124) );
  INV_X1 U19192 ( .A(n16124), .ZN(n16129) );
  OAI211_X1 U19193 ( .C1(n16127), .C2(n16126), .A(n19094), .B(n16125), .ZN(
        n16128) );
  NAND4_X1 U19194 ( .A1(n16131), .A2(n16130), .A3(n16129), .A4(n16128), .ZN(
        P2_U2829) );
  AOI22_X1 U19195 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19114), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19102), .ZN(n16142) );
  AOI22_X1 U19196 ( .A1(n16132), .A2(n19039), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n19107), .ZN(n16141) );
  OAI22_X1 U19197 ( .A1(n16134), .A2(n19109), .B1(n16133), .B2(n19085), .ZN(
        n16135) );
  INV_X1 U19198 ( .A(n16135), .ZN(n16140) );
  OAI211_X1 U19199 ( .C1(n16138), .C2(n16137), .A(n19094), .B(n16136), .ZN(
        n16139) );
  NAND4_X1 U19200 ( .A1(n16142), .A2(n16141), .A3(n16140), .A4(n16139), .ZN(
        P2_U2830) );
  INV_X1 U19201 ( .A(n16143), .ZN(n16148) );
  OAI22_X1 U19202 ( .A1(n19919), .A2(n19049), .B1(n10045), .B2(n19072), .ZN(
        n16144) );
  AOI21_X1 U19203 ( .B1(n19107), .B2(P2_EBX_REG_23__SCAN_IN), .A(n16144), .ZN(
        n16145) );
  OAI21_X1 U19204 ( .B1(n16146), .B2(n19109), .A(n16145), .ZN(n16147) );
  AOI21_X1 U19205 ( .B1(n16148), .B2(n19039), .A(n16147), .ZN(n16153) );
  OAI211_X1 U19206 ( .C1(n16151), .C2(n16150), .A(n19094), .B(n16149), .ZN(
        n16152) );
  OAI211_X1 U19207 ( .C1(n19085), .C2(n16154), .A(n16153), .B(n16152), .ZN(
        P2_U2832) );
  AOI22_X1 U19208 ( .A1(n16165), .A2(n19146), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19178), .ZN(n16159) );
  AOI22_X1 U19209 ( .A1(n19120), .A2(BUF1_REG_22__SCAN_IN), .B1(n19121), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16158) );
  AOI22_X1 U19210 ( .A1(n16156), .A2(n19181), .B1(n19179), .B2(n16155), .ZN(
        n16157) );
  NAND3_X1 U19211 ( .A1(n16159), .A2(n16158), .A3(n16157), .ZN(P2_U2897) );
  AOI22_X1 U19212 ( .A1(n16165), .A2(n19157), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19178), .ZN(n16163) );
  AOI22_X1 U19213 ( .A1(n19120), .A2(BUF1_REG_20__SCAN_IN), .B1(n19121), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16162) );
  AOI22_X1 U19214 ( .A1(n16160), .A2(n19181), .B1(n19179), .B2(n18947), .ZN(
        n16161) );
  NAND3_X1 U19215 ( .A1(n16163), .A2(n16162), .A3(n16161), .ZN(P2_U2899) );
  AOI22_X1 U19216 ( .A1(n16165), .A2(n16164), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19178), .ZN(n16169) );
  AOI22_X1 U19217 ( .A1(n19120), .A2(BUF1_REG_18__SCAN_IN), .B1(n19121), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16168) );
  AOI22_X1 U19218 ( .A1(n16166), .A2(n19181), .B1(n19179), .B2(n16291), .ZN(
        n16167) );
  NAND3_X1 U19219 ( .A1(n16169), .A2(n16168), .A3(n16167), .ZN(P2_U2901) );
  AOI22_X1 U19220 ( .A1(n19245), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19235), .ZN(n16173) );
  AOI222_X1 U19221 ( .A1(n16171), .A2(n19246), .B1(n19255), .B2(n16170), .C1(
        n19248), .C2(n10250), .ZN(n16172) );
  OAI211_X1 U19222 ( .C1(n19253), .C2(n16174), .A(n16173), .B(n16172), .ZN(
        P2_U2992) );
  AOI22_X1 U19223 ( .A1(n19245), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19235), .ZN(n16185) );
  INV_X1 U19224 ( .A(n16176), .ZN(n16179) );
  AND2_X1 U19225 ( .A1(n16176), .A2(n16175), .ZN(n16177) );
  OAI22_X1 U19226 ( .A1(n16180), .A2(n16179), .B1(n16178), .B2(n16177), .ZN(
        n16297) );
  INV_X1 U19227 ( .A(n16181), .ZN(n16295) );
  AOI21_X1 U19228 ( .B1(n16183), .B2(n16182), .A(n15213), .ZN(n16293) );
  AOI222_X1 U19229 ( .A1(n16297), .A2(n19246), .B1(n19255), .B2(n16295), .C1(
        n19248), .C2(n16293), .ZN(n16184) );
  OAI211_X1 U19230 ( .C1(n19253), .C2(n16186), .A(n16185), .B(n16184), .ZN(
        P2_U2996) );
  NOR2_X1 U19231 ( .A1(n19253), .A2(n18988), .ZN(n16189) );
  OAI21_X1 U19232 ( .B1(n16275), .B2(n10048), .A(n16187), .ZN(n16188) );
  AOI211_X1 U19233 ( .C1(n16190), .C2(n19246), .A(n16189), .B(n16188), .ZN(
        n16197) );
  INV_X1 U19234 ( .A(n16191), .ZN(n16195) );
  OAI21_X1 U19235 ( .B1(n15223), .B2(n16193), .A(n16192), .ZN(n16194) );
  NAND3_X1 U19236 ( .A1(n16195), .A2(n19248), .A3(n16194), .ZN(n16196) );
  OAI211_X1 U19237 ( .C1(n18990), .C2(n14106), .A(n16197), .B(n16196), .ZN(
        P2_U2998) );
  AOI22_X1 U19238 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19235), .B1(n16268), 
        .B2(n19005), .ZN(n16203) );
  INV_X1 U19239 ( .A(n16198), .ZN(n16199) );
  OAI22_X1 U19240 ( .A1(n16200), .A2(n19237), .B1(n16260), .B2(n16199), .ZN(
        n16201) );
  AOI21_X1 U19241 ( .B1(n19255), .B2(n18995), .A(n16201), .ZN(n16202) );
  OAI211_X1 U19242 ( .C1(n16275), .C2(n18999), .A(n16203), .B(n16202), .ZN(
        P2_U2999) );
  AOI22_X1 U19243 ( .A1(n19245), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19235), .ZN(n16213) );
  INV_X1 U19244 ( .A(n16204), .ZN(n16209) );
  OAI21_X1 U19245 ( .B1(n16208), .B2(n16206), .A(n16205), .ZN(n16207) );
  OAI21_X1 U19246 ( .B1(n16209), .B2(n16208), .A(n16207), .ZN(n16317) );
  OAI21_X1 U19247 ( .B1(n16210), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15223), .ZN(n16315) );
  OAI22_X1 U19248 ( .A1(n16315), .A2(n16260), .B1(n14106), .B2(n16312), .ZN(
        n16211) );
  AOI21_X1 U19249 ( .B1(n19246), .B2(n16317), .A(n16211), .ZN(n16212) );
  OAI211_X1 U19250 ( .C1(n19253), .C2(n16214), .A(n16213), .B(n16212), .ZN(
        P2_U3000) );
  AOI22_X1 U19251 ( .A1(n19245), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19235), .ZN(n16222) );
  NAND2_X1 U19252 ( .A1(n19255), .A2(n16215), .ZN(n16218) );
  NAND2_X1 U19253 ( .A1(n16216), .A2(n19246), .ZN(n16217) );
  OAI211_X1 U19254 ( .C1(n16219), .C2(n16260), .A(n16218), .B(n16217), .ZN(
        n16220) );
  INV_X1 U19255 ( .A(n16220), .ZN(n16221) );
  OAI211_X1 U19256 ( .C1(n19253), .C2(n16223), .A(n16222), .B(n16221), .ZN(
        P2_U3002) );
  AOI22_X1 U19257 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19235), .B1(n16268), 
        .B2(n19031), .ZN(n16229) );
  INV_X1 U19258 ( .A(n16224), .ZN(n16226) );
  OAI22_X1 U19259 ( .A1(n16226), .A2(n16260), .B1(n16225), .B2(n19237), .ZN(
        n16227) );
  AOI21_X1 U19260 ( .B1(n19255), .B2(n19032), .A(n16227), .ZN(n16228) );
  OAI211_X1 U19261 ( .C1(n16275), .C2(n16230), .A(n16229), .B(n16228), .ZN(
        P2_U3003) );
  AOI22_X1 U19262 ( .A1(n19245), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19235), .ZN(n16235) );
  OAI22_X1 U19263 ( .A1(n16231), .A2(n19237), .B1(n14106), .B2(n19043), .ZN(
        n16232) );
  AOI21_X1 U19264 ( .B1(n19248), .B2(n16233), .A(n16232), .ZN(n16234) );
  OAI211_X1 U19265 ( .C1(n19253), .C2(n19038), .A(n16235), .B(n16234), .ZN(
        P2_U3004) );
  AOI22_X1 U19266 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19235), .B1(n16268), 
        .B2(n19056), .ZN(n16240) );
  OAI22_X1 U19267 ( .A1(n16237), .A2(n16260), .B1(n19237), .B2(n16236), .ZN(
        n16238) );
  AOI21_X1 U19268 ( .B1(n19255), .B2(n19057), .A(n16238), .ZN(n16239) );
  OAI211_X1 U19269 ( .C1(n16275), .C2(n16241), .A(n16240), .B(n16239), .ZN(
        P2_U3005) );
  AOI22_X1 U19270 ( .A1(n19245), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19235), .ZN(n16249) );
  NAND2_X1 U19271 ( .A1(n16242), .A2(n19248), .ZN(n16245) );
  NAND2_X1 U19272 ( .A1(n16243), .A2(n19246), .ZN(n16244) );
  OAI211_X1 U19273 ( .C1(n14106), .C2(n16246), .A(n16245), .B(n16244), .ZN(
        n16247) );
  INV_X1 U19274 ( .A(n16247), .ZN(n16248) );
  OAI211_X1 U19275 ( .C1(n19253), .C2(n16250), .A(n16249), .B(n16248), .ZN(
        P2_U3006) );
  OAI22_X1 U19276 ( .A1(n16275), .A2(n16251), .B1(n19889), .B2(n19041), .ZN(
        n16252) );
  AOI21_X1 U19277 ( .B1(n16268), .B2(n16253), .A(n16252), .ZN(n16257) );
  AOI22_X1 U19278 ( .A1(n16255), .A2(n19246), .B1(n19255), .B2(n16254), .ZN(
        n16256) );
  OAI211_X1 U19279 ( .C1(n16260), .C2(n16258), .A(n16257), .B(n16256), .ZN(
        P2_U3007) );
  AOI22_X1 U19280 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19235), .B1(n16268), 
        .B2(n19079), .ZN(n16265) );
  INV_X1 U19281 ( .A(n16259), .ZN(n19080) );
  OAI22_X1 U19282 ( .A1(n16262), .A2(n19237), .B1(n16261), .B2(n16260), .ZN(
        n16263) );
  AOI21_X1 U19283 ( .B1(n19255), .B2(n19080), .A(n16263), .ZN(n16264) );
  OAI211_X1 U19284 ( .C1(n16275), .C2(n16266), .A(n16265), .B(n16264), .ZN(
        P2_U3009) );
  AOI22_X1 U19285 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19235), .B1(n16268), 
        .B2(n16267), .ZN(n16274) );
  NAND3_X1 U19286 ( .A1(n16269), .A2(n15553), .A3(n19248), .ZN(n16270) );
  OAI21_X1 U19287 ( .B1(n14106), .B2(n9814), .A(n16270), .ZN(n16271) );
  AOI21_X1 U19288 ( .B1(n16272), .B2(n19246), .A(n16271), .ZN(n16273) );
  OAI211_X1 U19289 ( .C1(n16276), .C2(n16275), .A(n16274), .B(n16273), .ZN(
        P2_U3011) );
  OAI22_X1 U19290 ( .A1(n16277), .A2(n18968), .B1(n19912), .B2(n19041), .ZN(
        n16278) );
  AOI221_X1 U19291 ( .B1(n16281), .B2(n16280), .C1(n16279), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16278), .ZN(n16285) );
  INV_X1 U19292 ( .A(n16282), .ZN(n18964) );
  AOI22_X1 U19293 ( .A1(n16283), .A2(n16294), .B1(n16296), .B2(n18964), .ZN(
        n16284) );
  OAI211_X1 U19294 ( .C1(n16287), .C2(n16286), .A(n16285), .B(n16284), .ZN(
        P2_U3027) );
  INV_X1 U19295 ( .A(n16288), .ZN(n16289) );
  OAI21_X1 U19296 ( .B1(n16299), .B2(n16290), .A(n16289), .ZN(n16292) );
  AOI22_X1 U19297 ( .A1(n16292), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n16307), .B2(n16291), .ZN(n16303) );
  AOI222_X1 U19298 ( .A1(n16297), .A2(n16318), .B1(n16296), .B2(n16295), .C1(
        n16294), .C2(n16293), .ZN(n16302) );
  NAND2_X1 U19299 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n19235), .ZN(n16301) );
  NAND3_X1 U19300 ( .A1(n16299), .A2(n16298), .A3(n16183), .ZN(n16300) );
  NAND4_X1 U19301 ( .A1(n16303), .A2(n16302), .A3(n16301), .A4(n16300), .ZN(
        P2_U3028) );
  NAND2_X1 U19302 ( .A1(n16321), .A2(n16304), .ZN(n16305) );
  NAND2_X1 U19303 ( .A1(n16306), .A2(n16305), .ZN(n16309) );
  AOI22_X1 U19304 ( .A1(n16307), .A2(n19126), .B1(n19076), .B2(
        P2_REIP_REG_14__SCAN_IN), .ZN(n16308) );
  OAI21_X1 U19305 ( .B1(n16310), .B2(n16309), .A(n16308), .ZN(n16311) );
  INV_X1 U19306 ( .A(n16311), .ZN(n16320) );
  OAI22_X1 U19307 ( .A1(n16315), .A2(n16314), .B1(n16313), .B2(n16312), .ZN(
        n16316) );
  AOI21_X1 U19308 ( .B1(n16318), .B2(n16317), .A(n16316), .ZN(n16319) );
  OAI211_X1 U19309 ( .C1(n16322), .C2(n16321), .A(n16320), .B(n16319), .ZN(
        P2_U3032) );
  AOI22_X1 U19310 ( .A1(n16351), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16323), .B2(n16330), .ZN(n16355) );
  MUX2_X1 U19311 ( .A(n16325), .B(n16324), .S(n16330), .Z(n16354) );
  OAI21_X1 U19312 ( .B1(n16332), .B2(n19987), .A(n19978), .ZN(n16329) );
  INV_X1 U19313 ( .A(n16326), .ZN(n16328) );
  NOR2_X1 U19314 ( .A1(n16355), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16335) );
  INV_X1 U19315 ( .A(n16335), .ZN(n16327) );
  AOI22_X1 U19316 ( .A1(n16329), .A2(n16328), .B1(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16327), .ZN(n16331) );
  OAI211_X1 U19317 ( .C1(n19617), .C2(n16332), .A(n16331), .B(n16330), .ZN(
        n16333) );
  AOI222_X1 U19318 ( .A1(n16354), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .B1(n16354), .B2(n16333), .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .C2(n16333), .ZN(n16336) );
  OAI221_X1 U19319 ( .B1(n16336), .B2(n16335), .C1(n16336), .C2(n19968), .A(
        n16334), .ZN(n16353) );
  AOI22_X1 U19320 ( .A1(n16340), .A2(n16339), .B1(n16338), .B2(n16337), .ZN(
        n16344) );
  NAND2_X1 U19321 ( .A1(n16342), .A2(n16341), .ZN(n16343) );
  AND2_X1 U19322 ( .A1(n16344), .A2(n16343), .ZN(n19996) );
  NAND2_X1 U19323 ( .A1(n16345), .A2(n19259), .ZN(n16349) );
  OAI21_X1 U19324 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16346), .ZN(n16348) );
  NAND4_X1 U19325 ( .A1(n19996), .A2(n16349), .A3(n16348), .A4(n16347), .ZN(
        n16350) );
  AOI21_X1 U19326 ( .B1(n16351), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16350), .ZN(n16352) );
  OAI211_X1 U19327 ( .C1(n16355), .C2(n16354), .A(n16353), .B(n16352), .ZN(
        n16360) );
  NOR3_X1 U19328 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18906), .A3(n16356), 
        .ZN(n16357) );
  AOI211_X1 U19329 ( .C1(n16359), .C2(n16360), .A(n16358), .B(n16357), .ZN(
        n16373) );
  OR2_X1 U19330 ( .A1(n16360), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16366) );
  NAND3_X1 U19331 ( .A1(n16363), .A2(n16362), .A3(n16361), .ZN(n16365) );
  NAND2_X1 U19332 ( .A1(n16365), .A2(n16364), .ZN(n16367) );
  INV_X1 U19333 ( .A(n16367), .ZN(n16368) );
  AOI22_X1 U19334 ( .A1(n16370), .A2(n16369), .B1(n19869), .B2(n16368), .ZN(
        n16371) );
  AOI22_X1 U19335 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19850), .B1(n16371), 
        .B2(n18906), .ZN(n16372) );
  OAI211_X1 U19336 ( .C1(n19994), .C2(n16374), .A(n16373), .B(n16372), .ZN(
        P2_U3176) );
  NOR2_X1 U19337 ( .A1(n19850), .A2(n18906), .ZN(n16375) );
  OAI21_X1 U19338 ( .B1(n16375), .B2(n19979), .A(n16374), .ZN(P2_U3593) );
  INV_X1 U19339 ( .A(n16377), .ZN(n16390) );
  INV_X1 U19340 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16575) );
  INV_X1 U19341 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17898) );
  NAND2_X1 U19342 ( .A1(n17868), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17849) );
  NAND4_X1 U19343 ( .A1(n17807), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17734) );
  NAND2_X1 U19344 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17737) );
  INV_X1 U19345 ( .A(n17737), .ZN(n16750) );
  NAND2_X1 U19346 ( .A1(n16750), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17697) );
  INV_X1 U19347 ( .A(n17697), .ZN(n16378) );
  NAND2_X1 U19348 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17698) );
  NAND2_X1 U19349 ( .A1(n17679), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17658) );
  NAND2_X1 U19350 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17660) );
  NAND2_X1 U19351 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17645), .ZN(
        n17623) );
  NAND2_X1 U19352 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17624) );
  NAND2_X1 U19353 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17580) );
  NAND2_X1 U19354 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16380) );
  INV_X1 U19355 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16589) );
  NAND2_X1 U19356 ( .A1(n18829), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18737) );
  OAI21_X1 U19357 ( .B1(n17898), .B2(n17680), .A(n18347), .ZN(n17696) );
  NAND2_X1 U19358 ( .A1(n16379), .A2(n17696), .ZN(n16393) );
  XNOR2_X1 U19359 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16382) );
  NOR2_X1 U19360 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17680), .ZN(
        n16409) );
  INV_X1 U19361 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16664) );
  INV_X1 U19362 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17634) );
  INV_X1 U19363 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16724) );
  NAND2_X1 U19364 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17679), .ZN(
        n16726) );
  NAND3_X1 U19365 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n17657), .ZN(n16694) );
  NAND2_X1 U19366 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17620), .ZN(
        n16567) );
  NOR2_X1 U19367 ( .A1(n17634), .A2(n16567), .ZN(n16566) );
  INV_X1 U19368 ( .A(n16566), .ZN(n16565) );
  NAND2_X1 U19369 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17577), .ZN(
        n16563) );
  NOR2_X1 U19370 ( .A1(n17580), .A2(n16563), .ZN(n17541) );
  NAND2_X1 U19371 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17541), .ZN(
        n16559) );
  NOR2_X1 U19372 ( .A1(n16380), .A2(n16559), .ZN(n16407) );
  NAND2_X1 U19373 ( .A1(n18608), .A2(n16381), .ZN(n16413) );
  OAI211_X1 U19374 ( .C1(n16407), .C2(n18737), .A(n17904), .B(n16413), .ZN(
        n16416) );
  NOR2_X1 U19375 ( .A1(n16409), .A2(n16416), .ZN(n16392) );
  OAI22_X1 U19376 ( .A1(n16393), .A2(n16382), .B1(n16392), .B2(n16575), .ZN(
        n16383) );
  AOI211_X1 U19377 ( .C1(n17755), .C2(n16891), .A(n16384), .B(n16383), .ZN(
        n16389) );
  INV_X1 U19378 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16579) );
  XNOR2_X1 U19379 ( .A(n16579), .B(n16408), .ZN(n16578) );
  OAI221_X1 U19380 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16393), .C1(
        n16579), .C2(n16392), .A(n16391), .ZN(n16394) );
  AOI21_X1 U19381 ( .B1(n17755), .B2(n16578), .A(n16394), .ZN(n16402) );
  OAI22_X1 U19382 ( .A1(n16405), .A2(n17730), .B1(n16395), .B2(n17908), .ZN(
        n16400) );
  INV_X1 U19383 ( .A(n17562), .ZN(n16399) );
  AOI22_X1 U19384 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16400), .B1(
        n16399), .B2(n16398), .ZN(n16401) );
  OAI211_X1 U19385 ( .C1(n16403), .C2(n17790), .A(n16402), .B(n16401), .ZN(
        P3_U2800) );
  INV_X1 U19386 ( .A(n16404), .ZN(n16429) );
  AOI211_X1 U19387 ( .C1(n16406), .C2(n16429), .A(n16405), .B(n17730), .ZN(
        n16415) );
  INV_X1 U19388 ( .A(n16407), .ZN(n16556) );
  AOI21_X1 U19389 ( .B1(n16589), .B2(n16556), .A(n16408), .ZN(n16588) );
  OAI21_X1 U19390 ( .B1(n16409), .B2(n17755), .A(n16588), .ZN(n16410) );
  OAI211_X1 U19391 ( .C1(n16413), .C2(n16412), .A(n16411), .B(n16410), .ZN(
        n16414) );
  AOI211_X1 U19392 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16416), .A(
        n16415), .B(n16414), .ZN(n16421) );
  NOR2_X1 U19393 ( .A1(n16418), .A2(n16417), .ZN(n16432) );
  OAI211_X1 U19394 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16432), .A(
        n17897), .B(n16419), .ZN(n16420) );
  OAI211_X1 U19395 ( .C1(n16422), .C2(n17790), .A(n16421), .B(n16420), .ZN(
        P3_U2801) );
  INV_X1 U19396 ( .A(n17559), .ZN(n16423) );
  OAI21_X1 U19397 ( .B1(n17558), .B2(n17777), .A(n16423), .ZN(n17551) );
  NOR3_X1 U19398 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16424), .A3(
        n17551), .ZN(n16426) );
  OAI22_X1 U19399 ( .A1(n17777), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n17540), .B2(n17814), .ZN(n17552) );
  INV_X1 U19400 ( .A(n17552), .ZN(n16425) );
  OAI221_X1 U19401 ( .B1(n16426), .B2(n17559), .C1(n16426), .C2(n16425), .A(
        n18139), .ZN(n16438) );
  AOI211_X1 U19402 ( .C1(n16427), .C2(n17558), .A(n17404), .B(n18662), .ZN(
        n16428) );
  NAND2_X1 U19403 ( .A1(n17552), .A2(n17551), .ZN(n17550) );
  AOI22_X1 U19404 ( .A1(n18137), .A2(n16429), .B1(n16428), .B2(n17550), .ZN(
        n16430) );
  OAI211_X1 U19405 ( .C1(n16432), .C2(n18198), .A(n16431), .B(n16430), .ZN(
        n16433) );
  NAND3_X1 U19406 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18221), .A3(
        n16433), .ZN(n16437) );
  NAND2_X1 U19407 ( .A1(n18122), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17544) );
  NAND2_X1 U19408 ( .A1(n17731), .A2(n18137), .ZN(n16434) );
  NAND2_X1 U19409 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18129) );
  OAI22_X1 U19410 ( .A1(n18195), .A2(n18701), .B1(n18190), .B2(n18129), .ZN(
        n18179) );
  NAND2_X1 U19411 ( .A1(n18091), .A2(n18179), .ZN(n18051) );
  OAI211_X1 U19412 ( .C1(n18090), .C2(n18198), .A(n16434), .B(n18051), .ZN(
        n18075) );
  NAND2_X1 U19413 ( .A1(n17966), .A2(n18075), .ZN(n17965) );
  NAND4_X1 U19414 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16435), .A3(
        n18020), .A4(n17540), .ZN(n16436) );
  NAND4_X1 U19415 ( .A1(n16438), .A2(n16437), .A3(n17544), .A4(n16436), .ZN(
        P3_U2834) );
  NOR3_X1 U19416 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16440) );
  NOR4_X1 U19417 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16439) );
  NAND4_X1 U19418 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16440), .A3(n16439), .A4(
        U215), .ZN(U213) );
  INV_X1 U19419 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19187) );
  INV_X1 U19420 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16442) );
  OAI222_X1 U19421 ( .A1(U212), .A2(n19187), .B1(n16488), .B2(n20220), .C1(
        U214), .C2(n16442), .ZN(U216) );
  INV_X1 U19422 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n16523) );
  INV_X1 U19423 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20214) );
  INV_X1 U19424 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19192) );
  OAI222_X1 U19425 ( .A1(U214), .A2(n16523), .B1(n16488), .B2(n20214), .C1(
        U212), .C2(n19192), .ZN(U217) );
  INV_X1 U19426 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20208) );
  INV_X2 U19427 ( .A(U212), .ZN(n16486) );
  AOI22_X1 U19428 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16485), .ZN(n16443) );
  OAI21_X1 U19429 ( .B1(n20208), .B2(n16488), .A(n16443), .ZN(U218) );
  INV_X1 U19430 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20201) );
  AOI22_X1 U19431 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16485), .ZN(n16444) );
  OAI21_X1 U19432 ( .B1(n20201), .B2(n16488), .A(n16444), .ZN(U219) );
  INV_X1 U19433 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20195) );
  AOI22_X1 U19434 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16485), .ZN(n16445) );
  OAI21_X1 U19435 ( .B1(n20195), .B2(n16488), .A(n16445), .ZN(U220) );
  INV_X1 U19436 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20189) );
  AOI22_X1 U19437 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16485), .ZN(n16446) );
  OAI21_X1 U19438 ( .B1(n20189), .B2(n16488), .A(n16446), .ZN(U221) );
  INV_X1 U19439 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20182) );
  AOI22_X1 U19440 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16485), .ZN(n16447) );
  OAI21_X1 U19441 ( .B1(n20182), .B2(n16488), .A(n16447), .ZN(U222) );
  INV_X1 U19442 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20167) );
  AOI22_X1 U19443 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16485), .ZN(n16448) );
  OAI21_X1 U19444 ( .B1(n20167), .B2(n16488), .A(n16448), .ZN(U223) );
  INV_X1 U19445 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20226) );
  AOI22_X1 U19446 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16485), .ZN(n16449) );
  OAI21_X1 U19447 ( .B1(n20226), .B2(n16488), .A(n16449), .ZN(U224) );
  INV_X1 U19448 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20216) );
  AOI22_X1 U19449 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16485), .ZN(n16450) );
  OAI21_X1 U19450 ( .B1(n20216), .B2(n16488), .A(n16450), .ZN(U225) );
  AOI22_X1 U19451 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16485), .ZN(n16451) );
  OAI21_X1 U19452 ( .B1(n20210), .B2(n16488), .A(n16451), .ZN(U226) );
  INV_X1 U19453 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20204) );
  AOI22_X1 U19454 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16485), .ZN(n16452) );
  OAI21_X1 U19455 ( .B1(n20204), .B2(n16488), .A(n16452), .ZN(U227) );
  AOI22_X1 U19456 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16485), .ZN(n16453) );
  OAI21_X1 U19457 ( .B1(n20196), .B2(n16488), .A(n16453), .ZN(U228) );
  INV_X1 U19458 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20191) );
  AOI22_X1 U19459 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16485), .ZN(n16454) );
  OAI21_X1 U19460 ( .B1(n20191), .B2(n16488), .A(n16454), .ZN(U229) );
  AOI22_X1 U19461 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16485), .ZN(n16455) );
  OAI21_X1 U19462 ( .B1(n20184), .B2(n16488), .A(n16455), .ZN(U230) );
  INV_X1 U19463 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20178) );
  AOI22_X1 U19464 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16485), .ZN(n16456) );
  OAI21_X1 U19465 ( .B1(n20178), .B2(n16488), .A(n16456), .ZN(U231) );
  INV_X1 U19466 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16458) );
  AOI22_X1 U19467 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16485), .ZN(n16457) );
  OAI21_X1 U19468 ( .B1(n16458), .B2(n16488), .A(n16457), .ZN(U232) );
  AOI22_X1 U19469 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16485), .ZN(n16459) );
  OAI21_X1 U19470 ( .B1(n16460), .B2(n16488), .A(n16459), .ZN(U233) );
  AOI22_X1 U19471 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16485), .ZN(n16461) );
  OAI21_X1 U19472 ( .B1(n13456), .B2(n16488), .A(n16461), .ZN(U234) );
  AOI22_X1 U19473 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16485), .ZN(n16462) );
  OAI21_X1 U19474 ( .B1(n16463), .B2(n16488), .A(n16462), .ZN(U235) );
  AOI22_X1 U19475 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16485), .ZN(n16464) );
  OAI21_X1 U19476 ( .B1(n13461), .B2(n16488), .A(n16464), .ZN(U236) );
  AOI22_X1 U19477 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16485), .ZN(n16465) );
  OAI21_X1 U19478 ( .B1(n16466), .B2(n16488), .A(n16465), .ZN(U237) );
  AOI22_X1 U19479 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16485), .ZN(n16467) );
  OAI21_X1 U19480 ( .B1(n16468), .B2(n16488), .A(n16467), .ZN(U238) );
  AOI22_X1 U19481 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16485), .ZN(n16469) );
  OAI21_X1 U19482 ( .B1(n16470), .B2(n16488), .A(n16469), .ZN(U239) );
  INV_X1 U19483 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16472) );
  AOI22_X1 U19484 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16485), .ZN(n16471) );
  OAI21_X1 U19485 ( .B1(n16472), .B2(n16488), .A(n16471), .ZN(U240) );
  AOI22_X1 U19486 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16485), .ZN(n16473) );
  OAI21_X1 U19487 ( .B1(n16474), .B2(n16488), .A(n16473), .ZN(U241) );
  INV_X1 U19488 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16476) );
  AOI22_X1 U19489 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16485), .ZN(n16475) );
  OAI21_X1 U19490 ( .B1(n16476), .B2(n16488), .A(n16475), .ZN(U242) );
  AOI22_X1 U19491 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16485), .ZN(n16477) );
  OAI21_X1 U19492 ( .B1(n16478), .B2(n16488), .A(n16477), .ZN(U243) );
  INV_X1 U19493 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16480) );
  AOI22_X1 U19494 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16485), .ZN(n16479) );
  OAI21_X1 U19495 ( .B1(n16480), .B2(n16488), .A(n16479), .ZN(U244) );
  INV_X1 U19496 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U19497 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16485), .ZN(n16481) );
  OAI21_X1 U19498 ( .B1(n16482), .B2(n16488), .A(n16481), .ZN(U245) );
  INV_X1 U19499 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16484) );
  AOI22_X1 U19500 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16485), .ZN(n16483) );
  OAI21_X1 U19501 ( .B1(n16484), .B2(n16488), .A(n16483), .ZN(U246) );
  INV_X1 U19502 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U19503 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16486), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16485), .ZN(n16487) );
  OAI21_X1 U19504 ( .B1(n16489), .B2(n16488), .A(n16487), .ZN(U247) );
  OAI22_X1 U19505 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16521), .ZN(n16490) );
  INV_X1 U19506 ( .A(n16490), .ZN(U251) );
  OAI22_X1 U19507 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16521), .ZN(n16491) );
  INV_X1 U19508 ( .A(n16491), .ZN(U252) );
  OAI22_X1 U19509 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16521), .ZN(n16492) );
  INV_X1 U19510 ( .A(n16492), .ZN(U253) );
  OAI22_X1 U19511 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16521), .ZN(n16493) );
  INV_X1 U19512 ( .A(n16493), .ZN(U254) );
  OAI22_X1 U19513 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16521), .ZN(n16494) );
  INV_X1 U19514 ( .A(n16494), .ZN(U255) );
  OAI22_X1 U19515 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16521), .ZN(n16495) );
  INV_X1 U19516 ( .A(n16495), .ZN(U256) );
  OAI22_X1 U19517 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16521), .ZN(n16496) );
  INV_X1 U19518 ( .A(n16496), .ZN(U257) );
  OAI22_X1 U19519 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16521), .ZN(n16497) );
  INV_X1 U19520 ( .A(n16497), .ZN(U258) );
  OAI22_X1 U19521 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16521), .ZN(n16498) );
  INV_X1 U19522 ( .A(n16498), .ZN(U259) );
  OAI22_X1 U19523 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16513), .ZN(n16499) );
  INV_X1 U19524 ( .A(n16499), .ZN(U260) );
  OAI22_X1 U19525 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16513), .ZN(n16500) );
  INV_X1 U19526 ( .A(n16500), .ZN(U261) );
  OAI22_X1 U19527 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16521), .ZN(n16501) );
  INV_X1 U19528 ( .A(n16501), .ZN(U262) );
  OAI22_X1 U19529 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16513), .ZN(n16502) );
  INV_X1 U19530 ( .A(n16502), .ZN(U263) );
  OAI22_X1 U19531 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16521), .ZN(n16503) );
  INV_X1 U19532 ( .A(n16503), .ZN(U264) );
  OAI22_X1 U19533 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16521), .ZN(n16504) );
  INV_X1 U19534 ( .A(n16504), .ZN(U265) );
  OAI22_X1 U19535 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16513), .ZN(n16505) );
  INV_X1 U19536 ( .A(n16505), .ZN(U266) );
  OAI22_X1 U19537 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16513), .ZN(n16506) );
  INV_X1 U19538 ( .A(n16506), .ZN(U267) );
  OAI22_X1 U19539 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16513), .ZN(n16507) );
  INV_X1 U19540 ( .A(n16507), .ZN(U268) );
  OAI22_X1 U19541 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16513), .ZN(n16508) );
  INV_X1 U19542 ( .A(n16508), .ZN(U269) );
  OAI22_X1 U19543 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16513), .ZN(n16509) );
  INV_X1 U19544 ( .A(n16509), .ZN(U270) );
  OAI22_X1 U19545 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16513), .ZN(n16510) );
  INV_X1 U19546 ( .A(n16510), .ZN(U271) );
  OAI22_X1 U19547 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16521), .ZN(n16511) );
  INV_X1 U19548 ( .A(n16511), .ZN(U272) );
  OAI22_X1 U19549 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16521), .ZN(n16512) );
  INV_X1 U19550 ( .A(n16512), .ZN(U273) );
  OAI22_X1 U19551 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16513), .ZN(n16514) );
  INV_X1 U19552 ( .A(n16514), .ZN(U274) );
  OAI22_X1 U19553 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16521), .ZN(n16515) );
  INV_X1 U19554 ( .A(n16515), .ZN(U275) );
  OAI22_X1 U19555 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16521), .ZN(n16516) );
  INV_X1 U19556 ( .A(n16516), .ZN(U276) );
  OAI22_X1 U19557 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16521), .ZN(n16517) );
  INV_X1 U19558 ( .A(n16517), .ZN(U277) );
  OAI22_X1 U19559 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16521), .ZN(n16518) );
  INV_X1 U19560 ( .A(n16518), .ZN(U278) );
  OAI22_X1 U19561 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16521), .ZN(n16519) );
  INV_X1 U19562 ( .A(n16519), .ZN(U279) );
  OAI22_X1 U19563 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16521), .ZN(n16520) );
  INV_X1 U19564 ( .A(n16520), .ZN(U280) );
  INV_X1 U19565 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19282) );
  AOI22_X1 U19566 ( .A1(n16521), .A2(n19192), .B1(n19282), .B2(U215), .ZN(U281) );
  INV_X1 U19567 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19289) );
  AOI22_X1 U19568 ( .A1(n16521), .A2(n19187), .B1(n19289), .B2(U215), .ZN(U282) );
  INV_X1 U19569 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n16522) );
  OAI222_X1 U19570 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n19192), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n16523), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n16522), .ZN(n16524) );
  INV_X2 U19571 ( .A(n20831), .ZN(n20832) );
  INV_X1 U19572 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18774) );
  INV_X1 U19573 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19896) );
  AOI22_X1 U19574 ( .A1(n20832), .A2(n18774), .B1(n19896), .B2(n20831), .ZN(
        U347) );
  INV_X1 U19575 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18772) );
  INV_X1 U19576 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U19577 ( .A1(n20832), .A2(n18772), .B1(n19894), .B2(n20831), .ZN(
        U348) );
  INV_X1 U19578 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18769) );
  INV_X1 U19579 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19892) );
  AOI22_X1 U19580 ( .A1(n20832), .A2(n18769), .B1(n19892), .B2(n20831), .ZN(
        U349) );
  INV_X1 U19581 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18768) );
  INV_X1 U19582 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19890) );
  AOI22_X1 U19583 ( .A1(n20832), .A2(n18768), .B1(n19890), .B2(n20831), .ZN(
        U350) );
  INV_X1 U19584 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18766) );
  INV_X1 U19585 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19888) );
  AOI22_X1 U19586 ( .A1(n20832), .A2(n18766), .B1(n19888), .B2(n20831), .ZN(
        U351) );
  INV_X1 U19587 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18764) );
  INV_X1 U19588 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19886) );
  AOI22_X1 U19589 ( .A1(n20832), .A2(n18764), .B1(n19886), .B2(n20831), .ZN(
        U352) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18762) );
  INV_X1 U19591 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U19592 ( .A1(n20832), .A2(n18762), .B1(n19885), .B2(n20831), .ZN(
        U353) );
  INV_X1 U19593 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18759) );
  AOI22_X1 U19594 ( .A1(n20832), .A2(n18759), .B1(n19883), .B2(n20831), .ZN(
        U354) );
  INV_X1 U19595 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18813) );
  INV_X1 U19596 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19932) );
  AOI22_X1 U19597 ( .A1(n20832), .A2(n18813), .B1(n19932), .B2(n16524), .ZN(
        U356) );
  INV_X1 U19598 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18810) );
  INV_X1 U19599 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19930) );
  AOI22_X1 U19600 ( .A1(n20832), .A2(n18810), .B1(n19930), .B2(n16524), .ZN(
        U357) );
  INV_X1 U19601 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18809) );
  INV_X1 U19602 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19927) );
  AOI22_X1 U19603 ( .A1(n20832), .A2(n18809), .B1(n19927), .B2(n20831), .ZN(
        U358) );
  INV_X1 U19604 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18807) );
  INV_X1 U19605 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19926) );
  AOI22_X1 U19606 ( .A1(n20832), .A2(n18807), .B1(n19926), .B2(n20831), .ZN(
        U359) );
  INV_X1 U19607 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18804) );
  INV_X1 U19608 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19924) );
  AOI22_X1 U19609 ( .A1(n20832), .A2(n18804), .B1(n19924), .B2(n20831), .ZN(
        U360) );
  INV_X1 U19610 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18802) );
  INV_X1 U19611 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19922) );
  AOI22_X1 U19612 ( .A1(n20832), .A2(n18802), .B1(n19922), .B2(n20831), .ZN(
        U361) );
  INV_X1 U19613 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18799) );
  INV_X1 U19614 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19920) );
  AOI22_X1 U19615 ( .A1(n20832), .A2(n18799), .B1(n19920), .B2(n20831), .ZN(
        U362) );
  INV_X1 U19616 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18798) );
  INV_X1 U19617 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19918) );
  AOI22_X1 U19618 ( .A1(n20832), .A2(n18798), .B1(n19918), .B2(n20831), .ZN(
        U363) );
  INV_X1 U19619 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18796) );
  INV_X1 U19620 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19916) );
  AOI22_X1 U19621 ( .A1(n20832), .A2(n18796), .B1(n19916), .B2(n20831), .ZN(
        U364) );
  INV_X1 U19622 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18758) );
  INV_X1 U19623 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U19624 ( .A1(n20832), .A2(n18758), .B1(n19881), .B2(n20831), .ZN(
        U365) );
  INV_X1 U19625 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18793) );
  INV_X1 U19626 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19914) );
  AOI22_X1 U19627 ( .A1(n20832), .A2(n18793), .B1(n19914), .B2(n16524), .ZN(
        U366) );
  INV_X1 U19628 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18792) );
  INV_X1 U19629 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19913) );
  AOI22_X1 U19630 ( .A1(n20832), .A2(n18792), .B1(n19913), .B2(n16524), .ZN(
        U367) );
  INV_X1 U19631 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18790) );
  INV_X1 U19632 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19911) );
  AOI22_X1 U19633 ( .A1(n20832), .A2(n18790), .B1(n19911), .B2(n16524), .ZN(
        U368) );
  INV_X1 U19634 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18787) );
  INV_X1 U19635 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19909) );
  AOI22_X1 U19636 ( .A1(n20832), .A2(n18787), .B1(n19909), .B2(n16524), .ZN(
        U369) );
  INV_X1 U19637 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18786) );
  INV_X1 U19638 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U19639 ( .A1(n20832), .A2(n18786), .B1(n19907), .B2(n16524), .ZN(
        U370) );
  INV_X1 U19640 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18784) );
  INV_X1 U19641 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U19642 ( .A1(n20832), .A2(n18784), .B1(n19905), .B2(n16524), .ZN(
        U371) );
  INV_X1 U19643 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18781) );
  INV_X1 U19644 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19903) );
  AOI22_X1 U19645 ( .A1(n20832), .A2(n18781), .B1(n19903), .B2(n20831), .ZN(
        U372) );
  INV_X1 U19646 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18780) );
  INV_X1 U19647 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U19648 ( .A1(n20832), .A2(n18780), .B1(n19901), .B2(n20831), .ZN(
        U373) );
  INV_X1 U19649 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18778) );
  INV_X1 U19650 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19899) );
  AOI22_X1 U19651 ( .A1(n20832), .A2(n18778), .B1(n19899), .B2(n20831), .ZN(
        U374) );
  INV_X1 U19652 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18776) );
  INV_X1 U19653 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U19654 ( .A1(n20832), .A2(n18776), .B1(n19897), .B2(n20831), .ZN(
        U375) );
  INV_X1 U19655 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18755) );
  INV_X1 U19656 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U19657 ( .A1(n20832), .A2(n18755), .B1(n19879), .B2(n20831), .ZN(
        U376) );
  INV_X1 U19658 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18752) );
  NOR2_X1 U19659 ( .A1(n18739), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18744) );
  OAI22_X1 U19660 ( .A1(n18752), .A2(n18744), .B1(n18739), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18825) );
  INV_X1 U19661 ( .A(n18825), .ZN(n18828) );
  AOI21_X1 U19662 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18828), .ZN(n16525) );
  INV_X1 U19663 ( .A(n16525), .ZN(P3_U2633) );
  INV_X1 U19664 ( .A(n18729), .ZN(n18719) );
  OAI21_X1 U19665 ( .B1(n16531), .B2(n17473), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16526) );
  OAI21_X1 U19666 ( .B1(n16527), .B2(n18719), .A(n16526), .ZN(P3_U2634) );
  INV_X1 U19667 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18754) );
  AOI21_X1 U19668 ( .B1(n18752), .B2(n18754), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16528) );
  AOI22_X1 U19669 ( .A1(n18821), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16528), 
        .B2(n18894), .ZN(P3_U2635) );
  OAI21_X1 U19670 ( .B1(n18740), .B2(BS16), .A(n18828), .ZN(n18826) );
  OAI21_X1 U19671 ( .B1(n18828), .B2(n18884), .A(n18826), .ZN(P3_U2636) );
  NOR3_X1 U19672 ( .A1(n16531), .A2(n16530), .A3(n16529), .ZN(n18711) );
  NOR2_X1 U19673 ( .A1(n18711), .A2(n18715), .ZN(n18873) );
  OAI21_X1 U19674 ( .B1(n18873), .B2(n16533), .A(n16532), .ZN(P3_U2637) );
  NOR4_X1 U19675 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16537) );
  NOR4_X1 U19676 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16536) );
  NOR4_X1 U19677 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16535) );
  NOR4_X1 U19678 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16534) );
  NAND4_X1 U19679 ( .A1(n16537), .A2(n16536), .A3(n16535), .A4(n16534), .ZN(
        n16543) );
  NOR4_X1 U19680 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16541) );
  AOI211_X1 U19681 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16540) );
  NOR4_X1 U19682 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16539) );
  NOR4_X1 U19683 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16538) );
  NAND4_X1 U19684 ( .A1(n16541), .A2(n16540), .A3(n16539), .A4(n16538), .ZN(
        n16542) );
  NOR2_X1 U19685 ( .A1(n16543), .A2(n16542), .ZN(n18867) );
  INV_X1 U19686 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16545) );
  NOR3_X1 U19687 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16546) );
  OAI21_X1 U19688 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16546), .A(n18867), .ZN(
        n16544) );
  OAI21_X1 U19689 ( .B1(n18867), .B2(n16545), .A(n16544), .ZN(P3_U2638) );
  INV_X1 U19690 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18863) );
  INV_X1 U19691 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18827) );
  AOI21_X1 U19692 ( .B1(n18863), .B2(n18827), .A(n16546), .ZN(n16548) );
  INV_X1 U19693 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16547) );
  INV_X1 U19694 ( .A(n18867), .ZN(n18870) );
  AOI22_X1 U19695 ( .A1(n18867), .A2(n16548), .B1(n16547), .B2(n18870), .ZN(
        P3_U2639) );
  NOR2_X1 U19696 ( .A1(n18832), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18556) );
  INV_X1 U19697 ( .A(n18556), .ZN(n18727) );
  NAND4_X1 U19698 ( .A1(n18718), .A2(n18829), .A3(n18884), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18733) );
  INV_X1 U19699 ( .A(n18733), .ZN(n16905) );
  NOR2_X1 U19700 ( .A1(n18144), .A2(n16905), .ZN(n16881) );
  AOI211_X1 U19701 ( .C1(n18883), .C2(n18885), .A(n18880), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18716) );
  INV_X1 U19702 ( .A(n16552), .ZN(n16555) );
  AOI211_X4 U19703 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18244), .A(n18716), .B(
        n16555), .ZN(n16932) );
  INV_X1 U19704 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18817) );
  INV_X1 U19705 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18811) );
  INV_X1 U19706 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18808) );
  INV_X1 U19707 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18806) );
  INV_X1 U19708 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18801) );
  INV_X1 U19709 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18782) );
  INV_X1 U19710 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18779) );
  INV_X1 U19711 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18775) );
  INV_X1 U19712 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18767) );
  INV_X1 U19713 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18765) );
  NAND3_X1 U19714 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16869) );
  NAND2_X1 U19715 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n16841) );
  NOR4_X1 U19716 ( .A1(n18767), .A2(n18765), .A3(n16869), .A4(n16841), .ZN(
        n16831) );
  NAND2_X1 U19717 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16831), .ZN(n16806) );
  NAND2_X1 U19718 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16787) );
  NOR3_X1 U19719 ( .A1(n18775), .A2(n16806), .A3(n16787), .ZN(n16780) );
  NAND2_X1 U19720 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16780), .ZN(n16760) );
  NOR3_X1 U19721 ( .A1(n18782), .A2(n18779), .A3(n16760), .ZN(n16713) );
  NAND4_X1 U19722 ( .A1(n16713), .A2(P3_REIP_REG_17__SCAN_IN), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n16668) );
  NAND3_X1 U19723 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n16660) );
  NAND2_X1 U19724 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16669) );
  NOR3_X1 U19725 ( .A1(n16668), .A2(n16660), .A3(n16669), .ZN(n16649) );
  NAND2_X1 U19726 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16649), .ZN(n16638) );
  NOR2_X1 U19727 ( .A1(n18801), .A2(n16638), .ZN(n16632) );
  NAND2_X1 U19728 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16632), .ZN(n16627) );
  NOR2_X1 U19729 ( .A1(n18806), .A2(n16627), .ZN(n16569) );
  NAND2_X1 U19730 ( .A1(n16912), .A2(n16569), .ZN(n16610) );
  NOR3_X1 U19731 ( .A1(n18811), .A2(n18808), .A3(n16610), .ZN(n16592) );
  NAND2_X1 U19732 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16592), .ZN(n16571) );
  NOR3_X1 U19733 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18817), .A3(n16571), 
        .ZN(n16553) );
  AOI21_X1 U19734 ( .B1(n16932), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16553), .ZN(
        n16574) );
  NAND2_X1 U19735 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18244), .ZN(n16554) );
  AOI211_X4 U19736 ( .C1(n18884), .C2(n18886), .A(n16555), .B(n16554), .ZN(
        n16931) );
  NOR3_X1 U19737 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16903) );
  INV_X1 U19738 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16897) );
  NAND2_X1 U19739 ( .A1(n16903), .A2(n16897), .ZN(n16896) );
  NOR2_X1 U19740 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16896), .ZN(n16870) );
  INV_X1 U19741 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17248) );
  NAND2_X1 U19742 ( .A1(n16870), .A2(n17248), .ZN(n16866) );
  NOR2_X1 U19743 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16866), .ZN(n16849) );
  INV_X1 U19744 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17245) );
  NAND2_X1 U19745 ( .A1(n16849), .A2(n17245), .ZN(n16844) );
  NAND2_X1 U19746 ( .A1(n16818), .A2(n16820), .ZN(n16802) );
  INV_X1 U19747 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16793) );
  NAND2_X1 U19748 ( .A1(n16801), .A2(n16793), .ZN(n16792) );
  INV_X1 U19749 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16771) );
  NAND2_X1 U19750 ( .A1(n16772), .A2(n16771), .ZN(n16768) );
  INV_X1 U19751 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16741) );
  NAND2_X1 U19752 ( .A1(n16754), .A2(n16741), .ZN(n16738) );
  NAND2_X1 U19753 ( .A1(n16731), .A2(n17085), .ZN(n16721) );
  NOR2_X1 U19754 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16721), .ZN(n16706) );
  INV_X1 U19755 ( .A(n16706), .ZN(n16692) );
  INV_X1 U19756 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17039) );
  NAND2_X1 U19757 ( .A1(n16685), .A2(n17039), .ZN(n16675) );
  NOR2_X1 U19758 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16675), .ZN(n16663) );
  NAND2_X1 U19759 ( .A1(n16663), .A2(n16940), .ZN(n16655) );
  NOR2_X1 U19760 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16655), .ZN(n16643) );
  NAND2_X1 U19761 ( .A1(n16643), .A2(n16942), .ZN(n16633) );
  NOR2_X1 U19762 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16633), .ZN(n16618) );
  INV_X1 U19763 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16614) );
  NAND2_X1 U19764 ( .A1(n16618), .A2(n16614), .ZN(n16613) );
  NOR2_X1 U19765 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16613), .ZN(n16598) );
  INV_X1 U19766 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16980) );
  NAND2_X1 U19767 ( .A1(n16598), .A2(n16980), .ZN(n16576) );
  NOR2_X1 U19768 ( .A1(n16924), .A2(n16576), .ZN(n16583) );
  INV_X1 U19769 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16973) );
  INV_X1 U19770 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16558) );
  NOR2_X1 U19771 ( .A1(n16558), .A2(n16559), .ZN(n16557) );
  OAI21_X1 U19772 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16557), .A(
        n16556), .ZN(n17546) );
  INV_X1 U19773 ( .A(n17546), .ZN(n16601) );
  AOI21_X1 U19774 ( .B1(n16558), .B2(n16559), .A(n16557), .ZN(n17556) );
  OAI21_X1 U19775 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17541), .A(
        n16559), .ZN(n16560) );
  INV_X1 U19776 ( .A(n16560), .ZN(n17567) );
  INV_X1 U19777 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17595) );
  NOR2_X1 U19778 ( .A1(n17595), .A2(n16563), .ZN(n16562) );
  INV_X1 U19779 ( .A(n17541), .ZN(n16561) );
  OAI21_X1 U19780 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16562), .A(
        n16561), .ZN(n17582) );
  INV_X1 U19781 ( .A(n17582), .ZN(n16630) );
  AOI21_X1 U19782 ( .B1(n17595), .B2(n16563), .A(n16562), .ZN(n17591) );
  OAI21_X1 U19783 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17577), .A(
        n16563), .ZN(n16564) );
  INV_X1 U19784 ( .A(n16564), .ZN(n17607) );
  AOI21_X1 U19785 ( .B1(n16664), .B2(n16565), .A(n17577), .ZN(n17622) );
  AOI21_X1 U19786 ( .B1(n17634), .B2(n16567), .A(n16566), .ZN(n17630) );
  OAI21_X1 U19787 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17620), .A(
        n16567), .ZN(n16568) );
  INV_X1 U19788 ( .A(n16568), .ZN(n17649) );
  NAND2_X1 U19789 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17719), .ZN(
        n16775) );
  NOR2_X1 U19790 ( .A1(n17697), .A2(n16775), .ZN(n17695) );
  NAND2_X1 U19791 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17695), .ZN(
        n16736) );
  INV_X1 U19792 ( .A(n16736), .ZN(n16727) );
  INV_X1 U19793 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16920) );
  NAND2_X1 U19794 ( .A1(n16727), .A2(n16920), .ZN(n16703) );
  NAND2_X1 U19795 ( .A1(n16891), .A2(n16703), .ZN(n16728) );
  OAI21_X1 U19796 ( .B1(n17620), .B2(n9865), .A(n16728), .ZN(n16682) );
  NOR2_X1 U19797 ( .A1(n17649), .A2(n16682), .ZN(n16681) );
  NOR2_X1 U19798 ( .A1(n16681), .A2(n9865), .ZN(n16674) );
  NOR2_X1 U19799 ( .A1(n17630), .A2(n16674), .ZN(n16673) );
  NOR2_X1 U19800 ( .A1(n16650), .A2(n9865), .ZN(n16642) );
  NOR2_X1 U19801 ( .A1(n17591), .A2(n16642), .ZN(n16641) );
  NOR2_X1 U19802 ( .A1(n16641), .A2(n9865), .ZN(n16629) );
  NOR2_X1 U19803 ( .A1(n16630), .A2(n16629), .ZN(n16628) );
  NOR2_X1 U19804 ( .A1(n16628), .A2(n9865), .ZN(n16620) );
  NOR2_X1 U19805 ( .A1(n17567), .A2(n16620), .ZN(n16619) );
  NOR2_X1 U19806 ( .A1(n16619), .A2(n9865), .ZN(n16609) );
  NOR2_X1 U19807 ( .A1(n17556), .A2(n16609), .ZN(n16608) );
  NOR2_X1 U19808 ( .A1(n16608), .A2(n9865), .ZN(n16600) );
  NOR2_X1 U19809 ( .A1(n16601), .A2(n16600), .ZN(n16599) );
  NOR2_X1 U19810 ( .A1(n16599), .A2(n9865), .ZN(n16587) );
  NOR2_X1 U19811 ( .A1(n16588), .A2(n16587), .ZN(n16586) );
  NAND2_X1 U19812 ( .A1(n16891), .A2(n16905), .ZN(n16919) );
  INV_X1 U19813 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18812) );
  NAND2_X1 U19814 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16570) );
  OR2_X1 U19815 ( .A1(n16925), .A2(n16569), .ZN(n16626) );
  NAND2_X1 U19816 ( .A1(n16936), .A2(n16626), .ZN(n16623) );
  AOI221_X1 U19817 ( .B1(n18812), .B2(n16912), .C1(n16570), .C2(n16912), .A(
        n16623), .ZN(n16597) );
  NOR2_X1 U19818 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16571), .ZN(n16581) );
  INV_X1 U19819 ( .A(n16581), .ZN(n16572) );
  AOI21_X1 U19820 ( .B1(n16597), .B2(n16572), .A(n18814), .ZN(n16573) );
  NAND2_X1 U19821 ( .A1(n16931), .A2(n16576), .ZN(n16593) );
  XOR2_X1 U19822 ( .A(n16578), .B(n16577), .Z(n16582) );
  OAI22_X1 U19823 ( .A1(n16597), .A2(n18817), .B1(n16579), .B2(n16918), .ZN(
        n16580) );
  AOI211_X1 U19824 ( .C1(n16582), .C2(n16905), .A(n16581), .B(n16580), .ZN(
        n16585) );
  OAI21_X1 U19825 ( .B1(n16932), .B2(n16583), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16584) );
  OAI211_X1 U19826 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16593), .A(n16585), .B(
        n16584), .ZN(P3_U2641) );
  AOI211_X1 U19827 ( .C1(n16588), .C2(n16587), .A(n16586), .B(n18733), .ZN(
        n16591) );
  OAI22_X1 U19828 ( .A1(n16589), .A2(n16918), .B1(n16879), .B2(n16980), .ZN(
        n16590) );
  AOI211_X1 U19829 ( .C1(n16592), .C2(n18812), .A(n16591), .B(n16590), .ZN(
        n16596) );
  INV_X1 U19830 ( .A(n16593), .ZN(n16594) );
  OAI21_X1 U19831 ( .B1(n16598), .B2(n16980), .A(n16594), .ZN(n16595) );
  OAI211_X1 U19832 ( .C1(n16597), .C2(n18812), .A(n16596), .B(n16595), .ZN(
        P3_U2642) );
  NAND2_X1 U19833 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n18811), .ZN(n16607) );
  AOI22_X1 U19834 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16902), .B1(
        n16932), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16606) );
  INV_X1 U19835 ( .A(n16623), .ZN(n16617) );
  OAI21_X1 U19836 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16610), .A(n16617), 
        .ZN(n16604) );
  AOI211_X1 U19837 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16613), .A(n16598), .B(
        n16924), .ZN(n16603) );
  AOI211_X1 U19838 ( .C1(n16601), .C2(n16600), .A(n16599), .B(n18733), .ZN(
        n16602) );
  AOI211_X1 U19839 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16604), .A(n16603), 
        .B(n16602), .ZN(n16605) );
  OAI211_X1 U19840 ( .C1(n16610), .C2(n16607), .A(n16606), .B(n16605), .ZN(
        P3_U2643) );
  AOI211_X1 U19841 ( .C1(n17556), .C2(n16609), .A(n16608), .B(n18733), .ZN(
        n16612) );
  OAI22_X1 U19842 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16610), .B1(n16614), 
        .B2(n16879), .ZN(n16611) );
  AOI211_X1 U19843 ( .C1(n16902), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16612), .B(n16611), .ZN(n16616) );
  OAI211_X1 U19844 ( .C1(n16618), .C2(n16614), .A(n16931), .B(n16613), .ZN(
        n16615) );
  OAI211_X1 U19845 ( .C1(n16617), .C2(n18808), .A(n16616), .B(n16615), .ZN(
        P3_U2644) );
  AOI22_X1 U19846 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16902), .B1(
        n16932), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16625) );
  AOI211_X1 U19847 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16633), .A(n16618), .B(
        n16924), .ZN(n16622) );
  AOI211_X1 U19848 ( .C1(n17567), .C2(n16620), .A(n16619), .B(n18733), .ZN(
        n16621) );
  AOI211_X1 U19849 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16623), .A(n16622), 
        .B(n16621), .ZN(n16624) );
  OAI211_X1 U19850 ( .C1(n16627), .C2(n16626), .A(n16625), .B(n16624), .ZN(
        P3_U2645) );
  AOI22_X1 U19851 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16902), .B1(
        n16932), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16637) );
  NOR2_X1 U19852 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16925), .ZN(n16639) );
  AOI21_X1 U19853 ( .B1(n16638), .B2(n16912), .A(n16901), .ZN(n16648) );
  INV_X1 U19854 ( .A(n16648), .ZN(n16654) );
  AOI211_X1 U19855 ( .C1(n16630), .C2(n16629), .A(n16628), .B(n18733), .ZN(
        n16631) );
  AOI221_X1 U19856 ( .B1(n16639), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16654), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n16631), .ZN(n16636) );
  INV_X1 U19857 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18803) );
  NAND3_X1 U19858 ( .A1(n16912), .A2(n16632), .A3(n18803), .ZN(n16635) );
  OAI211_X1 U19859 ( .C1(n16643), .C2(n16942), .A(n16931), .B(n16633), .ZN(
        n16634) );
  NAND4_X1 U19860 ( .A1(n16637), .A2(n16636), .A3(n16635), .A4(n16634), .ZN(
        P3_U2646) );
  INV_X1 U19861 ( .A(n16638), .ZN(n16640) );
  AOI22_X1 U19862 ( .A1(n16932), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16640), 
        .B2(n16639), .ZN(n16647) );
  AOI211_X1 U19863 ( .C1(n17591), .C2(n16642), .A(n16641), .B(n18733), .ZN(
        n16645) );
  AOI211_X1 U19864 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16655), .A(n16643), .B(
        n16924), .ZN(n16644) );
  AOI211_X1 U19865 ( .C1(n16902), .C2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16645), .B(n16644), .ZN(n16646) );
  OAI211_X1 U19866 ( .C1(n16648), .C2(n18801), .A(n16647), .B(n16646), .ZN(
        P3_U2647) );
  NAND2_X1 U19867 ( .A1(n16912), .A2(n16649), .ZN(n16658) );
  AOI211_X1 U19868 ( .C1(n17607), .C2(n16651), .A(n16650), .B(n18733), .ZN(
        n16653) );
  OAI22_X1 U19869 ( .A1(n10038), .A2(n16918), .B1(n16879), .B2(n16940), .ZN(
        n16652) );
  AOI211_X1 U19870 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16654), .A(n16653), 
        .B(n16652), .ZN(n16657) );
  OAI211_X1 U19871 ( .C1(n16663), .C2(n16940), .A(n16931), .B(n16655), .ZN(
        n16656) );
  OAI211_X1 U19872 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16658), .A(n16657), 
        .B(n16656), .ZN(P3_U2648) );
  NOR2_X1 U19873 ( .A1(n16912), .A2(n16901), .ZN(n16748) );
  INV_X1 U19874 ( .A(n16748), .ZN(n16935) );
  INV_X1 U19875 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18788) );
  NAND2_X1 U19876 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16714) );
  NOR2_X1 U19877 ( .A1(n18788), .A2(n16714), .ZN(n16659) );
  INV_X1 U19878 ( .A(n16713), .ZN(n16725) );
  NOR2_X1 U19879 ( .A1(n16901), .A2(n16725), .ZN(n16753) );
  AOI21_X1 U19880 ( .B1(n16659), .B2(n16753), .A(n16748), .ZN(n16720) );
  AOI21_X1 U19881 ( .B1(n16660), .B2(n16935), .A(n16720), .ZN(n16689) );
  INV_X1 U19882 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18797) );
  AOI211_X1 U19883 ( .C1(n17622), .C2(n16662), .A(n16661), .B(n18733), .ZN(
        n16667) );
  AOI211_X1 U19884 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16675), .A(n16663), .B(
        n16924), .ZN(n16666) );
  OAI22_X1 U19885 ( .A1(n16664), .A2(n16918), .B1(n16879), .B2(n17003), .ZN(
        n16665) );
  NOR3_X1 U19886 ( .A1(n16667), .A2(n16666), .A3(n16665), .ZN(n16671) );
  INV_X1 U19887 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18794) );
  NOR2_X1 U19888 ( .A1(n16925), .A2(n16668), .ZN(n16709) );
  NAND3_X1 U19889 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16709), .ZN(n16690) );
  NOR2_X1 U19890 ( .A1(n18794), .A2(n16690), .ZN(n16672) );
  OAI211_X1 U19891 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16672), .B(n16669), .ZN(n16670) );
  OAI211_X1 U19892 ( .C1(n16689), .C2(n18797), .A(n16671), .B(n16670), .ZN(
        P3_U2649) );
  INV_X1 U19893 ( .A(n16672), .ZN(n16680) );
  INV_X1 U19894 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18795) );
  AOI211_X1 U19895 ( .C1(n17630), .C2(n16674), .A(n16673), .B(n18733), .ZN(
        n16678) );
  OAI211_X1 U19896 ( .C1(n16685), .C2(n17039), .A(n16931), .B(n16675), .ZN(
        n16676) );
  OAI21_X1 U19897 ( .B1(n16918), .B2(n17634), .A(n16676), .ZN(n16677) );
  AOI211_X1 U19898 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16932), .A(n16678), .B(
        n16677), .ZN(n16679) );
  OAI221_X1 U19899 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16680), .C1(n18795), 
        .C2(n16689), .A(n16679), .ZN(P3_U2650) );
  AOI211_X1 U19900 ( .C1(n17649), .C2(n16682), .A(n16681), .B(n18733), .ZN(
        n16687) );
  OAI21_X1 U19901 ( .B1(n16691), .B2(n16683), .A(n16931), .ZN(n16684) );
  OAI22_X1 U19902 ( .A1(n16685), .A2(n16684), .B1(n16879), .B2(n16683), .ZN(
        n16686) );
  AOI211_X1 U19903 ( .C1(n16902), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16687), .B(n16686), .ZN(n16688) );
  OAI221_X1 U19904 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n16690), .C1(n18794), 
        .C2(n16689), .A(n16688), .ZN(P3_U2651) );
  AOI211_X1 U19905 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16692), .A(n16691), .B(
        n16924), .ZN(n16693) );
  AOI21_X1 U19906 ( .B1(n16902), .B2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16693), .ZN(n16701) );
  NAND2_X1 U19907 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17657), .ZN(
        n16702) );
  INV_X1 U19908 ( .A(n16702), .ZN(n16695) );
  OAI21_X1 U19909 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16695), .A(
        n16694), .ZN(n17663) );
  OAI21_X1 U19910 ( .B1(n16703), .B2(n16702), .A(n16891), .ZN(n16696) );
  XOR2_X1 U19911 ( .A(n17663), .B(n16696), .Z(n16697) );
  AOI22_X1 U19912 ( .A1(n16932), .A2(P3_EBX_REG_19__SCAN_IN), .B1(n16905), 
        .B2(n16697), .ZN(n16700) );
  INV_X1 U19913 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18791) );
  INV_X1 U19914 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18789) );
  XOR2_X1 U19915 ( .A(n18791), .B(n18789), .Z(n16698) );
  AOI22_X1 U19916 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16720), .B1(n16709), 
        .B2(n16698), .ZN(n16699) );
  NAND4_X1 U19917 ( .A1(n16701), .A2(n16700), .A3(n16699), .A4(n18221), .ZN(
        P3_U2652) );
  AOI22_X1 U19918 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16902), .B1(
        n16932), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16712) );
  OAI21_X1 U19919 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17657), .A(
        n16702), .ZN(n17668) );
  INV_X1 U19920 ( .A(n17657), .ZN(n16704) );
  OAI21_X1 U19921 ( .B1(n16704), .B2(n16703), .A(n16891), .ZN(n16705) );
  XOR2_X1 U19922 ( .A(n17668), .B(n16705), .Z(n16708) );
  AOI211_X1 U19923 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16721), .A(n16706), .B(
        n16924), .ZN(n16707) );
  AOI211_X1 U19924 ( .C1(n16905), .C2(n16708), .A(n18122), .B(n16707), .ZN(
        n16711) );
  AOI22_X1 U19925 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16720), .B1(n16709), 
        .B2(n18789), .ZN(n16710) );
  NAND3_X1 U19926 ( .A1(n16712), .A2(n16711), .A3(n16710), .ZN(P3_U2653) );
  NAND2_X1 U19927 ( .A1(n16912), .A2(n16713), .ZN(n16746) );
  NOR2_X1 U19928 ( .A1(n16714), .A2(n16746), .ZN(n16719) );
  AOI21_X1 U19929 ( .B1(n16724), .B2(n16726), .A(n17657), .ZN(n17681) );
  OAI21_X1 U19930 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16726), .A(
        n16891), .ZN(n16716) );
  OAI21_X1 U19931 ( .B1(n17681), .B2(n16716), .A(n18221), .ZN(n16715) );
  AOI21_X1 U19932 ( .B1(n17681), .B2(n16716), .A(n16715), .ZN(n16717) );
  OAI22_X1 U19933 ( .A1(n16881), .A2(n16717), .B1(n16879), .B2(n17085), .ZN(
        n16718) );
  AOI221_X1 U19934 ( .B1(n16720), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16719), 
        .C2(n18788), .A(n16718), .ZN(n16723) );
  OAI211_X1 U19935 ( .C1(n16731), .C2(n17085), .A(n16931), .B(n16721), .ZN(
        n16722) );
  OAI211_X1 U19936 ( .C1(n16918), .C2(n16724), .A(n16723), .B(n16722), .ZN(
        P3_U2654) );
  INV_X1 U19937 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18783) );
  AOI221_X1 U19938 ( .B1(n16725), .B2(n16912), .C1(n18783), .C2(n16912), .A(
        n16901), .ZN(n16747) );
  INV_X1 U19939 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18785) );
  INV_X1 U19940 ( .A(n16728), .ZN(n16737) );
  OAI21_X1 U19941 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16727), .A(
        n16726), .ZN(n17701) );
  INV_X1 U19942 ( .A(n17701), .ZN(n16729) );
  AOI221_X1 U19943 ( .B1(n16737), .B2(n16729), .C1(n16728), .C2(n17701), .A(
        n18733), .ZN(n16730) );
  AOI211_X1 U19944 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n16902), .A(
        n18122), .B(n16730), .ZN(n16735) );
  NOR3_X1 U19945 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18783), .A3(n16746), 
        .ZN(n16733) );
  AOI211_X1 U19946 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16738), .A(n16731), .B(
        n16924), .ZN(n16732) );
  AOI211_X1 U19947 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16932), .A(n16733), .B(
        n16732), .ZN(n16734) );
  OAI211_X1 U19948 ( .C1(n16747), .C2(n18785), .A(n16735), .B(n16734), .ZN(
        P3_U2655) );
  OAI21_X1 U19949 ( .B1(n9865), .B2(n16920), .A(n16905), .ZN(n16921) );
  OAI21_X1 U19950 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17695), .A(
        n16736), .ZN(n17708) );
  AOI211_X1 U19951 ( .C1(n16891), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16921), .B(n17708), .ZN(n16744) );
  NAND3_X1 U19952 ( .A1(n17708), .A2(n16905), .A3(n16737), .ZN(n16740) );
  OAI211_X1 U19953 ( .C1(n16754), .C2(n16741), .A(n16931), .B(n16738), .ZN(
        n16739) );
  NAND2_X1 U19954 ( .A1(n16740), .A2(n16739), .ZN(n16743) );
  INV_X1 U19955 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17712) );
  OAI22_X1 U19956 ( .A1(n17712), .A2(n16918), .B1(n16879), .B2(n16741), .ZN(
        n16742) );
  NOR4_X1 U19957 ( .A1(n18144), .A2(n16744), .A3(n16743), .A4(n16742), .ZN(
        n16745) );
  OAI221_X1 U19958 ( .B1(n16747), .B2(n18783), .C1(n16747), .C2(n16746), .A(
        n16745), .ZN(P3_U2656) );
  OR2_X1 U19959 ( .A1(n16748), .A2(n16753), .ZN(n16759) );
  INV_X1 U19960 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17721) );
  INV_X1 U19961 ( .A(n16775), .ZN(n17736) );
  NAND2_X1 U19962 ( .A1(n16750), .A2(n17736), .ZN(n16761) );
  AOI21_X1 U19963 ( .B1(n17721), .B2(n16761), .A(n17695), .ZN(n17723) );
  NOR2_X1 U19964 ( .A1(n17898), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16906) );
  INV_X1 U19965 ( .A(n16906), .ZN(n16892) );
  NOR2_X1 U19966 ( .A1(n17733), .A2(n16892), .ZN(n16852) );
  INV_X1 U19967 ( .A(n16852), .ZN(n16749) );
  OAI21_X1 U19968 ( .B1(n17734), .B2(n16749), .A(n16891), .ZN(n16777) );
  OAI21_X1 U19969 ( .B1(n16750), .B2(n9865), .A(n16777), .ZN(n16763) );
  OAI21_X1 U19970 ( .B1(n17723), .B2(n16763), .A(n16905), .ZN(n16751) );
  AOI21_X1 U19971 ( .B1(n17723), .B2(n16763), .A(n16751), .ZN(n16752) );
  AOI211_X1 U19972 ( .C1(n16932), .C2(P3_EBX_REG_14__SCAN_IN), .A(n18122), .B(
        n16752), .ZN(n16758) );
  NOR4_X1 U19973 ( .A1(n16753), .A2(n18779), .A3(n16925), .A4(n16760), .ZN(
        n16756) );
  AOI211_X1 U19974 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16768), .A(n16754), .B(
        n16924), .ZN(n16755) );
  AOI211_X1 U19975 ( .C1(n16902), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16756), .B(n16755), .ZN(n16757) );
  OAI211_X1 U19976 ( .C1(n18782), .C2(n16759), .A(n16758), .B(n16757), .ZN(
        P3_U2657) );
  OAI21_X1 U19977 ( .B1(n16780), .B2(n16925), .A(n16936), .ZN(n16791) );
  NOR2_X1 U19978 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16925), .ZN(n16779) );
  OR2_X1 U19979 ( .A1(n16925), .A2(n16760), .ZN(n16766) );
  INV_X1 U19980 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16776) );
  NOR2_X1 U19981 ( .A1(n16776), .A2(n16775), .ZN(n16774) );
  OAI21_X1 U19982 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16774), .A(
        n16761), .ZN(n17739) );
  AOI211_X1 U19983 ( .C1(n16891), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16921), .B(n17739), .ZN(n16762) );
  AOI211_X1 U19984 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16902), .A(
        n18122), .B(n16762), .ZN(n16765) );
  NAND3_X1 U19985 ( .A1(n16905), .A2(n17739), .A3(n16763), .ZN(n16764) );
  OAI211_X1 U19986 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16766), .A(n16765), 
        .B(n16764), .ZN(n16767) );
  AOI221_X1 U19987 ( .B1(n16791), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16779), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16767), .ZN(n16770) );
  OAI211_X1 U19988 ( .C1(n16772), .C2(n16771), .A(n16931), .B(n16768), .ZN(
        n16769) );
  OAI211_X1 U19989 ( .C1(n16771), .C2(n16879), .A(n16770), .B(n16769), .ZN(
        P3_U2658) );
  AOI211_X1 U19990 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16792), .A(n16772), .B(
        n16924), .ZN(n16773) );
  AOI21_X1 U19991 ( .B1(n16902), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16773), .ZN(n16783) );
  AOI21_X1 U19992 ( .B1(n16776), .B2(n16775), .A(n16774), .ZN(n17754) );
  XNOR2_X1 U19993 ( .A(n17754), .B(n16777), .ZN(n16778) );
  AOI22_X1 U19994 ( .A1(n16932), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n16905), 
        .B2(n16778), .ZN(n16782) );
  AOI22_X1 U19995 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16791), .B1(n16780), 
        .B2(n16779), .ZN(n16781) );
  NAND4_X1 U19996 ( .A1(n16783), .A2(n16782), .A3(n16781), .A4(n18221), .ZN(
        P3_U2659) );
  INV_X1 U19997 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16788) );
  NAND2_X1 U19998 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17768), .ZN(
        n16861) );
  NOR2_X1 U19999 ( .A1(n10034), .A2(n16861), .ZN(n16851) );
  NAND2_X1 U20000 ( .A1(n17807), .A2(n16851), .ZN(n16810) );
  INV_X1 U20001 ( .A(n16810), .ZN(n16827) );
  NAND2_X1 U20002 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16827), .ZN(
        n16797) );
  INV_X1 U20003 ( .A(n16797), .ZN(n16798) );
  NAND2_X1 U20004 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16798), .ZN(
        n16784) );
  AOI21_X1 U20005 ( .B1(n16788), .B2(n16784), .A(n17736), .ZN(n17763) );
  INV_X1 U20006 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17782) );
  NAND2_X1 U20007 ( .A1(n16798), .A2(n16920), .ZN(n16799) );
  OAI21_X1 U20008 ( .B1(n17782), .B2(n16799), .A(n16891), .ZN(n16786) );
  OAI21_X1 U20009 ( .B1(n17763), .B2(n16786), .A(n18221), .ZN(n16785) );
  AOI21_X1 U20010 ( .B1(n17763), .B2(n16786), .A(n16785), .ZN(n16796) );
  INV_X1 U20011 ( .A(n16806), .ZN(n16829) );
  NAND2_X1 U20012 ( .A1(n16912), .A2(n16829), .ZN(n16805) );
  OAI21_X1 U20013 ( .B1(n16787), .B2(n16805), .A(n18775), .ZN(n16790) );
  OAI22_X1 U20014 ( .A1(n16788), .A2(n16918), .B1(n16879), .B2(n16793), .ZN(
        n16789) );
  AOI21_X1 U20015 ( .B1(n16791), .B2(n16790), .A(n16789), .ZN(n16795) );
  OAI211_X1 U20016 ( .C1(n16801), .C2(n16793), .A(n16931), .B(n16792), .ZN(
        n16794) );
  OAI211_X1 U20017 ( .C1(n16881), .C2(n16796), .A(n16795), .B(n16794), .ZN(
        P3_U2660) );
  AOI22_X1 U20018 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16798), .B1(
        n16797), .B2(n17782), .ZN(n17784) );
  NAND2_X1 U20019 ( .A1(n16891), .A2(n16799), .ZN(n16811) );
  XNOR2_X1 U20020 ( .A(n17784), .B(n16811), .ZN(n16800) );
  AOI22_X1 U20021 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16902), .B1(
        n16905), .B2(n16800), .ZN(n16809) );
  INV_X1 U20022 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18771) );
  NOR3_X1 U20023 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18771), .A3(n16805), 
        .ZN(n16804) );
  AOI211_X1 U20024 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16802), .A(n16801), .B(
        n16924), .ZN(n16803) );
  AOI211_X1 U20025 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16932), .A(n16804), .B(
        n16803), .ZN(n16808) );
  NOR2_X1 U20026 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16805), .ZN(n16819) );
  AOI21_X1 U20027 ( .B1(n16806), .B2(n16912), .A(n16901), .ZN(n16824) );
  INV_X1 U20028 ( .A(n16824), .ZN(n16832) );
  OAI21_X1 U20029 ( .B1(n16819), .B2(n16832), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16807) );
  NAND4_X1 U20030 ( .A1(n16809), .A2(n16808), .A3(n18221), .A4(n16807), .ZN(
        P3_U2661) );
  INV_X1 U20031 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16814) );
  NAND2_X1 U20032 ( .A1(n16827), .A2(n16814), .ZN(n16812) );
  OAI22_X1 U20033 ( .A1(n16814), .A2(n16827), .B1(n16810), .B2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16813) );
  OAI22_X1 U20034 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16812), .B1(
        n16811), .B2(n16813), .ZN(n16816) );
  INV_X1 U20035 ( .A(n16813), .ZN(n17797) );
  NAND2_X1 U20036 ( .A1(n16905), .A2(n9865), .ZN(n16909) );
  OAI22_X1 U20037 ( .A1(n17797), .A2(n16909), .B1(n16814), .B2(n16918), .ZN(
        n16815) );
  AOI211_X1 U20038 ( .C1(n16905), .C2(n16816), .A(n18122), .B(n16815), .ZN(
        n16823) );
  AOI21_X1 U20039 ( .B1(n16931), .B2(n16818), .A(n16932), .ZN(n16817) );
  INV_X1 U20040 ( .A(n16817), .ZN(n16821) );
  NOR2_X1 U20041 ( .A1(n16818), .A2(n16924), .ZN(n16826) );
  AOI221_X1 U20042 ( .B1(n16821), .B2(P3_EBX_REG_9__SCAN_IN), .C1(n16826), 
        .C2(n16820), .A(n16819), .ZN(n16822) );
  OAI211_X1 U20043 ( .C1(n16824), .C2(n18771), .A(n16823), .B(n16822), .ZN(
        P3_U2662) );
  NAND2_X1 U20044 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16844), .ZN(n16825) );
  AOI22_X1 U20045 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16902), .B1(
        n16826), .B2(n16825), .ZN(n16835) );
  NAND2_X1 U20046 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16851), .ZN(
        n16836) );
  AOI21_X1 U20047 ( .B1(n17806), .B2(n16836), .A(n16827), .ZN(n17810) );
  OAI21_X1 U20048 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16836), .A(
        n16891), .ZN(n16839) );
  XNOR2_X1 U20049 ( .A(n17810), .B(n16839), .ZN(n16828) );
  AOI22_X1 U20050 ( .A1(n16932), .A2(P3_EBX_REG_8__SCAN_IN), .B1(n16905), .B2(
        n16828), .ZN(n16834) );
  NOR2_X1 U20051 ( .A1(n16829), .A2(n16925), .ZN(n16830) );
  AOI22_X1 U20052 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16832), .B1(n16831), 
        .B2(n16830), .ZN(n16833) );
  NAND4_X1 U20053 ( .A1(n16835), .A2(n16834), .A3(n16833), .A4(n18221), .ZN(
        P3_U2663) );
  AOI22_X1 U20054 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16902), .B1(
        n16932), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n16848) );
  OAI21_X1 U20055 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16851), .A(
        n16836), .ZN(n16837) );
  INV_X1 U20056 ( .A(n16837), .ZN(n17830) );
  OAI21_X1 U20057 ( .B1(n9865), .B2(n16852), .A(n17830), .ZN(n16838) );
  OAI21_X1 U20058 ( .B1(n17830), .B2(n16839), .A(n16838), .ZN(n16840) );
  AOI21_X1 U20059 ( .B1(n16905), .B2(n16840), .A(n18122), .ZN(n16847) );
  OAI21_X1 U20060 ( .B1(n16841), .B2(n16869), .A(n16912), .ZN(n16842) );
  NAND2_X1 U20061 ( .A1(n16842), .A2(n16936), .ZN(n16865) );
  INV_X1 U20062 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18763) );
  INV_X1 U20063 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18760) );
  NAND3_X1 U20064 ( .A1(n16912), .A2(P3_REIP_REG_1__SCAN_IN), .A3(
        P3_REIP_REG_2__SCAN_IN), .ZN(n16888) );
  NOR2_X1 U20065 ( .A1(n18760), .A2(n16888), .ZN(n16884) );
  NAND2_X1 U20066 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16884), .ZN(n16860) );
  NOR2_X1 U20067 ( .A1(n18763), .A2(n16860), .ZN(n16856) );
  XOR2_X1 U20068 ( .A(n18767), .B(n18765), .Z(n16843) );
  AOI22_X1 U20069 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16865), .B1(n16856), 
        .B2(n16843), .ZN(n16846) );
  OAI211_X1 U20070 ( .C1(n16849), .C2(n17245), .A(n16931), .B(n16844), .ZN(
        n16845) );
  NAND4_X1 U20071 ( .A1(n16848), .A2(n16847), .A3(n16846), .A4(n16845), .ZN(
        P3_U2664) );
  AOI211_X1 U20072 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16866), .A(n16849), .B(
        n16924), .ZN(n16850) );
  AOI21_X1 U20073 ( .B1(n16902), .B2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16850), .ZN(n16859) );
  AOI21_X1 U20074 ( .B1(n10034), .B2(n16861), .A(n16851), .ZN(n16853) );
  NOR3_X1 U20075 ( .A1(n16853), .A2(n16852), .A3(n16919), .ZN(n16855) );
  INV_X1 U20076 ( .A(n16853), .ZN(n17840) );
  AOI211_X1 U20077 ( .C1(n16891), .C2(n16861), .A(n16921), .B(n17840), .ZN(
        n16854) );
  AOI211_X1 U20078 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16932), .A(n16855), .B(
        n16854), .ZN(n16858) );
  AOI22_X1 U20079 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16865), .B1(n16856), 
        .B2(n18765), .ZN(n16857) );
  NAND4_X1 U20080 ( .A1(n16859), .A2(n16858), .A3(n16857), .A4(n18221), .ZN(
        P3_U2665) );
  NAND2_X1 U20081 ( .A1(n18763), .A2(n16860), .ZN(n16864) );
  NOR2_X1 U20082 ( .A1(n17898), .A2(n17849), .ZN(n16873) );
  OAI21_X1 U20083 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16873), .A(
        n16861), .ZN(n17853) );
  OAI21_X1 U20084 ( .B1(n17849), .B2(n16892), .A(n16891), .ZN(n16875) );
  XNOR2_X1 U20085 ( .A(n17853), .B(n16875), .ZN(n16862) );
  OAI22_X1 U20086 ( .A1(n16879), .A2(n17248), .B1(n18733), .B2(n16862), .ZN(
        n16863) );
  AOI211_X1 U20087 ( .C1(n16865), .C2(n16864), .A(n18122), .B(n16863), .ZN(
        n16868) );
  OAI211_X1 U20088 ( .C1(n16870), .C2(n17248), .A(n16931), .B(n16866), .ZN(
        n16867) );
  OAI211_X1 U20089 ( .C1(n16918), .C2(n17850), .A(n16868), .B(n16867), .ZN(
        P3_U2666) );
  INV_X1 U20090 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18761) );
  AOI21_X1 U20091 ( .B1(n16912), .B2(n16869), .A(n16901), .ZN(n16887) );
  AOI211_X1 U20092 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16896), .A(n16870), .B(
        n16924), .ZN(n16871) );
  AOI21_X1 U20093 ( .B1(n16902), .B2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16871), .ZN(n16886) );
  NOR2_X1 U20094 ( .A1(n18238), .A2(n18898), .ZN(n16934) );
  INV_X1 U20095 ( .A(n16934), .ZN(n18900) );
  AOI21_X1 U20096 ( .B1(n17218), .B2(n16872), .A(n18900), .ZN(n16883) );
  INV_X1 U20097 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16874) );
  NAND2_X1 U20098 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17868), .ZN(
        n16889) );
  AOI21_X1 U20099 ( .B1(n16874), .B2(n16889), .A(n16873), .ZN(n17869) );
  NAND2_X1 U20100 ( .A1(n17868), .A2(n16874), .ZN(n17864) );
  OAI22_X1 U20101 ( .A1(n17869), .A2(n16875), .B1(n16892), .B2(n17864), .ZN(
        n16876) );
  AOI211_X1 U20102 ( .C1(n17869), .C2(n9865), .A(n18122), .B(n16876), .ZN(
        n16880) );
  OAI22_X1 U20103 ( .A1(n16881), .A2(n16880), .B1(n16879), .B2(n16878), .ZN(
        n16882) );
  AOI211_X1 U20104 ( .C1(n16884), .C2(n18761), .A(n16883), .B(n16882), .ZN(
        n16885) );
  OAI211_X1 U20105 ( .C1(n18761), .C2(n16887), .A(n16886), .B(n16885), .ZN(
        P3_U2667) );
  AOI21_X1 U20106 ( .B1(n18760), .B2(n16888), .A(n16887), .ZN(n16895) );
  NOR2_X1 U20107 ( .A1(n17898), .A2(n17892), .ZN(n16890) );
  OAI21_X1 U20108 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16890), .A(
        n16889), .ZN(n17877) );
  OAI21_X1 U20109 ( .B1(n17892), .B2(n16892), .A(n16891), .ZN(n16908) );
  XNOR2_X1 U20110 ( .A(n17877), .B(n16908), .ZN(n16893) );
  OAI21_X1 U20111 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18672), .A(
        n17218), .ZN(n18834) );
  OAI22_X1 U20112 ( .A1(n18733), .A2(n16893), .B1(n18900), .B2(n18834), .ZN(
        n16894) );
  AOI211_X1 U20113 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16932), .A(n16895), .B(
        n16894), .ZN(n16899) );
  OAI211_X1 U20114 ( .C1(n16903), .C2(n16897), .A(n16931), .B(n16896), .ZN(
        n16898) );
  OAI211_X1 U20115 ( .C1(n16918), .C2(n16900), .A(n16899), .B(n16898), .ZN(
        P3_U2668) );
  AOI22_X1 U20116 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16902), .B1(
        P3_REIP_REG_2__SCAN_IN), .B2(n16901), .ZN(n16916) );
  INV_X1 U20117 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17277) );
  INV_X1 U20118 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17271) );
  NAND2_X1 U20119 ( .A1(n17277), .A2(n17271), .ZN(n16923) );
  AOI211_X1 U20120 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16923), .A(n16903), .B(
        n16924), .ZN(n16904) );
  AOI21_X1 U20121 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n16932), .A(n16904), .ZN(
        n16915) );
  AOI21_X1 U20122 ( .B1(n18849), .B2(n18670), .A(n18672), .ZN(n18845) );
  AOI22_X1 U20123 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17892), .B1(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17898), .ZN(n17888) );
  OAI21_X1 U20124 ( .B1(n16906), .B2(n17888), .A(n16905), .ZN(n16907) );
  OAI22_X1 U20125 ( .A1(n17888), .A2(n16909), .B1(n16908), .B2(n16907), .ZN(
        n16910) );
  AOI21_X1 U20126 ( .B1(n18845), .B2(n16934), .A(n16910), .ZN(n16914) );
  NAND2_X1 U20127 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16911) );
  OAI211_X1 U20128 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16912), .B(n16911), .ZN(n16913) );
  NAND4_X1 U20129 ( .A1(n16916), .A2(n16915), .A3(n16914), .A4(n16913), .ZN(
        P3_U2669) );
  AND2_X1 U20130 ( .A1(n16917), .A2(n18670), .ZN(n18853) );
  AOI22_X1 U20131 ( .A1(n16932), .A2(P3_EBX_REG_1__SCAN_IN), .B1(n18853), .B2(
        n16934), .ZN(n16930) );
  OAI21_X1 U20132 ( .B1(n16920), .B2(n16919), .A(n16918), .ZN(n16928) );
  OAI22_X1 U20133 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16921), .B1(
        n16936), .B2(n18863), .ZN(n16927) );
  NOR2_X1 U20134 ( .A1(n17277), .A2(n17271), .ZN(n17264) );
  INV_X1 U20135 ( .A(n17264), .ZN(n16922) );
  NAND2_X1 U20136 ( .A1(n16923), .A2(n16922), .ZN(n17273) );
  OAI22_X1 U20137 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16925), .B1(n16924), 
        .B2(n17273), .ZN(n16926) );
  AOI211_X1 U20138 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16928), .A(
        n16927), .B(n16926), .ZN(n16929) );
  NAND2_X1 U20139 ( .A1(n16930), .A2(n16929), .ZN(P3_U2670) );
  NOR2_X1 U20140 ( .A1(n16932), .A2(n16931), .ZN(n16939) );
  AOI22_X1 U20141 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16935), .B1(n16934), 
        .B2(n16933), .ZN(n16938) );
  NAND3_X1 U20142 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18896), .A3(
        n16936), .ZN(n16937) );
  OAI211_X1 U20143 ( .C1(n16939), .C2(n17277), .A(n16938), .B(n16937), .ZN(
        P3_U2671) );
  NOR2_X1 U20144 ( .A1(n16940), .A2(n17003), .ZN(n16944) );
  NAND2_X1 U20145 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16981), .ZN(n16941) );
  NAND2_X1 U20146 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17074), .ZN(n17038) );
  NOR4_X1 U20147 ( .A1(n16980), .A2(n16942), .A3(n16941), .A4(n17038), .ZN(
        n16943) );
  NAND4_X1 U20148 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16944), .A4(n16943), .ZN(n16972) );
  NOR2_X1 U20149 ( .A1(n16973), .A2(n16972), .ZN(n16971) );
  NAND2_X1 U20150 ( .A1(n17266), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16946) );
  NAND2_X1 U20151 ( .A1(n16971), .A2(n17402), .ZN(n16945) );
  OAI22_X1 U20152 ( .A1(n16971), .A2(n16946), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16945), .ZN(P3_U2672) );
  AOI22_X1 U20153 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17090), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16957) );
  INV_X1 U20154 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U20155 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20156 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16947) );
  OAI211_X1 U20157 ( .C1(n17191), .C2(n16949), .A(n16948), .B(n16947), .ZN(
        n16955) );
  AOI22_X1 U20158 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9800), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16953) );
  AOI22_X1 U20159 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16952) );
  AOI22_X1 U20160 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16951) );
  NAND2_X1 U20161 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n16950) );
  NAND4_X1 U20162 ( .A1(n16953), .A2(n16952), .A3(n16951), .A4(n16950), .ZN(
        n16954) );
  AOI211_X1 U20163 ( .C1(n17043), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n16955), .B(n16954), .ZN(n16956) );
  OAI211_X1 U20164 ( .C1(n17193), .C2(n17011), .A(n16957), .B(n16956), .ZN(
        n16977) );
  NAND2_X1 U20165 ( .A1(n16978), .A2(n16977), .ZN(n16976) );
  AOI22_X1 U20166 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17214), .ZN(n16969) );
  AOI22_X1 U20167 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17200), .ZN(n16968) );
  AOI22_X1 U20168 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16967) );
  OAI22_X1 U20169 ( .A1(n10239), .A2(n16959), .B1(n16958), .B2(n10240), .ZN(
        n16965) );
  AOI22_X1 U20170 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n17194), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n9800), .ZN(n16963) );
  AOI22_X1 U20171 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17063), .ZN(n16962) );
  AOI22_X1 U20172 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16961) );
  NAND2_X1 U20173 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17175), .ZN(
        n16960) );
  NAND4_X1 U20174 ( .A1(n16963), .A2(n16962), .A3(n16961), .A4(n16960), .ZN(
        n16964) );
  AOI211_X1 U20175 ( .C1(n17219), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n16965), .B(n16964), .ZN(n16966) );
  NAND4_X1 U20176 ( .A1(n16969), .A2(n16968), .A3(n16967), .A4(n16966), .ZN(
        n16970) );
  XNOR2_X1 U20177 ( .A(n16976), .B(n16970), .ZN(n17285) );
  AOI211_X1 U20178 ( .C1(n16973), .C2(n16972), .A(n16971), .B(n17275), .ZN(
        n16974) );
  AOI21_X1 U20179 ( .B1(n17275), .B2(n17285), .A(n16974), .ZN(n16975) );
  INV_X1 U20180 ( .A(n16975), .ZN(P3_U2673) );
  OAI21_X1 U20181 ( .B1(n16978), .B2(n16977), .A(n16976), .ZN(n17294) );
  NAND2_X1 U20182 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16979), .ZN(n16983) );
  NAND4_X1 U20183 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16997), .A3(n16981), 
        .A4(n16980), .ZN(n16982) );
  OAI211_X1 U20184 ( .C1(n17266), .C2(n17294), .A(n16983), .B(n16982), .ZN(
        P3_U2674) );
  OAI21_X1 U20185 ( .B1(n16988), .B2(n16985), .A(n16984), .ZN(n17303) );
  NAND3_X1 U20186 ( .A1(n16991), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17266), 
        .ZN(n16986) );
  OAI221_X1 U20187 ( .B1(n16991), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17266), 
        .C2(n17303), .A(n16986), .ZN(P3_U2676) );
  AOI21_X1 U20188 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17266), .A(n16997), .ZN(
        n16987) );
  INV_X1 U20189 ( .A(n16987), .ZN(n16990) );
  AOI21_X1 U20190 ( .B1(n16989), .B2(n16994), .A(n16988), .ZN(n17304) );
  AOI22_X1 U20191 ( .A1(n16991), .A2(n16990), .B1(n17304), .B2(n17275), .ZN(
        n16992) );
  INV_X1 U20192 ( .A(n16992), .ZN(P3_U2677) );
  INV_X1 U20193 ( .A(n16993), .ZN(n17002) );
  AOI21_X1 U20194 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17266), .A(n17002), .ZN(
        n16996) );
  OAI21_X1 U20195 ( .B1(n16998), .B2(n16995), .A(n16994), .ZN(n17313) );
  OAI22_X1 U20196 ( .A1(n16997), .A2(n16996), .B1(n17313), .B2(n17266), .ZN(
        P3_U2678) );
  AOI21_X1 U20197 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17266), .A(n17008), .ZN(
        n17001) );
  AOI21_X1 U20198 ( .B1(n16999), .B2(n17004), .A(n16998), .ZN(n17314) );
  INV_X1 U20199 ( .A(n17314), .ZN(n17000) );
  OAI22_X1 U20200 ( .A1(n17002), .A2(n17001), .B1(n17000), .B2(n17266), .ZN(
        P3_U2679) );
  NOR2_X1 U20201 ( .A1(n17003), .A2(n17009), .ZN(n17024) );
  AOI21_X1 U20202 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17266), .A(n17024), .ZN(
        n17007) );
  OAI21_X1 U20203 ( .B1(n17006), .B2(n17005), .A(n17004), .ZN(n17323) );
  OAI22_X1 U20204 ( .A1(n17008), .A2(n17007), .B1(n17323), .B2(n17266), .ZN(
        P3_U2680) );
  INV_X1 U20205 ( .A(n17009), .ZN(n17010) );
  AOI21_X1 U20206 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17266), .A(n17010), .ZN(
        n17023) );
  AOI22_X1 U20207 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20208 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17020) );
  AOI22_X1 U20209 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17019) );
  OAI22_X1 U20210 ( .A1(n17193), .A2(n17251), .B1(n17227), .B2(n17011), .ZN(
        n17017) );
  AOI22_X1 U20211 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20212 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20213 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17013) );
  NAND2_X1 U20214 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n17012) );
  NAND4_X1 U20215 ( .A1(n17015), .A2(n17014), .A3(n17013), .A4(n17012), .ZN(
        n17016) );
  AOI211_X1 U20216 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17017), .B(n17016), .ZN(n17018) );
  NAND4_X1 U20217 ( .A1(n17021), .A2(n17020), .A3(n17019), .A4(n17018), .ZN(
        n17324) );
  INV_X1 U20218 ( .A(n17324), .ZN(n17022) );
  OAI22_X1 U20219 ( .A1(n17024), .A2(n17023), .B1(n17022), .B2(n17266), .ZN(
        P3_U2681) );
  AOI22_X1 U20220 ( .A1(n9799), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17025) );
  OAI21_X1 U20221 ( .B1(n12780), .B2(n17026), .A(n17025), .ZN(n17037) );
  AOI22_X1 U20222 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20223 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17027) );
  OAI21_X1 U20224 ( .B1(n17227), .B2(n17028), .A(n17027), .ZN(n17033) );
  AOI22_X1 U20225 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20226 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17029) );
  OAI211_X1 U20227 ( .C1(n17216), .C2(n17031), .A(n17030), .B(n17029), .ZN(
        n17032) );
  AOI211_X1 U20228 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n17033), .B(n17032), .ZN(n17034) );
  OAI211_X1 U20229 ( .C1(n17193), .C2(n17253), .A(n17035), .B(n17034), .ZN(
        n17036) );
  AOI211_X1 U20230 ( .C1(n17223), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n17037), .B(n17036), .ZN(n17332) );
  AND2_X1 U20231 ( .A1(n17266), .A2(n17038), .ZN(n17056) );
  AOI22_X1 U20232 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17056), .B1(n17040), 
        .B2(n17039), .ZN(n17041) );
  OAI21_X1 U20233 ( .B1(n17332), .B2(n17266), .A(n17041), .ZN(P3_U2682) );
  AOI22_X1 U20234 ( .A1(n9800), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17042) );
  OAI21_X1 U20235 ( .B1(n10239), .B2(n17149), .A(n17042), .ZN(n17053) );
  AOI22_X1 U20236 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17051) );
  AOI22_X1 U20237 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17044) );
  OAI21_X1 U20238 ( .B1(n17218), .B2(n17140), .A(n17044), .ZN(n17049) );
  INV_X1 U20239 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17047) );
  AOI22_X1 U20240 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20241 ( .A1(n17219), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17045) );
  OAI211_X1 U20242 ( .C1(n17191), .C2(n17047), .A(n17046), .B(n17045), .ZN(
        n17048) );
  AOI211_X1 U20243 ( .C1(n17175), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17049), .B(n17048), .ZN(n17050) );
  OAI211_X1 U20244 ( .C1(n17193), .C2(n17261), .A(n17051), .B(n17050), .ZN(
        n17052) );
  AOI211_X1 U20245 ( .C1(n17223), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n17053), .B(n17052), .ZN(n17340) );
  INV_X1 U20246 ( .A(n17055), .ZN(n17057) );
  OAI21_X1 U20247 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17057), .A(n17056), .ZN(
        n17058) );
  OAI21_X1 U20248 ( .B1(n17340), .B2(n17266), .A(n17058), .ZN(P3_U2683) );
  OAI21_X1 U20249 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17059), .A(n17266), .ZN(
        n17073) );
  AOI22_X1 U20250 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17060) );
  OAI21_X1 U20251 ( .B1(n9849), .B2(n17061), .A(n17060), .ZN(n17072) );
  INV_X1 U20252 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20253 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20254 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17062) );
  OAI21_X1 U20255 ( .B1(n17193), .B2(n17263), .A(n17062), .ZN(n17068) );
  AOI22_X1 U20256 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20257 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17064) );
  OAI211_X1 U20258 ( .C1(n17227), .C2(n17066), .A(n17065), .B(n17064), .ZN(
        n17067) );
  AOI211_X1 U20259 ( .C1(n17206), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n17068), .B(n17067), .ZN(n17069) );
  OAI211_X1 U20260 ( .C1(n12737), .C2(n17158), .A(n17070), .B(n17069), .ZN(
        n17071) );
  AOI211_X1 U20261 ( .C1(n15615), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17072), .B(n17071), .ZN(n17344) );
  OAI22_X1 U20262 ( .A1(n17074), .A2(n17073), .B1(n17344), .B2(n17266), .ZN(
        P3_U2684) );
  NAND2_X1 U20263 ( .A1(n17266), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20264 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17220), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20265 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17076) );
  AOI22_X1 U20266 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17075) );
  OAI211_X1 U20267 ( .C1(n17218), .C2(n17174), .A(n17076), .B(n17075), .ZN(
        n17082) );
  AOI22_X1 U20268 ( .A1(n9800), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17080) );
  AOI22_X1 U20269 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20270 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17078) );
  NAND2_X1 U20271 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n17077) );
  NAND4_X1 U20272 ( .A1(n17080), .A2(n17079), .A3(n17078), .A4(n17077), .ZN(
        n17081) );
  AOI211_X1 U20273 ( .C1(n17043), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17082), .B(n17081), .ZN(n17083) );
  OAI211_X1 U20274 ( .C1(n12737), .C2(n17186), .A(n17084), .B(n17083), .ZN(
        n17345) );
  NOR4_X1 U20275 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17085), .A3(n17103), .A4(
        n17272), .ZN(n17086) );
  AOI21_X1 U20276 ( .B1(n17275), .B2(n17345), .A(n17086), .ZN(n17087) );
  OAI21_X1 U20277 ( .B1(n17089), .B2(n17088), .A(n17087), .ZN(P3_U2685) );
  AOI22_X1 U20278 ( .A1(n17090), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17091) );
  OAI21_X1 U20279 ( .B1(n12737), .B2(n17192), .A(n17091), .ZN(n17102) );
  AOI22_X1 U20280 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17100) );
  OAI22_X1 U20281 ( .A1(n10240), .A2(n17093), .B1(n9849), .B2(n17092), .ZN(
        n17098) );
  AOI22_X1 U20282 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20283 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U20284 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17043), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17094) );
  NAND3_X1 U20285 ( .A1(n17096), .A2(n17095), .A3(n17094), .ZN(n17097) );
  AOI211_X1 U20286 ( .C1(n17195), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n17098), .B(n17097), .ZN(n17099) );
  OAI211_X1 U20287 ( .C1(n17193), .C2(n17270), .A(n17100), .B(n17099), .ZN(
        n17101) );
  AOI211_X1 U20288 ( .C1(n9803), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n17102), .B(n17101), .ZN(n17355) );
  NOR2_X1 U20289 ( .A1(n17103), .A2(n17272), .ZN(n17106) );
  NAND2_X1 U20290 ( .A1(n17402), .A2(n17103), .ZN(n17122) );
  INV_X1 U20291 ( .A(n17122), .ZN(n17105) );
  INV_X1 U20292 ( .A(n17257), .ZN(n17278) );
  NAND2_X1 U20293 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17278), .ZN(n17104) );
  OAI22_X1 U20294 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17106), .B1(n17105), 
        .B2(n17104), .ZN(n17107) );
  OAI21_X1 U20295 ( .B1(n17355), .B2(n17266), .A(n17107), .ZN(P3_U2686) );
  NAND2_X1 U20296 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17136), .ZN(n17121) );
  AOI22_X1 U20297 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17108) );
  OAI21_X1 U20298 ( .B1(n9849), .B2(n17109), .A(n17108), .ZN(n17119) );
  AOI22_X1 U20299 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20300 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17110) );
  OAI21_X1 U20301 ( .B1(n17227), .B2(n17217), .A(n17110), .ZN(n17115) );
  AOI22_X1 U20302 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20303 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17111) );
  OAI211_X1 U20304 ( .C1(n17216), .C2(n17113), .A(n17112), .B(n17111), .ZN(
        n17114) );
  AOI211_X1 U20305 ( .C1(n17206), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17115), .B(n17114), .ZN(n17116) );
  OAI211_X1 U20306 ( .C1(n12780), .C2(n17215), .A(n17117), .B(n17116), .ZN(
        n17118) );
  AOI211_X1 U20307 ( .C1(n15615), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17119), .B(n17118), .ZN(n17361) );
  INV_X1 U20308 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17120) );
  NAND2_X1 U20309 ( .A1(n17266), .A2(n17121), .ZN(n17137) );
  OAI222_X1 U20310 ( .A1(n17122), .A2(n17121), .B1(n17266), .B2(n17361), .C1(
        n17120), .C2(n17137), .ZN(P3_U2687) );
  AOI22_X1 U20311 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17194), .ZN(n17123) );
  OAI21_X1 U20312 ( .B1(n12780), .B2(n17124), .A(n17123), .ZN(n17135) );
  AOI22_X1 U20313 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17222), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20314 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17125) );
  OAI21_X1 U20315 ( .B1(n17247), .B2(n17227), .A(n17125), .ZN(n17130) );
  AOI22_X1 U20316 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17219), .ZN(n17127) );
  AOI22_X1 U20317 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9800), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17126) );
  OAI211_X1 U20318 ( .C1(n17128), .C2(n17216), .A(n17127), .B(n17126), .ZN(
        n17129) );
  AOI211_X1 U20319 ( .C1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .C2(n17206), .A(
        n17130), .B(n17129), .ZN(n17131) );
  OAI211_X1 U20320 ( .C1(n17133), .C2(n10239), .A(n17132), .B(n17131), .ZN(
        n17134) );
  AOI211_X1 U20321 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n17135), .B(n17134), .ZN(n17366) );
  NOR2_X1 U20322 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17136), .ZN(n17138) );
  OAI22_X1 U20323 ( .A1(n17366), .A2(n17266), .B1(n17138), .B2(n17137), .ZN(
        P3_U2688) );
  AOI22_X1 U20324 ( .A1(n9800), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17139) );
  OAI21_X1 U20325 ( .B1(n12697), .B2(n17140), .A(n17139), .ZN(n17152) );
  AOI22_X1 U20326 ( .A1(n17196), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17148) );
  OAI22_X1 U20327 ( .A1(n17193), .A2(n17141), .B1(n17227), .B2(n17261), .ZN(
        n17146) );
  AOI22_X1 U20328 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17144) );
  AOI22_X1 U20329 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20330 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17142) );
  NAND3_X1 U20331 ( .A1(n17144), .A2(n17143), .A3(n17142), .ZN(n17145) );
  AOI211_X1 U20332 ( .C1(n17229), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17146), .B(n17145), .ZN(n17147) );
  OAI211_X1 U20333 ( .C1(n17150), .C2(n17149), .A(n17148), .B(n17147), .ZN(
        n17151) );
  AOI211_X1 U20334 ( .C1(n17153), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n17152), .B(n17151), .ZN(n17379) );
  NAND3_X1 U20335 ( .A1(n17155), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17266), 
        .ZN(n17154) );
  OAI221_X1 U20336 ( .B1(n17155), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17266), 
        .C2(n17379), .A(n17154), .ZN(P3_U2691) );
  AOI22_X1 U20337 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17156) );
  OAI21_X1 U20338 ( .B1(n12737), .B2(n17157), .A(n17156), .ZN(n17168) );
  INV_X1 U20339 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17166) );
  AOI22_X1 U20340 ( .A1(n17235), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17165) );
  OAI22_X1 U20341 ( .A1(n17193), .A2(n17158), .B1(n17227), .B2(n17263), .ZN(
        n17163) );
  AOI22_X1 U20342 ( .A1(n12723), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20343 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20344 ( .A1(n17206), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17229), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17159) );
  NAND3_X1 U20345 ( .A1(n17161), .A2(n17160), .A3(n17159), .ZN(n17162) );
  AOI211_X1 U20346 ( .C1(n17175), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17163), .B(n17162), .ZN(n17164) );
  OAI211_X1 U20347 ( .C1(n12697), .C2(n17166), .A(n17165), .B(n17164), .ZN(
        n17167) );
  AOI211_X1 U20348 ( .C1(n9803), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17168), .B(n17167), .ZN(n17383) );
  INV_X1 U20349 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17189) );
  NOR2_X1 U20350 ( .A1(n17189), .A2(n17172), .ZN(n17170) );
  OAI22_X1 U20351 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17170), .B1(n17169), 
        .B2(n17172), .ZN(n17171) );
  AOI22_X1 U20352 ( .A1(n17275), .A2(n17383), .B1(n17171), .B2(n17266), .ZN(
        P3_U2692) );
  NAND2_X1 U20353 ( .A1(n17266), .A2(n17172), .ZN(n17212) );
  AOI22_X1 U20354 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15615), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20355 ( .A1(n17200), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17221), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17173) );
  OAI21_X1 U20356 ( .B1(n12697), .B2(n17174), .A(n17173), .ZN(n17183) );
  AOI22_X1 U20357 ( .A1(n17175), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17181) );
  INV_X1 U20358 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20359 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17177) );
  AOI22_X1 U20360 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17176) );
  OAI211_X1 U20361 ( .C1(n17218), .C2(n17178), .A(n17177), .B(n17176), .ZN(
        n17179) );
  AOI21_X1 U20362 ( .B1(n17229), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17179), .ZN(n17180) );
  OAI211_X1 U20363 ( .C1(n17227), .C2(n17267), .A(n17181), .B(n17180), .ZN(
        n17182) );
  AOI211_X1 U20364 ( .C1(n9800), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17183), .B(n17182), .ZN(n17184) );
  OAI211_X1 U20365 ( .C1(n17193), .C2(n17186), .A(n17185), .B(n17184), .ZN(
        n17387) );
  AOI22_X1 U20366 ( .A1(n17275), .A2(n17387), .B1(n17187), .B2(n17189), .ZN(
        n17188) );
  OAI21_X1 U20367 ( .B1(n17189), .B2(n17212), .A(n17188), .ZN(P3_U2693) );
  OAI22_X1 U20368 ( .A1(n17193), .A2(n17192), .B1(n17191), .B2(n17190), .ZN(
        n17211) );
  AOI22_X1 U20369 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20370 ( .A1(n17195), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20371 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17196), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17197) );
  OAI21_X1 U20372 ( .B1(n17199), .B2(n17198), .A(n17197), .ZN(n17205) );
  AOI22_X1 U20373 ( .A1(n9799), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17200), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17203) );
  AOI22_X1 U20374 ( .A1(n17201), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17202) );
  OAI211_X1 U20375 ( .C1(n17227), .C2(n17270), .A(n17203), .B(n17202), .ZN(
        n17204) );
  AOI211_X1 U20376 ( .C1(n17206), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n17205), .B(n17204), .ZN(n17207) );
  NAND3_X1 U20377 ( .A1(n17209), .A2(n17208), .A3(n17207), .ZN(n17210) );
  AOI211_X1 U20378 ( .C1(n17175), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n17211), .B(n17210), .ZN(n17392) );
  NOR2_X1 U20379 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17242), .ZN(n17213) );
  OAI22_X1 U20380 ( .A1(n17392), .A2(n17266), .B1(n17213), .B2(n17212), .ZN(
        P3_U2694) );
  AOI22_X1 U20381 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17063), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20382 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17214), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17237) );
  OAI22_X1 U20383 ( .A1(n17218), .A2(n17217), .B1(n17216), .B2(n17215), .ZN(
        n17234) );
  AOI22_X1 U20384 ( .A1(n17220), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17219), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U20385 ( .A1(n15615), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17194), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20386 ( .A1(n17223), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9799), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17224) );
  OAI211_X1 U20387 ( .C1(n17227), .C2(n17226), .A(n17225), .B(n17224), .ZN(
        n17228) );
  AOI21_X1 U20388 ( .B1(n17229), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17228), .ZN(n17230) );
  OAI211_X1 U20389 ( .C1(n9849), .C2(n17232), .A(n17231), .B(n17230), .ZN(
        n17233) );
  AOI211_X1 U20390 ( .C1(n17235), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n17234), .B(n17233), .ZN(n17236) );
  NAND3_X1 U20391 ( .A1(n17238), .A2(n17237), .A3(n17236), .ZN(n17397) );
  INV_X1 U20392 ( .A(n17397), .ZN(n17243) );
  NOR2_X1 U20393 ( .A1(n18272), .A2(n17239), .ZN(n17240) );
  AOI21_X1 U20394 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17266), .A(n17240), .ZN(
        n17241) );
  OAI22_X1 U20395 ( .A1(n17243), .A2(n17266), .B1(n17242), .B2(n17241), .ZN(
        P3_U2695) );
  NAND3_X1 U20396 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17252), .ZN(n17249) );
  OAI21_X1 U20397 ( .B1(n17275), .B2(n17245), .A(n17249), .ZN(n17244) );
  OAI221_X1 U20398 ( .B1(n17402), .B2(n17249), .C1(n17249), .C2(n17245), .A(
        n17244), .ZN(n17246) );
  OAI21_X1 U20399 ( .B1(n17247), .B2(n17266), .A(n17246), .ZN(P3_U2696) );
  INV_X1 U20400 ( .A(n17252), .ZN(n17258) );
  NOR2_X1 U20401 ( .A1(n17248), .A2(n17258), .ZN(n17255) );
  OAI211_X1 U20402 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17255), .A(n17249), .B(
        n17266), .ZN(n17250) );
  OAI21_X1 U20403 ( .B1(n17266), .B2(n17251), .A(n17250), .ZN(P3_U2697) );
  OAI21_X1 U20404 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17252), .A(n17266), .ZN(
        n17254) );
  OAI22_X1 U20405 ( .A1(n17255), .A2(n17254), .B1(n17253), .B2(n17266), .ZN(
        P3_U2698) );
  NOR2_X1 U20406 ( .A1(n17257), .A2(n17256), .ZN(n17259) );
  OAI21_X1 U20407 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17259), .A(n17258), .ZN(
        n17260) );
  AOI22_X1 U20408 ( .A1(n17275), .A2(n17261), .B1(n17260), .B2(n17266), .ZN(
        P3_U2699) );
  NAND3_X1 U20409 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17264), .A3(n17274), .ZN(
        n17265) );
  NAND3_X1 U20410 ( .A1(n17265), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17266), .ZN(
        n17262) );
  OAI221_X1 U20411 ( .B1(n17265), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17266), 
        .C2(n17263), .A(n17262), .ZN(P3_U2700) );
  AOI21_X1 U20412 ( .B1(n17278), .B2(n17264), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17269) );
  NAND2_X1 U20413 ( .A1(n17266), .A2(n17265), .ZN(n17268) );
  OAI22_X1 U20414 ( .A1(n17269), .A2(n17268), .B1(n17267), .B2(n17266), .ZN(
        P3_U2701) );
  OAI222_X1 U20415 ( .A1(n17273), .A2(n17272), .B1(n17271), .B2(n17278), .C1(
        n17270), .C2(n17266), .ZN(P3_U2702) );
  AOI22_X1 U20416 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17275), .B1(
        n17274), .B2(n17277), .ZN(n17276) );
  OAI21_X1 U20417 ( .B1(n17278), .B2(n17277), .A(n17276), .ZN(P3_U2703) );
  INV_X1 U20418 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17498) );
  INV_X1 U20419 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17495) );
  INV_X1 U20420 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17506) );
  INV_X1 U20421 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17510) );
  INV_X1 U20422 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17508) );
  NAND4_X1 U20423 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n17280) );
  NOR3_X1 U20424 ( .A1(n17510), .A2(n17508), .A3(n17280), .ZN(n17368) );
  INV_X1 U20425 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17520) );
  NAND2_X1 U20426 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .ZN(n17374) );
  NOR2_X1 U20427 ( .A1(n17520), .A2(n17374), .ZN(n17281) );
  NAND4_X1 U20428 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(n17281), .ZN(n17369) );
  INV_X1 U20429 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17539) );
  NAND2_X1 U20430 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n17325) );
  NAND2_X1 U20431 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17316), .ZN(n17315) );
  NAND2_X1 U20432 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17296), .ZN(n17291) );
  INV_X1 U20433 ( .A(n17291), .ZN(n17287) );
  NAND2_X1 U20434 ( .A1(n17287), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17284) );
  NAND2_X1 U20435 ( .A1(n18267), .A2(n17428), .ZN(n17331) );
  NAND2_X1 U20436 ( .A1(n17422), .A2(n17291), .ZN(n17290) );
  OAI21_X1 U20437 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17326), .A(n17290), .ZN(
        n17282) );
  AOI22_X1 U20438 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17356), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17282), .ZN(n17283) );
  OAI21_X1 U20439 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17284), .A(n17283), .ZN(
        P3_U2704) );
  INV_X1 U20440 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17502) );
  AOI22_X1 U20441 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n17356), .B1(n17424), .B2(
        n17285), .ZN(n17289) );
  NAND2_X1 U20442 ( .A1(n17286), .A2(n17428), .ZN(n17350) );
  AOI22_X1 U20443 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17357), .B1(n17287), .B2(
        n17502), .ZN(n17288) );
  OAI211_X1 U20444 ( .C1(n17290), .C2(n17502), .A(n17289), .B(n17288), .ZN(
        P3_U2705) );
  AOI22_X1 U20445 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17356), .ZN(n17293) );
  OAI211_X1 U20446 ( .C1(n17296), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17422), .B(
        n17291), .ZN(n17292) );
  OAI211_X1 U20447 ( .C1(n17294), .C2(n17433), .A(n17293), .B(n17292), .ZN(
        P3_U2706) );
  INV_X1 U20448 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U20449 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n17356), .B1(n17424), .B2(
        n17295), .ZN(n17299) );
  AOI211_X1 U20450 ( .C1(n17498), .C2(n17300), .A(n17296), .B(n17428), .ZN(
        n17297) );
  INV_X1 U20451 ( .A(n17297), .ZN(n17298) );
  OAI211_X1 U20452 ( .C1(n17350), .C2(n17382), .A(n17299), .B(n17298), .ZN(
        P3_U2707) );
  AOI22_X1 U20453 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17356), .ZN(n17302) );
  OAI211_X1 U20454 ( .C1(n9878), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17422), .B(
        n17300), .ZN(n17301) );
  OAI211_X1 U20455 ( .C1(n17303), .C2(n17433), .A(n17302), .B(n17301), .ZN(
        P3_U2708) );
  INV_X1 U20456 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20457 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n17356), .B1(n17424), .B2(
        n17304), .ZN(n17307) );
  AOI211_X1 U20458 ( .C1(n17495), .C2(n17309), .A(n9878), .B(n17428), .ZN(
        n17305) );
  INV_X1 U20459 ( .A(n17305), .ZN(n17306) );
  OAI211_X1 U20460 ( .C1(n17350), .C2(n17308), .A(n17307), .B(n17306), .ZN(
        P3_U2709) );
  AOI22_X1 U20461 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17356), .ZN(n17312) );
  OAI211_X1 U20462 ( .C1(n17310), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17422), .B(
        n17309), .ZN(n17311) );
  OAI211_X1 U20463 ( .C1(n17313), .C2(n17433), .A(n17312), .B(n17311), .ZN(
        P3_U2710) );
  INV_X1 U20464 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U20465 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n17356), .B1(n17424), .B2(
        n17314), .ZN(n17318) );
  OAI211_X1 U20466 ( .C1(n17316), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17422), .B(
        n17315), .ZN(n17317) );
  OAI211_X1 U20467 ( .C1(n17350), .C2(n17401), .A(n17318), .B(n17317), .ZN(
        P3_U2711) );
  AOI22_X1 U20468 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17356), .ZN(n17322) );
  OAI211_X1 U20469 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17320), .A(n17422), .B(
        n17319), .ZN(n17321) );
  OAI211_X1 U20470 ( .C1(n17323), .C2(n17433), .A(n17322), .B(n17321), .ZN(
        P3_U2712) );
  AOI22_X1 U20471 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17356), .B1(n17424), .B2(
        n17324), .ZN(n17330) );
  NAND2_X1 U20472 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17346), .ZN(n17341) );
  NAND2_X1 U20473 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17337), .ZN(n17336) );
  NAND2_X1 U20474 ( .A1(n17422), .A2(n17336), .ZN(n17335) );
  OAI21_X1 U20475 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17326), .A(n17335), .ZN(
        n17328) );
  NOR2_X1 U20476 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17336), .ZN(n17327) );
  AOI22_X1 U20477 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17328), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17327), .ZN(n17329) );
  OAI211_X1 U20478 ( .C1(n18269), .C2(n17350), .A(n17330), .B(n17329), .ZN(
        P3_U2713) );
  INV_X1 U20479 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17486) );
  INV_X1 U20480 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19279) );
  OAI22_X1 U20481 ( .A1(n17332), .A2(n17433), .B1(n19279), .B2(n17331), .ZN(
        n17333) );
  AOI21_X1 U20482 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17357), .A(n17333), .ZN(
        n17334) );
  OAI221_X1 U20483 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17336), .C1(n17486), 
        .C2(n17335), .A(n17334), .ZN(P3_U2714) );
  AOI22_X1 U20484 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17356), .ZN(n17339) );
  OAI211_X1 U20485 ( .C1(n17337), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17422), .B(
        n17336), .ZN(n17338) );
  OAI211_X1 U20486 ( .C1(n17340), .C2(n17433), .A(n17339), .B(n17338), .ZN(
        P3_U2715) );
  AOI22_X1 U20487 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17356), .ZN(n17343) );
  OAI211_X1 U20488 ( .C1(n17346), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17422), .B(
        n17341), .ZN(n17342) );
  OAI211_X1 U20489 ( .C1(n17344), .C2(n17433), .A(n17343), .B(n17342), .ZN(
        P3_U2716) );
  INV_X1 U20490 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18249) );
  AOI22_X1 U20491 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17356), .B1(n17424), .B2(
        n17345), .ZN(n17349) );
  INV_X1 U20492 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17480) );
  INV_X1 U20493 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17478) );
  OR2_X1 U20494 ( .A1(n17478), .A2(n17358), .ZN(n17351) );
  AOI211_X1 U20495 ( .C1(n17480), .C2(n17351), .A(n17346), .B(n17428), .ZN(
        n17347) );
  INV_X1 U20496 ( .A(n17347), .ZN(n17348) );
  OAI211_X1 U20497 ( .C1(n17350), .C2(n18249), .A(n17349), .B(n17348), .ZN(
        P3_U2717) );
  AOI22_X1 U20498 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17356), .ZN(n17354) );
  INV_X1 U20499 ( .A(n17358), .ZN(n17352) );
  OAI211_X1 U20500 ( .C1(n17352), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17422), .B(
        n17351), .ZN(n17353) );
  OAI211_X1 U20501 ( .C1(n17355), .C2(n17433), .A(n17354), .B(n17353), .ZN(
        P3_U2718) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17357), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17356), .ZN(n17360) );
  OAI211_X1 U20503 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17362), .A(n17422), .B(
        n17358), .ZN(n17359) );
  OAI211_X1 U20504 ( .C1(n17361), .C2(n17433), .A(n17360), .B(n17359), .ZN(
        P3_U2719) );
  AOI21_X1 U20505 ( .B1(n17539), .B2(n17363), .A(n17362), .ZN(n17364) );
  AOI22_X1 U20506 ( .A1(n17431), .A2(BUF2_REG_15__SCAN_IN), .B1(n17364), .B2(
        n17422), .ZN(n17365) );
  OAI21_X1 U20507 ( .B1(n17366), .B2(n17433), .A(n17365), .ZN(P3_U2720) );
  INV_X1 U20508 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17534) );
  NOR3_X1 U20509 ( .A1(n17428), .A2(n17367), .A3(n17534), .ZN(n17371) );
  NAND3_X1 U20510 ( .A1(n17402), .A2(n9874), .A3(n17368), .ZN(n17396) );
  NOR3_X1 U20511 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17369), .A3(n17396), .ZN(
        n17370) );
  AOI211_X1 U20512 ( .C1(n17431), .C2(BUF2_REG_14__SCAN_IN), .A(n17371), .B(
        n17370), .ZN(n17372) );
  OAI21_X1 U20513 ( .B1(n17373), .B2(n17433), .A(n17372), .ZN(P3_U2721) );
  NOR2_X1 U20514 ( .A1(n17520), .A2(n17396), .ZN(n17391) );
  NAND2_X1 U20515 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17391), .ZN(n17388) );
  NOR2_X1 U20516 ( .A1(n17374), .A2(n17388), .ZN(n17385) );
  NAND2_X1 U20517 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17385), .ZN(n17378) );
  NAND3_X1 U20518 ( .A1(n17422), .A2(P3_EAX_REG_13__SCAN_IN), .A3(n17378), 
        .ZN(n17377) );
  AOI22_X1 U20519 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17431), .B1(n17424), .B2(
        n17375), .ZN(n17376) );
  OAI211_X1 U20520 ( .C1(P3_EAX_REG_13__SCAN_IN), .C2(n17378), .A(n17377), .B(
        n17376), .ZN(P3_U2722) );
  INV_X1 U20521 ( .A(n17378), .ZN(n17381) );
  AOI21_X1 U20522 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17422), .A(n17385), .ZN(
        n17380) );
  OAI222_X1 U20523 ( .A1(n17421), .A2(n17382), .B1(n17381), .B2(n17380), .C1(
        n17433), .C2(n17379), .ZN(P3_U2723) );
  INV_X1 U20524 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17386) );
  INV_X1 U20525 ( .A(n17388), .ZN(n17394) );
  AOI22_X1 U20526 ( .A1(n17394), .A2(P3_EAX_REG_10__SCAN_IN), .B1(
        P3_EAX_REG_11__SCAN_IN), .B2(n17422), .ZN(n17384) );
  OAI222_X1 U20527 ( .A1(n17421), .A2(n17386), .B1(n17385), .B2(n17384), .C1(
        n17433), .C2(n17383), .ZN(P3_U2724) );
  AOI22_X1 U20528 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17431), .B1(n17424), .B2(
        n17387), .ZN(n17390) );
  INV_X1 U20529 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17524) );
  OAI221_X1 U20530 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n17394), .C1(n17524), 
        .C2(n17388), .A(n17422), .ZN(n17389) );
  NAND2_X1 U20531 ( .A1(n17390), .A2(n17389), .ZN(P3_U2725) );
  INV_X1 U20532 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17395) );
  AOI21_X1 U20533 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17422), .A(n17391), .ZN(
        n17393) );
  OAI222_X1 U20534 ( .A1(n17421), .A2(n17395), .B1(n17394), .B2(n17393), .C1(
        n17433), .C2(n17392), .ZN(P3_U2726) );
  INV_X1 U20535 ( .A(n17396), .ZN(n17406) );
  AOI22_X1 U20536 ( .A1(n17424), .A2(n17397), .B1(n17406), .B2(n17520), .ZN(
        n17400) );
  NAND3_X1 U20537 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17422), .A3(n17398), .ZN(
        n17399) );
  OAI211_X1 U20538 ( .C1(n17421), .C2(n17401), .A(n17400), .B(n17399), .ZN(
        P3_U2727) );
  INV_X1 U20539 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18274) );
  INV_X1 U20540 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17516) );
  INV_X1 U20541 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17512) );
  NAND2_X1 U20542 ( .A1(n17402), .A2(n9874), .ZN(n17403) );
  NAND2_X1 U20543 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17427), .ZN(n17414) );
  NOR2_X1 U20544 ( .A1(n17512), .A2(n17414), .ZN(n17417) );
  NAND2_X1 U20545 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17417), .ZN(n17407) );
  NOR2_X1 U20546 ( .A1(n17516), .A2(n17407), .ZN(n17409) );
  AOI21_X1 U20547 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17422), .A(n17409), .ZN(
        n17405) );
  OAI222_X1 U20548 ( .A1(n17421), .A2(n18274), .B1(n17406), .B2(n17405), .C1(
        n17433), .C2(n17404), .ZN(P3_U2728) );
  INV_X1 U20549 ( .A(n17407), .ZN(n17413) );
  AOI21_X1 U20550 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17422), .A(n17413), .ZN(
        n17410) );
  OAI222_X1 U20551 ( .A1(n17421), .A2(n18269), .B1(n17410), .B2(n17409), .C1(
        n17433), .C2(n17408), .ZN(P3_U2729) );
  INV_X1 U20552 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18263) );
  AOI21_X1 U20553 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17422), .A(n17417), .ZN(
        n17412) );
  OAI222_X1 U20554 ( .A1(n18263), .A2(n17421), .B1(n17413), .B2(n17412), .C1(
        n17433), .C2(n17411), .ZN(P3_U2730) );
  INV_X1 U20555 ( .A(n17414), .ZN(n17420) );
  AOI21_X1 U20556 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17422), .A(n17420), .ZN(
        n17416) );
  OAI222_X1 U20557 ( .A1(n18259), .A2(n17421), .B1(n17417), .B2(n17416), .C1(
        n17433), .C2(n17415), .ZN(P3_U2731) );
  INV_X1 U20558 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18254) );
  AOI21_X1 U20559 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17422), .A(n17427), .ZN(
        n17419) );
  OAI222_X1 U20560 ( .A1(n18254), .A2(n17421), .B1(n17420), .B2(n17419), .C1(
        n17433), .C2(n17418), .ZN(P3_U2732) );
  OAI21_X1 U20561 ( .B1(n9874), .B2(P3_EAX_REG_2__SCAN_IN), .A(n17422), .ZN(
        n17426) );
  AOI22_X1 U20562 ( .A1(n17431), .A2(BUF2_REG_2__SCAN_IN), .B1(n17424), .B2(
        n17423), .ZN(n17425) );
  OAI21_X1 U20563 ( .B1(n17427), .B2(n17426), .A(n17425), .ZN(P3_U2733) );
  AOI211_X1 U20564 ( .C1(n17506), .C2(n17429), .A(n17428), .B(n9874), .ZN(
        n17430) );
  AOI21_X1 U20565 ( .B1(n17431), .B2(BUF2_REG_1__SCAN_IN), .A(n17430), .ZN(
        n17432) );
  OAI21_X1 U20566 ( .B1(n17434), .B2(n17433), .A(n17432), .ZN(P3_U2734) );
  OR2_X1 U20567 ( .A1(n18842), .A2(n18737), .ZN(n18879) );
  NOR2_X4 U20569 ( .A1(n18720), .A2(n17454), .ZN(n17451) );
  AND2_X1 U20570 ( .A1(n17451), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AOI22_X1 U20571 ( .A1(n18720), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17451), .ZN(n17437) );
  OAI21_X1 U20572 ( .B1(n17502), .B2(n17453), .A(n17437), .ZN(P3_U2737) );
  INV_X1 U20573 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U20574 ( .A1(n18720), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17438) );
  OAI21_X1 U20575 ( .B1(n17500), .B2(n17453), .A(n17438), .ZN(P3_U2738) );
  AOI22_X1 U20576 ( .A1(n18720), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17439) );
  OAI21_X1 U20577 ( .B1(n17498), .B2(n17453), .A(n17439), .ZN(P3_U2739) );
  AOI22_X1 U20578 ( .A1(n18720), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17440) );
  OAI21_X1 U20579 ( .B1(n10067), .B2(n17453), .A(n17440), .ZN(P3_U2740) );
  AOI22_X1 U20580 ( .A1(n18720), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17441) );
  OAI21_X1 U20581 ( .B1(n17495), .B2(n17453), .A(n17441), .ZN(P3_U2741) );
  AOI22_X1 U20582 ( .A1(n18720), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17442) );
  OAI21_X1 U20583 ( .B1(n10066), .B2(n17453), .A(n17442), .ZN(P3_U2742) );
  INV_X1 U20584 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U20585 ( .A1(n18720), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17443) );
  OAI21_X1 U20586 ( .B1(n17492), .B2(n17453), .A(n17443), .ZN(P3_U2743) );
  INV_X1 U20587 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17490) );
  AOI22_X1 U20589 ( .A1(n18720), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17444) );
  OAI21_X1 U20590 ( .B1(n17490), .B2(n17453), .A(n17444), .ZN(P3_U2744) );
  INV_X1 U20591 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U20592 ( .A1(n18720), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17445) );
  OAI21_X1 U20593 ( .B1(n17488), .B2(n17453), .A(n17445), .ZN(P3_U2745) );
  AOI22_X1 U20594 ( .A1(n18720), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17446) );
  OAI21_X1 U20595 ( .B1(n17486), .B2(n17453), .A(n17446), .ZN(P3_U2746) );
  INV_X1 U20596 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U20597 ( .A1(n18720), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20598 ( .B1(n17484), .B2(n17453), .A(n17447), .ZN(P3_U2747) );
  INV_X1 U20599 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U20600 ( .A1(n18720), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17448) );
  OAI21_X1 U20601 ( .B1(n17482), .B2(n17453), .A(n17448), .ZN(P3_U2748) );
  AOI22_X1 U20602 ( .A1(n18720), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U20603 ( .B1(n17480), .B2(n17453), .A(n17449), .ZN(P3_U2749) );
  AOI22_X1 U20604 ( .A1(n18720), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17450) );
  OAI21_X1 U20605 ( .B1(n17478), .B2(n17453), .A(n17450), .ZN(P3_U2750) );
  AOI22_X1 U20606 ( .A1(n18720), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U20607 ( .B1(n10064), .B2(n17453), .A(n17452), .ZN(P3_U2751) );
  AOI22_X1 U20608 ( .A1(n18720), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17455) );
  OAI21_X1 U20609 ( .B1(n17539), .B2(n17472), .A(n17455), .ZN(P3_U2752) );
  AOI22_X1 U20610 ( .A1(n18720), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17456) );
  OAI21_X1 U20611 ( .B1(n17534), .B2(n17472), .A(n17456), .ZN(P3_U2753) );
  INV_X1 U20612 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17532) );
  AOI22_X1 U20613 ( .A1(n18720), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17457) );
  OAI21_X1 U20614 ( .B1(n17532), .B2(n17472), .A(n17457), .ZN(P3_U2754) );
  INV_X1 U20615 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17530) );
  AOI22_X1 U20616 ( .A1(n18720), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17458) );
  OAI21_X1 U20617 ( .B1(n17530), .B2(n17472), .A(n17458), .ZN(P3_U2755) );
  INV_X1 U20618 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17526) );
  AOI22_X1 U20619 ( .A1(n18720), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U20620 ( .B1(n17526), .B2(n17472), .A(n17459), .ZN(P3_U2756) );
  AOI22_X1 U20621 ( .A1(n18720), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17460) );
  OAI21_X1 U20622 ( .B1(n17524), .B2(n17472), .A(n17460), .ZN(P3_U2757) );
  INV_X1 U20623 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17522) );
  AOI22_X1 U20624 ( .A1(n18720), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17461) );
  OAI21_X1 U20625 ( .B1(n17522), .B2(n17472), .A(n17461), .ZN(P3_U2758) );
  AOI22_X1 U20626 ( .A1(n18720), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17462) );
  OAI21_X1 U20627 ( .B1(n17520), .B2(n17472), .A(n17462), .ZN(P3_U2759) );
  INV_X1 U20628 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17518) );
  AOI22_X1 U20629 ( .A1(n18720), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17463) );
  OAI21_X1 U20630 ( .B1(n17518), .B2(n17472), .A(n17463), .ZN(P3_U2760) );
  AOI22_X1 U20631 ( .A1(n18720), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17464) );
  OAI21_X1 U20632 ( .B1(n17516), .B2(n17472), .A(n17464), .ZN(P3_U2761) );
  INV_X1 U20633 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U20634 ( .A1(n18720), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17465) );
  OAI21_X1 U20635 ( .B1(n17514), .B2(n17472), .A(n17465), .ZN(P3_U2762) );
  AOI22_X1 U20636 ( .A1(n18720), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20637 ( .B1(n17512), .B2(n17472), .A(n17466), .ZN(P3_U2763) );
  AOI22_X1 U20638 ( .A1(n18720), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17467) );
  OAI21_X1 U20639 ( .B1(n17510), .B2(n17472), .A(n17467), .ZN(P3_U2764) );
  AOI22_X1 U20640 ( .A1(n18720), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17468) );
  OAI21_X1 U20641 ( .B1(n17508), .B2(n17472), .A(n17468), .ZN(P3_U2765) );
  AOI22_X1 U20642 ( .A1(n18720), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U20643 ( .B1(n17506), .B2(n17472), .A(n17469), .ZN(P3_U2766) );
  AOI22_X1 U20644 ( .A1(n18720), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17451), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17471) );
  OAI21_X1 U20645 ( .B1(n17504), .B2(n17472), .A(n17471), .ZN(P3_U2767) );
  NAND2_X2 U20646 ( .A1(n18885), .A2(n17475), .ZN(n17538) );
  AOI22_X1 U20647 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17536), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17527), .ZN(n17476) );
  OAI21_X1 U20648 ( .B1(n10064), .B2(n17538), .A(n17476), .ZN(P3_U2768) );
  AOI22_X1 U20649 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17536), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17527), .ZN(n17477) );
  OAI21_X1 U20650 ( .B1(n17478), .B2(n17538), .A(n17477), .ZN(P3_U2769) );
  AOI22_X1 U20651 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17536), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17527), .ZN(n17479) );
  OAI21_X1 U20652 ( .B1(n17480), .B2(n17538), .A(n17479), .ZN(P3_U2770) );
  AOI22_X1 U20653 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17527), .ZN(n17481) );
  OAI21_X1 U20654 ( .B1(n17482), .B2(n17538), .A(n17481), .ZN(P3_U2771) );
  AOI22_X1 U20655 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17527), .ZN(n17483) );
  OAI21_X1 U20656 ( .B1(n17484), .B2(n17538), .A(n17483), .ZN(P3_U2772) );
  AOI22_X1 U20657 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17527), .ZN(n17485) );
  OAI21_X1 U20658 ( .B1(n17486), .B2(n17538), .A(n17485), .ZN(P3_U2773) );
  AOI22_X1 U20659 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17527), .ZN(n17487) );
  OAI21_X1 U20660 ( .B1(n17488), .B2(n17538), .A(n17487), .ZN(P3_U2774) );
  AOI22_X1 U20661 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17527), .ZN(n17489) );
  OAI21_X1 U20662 ( .B1(n17490), .B2(n17538), .A(n17489), .ZN(P3_U2775) );
  AOI22_X1 U20663 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17527), .ZN(n17491) );
  OAI21_X1 U20664 ( .B1(n17492), .B2(n17538), .A(n17491), .ZN(P3_U2776) );
  AOI22_X1 U20665 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17527), .ZN(n17493) );
  OAI21_X1 U20666 ( .B1(n10066), .B2(n17538), .A(n17493), .ZN(P3_U2777) );
  AOI22_X1 U20667 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17527), .ZN(n17494) );
  OAI21_X1 U20668 ( .B1(n17495), .B2(n17538), .A(n17494), .ZN(P3_U2778) );
  AOI22_X1 U20669 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17528), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17527), .ZN(n17496) );
  OAI21_X1 U20670 ( .B1(n10067), .B2(n17538), .A(n17496), .ZN(P3_U2779) );
  AOI22_X1 U20671 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17536), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17527), .ZN(n17497) );
  OAI21_X1 U20672 ( .B1(n17498), .B2(n17538), .A(n17497), .ZN(P3_U2780) );
  AOI22_X1 U20673 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17536), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17527), .ZN(n17499) );
  OAI21_X1 U20674 ( .B1(n17500), .B2(n17538), .A(n17499), .ZN(P3_U2781) );
  AOI22_X1 U20675 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17536), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17527), .ZN(n17501) );
  OAI21_X1 U20676 ( .B1(n17502), .B2(n17538), .A(n17501), .ZN(P3_U2782) );
  AOI22_X1 U20677 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17527), .ZN(n17503) );
  OAI21_X1 U20678 ( .B1(n17504), .B2(n17538), .A(n17503), .ZN(P3_U2783) );
  AOI22_X1 U20679 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17527), .ZN(n17505) );
  OAI21_X1 U20680 ( .B1(n17506), .B2(n17538), .A(n17505), .ZN(P3_U2784) );
  AOI22_X1 U20681 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17527), .ZN(n17507) );
  OAI21_X1 U20682 ( .B1(n17508), .B2(n17538), .A(n17507), .ZN(P3_U2785) );
  AOI22_X1 U20683 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17527), .ZN(n17509) );
  OAI21_X1 U20684 ( .B1(n17510), .B2(n17538), .A(n17509), .ZN(P3_U2786) );
  AOI22_X1 U20685 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17535), .ZN(n17511) );
  OAI21_X1 U20686 ( .B1(n17512), .B2(n17538), .A(n17511), .ZN(P3_U2787) );
  AOI22_X1 U20687 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17535), .ZN(n17513) );
  OAI21_X1 U20688 ( .B1(n17514), .B2(n17538), .A(n17513), .ZN(P3_U2788) );
  AOI22_X1 U20689 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17535), .ZN(n17515) );
  OAI21_X1 U20690 ( .B1(n17516), .B2(n17538), .A(n17515), .ZN(P3_U2789) );
  AOI22_X1 U20691 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17535), .ZN(n17517) );
  OAI21_X1 U20692 ( .B1(n17518), .B2(n17538), .A(n17517), .ZN(P3_U2790) );
  AOI22_X1 U20693 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17535), .ZN(n17519) );
  OAI21_X1 U20694 ( .B1(n17520), .B2(n17538), .A(n17519), .ZN(P3_U2791) );
  AOI22_X1 U20695 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17535), .ZN(n17521) );
  OAI21_X1 U20696 ( .B1(n17522), .B2(n17538), .A(n17521), .ZN(P3_U2792) );
  AOI22_X1 U20697 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17528), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17527), .ZN(n17523) );
  OAI21_X1 U20698 ( .B1(n17524), .B2(n17538), .A(n17523), .ZN(P3_U2793) );
  AOI22_X1 U20699 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17535), .ZN(n17525) );
  OAI21_X1 U20700 ( .B1(n17526), .B2(n17538), .A(n17525), .ZN(P3_U2794) );
  AOI22_X1 U20701 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17528), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17527), .ZN(n17529) );
  OAI21_X1 U20702 ( .B1(n17530), .B2(n17538), .A(n17529), .ZN(P3_U2795) );
  AOI22_X1 U20703 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17535), .ZN(n17531) );
  OAI21_X1 U20704 ( .B1(n17532), .B2(n17538), .A(n17531), .ZN(P3_U2796) );
  AOI22_X1 U20705 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17535), .ZN(n17533) );
  OAI21_X1 U20706 ( .B1(n17534), .B2(n17538), .A(n17533), .ZN(P3_U2797) );
  AOI22_X1 U20707 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17536), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17535), .ZN(n17537) );
  OAI21_X1 U20708 ( .B1(n17539), .B2(n17538), .A(n17537), .ZN(P3_U2798) );
  NAND2_X1 U20709 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17540), .ZN(
        n17555) );
  INV_X1 U20710 ( .A(n17696), .ZN(n17659) );
  NOR3_X1 U20711 ( .A1(n17659), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        n17543), .ZN(n17549) );
  NOR2_X1 U20712 ( .A1(n17816), .A2(n17897), .ZN(n17650) );
  OAI22_X1 U20713 ( .A1(n17914), .A2(n17730), .B1(n17913), .B2(n17908), .ZN(
        n17574) );
  NOR2_X1 U20714 ( .A1(n17923), .A2(n17574), .ZN(n17561) );
  NOR3_X1 U20715 ( .A1(n17650), .A2(n17561), .A3(n17540), .ZN(n17548) );
  NOR3_X1 U20716 ( .A1(n17659), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17543), .ZN(n17563) );
  OAI21_X1 U20717 ( .B1(n17541), .B2(n18737), .A(n17904), .ZN(n17542) );
  AOI21_X1 U20718 ( .B1(n17866), .B2(n17543), .A(n17542), .ZN(n17571) );
  OAI21_X1 U20719 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17680), .A(
        n17571), .ZN(n17557) );
  OAI21_X1 U20720 ( .B1(n17563), .B2(n17557), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17545) );
  OAI211_X1 U20721 ( .C1(n17740), .C2(n17546), .A(n17545), .B(n17544), .ZN(
        n17547) );
  AOI211_X1 U20722 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17549), .A(
        n17548), .B(n17547), .ZN(n17554) );
  OAI211_X1 U20723 ( .C1(n17552), .C2(n17551), .A(n17815), .B(n17550), .ZN(
        n17553) );
  OAI211_X1 U20724 ( .C1(n17562), .C2(n17555), .A(n17554), .B(n17553), .ZN(
        P3_U2802) );
  AOI22_X1 U20725 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17557), .B1(
        n17755), .B2(n17556), .ZN(n17564) );
  NOR2_X1 U20726 ( .A1(n17559), .A2(n17558), .ZN(n17560) );
  XOR2_X1 U20727 ( .A(n17777), .B(n17560), .Z(n17919) );
  AOI21_X1 U20728 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17566), .A(
        n17565), .ZN(n17931) );
  NOR4_X1 U20729 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17941), .A3(
        n17933), .A4(n17705), .ZN(n17573) );
  AOI21_X1 U20730 ( .B1(n18608), .B2(n9914), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17570) );
  INV_X1 U20731 ( .A(n17680), .ZN(n17568) );
  OAI21_X1 U20732 ( .B1(n17755), .B2(n17568), .A(n17567), .ZN(n17569) );
  NAND2_X1 U20733 ( .A1(n18122), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17929) );
  OAI211_X1 U20734 ( .C1(n17571), .C2(n17570), .A(n17569), .B(n17929), .ZN(
        n17572) );
  AOI211_X1 U20735 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17574), .A(
        n17573), .B(n17572), .ZN(n17575) );
  OAI21_X1 U20736 ( .B1(n17931), .B2(n17790), .A(n17575), .ZN(P3_U2804) );
  NOR2_X1 U20737 ( .A1(n18042), .A2(n17590), .ZN(n17951) );
  NAND2_X1 U20738 ( .A1(n17951), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17576) );
  XOR2_X1 U20739 ( .A(n17576), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17936) );
  OAI21_X1 U20740 ( .B1(n17577), .B2(n18737), .A(n17904), .ZN(n17578) );
  AOI21_X1 U20741 ( .B1(n18608), .B2(n17579), .A(n17578), .ZN(n17610) );
  OAI21_X1 U20742 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17680), .A(
        n17610), .ZN(n17594) );
  NOR2_X1 U20743 ( .A1(n17659), .A2(n17579), .ZN(n17596) );
  OAI211_X1 U20744 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17596), .B(n17580), .ZN(n17581) );
  NAND2_X1 U20745 ( .A1(n18122), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17943) );
  OAI211_X1 U20746 ( .C1(n17740), .C2(n17582), .A(n17581), .B(n17943), .ZN(
        n17588) );
  NOR2_X1 U20747 ( .A1(n17618), .A2(n17590), .ZN(n17947) );
  NAND2_X1 U20748 ( .A1(n17947), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17583) );
  XOR2_X1 U20749 ( .A(n17583), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17935) );
  OAI21_X1 U20750 ( .B1(n17777), .B2(n17585), .A(n17584), .ZN(n17586) );
  XOR2_X1 U20751 ( .A(n17586), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17940) );
  OAI22_X1 U20752 ( .A1(n17730), .A2(n17935), .B1(n17790), .B2(n17940), .ZN(
        n17587) );
  AOI211_X1 U20753 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17594), .A(
        n17588), .B(n17587), .ZN(n17589) );
  OAI21_X1 U20754 ( .B1(n17908), .B2(n17936), .A(n17589), .ZN(P3_U2805) );
  OR2_X1 U20755 ( .A1(n17590), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17958) );
  AOI22_X1 U20756 ( .A1(n18122), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17755), 
        .B2(n17591), .ZN(n17592) );
  INV_X1 U20757 ( .A(n17592), .ZN(n17593) );
  AOI221_X1 U20758 ( .B1(n17596), .B2(n17595), .C1(n17594), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17593), .ZN(n17601) );
  OAI22_X1 U20759 ( .A1(n17951), .A2(n17908), .B1(n17947), .B2(n17730), .ZN(
        n17612) );
  OAI21_X1 U20760 ( .B1(n17599), .B2(n17598), .A(n17597), .ZN(n17946) );
  AOI22_X1 U20761 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17612), .B1(
        n17815), .B2(n17946), .ZN(n17600) );
  OAI211_X1 U20762 ( .C1(n17705), .C2(n17958), .A(n17601), .B(n17600), .ZN(
        P3_U2806) );
  OAI22_X1 U20763 ( .A1(n17615), .A2(n17602), .B1(n17814), .B2(n17974), .ZN(
        n17603) );
  NOR2_X1 U20764 ( .A1(n17603), .A2(n17651), .ZN(n17604) );
  XOR2_X1 U20765 ( .A(n17604), .B(n17952), .Z(n17964) );
  INV_X1 U20766 ( .A(n17666), .ZN(n17643) );
  NOR2_X1 U20767 ( .A1(n17605), .A2(n17643), .ZN(n17613) );
  AOI21_X1 U20768 ( .B1(n18608), .B2(n17606), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17609) );
  OAI21_X1 U20769 ( .B1(n17755), .B2(n17568), .A(n17607), .ZN(n17608) );
  NAND2_X1 U20770 ( .A1(n18122), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17963) );
  OAI211_X1 U20771 ( .C1(n17610), .C2(n17609), .A(n17608), .B(n17963), .ZN(
        n17611) );
  AOI221_X1 U20772 ( .B1(n17613), .B2(n17952), .C1(n17612), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17611), .ZN(n17614) );
  OAI21_X1 U20773 ( .B1(n17790), .B2(n17964), .A(n17614), .ZN(P3_U2807) );
  INV_X1 U20774 ( .A(n17615), .ZN(n17616) );
  AOI221_X1 U20775 ( .B1(n17692), .B2(n17616), .C1(n17972), .C2(n17616), .A(
        n17651), .ZN(n17617) );
  XOR2_X1 U20776 ( .A(n17974), .B(n17617), .Z(n17981) );
  NOR2_X1 U20777 ( .A1(n17972), .A2(n17705), .ZN(n17628) );
  AOI22_X1 U20778 ( .A1(n17816), .A2(n17618), .B1(n17897), .B2(n18042), .ZN(
        n17704) );
  OAI21_X1 U20779 ( .B1(n17619), .B2(n17650), .A(n17704), .ZN(n17640) );
  OAI21_X1 U20780 ( .B1(n17620), .B2(n18737), .A(n17904), .ZN(n17621) );
  AOI21_X1 U20781 ( .B1(n17866), .B2(n17623), .A(n17621), .ZN(n17647) );
  OAI21_X1 U20782 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17680), .A(
        n17647), .ZN(n17633) );
  AOI22_X1 U20783 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17633), .B1(
        n17755), .B2(n17622), .ZN(n17626) );
  NOR2_X1 U20784 ( .A1(n17659), .A2(n17623), .ZN(n17635) );
  OAI211_X1 U20785 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17635), .B(n17624), .ZN(n17625) );
  OAI211_X1 U20786 ( .C1(n18797), .C2(n18221), .A(n17626), .B(n17625), .ZN(
        n17627) );
  AOI221_X1 U20787 ( .B1(n17628), .B2(n17974), .C1(n17640), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17627), .ZN(n17629) );
  OAI21_X1 U20788 ( .B1(n17790), .B2(n17981), .A(n17629), .ZN(P3_U2808) );
  OR2_X1 U20789 ( .A1(n17638), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17990) );
  AOI22_X1 U20790 ( .A1(n18122), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17755), 
        .B2(n17630), .ZN(n17631) );
  INV_X1 U20791 ( .A(n17631), .ZN(n17632) );
  AOI221_X1 U20792 ( .B1(n17635), .B2(n17634), .C1(n17633), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17632), .ZN(n17642) );
  NAND3_X1 U20793 ( .A1(n17814), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17636), .ZN(n17655) );
  OAI22_X1 U20794 ( .A1(n17638), .A2(n17655), .B1(n17637), .B2(n17675), .ZN(
        n17639) );
  XOR2_X1 U20795 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17639), .Z(
        n17983) );
  AOI22_X1 U20796 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17640), .B1(
        n17815), .B2(n17983), .ZN(n17641) );
  OAI211_X1 U20797 ( .C1(n17643), .C2(n17990), .A(n17642), .B(n17641), .ZN(
        P3_U2809) );
  INV_X1 U20798 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18004) );
  NOR2_X1 U20799 ( .A1(n17968), .A2(n18004), .ZN(n17991) );
  NAND2_X1 U20800 ( .A1(n17991), .A2(n17644), .ZN(n17999) );
  AOI21_X1 U20801 ( .B1(n18608), .B2(n17645), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17646) );
  OAI22_X1 U20802 ( .A1(n17647), .A2(n17646), .B1(n18221), .B2(n18794), .ZN(
        n17648) );
  AOI221_X1 U20803 ( .B1(n17755), .B2(n17649), .C1(n17568), .C2(n17649), .A(
        n17648), .ZN(n17654) );
  OAI21_X1 U20804 ( .B1(n17650), .B2(n17991), .A(n17704), .ZN(n17665) );
  AOI221_X1 U20805 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17655), 
        .C1(n18004), .C2(n17673), .A(n17651), .ZN(n17652) );
  XOR2_X1 U20806 ( .A(n17652), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n17995) );
  AOI22_X1 U20807 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17665), .B1(
        n17815), .B2(n17995), .ZN(n17653) );
  OAI211_X1 U20808 ( .C1(n17705), .C2(n17999), .A(n17654), .B(n17653), .ZN(
        P3_U2810) );
  OAI21_X1 U20809 ( .B1(n17675), .B2(n17673), .A(n17655), .ZN(n17656) );
  XOR2_X1 U20810 ( .A(n17656), .B(n18004), .Z(n18000) );
  AOI21_X1 U20811 ( .B1(n17866), .B2(n17658), .A(n17891), .ZN(n17689) );
  OAI21_X1 U20812 ( .B1(n17657), .B2(n18737), .A(n17689), .ZN(n17670) );
  AOI22_X1 U20813 ( .A1(n18122), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17670), .ZN(n17662) );
  NOR2_X1 U20814 ( .A1(n17659), .A2(n17658), .ZN(n17672) );
  OAI211_X1 U20815 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17672), .B(n17660), .ZN(n17661) );
  OAI211_X1 U20816 ( .C1(n17740), .C2(n17663), .A(n17662), .B(n17661), .ZN(
        n17664) );
  AOI221_X1 U20817 ( .B1(n17666), .B2(n18004), .C1(n17665), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17664), .ZN(n17667) );
  OAI21_X1 U20818 ( .B1(n18000), .B2(n17790), .A(n17667), .ZN(P3_U2811) );
  NAND2_X1 U20819 ( .A1(n18009), .A2(n17674), .ZN(n18016) );
  INV_X1 U20820 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17671) );
  OAI22_X1 U20821 ( .A1(n18221), .A2(n18789), .B1(n17740), .B2(n17668), .ZN(
        n17669) );
  AOI221_X1 U20822 ( .B1(n17672), .B2(n17671), .C1(n17670), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17669), .ZN(n17678) );
  OAI21_X1 U20823 ( .B1(n18009), .B2(n17705), .A(n17704), .ZN(n17686) );
  OAI21_X1 U20824 ( .B1(n17777), .B2(n17674), .A(n17673), .ZN(n17676) );
  XOR2_X1 U20825 ( .A(n17676), .B(n17675), .Z(n18012) );
  AOI22_X1 U20826 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17686), .B1(
        n17815), .B2(n18012), .ZN(n17677) );
  OAI211_X1 U20827 ( .C1(n17705), .C2(n18016), .A(n17678), .B(n17677), .ZN(
        P3_U2812) );
  AOI21_X1 U20828 ( .B1(n17679), .B2(n18608), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17690) );
  AOI22_X1 U20829 ( .A1(n18122), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n17681), 
        .B2(n17899), .ZN(n17688) );
  AOI21_X1 U20830 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17683), .A(
        n17682), .ZN(n18024) );
  NOR2_X1 U20831 ( .A1(n18033), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18021) );
  INV_X1 U20832 ( .A(n18021), .ZN(n17684) );
  OAI22_X1 U20833 ( .A1(n18024), .A2(n17790), .B1(n17705), .B2(n17684), .ZN(
        n17685) );
  AOI21_X1 U20834 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17686), .A(
        n17685), .ZN(n17687) );
  OAI211_X1 U20835 ( .C1(n17690), .C2(n17689), .A(n17688), .B(n17687), .ZN(
        P3_U2813) );
  NAND4_X1 U20836 ( .A1(n17691), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n17814), .A4(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17776) );
  INV_X1 U20837 ( .A(n17776), .ZN(n17791) );
  AOI22_X1 U20838 ( .A1(n17791), .A2(n17966), .B1(n17692), .B2(n17777), .ZN(
        n17693) );
  XOR2_X1 U20839 ( .A(n18033), .B(n17693), .Z(n18030) );
  AOI21_X1 U20840 ( .B1(n17866), .B2(n17694), .A(n17891), .ZN(n17720) );
  OAI21_X1 U20841 ( .B1(n17695), .B2(n18737), .A(n17720), .ZN(n17711) );
  AOI22_X1 U20842 ( .A1(n18122), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17711), .ZN(n17700) );
  NAND2_X1 U20843 ( .A1(n17719), .A2(n17696), .ZN(n17758) );
  NOR2_X1 U20844 ( .A1(n17697), .A2(n17758), .ZN(n17713) );
  OAI211_X1 U20845 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17713), .B(n17698), .ZN(n17699) );
  OAI211_X1 U20846 ( .C1(n17701), .C2(n17740), .A(n17700), .B(n17699), .ZN(
        n17702) );
  AOI21_X1 U20847 ( .B1(n17815), .B2(n18030), .A(n17702), .ZN(n17703) );
  OAI221_X1 U20848 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17705), 
        .C1(n18033), .C2(n17704), .A(n17703), .ZN(P3_U2814) );
  NAND2_X1 U20849 ( .A1(n18052), .A2(n17791), .ZN(n17749) );
  NAND2_X1 U20850 ( .A1(n17777), .A2(n17706), .ZN(n17774) );
  NOR2_X1 U20851 ( .A1(n17785), .A2(n17774), .ZN(n17764) );
  INV_X1 U20852 ( .A(n17764), .ZN(n17750) );
  NOR2_X1 U20853 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17750), .ZN(
        n17753) );
  INV_X1 U20854 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17747) );
  NAND2_X1 U20855 ( .A1(n17753), .A2(n17747), .ZN(n17726) );
  NOR2_X1 U20856 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18080), .ZN(
        n18076) );
  AOI221_X1 U20857 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17749), 
        .C1(n18054), .C2(n17726), .A(n18076), .ZN(n17707) );
  XOR2_X1 U20858 ( .A(n18037), .B(n17707), .Z(n18049) );
  NOR2_X1 U20859 ( .A1(n18221), .A2(n18783), .ZN(n18047) );
  NOR3_X1 U20860 ( .A1(n18090), .A2(n18054), .A3(n18055), .ZN(n17724) );
  NOR2_X1 U20861 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17724), .ZN(
        n18043) );
  NAND2_X1 U20862 ( .A1(n17897), .A2(n18042), .ZN(n17709) );
  OAI22_X1 U20863 ( .A1(n18043), .A2(n17709), .B1(n17740), .B2(n17708), .ZN(
        n17710) );
  AOI211_X1 U20864 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17711), .A(
        n18047), .B(n17710), .ZN(n17716) );
  NOR2_X1 U20865 ( .A1(n18036), .A2(n17730), .ZN(n17714) );
  NAND2_X1 U20866 ( .A1(n17717), .A2(n18037), .ZN(n18040) );
  AOI22_X1 U20867 ( .A1(n17714), .A2(n18040), .B1(n17713), .B2(n17712), .ZN(
        n17715) );
  OAI211_X1 U20868 ( .C1(n17790), .C2(n18049), .A(n17716), .B(n17715), .ZN(
        P3_U2815) );
  OAI21_X1 U20869 ( .B1(n17718), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17717), .ZN(n18050) );
  NAND2_X1 U20870 ( .A1(n18608), .A2(n17719), .ZN(n17769) );
  AOI221_X1 U20871 ( .B1(n17737), .B2(n17721), .C1(n17769), .C2(n17721), .A(
        n17720), .ZN(n17722) );
  NOR2_X1 U20872 ( .A1(n18221), .A2(n18782), .ZN(n18061) );
  AOI211_X1 U20873 ( .C1(n17723), .C2(n17899), .A(n17722), .B(n18061), .ZN(
        n17729) );
  OR2_X1 U20874 ( .A1(n18055), .A2(n18090), .ZN(n17725) );
  AOI21_X1 U20875 ( .B1(n18054), .B2(n17725), .A(n17724), .ZN(n18063) );
  AOI21_X1 U20876 ( .B1(n17726), .B2(n17749), .A(n18076), .ZN(n17727) );
  XOR2_X1 U20877 ( .A(n17727), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18062) );
  AOI22_X1 U20878 ( .A1(n17897), .A2(n18063), .B1(n17815), .B2(n18062), .ZN(
        n17728) );
  OAI211_X1 U20879 ( .C1(n17730), .C2(n18050), .A(n17729), .B(n17728), .ZN(
        P3_U2816) );
  NAND2_X1 U20880 ( .A1(n17731), .A2(n18052), .ZN(n18068) );
  NAND2_X1 U20881 ( .A1(n17732), .A2(n18052), .ZN(n18067) );
  AOI22_X1 U20882 ( .A1(n17816), .A2(n18068), .B1(n17897), .B2(n18067), .ZN(
        n17761) );
  AOI21_X1 U20883 ( .B1(n17866), .B2(n17733), .A(n17891), .ZN(n17827) );
  NAND2_X1 U20884 ( .A1(n17866), .A2(n17734), .ZN(n17735) );
  OAI211_X1 U20885 ( .C1(n17736), .C2(n18737), .A(n17827), .B(n17735), .ZN(
        n17756) );
  NOR2_X1 U20886 ( .A1(n18221), .A2(n18779), .ZN(n17742) );
  OAI21_X1 U20887 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17737), .ZN(n17738) );
  OAI22_X1 U20888 ( .A1(n17740), .A2(n17739), .B1(n17758), .B2(n17738), .ZN(
        n17741) );
  AOI211_X1 U20889 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17756), .A(
        n17742), .B(n17741), .ZN(n17746) );
  INV_X1 U20890 ( .A(n17743), .ZN(n17751) );
  OAI21_X1 U20891 ( .B1(n17751), .B2(n17750), .A(n17749), .ZN(n17744) );
  XOR2_X1 U20892 ( .A(n17744), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18077) );
  NOR2_X1 U20893 ( .A1(n17802), .A2(n18096), .ZN(n17748) );
  AOI22_X1 U20894 ( .A1(n17815), .A2(n18077), .B1(n18076), .B2(n17748), .ZN(
        n17745) );
  OAI211_X1 U20895 ( .C1(n17761), .C2(n17747), .A(n17746), .B(n17745), .ZN(
        P3_U2817) );
  INV_X1 U20896 ( .A(n17748), .ZN(n17762) );
  NOR2_X1 U20897 ( .A1(n17766), .A2(n17776), .ZN(n17775) );
  OAI211_X1 U20898 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17775), .A(
        n17749), .B(n17751), .ZN(n17752) );
  OAI22_X1 U20899 ( .A1(n17753), .A2(n17752), .B1(n17751), .B2(n17750), .ZN(
        n18084) );
  AOI22_X1 U20900 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17756), .B1(
        n17755), .B2(n17754), .ZN(n17757) );
  NAND2_X1 U20901 ( .A1(n18122), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18085) );
  OAI211_X1 U20902 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17758), .A(
        n17757), .B(n18085), .ZN(n17759) );
  AOI21_X1 U20903 ( .B1(n17815), .B2(n18084), .A(n17759), .ZN(n17760) );
  OAI221_X1 U20904 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17762), 
        .C1(n18080), .C2(n17761), .A(n17760), .ZN(P3_U2818) );
  AOI22_X1 U20905 ( .A1(n18122), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17763), 
        .B2(n17899), .ZN(n17773) );
  NOR2_X1 U20906 ( .A1(n17775), .A2(n17764), .ZN(n17765) );
  XNOR2_X1 U20907 ( .A(n17765), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18100) );
  NOR2_X1 U20908 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17766), .ZN(
        n18099) );
  AOI22_X1 U20909 ( .A1(n17815), .A2(n18100), .B1(n18099), .B2(n17767), .ZN(
        n17772) );
  NOR2_X1 U20910 ( .A1(n18094), .A2(n17802), .ZN(n17786) );
  AOI22_X1 U20911 ( .A1(n18089), .A2(n17816), .B1(n17897), .B2(n18090), .ZN(
        n17801) );
  INV_X1 U20912 ( .A(n17801), .ZN(n17787) );
  OAI21_X1 U20913 ( .B1(n17786), .B2(n17787), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17771) );
  NAND2_X1 U20914 ( .A1(n18608), .A2(n17768), .ZN(n17855) );
  NOR2_X1 U20915 ( .A1(n10034), .A2(n17855), .ZN(n17805) );
  NAND3_X1 U20916 ( .A1(n17807), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17805), .ZN(n17794) );
  NOR2_X1 U20917 ( .A1(n17782), .A2(n17794), .ZN(n17781) );
  INV_X1 U20918 ( .A(n17848), .ZN(n17900) );
  OAI211_X1 U20919 ( .C1(n17781), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17900), .B(n17769), .ZN(n17770) );
  NAND4_X1 U20920 ( .A1(n17773), .A2(n17772), .A3(n17771), .A4(n17770), .ZN(
        P3_U2819) );
  INV_X1 U20921 ( .A(n17774), .ZN(n17792) );
  NOR2_X1 U20922 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18125), .ZN(
        n18110) );
  AOI21_X1 U20923 ( .B1(n18110), .B2(n17776), .A(n17775), .ZN(n17780) );
  NAND4_X1 U20924 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17778), .A3(
        n17777), .A4(n18125), .ZN(n17779) );
  OAI211_X1 U20925 ( .C1(n17792), .C2(n17785), .A(n17780), .B(n17779), .ZN(
        n18112) );
  AOI211_X1 U20926 ( .C1(n17794), .C2(n17782), .A(n17848), .B(n17781), .ZN(
        n17783) );
  INV_X1 U20927 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18773) );
  NOR2_X1 U20928 ( .A1(n18221), .A2(n18773), .ZN(n18108) );
  AOI211_X1 U20929 ( .C1(n17784), .C2(n17899), .A(n17783), .B(n18108), .ZN(
        n17789) );
  AOI22_X1 U20930 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17787), .B1(
        n17786), .B2(n17785), .ZN(n17788) );
  OAI211_X1 U20931 ( .C1(n17790), .C2(n18112), .A(n17789), .B(n17788), .ZN(
        P3_U2820) );
  NOR2_X1 U20932 ( .A1(n17792), .A2(n17791), .ZN(n17793) );
  XOR2_X1 U20933 ( .A(n17793), .B(n18125), .Z(n18121) );
  NOR2_X1 U20934 ( .A1(n18221), .A2(n18771), .ZN(n17799) );
  INV_X1 U20935 ( .A(n17794), .ZN(n17796) );
  AOI22_X1 U20936 ( .A1(n17807), .A2(n17805), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17900), .ZN(n17795) );
  OAI22_X1 U20937 ( .A1(n17889), .A2(n17797), .B1(n17796), .B2(n17795), .ZN(
        n17798) );
  AOI211_X1 U20938 ( .C1(n17815), .C2(n18121), .A(n17799), .B(n17798), .ZN(
        n17800) );
  OAI221_X1 U20939 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17802), .C1(
        n18125), .C2(n17801), .A(n17800), .ZN(P3_U2821) );
  AOI21_X1 U20940 ( .B1(n17804), .B2(n18132), .A(n17803), .ZN(n18140) );
  AOI22_X1 U20941 ( .A1(n17897), .A2(n18140), .B1(n18144), .B2(
        P3_REIP_REG_8__SCAN_IN), .ZN(n17819) );
  INV_X1 U20942 ( .A(n17805), .ZN(n17843) );
  OAI21_X1 U20943 ( .B1(n17828), .B2(n17843), .A(n17806), .ZN(n17809) );
  OAI21_X1 U20944 ( .B1(n17807), .B2(n18347), .A(n17827), .ZN(n17808) );
  AOI22_X1 U20945 ( .A1(n17810), .A2(n17899), .B1(n17809), .B2(n17808), .ZN(
        n17818) );
  INV_X1 U20946 ( .A(n17811), .ZN(n17812) );
  AOI21_X1 U20947 ( .B1(n17814), .B2(n17813), .A(n17812), .ZN(n18138) );
  AOI22_X1 U20948 ( .A1(n17816), .A2(n18136), .B1(n17815), .B2(n18138), .ZN(
        n17817) );
  NAND3_X1 U20949 ( .A1(n17819), .A2(n17818), .A3(n17817), .ZN(P3_U2822) );
  OAI21_X1 U20950 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17820), .A(
        n17821), .ZN(n18152) );
  OAI21_X1 U20951 ( .B1(n17824), .B2(n17823), .A(n17822), .ZN(n17825) );
  XOR2_X1 U20952 ( .A(n17825), .B(n18147), .Z(n18148) );
  AOI22_X1 U20953 ( .A1(n17897), .A2(n18148), .B1(n18144), .B2(
        P3_REIP_REG_7__SCAN_IN), .ZN(n17826) );
  OAI221_X1 U20954 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17843), .C1(
        n17828), .C2(n17827), .A(n17826), .ZN(n17829) );
  AOI21_X1 U20955 ( .B1(n17830), .B2(n17899), .A(n17829), .ZN(n17831) );
  OAI21_X1 U20956 ( .B1(n17907), .B2(n18152), .A(n17831), .ZN(P3_U2823) );
  OAI21_X1 U20957 ( .B1(n17834), .B2(n17833), .A(n17832), .ZN(n18157) );
  OAI21_X1 U20958 ( .B1(n17848), .B2(n10034), .A(n17855), .ZN(n17842) );
  AOI22_X1 U20959 ( .A1(n17837), .A2(n17845), .B1(n17836), .B2(n17835), .ZN(
        n17838) );
  XOR2_X1 U20960 ( .A(n17839), .B(n17838), .Z(n18163) );
  OAI22_X1 U20961 ( .A1(n17889), .A2(n17840), .B1(n18163), .B2(n17908), .ZN(
        n17841) );
  AOI21_X1 U20962 ( .B1(n17843), .B2(n17842), .A(n17841), .ZN(n17844) );
  NAND2_X1 U20963 ( .A1(n18122), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18161) );
  OAI211_X1 U20964 ( .C1(n17907), .C2(n18157), .A(n17844), .B(n18161), .ZN(
        P3_U2824) );
  OAI21_X1 U20965 ( .B1(n17847), .B2(n17846), .A(n17845), .ZN(n18164) );
  AOI221_X1 U20966 ( .B1(n17891), .B2(n17850), .C1(n17849), .C2(n17850), .A(
        n17848), .ZN(n17856) );
  OAI21_X1 U20967 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17852), .A(
        n17851), .ZN(n18171) );
  OAI22_X1 U20968 ( .A1(n17889), .A2(n17853), .B1(n17907), .B2(n18171), .ZN(
        n17854) );
  AOI21_X1 U20969 ( .B1(n17856), .B2(n17855), .A(n17854), .ZN(n17857) );
  NAND2_X1 U20970 ( .A1(n18144), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18169) );
  OAI211_X1 U20971 ( .C1(n17908), .C2(n18164), .A(n17857), .B(n18169), .ZN(
        P3_U2825) );
  OAI21_X1 U20972 ( .B1(n17860), .B2(n17859), .A(n17858), .ZN(n18172) );
  OAI21_X1 U20973 ( .B1(n17863), .B2(n17862), .A(n17861), .ZN(n18178) );
  OAI22_X1 U20974 ( .A1(n17907), .A2(n18178), .B1(n18347), .B2(n17864), .ZN(
        n17865) );
  AOI21_X1 U20975 ( .B1(n18122), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17865), .ZN(
        n17871) );
  INV_X1 U20976 ( .A(n17866), .ZN(n17867) );
  OAI21_X1 U20977 ( .B1(n17868), .B2(n17867), .A(n17904), .ZN(n17880) );
  AOI22_X1 U20978 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17880), .B1(
        n17869), .B2(n17899), .ZN(n17870) );
  OAI211_X1 U20979 ( .C1(n17908), .C2(n18172), .A(n17871), .B(n17870), .ZN(
        P3_U2826) );
  OAI21_X1 U20980 ( .B1(n17874), .B2(n17873), .A(n17872), .ZN(n18180) );
  NOR2_X1 U20981 ( .A1(n17891), .A2(n17892), .ZN(n17879) );
  OAI21_X1 U20982 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17876), .A(
        n17875), .ZN(n18187) );
  OAI22_X1 U20983 ( .A1(n17889), .A2(n17877), .B1(n17907), .B2(n18187), .ZN(
        n17878) );
  AOI221_X1 U20984 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17880), .C1(
        n17879), .C2(n17880), .A(n17878), .ZN(n17881) );
  NAND2_X1 U20985 ( .A1(n18144), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18185) );
  OAI211_X1 U20986 ( .C1(n17908), .C2(n18180), .A(n17881), .B(n18185), .ZN(
        P3_U2827) );
  OAI21_X1 U20987 ( .B1(n17884), .B2(n17883), .A(n17882), .ZN(n18199) );
  OAI21_X1 U20988 ( .B1(n17887), .B2(n17886), .A(n17885), .ZN(n18204) );
  OAI22_X1 U20989 ( .A1(n17889), .A2(n17888), .B1(n17907), .B2(n18204), .ZN(
        n17890) );
  AOI221_X1 U20990 ( .B1(n18608), .B2(n17892), .C1(n17891), .C2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17890), .ZN(n17893) );
  NAND2_X1 U20991 ( .A1(n18144), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18202) );
  OAI211_X1 U20992 ( .C1(n17908), .C2(n18199), .A(n17893), .B(n18202), .ZN(
        P3_U2828) );
  OAI21_X1 U20993 ( .B1(n17903), .B2(n17895), .A(n17894), .ZN(n18215) );
  NAND2_X1 U20994 ( .A1(n18859), .A2(n10256), .ZN(n17896) );
  XNOR2_X1 U20995 ( .A(n17896), .B(n17895), .ZN(n18211) );
  AOI22_X1 U20996 ( .A1(n17897), .A2(n18211), .B1(n18144), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17902) );
  AOI22_X1 U20997 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17900), .B1(
        n17899), .B2(n17898), .ZN(n17901) );
  OAI211_X1 U20998 ( .C1(n17907), .C2(n18215), .A(n17902), .B(n17901), .ZN(
        P3_U2829) );
  AOI21_X1 U20999 ( .B1(n10256), .B2(n18859), .A(n17903), .ZN(n18219) );
  INV_X1 U21000 ( .A(n18219), .ZN(n18217) );
  NAND3_X1 U21001 ( .A1(n18842), .A2(n18737), .A3(n17904), .ZN(n17905) );
  AOI22_X1 U21002 ( .A1(n18122), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17905), .ZN(n17906) );
  OAI221_X1 U21003 ( .B1(n18219), .B2(n17908), .C1(n18217), .C2(n17907), .A(
        n17906), .ZN(P3_U2830) );
  NOR2_X1 U21004 ( .A1(n17909), .A2(n17965), .ZN(n17918) );
  NOR2_X1 U21005 ( .A1(n17953), .A2(n17924), .ZN(n17912) );
  NAND2_X1 U21006 ( .A1(n18691), .A2(n18859), .ZN(n18188) );
  INV_X1 U21007 ( .A(n18188), .ZN(n17911) );
  NOR2_X1 U21008 ( .A1(n18691), .A2(n18682), .ZN(n18189) );
  INV_X1 U21009 ( .A(n18189), .ZN(n18130) );
  OAI21_X1 U21010 ( .B1(n17911), .B2(n17910), .A(n18130), .ZN(n17949) );
  AOI21_X1 U21011 ( .B1(n17912), .B2(n17949), .A(n18133), .ZN(n17939) );
  INV_X1 U21012 ( .A(n18137), .ZN(n18035) );
  OAI22_X1 U21013 ( .A1(n17914), .A2(n18035), .B1(n17913), .B2(n18198), .ZN(
        n17915) );
  AOI211_X1 U21014 ( .C1(n18131), .C2(n17916), .A(n17939), .B(n17915), .ZN(
        n17925) );
  INV_X1 U21015 ( .A(n17925), .ZN(n17917) );
  MUX2_X1 U21016 ( .A(n17918), .B(n17917), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17920) );
  AOI22_X1 U21017 ( .A1(n18206), .A2(n17920), .B1(n18139), .B2(n17919), .ZN(
        n17922) );
  NAND2_X1 U21018 ( .A1(n18144), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17921) );
  OAI211_X1 U21019 ( .C1(n18207), .C2(n17923), .A(n17922), .B(n17921), .ZN(
        P3_U2835) );
  INV_X1 U21020 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17927) );
  OR4_X1 U21021 ( .A1(n17959), .A2(n17924), .A3(n17941), .A4(n17965), .ZN(
        n17926) );
  AOI211_X1 U21022 ( .C1(n17927), .C2(n17926), .A(n17925), .B(n18222), .ZN(
        n17928) );
  AOI21_X1 U21023 ( .B1(n18201), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17928), .ZN(n17930) );
  OAI211_X1 U21024 ( .C1(n17931), .C2(n18113), .A(n17930), .B(n17929), .ZN(
        P3_U2836) );
  INV_X1 U21025 ( .A(n18179), .ZN(n18154) );
  INV_X1 U21026 ( .A(n18091), .ZN(n17932) );
  NOR4_X1 U21027 ( .A1(n18154), .A2(n17934), .A3(n17933), .A4(n17932), .ZN(
        n17938) );
  OAI22_X1 U21028 ( .A1(n18198), .A2(n17936), .B1(n18035), .B2(n17935), .ZN(
        n17937) );
  AOI221_X1 U21029 ( .B1(n17939), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17938), .C2(n17941), .A(n17937), .ZN(n17945) );
  OAI22_X1 U21030 ( .A1(n17941), .A2(n18207), .B1(n18113), .B2(n17940), .ZN(
        n17942) );
  INV_X1 U21031 ( .A(n17942), .ZN(n17944) );
  OAI211_X1 U21032 ( .C1(n17945), .C2(n18222), .A(n17944), .B(n17943), .ZN(
        P3_U2837) );
  AOI22_X1 U21033 ( .A1(n18122), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18139), 
        .B2(n17946), .ZN(n17957) );
  INV_X1 U21034 ( .A(n17947), .ZN(n17948) );
  AOI21_X1 U21035 ( .B1(n18137), .B2(n17948), .A(n18201), .ZN(n17950) );
  OAI211_X1 U21036 ( .C1(n17951), .C2(n18198), .A(n17950), .B(n17949), .ZN(
        n17955) );
  NOR3_X1 U21037 ( .A1(n17953), .A2(n17952), .A3(n17955), .ZN(n17954) );
  NOR2_X1 U21038 ( .A1(n18144), .A2(n17954), .ZN(n17960) );
  OAI211_X1 U21039 ( .C1(n18131), .C2(n17955), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17960), .ZN(n17956) );
  OAI211_X1 U21040 ( .C1(n17958), .C2(n18034), .A(n17957), .B(n17956), .ZN(
        P3_U2838) );
  NOR2_X1 U21041 ( .A1(n17959), .A2(n17965), .ZN(n17961) );
  OAI221_X1 U21042 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17961), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18207), .A(n17960), .ZN(
        n17962) );
  OAI211_X1 U21043 ( .C1(n17964), .C2(n18113), .A(n17963), .B(n17962), .ZN(
        P3_U2839) );
  AOI221_X1 U21044 ( .B1(n17972), .B2(n17974), .C1(n17965), .C2(n17974), .A(
        n18222), .ZN(n17978) );
  NOR2_X1 U21045 ( .A1(n18665), .A2(n18137), .ZN(n18093) );
  INV_X1 U21046 ( .A(n18093), .ZN(n17971) );
  NOR2_X1 U21047 ( .A1(n18673), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17970) );
  NOR3_X1 U21048 ( .A1(n18193), .A2(n18843), .A3(n18859), .ZN(n18194) );
  NAND3_X1 U21049 ( .A1(n17966), .A2(n18091), .A3(n18194), .ZN(n18026) );
  AOI21_X1 U21050 ( .B1(n18006), .B2(n17991), .A(n18673), .ZN(n17967) );
  AOI221_X1 U21051 ( .B1(n17968), .B2(n18691), .C1(n18026), .C2(n18691), .A(
        n17967), .ZN(n17969) );
  OAI221_X1 U21052 ( .B1(n18701), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), 
        .C1(n18701), .C2(n18008), .A(n17969), .ZN(n17993) );
  AOI211_X1 U21053 ( .C1(n17972), .C2(n17971), .A(n17970), .B(n17993), .ZN(
        n17985) );
  INV_X1 U21054 ( .A(n18057), .ZN(n18205) );
  INV_X1 U21055 ( .A(n18042), .ZN(n17973) );
  OAI22_X1 U21056 ( .A1(n18036), .A2(n18035), .B1(n17973), .B2(n18198), .ZN(
        n17984) );
  AOI211_X1 U21057 ( .C1(n18205), .C2(n17975), .A(n17974), .B(n17984), .ZN(
        n17976) );
  OAI211_X1 U21058 ( .C1(n18673), .C2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n17985), .B(n17976), .ZN(n17977) );
  AOI22_X1 U21059 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18201), .B1(
        n17978), .B2(n17977), .ZN(n17980) );
  NAND2_X1 U21060 ( .A1(n18122), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17979) );
  OAI211_X1 U21061 ( .C1(n17981), .C2(n18113), .A(n17980), .B(n17979), .ZN(
        P3_U2840) );
  NAND2_X1 U21062 ( .A1(n17982), .A2(n18020), .ZN(n18005) );
  AOI22_X1 U21063 ( .A1(n18122), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18139), 
        .B2(n17983), .ZN(n17989) );
  NOR2_X1 U21064 ( .A1(n18222), .A2(n17984), .ZN(n18007) );
  OAI211_X1 U21065 ( .C1(n18057), .C2(n17986), .A(n18007), .B(n17985), .ZN(
        n17987) );
  NAND3_X1 U21066 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18221), .A3(
        n17987), .ZN(n17988) );
  OAI211_X1 U21067 ( .C1(n18005), .C2(n17990), .A(n17989), .B(n17988), .ZN(
        P3_U2841) );
  NAND2_X1 U21068 ( .A1(n18205), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17994) );
  OAI21_X1 U21069 ( .B1(n17991), .B2(n18093), .A(n18007), .ZN(n17992) );
  OAI21_X1 U21070 ( .B1(n17993), .B2(n17992), .A(n18221), .ZN(n18003) );
  OAI21_X1 U21071 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17994), .A(
        n18003), .ZN(n17996) );
  AOI22_X1 U21072 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17996), .B1(
        n18139), .B2(n17995), .ZN(n17998) );
  NAND2_X1 U21073 ( .A1(n18122), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17997) );
  OAI211_X1 U21074 ( .C1(n17999), .C2(n18034), .A(n17998), .B(n17997), .ZN(
        P3_U2842) );
  OAI22_X1 U21075 ( .A1(n18221), .A2(n18791), .B1(n18113), .B2(n18000), .ZN(
        n18001) );
  INV_X1 U21076 ( .A(n18001), .ZN(n18002) );
  OAI221_X1 U21077 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18005), 
        .C1(n18004), .C2(n18003), .A(n18002), .ZN(P3_U2843) );
  NAND3_X1 U21078 ( .A1(n18006), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18188), .ZN(n18011) );
  INV_X1 U21079 ( .A(n18007), .ZN(n18029) );
  OAI22_X1 U21080 ( .A1(n18009), .A2(n18093), .B1(n18008), .B2(n18701), .ZN(
        n18010) );
  AOI211_X1 U21081 ( .C1(n18130), .C2(n18011), .A(n18029), .B(n18010), .ZN(
        n18018) );
  AOI221_X1 U21082 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18018), 
        .C1(n18189), .C2(n18018), .A(n18122), .ZN(n18013) );
  AOI22_X1 U21083 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18013), .B1(
        n18139), .B2(n18012), .ZN(n18015) );
  NAND2_X1 U21084 ( .A1(n18122), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18014) );
  OAI211_X1 U21085 ( .C1(n18016), .C2(n18034), .A(n18015), .B(n18014), .ZN(
        P3_U2844) );
  NOR3_X1 U21086 ( .A1(n18122), .A2(n18018), .A3(n18017), .ZN(n18019) );
  AOI21_X1 U21087 ( .B1(n18021), .B2(n18020), .A(n18019), .ZN(n18023) );
  NAND2_X1 U21088 ( .A1(n18122), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18022) );
  OAI211_X1 U21089 ( .C1(n18024), .C2(n18113), .A(n18023), .B(n18022), .ZN(
        P3_U2845) );
  AND2_X1 U21090 ( .A1(n18682), .A2(n18025), .ZN(n18116) );
  AOI21_X1 U21091 ( .B1(n18667), .B2(n18114), .A(n18116), .ZN(n18070) );
  OAI21_X1 U21092 ( .B1(n18037), .B2(n18691), .A(n18026), .ZN(n18027) );
  OAI211_X1 U21093 ( .C1(n18073), .C2(n18028), .A(n18070), .B(n18027), .ZN(
        n18039) );
  OAI221_X1 U21094 ( .B1(n18029), .B2(n18131), .C1(n18029), .C2(n18039), .A(
        n18221), .ZN(n18032) );
  AOI22_X1 U21095 ( .A1(n18122), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18139), 
        .B2(n18030), .ZN(n18031) );
  OAI221_X1 U21096 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18034), 
        .C1(n18033), .C2(n18032), .A(n18031), .ZN(P3_U2846) );
  NOR2_X1 U21097 ( .A1(n18036), .A2(n18035), .ZN(n18041) );
  NAND2_X1 U21098 ( .A1(n18037), .A2(n18051), .ZN(n18038) );
  AOI22_X1 U21099 ( .A1(n18041), .A2(n18040), .B1(n18039), .B2(n18038), .ZN(
        n18045) );
  NAND2_X1 U21100 ( .A1(n18665), .A2(n18042), .ZN(n18044) );
  AOI211_X1 U21101 ( .C1(n18045), .C2(n18044), .A(n18043), .B(n18222), .ZN(
        n18046) );
  AOI211_X1 U21102 ( .C1(n18201), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18047), .B(n18046), .ZN(n18048) );
  OAI21_X1 U21103 ( .B1(n18113), .B2(n18049), .A(n18048), .ZN(P3_U2847) );
  INV_X1 U21104 ( .A(n18050), .ZN(n18060) );
  OAI21_X1 U21105 ( .B1(n18055), .B2(n18051), .A(n18054), .ZN(n18059) );
  NAND3_X1 U21106 ( .A1(n18052), .A2(n18091), .A3(n18194), .ZN(n18082) );
  NAND2_X1 U21107 ( .A1(n18691), .A2(n18082), .ZN(n18072) );
  OAI211_X1 U21108 ( .C1(n18052), .C2(n18701), .A(n18070), .B(n18072), .ZN(
        n18053) );
  AOI211_X1 U21109 ( .C1(n18682), .C2(n18055), .A(n18054), .B(n18053), .ZN(
        n18056) );
  OAI21_X1 U21110 ( .B1(n18057), .B2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n18056), .ZN(n18058) );
  AOI22_X1 U21111 ( .A1(n18137), .A2(n18060), .B1(n18059), .B2(n18058), .ZN(
        n18066) );
  AOI21_X1 U21112 ( .B1(n18201), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18061), .ZN(n18065) );
  AOI22_X1 U21113 ( .A1(n18218), .A2(n18063), .B1(n18139), .B2(n18062), .ZN(
        n18064) );
  OAI211_X1 U21114 ( .C1(n18066), .C2(n18222), .A(n18065), .B(n18064), .ZN(
        P3_U2848) );
  INV_X1 U21115 ( .A(n18067), .ZN(n18071) );
  AOI22_X1 U21116 ( .A1(n18137), .A2(n18068), .B1(n18096), .B2(n18103), .ZN(
        n18069) );
  OAI211_X1 U21117 ( .C1(n18071), .C2(n18198), .A(n18070), .B(n18069), .ZN(
        n18081) );
  OAI211_X1 U21118 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18073), .A(
        n18206), .B(n18072), .ZN(n18074) );
  OAI21_X1 U21119 ( .B1(n18081), .B2(n18074), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18079) );
  NAND2_X1 U21120 ( .A1(n18206), .A2(n18075), .ZN(n18126) );
  NOR2_X1 U21121 ( .A1(n18096), .A2(n18126), .ZN(n18083) );
  AOI22_X1 U21122 ( .A1(n18139), .A2(n18077), .B1(n18076), .B2(n18083), .ZN(
        n18078) );
  OAI221_X1 U21123 ( .B1(n18122), .B2(n18079), .C1(n18221), .C2(n18779), .A(
        n18078), .ZN(P3_U2849) );
  AOI211_X1 U21124 ( .C1(n18082), .C2(n18691), .A(n18081), .B(n18080), .ZN(
        n18088) );
  AOI21_X1 U21125 ( .B1(n18206), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18083), .ZN(n18087) );
  AOI22_X1 U21126 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18201), .B1(
        n18139), .B2(n18084), .ZN(n18086) );
  OAI211_X1 U21127 ( .C1(n18088), .C2(n18087), .A(n18086), .B(n18085), .ZN(
        P3_U2850) );
  AOI22_X1 U21128 ( .A1(n18665), .A2(n18090), .B1(n18137), .B2(n18089), .ZN(
        n18119) );
  NAND2_X1 U21129 ( .A1(n18091), .A2(n18194), .ZN(n18115) );
  OAI21_X1 U21130 ( .B1(n18125), .B2(n18115), .A(n18691), .ZN(n18092) );
  OAI211_X1 U21131 ( .C1(n18094), .C2(n18093), .A(n18119), .B(n18092), .ZN(
        n18095) );
  AOI211_X1 U21132 ( .C1(n18667), .C2(n18114), .A(n18201), .B(n18095), .ZN(
        n18106) );
  NAND2_X1 U21133 ( .A1(n18096), .A2(n18103), .ZN(n18097) );
  OAI211_X1 U21134 ( .C1(n18679), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18106), .B(n18097), .ZN(n18098) );
  OAI21_X1 U21135 ( .B1(n18116), .B2(n18098), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18102) );
  INV_X1 U21136 ( .A(n18126), .ZN(n18109) );
  AOI22_X1 U21137 ( .A1(n18139), .A2(n18100), .B1(n18109), .B2(n18099), .ZN(
        n18101) );
  OAI221_X1 U21138 ( .B1(n18122), .B2(n18102), .C1(n18221), .C2(n18775), .A(
        n18101), .ZN(P3_U2851) );
  OAI21_X1 U21139 ( .B1(n18116), .B2(n18125), .A(n18103), .ZN(n18105) );
  AOI211_X1 U21140 ( .C1(n18106), .C2(n18105), .A(n18122), .B(n18104), .ZN(
        n18107) );
  AOI211_X1 U21141 ( .C1(n18110), .C2(n18109), .A(n18108), .B(n18107), .ZN(
        n18111) );
  OAI21_X1 U21142 ( .B1(n18113), .B2(n18112), .A(n18111), .ZN(P3_U2852) );
  NAND2_X1 U21143 ( .A1(n18667), .A2(n18114), .ZN(n18118) );
  OAI21_X1 U21144 ( .B1(n18116), .B2(n18691), .A(n18115), .ZN(n18117) );
  NAND4_X1 U21145 ( .A1(n18206), .A2(n18119), .A3(n18118), .A4(n18117), .ZN(
        n18120) );
  NAND2_X1 U21146 ( .A1(n18221), .A2(n18120), .ZN(n18124) );
  AOI22_X1 U21147 ( .A1(n18122), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18139), 
        .B2(n18121), .ZN(n18123) );
  OAI221_X1 U21148 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18126), .C1(
        n18125), .C2(n18124), .A(n18123), .ZN(P3_U2853) );
  OAI211_X1 U21149 ( .C1(n18701), .C2(n18127), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18188), .ZN(n18128) );
  AOI21_X1 U21150 ( .B1(n18130), .B2(n18129), .A(n18128), .ZN(n18183) );
  NAND3_X1 U21151 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n18183), .ZN(n18155) );
  AOI221_X1 U21152 ( .B1(n18158), .B2(n18131), .C1(n18155), .C2(n18131), .A(
        n18147), .ZN(n18145) );
  NOR3_X1 U21153 ( .A1(n18133), .A2(n18145), .A3(n18132), .ZN(n18135) );
  NOR4_X1 U21154 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18154), .A3(
        n18147), .A4(n18146), .ZN(n18134) );
  AOI211_X1 U21155 ( .C1(n18137), .C2(n18136), .A(n18135), .B(n18134), .ZN(
        n18143) );
  AOI22_X1 U21156 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18201), .B1(
        n18144), .B2(P3_REIP_REG_8__SCAN_IN), .ZN(n18142) );
  AOI22_X1 U21157 ( .A1(n18218), .A2(n18140), .B1(n18139), .B2(n18138), .ZN(
        n18141) );
  OAI211_X1 U21158 ( .C1(n18143), .C2(n18222), .A(n18142), .B(n18141), .ZN(
        P3_U2854) );
  AOI22_X1 U21159 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18201), .B1(
        n18144), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n18151) );
  AOI221_X1 U21160 ( .B1(n18154), .B2(n18147), .C1(n18146), .C2(n18147), .A(
        n18145), .ZN(n18149) );
  AOI22_X1 U21161 ( .A1(n18206), .A2(n18149), .B1(n18218), .B2(n18148), .ZN(
        n18150) );
  OAI211_X1 U21162 ( .C1(n18214), .C2(n18152), .A(n18151), .B(n18150), .ZN(
        P3_U2855) );
  NAND3_X1 U21163 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18153) );
  NOR4_X1 U21164 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18154), .A3(
        n18222), .A4(n18153), .ZN(n18160) );
  AOI21_X1 U21165 ( .B1(n18156), .B2(n18155), .A(n18201), .ZN(n18166) );
  OAI22_X1 U21166 ( .A1(n18166), .A2(n18158), .B1(n18214), .B2(n18157), .ZN(
        n18159) );
  NOR2_X1 U21167 ( .A1(n18160), .A2(n18159), .ZN(n18162) );
  OAI211_X1 U21168 ( .C1(n18163), .C2(n18181), .A(n18162), .B(n18161), .ZN(
        P3_U2856) );
  NAND3_X1 U21169 ( .A1(n18206), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18179), .ZN(n18173) );
  NOR2_X1 U21170 ( .A1(n18173), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18168) );
  INV_X1 U21171 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18165) );
  OAI22_X1 U21172 ( .A1(n18166), .A2(n18165), .B1(n18181), .B2(n18164), .ZN(
        n18167) );
  AOI21_X1 U21173 ( .B1(n18168), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n18167), .ZN(n18170) );
  OAI211_X1 U21174 ( .C1(n18171), .C2(n18214), .A(n18170), .B(n18169), .ZN(
        P3_U2857) );
  OAI21_X1 U21175 ( .B1(n18183), .B2(n18208), .A(n18207), .ZN(n18175) );
  OAI22_X1 U21176 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18173), .B1(
        n18172), .B2(n18181), .ZN(n18174) );
  AOI21_X1 U21177 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18175), .A(
        n18174), .ZN(n18177) );
  NAND2_X1 U21178 ( .A1(n18122), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18176) );
  OAI211_X1 U21179 ( .C1(n18214), .C2(n18178), .A(n18177), .B(n18176), .ZN(
        P3_U2858) );
  OAI21_X1 U21180 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18179), .A(
        n18206), .ZN(n18182) );
  OAI22_X1 U21181 ( .A1(n18183), .A2(n18182), .B1(n18181), .B2(n18180), .ZN(
        n18184) );
  AOI21_X1 U21182 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18201), .A(
        n18184), .ZN(n18186) );
  OAI211_X1 U21183 ( .C1(n18187), .C2(n18214), .A(n18186), .B(n18185), .ZN(
        P3_U2859) );
  OAI21_X1 U21184 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18189), .A(
        n18188), .ZN(n18192) );
  OAI21_X1 U21185 ( .B1(n18843), .B2(n18190), .A(n18193), .ZN(n18191) );
  OAI21_X1 U21186 ( .B1(n18193), .B2(n18192), .A(n18191), .ZN(n18197) );
  OAI21_X1 U21187 ( .B1(n18195), .B2(n18194), .A(n18667), .ZN(n18196) );
  OAI211_X1 U21188 ( .C1(n18199), .C2(n18198), .A(n18197), .B(n18196), .ZN(
        n18200) );
  AOI22_X1 U21189 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18201), .B1(
        n18206), .B2(n18200), .ZN(n18203) );
  OAI211_X1 U21190 ( .C1(n18204), .C2(n18214), .A(n18203), .B(n18202), .ZN(
        P3_U2860) );
  NAND3_X1 U21191 ( .A1(n18206), .A2(n18205), .A3(n18859), .ZN(n18224) );
  AOI21_X1 U21192 ( .B1(n18207), .B2(n18224), .A(n18843), .ZN(n18210) );
  AOI211_X1 U21193 ( .C1(n18673), .C2(n18859), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18208), .ZN(n18209) );
  AOI211_X1 U21194 ( .C1(n18218), .C2(n18211), .A(n18210), .B(n18209), .ZN(
        n18213) );
  NAND2_X1 U21195 ( .A1(n18122), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18212) );
  OAI211_X1 U21196 ( .C1(n18215), .C2(n18214), .A(n18213), .B(n18212), .ZN(
        P3_U2861) );
  INV_X1 U21197 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18869) );
  NOR2_X1 U21198 ( .A1(n18221), .A2(n18869), .ZN(n18216) );
  AOI221_X1 U21199 ( .B1(n18220), .B2(n18219), .C1(n18218), .C2(n18217), .A(
        n18216), .ZN(n18225) );
  OAI211_X1 U21200 ( .C1(n18682), .C2(n18222), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18221), .ZN(n18223) );
  NAND3_X1 U21201 ( .A1(n18225), .A2(n18224), .A3(n18223), .ZN(P3_U2862) );
  OAI211_X1 U21202 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18226), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18726)
         );
  AOI21_X1 U21203 ( .B1(n18726), .B2(n18279), .A(n18227), .ZN(n18228) );
  INV_X1 U21204 ( .A(n18228), .ZN(n18229) );
  OAI221_X1 U21205 ( .B1(n18683), .B2(n18877), .C1(n18683), .C2(n18233), .A(
        n18229), .ZN(P3_U2863) );
  INV_X1 U21206 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18707) );
  NAND2_X1 U21207 ( .A1(n18235), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18506) );
  INV_X1 U21208 ( .A(n18506), .ZN(n18528) );
  NAND2_X1 U21209 ( .A1(n18707), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18391) );
  INV_X1 U21210 ( .A(n18391), .ZN(n18418) );
  NOR2_X1 U21211 ( .A1(n18528), .A2(n18418), .ZN(n18231) );
  OAI22_X1 U21212 ( .A1(n18232), .A2(n18707), .B1(n18231), .B2(n18230), .ZN(
        P3_U2866) );
  NOR2_X1 U21213 ( .A1(n18234), .A2(n18233), .ZN(P3_U2867) );
  NOR2_X1 U21214 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18687) );
  NAND2_X1 U21215 ( .A1(n18235), .A2(n18707), .ZN(n18322) );
  INV_X1 U21216 ( .A(n18322), .ZN(n18324) );
  NAND2_X1 U21217 ( .A1(n18687), .A2(n18324), .ZN(n18299) );
  NOR2_X1 U21218 ( .A1(n18237), .A2(n18236), .ZN(n18273) );
  NAND2_X1 U21219 ( .A1(n18273), .A2(n18238), .ZN(n18612) );
  NAND2_X1 U21220 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18241) );
  NOR2_X1 U21221 ( .A1(n18241), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18607) );
  NAND2_X1 U21222 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18607), .ZN(
        n18577) );
  INV_X1 U21223 ( .A(n18577), .ZN(n18654) );
  AND2_X1 U21224 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18608), .ZN(n18609) );
  AND2_X1 U21225 ( .A1(n18532), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18603) );
  NOR2_X1 U21226 ( .A1(n18707), .A2(n18416), .ZN(n18606) );
  NAND2_X1 U21227 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18606), .ZN(
        n18659) );
  NAND2_X1 U21228 ( .A1(n18659), .A2(n18299), .ZN(n18300) );
  AND2_X1 U21229 ( .A1(n18727), .A2(n18300), .ZN(n18275) );
  AOI22_X1 U21230 ( .A1(n18654), .A2(n18609), .B1(n18603), .B2(n18275), .ZN(
        n18243) );
  NAND2_X1 U21231 ( .A1(n18683), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18482) );
  INV_X1 U21232 ( .A(n18482), .ZN(n18239) );
  NOR2_X1 U21233 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18683), .ZN(
        n18459) );
  NOR2_X1 U21234 ( .A1(n18239), .A2(n18459), .ZN(n18530) );
  NOR2_X1 U21235 ( .A1(n18530), .A2(n18241), .ZN(n18582) );
  AOI21_X1 U21236 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18346), .ZN(n18579) );
  AOI22_X1 U21237 ( .A1(n18608), .A2(n18582), .B1(n18579), .B2(n18300), .ZN(
        n18276) );
  INV_X1 U21238 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18240) );
  NOR2_X2 U21239 ( .A1(n18347), .A2(n18240), .ZN(n18604) );
  NOR2_X2 U21240 ( .A1(n18241), .A2(n18482), .ZN(n18578) );
  AOI22_X1 U21241 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18276), .B1(
        n18604), .B2(n18578), .ZN(n18242) );
  OAI211_X1 U21242 ( .C1(n18299), .C2(n18612), .A(n18243), .B(n18242), .ZN(
        P3_U2868) );
  NAND2_X1 U21243 ( .A1(n18273), .A2(n18244), .ZN(n18618) );
  AND2_X1 U21244 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18608), .ZN(n18615) );
  AND2_X1 U21245 ( .A1(n18532), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18613) );
  AOI22_X1 U21246 ( .A1(n18654), .A2(n18615), .B1(n18275), .B2(n18613), .ZN(
        n18246) );
  NOR2_X2 U21247 ( .A1(n18347), .A2(n14204), .ZN(n18614) );
  AOI22_X1 U21248 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18276), .B1(
        n18578), .B2(n18614), .ZN(n18245) );
  OAI211_X1 U21249 ( .C1(n18299), .C2(n18618), .A(n18246), .B(n18245), .ZN(
        P3_U2869) );
  NAND2_X1 U21250 ( .A1(n18273), .A2(n18247), .ZN(n18624) );
  INV_X1 U21251 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18248) );
  NOR2_X2 U21252 ( .A1(n18347), .A2(n18248), .ZN(n18620) );
  NOR2_X2 U21253 ( .A1(n18346), .A2(n18249), .ZN(n18619) );
  AOI22_X1 U21254 ( .A1(n18578), .A2(n18620), .B1(n18275), .B2(n18619), .ZN(
        n18251) );
  AND2_X1 U21255 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18608), .ZN(n18621) );
  AOI22_X1 U21256 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18276), .B1(
        n18654), .B2(n18621), .ZN(n18250) );
  OAI211_X1 U21257 ( .C1(n18299), .C2(n18624), .A(n18251), .B(n18250), .ZN(
        P3_U2870) );
  NAND2_X1 U21258 ( .A1(n18273), .A2(n18252), .ZN(n18630) );
  INV_X1 U21259 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18253) );
  NOR2_X2 U21260 ( .A1(n18253), .A2(n18347), .ZN(n18625) );
  NOR2_X2 U21261 ( .A1(n18346), .A2(n18254), .ZN(n18626) );
  AOI22_X1 U21262 ( .A1(n18654), .A2(n18625), .B1(n18275), .B2(n18626), .ZN(
        n18256) );
  AND2_X1 U21263 ( .A1(n18608), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18627) );
  AOI22_X1 U21264 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18276), .B1(
        n18578), .B2(n18627), .ZN(n18255) );
  OAI211_X1 U21265 ( .C1(n18299), .C2(n18630), .A(n18256), .B(n18255), .ZN(
        P3_U2871) );
  NAND2_X1 U21266 ( .A1(n18273), .A2(n18257), .ZN(n18636) );
  INV_X1 U21267 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18258) );
  NOR2_X2 U21268 ( .A1(n18258), .A2(n18347), .ZN(n18632) );
  NOR2_X2 U21269 ( .A1(n18346), .A2(n18259), .ZN(n18631) );
  AOI22_X1 U21270 ( .A1(n18654), .A2(n18632), .B1(n18275), .B2(n18631), .ZN(
        n18261) );
  AND2_X1 U21271 ( .A1(n18608), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18633) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18276), .B1(
        n18578), .B2(n18633), .ZN(n18260) );
  OAI211_X1 U21273 ( .C1(n18299), .C2(n18636), .A(n18261), .B(n18260), .ZN(
        P3_U2872) );
  NAND2_X1 U21274 ( .A1(n18273), .A2(n18262), .ZN(n18642) );
  NOR2_X2 U21275 ( .A1(n18347), .A2(n19279), .ZN(n18639) );
  NOR2_X2 U21276 ( .A1(n18346), .A2(n18263), .ZN(n18637) );
  AOI22_X1 U21277 ( .A1(n18578), .A2(n18639), .B1(n18275), .B2(n18637), .ZN(
        n18266) );
  INV_X1 U21278 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18264) );
  NOR2_X2 U21279 ( .A1(n18264), .A2(n18347), .ZN(n18638) );
  AOI22_X1 U21280 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18276), .B1(
        n18654), .B2(n18638), .ZN(n18265) );
  OAI211_X1 U21281 ( .C1(n18299), .C2(n18642), .A(n18266), .B(n18265), .ZN(
        P3_U2873) );
  NAND2_X1 U21282 ( .A1(n18273), .A2(n18267), .ZN(n18648) );
  INV_X1 U21283 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18268) );
  NOR2_X2 U21284 ( .A1(n18268), .A2(n18347), .ZN(n18645) );
  NOR2_X2 U21285 ( .A1(n18269), .A2(n18346), .ZN(n18643) );
  AOI22_X1 U21286 ( .A1(n18578), .A2(n18645), .B1(n18275), .B2(n18643), .ZN(
        n18271) );
  NOR2_X2 U21287 ( .A1(n19282), .A2(n18347), .ZN(n18644) );
  AOI22_X1 U21288 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18276), .B1(
        n18654), .B2(n18644), .ZN(n18270) );
  OAI211_X1 U21289 ( .C1(n18299), .C2(n18648), .A(n18271), .B(n18270), .ZN(
        P3_U2874) );
  NAND2_X1 U21290 ( .A1(n18273), .A2(n18272), .ZN(n18658) );
  NOR2_X2 U21291 ( .A1(n18347), .A2(n19289), .ZN(n18650) );
  NOR2_X2 U21292 ( .A1(n18274), .A2(n18346), .ZN(n18652) );
  AOI22_X1 U21293 ( .A1(n18654), .A2(n18650), .B1(n18275), .B2(n18652), .ZN(
        n18278) );
  NOR2_X2 U21294 ( .A1(n15048), .A2(n18347), .ZN(n18653) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18276), .B1(
        n18578), .B2(n18653), .ZN(n18277) );
  OAI211_X1 U21296 ( .C1(n18299), .C2(n18658), .A(n18278), .B(n18277), .ZN(
        P3_U2875) );
  NAND2_X1 U21297 ( .A1(n18324), .A2(n18459), .ZN(n18325) );
  INV_X1 U21298 ( .A(n18659), .ZN(n18317) );
  NAND2_X1 U21299 ( .A1(n18684), .A2(n18727), .ZN(n18461) );
  NOR2_X1 U21300 ( .A1(n18322), .A2(n18461), .ZN(n18295) );
  AOI22_X1 U21301 ( .A1(n18317), .A2(n18604), .B1(n18603), .B2(n18295), .ZN(
        n18282) );
  INV_X1 U21302 ( .A(n18279), .ZN(n18280) );
  NOR2_X1 U21303 ( .A1(n18346), .A2(n18280), .ZN(n18605) );
  INV_X1 U21304 ( .A(n18605), .ZN(n18323) );
  NOR2_X1 U21305 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18323), .ZN(
        n18370) );
  AOI22_X1 U21306 ( .A1(n18608), .A2(n18606), .B1(n18324), .B2(n18370), .ZN(
        n18296) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18296), .B1(
        n18578), .B2(n18609), .ZN(n18281) );
  OAI211_X1 U21308 ( .C1(n18612), .C2(n18325), .A(n18282), .B(n18281), .ZN(
        P3_U2876) );
  AOI22_X1 U21309 ( .A1(n18317), .A2(n18614), .B1(n18613), .B2(n18295), .ZN(
        n18284) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18296), .B1(
        n18578), .B2(n18615), .ZN(n18283) );
  OAI211_X1 U21311 ( .C1(n18618), .C2(n18325), .A(n18284), .B(n18283), .ZN(
        P3_U2877) );
  AOI22_X1 U21312 ( .A1(n18317), .A2(n18620), .B1(n18619), .B2(n18295), .ZN(
        n18286) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18296), .B1(
        n18578), .B2(n18621), .ZN(n18285) );
  OAI211_X1 U21314 ( .C1(n18624), .C2(n18325), .A(n18286), .B(n18285), .ZN(
        P3_U2878) );
  AOI22_X1 U21315 ( .A1(n18578), .A2(n18625), .B1(n18626), .B2(n18295), .ZN(
        n18288) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18296), .B1(
        n18317), .B2(n18627), .ZN(n18287) );
  OAI211_X1 U21317 ( .C1(n18630), .C2(n18325), .A(n18288), .B(n18287), .ZN(
        P3_U2879) );
  AOI22_X1 U21318 ( .A1(n18317), .A2(n18633), .B1(n18631), .B2(n18295), .ZN(
        n18290) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18296), .B1(
        n18578), .B2(n18632), .ZN(n18289) );
  OAI211_X1 U21320 ( .C1(n18636), .C2(n18325), .A(n18290), .B(n18289), .ZN(
        P3_U2880) );
  AOI22_X1 U21321 ( .A1(n18578), .A2(n18638), .B1(n18637), .B2(n18295), .ZN(
        n18292) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18296), .B1(
        n18317), .B2(n18639), .ZN(n18291) );
  OAI211_X1 U21323 ( .C1(n18642), .C2(n18325), .A(n18292), .B(n18291), .ZN(
        P3_U2881) );
  AOI22_X1 U21324 ( .A1(n18317), .A2(n18645), .B1(n18643), .B2(n18295), .ZN(
        n18294) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18296), .B1(
        n18578), .B2(n18644), .ZN(n18293) );
  OAI211_X1 U21326 ( .C1(n18648), .C2(n18325), .A(n18294), .B(n18293), .ZN(
        P3_U2882) );
  AOI22_X1 U21327 ( .A1(n18317), .A2(n18653), .B1(n18652), .B2(n18295), .ZN(
        n18298) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18296), .B1(
        n18578), .B2(n18650), .ZN(n18297) );
  OAI211_X1 U21329 ( .C1(n18658), .C2(n18325), .A(n18298), .B(n18297), .ZN(
        P3_U2883) );
  NOR2_X2 U21330 ( .A1(n18322), .A2(n18482), .ZN(n18386) );
  INV_X1 U21331 ( .A(n18386), .ZN(n18321) );
  INV_X1 U21332 ( .A(n18299), .ZN(n18341) );
  NAND2_X1 U21333 ( .A1(n18325), .A2(n18321), .ZN(n18301) );
  INV_X1 U21334 ( .A(n18301), .ZN(n18348) );
  NOR2_X1 U21335 ( .A1(n18556), .A2(n18348), .ZN(n18316) );
  AOI22_X1 U21336 ( .A1(n18341), .A2(n18604), .B1(n18603), .B2(n18316), .ZN(
        n18303) );
  OAI221_X1 U21337 ( .B1(n18301), .B2(n18581), .C1(n18301), .C2(n18300), .A(
        n18579), .ZN(n18318) );
  AOI22_X1 U21338 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18318), .B1(
        n18317), .B2(n18609), .ZN(n18302) );
  OAI211_X1 U21339 ( .C1(n18612), .C2(n18321), .A(n18303), .B(n18302), .ZN(
        P3_U2884) );
  AOI22_X1 U21340 ( .A1(n18341), .A2(n18614), .B1(n18613), .B2(n18316), .ZN(
        n18305) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18318), .B1(
        n18317), .B2(n18615), .ZN(n18304) );
  OAI211_X1 U21342 ( .C1(n18618), .C2(n18321), .A(n18305), .B(n18304), .ZN(
        P3_U2885) );
  AOI22_X1 U21343 ( .A1(n18317), .A2(n18621), .B1(n18619), .B2(n18316), .ZN(
        n18307) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18318), .B1(
        n18341), .B2(n18620), .ZN(n18306) );
  OAI211_X1 U21345 ( .C1(n18624), .C2(n18321), .A(n18307), .B(n18306), .ZN(
        P3_U2886) );
  AOI22_X1 U21346 ( .A1(n18317), .A2(n18625), .B1(n18626), .B2(n18316), .ZN(
        n18309) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18318), .B1(
        n18341), .B2(n18627), .ZN(n18308) );
  OAI211_X1 U21348 ( .C1(n18630), .C2(n18321), .A(n18309), .B(n18308), .ZN(
        P3_U2887) );
  AOI22_X1 U21349 ( .A1(n18317), .A2(n18632), .B1(n18631), .B2(n18316), .ZN(
        n18311) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18318), .B1(
        n18341), .B2(n18633), .ZN(n18310) );
  OAI211_X1 U21351 ( .C1(n18636), .C2(n18321), .A(n18311), .B(n18310), .ZN(
        P3_U2888) );
  AOI22_X1 U21352 ( .A1(n18317), .A2(n18638), .B1(n18637), .B2(n18316), .ZN(
        n18313) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18318), .B1(
        n18341), .B2(n18639), .ZN(n18312) );
  OAI211_X1 U21354 ( .C1(n18642), .C2(n18321), .A(n18313), .B(n18312), .ZN(
        P3_U2889) );
  AOI22_X1 U21355 ( .A1(n18317), .A2(n18644), .B1(n18643), .B2(n18316), .ZN(
        n18315) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18318), .B1(
        n18341), .B2(n18645), .ZN(n18314) );
  OAI211_X1 U21357 ( .C1(n18648), .C2(n18321), .A(n18315), .B(n18314), .ZN(
        P3_U2890) );
  AOI22_X1 U21358 ( .A1(n18341), .A2(n18653), .B1(n18652), .B2(n18316), .ZN(
        n18320) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18318), .B1(
        n18317), .B2(n18650), .ZN(n18319) );
  OAI211_X1 U21360 ( .C1(n18658), .C2(n18321), .A(n18320), .B(n18319), .ZN(
        P3_U2891) );
  NOR2_X1 U21361 ( .A1(n18684), .A2(n18322), .ZN(n18371) );
  NAND2_X1 U21362 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18371), .ZN(
        n18345) );
  AND2_X1 U21363 ( .A1(n18727), .A2(n18371), .ZN(n18340) );
  AOI22_X1 U21364 ( .A1(n18341), .A2(n18609), .B1(n18603), .B2(n18340), .ZN(
        n18327) );
  AOI21_X1 U21365 ( .B1(n18684), .B2(n18393), .A(n18323), .ZN(n18417) );
  NAND2_X1 U21366 ( .A1(n18324), .A2(n18417), .ZN(n18342) );
  INV_X1 U21367 ( .A(n18325), .ZN(n18365) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18342), .B1(
        n18604), .B2(n18365), .ZN(n18326) );
  OAI211_X1 U21369 ( .C1(n18612), .C2(n18345), .A(n18327), .B(n18326), .ZN(
        P3_U2892) );
  AOI22_X1 U21370 ( .A1(n18614), .A2(n18365), .B1(n18613), .B2(n18340), .ZN(
        n18329) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18342), .B1(
        n18341), .B2(n18615), .ZN(n18328) );
  OAI211_X1 U21372 ( .C1(n18618), .C2(n18345), .A(n18329), .B(n18328), .ZN(
        P3_U2893) );
  AOI22_X1 U21373 ( .A1(n18341), .A2(n18621), .B1(n18619), .B2(n18340), .ZN(
        n18331) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18342), .B1(
        n18620), .B2(n18365), .ZN(n18330) );
  OAI211_X1 U21375 ( .C1(n18624), .C2(n18345), .A(n18331), .B(n18330), .ZN(
        P3_U2894) );
  AOI22_X1 U21376 ( .A1(n18341), .A2(n18625), .B1(n18626), .B2(n18340), .ZN(
        n18333) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18342), .B1(
        n18627), .B2(n18365), .ZN(n18332) );
  OAI211_X1 U21378 ( .C1(n18630), .C2(n18345), .A(n18333), .B(n18332), .ZN(
        P3_U2895) );
  AOI22_X1 U21379 ( .A1(n18633), .A2(n18365), .B1(n18631), .B2(n18340), .ZN(
        n18335) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18342), .B1(
        n18341), .B2(n18632), .ZN(n18334) );
  OAI211_X1 U21381 ( .C1(n18636), .C2(n18345), .A(n18335), .B(n18334), .ZN(
        P3_U2896) );
  AOI22_X1 U21382 ( .A1(n18341), .A2(n18638), .B1(n18637), .B2(n18340), .ZN(
        n18337) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18342), .B1(
        n18639), .B2(n18365), .ZN(n18336) );
  OAI211_X1 U21384 ( .C1(n18642), .C2(n18345), .A(n18337), .B(n18336), .ZN(
        P3_U2897) );
  AOI22_X1 U21385 ( .A1(n18341), .A2(n18644), .B1(n18643), .B2(n18340), .ZN(
        n18339) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18342), .B1(
        n18645), .B2(n18365), .ZN(n18338) );
  OAI211_X1 U21387 ( .C1(n18648), .C2(n18345), .A(n18339), .B(n18338), .ZN(
        P3_U2898) );
  AOI22_X1 U21388 ( .A1(n18341), .A2(n18650), .B1(n18652), .B2(n18340), .ZN(
        n18344) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18342), .B1(
        n18653), .B2(n18365), .ZN(n18343) );
  OAI211_X1 U21390 ( .C1(n18658), .C2(n18345), .A(n18344), .B(n18343), .ZN(
        P3_U2899) );
  NAND2_X1 U21391 ( .A1(n18687), .A2(n18418), .ZN(n18369) );
  INV_X1 U21392 ( .A(n18345), .ZN(n18411) );
  INV_X1 U21393 ( .A(n18369), .ZN(n18435) );
  NOR2_X1 U21394 ( .A1(n18411), .A2(n18435), .ZN(n18394) );
  NOR2_X1 U21395 ( .A1(n18556), .A2(n18394), .ZN(n18364) );
  AOI22_X1 U21396 ( .A1(n18604), .A2(n18386), .B1(n18603), .B2(n18364), .ZN(
        n18351) );
  OAI22_X1 U21397 ( .A1(n18348), .A2(n18347), .B1(n18394), .B2(n18346), .ZN(
        n18349) );
  OAI21_X1 U21398 ( .B1(n18435), .B2(n18832), .A(n18349), .ZN(n18366) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18366), .B1(
        n18609), .B2(n18365), .ZN(n18350) );
  OAI211_X1 U21400 ( .C1(n18612), .C2(n18369), .A(n18351), .B(n18350), .ZN(
        P3_U2900) );
  AOI22_X1 U21401 ( .A1(n18615), .A2(n18365), .B1(n18613), .B2(n18364), .ZN(
        n18353) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18366), .B1(
        n18614), .B2(n18386), .ZN(n18352) );
  OAI211_X1 U21403 ( .C1(n18618), .C2(n18369), .A(n18353), .B(n18352), .ZN(
        P3_U2901) );
  AOI22_X1 U21404 ( .A1(n18620), .A2(n18386), .B1(n18619), .B2(n18364), .ZN(
        n18355) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18366), .B1(
        n18621), .B2(n18365), .ZN(n18354) );
  OAI211_X1 U21406 ( .C1(n18624), .C2(n18369), .A(n18355), .B(n18354), .ZN(
        P3_U2902) );
  AOI22_X1 U21407 ( .A1(n18626), .A2(n18364), .B1(n18625), .B2(n18365), .ZN(
        n18357) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18366), .B1(
        n18627), .B2(n18386), .ZN(n18356) );
  OAI211_X1 U21409 ( .C1(n18630), .C2(n18369), .A(n18357), .B(n18356), .ZN(
        P3_U2903) );
  AOI22_X1 U21410 ( .A1(n18632), .A2(n18365), .B1(n18631), .B2(n18364), .ZN(
        n18359) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18366), .B1(
        n18633), .B2(n18386), .ZN(n18358) );
  OAI211_X1 U21412 ( .C1(n18636), .C2(n18369), .A(n18359), .B(n18358), .ZN(
        P3_U2904) );
  AOI22_X1 U21413 ( .A1(n18639), .A2(n18386), .B1(n18637), .B2(n18364), .ZN(
        n18361) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18366), .B1(
        n18638), .B2(n18365), .ZN(n18360) );
  OAI211_X1 U21415 ( .C1(n18642), .C2(n18369), .A(n18361), .B(n18360), .ZN(
        P3_U2905) );
  AOI22_X1 U21416 ( .A1(n18644), .A2(n18365), .B1(n18643), .B2(n18364), .ZN(
        n18363) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18366), .B1(
        n18645), .B2(n18386), .ZN(n18362) );
  OAI211_X1 U21418 ( .C1(n18648), .C2(n18369), .A(n18363), .B(n18362), .ZN(
        P3_U2906) );
  AOI22_X1 U21419 ( .A1(n18653), .A2(n18386), .B1(n18652), .B2(n18364), .ZN(
        n18368) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18366), .B1(
        n18650), .B2(n18365), .ZN(n18367) );
  OAI211_X1 U21421 ( .C1(n18658), .C2(n18369), .A(n18368), .B(n18367), .ZN(
        P3_U2907) );
  NAND2_X1 U21422 ( .A1(n18418), .A2(n18459), .ZN(n18419) );
  NOR2_X1 U21423 ( .A1(n18391), .A2(n18461), .ZN(n18387) );
  AOI22_X1 U21424 ( .A1(n18604), .A2(n18411), .B1(n18603), .B2(n18387), .ZN(
        n18373) );
  AOI22_X1 U21425 ( .A1(n18608), .A2(n18371), .B1(n18418), .B2(n18370), .ZN(
        n18388) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18388), .B1(
        n18609), .B2(n18386), .ZN(n18372) );
  OAI211_X1 U21427 ( .C1(n18612), .C2(n18419), .A(n18373), .B(n18372), .ZN(
        P3_U2908) );
  AOI22_X1 U21428 ( .A1(n18615), .A2(n18386), .B1(n18613), .B2(n18387), .ZN(
        n18375) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18388), .B1(
        n18614), .B2(n18411), .ZN(n18374) );
  OAI211_X1 U21430 ( .C1(n18618), .C2(n18419), .A(n18375), .B(n18374), .ZN(
        P3_U2909) );
  AOI22_X1 U21431 ( .A1(n18620), .A2(n18411), .B1(n18619), .B2(n18387), .ZN(
        n18377) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18388), .B1(
        n18621), .B2(n18386), .ZN(n18376) );
  OAI211_X1 U21433 ( .C1(n18624), .C2(n18419), .A(n18377), .B(n18376), .ZN(
        P3_U2910) );
  AOI22_X1 U21434 ( .A1(n18626), .A2(n18387), .B1(n18625), .B2(n18386), .ZN(
        n18379) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18388), .B1(
        n18627), .B2(n18411), .ZN(n18378) );
  OAI211_X1 U21436 ( .C1(n18630), .C2(n18419), .A(n18379), .B(n18378), .ZN(
        P3_U2911) );
  AOI22_X1 U21437 ( .A1(n18632), .A2(n18386), .B1(n18631), .B2(n18387), .ZN(
        n18381) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18388), .B1(
        n18633), .B2(n18411), .ZN(n18380) );
  OAI211_X1 U21439 ( .C1(n18636), .C2(n18419), .A(n18381), .B(n18380), .ZN(
        P3_U2912) );
  AOI22_X1 U21440 ( .A1(n18638), .A2(n18386), .B1(n18637), .B2(n18387), .ZN(
        n18383) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18388), .B1(
        n18639), .B2(n18411), .ZN(n18382) );
  OAI211_X1 U21442 ( .C1(n18642), .C2(n18419), .A(n18383), .B(n18382), .ZN(
        P3_U2913) );
  AOI22_X1 U21443 ( .A1(n18645), .A2(n18411), .B1(n18643), .B2(n18387), .ZN(
        n18385) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18388), .B1(
        n18644), .B2(n18386), .ZN(n18384) );
  OAI211_X1 U21445 ( .C1(n18648), .C2(n18419), .A(n18385), .B(n18384), .ZN(
        P3_U2914) );
  AOI22_X1 U21446 ( .A1(n18652), .A2(n18387), .B1(n18650), .B2(n18386), .ZN(
        n18390) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18388), .B1(
        n18653), .B2(n18411), .ZN(n18389) );
  OAI211_X1 U21448 ( .C1(n18658), .C2(n18419), .A(n18390), .B(n18389), .ZN(
        P3_U2915) );
  NOR2_X2 U21449 ( .A1(n18391), .A2(n18482), .ZN(n18477) );
  INV_X1 U21450 ( .A(n18477), .ZN(n18415) );
  NAND2_X1 U21451 ( .A1(n18419), .A2(n18415), .ZN(n18439) );
  INV_X1 U21452 ( .A(n18439), .ZN(n18392) );
  NOR2_X1 U21453 ( .A1(n18556), .A2(n18392), .ZN(n18410) );
  AOI22_X1 U21454 ( .A1(n18609), .A2(n18411), .B1(n18603), .B2(n18410), .ZN(
        n18397) );
  OAI21_X1 U21455 ( .B1(n18394), .B2(n18393), .A(n18392), .ZN(n18395) );
  OAI211_X1 U21456 ( .C1(n18477), .C2(n18832), .A(n18532), .B(n18395), .ZN(
        n18412) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18412), .B1(
        n18604), .B2(n18435), .ZN(n18396) );
  OAI211_X1 U21458 ( .C1(n18612), .C2(n18415), .A(n18397), .B(n18396), .ZN(
        P3_U2916) );
  AOI22_X1 U21459 ( .A1(n18614), .A2(n18435), .B1(n18613), .B2(n18410), .ZN(
        n18399) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18412), .B1(
        n18615), .B2(n18411), .ZN(n18398) );
  OAI211_X1 U21461 ( .C1(n18618), .C2(n18415), .A(n18399), .B(n18398), .ZN(
        P3_U2917) );
  AOI22_X1 U21462 ( .A1(n18621), .A2(n18411), .B1(n18619), .B2(n18410), .ZN(
        n18401) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18412), .B1(
        n18620), .B2(n18435), .ZN(n18400) );
  OAI211_X1 U21464 ( .C1(n18624), .C2(n18415), .A(n18401), .B(n18400), .ZN(
        P3_U2918) );
  AOI22_X1 U21465 ( .A1(n18626), .A2(n18410), .B1(n18625), .B2(n18411), .ZN(
        n18403) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18412), .B1(
        n18627), .B2(n18435), .ZN(n18402) );
  OAI211_X1 U21467 ( .C1(n18630), .C2(n18415), .A(n18403), .B(n18402), .ZN(
        P3_U2919) );
  AOI22_X1 U21468 ( .A1(n18632), .A2(n18411), .B1(n18631), .B2(n18410), .ZN(
        n18405) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18412), .B1(
        n18633), .B2(n18435), .ZN(n18404) );
  OAI211_X1 U21470 ( .C1(n18636), .C2(n18415), .A(n18405), .B(n18404), .ZN(
        P3_U2920) );
  AOI22_X1 U21471 ( .A1(n18638), .A2(n18411), .B1(n18637), .B2(n18410), .ZN(
        n18407) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18412), .B1(
        n18639), .B2(n18435), .ZN(n18406) );
  OAI211_X1 U21473 ( .C1(n18642), .C2(n18415), .A(n18407), .B(n18406), .ZN(
        P3_U2921) );
  AOI22_X1 U21474 ( .A1(n18644), .A2(n18411), .B1(n18643), .B2(n18410), .ZN(
        n18409) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18412), .B1(
        n18645), .B2(n18435), .ZN(n18408) );
  OAI211_X1 U21476 ( .C1(n18648), .C2(n18415), .A(n18409), .B(n18408), .ZN(
        P3_U2922) );
  AOI22_X1 U21477 ( .A1(n18653), .A2(n18435), .B1(n18652), .B2(n18410), .ZN(
        n18414) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18412), .B1(
        n18650), .B2(n18411), .ZN(n18413) );
  OAI211_X1 U21479 ( .C1(n18658), .C2(n18415), .A(n18414), .B(n18413), .ZN(
        P3_U2923) );
  NOR2_X1 U21480 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18416), .ZN(
        n18462) );
  NAND2_X1 U21481 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18462), .ZN(
        n18460) );
  AND2_X1 U21482 ( .A1(n18727), .A2(n18462), .ZN(n18434) );
  AOI22_X1 U21483 ( .A1(n18609), .A2(n18435), .B1(n18603), .B2(n18434), .ZN(
        n18421) );
  NAND2_X1 U21484 ( .A1(n18418), .A2(n18417), .ZN(n18436) );
  INV_X1 U21485 ( .A(n18419), .ZN(n18454) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18436), .B1(
        n18604), .B2(n18454), .ZN(n18420) );
  OAI211_X1 U21487 ( .C1(n18612), .C2(n18460), .A(n18421), .B(n18420), .ZN(
        P3_U2924) );
  AOI22_X1 U21488 ( .A1(n18615), .A2(n18435), .B1(n18613), .B2(n18434), .ZN(
        n18423) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18436), .B1(
        n18614), .B2(n18454), .ZN(n18422) );
  OAI211_X1 U21490 ( .C1(n18618), .C2(n18460), .A(n18423), .B(n18422), .ZN(
        P3_U2925) );
  AOI22_X1 U21491 ( .A1(n18621), .A2(n18435), .B1(n18619), .B2(n18434), .ZN(
        n18425) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18436), .B1(
        n18620), .B2(n18454), .ZN(n18424) );
  OAI211_X1 U21493 ( .C1(n18624), .C2(n18460), .A(n18425), .B(n18424), .ZN(
        P3_U2926) );
  AOI22_X1 U21494 ( .A1(n18627), .A2(n18454), .B1(n18626), .B2(n18434), .ZN(
        n18427) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18436), .B1(
        n18625), .B2(n18435), .ZN(n18426) );
  OAI211_X1 U21496 ( .C1(n18630), .C2(n18460), .A(n18427), .B(n18426), .ZN(
        P3_U2927) );
  AOI22_X1 U21497 ( .A1(n18632), .A2(n18435), .B1(n18631), .B2(n18434), .ZN(
        n18429) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18436), .B1(
        n18633), .B2(n18454), .ZN(n18428) );
  OAI211_X1 U21499 ( .C1(n18636), .C2(n18460), .A(n18429), .B(n18428), .ZN(
        P3_U2928) );
  AOI22_X1 U21500 ( .A1(n18639), .A2(n18454), .B1(n18637), .B2(n18434), .ZN(
        n18431) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18436), .B1(
        n18638), .B2(n18435), .ZN(n18430) );
  OAI211_X1 U21502 ( .C1(n18642), .C2(n18460), .A(n18431), .B(n18430), .ZN(
        P3_U2929) );
  AOI22_X1 U21503 ( .A1(n18644), .A2(n18435), .B1(n18643), .B2(n18434), .ZN(
        n18433) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18436), .B1(
        n18645), .B2(n18454), .ZN(n18432) );
  OAI211_X1 U21505 ( .C1(n18648), .C2(n18460), .A(n18433), .B(n18432), .ZN(
        P3_U2930) );
  AOI22_X1 U21506 ( .A1(n18653), .A2(n18454), .B1(n18652), .B2(n18434), .ZN(
        n18438) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18436), .B1(
        n18650), .B2(n18435), .ZN(n18437) );
  OAI211_X1 U21508 ( .C1(n18658), .C2(n18460), .A(n18438), .B(n18437), .ZN(
        P3_U2931) );
  NAND2_X1 U21509 ( .A1(n18687), .A2(n18528), .ZN(n18483) );
  NAND2_X1 U21510 ( .A1(n18460), .A2(n18483), .ZN(n18484) );
  AND2_X1 U21511 ( .A1(n18727), .A2(n18484), .ZN(n18455) );
  AOI22_X1 U21512 ( .A1(n18609), .A2(n18454), .B1(n18603), .B2(n18455), .ZN(
        n18441) );
  OAI221_X1 U21513 ( .B1(n18484), .B2(n18581), .C1(n18484), .C2(n18439), .A(
        n18579), .ZN(n18456) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18456), .B1(
        n18604), .B2(n18477), .ZN(n18440) );
  OAI211_X1 U21515 ( .C1(n18612), .C2(n18483), .A(n18441), .B(n18440), .ZN(
        P3_U2932) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18456), .B1(
        n18613), .B2(n18455), .ZN(n18443) );
  AOI22_X1 U21517 ( .A1(n18614), .A2(n18477), .B1(n18615), .B2(n18454), .ZN(
        n18442) );
  OAI211_X1 U21518 ( .C1(n18618), .C2(n18483), .A(n18443), .B(n18442), .ZN(
        P3_U2933) );
  AOI22_X1 U21519 ( .A1(n18620), .A2(n18477), .B1(n18619), .B2(n18455), .ZN(
        n18445) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18456), .B1(
        n18621), .B2(n18454), .ZN(n18444) );
  OAI211_X1 U21521 ( .C1(n18624), .C2(n18483), .A(n18445), .B(n18444), .ZN(
        P3_U2934) );
  AOI22_X1 U21522 ( .A1(n18627), .A2(n18477), .B1(n18626), .B2(n18455), .ZN(
        n18447) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18456), .B1(
        n18625), .B2(n18454), .ZN(n18446) );
  OAI211_X1 U21524 ( .C1(n18630), .C2(n18483), .A(n18447), .B(n18446), .ZN(
        P3_U2935) );
  AOI22_X1 U21525 ( .A1(n18633), .A2(n18477), .B1(n18631), .B2(n18455), .ZN(
        n18449) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18456), .B1(
        n18632), .B2(n18454), .ZN(n18448) );
  OAI211_X1 U21527 ( .C1(n18636), .C2(n18483), .A(n18449), .B(n18448), .ZN(
        P3_U2936) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18456), .B1(
        n18637), .B2(n18455), .ZN(n18451) );
  AOI22_X1 U21529 ( .A1(n18638), .A2(n18454), .B1(n18639), .B2(n18477), .ZN(
        n18450) );
  OAI211_X1 U21530 ( .C1(n18642), .C2(n18483), .A(n18451), .B(n18450), .ZN(
        P3_U2937) );
  AOI22_X1 U21531 ( .A1(n18645), .A2(n18477), .B1(n18643), .B2(n18455), .ZN(
        n18453) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18456), .B1(
        n18644), .B2(n18454), .ZN(n18452) );
  OAI211_X1 U21533 ( .C1(n18648), .C2(n18483), .A(n18453), .B(n18452), .ZN(
        P3_U2938) );
  AOI22_X1 U21534 ( .A1(n18652), .A2(n18455), .B1(n18650), .B2(n18454), .ZN(
        n18458) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18456), .B1(
        n18653), .B2(n18477), .ZN(n18457) );
  OAI211_X1 U21536 ( .C1(n18658), .C2(n18483), .A(n18458), .B(n18457), .ZN(
        P3_U2939) );
  NAND2_X1 U21537 ( .A1(n18528), .A2(n18459), .ZN(n18507) );
  INV_X1 U21538 ( .A(n18460), .ZN(n18501) );
  NOR2_X1 U21539 ( .A1(n18506), .A2(n18461), .ZN(n18478) );
  AOI22_X1 U21540 ( .A1(n18604), .A2(n18501), .B1(n18603), .B2(n18478), .ZN(
        n18464) );
  NOR2_X1 U21541 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18506), .ZN(
        n18508) );
  AOI22_X1 U21542 ( .A1(n18608), .A2(n18462), .B1(n18605), .B2(n18508), .ZN(
        n18479) );
  AOI22_X1 U21543 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18479), .B1(
        n18609), .B2(n18477), .ZN(n18463) );
  OAI211_X1 U21544 ( .C1(n18612), .C2(n18507), .A(n18464), .B(n18463), .ZN(
        P3_U2940) );
  AOI22_X1 U21545 ( .A1(n18615), .A2(n18477), .B1(n18613), .B2(n18478), .ZN(
        n18466) );
  AOI22_X1 U21546 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18479), .B1(
        n18614), .B2(n18501), .ZN(n18465) );
  OAI211_X1 U21547 ( .C1(n18618), .C2(n18507), .A(n18466), .B(n18465), .ZN(
        P3_U2941) );
  AOI22_X1 U21548 ( .A1(n18621), .A2(n18477), .B1(n18619), .B2(n18478), .ZN(
        n18468) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18479), .B1(
        n18620), .B2(n18501), .ZN(n18467) );
  OAI211_X1 U21550 ( .C1(n18624), .C2(n18507), .A(n18468), .B(n18467), .ZN(
        P3_U2942) );
  AOI22_X1 U21551 ( .A1(n18626), .A2(n18478), .B1(n18625), .B2(n18477), .ZN(
        n18470) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18479), .B1(
        n18627), .B2(n18501), .ZN(n18469) );
  OAI211_X1 U21553 ( .C1(n18630), .C2(n18507), .A(n18470), .B(n18469), .ZN(
        P3_U2943) );
  AOI22_X1 U21554 ( .A1(n18632), .A2(n18477), .B1(n18631), .B2(n18478), .ZN(
        n18472) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18479), .B1(
        n18633), .B2(n18501), .ZN(n18471) );
  OAI211_X1 U21556 ( .C1(n18636), .C2(n18507), .A(n18472), .B(n18471), .ZN(
        P3_U2944) );
  AOI22_X1 U21557 ( .A1(n18638), .A2(n18477), .B1(n18637), .B2(n18478), .ZN(
        n18474) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18479), .B1(
        n18639), .B2(n18501), .ZN(n18473) );
  OAI211_X1 U21559 ( .C1(n18642), .C2(n18507), .A(n18474), .B(n18473), .ZN(
        P3_U2945) );
  AOI22_X1 U21560 ( .A1(n18645), .A2(n18501), .B1(n18643), .B2(n18478), .ZN(
        n18476) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18479), .B1(
        n18644), .B2(n18477), .ZN(n18475) );
  OAI211_X1 U21562 ( .C1(n18648), .C2(n18507), .A(n18476), .B(n18475), .ZN(
        P3_U2946) );
  AOI22_X1 U21563 ( .A1(n18652), .A2(n18478), .B1(n18650), .B2(n18477), .ZN(
        n18481) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18479), .B1(
        n18653), .B2(n18501), .ZN(n18480) );
  OAI211_X1 U21565 ( .C1(n18658), .C2(n18507), .A(n18481), .B(n18480), .ZN(
        P3_U2947) );
  NOR2_X2 U21566 ( .A1(n18506), .A2(n18482), .ZN(n18573) );
  INV_X1 U21567 ( .A(n18573), .ZN(n18505) );
  INV_X1 U21568 ( .A(n18483), .ZN(n18523) );
  AOI21_X1 U21569 ( .B1(n18507), .B2(n18505), .A(n18556), .ZN(n18500) );
  AOI22_X1 U21570 ( .A1(n18604), .A2(n18523), .B1(n18603), .B2(n18500), .ZN(
        n18487) );
  NAND2_X1 U21571 ( .A1(n18507), .A2(n18505), .ZN(n18485) );
  OAI221_X1 U21572 ( .B1(n18485), .B2(n18581), .C1(n18485), .C2(n18484), .A(
        n18579), .ZN(n18502) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18502), .B1(
        n18609), .B2(n18501), .ZN(n18486) );
  OAI211_X1 U21574 ( .C1(n18612), .C2(n18505), .A(n18487), .B(n18486), .ZN(
        P3_U2948) );
  AOI22_X1 U21575 ( .A1(n18615), .A2(n18501), .B1(n18613), .B2(n18500), .ZN(
        n18489) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18502), .B1(
        n18614), .B2(n18523), .ZN(n18488) );
  OAI211_X1 U21577 ( .C1(n18618), .C2(n18505), .A(n18489), .B(n18488), .ZN(
        P3_U2949) );
  AOI22_X1 U21578 ( .A1(n18620), .A2(n18523), .B1(n18619), .B2(n18500), .ZN(
        n18491) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18502), .B1(
        n18621), .B2(n18501), .ZN(n18490) );
  OAI211_X1 U21580 ( .C1(n18624), .C2(n18505), .A(n18491), .B(n18490), .ZN(
        P3_U2950) );
  AOI22_X1 U21581 ( .A1(n18627), .A2(n18523), .B1(n18626), .B2(n18500), .ZN(
        n18493) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18502), .B1(
        n18625), .B2(n18501), .ZN(n18492) );
  OAI211_X1 U21583 ( .C1(n18630), .C2(n18505), .A(n18493), .B(n18492), .ZN(
        P3_U2951) );
  AOI22_X1 U21584 ( .A1(n18633), .A2(n18523), .B1(n18631), .B2(n18500), .ZN(
        n18495) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18502), .B1(
        n18632), .B2(n18501), .ZN(n18494) );
  OAI211_X1 U21586 ( .C1(n18636), .C2(n18505), .A(n18495), .B(n18494), .ZN(
        P3_U2952) );
  AOI22_X1 U21587 ( .A1(n18638), .A2(n18501), .B1(n18637), .B2(n18500), .ZN(
        n18497) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18502), .B1(
        n18639), .B2(n18523), .ZN(n18496) );
  OAI211_X1 U21589 ( .C1(n18642), .C2(n18505), .A(n18497), .B(n18496), .ZN(
        P3_U2953) );
  AOI22_X1 U21590 ( .A1(n18645), .A2(n18523), .B1(n18643), .B2(n18500), .ZN(
        n18499) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18502), .B1(
        n18644), .B2(n18501), .ZN(n18498) );
  OAI211_X1 U21592 ( .C1(n18648), .C2(n18505), .A(n18499), .B(n18498), .ZN(
        P3_U2954) );
  AOI22_X1 U21593 ( .A1(n18653), .A2(n18523), .B1(n18652), .B2(n18500), .ZN(
        n18504) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18502), .B1(
        n18650), .B2(n18501), .ZN(n18503) );
  OAI211_X1 U21595 ( .C1(n18658), .C2(n18505), .A(n18504), .B(n18503), .ZN(
        P3_U2955) );
  NOR2_X1 U21596 ( .A1(n18684), .A2(n18506), .ZN(n18557) );
  NAND2_X1 U21597 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18557), .ZN(
        n18554) );
  INV_X1 U21598 ( .A(n18507), .ZN(n18548) );
  AND2_X1 U21599 ( .A1(n18727), .A2(n18557), .ZN(n18524) );
  AOI22_X1 U21600 ( .A1(n18604), .A2(n18548), .B1(n18603), .B2(n18524), .ZN(
        n18510) );
  AOI22_X1 U21601 ( .A1(n18608), .A2(n18508), .B1(n18605), .B2(n18557), .ZN(
        n18525) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18525), .B1(
        n18609), .B2(n18523), .ZN(n18509) );
  OAI211_X1 U21603 ( .C1(n18612), .C2(n18554), .A(n18510), .B(n18509), .ZN(
        P3_U2956) );
  AOI22_X1 U21604 ( .A1(n18615), .A2(n18523), .B1(n18613), .B2(n18524), .ZN(
        n18512) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18525), .B1(
        n18614), .B2(n18548), .ZN(n18511) );
  OAI211_X1 U21606 ( .C1(n18618), .C2(n18554), .A(n18512), .B(n18511), .ZN(
        P3_U2957) );
  AOI22_X1 U21607 ( .A1(n18621), .A2(n18523), .B1(n18619), .B2(n18524), .ZN(
        n18514) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18525), .B1(
        n18620), .B2(n18548), .ZN(n18513) );
  OAI211_X1 U21609 ( .C1(n18624), .C2(n18554), .A(n18514), .B(n18513), .ZN(
        P3_U2958) );
  AOI22_X1 U21610 ( .A1(n18626), .A2(n18524), .B1(n18625), .B2(n18523), .ZN(
        n18516) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18525), .B1(
        n18627), .B2(n18548), .ZN(n18515) );
  OAI211_X1 U21612 ( .C1(n18630), .C2(n18554), .A(n18516), .B(n18515), .ZN(
        P3_U2959) );
  AOI22_X1 U21613 ( .A1(n18632), .A2(n18523), .B1(n18631), .B2(n18524), .ZN(
        n18518) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18525), .B1(
        n18633), .B2(n18548), .ZN(n18517) );
  OAI211_X1 U21615 ( .C1(n18636), .C2(n18554), .A(n18518), .B(n18517), .ZN(
        P3_U2960) );
  AOI22_X1 U21616 ( .A1(n18639), .A2(n18548), .B1(n18637), .B2(n18524), .ZN(
        n18520) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18525), .B1(
        n18638), .B2(n18523), .ZN(n18519) );
  OAI211_X1 U21618 ( .C1(n18642), .C2(n18554), .A(n18520), .B(n18519), .ZN(
        P3_U2961) );
  AOI22_X1 U21619 ( .A1(n18644), .A2(n18523), .B1(n18643), .B2(n18524), .ZN(
        n18522) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18525), .B1(
        n18645), .B2(n18548), .ZN(n18521) );
  OAI211_X1 U21621 ( .C1(n18648), .C2(n18554), .A(n18522), .B(n18521), .ZN(
        P3_U2962) );
  AOI22_X1 U21622 ( .A1(n18652), .A2(n18524), .B1(n18650), .B2(n18523), .ZN(
        n18527) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18525), .B1(
        n18653), .B2(n18548), .ZN(n18526) );
  OAI211_X1 U21624 ( .C1(n18658), .C2(n18554), .A(n18527), .B(n18526), .ZN(
        P3_U2963) );
  INV_X1 U21625 ( .A(n18607), .ZN(n18555) );
  NOR2_X2 U21626 ( .A1(n18555), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18649) );
  INV_X1 U21627 ( .A(n18649), .ZN(n18553) );
  NAND2_X1 U21628 ( .A1(n18581), .A2(n18528), .ZN(n18529) );
  NAND2_X1 U21629 ( .A1(n18554), .A2(n18553), .ZN(n18580) );
  INV_X1 U21630 ( .A(n18580), .ZN(n18533) );
  OAI21_X1 U21631 ( .B1(n18530), .B2(n18529), .A(n18533), .ZN(n18531) );
  OAI211_X1 U21632 ( .C1(n18649), .C2(n18832), .A(n18532), .B(n18531), .ZN(
        n18550) );
  NOR2_X1 U21633 ( .A1(n18556), .A2(n18533), .ZN(n18549) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18550), .B1(
        n18603), .B2(n18549), .ZN(n18535) );
  AOI22_X1 U21635 ( .A1(n18604), .A2(n18573), .B1(n18609), .B2(n18548), .ZN(
        n18534) );
  OAI211_X1 U21636 ( .C1(n18612), .C2(n18553), .A(n18535), .B(n18534), .ZN(
        P3_U2964) );
  AOI22_X1 U21637 ( .A1(n18615), .A2(n18548), .B1(n18613), .B2(n18549), .ZN(
        n18537) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18550), .B1(
        n18614), .B2(n18573), .ZN(n18536) );
  OAI211_X1 U21639 ( .C1(n18618), .C2(n18553), .A(n18537), .B(n18536), .ZN(
        P3_U2965) );
  AOI22_X1 U21640 ( .A1(n18621), .A2(n18548), .B1(n18619), .B2(n18549), .ZN(
        n18539) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18550), .B1(
        n18620), .B2(n18573), .ZN(n18538) );
  OAI211_X1 U21642 ( .C1(n18624), .C2(n18553), .A(n18539), .B(n18538), .ZN(
        P3_U2966) );
  AOI22_X1 U21643 ( .A1(n18626), .A2(n18549), .B1(n18625), .B2(n18548), .ZN(
        n18541) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18550), .B1(
        n18627), .B2(n18573), .ZN(n18540) );
  OAI211_X1 U21645 ( .C1(n18630), .C2(n18553), .A(n18541), .B(n18540), .ZN(
        P3_U2967) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18550), .B1(
        n18631), .B2(n18549), .ZN(n18543) );
  AOI22_X1 U21647 ( .A1(n18633), .A2(n18573), .B1(n18632), .B2(n18548), .ZN(
        n18542) );
  OAI211_X1 U21648 ( .C1(n18636), .C2(n18553), .A(n18543), .B(n18542), .ZN(
        P3_U2968) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18550), .B1(
        n18637), .B2(n18549), .ZN(n18545) );
  AOI22_X1 U21650 ( .A1(n18638), .A2(n18548), .B1(n18639), .B2(n18573), .ZN(
        n18544) );
  OAI211_X1 U21651 ( .C1(n18642), .C2(n18553), .A(n18545), .B(n18544), .ZN(
        P3_U2969) );
  AOI22_X1 U21652 ( .A1(n18644), .A2(n18548), .B1(n18643), .B2(n18549), .ZN(
        n18547) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18550), .B1(
        n18645), .B2(n18573), .ZN(n18546) );
  OAI211_X1 U21654 ( .C1(n18648), .C2(n18553), .A(n18547), .B(n18546), .ZN(
        P3_U2970) );
  AOI22_X1 U21655 ( .A1(n18652), .A2(n18549), .B1(n18650), .B2(n18548), .ZN(
        n18552) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18550), .B1(
        n18653), .B2(n18573), .ZN(n18551) );
  OAI211_X1 U21657 ( .C1(n18658), .C2(n18553), .A(n18552), .B(n18551), .ZN(
        P3_U2971) );
  INV_X1 U21658 ( .A(n18554), .ZN(n18597) );
  NOR2_X1 U21659 ( .A1(n18556), .A2(n18555), .ZN(n18572) );
  AOI22_X1 U21660 ( .A1(n18604), .A2(n18597), .B1(n18603), .B2(n18572), .ZN(
        n18559) );
  AOI22_X1 U21661 ( .A1(n18608), .A2(n18557), .B1(n18607), .B2(n18605), .ZN(
        n18574) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18574), .B1(
        n18609), .B2(n18573), .ZN(n18558) );
  OAI211_X1 U21663 ( .C1(n18612), .C2(n18577), .A(n18559), .B(n18558), .ZN(
        P3_U2972) );
  AOI22_X1 U21664 ( .A1(n18615), .A2(n18573), .B1(n18613), .B2(n18572), .ZN(
        n18561) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18574), .B1(
        n18614), .B2(n18597), .ZN(n18560) );
  OAI211_X1 U21666 ( .C1(n18577), .C2(n18618), .A(n18561), .B(n18560), .ZN(
        P3_U2973) );
  AOI22_X1 U21667 ( .A1(n18621), .A2(n18573), .B1(n18619), .B2(n18572), .ZN(
        n18563) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18574), .B1(
        n18620), .B2(n18597), .ZN(n18562) );
  OAI211_X1 U21669 ( .C1(n18577), .C2(n18624), .A(n18563), .B(n18562), .ZN(
        P3_U2974) );
  AOI22_X1 U21670 ( .A1(n18626), .A2(n18572), .B1(n18625), .B2(n18573), .ZN(
        n18565) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18574), .B1(
        n18627), .B2(n18597), .ZN(n18564) );
  OAI211_X1 U21672 ( .C1(n18577), .C2(n18630), .A(n18565), .B(n18564), .ZN(
        P3_U2975) );
  AOI22_X1 U21673 ( .A1(n18632), .A2(n18573), .B1(n18631), .B2(n18572), .ZN(
        n18567) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18574), .B1(
        n18633), .B2(n18597), .ZN(n18566) );
  OAI211_X1 U21675 ( .C1(n18577), .C2(n18636), .A(n18567), .B(n18566), .ZN(
        P3_U2976) );
  AOI22_X1 U21676 ( .A1(n18638), .A2(n18573), .B1(n18637), .B2(n18572), .ZN(
        n18569) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18574), .B1(
        n18639), .B2(n18597), .ZN(n18568) );
  OAI211_X1 U21678 ( .C1(n18577), .C2(n18642), .A(n18569), .B(n18568), .ZN(
        P3_U2977) );
  AOI22_X1 U21679 ( .A1(n18644), .A2(n18573), .B1(n18643), .B2(n18572), .ZN(
        n18571) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18574), .B1(
        n18645), .B2(n18597), .ZN(n18570) );
  OAI211_X1 U21681 ( .C1(n18577), .C2(n18648), .A(n18571), .B(n18570), .ZN(
        P3_U2978) );
  AOI22_X1 U21682 ( .A1(n18653), .A2(n18597), .B1(n18652), .B2(n18572), .ZN(
        n18576) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18574), .B1(
        n18650), .B2(n18573), .ZN(n18575) );
  OAI211_X1 U21684 ( .C1(n18577), .C2(n18658), .A(n18576), .B(n18575), .ZN(
        P3_U2979) );
  INV_X1 U21685 ( .A(n18578), .ZN(n18602) );
  AND2_X1 U21686 ( .A1(n18727), .A2(n18582), .ZN(n18598) );
  AOI22_X1 U21687 ( .A1(n18609), .A2(n18597), .B1(n18603), .B2(n18598), .ZN(
        n18584) );
  OAI221_X1 U21688 ( .B1(n18582), .B2(n18581), .C1(n18582), .C2(n18580), .A(
        n18579), .ZN(n18599) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18599), .B1(
        n18604), .B2(n18649), .ZN(n18583) );
  OAI211_X1 U21690 ( .C1(n18602), .C2(n18612), .A(n18584), .B(n18583), .ZN(
        P3_U2980) );
  AOI22_X1 U21691 ( .A1(n18615), .A2(n18597), .B1(n18613), .B2(n18598), .ZN(
        n18586) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18599), .B1(
        n18614), .B2(n18649), .ZN(n18585) );
  OAI211_X1 U21693 ( .C1(n18602), .C2(n18618), .A(n18586), .B(n18585), .ZN(
        P3_U2981) );
  AOI22_X1 U21694 ( .A1(n18621), .A2(n18597), .B1(n18619), .B2(n18598), .ZN(
        n18588) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18599), .B1(
        n18620), .B2(n18649), .ZN(n18587) );
  OAI211_X1 U21696 ( .C1(n18602), .C2(n18624), .A(n18588), .B(n18587), .ZN(
        P3_U2982) );
  AOI22_X1 U21697 ( .A1(n18626), .A2(n18598), .B1(n18625), .B2(n18597), .ZN(
        n18590) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18599), .B1(
        n18627), .B2(n18649), .ZN(n18589) );
  OAI211_X1 U21699 ( .C1(n18602), .C2(n18630), .A(n18590), .B(n18589), .ZN(
        P3_U2983) );
  AOI22_X1 U21700 ( .A1(n18633), .A2(n18649), .B1(n18631), .B2(n18598), .ZN(
        n18592) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18599), .B1(
        n18632), .B2(n18597), .ZN(n18591) );
  OAI211_X1 U21702 ( .C1(n18602), .C2(n18636), .A(n18592), .B(n18591), .ZN(
        P3_U2984) );
  AOI22_X1 U21703 ( .A1(n18638), .A2(n18597), .B1(n18637), .B2(n18598), .ZN(
        n18594) );
  AOI22_X1 U21704 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18599), .B1(
        n18639), .B2(n18649), .ZN(n18593) );
  OAI211_X1 U21705 ( .C1(n18602), .C2(n18642), .A(n18594), .B(n18593), .ZN(
        P3_U2985) );
  AOI22_X1 U21706 ( .A1(n18645), .A2(n18649), .B1(n18643), .B2(n18598), .ZN(
        n18596) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18599), .B1(
        n18644), .B2(n18597), .ZN(n18595) );
  OAI211_X1 U21708 ( .C1(n18602), .C2(n18648), .A(n18596), .B(n18595), .ZN(
        P3_U2986) );
  AOI22_X1 U21709 ( .A1(n18652), .A2(n18598), .B1(n18650), .B2(n18597), .ZN(
        n18601) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18599), .B1(
        n18653), .B2(n18649), .ZN(n18600) );
  OAI211_X1 U21711 ( .C1(n18602), .C2(n18658), .A(n18601), .B(n18600), .ZN(
        P3_U2987) );
  AND2_X1 U21712 ( .A1(n18727), .A2(n18606), .ZN(n18651) );
  AOI22_X1 U21713 ( .A1(n18604), .A2(n18654), .B1(n18603), .B2(n18651), .ZN(
        n18611) );
  AOI22_X1 U21714 ( .A1(n18608), .A2(n18607), .B1(n18606), .B2(n18605), .ZN(
        n18655) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18655), .B1(
        n18609), .B2(n18649), .ZN(n18610) );
  OAI211_X1 U21716 ( .C1(n18659), .C2(n18612), .A(n18611), .B(n18610), .ZN(
        P3_U2988) );
  AOI22_X1 U21717 ( .A1(n18654), .A2(n18614), .B1(n18613), .B2(n18651), .ZN(
        n18617) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18655), .B1(
        n18615), .B2(n18649), .ZN(n18616) );
  OAI211_X1 U21719 ( .C1(n18659), .C2(n18618), .A(n18617), .B(n18616), .ZN(
        P3_U2989) );
  AOI22_X1 U21720 ( .A1(n18654), .A2(n18620), .B1(n18619), .B2(n18651), .ZN(
        n18623) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18655), .B1(
        n18621), .B2(n18649), .ZN(n18622) );
  OAI211_X1 U21722 ( .C1(n18659), .C2(n18624), .A(n18623), .B(n18622), .ZN(
        P3_U2990) );
  AOI22_X1 U21723 ( .A1(n18626), .A2(n18651), .B1(n18625), .B2(n18649), .ZN(
        n18629) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18627), .ZN(n18628) );
  OAI211_X1 U21725 ( .C1(n18659), .C2(n18630), .A(n18629), .B(n18628), .ZN(
        P3_U2991) );
  AOI22_X1 U21726 ( .A1(n18632), .A2(n18649), .B1(n18631), .B2(n18651), .ZN(
        n18635) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18633), .ZN(n18634) );
  OAI211_X1 U21728 ( .C1(n18659), .C2(n18636), .A(n18635), .B(n18634), .ZN(
        P3_U2992) );
  AOI22_X1 U21729 ( .A1(n18638), .A2(n18649), .B1(n18637), .B2(n18651), .ZN(
        n18641) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18639), .ZN(n18640) );
  OAI211_X1 U21731 ( .C1(n18659), .C2(n18642), .A(n18641), .B(n18640), .ZN(
        P3_U2993) );
  AOI22_X1 U21732 ( .A1(n18644), .A2(n18649), .B1(n18643), .B2(n18651), .ZN(
        n18647) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18645), .ZN(n18646) );
  OAI211_X1 U21734 ( .C1(n18659), .C2(n18648), .A(n18647), .B(n18646), .ZN(
        P3_U2994) );
  AOI22_X1 U21735 ( .A1(n18652), .A2(n18651), .B1(n18650), .B2(n18649), .ZN(
        n18657) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18653), .ZN(n18656) );
  OAI211_X1 U21737 ( .C1(n18659), .C2(n18658), .A(n18657), .B(n18656), .ZN(
        P3_U2995) );
  OAI22_X1 U21738 ( .A1(n18663), .A2(n18662), .B1(n18661), .B2(n18660), .ZN(
        n18664) );
  AOI221_X1 U21739 ( .B1(n18667), .B2(n18666), .C1(n18665), .C2(n18666), .A(
        n18664), .ZN(n18875) );
  AOI211_X1 U21740 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18703), .A(
        n18669), .B(n18668), .ZN(n18714) );
  INV_X1 U21741 ( .A(n18703), .ZN(n18702) );
  AOI22_X1 U21742 ( .A1(n18849), .A2(n18670), .B1(n18697), .B2(n18682), .ZN(
        n18671) );
  OAI21_X1 U21743 ( .B1(n18672), .B2(n18690), .A(n18671), .ZN(n18838) );
  NOR2_X1 U21744 ( .A1(n18839), .A2(n18838), .ZN(n18677) );
  NOR2_X1 U21745 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18689), .ZN(
        n18675) );
  NAND2_X1 U21746 ( .A1(n18673), .A2(n16933), .ZN(n18680) );
  INV_X1 U21747 ( .A(n18680), .ZN(n18674) );
  OAI22_X1 U21748 ( .A1(n18675), .A2(n18701), .B1(n18674), .B2(n18697), .ZN(
        n18835) );
  AOI21_X1 U21749 ( .B1(n18835), .B2(n18702), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18676) );
  AOI21_X1 U21750 ( .B1(n18702), .B2(n18677), .A(n18676), .ZN(n18710) );
  NAND2_X1 U21751 ( .A1(n18679), .A2(n18678), .ZN(n18681) );
  AOI22_X1 U21752 ( .A1(n18853), .A2(n18681), .B1(n12687), .B2(n18680), .ZN(
        n18850) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18682), .B1(
        n18681), .B2(n16933), .ZN(n18685) );
  INV_X1 U21754 ( .A(n18685), .ZN(n18857) );
  NOR3_X1 U21755 ( .A1(n18684), .A2(n18683), .A3(n18857), .ZN(n18686) );
  OAI22_X1 U21756 ( .A1(n18850), .A2(n18686), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18685), .ZN(n18688) );
  AOI21_X1 U21757 ( .B1(n18688), .B2(n18702), .A(n18687), .ZN(n18705) );
  NOR2_X1 U21758 ( .A1(n18689), .A2(n18849), .ZN(n18696) );
  OAI21_X1 U21759 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18693), .A(
        n18690), .ZN(n18695) );
  NAND2_X1 U21760 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18691), .ZN(
        n18692) );
  AOI211_X1 U21761 ( .C1(n18693), .C2(n18692), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n12687), .ZN(n18694) );
  AOI21_X1 U21762 ( .B1(n18696), .B2(n18695), .A(n18694), .ZN(n18700) );
  OAI211_X1 U21763 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18698), .B(n18697), .ZN(
        n18699) );
  OAI211_X1 U21764 ( .C1(n18845), .C2(n18701), .A(n18700), .B(n18699), .ZN(
        n18847) );
  AOI22_X1 U21765 ( .A1(n18703), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18847), .B2(n18702), .ZN(n18706) );
  OR2_X1 U21766 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18706), .ZN(
        n18704) );
  AOI221_X1 U21767 ( .B1(n18705), .B2(n18704), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18706), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18709) );
  OAI21_X1 U21768 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18706), .ZN(n18708) );
  AOI222_X1 U21769 ( .A1(n18710), .A2(n18709), .B1(n18710), .B2(n18708), .C1(
        n18709), .C2(n18707), .ZN(n18713) );
  OAI21_X1 U21770 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18711), .ZN(n18712) );
  NAND4_X1 U21771 ( .A1(n18875), .A2(n18714), .A3(n18713), .A4(n18712), .ZN(
        n18724) );
  AOI211_X1 U21772 ( .C1(n18717), .C2(n18716), .A(n18715), .B(n18724), .ZN(
        n18830) );
  AOI21_X1 U21773 ( .B1(n18880), .B2(n18718), .A(n18830), .ZN(n18728) );
  NOR2_X1 U21774 ( .A1(n18719), .A2(n18727), .ZN(n18723) );
  NAND2_X1 U21775 ( .A1(n18880), .A2(n18720), .ZN(n18732) );
  INV_X1 U21776 ( .A(n18732), .ZN(n18721) );
  AOI211_X1 U21777 ( .C1(n18856), .C2(n18888), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18721), .ZN(n18722) );
  AOI211_X1 U21778 ( .C1(n18878), .C2(n18724), .A(n18723), .B(n18722), .ZN(
        n18725) );
  OAI221_X1 U21779 ( .B1(n18829), .B2(n18728), .C1(n18829), .C2(n18726), .A(
        n18725), .ZN(P3_U2996) );
  NOR4_X1 U21780 ( .A1(n18829), .A2(n18842), .A3(n18886), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18735) );
  INV_X1 U21781 ( .A(n18735), .ZN(n18731) );
  NAND3_X1 U21782 ( .A1(n18729), .A2(n18728), .A3(n18727), .ZN(n18730) );
  NAND4_X1 U21783 ( .A1(n18733), .A2(n18732), .A3(n18731), .A4(n18730), .ZN(
        P3_U2997) );
  OAI21_X1 U21784 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18734), .ZN(n18736) );
  AOI21_X1 U21785 ( .B1(n18737), .B2(n18736), .A(n18735), .ZN(P3_U2998) );
  AND2_X1 U21786 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18738), .ZN(
        P3_U2999) );
  AND2_X1 U21787 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18738), .ZN(
        P3_U3000) );
  AND2_X1 U21788 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18738), .ZN(
        P3_U3001) );
  AND2_X1 U21789 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18738), .ZN(
        P3_U3002) );
  AND2_X1 U21790 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18738), .ZN(
        P3_U3003) );
  AND2_X1 U21791 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18738), .ZN(
        P3_U3004) );
  AND2_X1 U21792 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18738), .ZN(
        P3_U3005) );
  AND2_X1 U21793 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18738), .ZN(
        P3_U3006) );
  AND2_X1 U21794 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18738), .ZN(
        P3_U3007) );
  AND2_X1 U21795 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18738), .ZN(
        P3_U3008) );
  AND2_X1 U21796 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18738), .ZN(
        P3_U3009) );
  AND2_X1 U21797 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18738), .ZN(
        P3_U3010) );
  AND2_X1 U21798 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18738), .ZN(
        P3_U3011) );
  AND2_X1 U21799 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18738), .ZN(
        P3_U3012) );
  AND2_X1 U21800 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18738), .ZN(
        P3_U3013) );
  AND2_X1 U21801 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18738), .ZN(
        P3_U3014) );
  AND2_X1 U21802 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18738), .ZN(
        P3_U3015) );
  AND2_X1 U21803 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18738), .ZN(
        P3_U3016) );
  AND2_X1 U21804 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18738), .ZN(
        P3_U3017) );
  AND2_X1 U21805 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18738), .ZN(
        P3_U3018) );
  AND2_X1 U21806 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18738), .ZN(
        P3_U3019) );
  AND2_X1 U21807 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18738), .ZN(
        P3_U3020) );
  AND2_X1 U21808 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18738), .ZN(P3_U3021) );
  AND2_X1 U21809 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18825), .ZN(P3_U3022) );
  AND2_X1 U21810 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18825), .ZN(P3_U3023) );
  AND2_X1 U21811 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18825), .ZN(P3_U3024) );
  AND2_X1 U21812 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18825), .ZN(P3_U3025) );
  AND2_X1 U21813 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18825), .ZN(P3_U3026) );
  AND2_X1 U21814 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18825), .ZN(P3_U3027) );
  AND2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18825), .ZN(P3_U3028) );
  NOR2_X1 U21816 ( .A1(n18886), .A2(n18739), .ZN(n18746) );
  INV_X1 U21817 ( .A(n18746), .ZN(n18748) );
  OAI21_X1 U21818 ( .B1(n18740), .B2(n20988), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18742) );
  INV_X1 U21819 ( .A(NA), .ZN(n21052) );
  NOR3_X1 U21820 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .A3(n21052), .ZN(n18741) );
  AOI21_X1 U21821 ( .B1(n18894), .B2(n18742), .A(n18741), .ZN(n18743) );
  OAI221_X1 U21822 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(P3_STATE_REG_0__SCAN_IN), .C1(P3_STATE_REG_2__SCAN_IN), .C2(n18748), .A(n18743), .ZN(P3_U3029) );
  NAND2_X1 U21823 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n18747) );
  AOI22_X1 U21824 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18747), .B1(HOLD), 
        .B2(n18744), .ZN(n18745) );
  OAI211_X1 U21825 ( .C1(n18745), .C2(n18752), .A(n18748), .B(n18883), .ZN(
        P3_U3030) );
  AOI221_X1 U21826 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18752), .C1(n21052), 
        .C2(n18752), .A(n18746), .ZN(n18753) );
  INV_X1 U21827 ( .A(n18747), .ZN(n18750) );
  OAI22_X1 U21828 ( .A1(NA), .A2(n18748), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18749) );
  OAI22_X1 U21829 ( .A1(n18750), .A2(n18749), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18751) );
  OAI22_X1 U21830 ( .A1(n18753), .A2(n18754), .B1(n18752), .B2(n18751), .ZN(
        P3_U3031) );
  INV_X1 U21831 ( .A(n18894), .ZN(n18893) );
  INV_X1 U21832 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18757) );
  OAI222_X1 U21833 ( .A1(n18863), .A2(n9805), .B1(n18755), .B2(n18893), .C1(
        n18757), .C2(n18805), .ZN(P3_U3032) );
  OAI222_X1 U21834 ( .A1(n18805), .A2(n18760), .B1(n18758), .B2(n18815), .C1(
        n18757), .C2(n9805), .ZN(P3_U3033) );
  OAI222_X1 U21835 ( .A1(n18760), .A2(n9805), .B1(n18759), .B2(n18893), .C1(
        n18761), .C2(n18805), .ZN(P3_U3034) );
  OAI222_X1 U21836 ( .A1(n18805), .A2(n18763), .B1(n18762), .B2(n18815), .C1(
        n18761), .C2(n9805), .ZN(P3_U3035) );
  OAI222_X1 U21837 ( .A1(n18805), .A2(n18765), .B1(n18764), .B2(n18893), .C1(
        n18763), .C2(n9805), .ZN(P3_U3036) );
  OAI222_X1 U21838 ( .A1(n18805), .A2(n18767), .B1(n18766), .B2(n18893), .C1(
        n18765), .C2(n9805), .ZN(P3_U3037) );
  INV_X1 U21839 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18770) );
  OAI222_X1 U21840 ( .A1(n18805), .A2(n18770), .B1(n18768), .B2(n18821), .C1(
        n18767), .C2(n9805), .ZN(P3_U3038) );
  OAI222_X1 U21841 ( .A1(n18770), .A2(n9805), .B1(n18769), .B2(n18893), .C1(
        n18771), .C2(n18805), .ZN(P3_U3039) );
  OAI222_X1 U21842 ( .A1(n18805), .A2(n18773), .B1(n18772), .B2(n18893), .C1(
        n18771), .C2(n9805), .ZN(P3_U3040) );
  OAI222_X1 U21843 ( .A1(n18805), .A2(n18775), .B1(n18774), .B2(n18893), .C1(
        n18773), .C2(n9805), .ZN(P3_U3041) );
  INV_X1 U21844 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18777) );
  OAI222_X1 U21845 ( .A1(n18805), .A2(n18777), .B1(n18776), .B2(n18893), .C1(
        n18775), .C2(n9805), .ZN(P3_U3042) );
  OAI222_X1 U21846 ( .A1(n18805), .A2(n18779), .B1(n18778), .B2(n18893), .C1(
        n18777), .C2(n9805), .ZN(P3_U3043) );
  OAI222_X1 U21847 ( .A1(n18805), .A2(n18782), .B1(n18780), .B2(n18893), .C1(
        n18779), .C2(n9805), .ZN(P3_U3044) );
  OAI222_X1 U21848 ( .A1(n18782), .A2(n9805), .B1(n18781), .B2(n18893), .C1(
        n18783), .C2(n18805), .ZN(P3_U3045) );
  OAI222_X1 U21849 ( .A1(n18805), .A2(n18785), .B1(n18784), .B2(n18893), .C1(
        n18783), .C2(n9805), .ZN(P3_U3046) );
  OAI222_X1 U21850 ( .A1(n18805), .A2(n18788), .B1(n18786), .B2(n18893), .C1(
        n18785), .C2(n9805), .ZN(P3_U3047) );
  OAI222_X1 U21851 ( .A1(n18788), .A2(n9805), .B1(n18787), .B2(n18893), .C1(
        n18789), .C2(n18805), .ZN(P3_U3048) );
  OAI222_X1 U21852 ( .A1(n18805), .A2(n18791), .B1(n18790), .B2(n18893), .C1(
        n18789), .C2(n9805), .ZN(P3_U3049) );
  OAI222_X1 U21853 ( .A1(n18805), .A2(n18794), .B1(n18792), .B2(n18893), .C1(
        n18791), .C2(n9805), .ZN(P3_U3050) );
  OAI222_X1 U21854 ( .A1(n18794), .A2(n9805), .B1(n18793), .B2(n18893), .C1(
        n18795), .C2(n18805), .ZN(P3_U3051) );
  OAI222_X1 U21855 ( .A1(n18805), .A2(n18797), .B1(n18796), .B2(n18893), .C1(
        n18795), .C2(n9805), .ZN(P3_U3052) );
  INV_X1 U21856 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18800) );
  OAI222_X1 U21857 ( .A1(n18805), .A2(n18800), .B1(n18798), .B2(n18893), .C1(
        n18797), .C2(n9805), .ZN(P3_U3053) );
  OAI222_X1 U21858 ( .A1(n18800), .A2(n9805), .B1(n18799), .B2(n18815), .C1(
        n18801), .C2(n18805), .ZN(P3_U3054) );
  OAI222_X1 U21859 ( .A1(n18805), .A2(n18803), .B1(n18802), .B2(n18815), .C1(
        n18801), .C2(n9805), .ZN(P3_U3055) );
  OAI222_X1 U21860 ( .A1(n18805), .A2(n18806), .B1(n18804), .B2(n18815), .C1(
        n18803), .C2(n9805), .ZN(P3_U3056) );
  OAI222_X1 U21861 ( .A1(n18805), .A2(n18808), .B1(n18807), .B2(n18815), .C1(
        n18806), .C2(n9805), .ZN(P3_U3057) );
  OAI222_X1 U21862 ( .A1(n18805), .A2(n18811), .B1(n18809), .B2(n18815), .C1(
        n18808), .C2(n9805), .ZN(P3_U3058) );
  OAI222_X1 U21863 ( .A1(n18811), .A2(n9805), .B1(n18810), .B2(n18815), .C1(
        n18812), .C2(n18805), .ZN(P3_U3059) );
  OAI222_X1 U21864 ( .A1(n18805), .A2(n18817), .B1(n18813), .B2(n18815), .C1(
        n18812), .C2(n9805), .ZN(P3_U3060) );
  INV_X1 U21865 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18816) );
  OAI222_X1 U21866 ( .A1(n9805), .A2(n18817), .B1(n18816), .B2(n18815), .C1(
        n18814), .C2(n18805), .ZN(P3_U3061) );
  OAI22_X1 U21867 ( .A1(n18894), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18893), .ZN(n18818) );
  INV_X1 U21868 ( .A(n18818), .ZN(P3_U3274) );
  OAI22_X1 U21869 ( .A1(n18894), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18893), .ZN(n18819) );
  INV_X1 U21870 ( .A(n18819), .ZN(P3_U3275) );
  OAI22_X1 U21871 ( .A1(n18894), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18893), .ZN(n18820) );
  INV_X1 U21872 ( .A(n18820), .ZN(P3_U3276) );
  OAI22_X1 U21873 ( .A1(n18894), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18821), .ZN(n18822) );
  INV_X1 U21874 ( .A(n18822), .ZN(P3_U3277) );
  INV_X1 U21875 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18824) );
  INV_X1 U21876 ( .A(n18826), .ZN(n18823) );
  AOI21_X1 U21877 ( .B1(n18825), .B2(n18824), .A(n18823), .ZN(P3_U3280) );
  OAI21_X1 U21878 ( .B1(n18828), .B2(n18827), .A(n18826), .ZN(P3_U3281) );
  NOR2_X1 U21879 ( .A1(n18830), .A2(n18829), .ZN(n18833) );
  OAI21_X1 U21880 ( .B1(n18833), .B2(n18832), .A(n18831), .ZN(P3_U3282) );
  INV_X1 U21881 ( .A(n18834), .ZN(n18837) );
  NOR2_X1 U21882 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18896), .ZN(
        n18836) );
  AOI22_X1 U21883 ( .A1(n18856), .A2(n18837), .B1(n18836), .B2(n18835), .ZN(
        n18841) );
  AOI21_X1 U21884 ( .B1(n18858), .B2(n18838), .A(n18862), .ZN(n18840) );
  OAI22_X1 U21885 ( .A1(n18862), .A2(n18841), .B1(n18840), .B2(n18839), .ZN(
        P3_U3285) );
  NOR2_X1 U21886 ( .A1(n18842), .A2(n18859), .ZN(n18851) );
  OAI22_X1 U21887 ( .A1(n18844), .A2(n18843), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18852) );
  INV_X1 U21888 ( .A(n18852), .ZN(n18846) );
  AOI222_X1 U21889 ( .A1(n18847), .A2(n18858), .B1(n18851), .B2(n18846), .C1(
        n18856), .C2(n18845), .ZN(n18848) );
  AOI22_X1 U21890 ( .A1(n18862), .A2(n18849), .B1(n18848), .B2(n18860), .ZN(
        P3_U3288) );
  INV_X1 U21891 ( .A(n18850), .ZN(n18854) );
  AOI222_X1 U21892 ( .A1(n18854), .A2(n18858), .B1(n18856), .B2(n18853), .C1(
        n18852), .C2(n18851), .ZN(n18855) );
  AOI22_X1 U21893 ( .A1(n18862), .A2(n12687), .B1(n18855), .B2(n18860), .ZN(
        P3_U3289) );
  AOI222_X1 U21894 ( .A1(n18859), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18858), 
        .B2(n18857), .C1(n16933), .C2(n18856), .ZN(n18861) );
  AOI22_X1 U21895 ( .A1(n18862), .A2(n16933), .B1(n18861), .B2(n18860), .ZN(
        P3_U3290) );
  AOI21_X1 U21896 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18864) );
  AOI22_X1 U21897 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18864), .B2(n18863), .ZN(n18866) );
  INV_X1 U21898 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18865) );
  AOI22_X1 U21899 ( .A1(n18867), .A2(n18866), .B1(n18865), .B2(n18870), .ZN(
        P3_U3292) );
  INV_X1 U21900 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18871) );
  NOR2_X1 U21901 ( .A1(n18870), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18868) );
  AOI22_X1 U21902 ( .A1(n18871), .A2(n18870), .B1(n18869), .B2(n18868), .ZN(
        P3_U3293) );
  INV_X1 U21903 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18872) );
  AOI22_X1 U21904 ( .A1(n18893), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18872), 
        .B2(n18894), .ZN(P3_U3294) );
  INV_X1 U21905 ( .A(n18873), .ZN(n18876) );
  NAND2_X1 U21906 ( .A1(n18876), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18874) );
  OAI21_X1 U21907 ( .B1(n18876), .B2(n18875), .A(n18874), .ZN(P3_U3295) );
  OAI22_X1 U21908 ( .A1(n18880), .A2(n18879), .B1(n18878), .B2(n18877), .ZN(
        n18881) );
  NOR2_X1 U21909 ( .A1(n18882), .A2(n18881), .ZN(n18892) );
  AOI21_X1 U21910 ( .B1(n18885), .B2(n18884), .A(n18883), .ZN(n18887) );
  OAI211_X1 U21911 ( .C1(n18897), .C2(n18887), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18886), .ZN(n18889) );
  AOI21_X1 U21912 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18889), .A(n18888), 
        .ZN(n18891) );
  NAND2_X1 U21913 ( .A1(n18892), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18890) );
  OAI21_X1 U21914 ( .B1(n18892), .B2(n18891), .A(n18890), .ZN(P3_U3296) );
  OAI22_X1 U21915 ( .A1(n18894), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18893), .ZN(n18895) );
  INV_X1 U21916 ( .A(n18895), .ZN(P3_U3297) );
  OAI21_X1 U21917 ( .B1(n18896), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18898), 
        .ZN(n18901) );
  OAI22_X1 U21918 ( .A1(n18901), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18898), 
        .B2(n18897), .ZN(n18899) );
  INV_X1 U21919 ( .A(n18899), .ZN(P3_U3298) );
  OAI21_X1 U21920 ( .B1(n18901), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18900), 
        .ZN(n18902) );
  INV_X1 U21921 ( .A(n18902), .ZN(P3_U3299) );
  INV_X1 U21922 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18908) );
  NAND2_X1 U21923 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19877), .ZN(n19867) );
  NAND2_X1 U21924 ( .A1(n18908), .A2(n18903), .ZN(n19864) );
  OAI21_X1 U21925 ( .B1(n18908), .B2(n19867), .A(n19864), .ZN(n19944) );
  AOI21_X1 U21926 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19944), .ZN(n18904) );
  INV_X1 U21927 ( .A(n18904), .ZN(P2_U2815) );
  INV_X1 U21928 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18909) );
  OAI22_X1 U21929 ( .A1(n18907), .A2(n18909), .B1(n18906), .B2(n18905), .ZN(
        P2_U2816) );
  INV_X1 U21930 ( .A(n19858), .ZN(n19872) );
  NAND2_X1 U21931 ( .A1(n18908), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20001) );
  AOI22_X1 U21932 ( .A1(n20000), .A2(n18909), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n20001), .ZN(n18910) );
  OAI21_X1 U21933 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19872), .A(n18910), 
        .ZN(P2_U2817) );
  OAI21_X1 U21934 ( .B1(n19858), .B2(BS16), .A(n19944), .ZN(n19942) );
  OAI21_X1 U21935 ( .B1(n19944), .B2(n19457), .A(n19942), .ZN(P2_U2818) );
  NOR4_X1 U21936 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18914) );
  NOR4_X1 U21937 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18913) );
  NOR4_X1 U21938 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18912) );
  NOR4_X1 U21939 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18911) );
  NAND4_X1 U21940 ( .A1(n18914), .A2(n18913), .A3(n18912), .A4(n18911), .ZN(
        n18920) );
  NOR4_X1 U21941 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18918) );
  AOI211_X1 U21942 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18917) );
  NOR4_X1 U21943 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18916) );
  NOR4_X1 U21944 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18915) );
  NAND4_X1 U21945 ( .A1(n18918), .A2(n18917), .A3(n18916), .A4(n18915), .ZN(
        n18919) );
  NOR2_X1 U21946 ( .A1(n18920), .A2(n18919), .ZN(n18931) );
  INV_X1 U21947 ( .A(n18931), .ZN(n18929) );
  NOR2_X1 U21948 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18929), .ZN(n18923) );
  INV_X1 U21949 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18921) );
  AOI22_X1 U21950 ( .A1(n18923), .A2(n18924), .B1(n18929), .B2(n18921), .ZN(
        P2_U2820) );
  OR3_X1 U21951 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18928) );
  INV_X1 U21952 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18922) );
  AOI22_X1 U21953 ( .A1(n18923), .A2(n18928), .B1(n18929), .B2(n18922), .ZN(
        P2_U2821) );
  INV_X1 U21954 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19943) );
  NAND2_X1 U21955 ( .A1(n18923), .A2(n19943), .ZN(n18927) );
  OAI21_X1 U21956 ( .B1(n19878), .B2(n18924), .A(n18931), .ZN(n18925) );
  OAI21_X1 U21957 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18931), .A(n18925), 
        .ZN(n18926) );
  OAI221_X1 U21958 ( .B1(n18927), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18927), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18926), .ZN(P2_U2822) );
  INV_X1 U21959 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18930) );
  OAI221_X1 U21960 ( .B1(n18931), .B2(n18930), .C1(n18929), .C2(n18928), .A(
        n18927), .ZN(P2_U2823) );
  INV_X1 U21961 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19915) );
  OAI22_X1 U21962 ( .A1(n18932), .A2(n19072), .B1(n19915), .B2(n19049), .ZN(
        n18934) );
  NOR2_X1 U21963 ( .A1(n19087), .A2(n14961), .ZN(n18933) );
  AOI211_X1 U21964 ( .C1(n18935), .C2(n19081), .A(n18934), .B(n18933), .ZN(
        n18936) );
  OAI21_X1 U21965 ( .B1(n18937), .B2(n19105), .A(n18936), .ZN(n18938) );
  INV_X1 U21966 ( .A(n18938), .ZN(n18943) );
  OAI211_X1 U21967 ( .C1(n18941), .C2(n18940), .A(n19094), .B(n18939), .ZN(
        n18942) );
  OAI211_X1 U21968 ( .C1(n19085), .C2(n18944), .A(n18943), .B(n18942), .ZN(
        P2_U2834) );
  AOI22_X1 U21969 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19102), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19114), .ZN(n18955) );
  AOI22_X1 U21970 ( .A1(n18945), .A2(n19039), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19107), .ZN(n18954) );
  INV_X1 U21971 ( .A(n18946), .ZN(n18948) );
  AOI22_X1 U21972 ( .A1(n18948), .A2(n19081), .B1(n18947), .B2(n19101), .ZN(
        n18953) );
  OAI211_X1 U21973 ( .C1(n18951), .C2(n18950), .A(n19094), .B(n18949), .ZN(
        n18952) );
  NAND4_X1 U21974 ( .A1(n18955), .A2(n18954), .A3(n18953), .A4(n18952), .ZN(
        P2_U2835) );
  OAI21_X1 U21975 ( .B1(n19912), .B2(n19049), .A(n19041), .ZN(n18960) );
  INV_X1 U21976 ( .A(n18956), .ZN(n18958) );
  OAI22_X1 U21977 ( .A1(n18958), .A2(n19105), .B1(n19072), .B2(n18957), .ZN(
        n18959) );
  AOI211_X1 U21978 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19107), .A(n18960), .B(
        n18959), .ZN(n18967) );
  NAND2_X1 U21979 ( .A1(n13929), .A2(n18961), .ZN(n18962) );
  XNOR2_X1 U21980 ( .A(n18963), .B(n18962), .ZN(n18965) );
  AOI22_X1 U21981 ( .A1(n18965), .A2(n19094), .B1(n18964), .B2(n19081), .ZN(
        n18966) );
  OAI211_X1 U21982 ( .C1(n18968), .C2(n19085), .A(n18967), .B(n18966), .ZN(
        P2_U2836) );
  INV_X1 U21983 ( .A(n19113), .ZN(n19023) );
  AOI211_X1 U21984 ( .C1(n18971), .C2(n18970), .A(n18969), .B(n19117), .ZN(
        n18977) );
  NAND2_X1 U21985 ( .A1(n18972), .A2(n19039), .ZN(n18975) );
  AOI22_X1 U21986 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19114), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19107), .ZN(n18974) );
  NAND2_X1 U21987 ( .A1(n19102), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n18973) );
  NAND4_X1 U21988 ( .A1(n18975), .A2(n18974), .A3(n19041), .A4(n18973), .ZN(
        n18976) );
  NOR2_X1 U21989 ( .A1(n18977), .A2(n18976), .ZN(n18982) );
  INV_X1 U21990 ( .A(n18978), .ZN(n18979) );
  AOI22_X1 U21991 ( .A1(n18980), .A2(n19081), .B1(n19101), .B2(n18979), .ZN(
        n18981) );
  OAI211_X1 U21992 ( .C1(n18983), .C2(n19023), .A(n18982), .B(n18981), .ZN(
        P2_U2838) );
  INV_X1 U21993 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n18984) );
  OAI22_X1 U21994 ( .A1(n18985), .A2(n19105), .B1(n19087), .B2(n18984), .ZN(
        n18986) );
  AOI211_X1 U21995 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19102), .A(n19235), 
        .B(n18986), .ZN(n18994) );
  OR2_X1 U21996 ( .A1(n19092), .A2(n18987), .ZN(n19004) );
  XOR2_X1 U21997 ( .A(n18988), .B(n19004), .Z(n18992) );
  OAI22_X1 U21998 ( .A1(n19109), .A2(n18990), .B1(n18989), .B2(n19085), .ZN(
        n18991) );
  AOI21_X1 U21999 ( .B1(n18992), .B2(n19094), .A(n18991), .ZN(n18993) );
  OAI211_X1 U22000 ( .C1(n10048), .C2(n19072), .A(n18994), .B(n18993), .ZN(
        P2_U2839) );
  INV_X1 U22001 ( .A(n18995), .ZN(n18998) );
  AOI21_X1 U22002 ( .B1(n19102), .B2(P2_REIP_REG_15__SCAN_IN), .A(n19076), 
        .ZN(n18997) );
  NAND2_X1 U22003 ( .A1(n19005), .A2(n19113), .ZN(n18996) );
  OAI211_X1 U22004 ( .C1(n19109), .C2(n18998), .A(n18997), .B(n18996), .ZN(
        n19002) );
  OAI22_X1 U22005 ( .A1(n19087), .A2(n19000), .B1(n18999), .B2(n19072), .ZN(
        n19001) );
  AOI211_X1 U22006 ( .C1(n19039), .C2(n19003), .A(n19002), .B(n19001), .ZN(
        n19009) );
  AOI211_X1 U22007 ( .C1(n19006), .C2(n19005), .A(n19048), .B(n19004), .ZN(
        n19007) );
  INV_X1 U22008 ( .A(n19007), .ZN(n19008) );
  OAI211_X1 U22009 ( .C1(n19085), .C2(n19125), .A(n19009), .B(n19008), .ZN(
        P2_U2840) );
  AOI211_X1 U22010 ( .C1(n19012), .C2(n19011), .A(n19010), .B(n19117), .ZN(
        n19018) );
  NAND2_X1 U22011 ( .A1(n19013), .A2(n19039), .ZN(n19016) );
  AOI22_X1 U22012 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19114), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19107), .ZN(n19015) );
  NAND2_X1 U22013 ( .A1(n19102), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n19014) );
  NAND4_X1 U22014 ( .A1(n19016), .A2(n19015), .A3(n19041), .A4(n19014), .ZN(
        n19017) );
  NOR2_X1 U22015 ( .A1(n19018), .A2(n19017), .ZN(n19022) );
  INV_X1 U22016 ( .A(n19130), .ZN(n19019) );
  AOI22_X1 U22017 ( .A1(n19020), .A2(n19081), .B1(n19101), .B2(n19019), .ZN(
        n19021) );
  OAI211_X1 U22018 ( .C1(n19024), .C2(n19023), .A(n19022), .B(n19021), .ZN(
        P2_U2842) );
  OAI21_X1 U22019 ( .B1(n10504), .B2(n19049), .A(n19041), .ZN(n19028) );
  OAI22_X1 U22020 ( .A1(n19026), .A2(n19105), .B1(n19087), .B2(n19025), .ZN(
        n19027) );
  AOI211_X1 U22021 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n19114), .A(
        n19028), .B(n19027), .ZN(n19035) );
  NAND2_X1 U22022 ( .A1(n13929), .A2(n19029), .ZN(n19030) );
  XNOR2_X1 U22023 ( .A(n19031), .B(n19030), .ZN(n19033) );
  AOI22_X1 U22024 ( .A1(n19033), .A2(n19094), .B1(n19032), .B2(n19081), .ZN(
        n19034) );
  OAI211_X1 U22025 ( .C1(n19135), .C2(n19085), .A(n19035), .B(n19034), .ZN(
        P2_U2844) );
  NOR2_X1 U22026 ( .A1(n19092), .A2(n19036), .ZN(n19037) );
  XOR2_X1 U22027 ( .A(n19038), .B(n19037), .Z(n19047) );
  AOI22_X1 U22028 ( .A1(n19040), .A2(n19039), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19107), .ZN(n19042) );
  OAI211_X1 U22029 ( .C1(n19895), .C2(n19049), .A(n19042), .B(n19041), .ZN(
        n19045) );
  OAI22_X1 U22030 ( .A1(n19109), .A2(n19043), .B1(n19138), .B2(n19085), .ZN(
        n19044) );
  AOI211_X1 U22031 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19114), .A(
        n19045), .B(n19044), .ZN(n19046) );
  OAI21_X1 U22032 ( .B1(n19048), .B2(n19047), .A(n19046), .ZN(P2_U2845) );
  OAI21_X1 U22033 ( .B1(n19893), .B2(n19049), .A(n19041), .ZN(n19053) );
  INV_X1 U22034 ( .A(n19050), .ZN(n19051) );
  OAI22_X1 U22035 ( .A1(n19051), .A2(n19105), .B1(n19087), .B2(n10887), .ZN(
        n19052) );
  AOI211_X1 U22036 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19114), .A(
        n19053), .B(n19052), .ZN(n19060) );
  NAND2_X1 U22037 ( .A1(n13929), .A2(n19054), .ZN(n19055) );
  XNOR2_X1 U22038 ( .A(n19056), .B(n19055), .ZN(n19058) );
  AOI22_X1 U22039 ( .A1(n19058), .A2(n19094), .B1(n19057), .B2(n19081), .ZN(
        n19059) );
  OAI211_X1 U22040 ( .C1(n19141), .C2(n19085), .A(n19060), .B(n19059), .ZN(
        P2_U2846) );
  OAI22_X1 U22041 ( .A1(n19087), .A2(n19062), .B1(n19061), .B2(n19105), .ZN(
        n19063) );
  AOI211_X1 U22042 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n19102), .A(n19076), .B(
        n19063), .ZN(n19071) );
  NOR2_X1 U22043 ( .A1(n19092), .A2(n19064), .ZN(n19065) );
  XNOR2_X1 U22044 ( .A(n19066), .B(n19065), .ZN(n19069) );
  OAI22_X1 U22045 ( .A1(n19148), .A2(n19085), .B1(n19067), .B2(n19109), .ZN(
        n19068) );
  AOI21_X1 U22046 ( .B1(n19069), .B2(n19094), .A(n19068), .ZN(n19070) );
  OAI211_X1 U22047 ( .C1(n10052), .C2(n19072), .A(n19071), .B(n19070), .ZN(
        P2_U2849) );
  AOI22_X1 U22048 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19114), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19107), .ZN(n19073) );
  OAI21_X1 U22049 ( .B1(n19105), .B2(n19074), .A(n19073), .ZN(n19075) );
  AOI211_X1 U22050 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19102), .A(n19076), .B(
        n19075), .ZN(n19084) );
  NAND2_X1 U22051 ( .A1(n13929), .A2(n19077), .ZN(n19078) );
  XNOR2_X1 U22052 ( .A(n19079), .B(n19078), .ZN(n19082) );
  AOI22_X1 U22053 ( .A1(n19082), .A2(n19094), .B1(n19081), .B2(n19080), .ZN(
        n19083) );
  OAI211_X1 U22054 ( .C1(n19085), .C2(n19155), .A(n19084), .B(n19083), .ZN(
        P2_U2850) );
  OAI22_X1 U22055 ( .A1(n19087), .A2(n10877), .B1(n19086), .B2(n19105), .ZN(
        n19088) );
  AOI211_X1 U22056 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19102), .A(n19235), .B(
        n19088), .ZN(n19100) );
  AOI22_X1 U22057 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19114), .B1(
        n19101), .B2(n19158), .ZN(n19099) );
  OAI22_X1 U22058 ( .A1(n19160), .A2(n19089), .B1(n19109), .B2(n19236), .ZN(
        n19090) );
  INV_X1 U22059 ( .A(n19090), .ZN(n19098) );
  INV_X1 U22060 ( .A(n19243), .ZN(n19096) );
  NOR2_X1 U22061 ( .A1(n19092), .A2(n19091), .ZN(n19095) );
  NAND2_X1 U22062 ( .A1(n19096), .A2(n19095), .ZN(n19093) );
  OAI211_X1 U22063 ( .C1(n19096), .C2(n19095), .A(n19094), .B(n19093), .ZN(
        n19097) );
  NAND4_X1 U22064 ( .A1(n19100), .A2(n19099), .A3(n19098), .A4(n19097), .ZN(
        P2_U2851) );
  AOI22_X1 U22065 ( .A1(n19102), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19101), 
        .B2(n19183), .ZN(n19103) );
  OAI21_X1 U22066 ( .B1(n19105), .B2(n19104), .A(n19103), .ZN(n19106) );
  AOI21_X1 U22067 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19107), .A(n19106), .ZN(
        n19108) );
  OAI21_X1 U22068 ( .B1(n19110), .B2(n19109), .A(n19108), .ZN(n19111) );
  AOI21_X1 U22069 ( .B1(n19520), .B2(n19112), .A(n19111), .ZN(n19116) );
  OAI21_X1 U22070 ( .B1(n19114), .B2(n19113), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19115) );
  OAI211_X1 U22071 ( .C1(n19118), .C2(n19117), .A(n19116), .B(n19115), .ZN(
        P2_U2855) );
  AOI22_X1 U22072 ( .A1(n19120), .A2(BUF1_REG_31__SCAN_IN), .B1(n19119), .B2(
        n19179), .ZN(n19123) );
  AOI22_X1 U22073 ( .A1(n19121), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19178), .ZN(n19122) );
  NAND2_X1 U22074 ( .A1(n19123), .A2(n19122), .ZN(P2_U2888) );
  OAI222_X1 U22075 ( .A1(n19125), .A2(n19156), .B1(n13450), .B2(n19147), .C1(
        n19124), .C2(n19186), .ZN(P2_U2904) );
  INV_X1 U22076 ( .A(n19126), .ZN(n19128) );
  AOI22_X1 U22077 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19178), .B1(n19228), 
        .B2(n19149), .ZN(n19127) );
  OAI21_X1 U22078 ( .B1(n19156), .B2(n19128), .A(n19127), .ZN(P2_U2905) );
  INV_X1 U22079 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19197) );
  OAI222_X1 U22080 ( .A1(n19130), .A2(n19156), .B1(n19197), .B2(n19147), .C1(
        n19186), .C2(n19129), .ZN(P2_U2906) );
  AOI22_X1 U22081 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19178), .B1(n19131), 
        .B2(n19149), .ZN(n19132) );
  OAI21_X1 U22082 ( .B1(n19156), .B2(n19133), .A(n19132), .ZN(P2_U2907) );
  INV_X1 U22083 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19201) );
  OAI222_X1 U22084 ( .A1(n19135), .A2(n19156), .B1(n19201), .B2(n19147), .C1(
        n19186), .C2(n19134), .ZN(P2_U2908) );
  AOI22_X1 U22085 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19178), .B1(n19136), 
        .B2(n19149), .ZN(n19137) );
  OAI21_X1 U22086 ( .B1(n19156), .B2(n19138), .A(n19137), .ZN(P2_U2909) );
  AOI22_X1 U22087 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19178), .B1(n19139), .B2(
        n19149), .ZN(n19140) );
  OAI21_X1 U22088 ( .B1(n19156), .B2(n19141), .A(n19140), .ZN(P2_U2910) );
  AOI22_X1 U22089 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19178), .B1(n19142), .B2(
        n19149), .ZN(n19143) );
  OAI21_X1 U22090 ( .B1(n19156), .B2(n19144), .A(n19143), .ZN(P2_U2911) );
  INV_X1 U22091 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19209) );
  OAI222_X1 U22092 ( .A1(n19145), .A2(n19156), .B1(n19209), .B2(n19147), .C1(
        n19186), .C2(n19294), .ZN(P2_U2912) );
  INV_X1 U22093 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19211) );
  INV_X1 U22094 ( .A(n19146), .ZN(n19284) );
  OAI222_X1 U22095 ( .A1(n19148), .A2(n19156), .B1(n19211), .B2(n19147), .C1(
        n19186), .C2(n19284), .ZN(P2_U2913) );
  AOI22_X1 U22096 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19178), .B1(n19150), .B2(
        n19149), .ZN(n19154) );
  AOI21_X1 U22097 ( .B1(n19962), .B2(n19961), .A(n19151), .ZN(n19167) );
  XNOR2_X1 U22098 ( .A(n19521), .B(n19957), .ZN(n19166) );
  NOR2_X1 U22099 ( .A1(n19167), .A2(n19166), .ZN(n19165) );
  AOI21_X1 U22100 ( .B1(n19521), .B2(n19957), .A(n19165), .ZN(n19152) );
  NOR2_X1 U22101 ( .A1(n19152), .A2(n19158), .ZN(n19159) );
  OR3_X1 U22102 ( .A1(n19159), .A2(n19160), .A3(n19174), .ZN(n19153) );
  OAI211_X1 U22103 ( .C1(n19156), .C2(n19155), .A(n19154), .B(n19153), .ZN(
        P2_U2914) );
  INV_X1 U22104 ( .A(n19157), .ZN(n19273) );
  AOI22_X1 U22105 ( .A1(n19179), .A2(n19158), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19178), .ZN(n19163) );
  XOR2_X1 U22106 ( .A(n19160), .B(n19159), .Z(n19161) );
  NAND2_X1 U22107 ( .A1(n19161), .A2(n19181), .ZN(n19162) );
  OAI211_X1 U22108 ( .C1(n19273), .C2(n19186), .A(n19163), .B(n19162), .ZN(
        P2_U2915) );
  INV_X1 U22109 ( .A(n19957), .ZN(n19164) );
  AOI22_X1 U22110 ( .A1(n19179), .A2(n19164), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19178), .ZN(n19170) );
  AOI21_X1 U22111 ( .B1(n19167), .B2(n19166), .A(n19165), .ZN(n19168) );
  OR2_X1 U22112 ( .A1(n19168), .A2(n19174), .ZN(n19169) );
  OAI211_X1 U22113 ( .C1(n19171), .C2(n19186), .A(n19170), .B(n19169), .ZN(
        P2_U2916) );
  AOI22_X1 U22114 ( .A1(n19179), .A2(n19976), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19178), .ZN(n19177) );
  AOI21_X1 U22115 ( .B1(n19180), .B2(n19173), .A(n19172), .ZN(n19175) );
  OR2_X1 U22116 ( .A1(n19175), .A2(n19174), .ZN(n19176) );
  OAI211_X1 U22117 ( .C1(n19265), .C2(n19186), .A(n19177), .B(n19176), .ZN(
        P2_U2918) );
  AOI22_X1 U22118 ( .A1(n19179), .A2(n19183), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19178), .ZN(n19185) );
  INV_X1 U22119 ( .A(n19180), .ZN(n19182) );
  OAI211_X1 U22120 ( .C1(n19520), .C2(n19183), .A(n19182), .B(n19181), .ZN(
        n19184) );
  OAI211_X1 U22121 ( .C1(n19260), .C2(n19186), .A(n19185), .B(n19184), .ZN(
        P2_U2919) );
  NOR2_X1 U22122 ( .A1(n19191), .A2(n19187), .ZN(P2_U2920) );
  INV_X1 U22123 ( .A(n19188), .ZN(n19189) );
  AOI22_X1 U22124 ( .A1(n19189), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n19224), .ZN(n19190) );
  OAI21_X1 U22125 ( .B1(n19192), .B2(n19191), .A(n19190), .ZN(P2_U2921) );
  AOI22_X1 U22126 ( .A1(n19224), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19193) );
  OAI21_X1 U22127 ( .B1(n13450), .B2(n19226), .A(n19193), .ZN(P2_U2936) );
  INV_X1 U22128 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19195) );
  AOI22_X1 U22129 ( .A1(n19224), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U22130 ( .B1(n19195), .B2(n19226), .A(n19194), .ZN(P2_U2937) );
  AOI22_X1 U22131 ( .A1(n19224), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19196) );
  OAI21_X1 U22132 ( .B1(n19197), .B2(n19226), .A(n19196), .ZN(P2_U2938) );
  AOI22_X1 U22133 ( .A1(n19224), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U22134 ( .B1(n19199), .B2(n19226), .A(n19198), .ZN(P2_U2939) );
  AOI22_X1 U22135 ( .A1(n19220), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U22136 ( .B1(n19201), .B2(n19226), .A(n19200), .ZN(P2_U2940) );
  AOI22_X1 U22137 ( .A1(n19220), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19202) );
  OAI21_X1 U22138 ( .B1(n19203), .B2(n19226), .A(n19202), .ZN(P2_U2941) );
  AOI22_X1 U22139 ( .A1(n19220), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19204) );
  OAI21_X1 U22140 ( .B1(n19205), .B2(n19226), .A(n19204), .ZN(P2_U2942) );
  AOI22_X1 U22141 ( .A1(n19220), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19206) );
  OAI21_X1 U22142 ( .B1(n19207), .B2(n19226), .A(n19206), .ZN(P2_U2943) );
  AOI22_X1 U22143 ( .A1(n19220), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19208) );
  OAI21_X1 U22144 ( .B1(n19209), .B2(n19226), .A(n19208), .ZN(P2_U2944) );
  AOI22_X1 U22145 ( .A1(n19220), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19210) );
  OAI21_X1 U22146 ( .B1(n19211), .B2(n19226), .A(n19210), .ZN(P2_U2945) );
  INV_X1 U22147 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19213) );
  AOI22_X1 U22148 ( .A1(n19220), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19212) );
  OAI21_X1 U22149 ( .B1(n19213), .B2(n19226), .A(n19212), .ZN(P2_U2946) );
  INV_X1 U22150 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19215) );
  AOI22_X1 U22151 ( .A1(n19220), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19214) );
  OAI21_X1 U22152 ( .B1(n19215), .B2(n19226), .A(n19214), .ZN(P2_U2947) );
  INV_X1 U22153 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19217) );
  AOI22_X1 U22154 ( .A1(n19220), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19216) );
  OAI21_X1 U22155 ( .B1(n19217), .B2(n19226), .A(n19216), .ZN(P2_U2948) );
  INV_X1 U22156 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19219) );
  AOI22_X1 U22157 ( .A1(n19220), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19218) );
  OAI21_X1 U22158 ( .B1(n19219), .B2(n19226), .A(n19218), .ZN(P2_U2949) );
  INV_X1 U22159 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19222) );
  AOI22_X1 U22160 ( .A1(n19220), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19221) );
  OAI21_X1 U22161 ( .B1(n19222), .B2(n19226), .A(n19221), .ZN(P2_U2950) );
  AOI22_X1 U22162 ( .A1(n19224), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19223), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19225) );
  OAI21_X1 U22163 ( .B1(n19227), .B2(n19226), .A(n19225), .ZN(P2_U2951) );
  AOI22_X1 U22164 ( .A1(n19232), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19231), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19230) );
  NAND2_X1 U22165 ( .A1(n19229), .A2(n19228), .ZN(n19233) );
  NAND2_X1 U22166 ( .A1(n19230), .A2(n19233), .ZN(P2_U2966) );
  AOI22_X1 U22167 ( .A1(n19232), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n19231), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19234) );
  NAND2_X1 U22168 ( .A1(n19234), .A2(n19233), .ZN(P2_U2981) );
  AOI22_X1 U22169 ( .A1(n19245), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19235), .ZN(n19242) );
  OAI22_X1 U22170 ( .A1(n19238), .A2(n19237), .B1(n14106), .B2(n19236), .ZN(
        n19239) );
  AOI21_X1 U22171 ( .B1(n19248), .B2(n19240), .A(n19239), .ZN(n19241) );
  OAI211_X1 U22172 ( .C1(n19253), .C2(n19243), .A(n19242), .B(n19241), .ZN(
        P2_U3010) );
  INV_X1 U22173 ( .A(n19244), .ZN(n19247) );
  AOI22_X1 U22174 ( .A1(n19247), .A2(n19246), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19245), .ZN(n19258) );
  NAND2_X1 U22175 ( .A1(n19249), .A2(n19248), .ZN(n19250) );
  OAI211_X1 U22176 ( .C1(n19253), .C2(n19252), .A(n19251), .B(n19250), .ZN(
        n19254) );
  AOI21_X1 U22177 ( .B1(n19256), .B2(n19255), .A(n19254), .ZN(n19257) );
  NAND2_X1 U22178 ( .A1(n19258), .A2(n19257), .ZN(P2_U3012) );
  INV_X1 U22179 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19263) );
  AOI22_X1 U22180 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19295), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19296), .ZN(n19800) );
  INV_X1 U22181 ( .A(n19800), .ZN(n19715) );
  NAND2_X1 U22182 ( .A1(n19259), .A2(n19291), .ZN(n19622) );
  AOI22_X1 U22183 ( .A1(n19842), .A2(n19715), .B1(n19293), .B2(n19788), .ZN(
        n19262) );
  NOR2_X2 U22184 ( .A1(n19260), .A2(n19495), .ZN(n19789) );
  AOI22_X1 U22185 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19295), .ZN(n19718) );
  AOI22_X1 U22186 ( .A1(n19789), .A2(n19297), .B1(n19323), .B2(n19797), .ZN(
        n19261) );
  OAI211_X1 U22187 ( .C1(n19300), .C2(n19263), .A(n19262), .B(n19261), .ZN(
        P2_U3048) );
  INV_X1 U22188 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19268) );
  AOI22_X2 U22189 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19295), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19296), .ZN(n19806) );
  INV_X1 U22190 ( .A(n19806), .ZN(n19759) );
  NAND2_X1 U22191 ( .A1(n19264), .A2(n19291), .ZN(n19634) );
  AOI22_X1 U22192 ( .A1(n19842), .A2(n19759), .B1(n19293), .B2(n19801), .ZN(
        n19267) );
  NOR2_X2 U22193 ( .A1(n19265), .A2(n19495), .ZN(n19802) );
  AOI22_X1 U22194 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19295), .ZN(n19762) );
  AOI22_X1 U22195 ( .A1(n19802), .A2(n19297), .B1(n19323), .B2(n19803), .ZN(
        n19266) );
  OAI211_X1 U22196 ( .C1(n19300), .C2(n19268), .A(n19267), .B(n19266), .ZN(
        P2_U3049) );
  INV_X1 U22197 ( .A(n19812), .ZN(n19721) );
  NAND2_X1 U22198 ( .A1(n13020), .A2(n19291), .ZN(n19639) );
  AOI22_X1 U22199 ( .A1(n19842), .A2(n19721), .B1(n19293), .B2(n19807), .ZN(
        n19271) );
  NOR2_X2 U22200 ( .A1(n19269), .A2(n19495), .ZN(n19808) );
  AOI22_X1 U22201 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19295), .ZN(n19724) );
  AOI22_X1 U22202 ( .A1(n19808), .A2(n19297), .B1(n19323), .B2(n19809), .ZN(
        n19270) );
  OAI211_X1 U22203 ( .C1(n19300), .C2(n19272), .A(n19271), .B(n19270), .ZN(
        P2_U3050) );
  AOI22_X1 U22204 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19295), .ZN(n19824) );
  INV_X1 U22205 ( .A(n19824), .ZN(n19729) );
  NAND2_X1 U22206 ( .A1(n10333), .A2(n19291), .ZN(n19649) );
  INV_X1 U22207 ( .A(n19649), .ZN(n19819) );
  AOI22_X1 U22208 ( .A1(n19842), .A2(n19729), .B1(n19293), .B2(n19819), .ZN(
        n19275) );
  NOR2_X2 U22209 ( .A1(n19273), .A2(n19495), .ZN(n19820) );
  AOI22_X1 U22210 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19295), .ZN(n19732) );
  INV_X1 U22211 ( .A(n19732), .ZN(n19821) );
  AOI22_X1 U22212 ( .A1(n19820), .A2(n19297), .B1(n19323), .B2(n19821), .ZN(
        n19274) );
  OAI211_X1 U22213 ( .C1(n19300), .C2(n19276), .A(n19275), .B(n19274), .ZN(
        P2_U3052) );
  AOI22_X1 U22214 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19295), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19296), .ZN(n19830) );
  AOI22_X1 U22215 ( .A1(n19842), .A2(n19769), .B1(n19293), .B2(n19825), .ZN(
        n19281) );
  NOR2_X2 U22216 ( .A1(n19278), .A2(n19495), .ZN(n19826) );
  AOI22_X1 U22217 ( .A1(n19826), .A2(n19297), .B1(n19323), .B2(n19827), .ZN(
        n19280) );
  OAI211_X1 U22218 ( .C1(n19300), .C2(n13606), .A(n19281), .B(n19280), .ZN(
        P2_U3053) );
  AND2_X1 U22219 ( .A1(n19283), .A2(n19291), .ZN(n19831) );
  AOI22_X1 U22220 ( .A1(n19842), .A2(n19735), .B1(n19293), .B2(n19831), .ZN(
        n19286) );
  NOR2_X2 U22221 ( .A1(n19284), .A2(n19495), .ZN(n19832) );
  AOI22_X1 U22222 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19295), .ZN(n19738) );
  AOI22_X1 U22223 ( .A1(n19832), .A2(n19297), .B1(n19323), .B2(n19833), .ZN(
        n19285) );
  OAI211_X1 U22224 ( .C1(n19300), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P2_U3054) );
  NAND2_X1 U22225 ( .A1(n19292), .A2(n19291), .ZN(n19666) );
  AOI22_X1 U22226 ( .A1(n19842), .A2(n19778), .B1(n19293), .B2(n19838), .ZN(
        n19299) );
  NOR2_X2 U22227 ( .A1(n19294), .A2(n19495), .ZN(n19839) );
  AOI22_X1 U22228 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19296), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19295), .ZN(n19784) );
  INV_X1 U22229 ( .A(n19784), .ZN(n19841) );
  AOI22_X1 U22230 ( .A1(n19839), .A2(n19297), .B1(n19323), .B2(n19841), .ZN(
        n19298) );
  OAI211_X1 U22231 ( .C1(n19300), .C2(n11973), .A(n19299), .B(n19298), .ZN(
        P2_U3055) );
  INV_X1 U22232 ( .A(n19301), .ZN(n19302) );
  NOR2_X1 U22233 ( .A1(n19559), .A2(n19360), .ZN(n19321) );
  NOR3_X1 U22234 ( .A1(n19302), .A2(n19321), .A3(n19851), .ZN(n19303) );
  AOI211_X2 U22235 ( .C1(n19304), .C2(n19851), .A(n19849), .B(n19303), .ZN(
        n19322) );
  AOI22_X1 U22236 ( .A1(n19322), .A2(n19789), .B1(n19788), .B2(n19321), .ZN(
        n19308) );
  NAND2_X1 U22237 ( .A1(n19521), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19954) );
  INV_X1 U22238 ( .A(n19954), .ZN(n19494) );
  INV_X1 U22239 ( .A(n19560), .ZN(n19522) );
  NAND2_X1 U22240 ( .A1(n19494), .A2(n19522), .ZN(n19305) );
  AOI21_X1 U22241 ( .B1(n19305), .B2(n19304), .A(n19303), .ZN(n19306) );
  OAI211_X1 U22242 ( .C1(n19321), .C2(n19979), .A(n19306), .B(n19795), .ZN(
        n19324) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19715), .ZN(n19307) );
  OAI211_X1 U22244 ( .C1(n19718), .C2(n19358), .A(n19308), .B(n19307), .ZN(
        P2_U3056) );
  AOI22_X1 U22245 ( .A1(n19322), .A2(n19802), .B1(n19801), .B2(n19321), .ZN(
        n19310) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19759), .ZN(n19309) );
  OAI211_X1 U22247 ( .C1(n19762), .C2(n19358), .A(n19310), .B(n19309), .ZN(
        P2_U3057) );
  AOI22_X1 U22248 ( .A1(n19322), .A2(n19808), .B1(n19807), .B2(n19321), .ZN(
        n19312) );
  AOI22_X1 U22249 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19721), .ZN(n19311) );
  OAI211_X1 U22250 ( .C1(n19724), .C2(n19358), .A(n19312), .B(n19311), .ZN(
        P2_U3058) );
  AOI22_X1 U22251 ( .A1(n19322), .A2(n19814), .B1(n19813), .B2(n19321), .ZN(
        n19314) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19725), .ZN(n19313) );
  OAI211_X1 U22253 ( .C1(n19728), .C2(n19358), .A(n19314), .B(n19313), .ZN(
        P2_U3059) );
  AOI22_X1 U22254 ( .A1(n19322), .A2(n19820), .B1(n19819), .B2(n19321), .ZN(
        n19316) );
  AOI22_X1 U22255 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19729), .ZN(n19315) );
  OAI211_X1 U22256 ( .C1(n19732), .C2(n19358), .A(n19316), .B(n19315), .ZN(
        P2_U3060) );
  AOI22_X1 U22257 ( .A1(n19322), .A2(n19826), .B1(n19825), .B2(n19321), .ZN(
        n19318) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19769), .ZN(n19317) );
  OAI211_X1 U22259 ( .C1(n19772), .C2(n19358), .A(n19318), .B(n19317), .ZN(
        P2_U3061) );
  AOI22_X1 U22260 ( .A1(n19322), .A2(n19832), .B1(n19831), .B2(n19321), .ZN(
        n19320) );
  AOI22_X1 U22261 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19735), .ZN(n19319) );
  OAI211_X1 U22262 ( .C1(n19738), .C2(n19358), .A(n19320), .B(n19319), .ZN(
        P2_U3062) );
  AOI22_X1 U22263 ( .A1(n19322), .A2(n19839), .B1(n19838), .B2(n19321), .ZN(
        n19326) );
  AOI22_X1 U22264 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19324), .B1(
        n19323), .B2(n19778), .ZN(n19325) );
  OAI211_X1 U22265 ( .C1(n19784), .C2(n19358), .A(n19326), .B(n19325), .ZN(
        P2_U3063) );
  NOR2_X1 U22266 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19978), .ZN(
        n19328) );
  AND2_X1 U22267 ( .A1(n19328), .A2(n19327), .ZN(n19353) );
  OAI21_X1 U22268 ( .B1(n19330), .B2(n19353), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19329) );
  OR2_X1 U22269 ( .A1(n19591), .A2(n19360), .ZN(n19333) );
  NAND2_X1 U22270 ( .A1(n19329), .A2(n19333), .ZN(n19354) );
  AOI22_X1 U22271 ( .A1(n19354), .A2(n19789), .B1(n19788), .B2(n19353), .ZN(
        n19339) );
  INV_X1 U22272 ( .A(n19330), .ZN(n19332) );
  INV_X1 U22273 ( .A(n19353), .ZN(n19331) );
  OAI21_X1 U22274 ( .B1(n19332), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19331), 
        .ZN(n19336) );
  OAI21_X1 U22275 ( .B1(n19384), .B2(n19348), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19334) );
  NAND2_X1 U22276 ( .A1(n19334), .A2(n19333), .ZN(n19335) );
  MUX2_X1 U22277 ( .A(n19336), .B(n19335), .S(n19945), .Z(n19337) );
  NAND2_X1 U22278 ( .A1(n19337), .A2(n19795), .ZN(n19355) );
  AOI22_X1 U22279 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19355), .B1(
        n19384), .B2(n19797), .ZN(n19338) );
  OAI211_X1 U22280 ( .C1(n19800), .C2(n19358), .A(n19339), .B(n19338), .ZN(
        P2_U3064) );
  AOI22_X1 U22281 ( .A1(n19354), .A2(n19802), .B1(n19801), .B2(n19353), .ZN(
        n19341) );
  AOI22_X1 U22282 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19355), .B1(
        n19384), .B2(n19803), .ZN(n19340) );
  OAI211_X1 U22283 ( .C1(n19806), .C2(n19358), .A(n19341), .B(n19340), .ZN(
        P2_U3065) );
  AOI22_X1 U22284 ( .A1(n19354), .A2(n19808), .B1(n19807), .B2(n19353), .ZN(
        n19343) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19355), .B1(
        n19384), .B2(n19809), .ZN(n19342) );
  OAI211_X1 U22286 ( .C1(n19812), .C2(n19358), .A(n19343), .B(n19342), .ZN(
        P2_U3066) );
  AOI22_X1 U22287 ( .A1(n19354), .A2(n19814), .B1(n19813), .B2(n19353), .ZN(
        n19345) );
  INV_X1 U22288 ( .A(n19728), .ZN(n19815) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19355), .B1(
        n19384), .B2(n19815), .ZN(n19344) );
  OAI211_X1 U22290 ( .C1(n19818), .C2(n19358), .A(n19345), .B(n19344), .ZN(
        P2_U3067) );
  AOI22_X1 U22291 ( .A1(n19354), .A2(n19820), .B1(n19819), .B2(n19353), .ZN(
        n19347) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19355), .B1(
        n19384), .B2(n19821), .ZN(n19346) );
  OAI211_X1 U22293 ( .C1(n19824), .C2(n19358), .A(n19347), .B(n19346), .ZN(
        P2_U3068) );
  AOI22_X1 U22294 ( .A1(n19354), .A2(n19826), .B1(n19825), .B2(n19353), .ZN(
        n19350) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19355), .B1(
        n19348), .B2(n19769), .ZN(n19349) );
  OAI211_X1 U22296 ( .C1(n19772), .C2(n19393), .A(n19350), .B(n19349), .ZN(
        P2_U3069) );
  AOI22_X1 U22297 ( .A1(n19354), .A2(n19832), .B1(n19831), .B2(n19353), .ZN(
        n19352) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19355), .B1(
        n19384), .B2(n19833), .ZN(n19351) );
  OAI211_X1 U22299 ( .C1(n19836), .C2(n19358), .A(n19352), .B(n19351), .ZN(
        P2_U3070) );
  AOI22_X1 U22300 ( .A1(n19354), .A2(n19839), .B1(n19838), .B2(n19353), .ZN(
        n19357) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19355), .B1(
        n19384), .B2(n19841), .ZN(n19356) );
  OAI211_X1 U22302 ( .C1(n19847), .C2(n19358), .A(n19357), .B(n19356), .ZN(
        P2_U3071) );
  NOR2_X1 U22303 ( .A1(n19617), .A2(n19360), .ZN(n19383) );
  INV_X1 U22304 ( .A(n19383), .ZN(n19387) );
  OAI22_X1 U22305 ( .A1(n19424), .A2(n19718), .B1(n19387), .B2(n19622), .ZN(
        n19359) );
  INV_X1 U22306 ( .A(n19359), .ZN(n19370) );
  OAI21_X1 U22307 ( .B1(n19954), .B2(n19946), .A(n19945), .ZN(n19368) );
  NOR2_X1 U22308 ( .A1(n19978), .A2(n19360), .ZN(n19364) );
  INV_X1 U22309 ( .A(n19361), .ZN(n19365) );
  OAI21_X1 U22310 ( .B1(n19365), .B2(n19851), .A(n19979), .ZN(n19362) );
  AOI21_X1 U22311 ( .B1(n19362), .B2(n19387), .A(n19495), .ZN(n19363) );
  OAI21_X1 U22312 ( .B1(n19368), .B2(n19364), .A(n19363), .ZN(n19390) );
  INV_X1 U22313 ( .A(n19364), .ZN(n19367) );
  OAI21_X1 U22314 ( .B1(n19365), .B2(n19383), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19366) );
  OAI21_X1 U22315 ( .B1(n19368), .B2(n19367), .A(n19366), .ZN(n19389) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19390), .B1(
        n19789), .B2(n19389), .ZN(n19369) );
  OAI211_X1 U22317 ( .C1(n19800), .C2(n19393), .A(n19370), .B(n19369), .ZN(
        P2_U3072) );
  OAI22_X1 U22318 ( .A1(n19424), .A2(n19762), .B1(n19387), .B2(n19634), .ZN(
        n19371) );
  INV_X1 U22319 ( .A(n19371), .ZN(n19373) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19390), .B1(
        n19802), .B2(n19389), .ZN(n19372) );
  OAI211_X1 U22321 ( .C1(n19806), .C2(n19393), .A(n19373), .B(n19372), .ZN(
        P2_U3073) );
  AOI22_X1 U22322 ( .A1(n19384), .A2(n19721), .B1(n19383), .B2(n19807), .ZN(
        n19375) );
  AOI22_X1 U22323 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19390), .B1(
        n19808), .B2(n19389), .ZN(n19374) );
  OAI211_X1 U22324 ( .C1(n19724), .C2(n19424), .A(n19375), .B(n19374), .ZN(
        P2_U3074) );
  AOI22_X1 U22325 ( .A1(n19416), .A2(n19815), .B1(n19813), .B2(n19383), .ZN(
        n19377) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19390), .B1(
        n19814), .B2(n19389), .ZN(n19376) );
  OAI211_X1 U22327 ( .C1(n19818), .C2(n19393), .A(n19377), .B(n19376), .ZN(
        P2_U3075) );
  OAI22_X1 U22328 ( .A1(n19393), .A2(n19824), .B1(n19387), .B2(n19649), .ZN(
        n19378) );
  INV_X1 U22329 ( .A(n19378), .ZN(n19380) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19390), .B1(
        n19820), .B2(n19389), .ZN(n19379) );
  OAI211_X1 U22331 ( .C1(n19732), .C2(n19424), .A(n19380), .B(n19379), .ZN(
        P2_U3076) );
  AOI22_X1 U22332 ( .A1(n19384), .A2(n19769), .B1(n19383), .B2(n19825), .ZN(
        n19382) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19390), .B1(
        n19826), .B2(n19389), .ZN(n19381) );
  OAI211_X1 U22334 ( .C1(n19772), .C2(n19424), .A(n19382), .B(n19381), .ZN(
        P2_U3077) );
  AOI22_X1 U22335 ( .A1(n19384), .A2(n19735), .B1(n19383), .B2(n19831), .ZN(
        n19386) );
  AOI22_X1 U22336 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19390), .B1(
        n19832), .B2(n19389), .ZN(n19385) );
  OAI211_X1 U22337 ( .C1(n19738), .C2(n19424), .A(n19386), .B(n19385), .ZN(
        P2_U3078) );
  OAI22_X1 U22338 ( .A1(n19424), .A2(n19784), .B1(n19387), .B2(n19666), .ZN(
        n19388) );
  INV_X1 U22339 ( .A(n19388), .ZN(n19392) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19390), .B1(
        n19839), .B2(n19389), .ZN(n19391) );
  OAI211_X1 U22341 ( .C1(n19847), .C2(n19393), .A(n19392), .B(n19391), .ZN(
        P2_U3079) );
  INV_X1 U22342 ( .A(n19394), .ZN(n19396) );
  NAND2_X1 U22343 ( .A1(n19396), .A2(n19395), .ZN(n19680) );
  NOR2_X1 U22344 ( .A1(n19680), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19403) );
  INV_X1 U22345 ( .A(n19403), .ZN(n19398) );
  NOR3_X1 U22346 ( .A1(n19968), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19426) );
  INV_X1 U22347 ( .A(n19426), .ZN(n19430) );
  NOR2_X1 U22348 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19430), .ZN(
        n19419) );
  OAI21_X1 U22349 ( .B1(n12438), .B2(n19419), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19397) );
  OAI21_X1 U22350 ( .B1(n19953), .B2(n19398), .A(n19397), .ZN(n19420) );
  AOI22_X1 U22351 ( .A1(n19420), .A2(n19789), .B1(n19788), .B2(n19419), .ZN(
        n19405) );
  AOI21_X1 U22352 ( .B1(n19424), .B2(n19448), .A(n19457), .ZN(n19402) );
  OAI21_X1 U22353 ( .B1(n12438), .B2(n19851), .A(n19979), .ZN(n19400) );
  INV_X1 U22354 ( .A(n19419), .ZN(n19399) );
  NAND2_X1 U22355 ( .A1(n19400), .A2(n19399), .ZN(n19401) );
  OAI211_X1 U22356 ( .C1(n19403), .C2(n19402), .A(n19401), .B(n19795), .ZN(
        n19421) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19421), .B1(
        n19451), .B2(n19797), .ZN(n19404) );
  OAI211_X1 U22358 ( .C1(n19800), .C2(n19424), .A(n19405), .B(n19404), .ZN(
        P2_U3080) );
  AOI22_X1 U22359 ( .A1(n19420), .A2(n19802), .B1(n19801), .B2(n19419), .ZN(
        n19407) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19421), .B1(
        n19451), .B2(n19803), .ZN(n19406) );
  OAI211_X1 U22361 ( .C1(n19806), .C2(n19424), .A(n19407), .B(n19406), .ZN(
        P2_U3081) );
  AOI22_X1 U22362 ( .A1(n19420), .A2(n19808), .B1(n19807), .B2(n19419), .ZN(
        n19409) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19421), .B1(
        n19451), .B2(n19809), .ZN(n19408) );
  OAI211_X1 U22364 ( .C1(n19812), .C2(n19424), .A(n19409), .B(n19408), .ZN(
        P2_U3082) );
  AOI22_X1 U22365 ( .A1(n19420), .A2(n19814), .B1(n19813), .B2(n19419), .ZN(
        n19411) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19421), .B1(
        n19416), .B2(n19725), .ZN(n19410) );
  OAI211_X1 U22367 ( .C1(n19728), .C2(n19448), .A(n19411), .B(n19410), .ZN(
        P2_U3083) );
  AOI22_X1 U22368 ( .A1(n19420), .A2(n19820), .B1(n19819), .B2(n19419), .ZN(
        n19413) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19421), .B1(
        n19416), .B2(n19729), .ZN(n19412) );
  OAI211_X1 U22370 ( .C1(n19732), .C2(n19448), .A(n19413), .B(n19412), .ZN(
        P2_U3084) );
  AOI22_X1 U22371 ( .A1(n19420), .A2(n19826), .B1(n19825), .B2(n19419), .ZN(
        n19415) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19421), .B1(
        n19416), .B2(n19769), .ZN(n19414) );
  OAI211_X1 U22373 ( .C1(n19772), .C2(n19448), .A(n19415), .B(n19414), .ZN(
        P2_U3085) );
  AOI22_X1 U22374 ( .A1(n19420), .A2(n19832), .B1(n19831), .B2(n19419), .ZN(
        n19418) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19421), .B1(
        n19416), .B2(n19735), .ZN(n19417) );
  OAI211_X1 U22376 ( .C1(n19738), .C2(n19448), .A(n19418), .B(n19417), .ZN(
        P2_U3086) );
  AOI22_X1 U22377 ( .A1(n19420), .A2(n19839), .B1(n19838), .B2(n19419), .ZN(
        n19423) );
  AOI22_X1 U22378 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19421), .B1(
        n19451), .B2(n19841), .ZN(n19422) );
  OAI211_X1 U22379 ( .C1(n19847), .C2(n19424), .A(n19423), .B(n19422), .ZN(
        P2_U3087) );
  NOR2_X1 U22380 ( .A1(n19987), .A2(n19430), .ZN(n19464) );
  AOI22_X1 U22381 ( .A1(n19451), .A2(n19715), .B1(n19464), .B2(n19788), .ZN(
        n19433) );
  OAI21_X1 U22382 ( .B1(n19954), .B2(n19709), .A(n19945), .ZN(n19431) );
  INV_X1 U22383 ( .A(n19464), .ZN(n19442) );
  OAI211_X1 U22384 ( .C1(n19427), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19442), 
        .B(n19953), .ZN(n19425) );
  OAI211_X1 U22385 ( .C1(n19431), .C2(n19426), .A(n19795), .B(n19425), .ZN(
        n19453) );
  INV_X1 U22386 ( .A(n19427), .ZN(n19428) );
  OAI21_X1 U22387 ( .B1(n19428), .B2(n19464), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19429) );
  OAI21_X1 U22388 ( .B1(n19431), .B2(n19430), .A(n19429), .ZN(n19452) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19453), .B1(
        n19789), .B2(n19452), .ZN(n19432) );
  OAI211_X1 U22390 ( .C1(n19718), .C2(n19482), .A(n19433), .B(n19432), .ZN(
        P2_U3088) );
  OAI22_X1 U22391 ( .A1(n19482), .A2(n19762), .B1(n19634), .B2(n19442), .ZN(
        n19434) );
  INV_X1 U22392 ( .A(n19434), .ZN(n19436) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19453), .B1(
        n19802), .B2(n19452), .ZN(n19435) );
  OAI211_X1 U22394 ( .C1(n19806), .C2(n19448), .A(n19436), .B(n19435), .ZN(
        P2_U3089) );
  OAI22_X1 U22395 ( .A1(n19482), .A2(n19724), .B1(n19442), .B2(n19639), .ZN(
        n19437) );
  INV_X1 U22396 ( .A(n19437), .ZN(n19439) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19453), .B1(
        n19808), .B2(n19452), .ZN(n19438) );
  OAI211_X1 U22398 ( .C1(n19812), .C2(n19448), .A(n19439), .B(n19438), .ZN(
        P2_U3090) );
  AOI22_X1 U22399 ( .A1(n19487), .A2(n19815), .B1(n19813), .B2(n19464), .ZN(
        n19441) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19453), .B1(
        n19814), .B2(n19452), .ZN(n19440) );
  OAI211_X1 U22401 ( .C1(n19818), .C2(n19448), .A(n19441), .B(n19440), .ZN(
        P2_U3091) );
  OAI22_X1 U22402 ( .A1(n19448), .A2(n19824), .B1(n19442), .B2(n19649), .ZN(
        n19443) );
  INV_X1 U22403 ( .A(n19443), .ZN(n19445) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19453), .B1(
        n19820), .B2(n19452), .ZN(n19444) );
  OAI211_X1 U22405 ( .C1(n19732), .C2(n19482), .A(n19445), .B(n19444), .ZN(
        P2_U3092) );
  AOI22_X1 U22406 ( .A1(n19487), .A2(n19827), .B1(n19464), .B2(n19825), .ZN(
        n19447) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19453), .B1(
        n19826), .B2(n19452), .ZN(n19446) );
  OAI211_X1 U22408 ( .C1(n19830), .C2(n19448), .A(n19447), .B(n19446), .ZN(
        P2_U3093) );
  AOI22_X1 U22409 ( .A1(n19451), .A2(n19735), .B1(n19464), .B2(n19831), .ZN(
        n19450) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19453), .B1(
        n19832), .B2(n19452), .ZN(n19449) );
  OAI211_X1 U22411 ( .C1(n19738), .C2(n19482), .A(n19450), .B(n19449), .ZN(
        P2_U3094) );
  AOI22_X1 U22412 ( .A1(n19451), .A2(n19778), .B1(n19464), .B2(n19838), .ZN(
        n19455) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19453), .B1(
        n19839), .B2(n19452), .ZN(n19454) );
  OAI211_X1 U22414 ( .C1(n19784), .C2(n19482), .A(n19455), .B(n19454), .ZN(
        P2_U3095) );
  AOI21_X1 U22415 ( .B1(n19482), .B2(n19519), .A(n19457), .ZN(n19458) );
  NOR2_X1 U22416 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19497), .ZN(
        n19485) );
  AOI221_X1 U22417 ( .B1(n19464), .B2(n19979), .C1(n19458), .C2(n19979), .A(
        n19485), .ZN(n19463) );
  INV_X1 U22418 ( .A(n19485), .ZN(n19459) );
  AND2_X1 U22419 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19459), .ZN(n19460) );
  NAND2_X1 U22420 ( .A1(n19461), .A2(n19460), .ZN(n19467) );
  NAND2_X1 U22421 ( .A1(n19467), .A2(n19795), .ZN(n19462) );
  INV_X1 U22422 ( .A(n19488), .ZN(n19471) );
  NOR2_X1 U22423 ( .A1(n19464), .A2(n19485), .ZN(n19465) );
  OAI21_X1 U22424 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19465), .A(n19851), 
        .ZN(n19466) );
  AOI22_X1 U22425 ( .A1(n19486), .A2(n19789), .B1(n19788), .B2(n19485), .ZN(
        n19469) );
  AOI22_X1 U22426 ( .A1(n19506), .A2(n19797), .B1(n19487), .B2(n19715), .ZN(
        n19468) );
  OAI211_X1 U22427 ( .C1(n19471), .C2(n19470), .A(n19469), .B(n19468), .ZN(
        P2_U3096) );
  AOI22_X1 U22428 ( .A1(n19486), .A2(n19802), .B1(n19801), .B2(n19485), .ZN(
        n19473) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19488), .B1(
        n19506), .B2(n19803), .ZN(n19472) );
  OAI211_X1 U22430 ( .C1(n19806), .C2(n19482), .A(n19473), .B(n19472), .ZN(
        P2_U3097) );
  AOI22_X1 U22431 ( .A1(n19486), .A2(n19808), .B1(n19807), .B2(n19485), .ZN(
        n19475) );
  AOI22_X1 U22432 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19488), .B1(
        n19506), .B2(n19809), .ZN(n19474) );
  OAI211_X1 U22433 ( .C1(n19812), .C2(n19482), .A(n19475), .B(n19474), .ZN(
        P2_U3098) );
  AOI22_X1 U22434 ( .A1(n19486), .A2(n19814), .B1(n19813), .B2(n19485), .ZN(
        n19477) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19725), .ZN(n19476) );
  OAI211_X1 U22436 ( .C1(n19728), .C2(n19519), .A(n19477), .B(n19476), .ZN(
        P2_U3099) );
  AOI22_X1 U22437 ( .A1(n19486), .A2(n19820), .B1(n19819), .B2(n19485), .ZN(
        n19479) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19488), .B1(
        n19506), .B2(n19821), .ZN(n19478) );
  OAI211_X1 U22439 ( .C1(n19824), .C2(n19482), .A(n19479), .B(n19478), .ZN(
        P2_U3100) );
  AOI22_X1 U22440 ( .A1(n19486), .A2(n19826), .B1(n19825), .B2(n19485), .ZN(
        n19481) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19488), .B1(
        n19506), .B2(n19827), .ZN(n19480) );
  OAI211_X1 U22442 ( .C1(n19830), .C2(n19482), .A(n19481), .B(n19480), .ZN(
        P2_U3101) );
  AOI22_X1 U22443 ( .A1(n19486), .A2(n19832), .B1(n19831), .B2(n19485), .ZN(
        n19484) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19735), .ZN(n19483) );
  OAI211_X1 U22445 ( .C1(n19738), .C2(n19519), .A(n19484), .B(n19483), .ZN(
        P2_U3102) );
  AOI22_X1 U22446 ( .A1(n19486), .A2(n19839), .B1(n19838), .B2(n19485), .ZN(
        n19490) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19488), .B1(
        n19487), .B2(n19778), .ZN(n19489) );
  OAI211_X1 U22448 ( .C1(n19784), .C2(n19519), .A(n19490), .B(n19489), .ZN(
        P2_U3103) );
  INV_X1 U22449 ( .A(n19492), .ZN(n19493) );
  NOR3_X1 U22450 ( .A1(n19493), .A2(n19530), .A3(n19851), .ZN(n19496) );
  AOI211_X2 U22451 ( .C1(n19497), .C2(n19851), .A(n19849), .B(n19496), .ZN(
        n19515) );
  AOI22_X1 U22452 ( .A1(n19515), .A2(n19789), .B1(n19530), .B2(n19788), .ZN(
        n19501) );
  INV_X1 U22453 ( .A(n19952), .ZN(n19790) );
  NAND2_X1 U22454 ( .A1(n19494), .A2(n19790), .ZN(n19498) );
  AOI211_X1 U22455 ( .C1(n19498), .C2(n19497), .A(n19496), .B(n19495), .ZN(
        n19499) );
  OAI21_X1 U22456 ( .B1(n19530), .B2(n19979), .A(n19499), .ZN(n19516) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19516), .B1(
        n19506), .B2(n19715), .ZN(n19500) );
  OAI211_X1 U22458 ( .C1(n19718), .C2(n19558), .A(n19501), .B(n19500), .ZN(
        P2_U3104) );
  AOI22_X1 U22459 ( .A1(n19515), .A2(n19802), .B1(n19530), .B2(n19801), .ZN(
        n19503) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19516), .B1(
        n19546), .B2(n19803), .ZN(n19502) );
  OAI211_X1 U22461 ( .C1(n19806), .C2(n19519), .A(n19503), .B(n19502), .ZN(
        P2_U3105) );
  AOI22_X1 U22462 ( .A1(n19515), .A2(n19808), .B1(n19530), .B2(n19807), .ZN(
        n19505) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19516), .B1(
        n19506), .B2(n19721), .ZN(n19504) );
  OAI211_X1 U22464 ( .C1(n19724), .C2(n19558), .A(n19505), .B(n19504), .ZN(
        P2_U3106) );
  AOI22_X1 U22465 ( .A1(n19515), .A2(n19814), .B1(n19530), .B2(n19813), .ZN(
        n19508) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19516), .B1(
        n19506), .B2(n19725), .ZN(n19507) );
  OAI211_X1 U22467 ( .C1(n19728), .C2(n19558), .A(n19508), .B(n19507), .ZN(
        P2_U3107) );
  AOI22_X1 U22468 ( .A1(n19515), .A2(n19820), .B1(n19530), .B2(n19819), .ZN(
        n19510) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19516), .B1(
        n19546), .B2(n19821), .ZN(n19509) );
  OAI211_X1 U22470 ( .C1(n19824), .C2(n19519), .A(n19510), .B(n19509), .ZN(
        P2_U3108) );
  AOI22_X1 U22471 ( .A1(n19515), .A2(n19826), .B1(n19530), .B2(n19825), .ZN(
        n19512) );
  AOI22_X1 U22472 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19516), .B1(
        n19546), .B2(n19827), .ZN(n19511) );
  OAI211_X1 U22473 ( .C1(n19830), .C2(n19519), .A(n19512), .B(n19511), .ZN(
        P2_U3109) );
  AOI22_X1 U22474 ( .A1(n19515), .A2(n19832), .B1(n19530), .B2(n19831), .ZN(
        n19514) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19516), .B1(
        n19546), .B2(n19833), .ZN(n19513) );
  OAI211_X1 U22476 ( .C1(n19836), .C2(n19519), .A(n19514), .B(n19513), .ZN(
        P2_U3110) );
  AOI22_X1 U22477 ( .A1(n19515), .A2(n19839), .B1(n19530), .B2(n19838), .ZN(
        n19518) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19516), .B1(
        n19546), .B2(n19841), .ZN(n19517) );
  OAI211_X1 U22479 ( .C1(n19847), .C2(n19519), .A(n19518), .B(n19517), .ZN(
        P2_U3111) );
  INV_X1 U22480 ( .A(n19744), .ZN(n19523) );
  NAND2_X1 U22481 ( .A1(n19968), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19619) );
  NOR2_X1 U22482 ( .A1(n19619), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19563) );
  INV_X1 U22483 ( .A(n19563), .ZN(n19565) );
  NOR2_X1 U22484 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19565), .ZN(
        n19549) );
  INV_X1 U22485 ( .A(n19549), .ZN(n19552) );
  OAI22_X1 U22486 ( .A1(n19589), .A2(n19718), .B1(n19622), .B2(n19552), .ZN(
        n19524) );
  INV_X1 U22487 ( .A(n19524), .ZN(n19534) );
  NAND2_X1 U22488 ( .A1(n19589), .A2(n19558), .ZN(n19525) );
  AOI21_X1 U22489 ( .B1(n19525), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19953), 
        .ZN(n19529) );
  OAI21_X1 U22490 ( .B1(n12379), .B2(n19851), .A(n19979), .ZN(n19526) );
  AOI21_X1 U22491 ( .B1(n19529), .B2(n19527), .A(n19526), .ZN(n19528) );
  OAI21_X1 U22492 ( .B1(n19530), .B2(n19549), .A(n19529), .ZN(n19532) );
  OAI21_X1 U22493 ( .B1(n12379), .B2(n19549), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19531) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19555), .B1(
        n19789), .B2(n19554), .ZN(n19533) );
  OAI211_X1 U22495 ( .C1(n19800), .C2(n19558), .A(n19534), .B(n19533), .ZN(
        P2_U3112) );
  OAI22_X1 U22496 ( .A1(n19589), .A2(n19762), .B1(n19634), .B2(n19552), .ZN(
        n19535) );
  INV_X1 U22497 ( .A(n19535), .ZN(n19537) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19802), .ZN(n19536) );
  OAI211_X1 U22499 ( .C1(n19806), .C2(n19558), .A(n19537), .B(n19536), .ZN(
        P2_U3113) );
  OAI22_X1 U22500 ( .A1(n19589), .A2(n19724), .B1(n19639), .B2(n19552), .ZN(
        n19538) );
  INV_X1 U22501 ( .A(n19538), .ZN(n19540) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19808), .ZN(n19539) );
  OAI211_X1 U22503 ( .C1(n19812), .C2(n19558), .A(n19540), .B(n19539), .ZN(
        P2_U3114) );
  AOI22_X1 U22504 ( .A1(n19546), .A2(n19725), .B1(n19813), .B2(n19549), .ZN(
        n19542) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19814), .ZN(n19541) );
  OAI211_X1 U22506 ( .C1(n19728), .C2(n19589), .A(n19542), .B(n19541), .ZN(
        P2_U3115) );
  OAI22_X1 U22507 ( .A1(n19558), .A2(n19824), .B1(n19649), .B2(n19552), .ZN(
        n19543) );
  INV_X1 U22508 ( .A(n19543), .ZN(n19545) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19820), .ZN(n19544) );
  OAI211_X1 U22510 ( .C1(n19732), .C2(n19589), .A(n19545), .B(n19544), .ZN(
        P2_U3116) );
  AOI22_X1 U22511 ( .A1(n19546), .A2(n19769), .B1(n19825), .B2(n19549), .ZN(
        n19548) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19826), .ZN(n19547) );
  OAI211_X1 U22513 ( .C1(n19772), .C2(n19589), .A(n19548), .B(n19547), .ZN(
        P2_U3117) );
  INV_X1 U22514 ( .A(n19589), .ZN(n19582) );
  AOI22_X1 U22515 ( .A1(n19582), .A2(n19833), .B1(n19831), .B2(n19549), .ZN(
        n19551) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19832), .ZN(n19550) );
  OAI211_X1 U22517 ( .C1(n19836), .C2(n19558), .A(n19551), .B(n19550), .ZN(
        P2_U3118) );
  OAI22_X1 U22518 ( .A1(n19589), .A2(n19784), .B1(n19666), .B2(n19552), .ZN(
        n19553) );
  INV_X1 U22519 ( .A(n19553), .ZN(n19557) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19555), .B1(
        n19554), .B2(n19839), .ZN(n19556) );
  OAI211_X1 U22521 ( .C1(n19847), .C2(n19558), .A(n19557), .B(n19556), .ZN(
        P2_U3119) );
  NOR2_X1 U22522 ( .A1(n19559), .A2(n19619), .ZN(n19592) );
  AOI22_X1 U22523 ( .A1(n19606), .A2(n19797), .B1(n19788), .B2(n19592), .ZN(
        n19568) );
  NAND2_X1 U22524 ( .A1(n19951), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19625) );
  OAI21_X1 U22525 ( .B1(n19625), .B2(n19560), .A(n19945), .ZN(n19566) );
  INV_X1 U22526 ( .A(n19592), .ZN(n19576) );
  OAI211_X1 U22527 ( .C1(n19561), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19576), 
        .B(n19953), .ZN(n19562) );
  OAI211_X1 U22528 ( .C1(n19566), .C2(n19563), .A(n19795), .B(n19562), .ZN(
        n19586) );
  OAI21_X1 U22529 ( .B1(n12352), .B2(n19592), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19564) );
  OAI21_X1 U22530 ( .B1(n19566), .B2(n19565), .A(n19564), .ZN(n19585) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19586), .B1(
        n19789), .B2(n19585), .ZN(n19567) );
  OAI211_X1 U22532 ( .C1(n19800), .C2(n19589), .A(n19568), .B(n19567), .ZN(
        P2_U3120) );
  AOI22_X1 U22533 ( .A1(n19606), .A2(n19803), .B1(n19801), .B2(n19592), .ZN(
        n19570) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19586), .B1(
        n19802), .B2(n19585), .ZN(n19569) );
  OAI211_X1 U22535 ( .C1(n19806), .C2(n19589), .A(n19570), .B(n19569), .ZN(
        P2_U3121) );
  AOI22_X1 U22536 ( .A1(n19606), .A2(n19809), .B1(n19807), .B2(n19592), .ZN(
        n19572) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19586), .B1(
        n19808), .B2(n19585), .ZN(n19571) );
  OAI211_X1 U22538 ( .C1(n19812), .C2(n19589), .A(n19572), .B(n19571), .ZN(
        P2_U3122) );
  OAI22_X1 U22539 ( .A1(n19589), .A2(n19818), .B1(n19644), .B2(n19576), .ZN(
        n19573) );
  INV_X1 U22540 ( .A(n19573), .ZN(n19575) );
  AOI22_X1 U22541 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19586), .B1(
        n19814), .B2(n19585), .ZN(n19574) );
  OAI211_X1 U22542 ( .C1(n19728), .C2(n19616), .A(n19575), .B(n19574), .ZN(
        P2_U3123) );
  OAI22_X1 U22543 ( .A1(n19589), .A2(n19824), .B1(n19649), .B2(n19576), .ZN(
        n19577) );
  INV_X1 U22544 ( .A(n19577), .ZN(n19579) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19586), .B1(
        n19820), .B2(n19585), .ZN(n19578) );
  OAI211_X1 U22546 ( .C1(n19732), .C2(n19616), .A(n19579), .B(n19578), .ZN(
        P2_U3124) );
  AOI22_X1 U22547 ( .A1(n19606), .A2(n19827), .B1(n19825), .B2(n19592), .ZN(
        n19581) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19586), .B1(
        n19826), .B2(n19585), .ZN(n19580) );
  OAI211_X1 U22549 ( .C1(n19830), .C2(n19589), .A(n19581), .B(n19580), .ZN(
        P2_U3125) );
  AOI22_X1 U22550 ( .A1(n19582), .A2(n19735), .B1(n19831), .B2(n19592), .ZN(
        n19584) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19586), .B1(
        n19832), .B2(n19585), .ZN(n19583) );
  OAI211_X1 U22552 ( .C1(n19738), .C2(n19616), .A(n19584), .B(n19583), .ZN(
        P2_U3126) );
  AOI22_X1 U22553 ( .A1(n19606), .A2(n19841), .B1(n19838), .B2(n19592), .ZN(
        n19588) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19586), .B1(
        n19839), .B2(n19585), .ZN(n19587) );
  OAI211_X1 U22555 ( .C1(n19847), .C2(n19589), .A(n19588), .B(n19587), .ZN(
        P2_U3127) );
  NOR3_X2 U22556 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19978), .A3(
        n19619), .ZN(n19611) );
  OAI21_X1 U22557 ( .B1(n12377), .B2(n19611), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19590) );
  OAI21_X1 U22558 ( .B1(n19619), .B2(n19591), .A(n19590), .ZN(n19612) );
  AOI22_X1 U22559 ( .A1(n19612), .A2(n19789), .B1(n19788), .B2(n19611), .ZN(
        n19597) );
  INV_X1 U22560 ( .A(n12377), .ZN(n19594) );
  AOI221_X1 U22561 ( .B1(n19670), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19606), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19592), .ZN(n19593) );
  AOI211_X1 U22562 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19594), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19593), .ZN(n19595) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19613), .B1(
        n19670), .B2(n19797), .ZN(n19596) );
  OAI211_X1 U22564 ( .C1(n19800), .C2(n19616), .A(n19597), .B(n19596), .ZN(
        P2_U3128) );
  AOI22_X1 U22565 ( .A1(n19612), .A2(n19802), .B1(n19801), .B2(n19611), .ZN(
        n19599) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19613), .B1(
        n19670), .B2(n19803), .ZN(n19598) );
  OAI211_X1 U22567 ( .C1(n19806), .C2(n19616), .A(n19599), .B(n19598), .ZN(
        P2_U3129) );
  AOI22_X1 U22568 ( .A1(n19612), .A2(n19808), .B1(n19807), .B2(n19611), .ZN(
        n19601) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19613), .B1(
        n19670), .B2(n19809), .ZN(n19600) );
  OAI211_X1 U22570 ( .C1(n19812), .C2(n19616), .A(n19601), .B(n19600), .ZN(
        P2_U3130) );
  AOI22_X1 U22571 ( .A1(n19612), .A2(n19814), .B1(n19813), .B2(n19611), .ZN(
        n19603) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19613), .B1(
        n19606), .B2(n19725), .ZN(n19602) );
  OAI211_X1 U22573 ( .C1(n19728), .C2(n19664), .A(n19603), .B(n19602), .ZN(
        P2_U3131) );
  AOI22_X1 U22574 ( .A1(n19612), .A2(n19820), .B1(n19819), .B2(n19611), .ZN(
        n19605) );
  AOI22_X1 U22575 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19613), .B1(
        n19606), .B2(n19729), .ZN(n19604) );
  OAI211_X1 U22576 ( .C1(n19732), .C2(n19664), .A(n19605), .B(n19604), .ZN(
        P2_U3132) );
  AOI22_X1 U22577 ( .A1(n19612), .A2(n19826), .B1(n19825), .B2(n19611), .ZN(
        n19608) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19613), .B1(
        n19606), .B2(n19769), .ZN(n19607) );
  OAI211_X1 U22579 ( .C1(n19772), .C2(n19664), .A(n19608), .B(n19607), .ZN(
        P2_U3133) );
  AOI22_X1 U22580 ( .A1(n19612), .A2(n19832), .B1(n19831), .B2(n19611), .ZN(
        n19610) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19613), .B1(
        n19670), .B2(n19833), .ZN(n19609) );
  OAI211_X1 U22582 ( .C1(n19836), .C2(n19616), .A(n19610), .B(n19609), .ZN(
        P2_U3134) );
  AOI22_X1 U22583 ( .A1(n19612), .A2(n19839), .B1(n19838), .B2(n19611), .ZN(
        n19615) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19613), .B1(
        n19670), .B2(n19841), .ZN(n19614) );
  OAI211_X1 U22585 ( .C1(n19847), .C2(n19616), .A(n19615), .B(n19614), .ZN(
        P2_U3135) );
  NOR2_X1 U22586 ( .A1(n19617), .A2(n19619), .ZN(n19631) );
  OR2_X1 U22587 ( .A1(n19631), .A2(n19851), .ZN(n19618) );
  NOR2_X1 U22588 ( .A1(n12386), .A2(n19618), .ZN(n19627) );
  OR2_X1 U22589 ( .A1(n19978), .A2(n19619), .ZN(n19628) );
  INV_X1 U22590 ( .A(n19628), .ZN(n19620) );
  AOI21_X1 U22591 ( .B1(n19979), .B2(n19620), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19621) );
  INV_X1 U22592 ( .A(n19789), .ZN(n19623) );
  INV_X1 U22593 ( .A(n19631), .ZN(n19665) );
  OAI22_X1 U22594 ( .A1(n19668), .A2(n19623), .B1(n19622), .B2(n19665), .ZN(
        n19624) );
  INV_X1 U22595 ( .A(n19624), .ZN(n19633) );
  INV_X1 U22596 ( .A(n19625), .ZN(n19791) );
  INV_X1 U22597 ( .A(n19946), .ZN(n19626) );
  NAND2_X1 U22598 ( .A1(n19791), .A2(n19626), .ZN(n19629) );
  AOI21_X1 U22599 ( .B1(n19629), .B2(n19628), .A(n19627), .ZN(n19630) );
  OAI211_X1 U22600 ( .C1(n19631), .C2(n19979), .A(n19630), .B(n19795), .ZN(
        n19671) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19715), .ZN(n19632) );
  OAI211_X1 U22602 ( .C1(n19718), .C2(n19704), .A(n19633), .B(n19632), .ZN(
        P2_U3136) );
  INV_X1 U22603 ( .A(n19802), .ZN(n19635) );
  OAI22_X1 U22604 ( .A1(n19668), .A2(n19635), .B1(n19634), .B2(n19665), .ZN(
        n19636) );
  INV_X1 U22605 ( .A(n19636), .ZN(n19638) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19671), .B1(
        n19678), .B2(n19803), .ZN(n19637) );
  OAI211_X1 U22607 ( .C1(n19806), .C2(n19664), .A(n19638), .B(n19637), .ZN(
        P2_U3137) );
  INV_X1 U22608 ( .A(n19808), .ZN(n19640) );
  OAI22_X1 U22609 ( .A1(n19668), .A2(n19640), .B1(n19639), .B2(n19665), .ZN(
        n19641) );
  INV_X1 U22610 ( .A(n19641), .ZN(n19643) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19671), .B1(
        n19678), .B2(n19809), .ZN(n19642) );
  OAI211_X1 U22612 ( .C1(n19812), .C2(n19664), .A(n19643), .B(n19642), .ZN(
        P2_U3138) );
  INV_X1 U22613 ( .A(n19814), .ZN(n19645) );
  OAI22_X1 U22614 ( .A1(n19668), .A2(n19645), .B1(n19644), .B2(n19665), .ZN(
        n19646) );
  INV_X1 U22615 ( .A(n19646), .ZN(n19648) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19725), .ZN(n19647) );
  OAI211_X1 U22617 ( .C1(n19728), .C2(n19704), .A(n19648), .B(n19647), .ZN(
        P2_U3139) );
  INV_X1 U22618 ( .A(n19820), .ZN(n19650) );
  OAI22_X1 U22619 ( .A1(n19668), .A2(n19650), .B1(n19649), .B2(n19665), .ZN(
        n19651) );
  INV_X1 U22620 ( .A(n19651), .ZN(n19653) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19729), .ZN(n19652) );
  OAI211_X1 U22622 ( .C1(n19732), .C2(n19704), .A(n19653), .B(n19652), .ZN(
        P2_U3140) );
  INV_X1 U22623 ( .A(n19826), .ZN(n19655) );
  INV_X1 U22624 ( .A(n19825), .ZN(n19654) );
  OAI22_X1 U22625 ( .A1(n19668), .A2(n19655), .B1(n19654), .B2(n19665), .ZN(
        n19656) );
  INV_X1 U22626 ( .A(n19656), .ZN(n19658) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19671), .B1(
        n19678), .B2(n19827), .ZN(n19657) );
  OAI211_X1 U22628 ( .C1(n19830), .C2(n19664), .A(n19658), .B(n19657), .ZN(
        P2_U3141) );
  INV_X1 U22629 ( .A(n19832), .ZN(n19660) );
  INV_X1 U22630 ( .A(n19831), .ZN(n19659) );
  OAI22_X1 U22631 ( .A1(n19668), .A2(n19660), .B1(n19659), .B2(n19665), .ZN(
        n19661) );
  INV_X1 U22632 ( .A(n19661), .ZN(n19663) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19671), .B1(
        n19678), .B2(n19833), .ZN(n19662) );
  OAI211_X1 U22634 ( .C1(n19836), .C2(n19664), .A(n19663), .B(n19662), .ZN(
        P2_U3142) );
  INV_X1 U22635 ( .A(n19839), .ZN(n19667) );
  OAI22_X1 U22636 ( .A1(n19668), .A2(n19667), .B1(n19666), .B2(n19665), .ZN(
        n19669) );
  INV_X1 U22637 ( .A(n19669), .ZN(n19673) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19671), .B1(
        n19670), .B2(n19778), .ZN(n19672) );
  OAI211_X1 U22639 ( .C1(n19784), .C2(n19704), .A(n19673), .B(n19672), .ZN(
        P2_U3143) );
  INV_X1 U22640 ( .A(n19674), .ZN(n19677) );
  NAND3_X1 U22641 ( .A1(n19978), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19712) );
  NOR2_X1 U22642 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19712), .ZN(
        n19699) );
  OAI21_X1 U22643 ( .B1(n19675), .B2(n19699), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19676) );
  OAI21_X1 U22644 ( .B1(n19677), .B2(n19680), .A(n19676), .ZN(n19700) );
  AOI22_X1 U22645 ( .A1(n19700), .A2(n19789), .B1(n19788), .B2(n19699), .ZN(
        n19686) );
  OAI21_X1 U22646 ( .B1(n19678), .B2(n19740), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19679) );
  OAI21_X1 U22647 ( .B1(n19680), .B2(n19960), .A(n19679), .ZN(n19684) );
  INV_X1 U22648 ( .A(n19699), .ZN(n19681) );
  OAI211_X1 U22649 ( .C1(n19682), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19681), 
        .B(n19953), .ZN(n19683) );
  NAND3_X1 U22650 ( .A1(n19684), .A2(n19795), .A3(n19683), .ZN(n19701) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19701), .B1(
        n19740), .B2(n19797), .ZN(n19685) );
  OAI211_X1 U22652 ( .C1(n19800), .C2(n19704), .A(n19686), .B(n19685), .ZN(
        P2_U3144) );
  AOI22_X1 U22653 ( .A1(n19700), .A2(n19802), .B1(n19801), .B2(n19699), .ZN(
        n19688) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19701), .B1(
        n19740), .B2(n19803), .ZN(n19687) );
  OAI211_X1 U22655 ( .C1(n19806), .C2(n19704), .A(n19688), .B(n19687), .ZN(
        P2_U3145) );
  AOI22_X1 U22656 ( .A1(n19700), .A2(n19808), .B1(n19807), .B2(n19699), .ZN(
        n19690) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19701), .B1(
        n19740), .B2(n19809), .ZN(n19689) );
  OAI211_X1 U22658 ( .C1(n19812), .C2(n19704), .A(n19690), .B(n19689), .ZN(
        P2_U3146) );
  AOI22_X1 U22659 ( .A1(n19700), .A2(n19814), .B1(n19813), .B2(n19699), .ZN(
        n19692) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19701), .B1(
        n19740), .B2(n19815), .ZN(n19691) );
  OAI211_X1 U22661 ( .C1(n19818), .C2(n19704), .A(n19692), .B(n19691), .ZN(
        P2_U3147) );
  AOI22_X1 U22662 ( .A1(n19700), .A2(n19820), .B1(n19819), .B2(n19699), .ZN(
        n19694) );
  AOI22_X1 U22663 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19701), .B1(
        n19740), .B2(n19821), .ZN(n19693) );
  OAI211_X1 U22664 ( .C1(n19824), .C2(n19704), .A(n19694), .B(n19693), .ZN(
        P2_U3148) );
  AOI22_X1 U22665 ( .A1(n19700), .A2(n19826), .B1(n19825), .B2(n19699), .ZN(
        n19696) );
  AOI22_X1 U22666 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19701), .B1(
        n19740), .B2(n19827), .ZN(n19695) );
  OAI211_X1 U22667 ( .C1(n19830), .C2(n19704), .A(n19696), .B(n19695), .ZN(
        P2_U3149) );
  AOI22_X1 U22668 ( .A1(n19700), .A2(n19832), .B1(n19831), .B2(n19699), .ZN(
        n19698) );
  AOI22_X1 U22669 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19701), .B1(
        n19740), .B2(n19833), .ZN(n19697) );
  OAI211_X1 U22670 ( .C1(n19836), .C2(n19704), .A(n19698), .B(n19697), .ZN(
        P2_U3150) );
  AOI22_X1 U22671 ( .A1(n19700), .A2(n19839), .B1(n19838), .B2(n19699), .ZN(
        n19703) );
  AOI22_X1 U22672 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19701), .B1(
        n19740), .B2(n19841), .ZN(n19702) );
  OAI211_X1 U22673 ( .C1(n19847), .C2(n19704), .A(n19703), .B(n19702), .ZN(
        P2_U3151) );
  NOR2_X1 U22674 ( .A1(n19987), .A2(n19712), .ZN(n19749) );
  NOR3_X1 U22675 ( .A1(n19706), .A2(n19749), .A3(n19851), .ZN(n19711) );
  INV_X1 U22676 ( .A(n19712), .ZN(n19707) );
  AOI21_X1 U22677 ( .B1(n19979), .B2(n19707), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19708) );
  NOR2_X1 U22678 ( .A1(n19711), .A2(n19708), .ZN(n19739) );
  AOI22_X1 U22679 ( .A1(n19739), .A2(n19789), .B1(n19788), .B2(n19749), .ZN(
        n19717) );
  INV_X1 U22680 ( .A(n19709), .ZN(n19710) );
  NAND2_X1 U22681 ( .A1(n19791), .A2(n19710), .ZN(n19713) );
  AOI21_X1 U22682 ( .B1(n19713), .B2(n19712), .A(n19711), .ZN(n19714) );
  OAI211_X1 U22683 ( .C1(n19749), .C2(n19979), .A(n19714), .B(n19795), .ZN(
        n19741) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19715), .ZN(n19716) );
  OAI211_X1 U22685 ( .C1(n19718), .C2(n19776), .A(n19717), .B(n19716), .ZN(
        P2_U3152) );
  AOI22_X1 U22686 ( .A1(n19739), .A2(n19802), .B1(n19801), .B2(n19749), .ZN(
        n19720) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19759), .ZN(n19719) );
  OAI211_X1 U22688 ( .C1(n19762), .C2(n19776), .A(n19720), .B(n19719), .ZN(
        P2_U3153) );
  AOI22_X1 U22689 ( .A1(n19739), .A2(n19808), .B1(n19807), .B2(n19749), .ZN(
        n19723) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19721), .ZN(n19722) );
  OAI211_X1 U22691 ( .C1(n19724), .C2(n19776), .A(n19723), .B(n19722), .ZN(
        P2_U3154) );
  AOI22_X1 U22692 ( .A1(n19739), .A2(n19814), .B1(n19813), .B2(n19749), .ZN(
        n19727) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19725), .ZN(n19726) );
  OAI211_X1 U22694 ( .C1(n19728), .C2(n19776), .A(n19727), .B(n19726), .ZN(
        P2_U3155) );
  AOI22_X1 U22695 ( .A1(n19739), .A2(n19820), .B1(n19819), .B2(n19749), .ZN(
        n19731) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19729), .ZN(n19730) );
  OAI211_X1 U22697 ( .C1(n19732), .C2(n19776), .A(n19731), .B(n19730), .ZN(
        P2_U3156) );
  AOI22_X1 U22698 ( .A1(n19739), .A2(n19826), .B1(n19825), .B2(n19749), .ZN(
        n19734) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19769), .ZN(n19733) );
  OAI211_X1 U22700 ( .C1(n19772), .C2(n19776), .A(n19734), .B(n19733), .ZN(
        P2_U3157) );
  AOI22_X1 U22701 ( .A1(n19739), .A2(n19832), .B1(n19831), .B2(n19749), .ZN(
        n19737) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19735), .ZN(n19736) );
  OAI211_X1 U22703 ( .C1(n19738), .C2(n19776), .A(n19737), .B(n19736), .ZN(
        P2_U3158) );
  AOI22_X1 U22704 ( .A1(n19739), .A2(n19839), .B1(n19838), .B2(n19749), .ZN(
        n19743) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19778), .ZN(n19742) );
  OAI211_X1 U22706 ( .C1(n19784), .C2(n19776), .A(n19743), .B(n19742), .ZN(
        P2_U3159) );
  NAND2_X1 U22707 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19745), .ZN(
        n19793) );
  NOR2_X1 U22708 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19793), .ZN(
        n19777) );
  AOI22_X1 U22709 ( .A1(n19773), .A2(n19797), .B1(n19788), .B2(n19777), .ZN(
        n19758) );
  AOI21_X1 U22710 ( .B1(n19746), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19751) );
  NAND2_X1 U22711 ( .A1(n19846), .A2(n19945), .ZN(n19748) );
  INV_X1 U22712 ( .A(n19948), .ZN(n19747) );
  OAI21_X1 U22713 ( .B1(n19748), .B2(n19779), .A(n19747), .ZN(n19752) );
  NOR2_X1 U22714 ( .A1(n19777), .A2(n19749), .ZN(n19755) );
  NAND2_X1 U22715 ( .A1(n19752), .A2(n19755), .ZN(n19750) );
  OAI211_X1 U22716 ( .C1(n19777), .C2(n19751), .A(n19750), .B(n19795), .ZN(
        n19781) );
  INV_X1 U22717 ( .A(n19752), .ZN(n19756) );
  OAI21_X1 U22718 ( .B1(n19753), .B2(n19777), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19754) );
  AOI22_X1 U22719 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19781), .B1(
        n19789), .B2(n19780), .ZN(n19757) );
  OAI211_X1 U22720 ( .C1(n19800), .C2(n19776), .A(n19758), .B(n19757), .ZN(
        P2_U3160) );
  AOI22_X1 U22721 ( .A1(n19779), .A2(n19759), .B1(n19801), .B2(n19777), .ZN(
        n19761) );
  AOI22_X1 U22722 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19781), .B1(
        n19802), .B2(n19780), .ZN(n19760) );
  OAI211_X1 U22723 ( .C1(n19762), .C2(n19846), .A(n19761), .B(n19760), .ZN(
        P2_U3161) );
  AOI22_X1 U22724 ( .A1(n19773), .A2(n19809), .B1(n19807), .B2(n19777), .ZN(
        n19764) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19781), .B1(
        n19808), .B2(n19780), .ZN(n19763) );
  OAI211_X1 U22726 ( .C1(n19812), .C2(n19776), .A(n19764), .B(n19763), .ZN(
        P2_U3162) );
  AOI22_X1 U22727 ( .A1(n19773), .A2(n19815), .B1(n19813), .B2(n19777), .ZN(
        n19766) );
  AOI22_X1 U22728 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19781), .B1(
        n19814), .B2(n19780), .ZN(n19765) );
  OAI211_X1 U22729 ( .C1(n19818), .C2(n19776), .A(n19766), .B(n19765), .ZN(
        P2_U3163) );
  AOI22_X1 U22730 ( .A1(n19773), .A2(n19821), .B1(n19819), .B2(n19777), .ZN(
        n19768) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19781), .B1(
        n19820), .B2(n19780), .ZN(n19767) );
  OAI211_X1 U22732 ( .C1(n19824), .C2(n19776), .A(n19768), .B(n19767), .ZN(
        P2_U3164) );
  AOI22_X1 U22733 ( .A1(n19779), .A2(n19769), .B1(n19825), .B2(n19777), .ZN(
        n19771) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19781), .B1(
        n19826), .B2(n19780), .ZN(n19770) );
  OAI211_X1 U22735 ( .C1(n19772), .C2(n19846), .A(n19771), .B(n19770), .ZN(
        P2_U3165) );
  AOI22_X1 U22736 ( .A1(n19773), .A2(n19833), .B1(n19831), .B2(n19777), .ZN(
        n19775) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19781), .B1(
        n19832), .B2(n19780), .ZN(n19774) );
  OAI211_X1 U22738 ( .C1(n19836), .C2(n19776), .A(n19775), .B(n19774), .ZN(
        P2_U3166) );
  AOI22_X1 U22739 ( .A1(n19779), .A2(n19778), .B1(n19838), .B2(n19777), .ZN(
        n19783) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19781), .B1(
        n19839), .B2(n19780), .ZN(n19782) );
  OAI211_X1 U22741 ( .C1(n19784), .C2(n19846), .A(n19783), .B(n19782), .ZN(
        P2_U3167) );
  NOR3_X1 U22742 ( .A1(n19785), .A2(n19837), .A3(n19851), .ZN(n19792) );
  INV_X1 U22743 ( .A(n19793), .ZN(n19786) );
  AOI21_X1 U22744 ( .B1(n19979), .B2(n19786), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19787) );
  NOR2_X1 U22745 ( .A1(n19792), .A2(n19787), .ZN(n19840) );
  AOI22_X1 U22746 ( .A1(n19840), .A2(n19789), .B1(n19788), .B2(n19837), .ZN(
        n19799) );
  NAND2_X1 U22747 ( .A1(n19791), .A2(n19790), .ZN(n19794) );
  AOI21_X1 U22748 ( .B1(n19794), .B2(n19793), .A(n19792), .ZN(n19796) );
  OAI211_X1 U22749 ( .C1(n19837), .C2(n19979), .A(n19796), .B(n19795), .ZN(
        n19843) );
  AOI22_X1 U22750 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19843), .B1(
        n19842), .B2(n19797), .ZN(n19798) );
  OAI211_X1 U22751 ( .C1(n19800), .C2(n19846), .A(n19799), .B(n19798), .ZN(
        P2_U3168) );
  AOI22_X1 U22752 ( .A1(n19840), .A2(n19802), .B1(n19801), .B2(n19837), .ZN(
        n19805) );
  AOI22_X1 U22753 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19843), .B1(
        n19842), .B2(n19803), .ZN(n19804) );
  OAI211_X1 U22754 ( .C1(n19806), .C2(n19846), .A(n19805), .B(n19804), .ZN(
        P2_U3169) );
  AOI22_X1 U22755 ( .A1(n19840), .A2(n19808), .B1(n19807), .B2(n19837), .ZN(
        n19811) );
  AOI22_X1 U22756 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19843), .B1(
        n19842), .B2(n19809), .ZN(n19810) );
  OAI211_X1 U22757 ( .C1(n19812), .C2(n19846), .A(n19811), .B(n19810), .ZN(
        P2_U3170) );
  AOI22_X1 U22758 ( .A1(n19840), .A2(n19814), .B1(n19813), .B2(n19837), .ZN(
        n19817) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19843), .B1(
        n19842), .B2(n19815), .ZN(n19816) );
  OAI211_X1 U22760 ( .C1(n19818), .C2(n19846), .A(n19817), .B(n19816), .ZN(
        P2_U3171) );
  AOI22_X1 U22761 ( .A1(n19840), .A2(n19820), .B1(n19819), .B2(n19837), .ZN(
        n19823) );
  AOI22_X1 U22762 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19843), .B1(
        n19842), .B2(n19821), .ZN(n19822) );
  OAI211_X1 U22763 ( .C1(n19824), .C2(n19846), .A(n19823), .B(n19822), .ZN(
        P2_U3172) );
  AOI22_X1 U22764 ( .A1(n19840), .A2(n19826), .B1(n19825), .B2(n19837), .ZN(
        n19829) );
  AOI22_X1 U22765 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19843), .B1(
        n19842), .B2(n19827), .ZN(n19828) );
  OAI211_X1 U22766 ( .C1(n19830), .C2(n19846), .A(n19829), .B(n19828), .ZN(
        P2_U3173) );
  AOI22_X1 U22767 ( .A1(n19840), .A2(n19832), .B1(n19831), .B2(n19837), .ZN(
        n19835) );
  AOI22_X1 U22768 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19843), .B1(
        n19842), .B2(n19833), .ZN(n19834) );
  OAI211_X1 U22769 ( .C1(n19836), .C2(n19846), .A(n19835), .B(n19834), .ZN(
        P2_U3174) );
  AOI22_X1 U22770 ( .A1(n19840), .A2(n19839), .B1(n19838), .B2(n19837), .ZN(
        n19845) );
  AOI22_X1 U22771 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19843), .B1(
        n19842), .B2(n19841), .ZN(n19844) );
  OAI211_X1 U22772 ( .C1(n19847), .C2(n19846), .A(n19845), .B(n19844), .ZN(
        P2_U3175) );
  AOI21_X1 U22773 ( .B1(n19869), .B2(n19850), .A(n19848), .ZN(n19856) );
  AOI211_X1 U22774 ( .C1(n19851), .C2(n19869), .A(n19850), .B(n19849), .ZN(
        n19852) );
  INV_X1 U22775 ( .A(n19852), .ZN(n19853) );
  OAI22_X1 U22776 ( .A1(n19856), .A2(n19855), .B1(n19854), .B2(n19853), .ZN(
        P2_U3177) );
  AND2_X1 U22777 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19857), .ZN(
        P2_U3179) );
  AND2_X1 U22778 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19857), .ZN(
        P2_U3180) );
  AND2_X1 U22779 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19857), .ZN(
        P2_U3181) );
  AND2_X1 U22780 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19857), .ZN(
        P2_U3182) );
  AND2_X1 U22781 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19857), .ZN(
        P2_U3183) );
  AND2_X1 U22782 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19857), .ZN(
        P2_U3184) );
  AND2_X1 U22783 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19857), .ZN(
        P2_U3185) );
  AND2_X1 U22784 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19857), .ZN(
        P2_U3186) );
  AND2_X1 U22785 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19857), .ZN(
        P2_U3187) );
  AND2_X1 U22786 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19857), .ZN(
        P2_U3188) );
  AND2_X1 U22787 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19857), .ZN(
        P2_U3189) );
  AND2_X1 U22788 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19857), .ZN(
        P2_U3190) );
  AND2_X1 U22789 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19857), .ZN(
        P2_U3191) );
  AND2_X1 U22790 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19857), .ZN(
        P2_U3192) );
  AND2_X1 U22791 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19857), .ZN(
        P2_U3193) );
  AND2_X1 U22792 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19857), .ZN(
        P2_U3194) );
  AND2_X1 U22793 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19857), .ZN(
        P2_U3195) );
  AND2_X1 U22794 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19857), .ZN(
        P2_U3196) );
  AND2_X1 U22795 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19857), .ZN(
        P2_U3197) );
  AND2_X1 U22796 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19857), .ZN(
        P2_U3198) );
  AND2_X1 U22797 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19857), .ZN(
        P2_U3199) );
  AND2_X1 U22798 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19857), .ZN(
        P2_U3200) );
  AND2_X1 U22799 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19857), .ZN(P2_U3201) );
  AND2_X1 U22800 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19857), .ZN(P2_U3202) );
  AND2_X1 U22801 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19857), .ZN(P2_U3203) );
  AND2_X1 U22802 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19857), .ZN(P2_U3204) );
  AND2_X1 U22803 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19857), .ZN(P2_U3205) );
  AND2_X1 U22804 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19857), .ZN(P2_U3206) );
  AND2_X1 U22805 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19857), .ZN(P2_U3207) );
  AND2_X1 U22806 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19857), .ZN(P2_U3208) );
  NAND2_X1 U22807 ( .A1(n19869), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19871) );
  NAND3_X1 U22808 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19871), .ZN(n19860) );
  AOI211_X1 U22809 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20988), .A(
        n19858), .B(n20000), .ZN(n19859) );
  NOR2_X1 U22810 ( .A1(n21052), .A2(n19864), .ZN(n19876) );
  AOI211_X1 U22811 ( .C1(n19877), .C2(n19860), .A(n19859), .B(n19876), .ZN(
        n19861) );
  INV_X1 U22812 ( .A(n19861), .ZN(P2_U3209) );
  INV_X1 U22813 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19862) );
  AOI21_X1 U22814 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20988), .A(n19877), 
        .ZN(n19868) );
  NOR2_X1 U22815 ( .A1(n19862), .A2(n19868), .ZN(n19865) );
  AOI21_X1 U22816 ( .B1(n19865), .B2(n19864), .A(n19863), .ZN(n19866) );
  OAI211_X1 U22817 ( .C1(n20988), .C2(n19867), .A(n19866), .B(n19871), .ZN(
        P2_U3210) );
  AOI21_X1 U22818 ( .B1(n19870), .B2(n19869), .A(n19868), .ZN(n19875) );
  OAI22_X1 U22819 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19872), .B1(NA), 
        .B2(n19871), .ZN(n19873) );
  OAI211_X1 U22820 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19873), .ZN(n19874) );
  OAI21_X1 U22821 ( .B1(n19876), .B2(n19875), .A(n19874), .ZN(P2_U3211) );
  OAI222_X1 U22822 ( .A1(n19937), .A2(n19880), .B1(n19879), .B2(n20000), .C1(
        n19878), .C2(n19933), .ZN(P2_U3212) );
  OAI222_X1 U22823 ( .A1(n19937), .A2(n19882), .B1(n19881), .B2(n20000), .C1(
        n19880), .C2(n19933), .ZN(P2_U3213) );
  INV_X1 U22824 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19884) );
  OAI222_X1 U22825 ( .A1(n19937), .A2(n19884), .B1(n19883), .B2(n20000), .C1(
        n19882), .C2(n19933), .ZN(P2_U3214) );
  OAI222_X1 U22826 ( .A1(n19937), .A2(n14180), .B1(n19885), .B2(n20000), .C1(
        n19884), .C2(n19933), .ZN(P2_U3215) );
  OAI222_X1 U22827 ( .A1(n19937), .A2(n19887), .B1(n19886), .B2(n20000), .C1(
        n14180), .C2(n19933), .ZN(P2_U3216) );
  OAI222_X1 U22828 ( .A1(n19937), .A2(n19889), .B1(n19888), .B2(n20000), .C1(
        n19887), .C2(n19933), .ZN(P2_U3217) );
  INV_X1 U22829 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19891) );
  OAI222_X1 U22830 ( .A1(n19937), .A2(n19891), .B1(n19890), .B2(n20000), .C1(
        n19889), .C2(n19933), .ZN(P2_U3218) );
  OAI222_X1 U22831 ( .A1(n19937), .A2(n19893), .B1(n19892), .B2(n20000), .C1(
        n19891), .C2(n19933), .ZN(P2_U3219) );
  OAI222_X1 U22832 ( .A1(n19937), .A2(n19895), .B1(n19894), .B2(n20000), .C1(
        n19893), .C2(n19933), .ZN(P2_U3220) );
  OAI222_X1 U22833 ( .A1(n19937), .A2(n10504), .B1(n19896), .B2(n20000), .C1(
        n19895), .C2(n19933), .ZN(P2_U3221) );
  INV_X1 U22834 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19898) );
  OAI222_X1 U22835 ( .A1(n19937), .A2(n19898), .B1(n19897), .B2(n20000), .C1(
        n10504), .C2(n19933), .ZN(P2_U3222) );
  INV_X1 U22836 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19900) );
  OAI222_X1 U22837 ( .A1(n19937), .A2(n19900), .B1(n19899), .B2(n20000), .C1(
        n19898), .C2(n19933), .ZN(P2_U3223) );
  OAI222_X1 U22838 ( .A1(n19937), .A2(n19902), .B1(n19901), .B2(n20000), .C1(
        n19900), .C2(n19933), .ZN(P2_U3224) );
  OAI222_X1 U22839 ( .A1(n19937), .A2(n19904), .B1(n19903), .B2(n20000), .C1(
        n19902), .C2(n19933), .ZN(P2_U3225) );
  INV_X1 U22840 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19906) );
  OAI222_X1 U22841 ( .A1(n19937), .A2(n19906), .B1(n19905), .B2(n20000), .C1(
        n19904), .C2(n19933), .ZN(P2_U3226) );
  OAI222_X1 U22842 ( .A1(n19937), .A2(n19908), .B1(n19907), .B2(n20000), .C1(
        n19906), .C2(n19933), .ZN(P2_U3227) );
  INV_X1 U22843 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19910) );
  OAI222_X1 U22844 ( .A1(n19937), .A2(n19910), .B1(n19909), .B2(n20000), .C1(
        n19908), .C2(n19933), .ZN(P2_U3228) );
  OAI222_X1 U22845 ( .A1(n19937), .A2(n19912), .B1(n19911), .B2(n20000), .C1(
        n19910), .C2(n19933), .ZN(P2_U3229) );
  OAI222_X1 U22846 ( .A1(n19937), .A2(n15199), .B1(n19913), .B2(n20000), .C1(
        n19912), .C2(n19933), .ZN(P2_U3230) );
  OAI222_X1 U22847 ( .A1(n19937), .A2(n19915), .B1(n19914), .B2(n20000), .C1(
        n15199), .C2(n19933), .ZN(P2_U3231) );
  INV_X1 U22848 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19917) );
  OAI222_X1 U22849 ( .A1(n19937), .A2(n19917), .B1(n19916), .B2(n20000), .C1(
        n19915), .C2(n19933), .ZN(P2_U3232) );
  OAI222_X1 U22850 ( .A1(n19937), .A2(n19919), .B1(n19918), .B2(n20000), .C1(
        n19917), .C2(n19933), .ZN(P2_U3233) );
  INV_X1 U22851 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19921) );
  OAI222_X1 U22852 ( .A1(n19937), .A2(n19921), .B1(n19920), .B2(n20000), .C1(
        n19919), .C2(n19933), .ZN(P2_U3234) );
  OAI222_X1 U22853 ( .A1(n19937), .A2(n19923), .B1(n19922), .B2(n20000), .C1(
        n19921), .C2(n19933), .ZN(P2_U3235) );
  INV_X1 U22854 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19925) );
  OAI222_X1 U22855 ( .A1(n19937), .A2(n19925), .B1(n19924), .B2(n20000), .C1(
        n19923), .C2(n19933), .ZN(P2_U3236) );
  INV_X1 U22856 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19928) );
  OAI222_X1 U22857 ( .A1(n19937), .A2(n19928), .B1(n19926), .B2(n20000), .C1(
        n19925), .C2(n19933), .ZN(P2_U3237) );
  INV_X1 U22858 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19929) );
  OAI222_X1 U22859 ( .A1(n19933), .A2(n19928), .B1(n19927), .B2(n20000), .C1(
        n19929), .C2(n19937), .ZN(P2_U3238) );
  OAI222_X1 U22860 ( .A1(n19937), .A2(n19931), .B1(n19930), .B2(n20000), .C1(
        n19929), .C2(n19933), .ZN(P2_U3239) );
  INV_X1 U22861 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19934) );
  OAI222_X1 U22862 ( .A1(n19937), .A2(n19934), .B1(n19932), .B2(n20000), .C1(
        n19931), .C2(n19933), .ZN(P2_U3240) );
  INV_X1 U22863 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19936) );
  INV_X1 U22864 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19935) );
  OAI222_X1 U22865 ( .A1(n19937), .A2(n19936), .B1(n19935), .B2(n20000), .C1(
        n19934), .C2(n19933), .ZN(P2_U3241) );
  OAI22_X1 U22866 ( .A1(n20001), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20000), .ZN(n19938) );
  INV_X1 U22867 ( .A(n19938), .ZN(P2_U3585) );
  MUX2_X1 U22868 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20001), .Z(P2_U3586) );
  OAI22_X1 U22869 ( .A1(n20001), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20000), .ZN(n19939) );
  INV_X1 U22870 ( .A(n19939), .ZN(P2_U3587) );
  OAI22_X1 U22871 ( .A1(n20001), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20000), .ZN(n19940) );
  INV_X1 U22872 ( .A(n19940), .ZN(P2_U3588) );
  OAI21_X1 U22873 ( .B1(n19944), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19942), 
        .ZN(n19941) );
  INV_X1 U22874 ( .A(n19941), .ZN(P2_U3591) );
  OAI21_X1 U22875 ( .B1(n19944), .B2(n19943), .A(n19942), .ZN(P2_U3592) );
  NAND2_X1 U22876 ( .A1(n19945), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19973) );
  NOR2_X1 U22877 ( .A1(n19946), .A2(n19973), .ZN(n19963) );
  OR2_X1 U22878 ( .A1(n19974), .A2(n19953), .ZN(n19950) );
  NOR2_X1 U22879 ( .A1(n19948), .A2(n19947), .ZN(n19949) );
  NAND2_X1 U22880 ( .A1(n19950), .A2(n19949), .ZN(n19965) );
  OAI21_X1 U22881 ( .B1(n19963), .B2(n19965), .A(n19951), .ZN(n19956) );
  OR3_X1 U22882 ( .A1(n19954), .A2(n19953), .A3(n19952), .ZN(n19955) );
  OAI211_X1 U22883 ( .C1(n19957), .C2(n19979), .A(n19956), .B(n19955), .ZN(
        n19958) );
  INV_X1 U22884 ( .A(n19958), .ZN(n19959) );
  AOI22_X1 U22885 ( .A1(n19988), .A2(n19960), .B1(n19959), .B2(n19985), .ZN(
        P2_U3602) );
  INV_X1 U22886 ( .A(n19961), .ZN(n19966) );
  NOR2_X1 U22887 ( .A1(n19962), .A2(n19979), .ZN(n19964) );
  AOI211_X1 U22888 ( .C1(n19966), .C2(n19965), .A(n19964), .B(n19963), .ZN(
        n19967) );
  AOI22_X1 U22889 ( .A1(n19988), .A2(n19968), .B1(n19967), .B2(n19985), .ZN(
        P2_U3603) );
  INV_X1 U22890 ( .A(n19969), .ZN(n19980) );
  AND2_X1 U22891 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19970) );
  OR3_X1 U22892 ( .A1(n19971), .A2(n19980), .A3(n19970), .ZN(n19972) );
  OAI21_X1 U22893 ( .B1(n19974), .B2(n19973), .A(n19972), .ZN(n19975) );
  AOI21_X1 U22894 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19976), .A(n19975), 
        .ZN(n19977) );
  AOI22_X1 U22895 ( .A1(n19988), .A2(n19978), .B1(n19977), .B2(n19985), .ZN(
        P2_U3604) );
  OAI22_X1 U22896 ( .A1(n19981), .A2(n19980), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19979), .ZN(n19982) );
  AOI21_X1 U22897 ( .B1(n19984), .B2(n19983), .A(n19982), .ZN(n19986) );
  AOI22_X1 U22898 ( .A1(n19988), .A2(n19987), .B1(n19986), .B2(n19985), .ZN(
        P2_U3605) );
  INV_X1 U22899 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19989) );
  AOI22_X1 U22900 ( .A1(n20000), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19989), 
        .B2(n20001), .ZN(P2_U3608) );
  INV_X1 U22901 ( .A(n19990), .ZN(n19999) );
  AOI22_X1 U22902 ( .A1(n19994), .A2(n19993), .B1(n19992), .B2(n19991), .ZN(
        n19995) );
  AND2_X1 U22903 ( .A1(n19996), .A2(n19995), .ZN(n19998) );
  NAND2_X1 U22904 ( .A1(n19999), .A2(P2_MORE_REG_SCAN_IN), .ZN(n19997) );
  OAI21_X1 U22905 ( .B1(n19999), .B2(n19998), .A(n19997), .ZN(P2_U3609) );
  OAI22_X1 U22906 ( .A1(n20001), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20000), .ZN(n20002) );
  INV_X1 U22907 ( .A(n20002), .ZN(P2_U3611) );
  INV_X1 U22908 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20990) );
  NAND2_X1 U22909 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20749), .ZN(n20004) );
  AOI21_X1 U22910 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20004), .A(n20830), 
        .ZN(n20795) );
  INV_X1 U22911 ( .A(n20795), .ZN(n20791) );
  OAI21_X1 U22912 ( .B1(n20830), .B2(n20990), .A(n20791), .ZN(P1_U2802) );
  OAI21_X1 U22913 ( .B1(n20006), .B2(n20005), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20007) );
  OAI21_X1 U22914 ( .B1(n20008), .B2(n20169), .A(n20007), .ZN(P1_U2803) );
  INV_X2 U22915 ( .A(n20830), .ZN(n20829) );
  NOR2_X1 U22916 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20010) );
  OAI21_X1 U22917 ( .B1(n20010), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20829), .ZN(
        n20009) );
  OAI21_X1 U22918 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20829), .A(n20009), 
        .ZN(P1_U2804) );
  OAI21_X1 U22919 ( .B1(BS16), .B2(n20010), .A(n20795), .ZN(n20793) );
  OAI21_X1 U22920 ( .B1(n20795), .B2(n21140), .A(n20793), .ZN(P1_U2805) );
  AND2_X1 U22921 ( .A1(n20012), .A2(n20011), .ZN(n20812) );
  INV_X1 U22922 ( .A(n20812), .ZN(n20809) );
  AOI21_X1 U22923 ( .B1(n20809), .B2(P1_FLUSH_REG_SCAN_IN), .A(n20013), .ZN(
        n20014) );
  INV_X1 U22924 ( .A(n20014), .ZN(P1_U2806) );
  NOR4_X1 U22925 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20018) );
  NOR4_X1 U22926 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20017) );
  NOR4_X1 U22927 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20016) );
  NOR4_X1 U22928 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20015) );
  NAND4_X1 U22929 ( .A1(n20018), .A2(n20017), .A3(n20016), .A4(n20015), .ZN(
        n20024) );
  NOR4_X1 U22930 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20022) );
  AOI211_X1 U22931 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20021) );
  NOR4_X1 U22932 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20020) );
  NOR4_X1 U22933 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20019) );
  NAND4_X1 U22934 ( .A1(n20022), .A2(n20021), .A3(n20020), .A4(n20019), .ZN(
        n20023) );
  NOR2_X1 U22935 ( .A1(n20024), .A2(n20023), .ZN(n20805) );
  INV_X1 U22936 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21037) );
  INV_X1 U22937 ( .A(n20805), .ZN(n20807) );
  NOR2_X1 U22938 ( .A1(P1_DATAWIDTH_REG_1__SCAN_IN), .A2(n20807), .ZN(n20025)
         );
  INV_X1 U22939 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20792) );
  NAND3_X1 U22940 ( .A1(n20025), .A2(n14021), .A3(n20792), .ZN(n20027) );
  OAI221_X1 U22941 ( .B1(n20805), .B2(n21037), .C1(n20807), .C2(n13638), .A(
        n20027), .ZN(P1_U2807) );
  OAI21_X1 U22942 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(n20805), .ZN(n20026) );
  OAI21_X1 U22943 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n20805), .A(n20026), 
        .ZN(n20028) );
  NAND2_X1 U22944 ( .A1(n20028), .A2(n20027), .ZN(P1_U2808) );
  INV_X1 U22945 ( .A(n20029), .ZN(n20097) );
  OAI21_X1 U22946 ( .B1(n20097), .B2(n20031), .A(n20030), .ZN(n20042) );
  NOR3_X1 U22947 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20102), .A3(n20031), .ZN(
        n20032) );
  AOI211_X1 U22948 ( .C1(n20098), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20070), .B(n20032), .ZN(n20038) );
  NAND2_X1 U22949 ( .A1(n20113), .A2(n20048), .ZN(n20037) );
  INV_X1 U22950 ( .A(n20033), .ZN(n20034) );
  AOI22_X1 U22951 ( .A1(n20084), .A2(P1_EBX_REG_7__SCAN_IN), .B1(n20034), .B2(
        n20075), .ZN(n20036) );
  NAND2_X1 U22952 ( .A1(n20096), .A2(n20110), .ZN(n20035) );
  AND4_X1 U22953 ( .A1(n20038), .A2(n20037), .A3(n20036), .A4(n20035), .ZN(
        n20039) );
  OAI21_X1 U22954 ( .B1(n20040), .B2(n20042), .A(n20039), .ZN(P1_U2833) );
  INV_X1 U22955 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20940) );
  OAI22_X1 U22956 ( .A1(n20042), .A2(n20940), .B1(n20073), .B2(n20041), .ZN(
        n20043) );
  AOI211_X1 U22957 ( .C1(n20098), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20070), .B(n20043), .ZN(n20051) );
  INV_X1 U22958 ( .A(n20044), .ZN(n20049) );
  NAND4_X1 U22959 ( .A1(n20091), .A2(n20045), .A3(P1_REIP_REG_5__SCAN_IN), 
        .A4(n20940), .ZN(n20046) );
  OAI21_X1 U22960 ( .B1(n20103), .B2(n20907), .A(n20046), .ZN(n20047) );
  AOI21_X1 U22961 ( .B1(n20049), .B2(n20048), .A(n20047), .ZN(n20050) );
  OAI211_X1 U22962 ( .C1(n20052), .C2(n20109), .A(n20051), .B(n20050), .ZN(
        P1_U2834) );
  AOI21_X1 U22963 ( .B1(n20091), .B2(n20053), .A(n20097), .ZN(n20080) );
  OR3_X1 U22964 ( .A1(n20102), .A2(P1_REIP_REG_5__SCAN_IN), .A3(n20053), .ZN(
        n20060) );
  NAND2_X1 U22965 ( .A1(n20084), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n20059) );
  NAND2_X1 U22966 ( .A1(n20096), .A2(n20054), .ZN(n20058) );
  NAND2_X1 U22967 ( .A1(n20098), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n20056) );
  AND2_X1 U22968 ( .A1(n20056), .A2(n20055), .ZN(n20057) );
  AND4_X1 U22969 ( .A1(n20060), .A2(n20059), .A3(n20058), .A4(n20057), .ZN(
        n20063) );
  NAND2_X1 U22970 ( .A1(n20061), .A2(n20106), .ZN(n20062) );
  OAI211_X1 U22971 ( .C1(n20080), .C2(n20984), .A(n20063), .B(n20062), .ZN(
        n20064) );
  INV_X1 U22972 ( .A(n20064), .ZN(n20065) );
  OAI21_X1 U22973 ( .B1(n20066), .B2(n20109), .A(n20065), .ZN(P1_U2835) );
  AOI21_X1 U22974 ( .B1(n20091), .B2(n20067), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n20081) );
  NOR2_X1 U22975 ( .A1(n20101), .A2(n20068), .ZN(n20069) );
  AOI211_X1 U22976 ( .C1(n20098), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20070), .B(n20069), .ZN(n20071) );
  OAI21_X1 U22977 ( .B1(n20073), .B2(n20072), .A(n20071), .ZN(n20074) );
  AOI21_X1 U22978 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n20084), .A(n20074), .ZN(
        n20079) );
  AOI22_X1 U22979 ( .A1(n20077), .A2(n20106), .B1(n20076), .B2(n20075), .ZN(
        n20078) );
  OAI211_X1 U22980 ( .C1(n20081), .C2(n20080), .A(n20079), .B(n20078), .ZN(
        P1_U2836) );
  INV_X1 U22981 ( .A(n20101), .ZN(n20082) );
  INV_X1 U22982 ( .A(n13382), .ZN(n20161) );
  AOI22_X1 U22983 ( .A1(n20082), .A2(n20161), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20098), .ZN(n20089) );
  NAND2_X1 U22984 ( .A1(n20083), .A2(n20106), .ZN(n20088) );
  NAND2_X1 U22985 ( .A1(n20084), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n20087) );
  NAND2_X1 U22986 ( .A1(n20096), .A2(n20085), .ZN(n20086) );
  AND4_X1 U22987 ( .A1(n20089), .A2(n20088), .A3(n20087), .A4(n20086), .ZN(
        n20093) );
  OAI221_X1 U22988 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_REIP_REG_2__SCAN_IN), .C2(n20091), .A(n20090), .ZN(n20092) );
  OAI211_X1 U22989 ( .C1(n20109), .C2(n20094), .A(n20093), .B(n20092), .ZN(
        P1_U2838) );
  NAND2_X1 U22990 ( .A1(n20096), .A2(n20095), .ZN(n20100) );
  AOI22_X1 U22991 ( .A1(n20098), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20097), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20099) );
  OAI211_X1 U22992 ( .C1(n20101), .C2(n20493), .A(n20100), .B(n20099), .ZN(
        n20105) );
  OAI22_X1 U22993 ( .A1(n20103), .A2(n21056), .B1(P1_REIP_REG_1__SCAN_IN), 
        .B2(n20102), .ZN(n20104) );
  AOI211_X1 U22994 ( .C1(n20107), .C2(n20106), .A(n20105), .B(n20104), .ZN(
        n20108) );
  OAI21_X1 U22995 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20109), .A(
        n20108), .ZN(P1_U2839) );
  INV_X1 U22996 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21147) );
  AOI22_X1 U22997 ( .A1(n20113), .A2(n20112), .B1(n20111), .B2(n20110), .ZN(
        n20114) );
  OAI21_X1 U22998 ( .B1(n14492), .B2(n21147), .A(n20114), .ZN(P1_U2865) );
  AOI22_X1 U22999 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20118), .B1(n15757), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20115) );
  OAI21_X1 U23000 ( .B1(n20117), .B2(n20116), .A(n20115), .ZN(P1_U2921) );
  INV_X1 U23001 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20120) );
  AOI22_X1 U23002 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20119) );
  OAI21_X1 U23003 ( .B1(n20120), .B2(n20143), .A(n20119), .ZN(P1_U2922) );
  INV_X1 U23004 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U23005 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20121) );
  OAI21_X1 U23006 ( .B1(n20122), .B2(n20143), .A(n20121), .ZN(P1_U2923) );
  INV_X1 U23007 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20124) );
  AOI22_X1 U23008 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20123) );
  OAI21_X1 U23009 ( .B1(n20124), .B2(n20143), .A(n20123), .ZN(P1_U2924) );
  AOI22_X1 U23010 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20125) );
  OAI21_X1 U23011 ( .B1(n20126), .B2(n20143), .A(n20125), .ZN(P1_U2925) );
  INV_X1 U23012 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20128) );
  AOI22_X1 U23013 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20127) );
  OAI21_X1 U23014 ( .B1(n20128), .B2(n20143), .A(n20127), .ZN(P1_U2926) );
  INV_X1 U23015 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20130) );
  AOI22_X1 U23016 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20129) );
  OAI21_X1 U23017 ( .B1(n20130), .B2(n20143), .A(n20129), .ZN(P1_U2927) );
  AOI22_X1 U23018 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20131) );
  OAI21_X1 U23019 ( .B1(n20132), .B2(n20143), .A(n20131), .ZN(P1_U2928) );
  AOI22_X1 U23020 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20133) );
  OAI21_X1 U23021 ( .B1(n11233), .B2(n20143), .A(n20133), .ZN(P1_U2929) );
  AOI22_X1 U23022 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20134) );
  OAI21_X1 U23023 ( .B1(n11311), .B2(n20143), .A(n20134), .ZN(P1_U2930) );
  AOI22_X1 U23024 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20135) );
  OAI21_X1 U23025 ( .B1(n11300), .B2(n20143), .A(n20135), .ZN(P1_U2931) );
  AOI22_X1 U23026 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20136) );
  OAI21_X1 U23027 ( .B1(n20137), .B2(n20143), .A(n20136), .ZN(P1_U2932) );
  AOI22_X1 U23028 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20138) );
  OAI21_X1 U23029 ( .B1(n11282), .B2(n20143), .A(n20138), .ZN(P1_U2933) );
  AOI22_X1 U23030 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20139) );
  OAI21_X1 U23031 ( .B1(n11255), .B2(n20143), .A(n20139), .ZN(P1_U2934) );
  AOI22_X1 U23032 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20140) );
  OAI21_X1 U23033 ( .B1(n11261), .B2(n20143), .A(n20140), .ZN(P1_U2935) );
  AOI22_X1 U23034 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20141), .B1(n15757), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20142) );
  OAI21_X1 U23035 ( .B1(n11271), .B2(n20143), .A(n20142), .ZN(P1_U2936) );
  AOI22_X1 U23036 ( .A1(n20153), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20152), .ZN(n20145) );
  NAND2_X1 U23037 ( .A1(n20145), .A2(n20144), .ZN(P1_U2961) );
  AOI22_X1 U23038 ( .A1(n20153), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20152), .ZN(n20147) );
  NAND2_X1 U23039 ( .A1(n20147), .A2(n20146), .ZN(P1_U2962) );
  AOI22_X1 U23040 ( .A1(n20153), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20152), .ZN(n20149) );
  NAND2_X1 U23041 ( .A1(n20149), .A2(n20148), .ZN(P1_U2964) );
  AOI22_X1 U23042 ( .A1(n20153), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20152), .ZN(n20151) );
  NAND2_X1 U23043 ( .A1(n20151), .A2(n20150), .ZN(P1_U2965) );
  AOI22_X1 U23044 ( .A1(n20153), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20152), .ZN(n20155) );
  NAND2_X1 U23045 ( .A1(n20155), .A2(n20154), .ZN(P1_U2966) );
  NOR2_X1 U23046 ( .A1(n20157), .A2(n20156), .ZN(P1_U3032) );
  INV_X1 U23047 ( .A(n20257), .ZN(n20159) );
  INV_X1 U23048 ( .A(n20730), .ZN(n20158) );
  NAND2_X1 U23049 ( .A1(n20158), .A2(n20688), .ZN(n20160) );
  OAI21_X1 U23050 ( .B1(n20160), .B2(n20253), .A(n20568), .ZN(n20176) );
  OR2_X1 U23051 ( .A1(n20436), .A2(n20161), .ZN(n20295) );
  INV_X1 U23052 ( .A(n20493), .ZN(n20639) );
  NOR2_X1 U23053 ( .A1(n20295), .A2(n20639), .ZN(n20173) );
  NOR2_X1 U23054 ( .A1(n20171), .A2(n20813), .ZN(n20496) );
  INV_X1 U23055 ( .A(n20494), .ZN(n20162) );
  NOR2_X1 U23056 ( .A1(n20162), .A2(n20437), .ZN(n20327) );
  INV_X1 U23057 ( .A(n20682), .ZN(n20582) );
  INV_X1 U23058 ( .A(DATAI_24_), .ZN(n21012) );
  NOR2_X2 U23059 ( .A1(n20222), .A2(n9812), .ZN(n20681) );
  NOR3_X1 U23060 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20236) );
  NAND2_X1 U23061 ( .A1(n20610), .A2(n20236), .ZN(n20174) );
  INV_X1 U23062 ( .A(n20174), .ZN(n20223) );
  AOI22_X1 U23063 ( .A1(n20730), .A2(n20648), .B1(n20681), .B2(n20223), .ZN(
        n20180) );
  INV_X1 U23064 ( .A(n20171), .ZN(n20172) );
  NOR2_X1 U23065 ( .A1(n20172), .A2(n20813), .ZN(n20572) );
  INV_X1 U23066 ( .A(n20173), .ZN(n20175) );
  AOI22_X1 U23067 ( .A1(n20176), .A2(n20175), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20174), .ZN(n20177) );
  INV_X1 U23068 ( .A(DATAI_16_), .ZN(n21182) );
  OAI22_X1 U23069 ( .A1(n21182), .A2(n20224), .B1(n20178), .B2(n20225), .ZN(
        n20690) );
  AOI22_X1 U23070 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20227), .B1(
        n20253), .B2(n9943), .ZN(n20179) );
  OAI211_X1 U23071 ( .C1(n20230), .C2(n20582), .A(n20180), .B(n20179), .ZN(
        P1_U3033) );
  INV_X1 U23072 ( .A(DATAI_25_), .ZN(n21154) );
  OAI22_X1 U23073 ( .A1(n20182), .A2(n20225), .B1(n21154), .B2(n20224), .ZN(
        n20651) );
  NOR2_X2 U23074 ( .A1(n20222), .A2(n20183), .ZN(n20694) );
  AOI22_X1 U23075 ( .A1(n20730), .A2(n9923), .B1(n20694), .B2(n20223), .ZN(
        n20186) );
  OAI22_X1 U23076 ( .A1(n20184), .A2(n20225), .B1(n15894), .B2(n20224), .ZN(
        n20696) );
  AOI22_X1 U23077 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20227), .B1(
        n20253), .B2(n9937), .ZN(n20185) );
  OAI211_X1 U23078 ( .C1(n20230), .C2(n20585), .A(n20186), .B(n20185), .ZN(
        P1_U3034) );
  INV_X1 U23079 ( .A(n20700), .ZN(n20588) );
  INV_X1 U23080 ( .A(DATAI_26_), .ZN(n20188) );
  OAI22_X1 U23081 ( .A1(n20189), .A2(n20225), .B1(n20188), .B2(n20224), .ZN(
        n20654) );
  NOR2_X2 U23082 ( .A1(n20222), .A2(n20190), .ZN(n20699) );
  AOI22_X1 U23083 ( .A1(n20730), .A2(n9925), .B1(n20699), .B2(n20223), .ZN(
        n20193) );
  INV_X1 U23084 ( .A(DATAI_18_), .ZN(n21170) );
  OAI22_X1 U23085 ( .A1(n20191), .A2(n20225), .B1(n21170), .B2(n20224), .ZN(
        n20701) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20227), .B1(
        n20253), .B2(n9939), .ZN(n20192) );
  OAI211_X1 U23087 ( .C1(n20230), .C2(n20588), .A(n20193), .B(n20192), .ZN(
        P1_U3035) );
  INV_X1 U23088 ( .A(n20705), .ZN(n20591) );
  INV_X1 U23089 ( .A(DATAI_27_), .ZN(n21153) );
  OAI22_X1 U23090 ( .A1(n20195), .A2(n20225), .B1(n21153), .B2(n20224), .ZN(
        n20657) );
  NOR2_X2 U23091 ( .A1(n20222), .A2(n11030), .ZN(n20704) );
  AOI22_X1 U23092 ( .A1(n20730), .A2(n9945), .B1(n20704), .B2(n20223), .ZN(
        n20199) );
  INV_X1 U23093 ( .A(DATAI_19_), .ZN(n20197) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20227), .B1(
        n20253), .B2(n20706), .ZN(n20198) );
  OAI211_X1 U23095 ( .C1(n20230), .C2(n20591), .A(n20199), .B(n20198), .ZN(
        P1_U3036) );
  INV_X1 U23096 ( .A(n20710), .ZN(n20594) );
  INV_X1 U23097 ( .A(DATAI_28_), .ZN(n20861) );
  OAI22_X1 U23098 ( .A1(n20201), .A2(n20225), .B1(n20861), .B2(n20224), .ZN(
        n20661) );
  NOR2_X2 U23099 ( .A1(n20222), .A2(n20202), .ZN(n20709) );
  AOI22_X1 U23100 ( .A1(n20730), .A2(n9933), .B1(n20709), .B2(n20223), .ZN(
        n20206) );
  INV_X1 U23101 ( .A(DATAI_20_), .ZN(n20203) );
  OAI22_X1 U23102 ( .A1(n20204), .A2(n20225), .B1(n20203), .B2(n20224), .ZN(
        n20711) );
  AOI22_X1 U23103 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20227), .B1(
        n20253), .B2(n9929), .ZN(n20205) );
  OAI211_X1 U23104 ( .C1(n20230), .C2(n20594), .A(n20206), .B(n20205), .ZN(
        P1_U3037) );
  INV_X1 U23105 ( .A(n20715), .ZN(n20597) );
  INV_X1 U23106 ( .A(DATAI_29_), .ZN(n20973) );
  NOR2_X2 U23107 ( .A1(n20222), .A2(n20209), .ZN(n20714) );
  AOI22_X1 U23108 ( .A1(n20730), .A2(n20664), .B1(n20714), .B2(n20223), .ZN(
        n20212) );
  OAI22_X1 U23109 ( .A1(n15882), .A2(n20224), .B1(n20210), .B2(n20225), .ZN(
        n20716) );
  AOI22_X1 U23110 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20227), .B1(
        n20253), .B2(n9921), .ZN(n20211) );
  OAI211_X1 U23111 ( .C1(n20230), .C2(n20597), .A(n20212), .B(n20211), .ZN(
        P1_U3038) );
  INV_X1 U23112 ( .A(DATAI_30_), .ZN(n21144) );
  OAI22_X1 U23113 ( .A1(n20214), .A2(n20225), .B1(n21144), .B2(n20224), .ZN(
        n20667) );
  NOR2_X2 U23114 ( .A1(n20222), .A2(n20215), .ZN(n20720) );
  AOI22_X1 U23115 ( .A1(n20730), .A2(n9935), .B1(n20720), .B2(n20223), .ZN(
        n20218) );
  INV_X1 U23116 ( .A(DATAI_22_), .ZN(n21168) );
  OAI22_X1 U23117 ( .A1(n20216), .A2(n20225), .B1(n21168), .B2(n20224), .ZN(
        n20722) );
  AOI22_X1 U23118 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20227), .B1(
        n20253), .B2(n9931), .ZN(n20217) );
  OAI211_X1 U23119 ( .C1(n20230), .C2(n20600), .A(n20218), .B(n20217), .ZN(
        P1_U3039) );
  INV_X1 U23120 ( .A(n20728), .ZN(n20607) );
  INV_X1 U23121 ( .A(DATAI_31_), .ZN(n21011) );
  OAI22_X1 U23122 ( .A1(n21011), .A2(n20224), .B1(n20220), .B2(n20225), .ZN(
        n20672) );
  NOR2_X2 U23123 ( .A1(n20222), .A2(n20221), .ZN(n20725) );
  AOI22_X1 U23124 ( .A1(n20730), .A2(n9927), .B1(n20725), .B2(n20223), .ZN(
        n20229) );
  INV_X1 U23125 ( .A(DATAI_23_), .ZN(n21189) );
  OAI22_X1 U23126 ( .A1(n20226), .A2(n20225), .B1(n21189), .B2(n20224), .ZN(
        n20729) );
  AOI22_X1 U23127 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20227), .B1(
        n20253), .B2(n9941), .ZN(n20228) );
  OAI211_X1 U23128 ( .C1(n20230), .C2(n20607), .A(n20229), .B(n20228), .ZN(
        P1_U3040) );
  INV_X1 U23129 ( .A(n20295), .ZN(n20232) );
  INV_X1 U23130 ( .A(n20231), .ZN(n20611) );
  INV_X1 U23131 ( .A(n20236), .ZN(n20233) );
  NOR2_X1 U23132 ( .A1(n20610), .A2(n20233), .ZN(n20251) );
  AOI21_X1 U23133 ( .B1(n20232), .B2(n20611), .A(n20251), .ZN(n20234) );
  OAI22_X1 U23134 ( .A1(n20234), .A2(n20540), .B1(n20233), .B2(n20813), .ZN(
        n20252) );
  AOI22_X1 U23135 ( .A1(n20682), .A2(n20252), .B1(n20681), .B2(n20251), .ZN(
        n20238) );
  OAI211_X1 U23136 ( .C1(n20300), .C2(n21140), .A(n20688), .B(n20234), .ZN(
        n20235) );
  OAI211_X1 U23137 ( .C1(n20688), .C2(n20236), .A(n20687), .B(n20235), .ZN(
        n20254) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20648), .ZN(n20237) );
  OAI211_X1 U23139 ( .C1(n9942), .C2(n20287), .A(n20238), .B(n20237), .ZN(
        P1_U3041) );
  AOI22_X1 U23140 ( .A1(n20695), .A2(n20252), .B1(n20694), .B2(n20251), .ZN(
        n20240) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n9923), .ZN(n20239) );
  OAI211_X1 U23142 ( .C1(n9936), .C2(n20287), .A(n20240), .B(n20239), .ZN(
        P1_U3042) );
  AOI22_X1 U23143 ( .A1(n20700), .A2(n20252), .B1(n20699), .B2(n20251), .ZN(
        n20242) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n9925), .ZN(n20241) );
  OAI211_X1 U23145 ( .C1(n9938), .C2(n20287), .A(n20242), .B(n20241), .ZN(
        P1_U3043) );
  INV_X1 U23146 ( .A(n20706), .ZN(n20660) );
  AOI22_X1 U23147 ( .A1(n20705), .A2(n20252), .B1(n20704), .B2(n20251), .ZN(
        n20244) );
  AOI22_X1 U23148 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n9945), .ZN(n20243) );
  OAI211_X1 U23149 ( .C1(n20660), .C2(n20287), .A(n20244), .B(n20243), .ZN(
        P1_U3044) );
  AOI22_X1 U23150 ( .A1(n20710), .A2(n20252), .B1(n20709), .B2(n20251), .ZN(
        n20246) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n9933), .ZN(n20245) );
  OAI211_X1 U23152 ( .C1(n9928), .C2(n20287), .A(n20246), .B(n20245), .ZN(
        P1_U3045) );
  AOI22_X1 U23153 ( .A1(n20715), .A2(n20252), .B1(n20714), .B2(n20251), .ZN(
        n20248) );
  AOI22_X1 U23154 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n20664), .ZN(n20247) );
  OAI211_X1 U23155 ( .C1(n9920), .C2(n20287), .A(n20248), .B(n20247), .ZN(
        P1_U3046) );
  AOI22_X1 U23156 ( .A1(n20721), .A2(n20252), .B1(n20720), .B2(n20251), .ZN(
        n20250) );
  AOI22_X1 U23157 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n9935), .ZN(n20249) );
  OAI211_X1 U23158 ( .C1(n9930), .C2(n20287), .A(n20250), .B(n20249), .ZN(
        P1_U3047) );
  AOI22_X1 U23159 ( .A1(n20728), .A2(n20252), .B1(n20725), .B2(n20251), .ZN(
        n20256) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20254), .B1(
        n20253), .B2(n9927), .ZN(n20255) );
  OAI211_X1 U23161 ( .C1(n9940), .C2(n20287), .A(n20256), .B(n20255), .ZN(
        P1_U3048) );
  NAND2_X1 U23162 ( .A1(n20287), .A2(n20688), .ZN(n20258) );
  OAI21_X1 U23163 ( .B1(n20321), .B2(n20258), .A(n20568), .ZN(n20260) );
  NOR2_X1 U23164 ( .A1(n20295), .A2(n20493), .ZN(n20262) );
  NOR3_X1 U23165 ( .A1(n20259), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20293) );
  NAND2_X1 U23166 ( .A1(n20610), .A2(n20293), .ZN(n20285) );
  INV_X1 U23167 ( .A(n20285), .ZN(n20281) );
  AOI22_X1 U23168 ( .A1(n20321), .A2(n9943), .B1(n20681), .B2(n20281), .ZN(
        n20265) );
  INV_X1 U23169 ( .A(n20260), .ZN(n20263) );
  NOR2_X1 U23170 ( .A1(n9913), .A2(n20813), .ZN(n20384) );
  AOI21_X1 U23171 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20285), .A(n20384), 
        .ZN(n20261) );
  INV_X1 U23172 ( .A(n20287), .ZN(n20282) );
  AOI22_X1 U23173 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20289), .B1(
        n20282), .B2(n20648), .ZN(n20264) );
  OAI211_X1 U23174 ( .C1(n20292), .C2(n20582), .A(n20265), .B(n20264), .ZN(
        P1_U3049) );
  INV_X1 U23175 ( .A(n20694), .ZN(n20266) );
  OAI22_X1 U23176 ( .A1(n20287), .A2(n9922), .B1(n20266), .B2(n20285), .ZN(
        n20267) );
  INV_X1 U23177 ( .A(n20267), .ZN(n20269) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20289), .B1(
        n20321), .B2(n9937), .ZN(n20268) );
  OAI211_X1 U23179 ( .C1(n20292), .C2(n20585), .A(n20269), .B(n20268), .ZN(
        P1_U3050) );
  INV_X1 U23180 ( .A(n20699), .ZN(n20270) );
  OAI22_X1 U23181 ( .A1(n20287), .A2(n9924), .B1(n20270), .B2(n20285), .ZN(
        n20271) );
  INV_X1 U23182 ( .A(n20271), .ZN(n20273) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20289), .B1(
        n20321), .B2(n9939), .ZN(n20272) );
  OAI211_X1 U23184 ( .C1(n20292), .C2(n20588), .A(n20273), .B(n20272), .ZN(
        P1_U3051) );
  AOI22_X1 U23185 ( .A1(n20321), .A2(n20706), .B1(n20281), .B2(n20704), .ZN(
        n20275) );
  AOI22_X1 U23186 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20289), .B1(
        n20282), .B2(n9945), .ZN(n20274) );
  OAI211_X1 U23187 ( .C1(n20292), .C2(n20591), .A(n20275), .B(n20274), .ZN(
        P1_U3052) );
  AOI22_X1 U23188 ( .A1(n20321), .A2(n9929), .B1(n20709), .B2(n20281), .ZN(
        n20277) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20289), .B1(
        n20282), .B2(n9933), .ZN(n20276) );
  OAI211_X1 U23190 ( .C1(n20292), .C2(n20594), .A(n20277), .B(n20276), .ZN(
        P1_U3053) );
  INV_X1 U23191 ( .A(n20664), .ZN(n20719) );
  INV_X1 U23192 ( .A(n20714), .ZN(n20517) );
  OAI22_X1 U23193 ( .A1(n20287), .A2(n20719), .B1(n20517), .B2(n20285), .ZN(
        n20278) );
  INV_X1 U23194 ( .A(n20278), .ZN(n20280) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20289), .B1(
        n20321), .B2(n9921), .ZN(n20279) );
  OAI211_X1 U23196 ( .C1(n20292), .C2(n20597), .A(n20280), .B(n20279), .ZN(
        P1_U3054) );
  AOI22_X1 U23197 ( .A1(n20321), .A2(n9931), .B1(n20720), .B2(n20281), .ZN(
        n20284) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20289), .B1(
        n20282), .B2(n9935), .ZN(n20283) );
  OAI211_X1 U23199 ( .C1(n20292), .C2(n20600), .A(n20284), .B(n20283), .ZN(
        P1_U3055) );
  INV_X1 U23200 ( .A(n20725), .ZN(n20286) );
  OAI22_X1 U23201 ( .A1(n20287), .A2(n9926), .B1(n20286), .B2(n20285), .ZN(
        n20288) );
  INV_X1 U23202 ( .A(n20288), .ZN(n20291) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20289), .B1(
        n20321), .B2(n9941), .ZN(n20290) );
  OAI211_X1 U23204 ( .C1(n20292), .C2(n20607), .A(n20291), .B(n20290), .ZN(
        P1_U3056) );
  INV_X1 U23205 ( .A(n20293), .ZN(n20302) );
  NAND2_X1 U23206 ( .A1(n11269), .A2(n20294), .ZN(n20535) );
  OR2_X1 U23207 ( .A1(n20295), .A2(n20535), .ZN(n20297) );
  NOR2_X1 U23208 ( .A1(n20533), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20320) );
  INV_X1 U23209 ( .A(n20320), .ZN(n20296) );
  AND2_X1 U23210 ( .A1(n20297), .A2(n20296), .ZN(n20301) );
  OAI21_X1 U23211 ( .B1(n20300), .B2(n20684), .A(n20688), .ZN(n20305) );
  OAI22_X1 U23212 ( .A1(n20813), .A2(n20302), .B1(n20301), .B2(n20305), .ZN(
        n20299) );
  AOI22_X1 U23213 ( .A1(n20352), .A2(n9943), .B1(n20320), .B2(n20681), .ZN(
        n20307) );
  INV_X1 U23214 ( .A(n20301), .ZN(n20304) );
  INV_X1 U23215 ( .A(n20687), .ZN(n20539) );
  AOI21_X1 U23216 ( .B1(n20540), .B2(n20302), .A(n20539), .ZN(n20303) );
  OAI21_X1 U23217 ( .B1(n20305), .B2(n20304), .A(n20303), .ZN(n20322) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20648), .ZN(n20306) );
  OAI211_X1 U23219 ( .C1(n20325), .C2(n20582), .A(n20307), .B(n20306), .ZN(
        P1_U3057) );
  AOI22_X1 U23220 ( .A1(n20352), .A2(n9937), .B1(n20320), .B2(n20694), .ZN(
        n20309) );
  AOI22_X1 U23221 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n9923), .ZN(n20308) );
  OAI211_X1 U23222 ( .C1(n20325), .C2(n20585), .A(n20309), .B(n20308), .ZN(
        P1_U3058) );
  AOI22_X1 U23223 ( .A1(n20321), .A2(n9925), .B1(n20320), .B2(n20699), .ZN(
        n20311) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20322), .B1(
        n20352), .B2(n9939), .ZN(n20310) );
  OAI211_X1 U23225 ( .C1(n20325), .C2(n20588), .A(n20311), .B(n20310), .ZN(
        P1_U3059) );
  AOI22_X1 U23226 ( .A1(n20321), .A2(n9945), .B1(n20320), .B2(n20704), .ZN(
        n20313) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20322), .B1(
        n20352), .B2(n20706), .ZN(n20312) );
  OAI211_X1 U23228 ( .C1(n20325), .C2(n20591), .A(n20313), .B(n20312), .ZN(
        P1_U3060) );
  AOI22_X1 U23229 ( .A1(n20352), .A2(n9929), .B1(n20320), .B2(n20709), .ZN(
        n20315) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n9933), .ZN(n20314) );
  OAI211_X1 U23231 ( .C1(n20325), .C2(n20594), .A(n20315), .B(n20314), .ZN(
        P1_U3061) );
  AOI22_X1 U23232 ( .A1(n20321), .A2(n20664), .B1(n20320), .B2(n20714), .ZN(
        n20317) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20322), .B1(
        n20352), .B2(n9921), .ZN(n20316) );
  OAI211_X1 U23234 ( .C1(n20325), .C2(n20597), .A(n20317), .B(n20316), .ZN(
        P1_U3062) );
  AOI22_X1 U23235 ( .A1(n20352), .A2(n9931), .B1(n20320), .B2(n20720), .ZN(
        n20319) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n9935), .ZN(n20318) );
  OAI211_X1 U23237 ( .C1(n20325), .C2(n20600), .A(n20319), .B(n20318), .ZN(
        P1_U3063) );
  AOI22_X1 U23238 ( .A1(n20352), .A2(n9941), .B1(n20320), .B2(n20725), .ZN(
        n20324) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n9927), .ZN(n20323) );
  OAI211_X1 U23240 ( .C1(n20325), .C2(n20607), .A(n20324), .B(n20323), .ZN(
        P1_U3064) );
  INV_X1 U23241 ( .A(n20572), .ZN(n20640) );
  INV_X1 U23242 ( .A(n20327), .ZN(n20330) );
  NOR2_X1 U23243 ( .A1(n13382), .A2(n20328), .ZN(n20411) );
  NAND3_X1 U23244 ( .A1(n20411), .A2(n20688), .A3(n20493), .ZN(n20329) );
  OAI21_X1 U23245 ( .B1(n20640), .B2(n20330), .A(n20329), .ZN(n20351) );
  NOR3_X1 U23246 ( .A1(n20573), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20359) );
  INV_X1 U23247 ( .A(n20359), .ZN(n20356) );
  NOR2_X1 U23248 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20356), .ZN(
        n20350) );
  AOI22_X1 U23249 ( .A1(n20682), .A2(n20351), .B1(n20681), .B2(n20350), .ZN(
        n20337) );
  INV_X1 U23250 ( .A(n20352), .ZN(n20331) );
  AOI21_X1 U23251 ( .B1(n20331), .B2(n20379), .A(n21140), .ZN(n20332) );
  AOI21_X1 U23252 ( .B1(n20411), .B2(n20493), .A(n20332), .ZN(n20333) );
  NOR2_X1 U23253 ( .A1(n20333), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20335) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20648), .ZN(n20336) );
  OAI211_X1 U23255 ( .C1(n9942), .C2(n20379), .A(n20337), .B(n20336), .ZN(
        P1_U3065) );
  AOI22_X1 U23256 ( .A1(n20695), .A2(n20351), .B1(n20694), .B2(n20350), .ZN(
        n20339) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n9923), .ZN(n20338) );
  OAI211_X1 U23258 ( .C1(n9936), .C2(n20379), .A(n20339), .B(n20338), .ZN(
        P1_U3066) );
  AOI22_X1 U23259 ( .A1(n20700), .A2(n20351), .B1(n20699), .B2(n20350), .ZN(
        n20341) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n9925), .ZN(n20340) );
  OAI211_X1 U23261 ( .C1(n9938), .C2(n20379), .A(n20341), .B(n20340), .ZN(
        P1_U3067) );
  AOI22_X1 U23262 ( .A1(n20705), .A2(n20351), .B1(n20704), .B2(n20350), .ZN(
        n20343) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n9945), .ZN(n20342) );
  OAI211_X1 U23264 ( .C1(n20660), .C2(n20379), .A(n20343), .B(n20342), .ZN(
        P1_U3068) );
  AOI22_X1 U23265 ( .A1(n20710), .A2(n20351), .B1(n20709), .B2(n20350), .ZN(
        n20345) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n9933), .ZN(n20344) );
  OAI211_X1 U23267 ( .C1(n9928), .C2(n20379), .A(n20345), .B(n20344), .ZN(
        P1_U3069) );
  AOI22_X1 U23268 ( .A1(n20715), .A2(n20351), .B1(n20714), .B2(n20350), .ZN(
        n20347) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20664), .ZN(n20346) );
  OAI211_X1 U23270 ( .C1(n9920), .C2(n20379), .A(n20347), .B(n20346), .ZN(
        P1_U3070) );
  AOI22_X1 U23271 ( .A1(n20721), .A2(n20351), .B1(n20720), .B2(n20350), .ZN(
        n20349) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n9935), .ZN(n20348) );
  OAI211_X1 U23273 ( .C1(n9930), .C2(n20379), .A(n20349), .B(n20348), .ZN(
        P1_U3071) );
  AOI22_X1 U23274 ( .A1(n20728), .A2(n20351), .B1(n20725), .B2(n20350), .ZN(
        n20355) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n9927), .ZN(n20354) );
  OAI211_X1 U23276 ( .C1(n9940), .C2(n20379), .A(n20355), .B(n20354), .ZN(
        P1_U3072) );
  INV_X1 U23277 ( .A(n20648), .ZN(n20693) );
  NOR2_X1 U23278 ( .A1(n20610), .A2(n20356), .ZN(n20374) );
  AOI21_X1 U23279 ( .B1(n20411), .B2(n20611), .A(n20374), .ZN(n20357) );
  OAI22_X1 U23280 ( .A1(n20357), .A2(n20540), .B1(n20356), .B2(n20813), .ZN(
        n20375) );
  AOI22_X1 U23281 ( .A1(n20682), .A2(n20375), .B1(n20681), .B2(n20374), .ZN(
        n20361) );
  OAI211_X1 U23282 ( .C1(n20414), .C2(n21140), .A(n20688), .B(n20357), .ZN(
        n20358) );
  OAI211_X1 U23283 ( .C1(n20688), .C2(n20359), .A(n20687), .B(n20358), .ZN(
        n20376) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20376), .B1(
        n20403), .B2(n9943), .ZN(n20360) );
  OAI211_X1 U23285 ( .C1(n20693), .C2(n20379), .A(n20361), .B(n20360), .ZN(
        P1_U3073) );
  AOI22_X1 U23286 ( .A1(n20695), .A2(n20375), .B1(n20694), .B2(n20374), .ZN(
        n20363) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20376), .B1(
        n20403), .B2(n9937), .ZN(n20362) );
  OAI211_X1 U23288 ( .C1(n9922), .C2(n20379), .A(n20363), .B(n20362), .ZN(
        P1_U3074) );
  AOI22_X1 U23289 ( .A1(n20700), .A2(n20375), .B1(n20699), .B2(n20374), .ZN(
        n20365) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20376), .B1(
        n20403), .B2(n9939), .ZN(n20364) );
  OAI211_X1 U23291 ( .C1(n9924), .C2(n20379), .A(n20365), .B(n20364), .ZN(
        P1_U3075) );
  AOI22_X1 U23292 ( .A1(n20705), .A2(n20375), .B1(n20704), .B2(n20374), .ZN(
        n20367) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20376), .B1(
        n20403), .B2(n20706), .ZN(n20366) );
  OAI211_X1 U23294 ( .C1(n9944), .C2(n20379), .A(n20367), .B(n20366), .ZN(
        P1_U3076) );
  AOI22_X1 U23295 ( .A1(n20710), .A2(n20375), .B1(n20709), .B2(n20374), .ZN(
        n20369) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20376), .B1(
        n20403), .B2(n9929), .ZN(n20368) );
  OAI211_X1 U23297 ( .C1(n9932), .C2(n20379), .A(n20369), .B(n20368), .ZN(
        P1_U3077) );
  AOI22_X1 U23298 ( .A1(n20715), .A2(n20375), .B1(n20714), .B2(n20374), .ZN(
        n20371) );
  AOI22_X1 U23299 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20376), .B1(
        n20403), .B2(n9921), .ZN(n20370) );
  OAI211_X1 U23300 ( .C1(n20719), .C2(n20379), .A(n20371), .B(n20370), .ZN(
        P1_U3078) );
  AOI22_X1 U23301 ( .A1(n20721), .A2(n20375), .B1(n20720), .B2(n20374), .ZN(
        n20373) );
  AOI22_X1 U23302 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20376), .B1(
        n20403), .B2(n9931), .ZN(n20372) );
  OAI211_X1 U23303 ( .C1(n9934), .C2(n20379), .A(n20373), .B(n20372), .ZN(
        P1_U3079) );
  AOI22_X1 U23304 ( .A1(n20728), .A2(n20375), .B1(n20725), .B2(n20374), .ZN(
        n20378) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20376), .B1(
        n20403), .B2(n9941), .ZN(n20377) );
  OAI211_X1 U23306 ( .C1(n9926), .C2(n20379), .A(n20378), .B(n20377), .ZN(
        P1_U3080) );
  INV_X1 U23307 ( .A(n20432), .ZN(n20381) );
  NAND2_X1 U23308 ( .A1(n20381), .A2(n20688), .ZN(n20382) );
  OAI21_X1 U23309 ( .B1(n20382), .B2(n20403), .A(n20568), .ZN(n20386) );
  AND2_X1 U23310 ( .A1(n20411), .A2(n20639), .ZN(n20383) );
  NOR2_X1 U23311 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20412), .ZN(
        n20402) );
  AOI22_X1 U23312 ( .A1(n20403), .A2(n20648), .B1(n20681), .B2(n20402), .ZN(
        n20389) );
  INV_X1 U23313 ( .A(n20383), .ZN(n20385) );
  AOI21_X1 U23314 ( .B1(n20386), .B2(n20385), .A(n20384), .ZN(n20387) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20404), .B1(
        n20432), .B2(n9943), .ZN(n20388) );
  OAI211_X1 U23316 ( .C1(n20407), .C2(n20582), .A(n20389), .B(n20388), .ZN(
        P1_U3081) );
  AOI22_X1 U23317 ( .A1(n20403), .A2(n9923), .B1(n20694), .B2(n20402), .ZN(
        n20391) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20404), .B1(
        n20432), .B2(n9937), .ZN(n20390) );
  OAI211_X1 U23319 ( .C1(n20407), .C2(n20585), .A(n20391), .B(n20390), .ZN(
        P1_U3082) );
  AOI22_X1 U23320 ( .A1(n20403), .A2(n9925), .B1(n20699), .B2(n20402), .ZN(
        n20393) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20404), .B1(
        n20432), .B2(n9939), .ZN(n20392) );
  OAI211_X1 U23322 ( .C1(n20407), .C2(n20588), .A(n20393), .B(n20392), .ZN(
        P1_U3083) );
  AOI22_X1 U23323 ( .A1(n20403), .A2(n9945), .B1(n20704), .B2(n20402), .ZN(
        n20395) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20404), .B1(
        n20432), .B2(n20706), .ZN(n20394) );
  OAI211_X1 U23325 ( .C1(n20407), .C2(n20591), .A(n20395), .B(n20394), .ZN(
        P1_U3084) );
  AOI22_X1 U23326 ( .A1(n20432), .A2(n9929), .B1(n20709), .B2(n20402), .ZN(
        n20397) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20404), .B1(
        n20403), .B2(n9933), .ZN(n20396) );
  OAI211_X1 U23328 ( .C1(n20407), .C2(n20594), .A(n20397), .B(n20396), .ZN(
        P1_U3085) );
  AOI22_X1 U23329 ( .A1(n20432), .A2(n9921), .B1(n20714), .B2(n20402), .ZN(
        n20399) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20404), .B1(
        n20403), .B2(n20664), .ZN(n20398) );
  OAI211_X1 U23331 ( .C1(n20407), .C2(n20597), .A(n20399), .B(n20398), .ZN(
        P1_U3086) );
  AOI22_X1 U23332 ( .A1(n20432), .A2(n9931), .B1(n20720), .B2(n20402), .ZN(
        n20401) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20404), .B1(
        n20403), .B2(n9935), .ZN(n20400) );
  OAI211_X1 U23334 ( .C1(n20407), .C2(n20600), .A(n20401), .B(n20400), .ZN(
        P1_U3087) );
  AOI22_X1 U23335 ( .A1(n20403), .A2(n9927), .B1(n20725), .B2(n20402), .ZN(
        n20406) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20404), .B1(
        n20432), .B2(n9941), .ZN(n20405) );
  OAI211_X1 U23337 ( .C1(n20407), .C2(n20607), .A(n20406), .B(n20405), .ZN(
        P1_U3088) );
  INV_X1 U23338 ( .A(n20545), .ZN(n20408) );
  INV_X1 U23339 ( .A(n20535), .ZN(n20678) );
  INV_X1 U23340 ( .A(n20410), .ZN(n20430) );
  AOI21_X1 U23341 ( .B1(n20411), .B2(n20678), .A(n20430), .ZN(n20413) );
  OAI22_X1 U23342 ( .A1(n20413), .A2(n20540), .B1(n20412), .B2(n20813), .ZN(
        n20431) );
  AOI22_X1 U23343 ( .A1(n20682), .A2(n20431), .B1(n20430), .B2(n20681), .ZN(
        n20417) );
  OAI211_X1 U23344 ( .C1(n20414), .C2(n20684), .A(n20688), .B(n20413), .ZN(
        n20415) );
  OAI211_X1 U23345 ( .C1(n11169), .C2(n20688), .A(n20687), .B(n20415), .ZN(
        n20433) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20648), .ZN(n20416) );
  OAI211_X1 U23347 ( .C1(n9942), .C2(n20439), .A(n20417), .B(n20416), .ZN(
        P1_U3089) );
  AOI22_X1 U23348 ( .A1(n20695), .A2(n20431), .B1(n20430), .B2(n20694), .ZN(
        n20419) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n9923), .ZN(n20418) );
  OAI211_X1 U23350 ( .C1(n9936), .C2(n20439), .A(n20419), .B(n20418), .ZN(
        P1_U3090) );
  AOI22_X1 U23351 ( .A1(n20700), .A2(n20431), .B1(n20430), .B2(n20699), .ZN(
        n20421) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n9925), .ZN(n20420) );
  OAI211_X1 U23353 ( .C1(n9938), .C2(n20439), .A(n20421), .B(n20420), .ZN(
        P1_U3091) );
  AOI22_X1 U23354 ( .A1(n20705), .A2(n20431), .B1(n20430), .B2(n20704), .ZN(
        n20423) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n9945), .ZN(n20422) );
  OAI211_X1 U23356 ( .C1(n20660), .C2(n20439), .A(n20423), .B(n20422), .ZN(
        P1_U3092) );
  AOI22_X1 U23357 ( .A1(n20710), .A2(n20431), .B1(n20430), .B2(n20709), .ZN(
        n20425) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n9933), .ZN(n20424) );
  OAI211_X1 U23359 ( .C1(n9928), .C2(n20439), .A(n20425), .B(n20424), .ZN(
        P1_U3093) );
  AOI22_X1 U23360 ( .A1(n20715), .A2(n20431), .B1(n20430), .B2(n20714), .ZN(
        n20427) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n20664), .ZN(n20426) );
  OAI211_X1 U23362 ( .C1(n9920), .C2(n20439), .A(n20427), .B(n20426), .ZN(
        P1_U3094) );
  AOI22_X1 U23363 ( .A1(n20721), .A2(n20431), .B1(n20430), .B2(n20720), .ZN(
        n20429) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n9935), .ZN(n20428) );
  OAI211_X1 U23365 ( .C1(n9930), .C2(n20439), .A(n20429), .B(n20428), .ZN(
        P1_U3095) );
  AOI22_X1 U23366 ( .A1(n20728), .A2(n20431), .B1(n20430), .B2(n20725), .ZN(
        n20435) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20433), .B1(
        n20432), .B2(n9927), .ZN(n20434) );
  OAI211_X1 U23368 ( .C1(n9940), .C2(n20439), .A(n20435), .B(n20434), .ZN(
        P1_U3096) );
  NAND2_X1 U23369 ( .A1(n20436), .A2(n13382), .ZN(n20536) );
  INV_X1 U23370 ( .A(n20536), .ZN(n20464) );
  NOR3_X1 U23371 ( .A1(n15688), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20468) );
  INV_X1 U23372 ( .A(n20468), .ZN(n20465) );
  NOR2_X1 U23373 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20465), .ZN(
        n20458) );
  AOI21_X1 U23374 ( .B1(n20464), .B2(n20493), .A(n20458), .ZN(n20441) );
  INV_X1 U23375 ( .A(n20496), .ZN(n20438) );
  AND2_X1 U23376 ( .A1(n20437), .A2(n20494), .ZN(n20571) );
  INV_X1 U23377 ( .A(n20571), .ZN(n20575) );
  OAI22_X1 U23378 ( .A1(n20441), .A2(n20540), .B1(n20438), .B2(n20575), .ZN(
        n20459) );
  AOI22_X1 U23379 ( .A1(n20682), .A2(n20459), .B1(n20681), .B2(n20458), .ZN(
        n20445) );
  INV_X1 U23380 ( .A(n20489), .ZN(n20440) );
  OAI21_X1 U23381 ( .B1(n20440), .B2(n20460), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20442) );
  NAND2_X1 U23382 ( .A1(n20442), .A2(n20441), .ZN(n20443) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20648), .ZN(n20444) );
  OAI211_X1 U23384 ( .C1(n9942), .C2(n20489), .A(n20445), .B(n20444), .ZN(
        P1_U3097) );
  AOI22_X1 U23385 ( .A1(n20695), .A2(n20459), .B1(n20694), .B2(n20458), .ZN(
        n20447) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n9923), .ZN(n20446) );
  OAI211_X1 U23387 ( .C1(n9936), .C2(n20489), .A(n20447), .B(n20446), .ZN(
        P1_U3098) );
  AOI22_X1 U23388 ( .A1(n20700), .A2(n20459), .B1(n20699), .B2(n20458), .ZN(
        n20449) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n9925), .ZN(n20448) );
  OAI211_X1 U23390 ( .C1(n9938), .C2(n20489), .A(n20449), .B(n20448), .ZN(
        P1_U3099) );
  AOI22_X1 U23391 ( .A1(n20705), .A2(n20459), .B1(n20704), .B2(n20458), .ZN(
        n20451) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n9945), .ZN(n20450) );
  OAI211_X1 U23393 ( .C1(n20660), .C2(n20489), .A(n20451), .B(n20450), .ZN(
        P1_U3100) );
  AOI22_X1 U23394 ( .A1(n20710), .A2(n20459), .B1(n20709), .B2(n20458), .ZN(
        n20453) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n9933), .ZN(n20452) );
  OAI211_X1 U23396 ( .C1(n9928), .C2(n20489), .A(n20453), .B(n20452), .ZN(
        P1_U3101) );
  AOI22_X1 U23397 ( .A1(n20715), .A2(n20459), .B1(n20714), .B2(n20458), .ZN(
        n20455) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20664), .ZN(n20454) );
  OAI211_X1 U23399 ( .C1(n9920), .C2(n20489), .A(n20455), .B(n20454), .ZN(
        P1_U3102) );
  AOI22_X1 U23400 ( .A1(n20721), .A2(n20459), .B1(n20720), .B2(n20458), .ZN(
        n20457) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n9935), .ZN(n20456) );
  OAI211_X1 U23402 ( .C1(n9930), .C2(n20489), .A(n20457), .B(n20456), .ZN(
        P1_U3103) );
  AOI22_X1 U23403 ( .A1(n20728), .A2(n20459), .B1(n20725), .B2(n20458), .ZN(
        n20463) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n9927), .ZN(n20462) );
  OAI211_X1 U23405 ( .C1(n9940), .C2(n20489), .A(n20463), .B(n20462), .ZN(
        P1_U3104) );
  NOR2_X1 U23406 ( .A1(n20610), .A2(n20465), .ZN(n20484) );
  AOI21_X1 U23407 ( .B1(n20464), .B2(n20611), .A(n20484), .ZN(n20466) );
  OAI22_X1 U23408 ( .A1(n20466), .A2(n20540), .B1(n20465), .B2(n20813), .ZN(
        n20485) );
  AOI22_X1 U23409 ( .A1(n20682), .A2(n20485), .B1(n20681), .B2(n20484), .ZN(
        n20471) );
  INV_X1 U23410 ( .A(n20490), .ZN(n20546) );
  OAI211_X1 U23411 ( .C1(n20546), .C2(n21140), .A(n20688), .B(n20466), .ZN(
        n20467) );
  OAI211_X1 U23412 ( .C1(n20688), .C2(n20468), .A(n20687), .B(n20467), .ZN(
        n20486) );
  INV_X1 U23413 ( .A(n20616), .ZN(n20469) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20486), .B1(
        n20527), .B2(n9943), .ZN(n20470) );
  OAI211_X1 U23415 ( .C1(n20693), .C2(n20489), .A(n20471), .B(n20470), .ZN(
        P1_U3105) );
  AOI22_X1 U23416 ( .A1(n20695), .A2(n20485), .B1(n20694), .B2(n20484), .ZN(
        n20473) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20486), .B1(
        n20527), .B2(n9937), .ZN(n20472) );
  OAI211_X1 U23418 ( .C1(n9922), .C2(n20489), .A(n20473), .B(n20472), .ZN(
        P1_U3106) );
  AOI22_X1 U23419 ( .A1(n20700), .A2(n20485), .B1(n20699), .B2(n20484), .ZN(
        n20475) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20486), .B1(
        n20527), .B2(n9939), .ZN(n20474) );
  OAI211_X1 U23421 ( .C1(n9924), .C2(n20489), .A(n20475), .B(n20474), .ZN(
        P1_U3107) );
  AOI22_X1 U23422 ( .A1(n20705), .A2(n20485), .B1(n20704), .B2(n20484), .ZN(
        n20477) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20486), .B1(
        n20527), .B2(n20706), .ZN(n20476) );
  OAI211_X1 U23424 ( .C1(n9944), .C2(n20489), .A(n20477), .B(n20476), .ZN(
        P1_U3108) );
  AOI22_X1 U23425 ( .A1(n20710), .A2(n20485), .B1(n20709), .B2(n20484), .ZN(
        n20479) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20486), .B1(
        n20527), .B2(n9929), .ZN(n20478) );
  OAI211_X1 U23427 ( .C1(n9932), .C2(n20489), .A(n20479), .B(n20478), .ZN(
        P1_U3109) );
  AOI22_X1 U23428 ( .A1(n20715), .A2(n20485), .B1(n20714), .B2(n20484), .ZN(
        n20481) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20486), .B1(
        n20527), .B2(n9921), .ZN(n20480) );
  OAI211_X1 U23430 ( .C1(n20719), .C2(n20489), .A(n20481), .B(n20480), .ZN(
        P1_U3110) );
  AOI22_X1 U23431 ( .A1(n20721), .A2(n20485), .B1(n20720), .B2(n20484), .ZN(
        n20483) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20486), .B1(
        n20527), .B2(n9931), .ZN(n20482) );
  OAI211_X1 U23433 ( .C1(n9934), .C2(n20489), .A(n20483), .B(n20482), .ZN(
        P1_U3111) );
  AOI22_X1 U23434 ( .A1(n20728), .A2(n20485), .B1(n20725), .B2(n20484), .ZN(
        n20488) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20486), .B1(
        n20527), .B2(n9941), .ZN(n20487) );
  OAI211_X1 U23436 ( .C1(n9926), .C2(n20489), .A(n20488), .B(n20487), .ZN(
        P1_U3112) );
  INV_X1 U23437 ( .A(n20527), .ZN(n20491) );
  NAND3_X1 U23438 ( .A1(n20491), .A2(n20688), .A3(n20566), .ZN(n20492) );
  NAND2_X1 U23439 ( .A1(n20492), .A2(n20568), .ZN(n20497) );
  NOR2_X1 U23440 ( .A1(n20536), .A2(n20493), .ZN(n20501) );
  OR2_X1 U23441 ( .A1(n20494), .A2(n15688), .ZN(n20641) );
  INV_X1 U23442 ( .A(n20641), .ZN(n20495) );
  NAND3_X1 U23443 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n20573), .ZN(n20541) );
  NOR2_X1 U23444 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20541), .ZN(
        n20526) );
  AOI22_X1 U23445 ( .A1(n20527), .A2(n20648), .B1(n20681), .B2(n20526), .ZN(
        n20504) );
  INV_X1 U23446 ( .A(n20497), .ZN(n20502) );
  NAND2_X1 U23447 ( .A1(n20641), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20645) );
  OAI21_X1 U23448 ( .B1(n20579), .B2(n20526), .A(n20645), .ZN(n20498) );
  INV_X1 U23449 ( .A(n20498), .ZN(n20499) );
  OAI211_X1 U23450 ( .C1(n20502), .C2(n20501), .A(n20500), .B(n20499), .ZN(
        n20529) );
  INV_X1 U23451 ( .A(n20566), .ZN(n20528) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20529), .B1(
        n20528), .B2(n9943), .ZN(n20503) );
  OAI211_X1 U23453 ( .C1(n20532), .C2(n20582), .A(n20504), .B(n20503), .ZN(
        P1_U3113) );
  AOI22_X1 U23454 ( .A1(n20527), .A2(n9923), .B1(n20694), .B2(n20526), .ZN(
        n20506) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20529), .B1(
        n20528), .B2(n9937), .ZN(n20505) );
  OAI211_X1 U23456 ( .C1(n20532), .C2(n20585), .A(n20506), .B(n20505), .ZN(
        P1_U3114) );
  AOI22_X1 U23457 ( .A1(n20528), .A2(n9939), .B1(n20699), .B2(n20526), .ZN(
        n20508) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20529), .B1(
        n20527), .B2(n9925), .ZN(n20507) );
  OAI211_X1 U23459 ( .C1(n20532), .C2(n20588), .A(n20508), .B(n20507), .ZN(
        P1_U3115) );
  INV_X1 U23460 ( .A(n20526), .ZN(n20521) );
  INV_X1 U23461 ( .A(n20704), .ZN(n20509) );
  OAI22_X1 U23462 ( .A1(n20566), .A2(n20660), .B1(n20521), .B2(n20509), .ZN(
        n20510) );
  INV_X1 U23463 ( .A(n20510), .ZN(n20512) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20529), .B1(
        n20527), .B2(n9945), .ZN(n20511) );
  OAI211_X1 U23465 ( .C1(n20532), .C2(n20591), .A(n20512), .B(n20511), .ZN(
        P1_U3116) );
  INV_X1 U23466 ( .A(n20709), .ZN(n20513) );
  OAI22_X1 U23467 ( .A1(n20566), .A2(n9928), .B1(n20513), .B2(n20521), .ZN(
        n20514) );
  INV_X1 U23468 ( .A(n20514), .ZN(n20516) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20529), .B1(
        n20527), .B2(n9933), .ZN(n20515) );
  OAI211_X1 U23470 ( .C1(n20532), .C2(n20594), .A(n20516), .B(n20515), .ZN(
        P1_U3117) );
  OAI22_X1 U23471 ( .A1(n20566), .A2(n9920), .B1(n20517), .B2(n20521), .ZN(
        n20518) );
  INV_X1 U23472 ( .A(n20518), .ZN(n20520) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20529), .B1(
        n20527), .B2(n20664), .ZN(n20519) );
  OAI211_X1 U23474 ( .C1(n20532), .C2(n20597), .A(n20520), .B(n20519), .ZN(
        P1_U3118) );
  INV_X1 U23475 ( .A(n20720), .ZN(n20522) );
  OAI22_X1 U23476 ( .A1(n20566), .A2(n9930), .B1(n20522), .B2(n20521), .ZN(
        n20523) );
  INV_X1 U23477 ( .A(n20523), .ZN(n20525) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20529), .B1(
        n20527), .B2(n9935), .ZN(n20524) );
  OAI211_X1 U23479 ( .C1(n20532), .C2(n20600), .A(n20525), .B(n20524), .ZN(
        P1_U3119) );
  AOI22_X1 U23480 ( .A1(n20527), .A2(n9927), .B1(n20725), .B2(n20526), .ZN(
        n20531) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20529), .B1(
        n20528), .B2(n9941), .ZN(n20530) );
  OAI211_X1 U23482 ( .C1(n20532), .C2(n20607), .A(n20531), .B(n20530), .ZN(
        P1_U3120) );
  INV_X1 U23483 ( .A(n20533), .ZN(n20534) );
  NAND2_X1 U23484 ( .A1(n20534), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20538) );
  OAI21_X1 U23485 ( .B1(n20536), .B2(n20535), .A(n20538), .ZN(n20543) );
  INV_X1 U23486 ( .A(n20543), .ZN(n20537) );
  OAI22_X1 U23487 ( .A1(n20537), .A2(n20540), .B1(n20541), .B2(n20813), .ZN(
        n20562) );
  INV_X1 U23488 ( .A(n20538), .ZN(n20561) );
  AOI22_X1 U23489 ( .A1(n20682), .A2(n20562), .B1(n20561), .B2(n20681), .ZN(
        n20548) );
  AOI21_X1 U23490 ( .B1(n20546), .B2(n20688), .A(n20684), .ZN(n20544) );
  AOI21_X1 U23491 ( .B1(n20541), .B2(n20540), .A(n20539), .ZN(n20542) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20563), .B1(
        n20603), .B2(n9943), .ZN(n20547) );
  OAI211_X1 U23493 ( .C1(n20693), .C2(n20566), .A(n20548), .B(n20547), .ZN(
        P1_U3121) );
  AOI22_X1 U23494 ( .A1(n20695), .A2(n20562), .B1(n20561), .B2(n20694), .ZN(
        n20550) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20563), .B1(
        n20603), .B2(n9937), .ZN(n20549) );
  OAI211_X1 U23496 ( .C1(n9922), .C2(n20566), .A(n20550), .B(n20549), .ZN(
        P1_U3122) );
  AOI22_X1 U23497 ( .A1(n20700), .A2(n20562), .B1(n20561), .B2(n20699), .ZN(
        n20552) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20563), .B1(
        n20603), .B2(n9939), .ZN(n20551) );
  OAI211_X1 U23499 ( .C1(n9924), .C2(n20566), .A(n20552), .B(n20551), .ZN(
        P1_U3123) );
  AOI22_X1 U23500 ( .A1(n20705), .A2(n20562), .B1(n20561), .B2(n20704), .ZN(
        n20554) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20563), .B1(
        n20603), .B2(n20706), .ZN(n20553) );
  OAI211_X1 U23502 ( .C1(n9944), .C2(n20566), .A(n20554), .B(n20553), .ZN(
        P1_U3124) );
  AOI22_X1 U23503 ( .A1(n20710), .A2(n20562), .B1(n20561), .B2(n20709), .ZN(
        n20556) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20563), .B1(
        n20603), .B2(n9929), .ZN(n20555) );
  OAI211_X1 U23505 ( .C1(n9932), .C2(n20566), .A(n20556), .B(n20555), .ZN(
        P1_U3125) );
  AOI22_X1 U23506 ( .A1(n20715), .A2(n20562), .B1(n20561), .B2(n20714), .ZN(
        n20558) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20563), .B1(
        n20603), .B2(n9921), .ZN(n20557) );
  OAI211_X1 U23508 ( .C1(n20719), .C2(n20566), .A(n20558), .B(n20557), .ZN(
        P1_U3126) );
  AOI22_X1 U23509 ( .A1(n20721), .A2(n20562), .B1(n20561), .B2(n20720), .ZN(
        n20560) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20563), .B1(
        n20603), .B2(n9931), .ZN(n20559) );
  OAI211_X1 U23511 ( .C1(n9934), .C2(n20566), .A(n20560), .B(n20559), .ZN(
        P1_U3127) );
  AOI22_X1 U23512 ( .A1(n20728), .A2(n20562), .B1(n20561), .B2(n20725), .ZN(
        n20565) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20563), .B1(
        n20603), .B2(n9941), .ZN(n20564) );
  OAI211_X1 U23514 ( .C1(n9926), .C2(n20566), .A(n20565), .B(n20564), .ZN(
        P1_U3128) );
  NAND2_X1 U23515 ( .A1(n20636), .A2(n20688), .ZN(n20569) );
  OAI21_X1 U23516 ( .B1(n20603), .B2(n20569), .A(n20568), .ZN(n20577) );
  OR2_X1 U23517 ( .A1(n13382), .A2(n20570), .ZN(n20609) );
  NOR2_X1 U23518 ( .A1(n20609), .A2(n20639), .ZN(n20574) );
  NOR3_X1 U23519 ( .A1(n20573), .A2(n15688), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20615) );
  INV_X1 U23520 ( .A(n20615), .ZN(n20612) );
  NOR2_X1 U23521 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20612), .ZN(
        n20601) );
  AOI22_X1 U23522 ( .A1(n20602), .A2(n9943), .B1(n20681), .B2(n20601), .ZN(
        n20581) );
  INV_X1 U23523 ( .A(n20574), .ZN(n20576) );
  AOI22_X1 U23524 ( .A1(n20577), .A2(n20576), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20575), .ZN(n20578) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n20648), .ZN(n20580) );
  OAI211_X1 U23526 ( .C1(n20608), .C2(n20582), .A(n20581), .B(n20580), .ZN(
        P1_U3129) );
  AOI22_X1 U23527 ( .A1(n20602), .A2(n9937), .B1(n20694), .B2(n20601), .ZN(
        n20584) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n9923), .ZN(n20583) );
  OAI211_X1 U23529 ( .C1(n20608), .C2(n20585), .A(n20584), .B(n20583), .ZN(
        P1_U3130) );
  AOI22_X1 U23530 ( .A1(n20602), .A2(n9939), .B1(n20699), .B2(n20601), .ZN(
        n20587) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n9925), .ZN(n20586) );
  OAI211_X1 U23532 ( .C1(n20608), .C2(n20588), .A(n20587), .B(n20586), .ZN(
        P1_U3131) );
  AOI22_X1 U23533 ( .A1(n20602), .A2(n20706), .B1(n20704), .B2(n20601), .ZN(
        n20590) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n9945), .ZN(n20589) );
  OAI211_X1 U23535 ( .C1(n20608), .C2(n20591), .A(n20590), .B(n20589), .ZN(
        P1_U3132) );
  AOI22_X1 U23536 ( .A1(n20602), .A2(n9929), .B1(n20709), .B2(n20601), .ZN(
        n20593) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n9933), .ZN(n20592) );
  OAI211_X1 U23538 ( .C1(n20608), .C2(n20594), .A(n20593), .B(n20592), .ZN(
        P1_U3133) );
  AOI22_X1 U23539 ( .A1(n20602), .A2(n9921), .B1(n20714), .B2(n20601), .ZN(
        n20596) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n20664), .ZN(n20595) );
  OAI211_X1 U23541 ( .C1(n20608), .C2(n20597), .A(n20596), .B(n20595), .ZN(
        P1_U3134) );
  AOI22_X1 U23542 ( .A1(n20602), .A2(n9931), .B1(n20720), .B2(n20601), .ZN(
        n20599) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n9935), .ZN(n20598) );
  OAI211_X1 U23544 ( .C1(n20608), .C2(n20600), .A(n20599), .B(n20598), .ZN(
        P1_U3135) );
  AOI22_X1 U23545 ( .A1(n20602), .A2(n9941), .B1(n20725), .B2(n20601), .ZN(
        n20606) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20604), .B1(
        n20603), .B2(n9927), .ZN(n20605) );
  OAI211_X1 U23547 ( .C1(n20608), .C2(n20607), .A(n20606), .B(n20605), .ZN(
        P1_U3136) );
  INV_X1 U23548 ( .A(n20609), .ZN(n20679) );
  NOR2_X1 U23549 ( .A1(n20610), .A2(n20612), .ZN(n20631) );
  AOI21_X1 U23550 ( .B1(n20679), .B2(n20611), .A(n20631), .ZN(n20613) );
  OAI22_X1 U23551 ( .A1(n20613), .A2(n20540), .B1(n20612), .B2(n20813), .ZN(
        n20632) );
  AOI22_X1 U23552 ( .A1(n20682), .A2(n20632), .B1(n20681), .B2(n20631), .ZN(
        n20618) );
  OAI211_X1 U23553 ( .C1(n20685), .C2(n21140), .A(n20688), .B(n20613), .ZN(
        n20614) );
  OAI211_X1 U23554 ( .C1(n20688), .C2(n20615), .A(n20687), .B(n20614), .ZN(
        n20633) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20633), .B1(
        n20673), .B2(n9943), .ZN(n20617) );
  OAI211_X1 U23556 ( .C1(n20693), .C2(n20636), .A(n20618), .B(n20617), .ZN(
        P1_U3137) );
  AOI22_X1 U23557 ( .A1(n20695), .A2(n20632), .B1(n20694), .B2(n20631), .ZN(
        n20620) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20633), .B1(
        n20673), .B2(n9937), .ZN(n20619) );
  OAI211_X1 U23559 ( .C1(n9922), .C2(n20636), .A(n20620), .B(n20619), .ZN(
        P1_U3138) );
  AOI22_X1 U23560 ( .A1(n20700), .A2(n20632), .B1(n20699), .B2(n20631), .ZN(
        n20622) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20633), .B1(
        n20673), .B2(n9939), .ZN(n20621) );
  OAI211_X1 U23562 ( .C1(n9924), .C2(n20636), .A(n20622), .B(n20621), .ZN(
        P1_U3139) );
  AOI22_X1 U23563 ( .A1(n20705), .A2(n20632), .B1(n20704), .B2(n20631), .ZN(
        n20624) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20633), .B1(
        n20673), .B2(n20706), .ZN(n20623) );
  OAI211_X1 U23565 ( .C1(n9944), .C2(n20636), .A(n20624), .B(n20623), .ZN(
        P1_U3140) );
  AOI22_X1 U23566 ( .A1(n20710), .A2(n20632), .B1(n20709), .B2(n20631), .ZN(
        n20626) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20633), .B1(
        n20673), .B2(n9929), .ZN(n20625) );
  OAI211_X1 U23568 ( .C1(n9932), .C2(n20636), .A(n20626), .B(n20625), .ZN(
        P1_U3141) );
  AOI22_X1 U23569 ( .A1(n20715), .A2(n20632), .B1(n20714), .B2(n20631), .ZN(
        n20628) );
  AOI22_X1 U23570 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20633), .B1(
        n20673), .B2(n9921), .ZN(n20627) );
  OAI211_X1 U23571 ( .C1(n20719), .C2(n20636), .A(n20628), .B(n20627), .ZN(
        P1_U3142) );
  AOI22_X1 U23572 ( .A1(n20721), .A2(n20632), .B1(n20720), .B2(n20631), .ZN(
        n20630) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20633), .B1(
        n20673), .B2(n9931), .ZN(n20629) );
  OAI211_X1 U23574 ( .C1(n9934), .C2(n20636), .A(n20630), .B(n20629), .ZN(
        P1_U3143) );
  AOI22_X1 U23575 ( .A1(n20728), .A2(n20632), .B1(n20725), .B2(n20631), .ZN(
        n20635) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20633), .B1(
        n20673), .B2(n9941), .ZN(n20634) );
  OAI211_X1 U23577 ( .C1(n9926), .C2(n20636), .A(n20635), .B(n20634), .ZN(
        P1_U3144) );
  NAND2_X1 U23578 ( .A1(n20679), .A2(n20639), .ZN(n20643) );
  OAI22_X1 U23579 ( .A1(n20643), .A2(n20540), .B1(n20641), .B2(n20640), .ZN(
        n20671) );
  INV_X1 U23580 ( .A(n20689), .ZN(n20680) );
  NOR2_X1 U23581 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20680), .ZN(
        n20670) );
  AOI22_X1 U23582 ( .A1(n20682), .A2(n20671), .B1(n20681), .B2(n20670), .ZN(
        n20650) );
  INV_X1 U23583 ( .A(n20734), .ZN(n20642) );
  OAI21_X1 U23584 ( .B1(n20673), .B2(n20642), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20644) );
  AOI21_X1 U23585 ( .B1(n20644), .B2(n20643), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20647) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n20648), .ZN(n20649) );
  OAI211_X1 U23587 ( .C1(n9942), .C2(n20734), .A(n20650), .B(n20649), .ZN(
        P1_U3145) );
  AOI22_X1 U23588 ( .A1(n20695), .A2(n20671), .B1(n20694), .B2(n20670), .ZN(
        n20653) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n9923), .ZN(n20652) );
  OAI211_X1 U23590 ( .C1(n9936), .C2(n20734), .A(n20653), .B(n20652), .ZN(
        P1_U3146) );
  AOI22_X1 U23591 ( .A1(n20700), .A2(n20671), .B1(n20699), .B2(n20670), .ZN(
        n20656) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n9925), .ZN(n20655) );
  OAI211_X1 U23593 ( .C1(n9938), .C2(n20734), .A(n20656), .B(n20655), .ZN(
        P1_U3147) );
  AOI22_X1 U23594 ( .A1(n20705), .A2(n20671), .B1(n20704), .B2(n20670), .ZN(
        n20659) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n9945), .ZN(n20658) );
  OAI211_X1 U23596 ( .C1(n20660), .C2(n20734), .A(n20659), .B(n20658), .ZN(
        P1_U3148) );
  AOI22_X1 U23597 ( .A1(n20710), .A2(n20671), .B1(n20709), .B2(n20670), .ZN(
        n20663) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n9933), .ZN(n20662) );
  OAI211_X1 U23599 ( .C1(n9928), .C2(n20734), .A(n20663), .B(n20662), .ZN(
        P1_U3149) );
  AOI22_X1 U23600 ( .A1(n20715), .A2(n20671), .B1(n20714), .B2(n20670), .ZN(
        n20666) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n20664), .ZN(n20665) );
  OAI211_X1 U23602 ( .C1(n9920), .C2(n20734), .A(n20666), .B(n20665), .ZN(
        P1_U3150) );
  AOI22_X1 U23603 ( .A1(n20721), .A2(n20671), .B1(n20720), .B2(n20670), .ZN(
        n20669) );
  AOI22_X1 U23604 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n9935), .ZN(n20668) );
  OAI211_X1 U23605 ( .C1(n9930), .C2(n20734), .A(n20669), .B(n20668), .ZN(
        P1_U3151) );
  AOI22_X1 U23606 ( .A1(n20728), .A2(n20671), .B1(n20725), .B2(n20670), .ZN(
        n20676) );
  AOI22_X1 U23607 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20674), .B1(
        n20673), .B2(n9927), .ZN(n20675) );
  OAI211_X1 U23608 ( .C1(n9940), .C2(n20734), .A(n20676), .B(n20675), .ZN(
        P1_U3152) );
  INV_X1 U23609 ( .A(n20677), .ZN(n20726) );
  AOI21_X1 U23610 ( .B1(n20679), .B2(n20678), .A(n20726), .ZN(n20683) );
  OAI22_X1 U23611 ( .A1(n20683), .A2(n20540), .B1(n20813), .B2(n20680), .ZN(
        n20727) );
  AOI22_X1 U23612 ( .A1(n20682), .A2(n20727), .B1(n20726), .B2(n20681), .ZN(
        n20692) );
  OAI211_X1 U23613 ( .C1(n20685), .C2(n20684), .A(n20688), .B(n20683), .ZN(
        n20686) );
  OAI211_X1 U23614 ( .C1(n20689), .C2(n20688), .A(n20687), .B(n20686), .ZN(
        n20731) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20731), .B1(
        n20730), .B2(n9943), .ZN(n20691) );
  OAI211_X1 U23616 ( .C1(n20693), .C2(n20734), .A(n20692), .B(n20691), .ZN(
        P1_U3153) );
  AOI22_X1 U23617 ( .A1(n20695), .A2(n20727), .B1(n20726), .B2(n20694), .ZN(
        n20698) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20731), .B1(
        n20730), .B2(n9937), .ZN(n20697) );
  OAI211_X1 U23619 ( .C1(n9922), .C2(n20734), .A(n20698), .B(n20697), .ZN(
        P1_U3154) );
  AOI22_X1 U23620 ( .A1(n20700), .A2(n20727), .B1(n20726), .B2(n20699), .ZN(
        n20703) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20731), .B1(
        n20730), .B2(n9939), .ZN(n20702) );
  OAI211_X1 U23622 ( .C1(n9924), .C2(n20734), .A(n20703), .B(n20702), .ZN(
        P1_U3155) );
  AOI22_X1 U23623 ( .A1(n20705), .A2(n20727), .B1(n20726), .B2(n20704), .ZN(
        n20708) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20731), .B1(
        n20730), .B2(n20706), .ZN(n20707) );
  OAI211_X1 U23625 ( .C1(n9944), .C2(n20734), .A(n20708), .B(n20707), .ZN(
        P1_U3156) );
  AOI22_X1 U23626 ( .A1(n20710), .A2(n20727), .B1(n20726), .B2(n20709), .ZN(
        n20713) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20731), .B1(
        n20730), .B2(n9929), .ZN(n20712) );
  OAI211_X1 U23628 ( .C1(n9932), .C2(n20734), .A(n20713), .B(n20712), .ZN(
        P1_U3157) );
  AOI22_X1 U23629 ( .A1(n20715), .A2(n20727), .B1(n20726), .B2(n20714), .ZN(
        n20718) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20731), .B1(
        n20730), .B2(n9921), .ZN(n20717) );
  OAI211_X1 U23631 ( .C1(n20719), .C2(n20734), .A(n20718), .B(n20717), .ZN(
        P1_U3158) );
  AOI22_X1 U23632 ( .A1(n20721), .A2(n20727), .B1(n20726), .B2(n20720), .ZN(
        n20724) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20731), .B1(
        n20730), .B2(n9931), .ZN(n20723) );
  OAI211_X1 U23634 ( .C1(n9934), .C2(n20734), .A(n20724), .B(n20723), .ZN(
        P1_U3159) );
  AOI22_X1 U23635 ( .A1(n20728), .A2(n20727), .B1(n20726), .B2(n20725), .ZN(
        n20733) );
  AOI22_X1 U23636 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20731), .B1(
        n20730), .B2(n9941), .ZN(n20732) );
  OAI211_X1 U23637 ( .C1(n9926), .C2(n20734), .A(n20733), .B(n20732), .ZN(
        P1_U3160) );
  OAI221_X1 U23638 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20737), .C1(n20813), 
        .C2(n20736), .A(n20735), .ZN(P1_U3163) );
  AND2_X1 U23639 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20791), .ZN(
        P1_U3164) );
  AND2_X1 U23640 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20791), .ZN(
        P1_U3165) );
  AND2_X1 U23641 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20791), .ZN(
        P1_U3166) );
  AND2_X1 U23642 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20791), .ZN(
        P1_U3167) );
  AND2_X1 U23643 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20791), .ZN(
        P1_U3168) );
  AND2_X1 U23644 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20791), .ZN(
        P1_U3169) );
  AND2_X1 U23645 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20791), .ZN(
        P1_U3170) );
  AND2_X1 U23646 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20791), .ZN(
        P1_U3171) );
  AND2_X1 U23647 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20791), .ZN(
        P1_U3172) );
  AND2_X1 U23648 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20791), .ZN(
        P1_U3173) );
  AND2_X1 U23649 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20791), .ZN(
        P1_U3174) );
  AND2_X1 U23650 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20791), .ZN(
        P1_U3175) );
  AND2_X1 U23651 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20791), .ZN(
        P1_U3176) );
  AND2_X1 U23652 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20791), .ZN(
        P1_U3177) );
  AND2_X1 U23653 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20791), .ZN(
        P1_U3178) );
  AND2_X1 U23654 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20791), .ZN(
        P1_U3179) );
  AND2_X1 U23655 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20791), .ZN(
        P1_U3180) );
  AND2_X1 U23656 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20791), .ZN(
        P1_U3181) );
  AND2_X1 U23657 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20791), .ZN(
        P1_U3182) );
  AND2_X1 U23658 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20791), .ZN(
        P1_U3183) );
  AND2_X1 U23659 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20791), .ZN(
        P1_U3184) );
  AND2_X1 U23660 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20791), .ZN(
        P1_U3185) );
  AND2_X1 U23661 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20791), .ZN(P1_U3186) );
  AND2_X1 U23662 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20791), .ZN(P1_U3187) );
  AND2_X1 U23663 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20791), .ZN(P1_U3188) );
  AND2_X1 U23664 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20791), .ZN(P1_U3189) );
  AND2_X1 U23665 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20791), .ZN(P1_U3190) );
  AND2_X1 U23666 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20791), .ZN(P1_U3191) );
  AND2_X1 U23667 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20791), .ZN(P1_U3192) );
  AND2_X1 U23668 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20791), .ZN(P1_U3193) );
  OAI21_X1 U23669 ( .B1(n20748), .B2(n20820), .A(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20744) );
  INV_X1 U23670 ( .A(n20744), .ZN(n20741) );
  OAI22_X1 U23671 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21052), .B1(n20749), 
        .B2(n20988), .ZN(n20738) );
  NOR3_X1 U23672 ( .A1(n20739), .A2(n21175), .A3(n20738), .ZN(n20740) );
  OAI22_X1 U23673 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20741), .B1(n20830), 
        .B2(n20740), .ZN(P1_U3194) );
  NAND4_X1 U23674 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20814), .A3(
        P1_REQUESTPENDING_REG_SCAN_IN), .A4(n21052), .ZN(n20747) );
  NAND2_X1 U23675 ( .A1(n20814), .A2(n21052), .ZN(n20742) );
  OAI221_X1 U23676 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(
        n20742), .A(n20749), .ZN(n20743) );
  NAND3_X1 U23677 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(HOLD), .A3(n20743), .ZN(
        n20746) );
  OAI211_X1 U23678 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21052), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20744), .ZN(n20745) );
  OAI211_X1 U23679 ( .C1(n20748), .C2(n20747), .A(n20746), .B(n20745), .ZN(
        P1_U3196) );
  OR2_X1 U23680 ( .A1(n20829), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20769) );
  INV_X1 U23681 ( .A(n20769), .ZN(n20783) );
  NOR2_X1 U23682 ( .A1(n20749), .A2(n20829), .ZN(n20784) );
  INV_X1 U23683 ( .A(n20784), .ZN(n20767) );
  INV_X1 U23684 ( .A(n20767), .ZN(n20775) );
  AOI222_X1 U23685 ( .A1(n20783), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20775), .ZN(n20750) );
  INV_X1 U23686 ( .A(n20750), .ZN(P1_U3197) );
  AOI222_X1 U23687 ( .A1(n20775), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20783), .ZN(n20751) );
  INV_X1 U23688 ( .A(n20751), .ZN(P1_U3198) );
  OAI222_X1 U23689 ( .A1(n20767), .A2(n20912), .B1(n20752), .B2(n20830), .C1(
        n20962), .C2(n20769), .ZN(P1_U3199) );
  INV_X1 U23690 ( .A(n20769), .ZN(n20780) );
  AOI222_X1 U23691 ( .A1(n20775), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20780), .ZN(n20753) );
  INV_X1 U23692 ( .A(n20753), .ZN(P1_U3200) );
  AOI222_X1 U23693 ( .A1(n20780), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20775), .ZN(n20754) );
  INV_X1 U23694 ( .A(n20754), .ZN(P1_U3201) );
  AOI222_X1 U23695 ( .A1(n20775), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20780), .ZN(n20755) );
  INV_X1 U23696 ( .A(n20755), .ZN(P1_U3202) );
  AOI222_X1 U23697 ( .A1(n20775), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20780), .ZN(n20756) );
  INV_X1 U23698 ( .A(n20756), .ZN(P1_U3203) );
  AOI222_X1 U23699 ( .A1(n20783), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20775), .ZN(n20757) );
  INV_X1 U23700 ( .A(n20757), .ZN(P1_U3204) );
  AOI222_X1 U23701 ( .A1(n20783), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20775), .ZN(n20758) );
  INV_X1 U23702 ( .A(n20758), .ZN(P1_U3205) );
  AOI222_X1 U23703 ( .A1(n20783), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20775), .ZN(n20759) );
  INV_X1 U23704 ( .A(n20759), .ZN(P1_U3206) );
  AOI222_X1 U23705 ( .A1(n20780), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20775), .ZN(n20760) );
  INV_X1 U23706 ( .A(n20760), .ZN(P1_U3207) );
  AOI222_X1 U23707 ( .A1(n20784), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20780), .ZN(n20761) );
  INV_X1 U23708 ( .A(n20761), .ZN(P1_U3208) );
  AOI222_X1 U23709 ( .A1(n20784), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20783), .ZN(n20762) );
  INV_X1 U23710 ( .A(n20762), .ZN(P1_U3209) );
  AOI222_X1 U23711 ( .A1(n20780), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20775), .ZN(n20763) );
  INV_X1 U23712 ( .A(n20763), .ZN(P1_U3210) );
  AOI222_X1 U23713 ( .A1(n20784), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20783), .ZN(n20764) );
  INV_X1 U23714 ( .A(n20764), .ZN(P1_U3211) );
  AOI222_X1 U23715 ( .A1(n20775), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20783), .ZN(n20765) );
  INV_X1 U23716 ( .A(n20765), .ZN(P1_U3212) );
  INV_X1 U23717 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20918) );
  AOI22_X1 U23718 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20829), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20780), .ZN(n20766) );
  OAI21_X1 U23719 ( .B1(n20918), .B2(n20767), .A(n20766), .ZN(P1_U3213) );
  AOI22_X1 U23720 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20829), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n20784), .ZN(n20768) );
  OAI21_X1 U23721 ( .B1(n21157), .B2(n20769), .A(n20768), .ZN(P1_U3214) );
  AOI222_X1 U23722 ( .A1(n20775), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20783), .ZN(n20770) );
  INV_X1 U23723 ( .A(n20770), .ZN(P1_U3215) );
  AOI222_X1 U23724 ( .A1(n20783), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20775), .ZN(n20771) );
  INV_X1 U23725 ( .A(n20771), .ZN(P1_U3216) );
  AOI222_X1 U23726 ( .A1(n20780), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20775), .ZN(n20772) );
  INV_X1 U23727 ( .A(n20772), .ZN(P1_U3217) );
  AOI222_X1 U23728 ( .A1(n20775), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20783), .ZN(n20773) );
  INV_X1 U23729 ( .A(n20773), .ZN(P1_U3218) );
  AOI222_X1 U23730 ( .A1(n20775), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20783), .ZN(n20774) );
  INV_X1 U23731 ( .A(n20774), .ZN(P1_U3219) );
  AOI222_X1 U23732 ( .A1(n20775), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20783), .ZN(n20776) );
  INV_X1 U23733 ( .A(n20776), .ZN(P1_U3220) );
  AOI222_X1 U23734 ( .A1(n20780), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20784), .ZN(n20777) );
  INV_X1 U23735 ( .A(n20777), .ZN(P1_U3221) );
  AOI222_X1 U23736 ( .A1(n20784), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20783), .ZN(n20778) );
  INV_X1 U23737 ( .A(n20778), .ZN(P1_U3222) );
  AOI222_X1 U23738 ( .A1(n20783), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20784), .ZN(n20779) );
  INV_X1 U23739 ( .A(n20779), .ZN(P1_U3223) );
  AOI222_X1 U23740 ( .A1(n20780), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20784), .ZN(n20781) );
  INV_X1 U23741 ( .A(n20781), .ZN(P1_U3224) );
  AOI222_X1 U23742 ( .A1(n20784), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20783), .ZN(n20782) );
  INV_X1 U23743 ( .A(n20782), .ZN(P1_U3225) );
  AOI222_X1 U23744 ( .A1(n20784), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20829), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20783), .ZN(n20785) );
  INV_X1 U23745 ( .A(n20785), .ZN(P1_U3226) );
  OAI22_X1 U23746 ( .A1(n20829), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20830), .ZN(n20786) );
  INV_X1 U23747 ( .A(n20786), .ZN(P1_U3458) );
  OAI22_X1 U23748 ( .A1(n20829), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20830), .ZN(n20787) );
  INV_X1 U23749 ( .A(n20787), .ZN(P1_U3459) );
  OAI22_X1 U23750 ( .A1(n20829), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20830), .ZN(n20788) );
  INV_X1 U23751 ( .A(n20788), .ZN(P1_U3460) );
  OAI22_X1 U23752 ( .A1(n20829), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20830), .ZN(n20789) );
  INV_X1 U23753 ( .A(n20789), .ZN(P1_U3461) );
  INV_X1 U23754 ( .A(n20793), .ZN(n20790) );
  AOI21_X1 U23755 ( .B1(n20792), .B2(n20791), .A(n20790), .ZN(P1_U3464) );
  INV_X1 U23756 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20794) );
  OAI21_X1 U23757 ( .B1(n20795), .B2(n20794), .A(n20793), .ZN(P1_U3465) );
  AOI22_X1 U23758 ( .A1(n20799), .A2(n20798), .B1(n20797), .B2(n20796), .ZN(
        n20800) );
  INV_X1 U23759 ( .A(n20800), .ZN(n20802) );
  MUX2_X1 U23760 ( .A(n20802), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20801), .Z(P1_U3469) );
  INV_X1 U23761 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21014) );
  AOI21_X1 U23762 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(
        P1_REIP_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20803)
         );
  OAI221_X1 U23763 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20803), .C1(n13638), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20805), .ZN(n20804) );
  OAI21_X1 U23764 ( .B1(n20805), .B2(n21014), .A(n20804), .ZN(P1_U3481) );
  INV_X1 U23765 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20808) );
  NOR2_X1 U23766 ( .A1(n20807), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20806) );
  AOI22_X1 U23767 ( .A1(n20808), .A2(n20807), .B1(n14021), .B2(n20806), .ZN(
        P1_U3482) );
  AOI22_X1 U23768 ( .A1(n20830), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20966), 
        .B2(n20829), .ZN(P1_U3483) );
  INV_X1 U23769 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n20810) );
  AOI22_X1 U23770 ( .A1(n20812), .A2(n20811), .B1(n20810), .B2(n20809), .ZN(
        P1_U3484) );
  NOR2_X1 U23771 ( .A1(n20814), .A2(n20813), .ZN(n20817) );
  AOI211_X1 U23772 ( .C1(n20818), .C2(n20817), .A(n20816), .B(n20815), .ZN(
        n20828) );
  AOI21_X1 U23773 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20821), .A(n20819), 
        .ZN(n20824) );
  OAI211_X1 U23774 ( .C1(n20822), .C2(n20821), .A(P1_STATE2_REG_2__SCAN_IN), 
        .B(n20820), .ZN(n20823) );
  OAI21_X1 U23775 ( .B1(n20824), .B2(n20823), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n20827) );
  NOR2_X1 U23776 ( .A1(n20828), .A2(n20825), .ZN(n20826) );
  AOI22_X1 U23777 ( .A1(n21175), .A2(n20828), .B1(n20827), .B2(n20826), .ZN(
        P1_U3485) );
  AOI22_X1 U23778 ( .A1(n20830), .A2(n21188), .B1(n21156), .B2(n20829), .ZN(
        P1_U3486) );
  AOI22_X1 U23779 ( .A1(n20832), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n20831), .ZN(n21214) );
  OAI22_X1 U23780 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_g104), .B1(
        keyinput_g7), .B2(DATAI_25_), .ZN(n20833) );
  AOI221_X1 U23781 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_g104), .C1(
        DATAI_25_), .C2(keyinput_g7), .A(n20833), .ZN(n20840) );
  OAI22_X1 U23782 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_g52), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .ZN(n20834) );
  AOI221_X1 U23783 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_g52), .C1(
        keyinput_g63), .C2(P1_REIP_REG_20__SCAN_IN), .A(n20834), .ZN(n20839)
         );
  OAI22_X1 U23784 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_g55), .B1(
        keyinput_g6), .B2(DATAI_26_), .ZN(n20835) );
  AOI221_X1 U23785 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .C1(
        DATAI_26_), .C2(keyinput_g6), .A(n20835), .ZN(n20838) );
  OAI22_X1 U23786 ( .A1(DATAI_24_), .A2(keyinput_g8), .B1(keyinput_g0), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20836) );
  AOI221_X1 U23787 ( .B1(DATAI_24_), .B2(keyinput_g8), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_g0), .A(n20836), .ZN(n20837)
         );
  NAND4_X1 U23788 ( .A1(n20840), .A2(n20839), .A3(n20838), .A4(n20837), .ZN(
        n20869) );
  OAI22_X1 U23789 ( .A1(P1_EBX_REG_17__SCAN_IN), .A2(keyinput_g98), .B1(
        keyinput_g72), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n20841) );
  AOI221_X1 U23790 ( .B1(P1_EBX_REG_17__SCAN_IN), .B2(keyinput_g98), .C1(
        P1_REIP_REG_11__SCAN_IN), .C2(keyinput_g72), .A(n20841), .ZN(n20848)
         );
  OAI22_X1 U23791 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(keyinput_g69), .B1(
        DATAI_8_), .B2(keyinput_g24), .ZN(n20842) );
  AOI221_X1 U23792 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(keyinput_g69), .C1(
        keyinput_g24), .C2(DATAI_8_), .A(n20842), .ZN(n20847) );
  OAI22_X1 U23793 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_g88), .B1(READY2), .B2(keyinput_g37), .ZN(n20843) );
  AOI221_X1 U23794 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_g88), .C1(
        keyinput_g37), .C2(READY2), .A(n20843), .ZN(n20846) );
  OAI22_X1 U23795 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_g116), .B1(
        keyinput_g23), .B2(DATAI_9_), .ZN(n20844) );
  AOI221_X1 U23796 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_g116), .C1(
        DATAI_9_), .C2(keyinput_g23), .A(n20844), .ZN(n20845) );
  NAND4_X1 U23797 ( .A1(n20848), .A2(n20847), .A3(n20846), .A4(n20845), .ZN(
        n20868) );
  OAI22_X1 U23798 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(keyinput_g102), .B1(
        keyinput_g34), .B2(NA), .ZN(n20849) );
  AOI221_X1 U23799 ( .B1(P1_EBX_REG_13__SCAN_IN), .B2(keyinput_g102), .C1(NA), 
        .C2(keyinput_g34), .A(n20849), .ZN(n20856) );
  OAI22_X1 U23800 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        keyinput_g48), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20850) );
  AOI221_X1 U23801 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_g48), .A(n20850), .ZN(
        n20855) );
  OAI22_X1 U23802 ( .A1(P1_EBX_REG_26__SCAN_IN), .A2(keyinput_g89), .B1(
        keyinput_g108), .B2(P1_EBX_REG_7__SCAN_IN), .ZN(n20851) );
  AOI221_X1 U23803 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(keyinput_g89), .C1(
        P1_EBX_REG_7__SCAN_IN), .C2(keyinput_g108), .A(n20851), .ZN(n20854) );
  OAI22_X1 U23804 ( .A1(P1_EBX_REG_23__SCAN_IN), .A2(keyinput_g92), .B1(
        keyinput_g12), .B2(DATAI_20_), .ZN(n20852) );
  AOI221_X1 U23805 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(keyinput_g92), .C1(
        DATAI_20_), .C2(keyinput_g12), .A(n20852), .ZN(n20853) );
  NAND4_X1 U23806 ( .A1(n20856), .A2(n20855), .A3(n20854), .A4(n20853), .ZN(
        n20867) );
  OAI22_X1 U23807 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(keyinput_g114), .B1(
        DATAI_16_), .B2(keyinput_g16), .ZN(n20857) );
  AOI221_X1 U23808 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput_g114), .C1(
        keyinput_g16), .C2(DATAI_16_), .A(n20857), .ZN(n20865) );
  OAI22_X1 U23809 ( .A1(DATAI_19_), .A2(keyinput_g13), .B1(keyinput_g29), .B2(
        DATAI_3_), .ZN(n20858) );
  AOI221_X1 U23810 ( .B1(DATAI_19_), .B2(keyinput_g13), .C1(DATAI_3_), .C2(
        keyinput_g29), .A(n20858), .ZN(n20864) );
  OAI22_X1 U23811 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_g60), .B1(
        keyinput_g61), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n20859) );
  AOI221_X1 U23812 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_g61), .A(n20859), .ZN(n20863)
         );
  OAI22_X1 U23813 ( .A1(n20861), .A2(keyinput_g4), .B1(keyinput_g56), .B2(
        P1_REIP_REG_27__SCAN_IN), .ZN(n20860) );
  AOI221_X1 U23814 ( .B1(n20861), .B2(keyinput_g4), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_g56), .A(n20860), .ZN(n20862)
         );
  NAND4_X1 U23815 ( .A1(n20865), .A2(n20864), .A3(n20863), .A4(n20862), .ZN(
        n20866) );
  NOR4_X1 U23816 ( .A1(n20869), .A2(n20868), .A3(n20867), .A4(n20866), .ZN(
        n21004) );
  OAI22_X1 U23817 ( .A1(READY1), .A2(keyinput_g36), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(keyinput_g65), .ZN(n20870) );
  AOI221_X1 U23818 ( .B1(READY1), .B2(keyinput_g36), .C1(keyinput_g65), .C2(
        P1_REIP_REG_18__SCAN_IN), .A(n20870), .ZN(n20877) );
  OAI22_X1 U23819 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(keyinput_g107), .B1(
        keyinput_g20), .B2(DATAI_12_), .ZN(n20871) );
  AOI221_X1 U23820 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(keyinput_g107), .C1(
        DATAI_12_), .C2(keyinput_g20), .A(n20871), .ZN(n20876) );
  OAI22_X1 U23821 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(keyinput_g110), .B1(
        keyinput_g32), .B2(DATAI_0_), .ZN(n20872) );
  AOI221_X1 U23822 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput_g110), .C1(
        DATAI_0_), .C2(keyinput_g32), .A(n20872), .ZN(n20875) );
  OAI22_X1 U23823 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_g57), .B1(
        keyinput_g76), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n20873) );
  AOI221_X1 U23824 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(keyinput_g76), .A(n20873), .ZN(n20874) );
  NAND4_X1 U23825 ( .A1(n20877), .A2(n20876), .A3(n20875), .A4(n20874), .ZN(
        n21002) );
  OAI22_X1 U23826 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_g112), .B1(
        keyinput_g111), .B2(P1_EBX_REG_4__SCAN_IN), .ZN(n20878) );
  AOI221_X1 U23827 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_g112), .C1(
        P1_EBX_REG_4__SCAN_IN), .C2(keyinput_g111), .A(n20878), .ZN(n20903) );
  OAI22_X1 U23828 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_g101), .B1(
        keyinput_g74), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n20879) );
  AOI221_X1 U23829 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_g101), .C1(
        P1_REIP_REG_9__SCAN_IN), .C2(keyinput_g74), .A(n20879), .ZN(n20882) );
  OAI22_X1 U23830 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(keyinput_g105), .B1(
        keyinput_g45), .B2(P1_MORE_REG_SCAN_IN), .ZN(n20880) );
  AOI221_X1 U23831 ( .B1(P1_EBX_REG_10__SCAN_IN), .B2(keyinput_g105), .C1(
        P1_MORE_REG_SCAN_IN), .C2(keyinput_g45), .A(n20880), .ZN(n20881) );
  OAI211_X1 U23832 ( .C1(n15894), .C2(keyinput_g15), .A(n20882), .B(n20881), 
        .ZN(n20883) );
  AOI21_X1 U23833 ( .B1(n15894), .B2(keyinput_g15), .A(n20883), .ZN(n20902) );
  AOI22_X1 U23834 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(keyinput_g73), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(keyinput_g93), .ZN(n20884) );
  OAI221_X1 U23835 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(keyinput_g73), .C1(
        P1_EBX_REG_22__SCAN_IN), .C2(keyinput_g93), .A(n20884), .ZN(n20891) );
  AOI22_X1 U23836 ( .A1(DATAI_21_), .A2(keyinput_g11), .B1(DATAI_13_), .B2(
        keyinput_g19), .ZN(n20885) );
  OAI221_X1 U23837 ( .B1(DATAI_21_), .B2(keyinput_g11), .C1(DATAI_13_), .C2(
        keyinput_g19), .A(n20885), .ZN(n20890) );
  AOI22_X1 U23838 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_g62), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(keyinput_g127), .ZN(n20886) );
  OAI221_X1 U23839 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .C1(
        P1_EAX_REG_20__SCAN_IN), .C2(keyinput_g127), .A(n20886), .ZN(n20889)
         );
  AOI22_X1 U23840 ( .A1(DATAI_30_), .A2(keyinput_g2), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(keyinput_g68), .ZN(n20887) );
  OAI221_X1 U23841 ( .B1(DATAI_30_), .B2(keyinput_g2), .C1(
        P1_REIP_REG_15__SCAN_IN), .C2(keyinput_g68), .A(n20887), .ZN(n20888)
         );
  NOR4_X1 U23842 ( .A1(n20891), .A2(n20890), .A3(n20889), .A4(n20888), .ZN(
        n20901) );
  AOI22_X1 U23843 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput_g85), .ZN(n20892) );
  OAI221_X1 U23844 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput_g85), .A(n20892), .ZN(n20899) );
  AOI22_X1 U23845 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(keyinput_g64), .B1(
        P1_EBX_REG_2__SCAN_IN), .B2(keyinput_g113), .ZN(n20893) );
  OAI221_X1 U23846 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput_g64), .C1(
        P1_EBX_REG_2__SCAN_IN), .C2(keyinput_g113), .A(n20893), .ZN(n20898) );
  AOI22_X1 U23847 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g51), .B1(
        DATAI_6_), .B2(keyinput_g26), .ZN(n20894) );
  OAI221_X1 U23848 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g51), 
        .C1(DATAI_6_), .C2(keyinput_g26), .A(n20894), .ZN(n20897) );
  AOI22_X1 U23849 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_g46), .B1(
        DATAI_23_), .B2(keyinput_g9), .ZN(n20895) );
  OAI221_X1 U23850 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .C1(
        DATAI_23_), .C2(keyinput_g9), .A(n20895), .ZN(n20896) );
  NOR4_X1 U23851 ( .A1(n20899), .A2(n20898), .A3(n20897), .A4(n20896), .ZN(
        n20900) );
  NAND4_X1 U23852 ( .A1(n20903), .A2(n20902), .A3(n20901), .A4(n20900), .ZN(
        n21001) );
  INV_X1 U23853 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21173) );
  AOI22_X1 U23854 ( .A1(n21173), .A2(keyinput_g71), .B1(n20905), .B2(
        keyinput_g100), .ZN(n20904) );
  OAI221_X1 U23855 ( .B1(n21173), .B2(keyinput_g71), .C1(n20905), .C2(
        keyinput_g100), .A(n20904), .ZN(n20916) );
  AOI22_X1 U23856 ( .A1(n20908), .A2(keyinput_g54), .B1(n20907), .B2(
        keyinput_g109), .ZN(n20906) );
  OAI221_X1 U23857 ( .B1(n20908), .B2(keyinput_g54), .C1(n20907), .C2(
        keyinput_g109), .A(n20906), .ZN(n20915) );
  AOI22_X1 U23858 ( .A1(n14193), .A2(keyinput_g75), .B1(keyinput_g53), .B2(
        n20910), .ZN(n20909) );
  OAI221_X1 U23859 ( .B1(n14193), .B2(keyinput_g75), .C1(n20910), .C2(
        keyinput_g53), .A(n20909), .ZN(n20914) );
  AOI22_X1 U23860 ( .A1(n20912), .A2(keyinput_g80), .B1(n21011), .B2(
        keyinput_g1), .ZN(n20911) );
  OAI221_X1 U23861 ( .B1(n20912), .B2(keyinput_g80), .C1(n21011), .C2(
        keyinput_g1), .A(n20911), .ZN(n20913) );
  NOR4_X1 U23862 ( .A1(n20916), .A2(n20915), .A3(n20914), .A4(n20913), .ZN(
        n20951) );
  AOI22_X1 U23863 ( .A1(n20919), .A2(keyinput_g86), .B1(keyinput_g66), .B2(
        n20918), .ZN(n20917) );
  OAI221_X1 U23864 ( .B1(n20919), .B2(keyinput_g86), .C1(n20918), .C2(
        keyinput_g66), .A(n20917), .ZN(n20928) );
  AOI22_X1 U23865 ( .A1(n20921), .A2(keyinput_g106), .B1(n11581), .B2(
        keyinput_g124), .ZN(n20920) );
  OAI221_X1 U23866 ( .B1(n20921), .B2(keyinput_g106), .C1(n11581), .C2(
        keyinput_g124), .A(n20920), .ZN(n20927) );
  AOI22_X1 U23867 ( .A1(n21175), .A2(keyinput_g43), .B1(n14016), .B2(
        keyinput_g115), .ZN(n20922) );
  OAI221_X1 U23868 ( .B1(n21175), .B2(keyinput_g43), .C1(n14016), .C2(
        keyinput_g115), .A(n20922), .ZN(n20926) );
  AOI22_X1 U23869 ( .A1(n20924), .A2(keyinput_g87), .B1(keyinput_g50), .B2(
        n21014), .ZN(n20923) );
  OAI221_X1 U23870 ( .B1(n20924), .B2(keyinput_g87), .C1(n21014), .C2(
        keyinput_g50), .A(n20923), .ZN(n20925) );
  NOR4_X1 U23871 ( .A1(n20928), .A2(n20927), .A3(n20926), .A4(n20925), .ZN(
        n20950) );
  AOI22_X1 U23872 ( .A1(n11606), .A2(keyinput_g123), .B1(keyinput_g82), .B2(
        n13638), .ZN(n20929) );
  OAI221_X1 U23873 ( .B1(n11606), .B2(keyinput_g123), .C1(n13638), .C2(
        keyinput_g82), .A(n20929), .ZN(n20938) );
  AOI22_X1 U23874 ( .A1(n20931), .A2(keyinput_g67), .B1(n21128), .B2(
        keyinput_g91), .ZN(n20930) );
  OAI221_X1 U23875 ( .B1(n20931), .B2(keyinput_g67), .C1(n21128), .C2(
        keyinput_g91), .A(n20930), .ZN(n20937) );
  INV_X1 U23876 ( .A(DATAI_10_), .ZN(n20933) );
  AOI22_X1 U23877 ( .A1(n21176), .A2(keyinput_g126), .B1(keyinput_g22), .B2(
        n20933), .ZN(n20932) );
  OAI221_X1 U23878 ( .B1(n21176), .B2(keyinput_g126), .C1(n20933), .C2(
        keyinput_g22), .A(n20932), .ZN(n20936) );
  INV_X1 U23879 ( .A(DATAI_14_), .ZN(n21006) );
  AOI22_X1 U23880 ( .A1(n21006), .A2(keyinput_g18), .B1(n21050), .B2(
        keyinput_g99), .ZN(n20934) );
  OAI221_X1 U23881 ( .B1(n21006), .B2(keyinput_g18), .C1(n21050), .C2(
        keyinput_g99), .A(n20934), .ZN(n20935) );
  NOR4_X1 U23882 ( .A1(n20938), .A2(n20937), .A3(n20936), .A4(n20935), .ZN(
        n20949) );
  AOI22_X1 U23883 ( .A1(n20940), .A2(keyinput_g77), .B1(n21008), .B2(
        keyinput_g97), .ZN(n20939) );
  OAI221_X1 U23884 ( .B1(n20940), .B2(keyinput_g77), .C1(n21008), .C2(
        keyinput_g97), .A(n20939), .ZN(n20947) );
  AOI22_X1 U23885 ( .A1(n21191), .A2(keyinput_g81), .B1(n21140), .B2(
        keyinput_g44), .ZN(n20941) );
  OAI221_X1 U23886 ( .B1(n21191), .B2(keyinput_g81), .C1(n21140), .C2(
        keyinput_g44), .A(n20941), .ZN(n20946) );
  AOI22_X1 U23887 ( .A1(n21047), .A2(keyinput_g90), .B1(keyinput_g83), .B2(
        n14021), .ZN(n20942) );
  OAI221_X1 U23888 ( .B1(n21047), .B2(keyinput_g90), .C1(n14021), .C2(
        keyinput_g83), .A(n20942), .ZN(n20945) );
  INV_X1 U23889 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21079) );
  AOI22_X1 U23890 ( .A1(n21156), .A2(keyinput_g41), .B1(n21079), .B2(
        keyinput_g38), .ZN(n20943) );
  OAI221_X1 U23891 ( .B1(n21156), .B2(keyinput_g41), .C1(n21079), .C2(
        keyinput_g38), .A(n20943), .ZN(n20944) );
  NOR4_X1 U23892 ( .A1(n20947), .A2(n20946), .A3(n20945), .A4(n20944), .ZN(
        n20948) );
  NAND4_X1 U23893 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n21000) );
  INV_X1 U23894 ( .A(DATAI_4_), .ZN(n21015) );
  INV_X1 U23895 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21049) );
  AOI22_X1 U23896 ( .A1(n21015), .A2(keyinput_g28), .B1(keyinput_g40), .B2(
        n21049), .ZN(n20952) );
  OAI221_X1 U23897 ( .B1(n21015), .B2(keyinput_g28), .C1(n21049), .C2(
        keyinput_g40), .A(n20952), .ZN(n20960) );
  INV_X1 U23898 ( .A(DATAI_1_), .ZN(n21034) );
  AOI22_X1 U23899 ( .A1(n21026), .A2(keyinput_g94), .B1(keyinput_g31), .B2(
        n21034), .ZN(n20953) );
  OAI221_X1 U23900 ( .B1(n21026), .B2(keyinput_g94), .C1(n21034), .C2(
        keyinput_g31), .A(n20953), .ZN(n20959) );
  INV_X1 U23901 ( .A(DATAI_5_), .ZN(n21161) );
  AOI22_X1 U23902 ( .A1(n21161), .A2(keyinput_g27), .B1(n21153), .B2(
        keyinput_g5), .ZN(n20954) );
  OAI221_X1 U23903 ( .B1(n21161), .B2(keyinput_g27), .C1(n21153), .C2(
        keyinput_g5), .A(n20954), .ZN(n20958) );
  INV_X1 U23904 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20956) );
  AOI22_X1 U23905 ( .A1(n20956), .A2(keyinput_g58), .B1(n21141), .B2(
        keyinput_g122), .ZN(n20955) );
  OAI221_X1 U23906 ( .B1(n20956), .B2(keyinput_g58), .C1(n21141), .C2(
        keyinput_g122), .A(n20955), .ZN(n20957) );
  NOR4_X1 U23907 ( .A1(n20960), .A2(n20959), .A3(n20958), .A4(n20957), .ZN(
        n20998) );
  AOI22_X1 U23908 ( .A1(n21170), .A2(keyinput_g14), .B1(n20962), .B2(
        keyinput_g79), .ZN(n20961) );
  OAI221_X1 U23909 ( .B1(n21170), .B2(keyinput_g14), .C1(n20962), .C2(
        keyinput_g79), .A(n20961), .ZN(n20971) );
  INV_X1 U23910 ( .A(BS16), .ZN(n20964) );
  AOI22_X1 U23911 ( .A1(n20964), .A2(keyinput_g35), .B1(n11717), .B2(
        keyinput_g118), .ZN(n20963) );
  OAI221_X1 U23912 ( .B1(n20964), .B2(keyinput_g35), .C1(n11717), .C2(
        keyinput_g118), .A(n20963), .ZN(n20970) );
  AOI22_X1 U23913 ( .A1(n20966), .A2(keyinput_g47), .B1(n21172), .B2(
        keyinput_g70), .ZN(n20965) );
  OAI221_X1 U23914 ( .B1(n20966), .B2(keyinput_g47), .C1(n21172), .C2(
        keyinput_g70), .A(n20965), .ZN(n20969) );
  INV_X1 U23915 ( .A(DATAI_11_), .ZN(n21185) );
  AOI22_X1 U23916 ( .A1(n11695), .A2(keyinput_g119), .B1(keyinput_g21), .B2(
        n21185), .ZN(n20967) );
  OAI221_X1 U23917 ( .B1(n11695), .B2(keyinput_g119), .C1(n21185), .C2(
        keyinput_g21), .A(n20967), .ZN(n20968) );
  NOR4_X1 U23918 ( .A1(n20971), .A2(n20970), .A3(n20969), .A4(n20968), .ZN(
        n20997) );
  INV_X1 U23919 ( .A(DATAI_2_), .ZN(n21167) );
  AOI22_X1 U23920 ( .A1(n20973), .A2(keyinput_g3), .B1(keyinput_g30), .B2(
        n21167), .ZN(n20972) );
  OAI221_X1 U23921 ( .B1(n20973), .B2(keyinput_g3), .C1(n21167), .C2(
        keyinput_g30), .A(n20972), .ZN(n20982) );
  AOI22_X1 U23922 ( .A1(n20975), .A2(keyinput_g103), .B1(keyinput_g49), .B2(
        n21037), .ZN(n20974) );
  OAI221_X1 U23923 ( .B1(n20975), .B2(keyinput_g103), .C1(n21037), .C2(
        keyinput_g49), .A(n20974), .ZN(n20981) );
  AOI22_X1 U23924 ( .A1(n21168), .A2(keyinput_g10), .B1(n20977), .B2(
        keyinput_g95), .ZN(n20976) );
  OAI221_X1 U23925 ( .B1(n21168), .B2(keyinput_g10), .C1(n20977), .C2(
        keyinput_g95), .A(n20976), .ZN(n20980) );
  AOI22_X1 U23926 ( .A1(n11752), .A2(keyinput_g117), .B1(keyinput_g59), .B2(
        n21036), .ZN(n20978) );
  OAI221_X1 U23927 ( .B1(n11752), .B2(keyinput_g117), .C1(n21036), .C2(
        keyinput_g59), .A(n20978), .ZN(n20979) );
  NOR4_X1 U23928 ( .A1(n20982), .A2(n20981), .A3(n20980), .A4(n20979), .ZN(
        n20996) );
  INV_X1 U23929 ( .A(DATAI_7_), .ZN(n21039) );
  AOI22_X1 U23930 ( .A1(n20984), .A2(keyinput_g78), .B1(keyinput_g25), .B2(
        n21039), .ZN(n20983) );
  OAI221_X1 U23931 ( .B1(n20984), .B2(keyinput_g78), .C1(n21039), .C2(
        keyinput_g25), .A(n20983), .ZN(n20994) );
  AOI22_X1 U23932 ( .A1(n20986), .A2(keyinput_g84), .B1(n21186), .B2(
        keyinput_g96), .ZN(n20985) );
  OAI221_X1 U23933 ( .B1(n20986), .B2(keyinput_g84), .C1(n21186), .C2(
        keyinput_g96), .A(n20985), .ZN(n20993) );
  AOI22_X1 U23934 ( .A1(n20988), .A2(keyinput_g33), .B1(n11671), .B2(
        keyinput_g120), .ZN(n20987) );
  OAI221_X1 U23935 ( .B1(n20988), .B2(keyinput_g33), .C1(n11671), .C2(
        keyinput_g120), .A(n20987), .ZN(n20992) );
  AOI22_X1 U23936 ( .A1(n20990), .A2(keyinput_g39), .B1(n11652), .B2(
        keyinput_g121), .ZN(n20989) );
  OAI221_X1 U23937 ( .B1(n20990), .B2(keyinput_g39), .C1(n11652), .C2(
        keyinput_g121), .A(n20989), .ZN(n20991) );
  NOR4_X1 U23938 ( .A1(n20994), .A2(n20993), .A3(n20992), .A4(n20991), .ZN(
        n20995) );
  NAND4_X1 U23939 ( .A1(n20998), .A2(n20997), .A3(n20996), .A4(n20995), .ZN(
        n20999) );
  NOR4_X1 U23940 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21003) );
  AOI22_X1 U23941 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(keyinput_g125), .B1(
        n21004), .B2(n21003), .ZN(n21212) );
  INV_X1 U23942 ( .A(keyinput_f125), .ZN(n21210) );
  AOI22_X1 U23943 ( .A1(n21006), .A2(keyinput_f18), .B1(keyinput_f17), .B2(
        n13439), .ZN(n21005) );
  OAI221_X1 U23944 ( .B1(n21006), .B2(keyinput_f18), .C1(n13439), .C2(
        keyinput_f17), .A(n21005), .ZN(n21019) );
  INV_X1 U23945 ( .A(DATAI_9_), .ZN(n21009) );
  AOI22_X1 U23946 ( .A1(n21009), .A2(keyinput_f23), .B1(n21008), .B2(
        keyinput_f97), .ZN(n21007) );
  OAI221_X1 U23947 ( .B1(n21009), .B2(keyinput_f23), .C1(n21008), .C2(
        keyinput_f97), .A(n21007), .ZN(n21018) );
  AOI22_X1 U23948 ( .A1(n21012), .A2(keyinput_f8), .B1(n21011), .B2(
        keyinput_f1), .ZN(n21010) );
  OAI221_X1 U23949 ( .B1(n21012), .B2(keyinput_f8), .C1(n21011), .C2(
        keyinput_f1), .A(n21010), .ZN(n21017) );
  AOI22_X1 U23950 ( .A1(n21015), .A2(keyinput_f28), .B1(keyinput_f50), .B2(
        n21014), .ZN(n21013) );
  OAI221_X1 U23951 ( .B1(n21015), .B2(keyinput_f28), .C1(n21014), .C2(
        keyinput_f50), .A(n21013), .ZN(n21016) );
  NOR4_X1 U23952 ( .A1(n21019), .A2(n21018), .A3(n21017), .A4(n21016), .ZN(
        n21208) );
  INV_X1 U23953 ( .A(DATAI_12_), .ZN(n21022) );
  INV_X1 U23954 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21021) );
  AOI22_X1 U23955 ( .A1(n21022), .A2(keyinput_f20), .B1(n21021), .B2(
        keyinput_f110), .ZN(n21020) );
  OAI221_X1 U23956 ( .B1(n21022), .B2(keyinput_f20), .C1(n21021), .C2(
        keyinput_f110), .A(n21020), .ZN(n21031) );
  AOI22_X1 U23957 ( .A1(n21024), .A2(keyinput_f85), .B1(keyinput_f61), .B2(
        n14632), .ZN(n21023) );
  OAI221_X1 U23958 ( .B1(n21024), .B2(keyinput_f85), .C1(n14632), .C2(
        keyinput_f61), .A(n21023), .ZN(n21030) );
  AOI22_X1 U23959 ( .A1(n11581), .A2(keyinput_f124), .B1(keyinput_f94), .B2(
        n21026), .ZN(n21025) );
  OAI221_X1 U23960 ( .B1(n11581), .B2(keyinput_f124), .C1(n21026), .C2(
        keyinput_f94), .A(n21025), .ZN(n21029) );
  AOI22_X1 U23961 ( .A1(n15882), .A2(keyinput_f11), .B1(n13972), .B2(
        keyinput_f112), .ZN(n21027) );
  OAI221_X1 U23962 ( .B1(n15882), .B2(keyinput_f11), .C1(n13972), .C2(
        keyinput_f112), .A(n21027), .ZN(n21028) );
  NOR4_X1 U23963 ( .A1(n21031), .A2(n21030), .A3(n21029), .A4(n21028), .ZN(
        n21207) );
  INV_X1 U23964 ( .A(READY2), .ZN(n21033) );
  AOI22_X1 U23965 ( .A1(n21034), .A2(keyinput_f31), .B1(keyinput_f37), .B2(
        n21033), .ZN(n21032) );
  OAI221_X1 U23966 ( .B1(n21034), .B2(keyinput_f31), .C1(n21033), .C2(
        keyinput_f37), .A(n21032), .ZN(n21064) );
  AOI22_X1 U23967 ( .A1(n21036), .A2(keyinput_f59), .B1(keyinput_f15), .B2(
        n15894), .ZN(n21035) );
  OAI221_X1 U23968 ( .B1(n21036), .B2(keyinput_f59), .C1(n15894), .C2(
        keyinput_f15), .A(n21035), .ZN(n21063) );
  INV_X1 U23969 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21044) );
  XNOR2_X1 U23970 ( .A(keyinput_f49), .B(n21037), .ZN(n21042) );
  AOI22_X1 U23971 ( .A1(n21040), .A2(keyinput_f57), .B1(keyinput_f25), .B2(
        n21039), .ZN(n21038) );
  OAI221_X1 U23972 ( .B1(n21040), .B2(keyinput_f57), .C1(n21039), .C2(
        keyinput_f25), .A(n21038), .ZN(n21041) );
  AOI211_X1 U23973 ( .C1(n21044), .C2(keyinput_f116), .A(n21042), .B(n21041), 
        .ZN(n21043) );
  OAI21_X1 U23974 ( .B1(n21044), .B2(keyinput_f116), .A(n21043), .ZN(n21062)
         );
  OAI22_X1 U23975 ( .A1(n21047), .A2(keyinput_f90), .B1(n21046), .B2(
        keyinput_f56), .ZN(n21045) );
  AOI221_X1 U23976 ( .B1(n21047), .B2(keyinput_f90), .C1(keyinput_f56), .C2(
        n21046), .A(n21045), .ZN(n21060) );
  OAI22_X1 U23977 ( .A1(n21050), .A2(keyinput_f99), .B1(n21049), .B2(
        keyinput_f40), .ZN(n21048) );
  AOI221_X1 U23978 ( .B1(n21050), .B2(keyinput_f99), .C1(keyinput_f40), .C2(
        n21049), .A(n21048), .ZN(n21059) );
  OAI22_X1 U23979 ( .A1(n21053), .A2(keyinput_f72), .B1(n21052), .B2(
        keyinput_f34), .ZN(n21051) );
  AOI221_X1 U23980 ( .B1(n21053), .B2(keyinput_f72), .C1(keyinput_f34), .C2(
        n21052), .A(n21051), .ZN(n21058) );
  INV_X1 U23981 ( .A(DATAI_8_), .ZN(n21055) );
  OAI22_X1 U23982 ( .A1(n21056), .A2(keyinput_f114), .B1(n21055), .B2(
        keyinput_f24), .ZN(n21054) );
  AOI221_X1 U23983 ( .B1(n21056), .B2(keyinput_f114), .C1(keyinput_f24), .C2(
        n21055), .A(n21054), .ZN(n21057) );
  NAND4_X1 U23984 ( .A1(n21060), .A2(n21059), .A3(n21058), .A4(n21057), .ZN(
        n21061) );
  NOR4_X1 U23985 ( .A1(n21064), .A2(n21063), .A3(n21062), .A4(n21061), .ZN(
        n21206) );
  OAI22_X1 U23986 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(keyinput_f78), .B1(
        keyinput_f42), .B2(P1_D_C_N_REG_SCAN_IN), .ZN(n21065) );
  AOI221_X1 U23987 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(keyinput_f78), .C1(
        P1_D_C_N_REG_SCAN_IN), .C2(keyinput_f42), .A(n21065), .ZN(n21072) );
  OAI22_X1 U23988 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(keyinput_f113), .B1(
        keyinput_f12), .B2(DATAI_20_), .ZN(n21066) );
  AOI221_X1 U23989 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(keyinput_f113), .C1(
        DATAI_20_), .C2(keyinput_f12), .A(n21066), .ZN(n21071) );
  OAI22_X1 U23990 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_f88), .B1(
        keyinput_f63), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n21067) );
  AOI221_X1 U23991 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_f88), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_f63), .A(n21067), .ZN(n21070)
         );
  OAI22_X1 U23992 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(keyinput_f84), .B1(
        DATAI_3_), .B2(keyinput_f29), .ZN(n21068) );
  AOI221_X1 U23993 ( .B1(P1_EBX_REG_31__SCAN_IN), .B2(keyinput_f84), .C1(
        keyinput_f29), .C2(DATAI_3_), .A(n21068), .ZN(n21069) );
  NAND4_X1 U23994 ( .A1(n21072), .A2(n21071), .A3(n21070), .A4(n21069), .ZN(
        n21204) );
  OAI22_X1 U23995 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(keyinput_f109), .B1(
        keyinput_f79), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n21073) );
  AOI221_X1 U23996 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(keyinput_f109), .C1(
        P1_REIP_REG_4__SCAN_IN), .C2(keyinput_f79), .A(n21073), .ZN(n21099) );
  OAI22_X1 U23997 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_f104), .B1(
        keyinput_f80), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n21074) );
  AOI221_X1 U23998 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_f104), .C1(
        P1_REIP_REG_3__SCAN_IN), .C2(keyinput_f80), .A(n21074), .ZN(n21077) );
  OAI22_X1 U23999 ( .A1(P1_EBX_REG_29__SCAN_IN), .A2(keyinput_f86), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(keyinput_f75), .ZN(n21075) );
  AOI221_X1 U24000 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(keyinput_f86), .C1(
        keyinput_f75), .C2(P1_REIP_REG_8__SCAN_IN), .A(n21075), .ZN(n21076) );
  OAI211_X1 U24001 ( .C1(n21079), .C2(keyinput_f38), .A(n21077), .B(n21076), 
        .ZN(n21078) );
  AOI21_X1 U24002 ( .B1(n21079), .B2(keyinput_f38), .A(n21078), .ZN(n21098) );
  AOI22_X1 U24003 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(keyinput_f111), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(keyinput_f103), .ZN(n21080) );
  OAI221_X1 U24004 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(keyinput_f111), .C1(
        P1_EBX_REG_12__SCAN_IN), .C2(keyinput_f103), .A(n21080), .ZN(n21087)
         );
  AOI22_X1 U24005 ( .A1(DATAI_28_), .A2(keyinput_f4), .B1(
        P1_EBX_REG_13__SCAN_IN), .B2(keyinput_f102), .ZN(n21081) );
  OAI221_X1 U24006 ( .B1(DATAI_28_), .B2(keyinput_f4), .C1(
        P1_EBX_REG_13__SCAN_IN), .C2(keyinput_f102), .A(n21081), .ZN(n21086)
         );
  AOI22_X1 U24007 ( .A1(DATAI_6_), .A2(keyinput_f26), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(keyinput_f82), .ZN(n21082) );
  OAI221_X1 U24008 ( .B1(DATAI_6_), .B2(keyinput_f26), .C1(
        P1_REIP_REG_1__SCAN_IN), .C2(keyinput_f82), .A(n21082), .ZN(n21085) );
  AOI22_X1 U24009 ( .A1(keyinput_f51), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        DATAI_10_), .B2(keyinput_f22), .ZN(n21083) );
  OAI221_X1 U24010 ( .B1(keyinput_f51), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), 
        .C1(DATAI_10_), .C2(keyinput_f22), .A(n21083), .ZN(n21084) );
  NOR4_X1 U24011 ( .A1(n21087), .A2(n21086), .A3(n21085), .A4(n21084), .ZN(
        n21097) );
  AOI22_X1 U24012 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_f39), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(keyinput_f67), .ZN(n21088) );
  OAI221_X1 U24013 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_f39), .C1(
        P1_REIP_REG_16__SCAN_IN), .C2(keyinput_f67), .A(n21088), .ZN(n21095)
         );
  AOI22_X1 U24014 ( .A1(keyinput_f33), .A2(HOLD), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(keyinput_f100), .ZN(n21089) );
  OAI221_X1 U24015 ( .B1(keyinput_f33), .B2(HOLD), .C1(P1_EBX_REG_15__SCAN_IN), 
        .C2(keyinput_f100), .A(n21089), .ZN(n21094) );
  AOI22_X1 U24016 ( .A1(DATAI_0_), .A2(keyinput_f32), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_f62), .ZN(n21090) );
  OAI221_X1 U24017 ( .B1(DATAI_0_), .B2(keyinput_f32), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_f62), .A(n21090), .ZN(n21093)
         );
  AOI22_X1 U24018 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_f53), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(keyinput_f101), .ZN(n21091) );
  OAI221_X1 U24019 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .C1(
        P1_EBX_REG_14__SCAN_IN), .C2(keyinput_f101), .A(n21091), .ZN(n21092)
         );
  NOR4_X1 U24020 ( .A1(n21095), .A2(n21094), .A3(n21093), .A4(n21092), .ZN(
        n21096) );
  NAND4_X1 U24021 ( .A1(n21099), .A2(n21098), .A3(n21097), .A4(n21096), .ZN(
        n21203) );
  AOI22_X1 U24022 ( .A1(keyinput_f35), .A2(BS16), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(keyinput_f87), .ZN(n21100) );
  OAI221_X1 U24023 ( .B1(keyinput_f35), .B2(BS16), .C1(P1_EBX_REG_28__SCAN_IN), 
        .C2(keyinput_f87), .A(n21100), .ZN(n21107) );
  AOI22_X1 U24024 ( .A1(keyinput_f47), .A2(P1_W_R_N_REG_SCAN_IN), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(keyinput_f74), .ZN(n21101) );
  OAI221_X1 U24025 ( .B1(keyinput_f47), .B2(P1_W_R_N_REG_SCAN_IN), .C1(
        P1_REIP_REG_9__SCAN_IN), .C2(keyinput_f74), .A(n21101), .ZN(n21106) );
  AOI22_X1 U24026 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_f46), .B1(
        P1_EBX_REG_17__SCAN_IN), .B2(keyinput_f98), .ZN(n21102) );
  OAI221_X1 U24027 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .C1(
        P1_EBX_REG_17__SCAN_IN), .C2(keyinput_f98), .A(n21102), .ZN(n21105) );
  AOI22_X1 U24028 ( .A1(P1_EBX_REG_10__SCAN_IN), .A2(keyinput_f105), .B1(
        P1_EBX_REG_26__SCAN_IN), .B2(keyinput_f89), .ZN(n21103) );
  OAI221_X1 U24029 ( .B1(P1_EBX_REG_10__SCAN_IN), .B2(keyinput_f105), .C1(
        P1_EBX_REG_26__SCAN_IN), .C2(keyinput_f89), .A(n21103), .ZN(n21104) );
  NOR4_X1 U24030 ( .A1(n21107), .A2(n21106), .A3(n21105), .A4(n21104), .ZN(
        n21136) );
  AOI22_X1 U24031 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(keyinput_f106), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(keyinput_f107), .ZN(n21108) );
  OAI221_X1 U24032 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(keyinput_f106), .C1(
        P1_EBX_REG_8__SCAN_IN), .C2(keyinput_f107), .A(n21108), .ZN(n21115) );
  AOI22_X1 U24033 ( .A1(P1_EBX_REG_23__SCAN_IN), .A2(keyinput_f92), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(keyinput_f123), .ZN(n21109) );
  OAI221_X1 U24034 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(keyinput_f92), .C1(
        P1_EAX_REG_24__SCAN_IN), .C2(keyinput_f123), .A(n21109), .ZN(n21114)
         );
  AOI22_X1 U24035 ( .A1(DATAI_13_), .A2(keyinput_f19), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(keyinput_f121), .ZN(n21110) );
  OAI221_X1 U24036 ( .B1(DATAI_13_), .B2(keyinput_f19), .C1(
        P1_EAX_REG_26__SCAN_IN), .C2(keyinput_f121), .A(n21110), .ZN(n21113)
         );
  AOI22_X1 U24037 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(keyinput_f83), .B1(
        DATAI_29_), .B2(keyinput_f3), .ZN(n21111) );
  OAI221_X1 U24038 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(keyinput_f83), .C1(
        DATAI_29_), .C2(keyinput_f3), .A(n21111), .ZN(n21112) );
  NOR4_X1 U24039 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21135) );
  AOI22_X1 U24040 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_f45), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(keyinput_f65), .ZN(n21116) );
  OAI221_X1 U24041 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_f45), .C1(
        P1_REIP_REG_18__SCAN_IN), .C2(keyinput_f65), .A(n21116), .ZN(n21123)
         );
  AOI22_X1 U24042 ( .A1(DATAI_26_), .A2(keyinput_f6), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_f54), .ZN(n21117) );
  OAI221_X1 U24043 ( .B1(DATAI_26_), .B2(keyinput_f6), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_f54), .A(n21117), .ZN(n21122)
         );
  AOI22_X1 U24044 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(keyinput_f66), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_f118), .ZN(n21118) );
  OAI221_X1 U24045 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(keyinput_f66), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_f118), .A(n21118), .ZN(n21121)
         );
  AOI22_X1 U24046 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(keyinput_f73), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(keyinput_f76), .ZN(n21119) );
  OAI221_X1 U24047 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(keyinput_f73), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(keyinput_f76), .A(n21119), .ZN(n21120) );
  NOR4_X1 U24048 ( .A1(n21123), .A2(n21122), .A3(n21121), .A4(n21120), .ZN(
        n21134) );
  AOI22_X1 U24049 ( .A1(READY1), .A2(keyinput_f36), .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_f120), .ZN(n21124) );
  OAI221_X1 U24050 ( .B1(READY1), .B2(keyinput_f36), .C1(
        P1_EAX_REG_27__SCAN_IN), .C2(keyinput_f120), .A(n21124), .ZN(n21132)
         );
  AOI22_X1 U24051 ( .A1(DATAI_19_), .A2(keyinput_f13), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .ZN(n21125) );
  OAI221_X1 U24052 ( .B1(DATAI_19_), .B2(keyinput_f13), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_f58), .A(n21125), .ZN(n21131)
         );
  AOI22_X1 U24053 ( .A1(P1_EBX_REG_20__SCAN_IN), .A2(keyinput_f95), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(keyinput_f93), .ZN(n21126) );
  OAI221_X1 U24054 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(keyinput_f95), .C1(
        P1_EBX_REG_22__SCAN_IN), .C2(keyinput_f93), .A(n21126), .ZN(n21130) );
  AOI22_X1 U24055 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(keyinput_f77), .B1(n21128), .B2(keyinput_f91), .ZN(n21127) );
  OAI221_X1 U24056 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(keyinput_f77), .C1(
        n21128), .C2(keyinput_f91), .A(n21127), .ZN(n21129) );
  NOR4_X1 U24057 ( .A1(n21132), .A2(n21131), .A3(n21130), .A4(n21129), .ZN(
        n21133) );
  NAND4_X1 U24058 ( .A1(n21136), .A2(n21135), .A3(n21134), .A4(n21133), .ZN(
        n21202) );
  AOI22_X1 U24059 ( .A1(n14016), .A2(keyinput_f115), .B1(keyinput_f68), .B2(
        n21138), .ZN(n21137) );
  OAI221_X1 U24060 ( .B1(n14016), .B2(keyinput_f115), .C1(n21138), .C2(
        keyinput_f68), .A(n21137), .ZN(n21151) );
  AOI22_X1 U24061 ( .A1(n21141), .A2(keyinput_f122), .B1(n21140), .B2(
        keyinput_f44), .ZN(n21139) );
  OAI221_X1 U24062 ( .B1(n21141), .B2(keyinput_f122), .C1(n21140), .C2(
        keyinput_f44), .A(n21139), .ZN(n21150) );
  INV_X1 U24063 ( .A(keyinput_f48), .ZN(n21143) );
  AOI22_X1 U24064 ( .A1(n21144), .A2(keyinput_f2), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(n21143), .ZN(n21142) );
  OAI221_X1 U24065 ( .B1(n21144), .B2(keyinput_f2), .C1(n21143), .C2(
        P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21142), .ZN(n21149) );
  INV_X1 U24066 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21146) );
  AOI22_X1 U24067 ( .A1(n21147), .A2(keyinput_f108), .B1(keyinput_f55), .B2(
        n21146), .ZN(n21145) );
  OAI221_X1 U24068 ( .B1(n21147), .B2(keyinput_f108), .C1(n21146), .C2(
        keyinput_f55), .A(n21145), .ZN(n21148) );
  NOR4_X1 U24069 ( .A1(n21151), .A2(n21150), .A3(n21149), .A4(n21148), .ZN(
        n21200) );
  AOI22_X1 U24070 ( .A1(n21154), .A2(keyinput_f7), .B1(n21153), .B2(
        keyinput_f5), .ZN(n21152) );
  OAI221_X1 U24071 ( .B1(n21154), .B2(keyinput_f7), .C1(n21153), .C2(
        keyinput_f5), .A(n21152), .ZN(n21165) );
  AOI22_X1 U24072 ( .A1(n21157), .A2(keyinput_f64), .B1(keyinput_f41), .B2(
        n21156), .ZN(n21155) );
  OAI221_X1 U24073 ( .B1(n21157), .B2(keyinput_f64), .C1(n21156), .C2(
        keyinput_f41), .A(n21155), .ZN(n21164) );
  AOI22_X1 U24074 ( .A1(n21159), .A2(keyinput_f60), .B1(keyinput_f69), .B2(
        n14256), .ZN(n21158) );
  OAI221_X1 U24075 ( .B1(n21159), .B2(keyinput_f60), .C1(n14256), .C2(
        keyinput_f69), .A(n21158), .ZN(n21163) );
  AOI22_X1 U24076 ( .A1(n11752), .A2(keyinput_f117), .B1(keyinput_f27), .B2(
        n21161), .ZN(n21160) );
  OAI221_X1 U24077 ( .B1(n11752), .B2(keyinput_f117), .C1(n21161), .C2(
        keyinput_f27), .A(n21160), .ZN(n21162) );
  NOR4_X1 U24078 ( .A1(n21165), .A2(n21164), .A3(n21163), .A4(n21162), .ZN(
        n21199) );
  AOI22_X1 U24079 ( .A1(n21168), .A2(keyinput_f10), .B1(keyinput_f30), .B2(
        n21167), .ZN(n21166) );
  OAI221_X1 U24080 ( .B1(n21168), .B2(keyinput_f10), .C1(n21167), .C2(
        keyinput_f30), .A(n21166), .ZN(n21180) );
  AOI22_X1 U24081 ( .A1(n11695), .A2(keyinput_f119), .B1(keyinput_f14), .B2(
        n21170), .ZN(n21169) );
  OAI221_X1 U24082 ( .B1(n11695), .B2(keyinput_f119), .C1(n21170), .C2(
        keyinput_f14), .A(n21169), .ZN(n21179) );
  AOI22_X1 U24083 ( .A1(n21173), .A2(keyinput_f71), .B1(n21172), .B2(
        keyinput_f70), .ZN(n21171) );
  OAI221_X1 U24084 ( .B1(n21173), .B2(keyinput_f71), .C1(n21172), .C2(
        keyinput_f70), .A(n21171), .ZN(n21178) );
  AOI22_X1 U24085 ( .A1(n21176), .A2(keyinput_f126), .B1(keyinput_f43), .B2(
        n21175), .ZN(n21174) );
  OAI221_X1 U24086 ( .B1(n21176), .B2(keyinput_f126), .C1(n21175), .C2(
        keyinput_f43), .A(n21174), .ZN(n21177) );
  NOR4_X1 U24087 ( .A1(n21180), .A2(n21179), .A3(n21178), .A4(n21177), .ZN(
        n21198) );
  AOI22_X1 U24088 ( .A1(n21183), .A2(keyinput_f52), .B1(keyinput_f16), .B2(
        n21182), .ZN(n21181) );
  OAI221_X1 U24089 ( .B1(n21183), .B2(keyinput_f52), .C1(n21182), .C2(
        keyinput_f16), .A(n21181), .ZN(n21196) );
  AOI22_X1 U24090 ( .A1(n21186), .A2(keyinput_f96), .B1(keyinput_f21), .B2(
        n21185), .ZN(n21184) );
  OAI221_X1 U24091 ( .B1(n21186), .B2(keyinput_f96), .C1(n21185), .C2(
        keyinput_f21), .A(n21184), .ZN(n21195) );
  AOI22_X1 U24092 ( .A1(n21189), .A2(keyinput_f9), .B1(keyinput_f0), .B2(
        n21188), .ZN(n21187) );
  OAI221_X1 U24093 ( .B1(n21189), .B2(keyinput_f9), .C1(n21188), .C2(
        keyinput_f0), .A(n21187), .ZN(n21194) );
  AOI22_X1 U24094 ( .A1(n21192), .A2(keyinput_f127), .B1(keyinput_f81), .B2(
        n21191), .ZN(n21190) );
  OAI221_X1 U24095 ( .B1(n21192), .B2(keyinput_f127), .C1(n21191), .C2(
        keyinput_f81), .A(n21190), .ZN(n21193) );
  NOR4_X1 U24096 ( .A1(n21196), .A2(n21195), .A3(n21194), .A4(n21193), .ZN(
        n21197) );
  NAND4_X1 U24097 ( .A1(n21200), .A2(n21199), .A3(n21198), .A4(n21197), .ZN(
        n21201) );
  NOR4_X1 U24098 ( .A1(n21204), .A2(n21203), .A3(n21202), .A4(n21201), .ZN(
        n21205) );
  NAND4_X1 U24099 ( .A1(n21208), .A2(n21207), .A3(n21206), .A4(n21205), .ZN(
        n21209) );
  OAI221_X1 U24100 ( .B1(P1_EAX_REG_22__SCAN_IN), .B2(n21210), .C1(n11553), 
        .C2(keyinput_f125), .A(n21209), .ZN(n21211) );
  OAI211_X1 U24101 ( .C1(P1_EAX_REG_22__SCAN_IN), .C2(keyinput_g125), .A(
        n21212), .B(n21211), .ZN(n21213) );
  XOR2_X1 U24102 ( .A(n21214), .B(n21213), .Z(U355) );
  AND2_X1 U13912 ( .A1(n13737), .A2(n10921), .ZN(n11115) );
  CLKBUF_X2 U12502 ( .A(n10431), .Z(n13446) );
  INV_X2 U11269 ( .A(n12697), .ZN(n17195) );
  INV_X1 U15683 ( .A(n10240), .ZN(n17235) );
  NAND2_X2 U11274 ( .A1(n10938), .A2(n10937), .ZN(n11031) );
  INV_X4 U15677 ( .A(n17199), .ZN(n17223) );
  CLKBUF_X1 U11255 ( .A(n10992), .Z(n11741) );
  CLKBUF_X1 U11279 ( .A(n10972), .Z(n11569) );
  AND2_X1 U11280 ( .A1(n9814), .A2(n12330), .ZN(n12319) );
  CLKBUF_X2 U11296 ( .A(n10335), .Z(n10593) );
  NAND2_X1 U11303 ( .A1(n20294), .A2(n11155), .ZN(n11158) );
  NOR2_X1 U11316 ( .A1(n11047), .A2(n11009), .ZN(n13253) );
  CLKBUF_X1 U11353 ( .A(n20170), .Z(n9812) );
  CLKBUF_X1 U11359 ( .A(n11043), .Z(n20202) );
  INV_X1 U11375 ( .A(n10587), .ZN(n19277) );
  CLKBUF_X1 U11605 ( .A(n10257), .Z(n17193) );
  CLKBUF_X1 U12223 ( .A(n11067), .Z(n15708) );
  INV_X1 U12405 ( .A(n18244), .ZN(n18885) );
  NAND2_X1 U12441 ( .A1(n18668), .A2(n18878), .ZN(n16532) );
  CLKBUF_X1 U12540 ( .A(n16513), .Z(n16521) );
  INV_X2 U12728 ( .A(n18879), .ZN(n18720) );
  CLKBUF_X1 U12781 ( .A(n17528), .Z(n17536) );
endmodule

