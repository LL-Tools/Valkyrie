

module b15_C_SARLock_k_64_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2963, n2964, n2965, n2966, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671;

  OR2_X1 U3412 ( .A1(n5559), .A2(n3048), .ZN(n3045) );
  NAND2_X1 U3413 ( .A1(n3448), .A2(n3447), .ZN(n3475) );
  NOR2_X1 U3414 ( .A1(n3429), .A2(n3410), .ZN(n3421) );
  OR2_X1 U3415 ( .A1(n3612), .A2(n5373), .ZN(n3601) );
  NAND2_X2 U3416 ( .A1(n4590), .A2(n3224), .ZN(n3612) );
  CLKBUF_X2 U3418 ( .A(n3195), .Z(n3390) );
  INV_X2 U3419 ( .A(n3222), .ZN(n3224) );
  CLKBUF_X2 U3420 ( .A(n3188), .Z(n4169) );
  INV_X1 U3421 ( .A(n4368), .ZN(n3155) );
  AND4_X1 U3422 ( .A1(n3122), .A2(n3121), .A3(n3120), .A4(n3119), .ZN(n4368)
         );
  INV_X1 U3423 ( .A(n3231), .ZN(n4612) );
  AND2_X1 U3424 ( .A1(n4538), .A2(n4553), .ZN(n3195) );
  AND2_X2 U3425 ( .A1(n5276), .A2(n4537), .ZN(n3186) );
  AND2_X2 U3426 ( .A1(n4538), .A2(n5274), .ZN(n3189) );
  INV_X1 U3427 ( .A(n3601), .ZN(n3609) );
  NAND2_X1 U3428 ( .A1(n3389), .A2(n6192), .ZN(n3429) );
  AND2_X1 U3429 ( .A1(n3166), .A2(n3219), .ZN(n3167) );
  AND3_X1 U3430 ( .A1(n4590), .A2(n4585), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3505) );
  NAND2_X1 U3431 ( .A1(n4369), .A2(n2992), .ZN(n3606) );
  XNOR2_X1 U3432 ( .A(n3429), .B(n3432), .ZN(n3737) );
  AND4_X1 U3433 ( .A1(n3106), .A2(n3105), .A3(n3104), .A4(n3103), .ZN(n3122)
         );
  AND4_X1 U3434 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n4370)
         );
  AND2_X1 U3435 ( .A1(n4269), .A2(n3222), .ZN(n5082) );
  INV_X1 U3436 ( .A(n5928), .ZN(n5952) );
  OAI21_X1 U3437 ( .B1(n5315), .B2(n4214), .A(n4230), .ZN(n4233) );
  AND2_X4 U3438 ( .A1(n4537), .A2(n5274), .ZN(n3194) );
  AND2_X4 U3439 ( .A1(n5292), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4537)
         );
  NOR2_X2 U3440 ( .A1(n5547), .A2(n5540), .ZN(n5523) );
  NAND2_X2 U3441 ( .A1(n5549), .A2(n5548), .ZN(n5547) );
  OAI21_X2 U3442 ( .B1(n4575), .B2(n3472), .A(n3328), .ZN(n6031) );
  NAND2_X1 U3443 ( .A1(n6015), .A2(n6014), .ZN(n6013) );
  NAND2_X1 U3444 ( .A1(n4848), .A2(n3428), .ZN(n6015) );
  NAND2_X2 U34450 ( .A1(n3475), .A2(n3474), .ZN(n5581) );
  AOI21_X1 U34470 ( .B1(n3330), .B2(n3329), .A(n3471), .ZN(n3342) );
  INV_X1 U34480 ( .A(n3612), .ZN(n4422) );
  AND2_X2 U3449 ( .A1(n3068), .A2(n3067), .ZN(n3222) );
  INV_X1 U3450 ( .A(n4370), .ZN(n4585) );
  AND4_X1 U34510 ( .A1(n3096), .A2(n3095), .A3(n3094), .A4(n3093), .ZN(n3102)
         );
  AND4_X1 U34520 ( .A1(n3100), .A2(n3099), .A3(n3098), .A4(n3097), .ZN(n3101)
         );
  BUF_X2 U34530 ( .A(n3189), .Z(n4188) );
  BUF_X2 U3454 ( .A(n3186), .Z(n4168) );
  CLKBUF_X2 U34550 ( .A(n4081), .Z(n3366) );
  BUF_X2 U34560 ( .A(n3286), .Z(n2964) );
  CLKBUF_X2 U3457 ( .A(n3280), .Z(n4193) );
  CLKBUF_X2 U3458 ( .A(n3187), .Z(n4195) );
  CLKBUF_X2 U34590 ( .A(n3198), .Z(n4194) );
  INV_X2 U34600 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5292) );
  INV_X2 U34610 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4539) );
  INV_X2 U34620 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3075) );
  OAI21_X1 U34630 ( .B1(n4308), .B2(n5805), .A(n4307), .ZN(n3003) );
  XNOR2_X1 U34640 ( .A(n4221), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4308)
         );
  NAND2_X1 U34650 ( .A1(n4220), .A2(n4219), .ZN(n4221) );
  NOR2_X1 U3466 ( .A1(n5493), .A2(n5595), .ZN(n4216) );
  NOR3_X1 U3467 ( .A1(n4217), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5581), 
        .ZN(n5494) );
  NAND2_X1 U34680 ( .A1(n3045), .A2(n3043), .ZN(n5493) );
  NAND2_X1 U34690 ( .A1(n3035), .A2(n5186), .ZN(n5788) );
  OR2_X1 U34700 ( .A1(n4864), .A2(n2974), .ZN(n3039) );
  AND2_X1 U34710 ( .A1(n4569), .A2(n3748), .ZN(n3013) );
  INV_X1 U34720 ( .A(n5581), .ZN(n5776) );
  XNOR2_X1 U34730 ( .A(n3475), .B(n3462), .ZN(n3752) );
  INV_X1 U34740 ( .A(n3450), .ZN(n3448) );
  NOR2_X1 U3475 ( .A1(n4953), .A2(n4914), .ZN(n6170) );
  NAND2_X1 U3476 ( .A1(n3385), .A2(n3384), .ZN(n3386) );
  CLKBUF_X1 U3477 ( .A(n4576), .Z(n4577) );
  NAND2_X2 U3478 ( .A1(n3379), .A2(n3378), .ZN(n6192) );
  OAI21_X1 U3479 ( .B1(n4564), .B2(n3472), .A(n3337), .ZN(n4346) );
  NAND2_X1 U3481 ( .A1(n4533), .A2(n6379), .ZN(n3379) );
  XNOR2_X1 U3482 ( .A(n4554), .B(n4555), .ZN(n4533) );
  NAND2_X1 U3483 ( .A1(n3319), .A2(n3318), .ZN(n3343) );
  XNOR2_X1 U3484 ( .A(n3266), .B(n3265), .ZN(n3322) );
  NAND2_X1 U3485 ( .A1(n5458), .A2(n4502), .ZN(n5760) );
  NAND2_X1 U3486 ( .A1(n3267), .A2(n3268), .ZN(n3314) );
  NAND2_X1 U3487 ( .A1(n3215), .A2(n3214), .ZN(n3267) );
  NAND3_X1 U3488 ( .A1(n3247), .A2(n3246), .A3(n3245), .ZN(n3313) );
  AND2_X1 U3489 ( .A1(n4415), .A2(n4590), .ZN(n4326) );
  NAND2_X1 U3490 ( .A1(n3154), .A2(n3217), .ZN(n3168) );
  AND4_X1 U3491 ( .A1(n3584), .A2(n4542), .A3(n3221), .A4(n3220), .ZN(n3228)
         );
  AND2_X1 U3492 ( .A1(n3234), .A2(n3233), .ZN(n4415) );
  NOR2_X1 U3493 ( .A1(n4413), .A2(n4500), .ZN(n3678) );
  CLKBUF_X3 U3494 ( .A(n3581), .Z(n5373) );
  AND2_X1 U3495 ( .A1(n4603), .A2(n3224), .ZN(n3581) );
  OR2_X1 U3496 ( .A1(n3508), .A2(n4590), .ZN(n3229) );
  AND2_X2 U3497 ( .A1(n3222), .A2(n4590), .ZN(n4351) );
  OR2_X1 U3498 ( .A1(n3292), .A2(n3291), .ZN(n3466) );
  OR2_X1 U3499 ( .A1(n3279), .A2(n3278), .ZN(n3346) );
  NAND4_X2 U3500 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n4590)
         );
  NAND2_X2 U3501 ( .A1(n3165), .A2(n3164), .ZN(n4603) );
  AND4_X1 U3502 ( .A1(n3114), .A2(n3113), .A3(n3112), .A4(n3111), .ZN(n3120)
         );
  AND4_X1 U3503 ( .A1(n3074), .A2(n3073), .A3(n3072), .A4(n3071), .ZN(n3092)
         );
  AND4_X1 U3504 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3067)
         );
  AND2_X1 U3505 ( .A1(n2978), .A2(n3163), .ZN(n3164) );
  AND4_X1 U3506 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3206)
         );
  AND4_X1 U3507 ( .A1(n3159), .A2(n3158), .A3(n3157), .A4(n3156), .ZN(n3165)
         );
  AND4_X1 U3508 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3203)
         );
  AND4_X1 U3509 ( .A1(n3083), .A2(n3082), .A3(n3081), .A4(n3080), .ZN(n3090)
         );
  AND4_X1 U3510 ( .A1(n3110), .A2(n3109), .A3(n3108), .A4(n3107), .ZN(n3121)
         );
  AND4_X1 U3511 ( .A1(n3079), .A2(n3078), .A3(n3077), .A4(n3076), .ZN(n3091)
         );
  AND4_X1 U3512 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3152)
         );
  AND4_X1 U3513 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3204)
         );
  AND4_X1 U3514 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3151)
         );
  AND4_X1 U3515 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3153)
         );
  AND4_X1 U3516 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3150)
         );
  AND4_X1 U3517 ( .A1(n3118), .A2(n3117), .A3(n3116), .A4(n3115), .ZN(n3119)
         );
  AND4_X1 U3518 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3205)
         );
  BUF_X2 U3519 ( .A(n3197), .Z(n4196) );
  BUF_X2 U3520 ( .A(n3257), .Z(n4186) );
  BUF_X2 U3521 ( .A(n3269), .Z(n4541) );
  INV_X2 U3522 ( .A(n5579), .ZN(n2963) );
  BUF_X2 U3523 ( .A(n3196), .Z(n4187) );
  AND2_X2 U3524 ( .A1(n4537), .A2(n4553), .ZN(n3196) );
  AND2_X2 U3525 ( .A1(n5276), .A2(n4551), .ZN(n4081) );
  AND2_X2 U3526 ( .A1(n4537), .A2(n4521), .ZN(n3257) );
  NOR2_X2 U3527 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3084) );
  AND2_X2 U3528 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4521) );
  OR2_X2 U3529 ( .A1(n4233), .A2(n5579), .ZN(n2975) );
  BUF_X2 U3530 ( .A(n4213), .Z(n5315) );
  AOI22_X2 U3531 ( .A1(n3495), .A2(n5553), .B1(n5776), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5549) );
  NOR2_X2 U3532 ( .A1(n5560), .A2(n3494), .ZN(n3495) );
  AND2_X2 U3533 ( .A1(n4539), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4538)
         );
  XNOR2_X1 U3534 ( .A(n3344), .B(n3343), .ZN(n4576) );
  AND2_X1 U3535 ( .A1(n4603), .A2(n4368), .ZN(n3347) );
  NAND2_X1 U3536 ( .A1(n3322), .A2(n3321), .ZN(n3388) );
  AND2_X4 U3537 ( .A1(n3075), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5274)
         );
  NOR2_X2 U3538 ( .A1(n3034), .A2(n3229), .ZN(n3555) );
  AND2_X2 U3539 ( .A1(n5276), .A2(n4538), .ZN(n3285) );
  NAND2_X2 U3540 ( .A1(n3388), .A2(n3325), .ZN(n4575) );
  NAND2_X1 U3541 ( .A1(n3062), .A2(n2971), .ZN(n5179) );
  NAND2_X2 U3542 ( .A1(n5788), .A2(n5787), .ZN(n3487) );
  NAND2_X4 U3543 ( .A1(n3102), .A2(n3101), .ZN(n3207) );
  NOR2_X4 U3544 ( .A1(n5198), .A2(n5237), .ZN(n5238) );
  NAND2_X2 U3545 ( .A1(n5200), .A2(n5199), .ZN(n5198) );
  NOR2_X2 U3546 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n5559), .ZN(n5560)
         );
  NAND2_X2 U3547 ( .A1(n3492), .A2(n3491), .ZN(n5559) );
  AND2_X1 U3548 ( .A1(n5276), .A2(n4551), .ZN(n2965) );
  AND2_X1 U3549 ( .A1(n4538), .A2(n4553), .ZN(n2966) );
  XNOR2_X2 U3551 ( .A(n3388), .B(n6192), .ZN(n3717) );
  INV_X1 U3552 ( .A(n4342), .ZN(n3029) );
  INV_X1 U3553 ( .A(n5405), .ZN(n4122) );
  OR2_X1 U3554 ( .A1(n5570), .A2(n3489), .ZN(n3057) );
  NAND2_X1 U3555 ( .A1(n5115), .A2(n5113), .ZN(n3062) );
  NAND2_X1 U3556 ( .A1(n4576), .A2(n3814), .ZN(n3032) );
  INV_X1 U3557 ( .A(n3702), .ZN(n3031) );
  AOI21_X1 U3558 ( .B1(n4342), .B2(n3028), .A(n2972), .ZN(n3027) );
  OAI21_X1 U3559 ( .B1(n3030), .B2(n6285), .A(n3029), .ZN(n3024) );
  NOR2_X1 U3560 ( .A1(n3044), .A2(n5509), .ZN(n3043) );
  INV_X1 U3561 ( .A(n3046), .ZN(n3044) );
  NAND2_X1 U3562 ( .A1(n3010), .A2(n3331), .ZN(n3330) );
  NAND2_X1 U3563 ( .A1(n3434), .A2(n3433), .ZN(n3450) );
  AND2_X1 U3564 ( .A1(n3432), .A2(n3431), .ZN(n3433) );
  OR2_X1 U3565 ( .A1(n3307), .A2(n3306), .ZN(n3345) );
  NAND2_X1 U3566 ( .A1(n2970), .A2(n4585), .ZN(n3217) );
  INV_X1 U3567 ( .A(n5355), .ZN(n4005) );
  NOR2_X1 U3568 ( .A1(n3063), .A2(n3019), .ZN(n3018) );
  INV_X1 U3569 ( .A(n5384), .ZN(n3019) );
  INV_X1 U3570 ( .A(n4662), .ZN(n3015) );
  INV_X1 U3571 ( .A(n3033), .ZN(n3030) );
  AND2_X1 U3572 ( .A1(n5519), .A2(n2981), .ZN(n3049) );
  NAND2_X1 U3573 ( .A1(n2985), .A2(n5220), .ZN(n3054) );
  NAND2_X1 U3574 ( .A1(n2994), .A2(n4573), .ZN(n2993) );
  INV_X1 U3575 ( .A(n2995), .ZN(n2994) );
  INV_X1 U3576 ( .A(n4269), .ZN(n2992) );
  OR2_X1 U3577 ( .A1(n3263), .A2(n3262), .ZN(n3264) );
  NAND2_X1 U3578 ( .A1(n4370), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U3579 ( .A1(n3061), .A2(n6379), .ZN(n3059) );
  INV_X1 U3580 ( .A(n3217), .ZN(n3554) );
  NAND2_X1 U3581 ( .A1(n3363), .A2(n3362), .ZN(n4555) );
  NAND2_X1 U3582 ( .A1(n3286), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3174)
         );
  AND2_X1 U3583 ( .A1(n5100), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5087) );
  INV_X1 U3584 ( .A(n5082), .ZN(n4492) );
  OR2_X1 U3585 ( .A1(n4442), .A2(n4329), .ZN(n4349) );
  OR2_X1 U3586 ( .A1(n4121), .A2(n4120), .ZN(n5405) );
  NAND2_X1 U3587 ( .A1(n5238), .A2(n5384), .ZN(n5443) );
  AND2_X1 U3588 ( .A1(n3743), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3753)
         );
  INV_X1 U3589 ( .A(n4507), .ZN(n3726) );
  INV_X1 U3590 ( .A(n3731), .ZN(n4212) );
  NAND2_X1 U3591 ( .A1(n4564), .A2(n2970), .ZN(n3033) );
  AOI21_X1 U3592 ( .B1(n6278), .B2(n3814), .A(n3706), .ZN(n4342) );
  NOR2_X2 U3593 ( .A1(n3000), .A2(n2999), .ZN(n4301) );
  INV_X1 U3594 ( .A(n5318), .ZN(n2999) );
  AND2_X1 U3595 ( .A1(n5569), .A2(n3490), .ZN(n3491) );
  NOR2_X1 U3596 ( .A1(n5219), .A2(n3056), .ZN(n3055) );
  INV_X1 U3597 ( .A(n3486), .ZN(n3056) );
  NAND2_X1 U3598 ( .A1(n5110), .A2(n5109), .ZN(n5169) );
  NAND2_X1 U3599 ( .A1(n6013), .A2(n3041), .ZN(n3040) );
  NOR2_X1 U3600 ( .A1(n2974), .A2(n3042), .ZN(n3041) );
  INV_X1 U3601 ( .A(n3459), .ZN(n3042) );
  XNOR2_X1 U3602 ( .A(n3342), .B(n3341), .ZN(n3344) );
  INV_X1 U3603 ( .A(n3703), .ZN(n6278) );
  OR2_X1 U3604 ( .A1(n3553), .A2(n3552), .ZN(n4404) );
  AND2_X1 U3605 ( .A1(n5458), .A2(n4503), .ZN(n5967) );
  AND2_X1 U3606 ( .A1(n5458), .A2(n4504), .ZN(n5971) );
  INV_X1 U3607 ( .A(n5458), .ZN(n5970) );
  NOR2_X1 U3608 ( .A1(n3224), .A2(n3562), .ZN(n3235) );
  CLKBUF_X2 U3609 ( .A(n3285), .Z(n3436) );
  OR2_X1 U3610 ( .A1(n3420), .A2(n3419), .ZN(n3451) );
  OR2_X1 U3611 ( .A1(n3446), .A2(n3445), .ZN(n3464) );
  NAND2_X1 U3612 ( .A1(n4370), .A2(n3207), .ZN(n3508) );
  AND2_X1 U3613 ( .A1(n3537), .A2(n3536), .ZN(n3565) );
  OAI211_X1 U3614 ( .C1(n3212), .C2(n4585), .A(n4371), .B(n3232), .ZN(n3582)
         );
  NAND2_X1 U3615 ( .A1(n3207), .A2(n3231), .ZN(n3212) );
  NAND2_X1 U3616 ( .A1(n4122), .A2(n3023), .ZN(n3022) );
  INV_X1 U3617 ( .A(n4312), .ZN(n3023) );
  NOR2_X1 U3618 ( .A1(n6634), .A2(n4071), .ZN(n4072) );
  NAND2_X1 U3619 ( .A1(n5238), .A2(n2984), .ZN(n5355) );
  INV_X1 U3620 ( .A(n5105), .ZN(n3020) );
  INV_X1 U3621 ( .A(n4387), .ZN(n3713) );
  AOI21_X1 U3622 ( .B1(n3049), .B2(n3047), .A(n2983), .ZN(n3046) );
  INV_X1 U3623 ( .A(n4053), .ZN(n3047) );
  INV_X1 U3624 ( .A(n3049), .ZN(n3048) );
  NAND2_X1 U3625 ( .A1(n3616), .A2(n2996), .ZN(n2995) );
  INV_X1 U3626 ( .A(n5920), .ZN(n2996) );
  NAND2_X1 U3627 ( .A1(n2973), .A2(n6127), .ZN(n3605) );
  AOI21_X1 U3628 ( .B1(n3609), .B2(n3603), .A(n3602), .ZN(n3604) );
  AND2_X1 U3629 ( .A1(n3207), .A2(n3224), .ZN(n3504) );
  NAND2_X1 U3630 ( .A1(n4580), .A2(n6379), .ZN(n3319) );
  OR2_X1 U3631 ( .A1(n3377), .A2(n3376), .ZN(n3403) );
  INV_X1 U3632 ( .A(n3550), .ZN(n3566) );
  NAND2_X1 U3633 ( .A1(n3577), .A2(n3581), .ZN(n4412) );
  AND2_X1 U3634 ( .A1(n3359), .A2(n5257), .ZN(n4736) );
  INV_X1 U3635 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6345) );
  AND2_X1 U3636 ( .A1(n3250), .A2(n6273), .ZN(n4586) );
  AOI21_X1 U3637 ( .B1(n6390), .B2(n4562), .A(n5287), .ZN(n4584) );
  INV_X1 U3638 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6351) );
  AND2_X1 U3639 ( .A1(n3347), .A2(n4499), .ZN(n3233) );
  NAND2_X1 U3640 ( .A1(n4269), .A2(n3224), .ZN(n5085) );
  NAND2_X1 U3641 ( .A1(n5417), .A2(n2997), .ZN(n5334) );
  AND2_X1 U3642 ( .A1(n5407), .A2(n2998), .ZN(n2997) );
  INV_X1 U3643 ( .A(n4314), .ZN(n2998) );
  NAND2_X1 U3644 ( .A1(n5417), .A2(n5407), .ZN(n5409) );
  INV_X1 U3645 ( .A(n4497), .ZN(n4475) );
  OR2_X1 U3646 ( .A1(n4165), .A2(n5326), .ZN(n4222) );
  NOR2_X1 U3647 ( .A1(n4140), .A2(n5504), .ZN(n4159) );
  NAND2_X1 U3648 ( .A1(n4310), .A2(n5333), .ZN(n5314) );
  NAND2_X1 U3649 ( .A1(n4116), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4140)
         );
  INV_X1 U3650 ( .A(n5404), .ZN(n3021) );
  NAND2_X1 U3651 ( .A1(n4057), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4071)
         );
  NOR2_X1 U3652 ( .A1(n3947), .A2(n3946), .ZN(n3948) );
  CLKBUF_X1 U3653 ( .A(n5355), .Z(n5538) );
  INV_X1 U3654 ( .A(n3018), .ZN(n3016) );
  INV_X1 U3655 ( .A(n5238), .ZN(n3017) );
  NAND2_X1 U3656 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n3897), .ZN(n3947)
         );
  NOR2_X1 U3657 ( .A1(n3883), .A2(n3867), .ZN(n3896) );
  AND2_X1 U3658 ( .A1(n3834), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3835)
         );
  NOR2_X1 U3659 ( .A1(n3817), .A2(n5888), .ZN(n3834) );
  CLKBUF_X1 U3660 ( .A(n5144), .Z(n5174) );
  AND2_X1 U3661 ( .A1(n3753), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3769)
         );
  CLKBUF_X1 U3662 ( .A(n4906), .Z(n4907) );
  AOI21_X1 U3663 ( .B1(n3752), .B2(n3814), .A(n3751), .ZN(n4857) );
  NOR2_X1 U3664 ( .A1(n3742), .A2(n4852), .ZN(n3743) );
  AOI21_X1 U3665 ( .B1(n3747), .B2(n3814), .A(n3746), .ZN(n4859) );
  AND2_X1 U3666 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3718), .ZN(n3733)
         );
  AOI21_X1 U3667 ( .B1(n3717), .B2(n3814), .A(n3725), .ZN(n4507) );
  NAND2_X1 U3668 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3719) );
  AOI21_X1 U3669 ( .B1(n4734), .B2(n3814), .A(n4226), .ZN(n4434) );
  INV_X1 U3670 ( .A(n2973), .ZN(n4304) );
  NAND2_X1 U3671 ( .A1(n3045), .A2(n3046), .ZN(n5481) );
  OR2_X1 U3672 ( .A1(n5653), .A2(n3676), .ZN(n5413) );
  NOR3_X1 U3673 ( .A1(n5776), .A2(n5524), .A3(n5661), .ZN(n5525) );
  AND2_X1 U3674 ( .A1(n5357), .A2(n3664), .ZN(n5425) );
  NAND2_X1 U3675 ( .A1(n5425), .A2(n5424), .ZN(n5653) );
  NOR3_X1 U3676 ( .A1(n5446), .A2(n5445), .A3(n5376), .ZN(n5357) );
  OR2_X1 U3677 ( .A1(n5391), .A2(n5392), .ZN(n5446) );
  INV_X1 U3678 ( .A(n3053), .ZN(n3052) );
  OAI21_X1 U3679 ( .B1(n3055), .B2(n3054), .A(n3488), .ZN(n3053) );
  AND2_X1 U3680 ( .A1(n5209), .A2(n3649), .ZN(n5243) );
  NOR2_X1 U3681 ( .A1(n5175), .A2(n5176), .ZN(n5209) );
  OR2_X1 U3682 ( .A1(n5169), .A2(n5168), .ZN(n5175) );
  AND2_X1 U3683 ( .A1(n5114), .A2(n3481), .ZN(n2971) );
  NOR2_X1 U3684 ( .A1(n5899), .A2(n2977), .ZN(n5110) );
  INV_X1 U3685 ( .A(n3630), .ZN(n3001) );
  OR2_X1 U3686 ( .A1(n5581), .A2(n6050), .ZN(n5114) );
  NAND2_X1 U3687 ( .A1(n3631), .A2(n3630), .ZN(n5049) );
  AND2_X1 U3688 ( .A1(n3629), .A2(n3628), .ZN(n4910) );
  AND2_X1 U3689 ( .A1(n3624), .A2(n3623), .ZN(n5898) );
  INV_X1 U3690 ( .A(n5899), .ZN(n3631) );
  OR2_X1 U3691 ( .A1(n4509), .A2(n4508), .ZN(n5919) );
  INV_X1 U3692 ( .A(n3268), .ZN(n3012) );
  OAI211_X1 U3693 ( .C1(n3060), .C2(n3059), .A(n2976), .B(n3058), .ZN(n3266)
         );
  INV_X1 U3694 ( .A(n3323), .ZN(n3321) );
  AND2_X2 U3695 ( .A1(n3070), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5276)
         );
  NAND2_X1 U3696 ( .A1(n3218), .A2(n3554), .ZN(n4542) );
  NOR2_X1 U3697 ( .A1(n6136), .A2(n4577), .ZN(n4827) );
  OR2_X1 U3698 ( .A1(n6190), .A2(n4577), .ZN(n4953) );
  AND2_X1 U3699 ( .A1(n4683), .A2(n6284), .ZN(n4686) );
  INV_X1 U3700 ( .A(n4737), .ZN(n4628) );
  NOR2_X1 U3701 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4584), .ZN(n4737) );
  AND2_X1 U3702 ( .A1(n6374), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3570) );
  OR2_X1 U3703 ( .A1(n4324), .A2(n6384), .ZN(n4340) );
  INV_X1 U3704 ( .A(n5927), .ZN(n5939) );
  NAND2_X1 U3705 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5909), .ZN(n5897) );
  INV_X1 U3706 ( .A(n5880), .ZN(n5907) );
  AND2_X1 U3707 ( .A1(n5087), .A2(n4265), .ZN(n5943) );
  AND2_X1 U3708 ( .A1(n5938), .A2(n4274), .ZN(n5909) );
  AND2_X1 U3709 ( .A1(n5100), .A2(n4261), .ZN(n5928) );
  AND2_X1 U3710 ( .A1(n5100), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5927) );
  AND2_X1 U3711 ( .A1(n5305), .A2(n4259), .ZN(n5944) );
  INV_X1 U3712 ( .A(n5455), .ZN(n5955) );
  AND2_X1 U3713 ( .A1(n4375), .A2(n4494), .ZN(n5959) );
  INV_X1 U3714 ( .A(n5740), .ZN(n5764) );
  OR2_X1 U3715 ( .A1(n5967), .A2(n5971), .ZN(n5240) );
  NAND2_X1 U3716 ( .A1(n4498), .A2(n4497), .ZN(n5458) );
  INV_X1 U3717 ( .A(n5240), .ZN(n4944) );
  CLKBUF_X1 U3718 ( .A(n6001), .Z(n6486) );
  NOR2_X1 U3719 ( .A1(n5732), .A2(n5579), .ZN(n4048) );
  AND2_X1 U3720 ( .A1(n5435), .A2(n5434), .ZN(n5960) );
  NAND2_X1 U3721 ( .A1(n3007), .A2(n3852), .ZN(n5194) );
  INV_X1 U3722 ( .A(n3008), .ZN(n3007) );
  NOR2_X1 U3723 ( .A1(n4506), .A2(n4662), .ZN(n4570) );
  INV_X1 U3724 ( .A(n5574), .ZN(n6030) );
  NAND2_X1 U3725 ( .A1(n3026), .A2(n3025), .ZN(n4388) );
  NAND2_X1 U3726 ( .A1(n3032), .A2(n3702), .ZN(n4389) );
  NAND2_X1 U3727 ( .A1(n4342), .A2(n4212), .ZN(n3025) );
  AND2_X1 U3728 ( .A1(n5325), .A2(n5324), .ZN(n5610) );
  XNOR2_X1 U3729 ( .A(n5495), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5613)
         );
  AND2_X1 U3730 ( .A1(n3050), .A2(n2981), .ZN(n5520) );
  AND2_X1 U3731 ( .A1(n4293), .A2(n4292), .ZN(n5645) );
  NAND2_X1 U3732 ( .A1(n3487), .A2(n3055), .ZN(n3051) );
  NAND2_X1 U3733 ( .A1(n3038), .A2(n3036), .ZN(n5062) );
  NAND2_X1 U3734 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  INV_X1 U3735 ( .A(n6164), .ZN(n6135) );
  INV_X1 U3736 ( .A(n6174), .ZN(n6159) );
  INV_X1 U3737 ( .A(n6185), .ZN(n5038) );
  INV_X1 U3738 ( .A(n6272), .ZN(n6236) );
  INV_X1 U3739 ( .A(n5008), .ZN(n6275) );
  INV_X1 U3740 ( .A(n4767), .ZN(n5254) );
  OR2_X1 U3741 ( .A1(n4630), .A2(n4980), .ZN(n6496) );
  CLKBUF_X1 U3742 ( .A(n6482), .Z(n6448) );
  NOR3_X1 U3743 ( .A1(n4289), .A2(n4288), .A3(n4287), .ZN(n4290) );
  AND2_X1 U3744 ( .A1(n5303), .A2(n6452), .ZN(n4287) );
  OAI21_X1 U3745 ( .B1(n5399), .B2(n6089), .A(n3002), .ZN(U2987) );
  INV_X1 U3746 ( .A(n3003), .ZN(n3002) );
  AND2_X2 U3747 ( .A1(n3084), .A2(n4553), .ZN(n3187) );
  INV_X2 U3748 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6285) );
  AND2_X2 U3749 ( .A1(n3084), .A2(n4521), .ZN(n3198) );
  NAND2_X1 U3750 ( .A1(n3011), .A2(n3314), .ZN(n3703) );
  AND2_X2 U3751 ( .A1(n4538), .A2(n4521), .ZN(n3269) );
  NOR2_X1 U3752 ( .A1(n3017), .A2(n3016), .ZN(n5354) );
  AND2_X1 U3753 ( .A1(n3232), .A2(n3231), .ZN(n2970) );
  AOI21_X1 U3754 ( .B1(n3243), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3251), 
        .ZN(n3252) );
  AND2_X1 U3755 ( .A1(n3702), .A2(n3880), .ZN(n2972) );
  OAI21_X1 U3756 ( .B1(n3060), .B2(n3061), .A(n4554), .ZN(n4529) );
  AND2_X1 U3757 ( .A1(n3785), .A2(n2982), .ZN(n5106) );
  AND2_X1 U3758 ( .A1(n5317), .A2(n3606), .ZN(n2973) );
  AND2_X1 U3759 ( .A1(n3470), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n2974)
         );
  AND2_X2 U3760 ( .A1(n4521), .A2(n4551), .ZN(n3280) );
  AND2_X1 U3761 ( .A1(n4079), .A2(n5347), .ZN(n5348) );
  INV_X1 U3762 ( .A(n3000), .ZN(n5323) );
  OR2_X1 U3763 ( .A1(n5334), .A2(n5335), .ZN(n3000) );
  NOR2_X1 U3764 ( .A1(n4035), .A2(n4034), .ZN(n4079) );
  NAND2_X1 U3765 ( .A1(n3050), .A2(n3049), .ZN(n4217) );
  NAND2_X1 U3766 ( .A1(n5348), .A2(n5412), .ZN(n5404) );
  OR2_X1 U3767 ( .A1(n3380), .A2(n3365), .ZN(n2976) );
  OR2_X1 U3768 ( .A1(n3001), .A2(n5048), .ZN(n2977) );
  AND4_X1 U3769 ( .A1(n3092), .A2(n3091), .A3(n3090), .A4(n3089), .ZN(n3231)
         );
  AND3_X1 U3770 ( .A1(n3162), .A2(n3161), .A3(n3160), .ZN(n2978) );
  NAND2_X1 U3771 ( .A1(n3021), .A2(n4122), .ZN(n4309) );
  AND2_X1 U3772 ( .A1(n3203), .A2(n3204), .ZN(n2979) );
  BUF_X1 U3773 ( .A(n3969), .Z(n3371) );
  OR2_X1 U3774 ( .A1(n3232), .A2(n6285), .ZN(n2980) );
  OR2_X1 U3775 ( .A1(n5581), .A2(n4052), .ZN(n2981) );
  AND2_X1 U3776 ( .A1(n3248), .A2(n3313), .ZN(n3060) );
  NAND2_X1 U3777 ( .A1(n3785), .A2(n3784), .ZN(n5044) );
  INV_X1 U3778 ( .A(n3880), .ZN(n3814) );
  NAND2_X1 U3779 ( .A1(n3051), .A2(n5220), .ZN(n5580) );
  NAND2_X1 U3780 ( .A1(n3487), .A2(n3486), .ZN(n5218) );
  AND2_X1 U3781 ( .A1(n3784), .A2(n3020), .ZN(n2982) );
  AND2_X1 U3782 ( .A1(n5581), .A2(n5636), .ZN(n2983) );
  AND2_X1 U3783 ( .A1(n3018), .A2(n5356), .ZN(n2984) );
  OR2_X1 U3784 ( .A1(n5581), .A2(n5707), .ZN(n2985) );
  INV_X1 U3785 ( .A(n3004), .ZN(n5448) );
  NOR2_X1 U3786 ( .A1(n5446), .A2(n5445), .ZN(n3004) );
  NOR2_X1 U3787 ( .A1(n5537), .A2(n5536), .ZN(n2986) );
  AND2_X1 U3788 ( .A1(n2982), .A2(n5145), .ZN(n2987) );
  AND2_X1 U3789 ( .A1(n3852), .A2(n3840), .ZN(n2988) );
  INV_X1 U3790 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6379) );
  INV_X1 U3791 ( .A(n4212), .ZN(n3028) );
  AND2_X1 U3792 ( .A1(n3682), .A2(n3680), .ZN(n6121) );
  NAND2_X2 U3793 ( .A1(n3334), .A2(n3333), .ZN(n4564) );
  NOR2_X1 U3794 ( .A1(n4509), .A2(n2995), .ZN(n2989) );
  OR2_X1 U3795 ( .A1(n5581), .A2(n3485), .ZN(n2990) );
  OAI211_X1 U3796 ( .C1(n3031), .C2(n4576), .A(n3024), .B(n3027), .ZN(n4387)
         );
  NAND2_X1 U3797 ( .A1(n3060), .A2(n3061), .ZN(n4554) );
  NOR2_X1 U3798 ( .A1(n4856), .A2(n4857), .ZN(n4905) );
  INV_X1 U3799 ( .A(n4506), .ZN(n3014) );
  AND2_X1 U3800 ( .A1(n3033), .A2(STATE2_REG_2__SCAN_IN), .ZN(n2991) );
  INV_X1 U3801 ( .A(n4508), .ZN(n3616) );
  AND3_X2 U3802 ( .A1(n2979), .A2(n3205), .A3(n3206), .ZN(n4269) );
  NOR2_X2 U3803 ( .A1(n4509), .A2(n2993), .ZN(n4572) );
  AND2_X2 U3804 ( .A1(n5274), .A2(n4551), .ZN(n3286) );
  AND2_X2 U3805 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U3806 ( .A1(n3243), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U3807 ( .A1(n3005), .A2(n3213), .ZN(n3243) );
  NAND2_X1 U3808 ( .A1(n3006), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3005) );
  NAND3_X1 U3809 ( .A1(n3211), .A2(n3210), .A3(n3227), .ZN(n3006) );
  NAND2_X1 U3810 ( .A1(n3840), .A2(n5195), .ZN(n3008) );
  NAND2_X2 U3811 ( .A1(n3852), .A2(n3008), .ZN(n5200) );
  NAND3_X1 U3812 ( .A1(n3011), .A2(n6379), .A3(n3314), .ZN(n3010) );
  NAND2_X1 U3813 ( .A1(n3009), .A2(n3012), .ZN(n3011) );
  INV_X1 U3814 ( .A(n3267), .ZN(n3009) );
  NAND3_X1 U3815 ( .A1(n3014), .A2(n3015), .A3(n3013), .ZN(n4856) );
  NAND3_X1 U3816 ( .A1(n3014), .A2(n4569), .A3(n3015), .ZN(n4568) );
  NAND2_X1 U3817 ( .A1(n3785), .A2(n2987), .ZN(n5144) );
  INV_X1 U3818 ( .A(n5144), .ZN(n3833) );
  NOR2_X2 U3819 ( .A1(n5404), .A2(n3022), .ZN(n4310) );
  NAND3_X1 U3820 ( .A1(n3029), .A2(n3033), .A3(STATE2_REG_2__SCAN_IN), .ZN(
        n3026) );
  NAND2_X1 U3821 ( .A1(n3034), .A2(n4269), .ZN(n3211) );
  NAND2_X1 U3822 ( .A1(n3034), .A2(n5082), .ZN(n3589) );
  NAND2_X2 U3823 ( .A1(n3167), .A2(n3168), .ZN(n3034) );
  NAND3_X1 U3824 ( .A1(n3484), .A2(n2990), .A3(n3483), .ZN(n3035) );
  NAND2_X1 U3825 ( .A1(n3484), .A2(n3483), .ZN(n5188) );
  NAND2_X1 U3826 ( .A1(n3037), .A2(n4864), .ZN(n3036) );
  INV_X1 U3827 ( .A(n6013), .ZN(n3037) );
  AOI21_X1 U3828 ( .B1(n4864), .B2(n3042), .A(n2974), .ZN(n3038) );
  NAND3_X1 U3829 ( .A1(n3040), .A2(n5061), .A3(n3039), .ZN(n5060) );
  NAND2_X1 U3830 ( .A1(n4865), .A2(n4864), .ZN(n4863) );
  NAND2_X1 U3831 ( .A1(n6013), .A2(n3459), .ZN(n4865) );
  NAND2_X1 U3832 ( .A1(n5559), .A2(n4053), .ZN(n3050) );
  OAI21_X2 U3833 ( .B1(n3487), .B2(n3054), .A(n3052), .ZN(n5568) );
  OR2_X2 U3834 ( .A1(n5568), .A2(n3057), .ZN(n3492) );
  NAND4_X1 U3835 ( .A1(n3248), .A2(n3313), .A3(n6379), .A4(n3252), .ZN(n3058)
         );
  INV_X1 U3836 ( .A(n3252), .ZN(n3061) );
  NAND2_X1 U3837 ( .A1(n3062), .A2(n5114), .ZN(n3482) );
  OR2_X1 U3838 ( .A1(n3717), .A2(n4734), .ZN(n6136) );
  NAND2_X1 U3839 ( .A1(n4005), .A2(n2986), .ZN(n4035) );
  NOR2_X1 U3841 ( .A1(n5523), .A2(n3496), .ZN(n3497) );
  AOI22_X1 U3842 ( .A1(n3186), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3843 ( .A1(n4213), .A2(n4214), .ZN(n4230) );
  OAI211_X1 U3844 ( .C1(n5602), .C2(n6011), .A(n4215), .B(n2975), .ZN(U2956)
         );
  NAND2_X1 U3845 ( .A1(n4850), .A2(n4849), .ZN(n4848) );
  OR2_X1 U3846 ( .A1(n5366), .A2(n5369), .ZN(n3063) );
  OR2_X1 U3847 ( .A1(n3244), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3064)
         );
  OR2_X1 U3848 ( .A1(n4304), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3065)
         );
  OR2_X1 U3849 ( .A1(n4304), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3066)
         );
  AND4_X1 U3850 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3068)
         );
  INV_X1 U3851 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3481) );
  OR2_X1 U3852 ( .A1(n5776), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3069)
         );
  NAND2_X1 U3853 ( .A1(n4572), .A2(n5898), .ZN(n5899) );
  NOR2_X1 U3854 ( .A1(n3209), .A2(n3582), .ZN(n3210) );
  NAND2_X1 U3855 ( .A1(n3212), .A2(n3505), .ZN(n3213) );
  AND3_X1 U3856 ( .A1(n3311), .A2(n3310), .A3(n3309), .ZN(n3341) );
  OR2_X1 U3857 ( .A1(n3400), .A2(n3399), .ZN(n3452) );
  NAND2_X1 U3858 ( .A1(n4326), .A2(n3236), .ZN(n3237) );
  NAND2_X1 U3859 ( .A1(n3212), .A2(n4603), .ZN(n3219) );
  AOI22_X1 U3860 ( .A1(n3195), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3201) );
  INV_X1 U3861 ( .A(n5046), .ZN(n3784) );
  INV_X1 U3862 ( .A(n3388), .ZN(n3389) );
  AND2_X1 U3863 ( .A1(n3317), .A2(n3466), .ZN(n3471) );
  INV_X1 U3864 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3603) );
  AND2_X1 U3865 ( .A1(n3543), .A2(n3542), .ZN(n3550) );
  AND2_X1 U3866 ( .A1(n3208), .A2(n4412), .ZN(n3227) );
  NAND2_X1 U3867 ( .A1(n3320), .A2(n3343), .ZN(n3323) );
  AND4_X1 U3868 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), .ZN(n3089)
         );
  AOI22_X1 U3869 ( .A1(n3195), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3127) );
  AND2_X1 U3870 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4072), .ZN(n4116)
         );
  INV_X1 U3871 ( .A(n4859), .ZN(n3748) );
  INV_X1 U3872 ( .A(n3449), .ZN(n3447) );
  INV_X1 U3873 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3070) );
  NAND2_X1 U3874 ( .A1(n3365), .A2(n3364), .ZN(n3544) );
  NAND2_X1 U3875 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  NAND2_X1 U3876 ( .A1(n4422), .A2(n5373), .ZN(n4300) );
  INV_X1 U3877 ( .A(n3979), .ZN(n3980) );
  OR2_X1 U3878 ( .A1(n3866), .A2(n5204), .ZN(n3883) );
  NOR2_X1 U3879 ( .A1(n3787), .A2(n3786), .ZN(n3802) );
  NOR2_X1 U3880 ( .A1(n4909), .A2(n4910), .ZN(n3630) );
  AND2_X1 U3881 ( .A1(n3615), .A2(n3614), .ZN(n4508) );
  AOI21_X1 U3882 ( .B1(n5309), .B2(REIP_REG_31__SCAN_IN), .A(n5308), .ZN(n5310) );
  AND2_X1 U3883 ( .A1(n3998), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4057)
         );
  NAND2_X1 U3884 ( .A1(n3769), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3787)
         );
  INV_X1 U3885 ( .A(n5931), .ZN(n5938) );
  INV_X1 U3886 ( .A(n5943), .ZN(n5924) );
  AND2_X1 U3887 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3980), .ZN(n3998)
         );
  NOR2_X1 U3888 ( .A1(n3914), .A2(n5854), .ZN(n3897) );
  NAND2_X1 U3889 ( .A1(n3356), .A2(n3355), .ZN(n3357) );
  NAND2_X1 U3890 ( .A1(n5494), .A2(n4218), .ZN(n4219) );
  NAND2_X1 U3891 ( .A1(n5581), .A2(n6050), .ZN(n5113) );
  AOI21_X1 U3892 ( .B1(n4386), .B2(n4385), .A(n3353), .ZN(n6032) );
  OR3_X1 U3893 ( .A1(n4442), .A2(n3573), .A3(n3155), .ZN(n3574) );
  OR2_X1 U3894 ( .A1(n4630), .A2(n4577), .ZN(n4797) );
  OAI21_X1 U3895 ( .B1(n5399), .B2(n5910), .A(n5310), .ZN(n5311) );
  NOR2_X1 U3896 ( .A1(n6431), .A2(n5857), .ZN(n5371) );
  NOR2_X1 U3897 ( .A1(n4275), .A2(n5897), .ZN(n5886) );
  OR4_X1 U3898 ( .A1(n6483), .A2(n6101), .A3(n6375), .A4(n6386), .ZN(n5100) );
  NAND2_X1 U3899 ( .A1(n5087), .A2(n4272), .ZN(n5931) );
  INV_X1 U3900 ( .A(n4440), .ZN(n4481) );
  NAND2_X1 U3901 ( .A1(n3835), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3866)
         );
  NAND2_X1 U3902 ( .A1(n3733), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3742)
         );
  NAND2_X1 U3903 ( .A1(n4404), .A2(n4494), .ZN(n4442) );
  OR2_X1 U3904 ( .A1(n5225), .A2(n4381), .ZN(n5674) );
  AND2_X1 U3905 ( .A1(n6043), .A2(n3685), .ZN(n5708) );
  INV_X1 U3906 ( .A(n5805), .ZN(n6129) );
  NAND2_X1 U3907 ( .A1(n3575), .A2(n3574), .ZN(n3682) );
  AND2_X1 U3908 ( .A1(n4404), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5287) );
  INV_X1 U3909 ( .A(n5028), .ZN(n4981) );
  INV_X1 U3910 ( .A(n4564), .ZN(n4914) );
  OAI21_X1 U3911 ( .B1(n6169), .B2(n6464), .A(n4921), .ZN(n6171) );
  NOR2_X1 U3912 ( .A1(n4953), .A2(n4564), .ZN(n6185) );
  INV_X1 U3913 ( .A(n6227), .ZN(n6209) );
  OR2_X1 U3914 ( .A1(n6277), .A2(n4577), .ZN(n4689) );
  INV_X1 U3915 ( .A(n6339), .ZN(n6318) );
  NOR2_X1 U3916 ( .A1(n4797), .A2(n4914), .ZN(n5267) );
  NOR2_X1 U3917 ( .A1(n6463), .A2(n4584), .ZN(n4616) );
  INV_X1 U3918 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U3919 ( .A1(n4349), .A2(n4340), .ZN(n6483) );
  INV_X1 U3920 ( .A(n5311), .ZN(n5312) );
  INV_X1 U3921 ( .A(n5944), .ZN(n5910) );
  NAND2_X1 U3922 ( .A1(n5100), .A2(n4235), .ZN(n5880) );
  NOR2_X1 U3923 ( .A1(n5974), .A2(n6486), .ZN(n5993) );
  INV_X1 U3924 ( .A(n5974), .ZN(n6004) );
  NOR2_X1 U3925 ( .A1(n4048), .A2(n4047), .ZN(n4049) );
  OR2_X1 U3926 ( .A1(n4442), .A2(n6360), .ZN(n6011) );
  AND2_X1 U3927 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  INV_X1 U3928 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4955) );
  OR2_X1 U3929 ( .A1(n6136), .A2(n4980), .ZN(n6164) );
  OR2_X1 U3930 ( .A1(n6136), .A2(n6189), .ZN(n6174) );
  OR2_X1 U3931 ( .A1(n6190), .A2(n4980), .ZN(n6227) );
  OR2_X1 U3932 ( .A1(n6190), .A2(n6189), .ZN(n6272) );
  OR2_X1 U3933 ( .A1(n4689), .A2(n4564), .ZN(n4876) );
  OR2_X1 U3934 ( .A1(n6277), .A2(n4980), .ZN(n6323) );
  OR2_X1 U3935 ( .A1(n6277), .A2(n6189), .ZN(n6339) );
  OAI21_X1 U3936 ( .B1(n4233), .B2(n5880), .A(n4290), .ZN(U2797) );
  OAI211_X1 U3937 ( .C1(n4308), .C2(n6011), .A(n4232), .B(n4231), .ZN(U2955)
         );
  NOR2_X4 U3938 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U3939 ( .A1(n2966), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3074) );
  NAND2_X1 U3940 ( .A1(n3285), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3073) );
  NAND2_X1 U3941 ( .A1(n2965), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3072)
         );
  NAND2_X1 U3942 ( .A1(n3269), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3071) );
  NAND2_X1 U3943 ( .A1(n3196), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3079) );
  NAND2_X1 U3944 ( .A1(n3257), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3078)
         );
  NAND2_X1 U3945 ( .A1(n3286), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3077)
         );
  AND2_X4 U3946 ( .A1(n5274), .A2(n3084), .ZN(n3969) );
  NAND2_X1 U3947 ( .A1(n3969), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3076) );
  NAND2_X1 U3948 ( .A1(n3186), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3083)
         );
  NAND2_X1 U3949 ( .A1(n3194), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3082) );
  NAND2_X1 U3950 ( .A1(n3198), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3081) );
  NAND2_X1 U3951 ( .A1(n3280), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3080)
         );
  NAND2_X1 U3952 ( .A1(n3189), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3953 ( .A1(n3187), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3087) );
  AND2_X2 U3954 ( .A1(n4553), .A2(n4551), .ZN(n3188) );
  NAND2_X1 U3955 ( .A1(n3188), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3086)
         );
  AND2_X2 U3956 ( .A1(n5276), .A2(n3084), .ZN(n3197) );
  NAND2_X1 U3957 ( .A1(n3197), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3085) );
  AOI22_X1 U3958 ( .A1(n2965), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3096) );
  AOI22_X1 U3959 ( .A1(n3285), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3095) );
  AOI22_X1 U3960 ( .A1(n3194), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3094) );
  AOI22_X1 U3961 ( .A1(n3197), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3093) );
  AOI22_X1 U3962 ( .A1(n2966), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3969), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3100) );
  AOI22_X1 U3963 ( .A1(n3189), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3099) );
  AOI22_X1 U3964 ( .A1(n3286), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3098) );
  NAND2_X2 U3965 ( .A1(n4612), .A2(n4499), .ZN(n4371) );
  NAND2_X1 U3966 ( .A1(n3186), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3106)
         );
  NAND2_X1 U3967 ( .A1(n3194), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U3968 ( .A1(n3198), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U3969 ( .A1(n3280), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3103)
         );
  NAND2_X1 U3970 ( .A1(n3189), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U3971 ( .A1(n3197), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3109) );
  NAND2_X1 U3972 ( .A1(n3188), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3108)
         );
  NAND2_X1 U3973 ( .A1(n3187), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3974 ( .A1(n3195), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3114) );
  NAND2_X1 U3975 ( .A1(n3285), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U3976 ( .A1(n4081), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3112)
         );
  NAND2_X1 U3977 ( .A1(n3269), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3111) );
  NAND2_X1 U3978 ( .A1(n3196), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3118) );
  NAND2_X1 U3979 ( .A1(n3257), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3117)
         );
  NAND2_X1 U3980 ( .A1(n3286), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3116)
         );
  NAND2_X1 U3981 ( .A1(n3969), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3115) );
  NAND2_X1 U3982 ( .A1(n4371), .A2(n4368), .ZN(n3133) );
  AOI22_X1 U3983 ( .A1(n3186), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U3984 ( .A1(n3269), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U3985 ( .A1(n3189), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3286), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3124) );
  AOI22_X1 U3986 ( .A1(n3194), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3123) );
  NAND4_X1 U3987 ( .A1(n3126), .A2(n3125), .A3(n3124), .A4(n3123), .ZN(n3132)
         );
  AOI22_X1 U3988 ( .A1(n4081), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U3989 ( .A1(n3969), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U3990 ( .A1(n3197), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3128) );
  NAND4_X1 U3991 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .ZN(n3131)
         );
  OR2_X2 U3992 ( .A1(n3132), .A2(n3131), .ZN(n3232) );
  NAND2_X1 U3993 ( .A1(n3133), .A2(n3232), .ZN(n3154) );
  NAND2_X1 U3994 ( .A1(n3187), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U3995 ( .A1(n3197), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U3996 ( .A1(n3188), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3135)
         );
  NAND2_X1 U3997 ( .A1(n3189), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U3998 ( .A1(n3195), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U3999 ( .A1(n3285), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3140) );
  NAND2_X1 U4000 ( .A1(n4081), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3139)
         );
  NAND2_X1 U4001 ( .A1(n3269), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U4002 ( .A1(n3186), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3145)
         );
  NAND2_X1 U4003 ( .A1(n3194), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U4004 ( .A1(n3198), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U4005 ( .A1(n3280), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3142)
         );
  NAND2_X1 U4006 ( .A1(n3196), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4007 ( .A1(n3257), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3148)
         );
  NAND2_X1 U4008 ( .A1(n3286), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3147)
         );
  NAND2_X1 U4009 ( .A1(n3969), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U4010 ( .A1(n2970), .A2(n3155), .ZN(n3166) );
  AOI22_X1 U4011 ( .A1(n3197), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4012 ( .A1(n4081), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3286), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4013 ( .A1(n3186), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4014 ( .A1(n3187), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4015 ( .A1(n3196), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3969), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4016 ( .A1(n3269), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4017 ( .A1(n3194), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4018 ( .A1(n3285), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U4019 ( .A1(n2966), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3172) );
  NAND2_X1 U4020 ( .A1(n3285), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4021 ( .A1(n4081), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3170)
         );
  NAND2_X1 U4022 ( .A1(n3269), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U4023 ( .A1(n3196), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4024 ( .A1(n3257), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3175)
         );
  NAND2_X1 U4025 ( .A1(n3969), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3173) );
  NAND2_X1 U4026 ( .A1(n3186), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3180)
         );
  NAND2_X1 U4027 ( .A1(n3194), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U4028 ( .A1(n3198), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3178) );
  NAND2_X1 U4029 ( .A1(n3280), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3177)
         );
  NAND2_X1 U4030 ( .A1(n3197), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U4031 ( .A1(n3189), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U4032 ( .A1(n3188), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3182)
         );
  NAND2_X1 U4033 ( .A1(n3187), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3181) );
  AND2_X1 U4034 ( .A1(n4370), .A2(n3232), .ZN(n3185) );
  NAND2_X1 U4035 ( .A1(n4371), .A2(n3185), .ZN(n3558) );
  AOI22_X1 U4036 ( .A1(n4081), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3969), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4037 ( .A1(n3186), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U4038 ( .A1(n3286), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4039 ( .A1(n3189), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3190) );
  AOI22_X1 U4040 ( .A1(n3285), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U4041 ( .A1(n3197), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4042 ( .A1(n3198), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4043 ( .A1(n3558), .A2(n4351), .ZN(n3208) );
  INV_X1 U4044 ( .A(n3508), .ZN(n3577) );
  INV_X1 U4045 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6399) );
  XNOR2_X1 U4046 ( .A(n6399), .B(STATE_REG_2__SCAN_IN), .ZN(n3562) );
  OAI211_X1 U4047 ( .C1(n3235), .C2(n3207), .A(n3347), .B(n5085), .ZN(n3209)
         );
  NOR2_X1 U4048 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5818) );
  NAND2_X1 U4049 ( .A1(n5818), .A2(n6379), .ZN(n4038) );
  MUX2_X1 U4050 ( .A(n3570), .B(n4038), .S(n4955), .Z(n3214) );
  NAND2_X1 U4051 ( .A1(n5085), .A2(n4368), .ZN(n3216) );
  NAND2_X1 U4052 ( .A1(n3229), .A2(n3216), .ZN(n3584) );
  INV_X1 U4053 ( .A(n4603), .ZN(n4369) );
  AND3_X1 U4054 ( .A1(n4368), .A2(n4369), .A3(n4269), .ZN(n3218) );
  NAND2_X1 U4055 ( .A1(n5818), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6385) );
  INV_X1 U4056 ( .A(n6385), .ZN(n3221) );
  NAND2_X1 U4057 ( .A1(n3219), .A2(n4351), .ZN(n3220) );
  NAND2_X1 U4058 ( .A1(n3212), .A2(n4585), .ZN(n3223) );
  NAND2_X1 U4059 ( .A1(n3223), .A2(n4603), .ZN(n3225) );
  OAI21_X1 U4060 ( .B1(n3582), .B2(n3225), .A(n3224), .ZN(n3226) );
  NAND4_X1 U4061 ( .A1(n3228), .A2(n3227), .A3(n3589), .A4(n3226), .ZN(n3268)
         );
  NAND2_X1 U4062 ( .A1(n3555), .A2(n3222), .ZN(n4557) );
  NOR2_X1 U4063 ( .A1(n3207), .A2(n4603), .ZN(n3230) );
  NAND3_X1 U4064 ( .A1(n3230), .A2(n4368), .A3(n5082), .ZN(n4413) );
  INV_X1 U4065 ( .A(n3232), .ZN(n5459) );
  NAND2_X1 U4066 ( .A1(n4612), .A2(n3232), .ZN(n4500) );
  INV_X1 U4067 ( .A(n3678), .ZN(n3238) );
  INV_X1 U4068 ( .A(n3558), .ZN(n3234) );
  INV_X1 U4069 ( .A(n3207), .ZN(n4499) );
  INV_X1 U4070 ( .A(n3235), .ZN(n3236) );
  NAND3_X1 U4071 ( .A1(n4557), .A2(n3238), .A3(n3237), .ZN(n3242) );
  INV_X1 U4072 ( .A(n4038), .ZN(n3361) );
  XNOR2_X1 U4073 ( .A(n4955), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4989)
         );
  NAND2_X1 U4074 ( .A1(n3361), .A2(n4989), .ZN(n3240) );
  INV_X1 U4075 ( .A(n3570), .ZN(n3360) );
  NAND2_X1 U4076 ( .A1(n3360), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4077 ( .A1(n3240), .A2(n3239), .ZN(n3244) );
  AND2_X1 U4078 ( .A1(n3064), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4079 ( .A1(n3242), .A2(n3241), .ZN(n3312) );
  NAND2_X1 U4080 ( .A1(n3314), .A2(n3312), .ZN(n3248) );
  NAND2_X1 U4081 ( .A1(n3242), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U4082 ( .A1(n3243), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3246) );
  INV_X1 U4083 ( .A(n3244), .ZN(n3245) );
  NAND2_X1 U4084 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U4085 ( .A1(n3249), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3250) );
  NOR2_X1 U4086 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6345), .ZN(n4979)
         );
  NAND2_X1 U4087 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4979), .ZN(n6273) );
  OAI22_X1 U4088 ( .A1(n4038), .A2(n4586), .B1(n3570), .B2(n6351), .ZN(n3251)
         );
  AOI22_X1 U4089 ( .A1(n4168), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4090 ( .A1(n3436), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4091 ( .A1(n4081), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4092 ( .A1(n4194), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3253) );
  NAND4_X1 U4093 ( .A1(n3256), .A2(n3255), .A3(n3254), .A4(n3253), .ZN(n3263)
         );
  AOI22_X1 U4094 ( .A1(n4187), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4095 ( .A1(n4196), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3260) );
  INV_X1 U4096 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6524) );
  AOI22_X1 U4097 ( .A1(n2964), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4098 ( .A1(n3187), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3258) );
  NAND4_X1 U4099 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(n3262)
         );
  INV_X1 U4100 ( .A(n3264), .ZN(n3380) );
  NAND2_X1 U4101 ( .A1(n4269), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3364) );
  INV_X1 U4102 ( .A(n3364), .ZN(n3308) );
  AOI22_X1 U4103 ( .A1(n3308), .A2(n3264), .B1(n3505), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4104 ( .A1(n4168), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4105 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n3197), .B1(n3189), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4106 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3194), .B1(n3198), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4107 ( .A1(n4541), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3270) );
  NAND4_X1 U4108 ( .A1(n3273), .A2(n3272), .A3(n3271), .A4(n3270), .ZN(n3279)
         );
  AOI22_X1 U4109 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n4081), .B1(n3257), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4110 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4187), .B1(n3371), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4111 ( .A1(n3436), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4112 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n2964), .B1(n4169), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3274) );
  NAND4_X1 U4113 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3278)
         );
  INV_X1 U4114 ( .A(n3346), .ZN(n3293) );
  AOI22_X1 U4115 ( .A1(n4168), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4116 ( .A1(n4081), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3257), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4117 ( .A1(n3197), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4118 ( .A1(n3435), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3281) );
  NAND4_X1 U4119 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3292)
         );
  AOI22_X1 U4120 ( .A1(n4541), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4121 ( .A1(n3436), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4122 ( .A1(n2964), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4123 ( .A1(n3189), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3287) );
  NAND4_X1 U4124 ( .A1(n3290), .A2(n3289), .A3(n3288), .A4(n3287), .ZN(n3291)
         );
  XNOR2_X1 U4125 ( .A(n3293), .B(n3466), .ZN(n3294) );
  INV_X1 U4126 ( .A(n3365), .ZN(n3317) );
  NAND2_X1 U4127 ( .A1(n3294), .A2(n3317), .ZN(n3331) );
  INV_X1 U4128 ( .A(n3505), .ZN(n3539) );
  INV_X1 U4129 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3297) );
  AOI21_X1 U4130 ( .B1(n4370), .B2(n3466), .A(n6379), .ZN(n3296) );
  NAND2_X1 U4131 ( .A1(n4269), .A2(n3346), .ZN(n3295) );
  OAI211_X1 U4132 ( .C1(n3539), .C2(n3297), .A(n3296), .B(n3295), .ZN(n3329)
         );
  INV_X1 U4133 ( .A(n3466), .ZN(n3476) );
  NAND2_X1 U4134 ( .A1(n3317), .A2(n3476), .ZN(n3311) );
  NAND2_X1 U4135 ( .A1(n3505), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4136 ( .A1(n4081), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4137 ( .A1(n4196), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4138 ( .A1(n4168), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4139 ( .A1(n4186), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3298) );
  NAND4_X1 U4140 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3307)
         );
  AOI22_X1 U4141 ( .A1(n3436), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4142 ( .A1(n4187), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4143 ( .A1(n2964), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3187), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4144 ( .A1(n3435), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3302) );
  NAND4_X1 U4145 ( .A1(n3305), .A2(n3304), .A3(n3303), .A4(n3302), .ZN(n3306)
         );
  NAND2_X1 U4146 ( .A1(n3308), .A2(n3345), .ZN(n3309) );
  NAND2_X1 U4147 ( .A1(n3342), .A2(n3341), .ZN(n3320) );
  NAND2_X1 U4148 ( .A1(n3313), .A2(n3312), .ZN(n3316) );
  INV_X1 U4149 ( .A(n3314), .ZN(n3315) );
  XNOR2_X2 U4150 ( .A(n3316), .B(n3315), .ZN(n4580) );
  NAND2_X1 U4151 ( .A1(n3317), .A2(n3345), .ZN(n3318) );
  INV_X1 U4152 ( .A(n3322), .ZN(n3324) );
  NAND2_X1 U4153 ( .A1(n3324), .A2(n3323), .ZN(n3325) );
  INV_X1 U4154 ( .A(n3504), .ZN(n3472) );
  NAND2_X1 U4155 ( .A1(n3345), .A2(n3346), .ZN(n3381) );
  XNOR2_X1 U4156 ( .A(n3381), .B(n3380), .ZN(n3327) );
  NAND2_X1 U4157 ( .A1(n4269), .A2(n4603), .ZN(n3335) );
  INV_X1 U4158 ( .A(n3335), .ZN(n3326) );
  AOI21_X1 U4159 ( .B1(n3327), .B2(n4351), .A(n3326), .ZN(n3328) );
  NAND2_X1 U4160 ( .A1(n6031), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3354)
         );
  INV_X1 U4161 ( .A(n3329), .ZN(n3332) );
  NAND2_X1 U4162 ( .A1(n3330), .A2(n3329), .ZN(n3334) );
  INV_X1 U4163 ( .A(n4351), .ZN(n6488) );
  OAI21_X1 U4164 ( .B1(n6488), .B2(n3346), .A(n3335), .ZN(n3336) );
  INV_X1 U4165 ( .A(n3336), .ZN(n3337) );
  NAND2_X1 U4166 ( .A1(n4346), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3338)
         );
  INV_X1 U4167 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U4168 ( .A1(n3338), .A2(n6127), .ZN(n3340) );
  AND2_X1 U4169 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4170 ( .A1(n4346), .A2(n3339), .ZN(n3352) );
  AND2_X1 U4171 ( .A1(n3340), .A2(n3352), .ZN(n4386) );
  NAND2_X1 U4172 ( .A1(n4576), .A2(n3504), .ZN(n3351) );
  OAI21_X1 U4173 ( .B1(n3346), .B2(n3345), .A(n3381), .ZN(n3348) );
  OAI211_X1 U4174 ( .C1(n3348), .C2(n6488), .A(n3347), .B(n3207), .ZN(n3349)
         );
  INV_X1 U4175 ( .A(n3349), .ZN(n3350) );
  NAND2_X1 U4176 ( .A1(n3351), .A2(n3350), .ZN(n4385) );
  INV_X1 U4177 ( .A(n3352), .ZN(n3353) );
  NAND2_X1 U4178 ( .A1(n3354), .A2(n6032), .ZN(n3358) );
  INV_X1 U4179 ( .A(n6031), .ZN(n3356) );
  INV_X1 U4180 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3355) );
  AND2_X1 U4181 ( .A1(n3358), .A2(n3357), .ZN(n4514) );
  NAND2_X1 U4182 ( .A1(n3243), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3363) );
  INV_X1 U4183 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6358) );
  NOR3_X1 U4184 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6351), .A3(n6345), 
        .ZN(n6199) );
  NAND2_X1 U4185 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6199), .ZN(n6195) );
  NAND2_X1 U4186 ( .A1(n6358), .A2(n6195), .ZN(n3359) );
  NAND3_X1 U4187 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4709) );
  INV_X1 U4188 ( .A(n4709), .ZN(n4633) );
  NAND2_X1 U4189 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4633), .ZN(n5257) );
  AOI22_X1 U4190 ( .A1(n3361), .A2(n4736), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3360), .ZN(n3362) );
  AOI22_X1 U4191 ( .A1(n4168), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4192 ( .A1(n3436), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4193 ( .A1(n2965), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4194 ( .A1(n4194), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3367) );
  NAND4_X1 U4195 ( .A1(n3370), .A2(n3369), .A3(n3368), .A4(n3367), .ZN(n3377)
         );
  AOI22_X1 U4196 ( .A1(n4187), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4197 ( .A1(n4196), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4198 ( .A1(n2964), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4199 ( .A1(n4195), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3372) );
  NAND4_X1 U4200 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3376)
         );
  AOI22_X1 U4201 ( .A1(n3544), .A2(n3403), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3505), .ZN(n3378) );
  NAND2_X1 U4202 ( .A1(n3717), .A2(n3504), .ZN(n3385) );
  NAND2_X1 U4203 ( .A1(n3381), .A2(n3380), .ZN(n3404) );
  INV_X1 U4204 ( .A(n3403), .ZN(n3382) );
  XNOR2_X1 U4205 ( .A(n3404), .B(n3382), .ZN(n3383) );
  NAND2_X1 U4206 ( .A1(n3383), .A2(n4351), .ZN(n3384) );
  INV_X1 U4207 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6099) );
  XNOR2_X1 U4208 ( .A(n3386), .B(n6099), .ZN(n4512) );
  NAND2_X1 U4209 ( .A1(n4514), .A2(n4512), .ZN(n4513) );
  NAND2_X1 U4210 ( .A1(n3386), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3387)
         );
  NAND2_X1 U4211 ( .A1(n4513), .A2(n3387), .ZN(n6021) );
  AOI22_X1 U4212 ( .A1(n4168), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4213 ( .A1(n3436), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4214 ( .A1(n2965), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4215 ( .A1(n4194), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4216 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3400)
         );
  AOI22_X1 U4217 ( .A1(n4187), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4218 ( .A1(n4196), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4219 ( .A1(n2964), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4220 ( .A1(n4195), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3395) );
  NAND4_X1 U4221 ( .A1(n3398), .A2(n3397), .A3(n3396), .A4(n3395), .ZN(n3399)
         );
  NAND2_X1 U4222 ( .A1(n3544), .A2(n3452), .ZN(n3402) );
  NAND2_X1 U4223 ( .A1(n3505), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3401) );
  NAND2_X1 U4224 ( .A1(n3402), .A2(n3401), .ZN(n3432) );
  NAND2_X1 U4225 ( .A1(n3737), .A2(n3504), .ZN(n3407) );
  NAND2_X1 U4226 ( .A1(n3404), .A2(n3403), .ZN(n3454) );
  XNOR2_X1 U4227 ( .A(n3454), .B(n3452), .ZN(n3405) );
  NAND2_X1 U4228 ( .A1(n3405), .A2(n4351), .ZN(n3406) );
  NAND2_X1 U4229 ( .A1(n3407), .A2(n3406), .ZN(n3408) );
  INV_X1 U4230 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6100) );
  XNOR2_X1 U4231 ( .A(n3408), .B(n6100), .ZN(n6022) );
  NAND2_X1 U4232 ( .A1(n6021), .A2(n6022), .ZN(n6023) );
  NAND2_X1 U4233 ( .A1(n3408), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3409)
         );
  NAND2_X1 U4234 ( .A1(n6023), .A2(n3409), .ZN(n4850) );
  INV_X1 U4235 ( .A(n3432), .ZN(n3410) );
  AOI22_X1 U4236 ( .A1(n4168), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3414) );
  INV_X1 U4237 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U4238 ( .A1(n3436), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4239 ( .A1(n4081), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4240 ( .A1(n4194), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3411) );
  NAND4_X1 U4241 ( .A1(n3414), .A2(n3413), .A3(n3412), .A4(n3411), .ZN(n3420)
         );
  AOI22_X1 U4242 ( .A1(n4187), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4243 ( .A1(n4196), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4244 ( .A1(n2964), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4245 ( .A1(n4195), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3415) );
  NAND4_X1 U4246 ( .A1(n3418), .A2(n3417), .A3(n3416), .A4(n3415), .ZN(n3419)
         );
  AOI22_X1 U4247 ( .A1(n3544), .A2(n3451), .B1(INSTQUEUE_REG_0__5__SCAN_IN), 
        .B2(n3505), .ZN(n3430) );
  XNOR2_X1 U4248 ( .A(n3421), .B(n3430), .ZN(n3738) );
  NAND2_X1 U4249 ( .A1(n3738), .A2(n3504), .ZN(n3426) );
  INV_X1 U4250 ( .A(n3452), .ZN(n3422) );
  OR2_X1 U4251 ( .A1(n3454), .A2(n3422), .ZN(n3423) );
  XNOR2_X1 U4252 ( .A(n3423), .B(n3451), .ZN(n3424) );
  NAND2_X1 U4253 ( .A1(n3424), .A2(n4351), .ZN(n3425) );
  NAND2_X1 U4254 ( .A1(n3426), .A2(n3425), .ZN(n3427) );
  INV_X1 U4255 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5121) );
  XNOR2_X1 U4256 ( .A(n3427), .B(n5121), .ZN(n4849) );
  NAND2_X1 U4257 ( .A1(n3427), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3428)
         );
  INV_X1 U4258 ( .A(n3429), .ZN(n3434) );
  INV_X1 U4259 ( .A(n3430), .ZN(n3431) );
  AOI22_X1 U4260 ( .A1(n4168), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4261 ( .A1(n3436), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4262 ( .A1(n3366), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4263 ( .A1(n4194), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3437) );
  NAND4_X1 U4264 ( .A1(n3440), .A2(n3439), .A3(n3438), .A4(n3437), .ZN(n3446)
         );
  AOI22_X1 U4265 ( .A1(n4187), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4266 ( .A1(n4196), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4267 ( .A1(n2964), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4268 ( .A1(n4195), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3441) );
  NAND4_X1 U4269 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3445)
         );
  AOI22_X1 U4270 ( .A1(n3544), .A2(n3464), .B1(n3505), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3449) );
  NAND2_X1 U4271 ( .A1(n3450), .A2(n3449), .ZN(n3747) );
  NAND3_X1 U4272 ( .A1(n3475), .A2(n3747), .A3(n3504), .ZN(n3457) );
  NAND2_X1 U4273 ( .A1(n3452), .A2(n3451), .ZN(n3453) );
  OR2_X1 U4274 ( .A1(n3454), .A2(n3453), .ZN(n3463) );
  XNOR2_X1 U4275 ( .A(n3463), .B(n3464), .ZN(n3455) );
  NAND2_X1 U4276 ( .A1(n3455), .A2(n4351), .ZN(n3456) );
  NAND2_X1 U4277 ( .A1(n3457), .A2(n3456), .ZN(n3458) );
  INV_X1 U4278 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5122) );
  XNOR2_X1 U4279 ( .A(n3458), .B(n5122), .ZN(n6014) );
  NAND2_X1 U4280 ( .A1(n3458), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3459)
         );
  INV_X1 U4281 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3461) );
  NAND2_X1 U4282 ( .A1(n3544), .A2(n3466), .ZN(n3460) );
  OAI21_X1 U4283 ( .B1(n3461), .B2(n3539), .A(n3460), .ZN(n3462) );
  NAND2_X1 U4284 ( .A1(n3752), .A2(n3504), .ZN(n3469) );
  INV_X1 U4285 ( .A(n3463), .ZN(n3465) );
  NAND2_X1 U4286 ( .A1(n3465), .A2(n3464), .ZN(n3477) );
  XNOR2_X1 U4287 ( .A(n3477), .B(n3466), .ZN(n3467) );
  NAND2_X1 U4288 ( .A1(n3467), .A2(n4351), .ZN(n3468) );
  NAND2_X1 U4289 ( .A1(n3469), .A2(n3468), .ZN(n3470) );
  INV_X1 U4290 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6074) );
  XNOR2_X1 U4291 ( .A(n3470), .B(n6074), .ZN(n4864) );
  INV_X1 U4292 ( .A(n3471), .ZN(n3473) );
  NOR2_X1 U4293 ( .A1(n3473), .A2(n3472), .ZN(n3474) );
  OR3_X1 U4294 ( .A1(n3477), .A2(n3476), .A3(n6488), .ZN(n3478) );
  NAND2_X1 U4295 ( .A1(n5581), .A2(n3478), .ZN(n3479) );
  INV_X1 U4296 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6066) );
  XNOR2_X1 U4297 ( .A(n3479), .B(n6066), .ZN(n5061) );
  NAND2_X1 U4298 ( .A1(n3479), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3480)
         );
  NAND2_X1 U4299 ( .A1(n5060), .A2(n3480), .ZN(n5115) );
  INV_X1 U4300 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6050) );
  OAI21_X2 U4301 ( .B1(n5179), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5776), 
        .ZN(n3484) );
  NAND3_X1 U4302 ( .A1(n3482), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3483) );
  INV_X1 U4303 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3485) );
  NAND2_X1 U4304 ( .A1(n5581), .A2(n3485), .ZN(n5186) );
  XNOR2_X1 U4305 ( .A(n5581), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5787)
         );
  INV_X1 U4306 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U4307 ( .A1(n5581), .A2(n3645), .ZN(n3486) );
  INV_X1 U4308 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6548) );
  AND2_X1 U4309 ( .A1(n5581), .A2(n6548), .ZN(n5219) );
  OR2_X1 U4310 ( .A1(n5581), .A2(n6548), .ZN(n5220) );
  INV_X1 U4311 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U4312 ( .A1(n5581), .A2(n5707), .ZN(n3488) );
  NAND2_X1 U4313 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3690) );
  AND2_X1 U4314 ( .A1(n5581), .A2(n3690), .ZN(n3489) );
  INV_X1 U4315 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5775) );
  AND2_X1 U4316 ( .A1(n5581), .A2(n5775), .ZN(n5570) );
  OR2_X1 U4317 ( .A1(n5581), .A2(n5775), .ZN(n5569) );
  OAI21_X1 U4318 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5776), .ZN(n3490) );
  INV_X1 U4319 ( .A(n3492), .ZN(n3493) );
  AOI21_X1 U4320 ( .B1(n3493), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5776), 
        .ZN(n3494) );
  XNOR2_X1 U4321 ( .A(n5581), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5553)
         );
  XNOR2_X1 U4322 ( .A(n5581), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5548)
         );
  INV_X1 U4323 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U4324 ( .A1(n5776), .A2(n5661), .ZN(n5540) );
  AND2_X1 U4325 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5655) );
  AND4_X1 U4326 ( .A1(n3495), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5655), 
        .A4(n5581), .ZN(n3496) );
  XNOR2_X1 U4327 ( .A(n3497), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3699)
         );
  NAND2_X1 U4328 ( .A1(n3222), .A2(n3207), .ZN(n3498) );
  NAND2_X1 U4329 ( .A1(n4492), .A2(n3498), .ZN(n3509) );
  INV_X1 U4330 ( .A(n3509), .ZN(n3525) );
  XNOR2_X1 U4331 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3503) );
  NAND2_X1 U4332 ( .A1(n4955), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3506) );
  INV_X1 U4333 ( .A(n3506), .ZN(n3499) );
  NAND2_X1 U4334 ( .A1(n3503), .A2(n3499), .ZN(n3501) );
  NAND2_X1 U4335 ( .A1(n6345), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3500) );
  NAND2_X1 U4336 ( .A1(n3501), .A2(n3500), .ZN(n3528) );
  XNOR2_X1 U4337 ( .A(n5292), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3526)
         );
  XNOR2_X1 U4338 ( .A(n3528), .B(n3526), .ZN(n3564) );
  NAND2_X1 U4339 ( .A1(n3544), .A2(n3564), .ZN(n3524) );
  NAND2_X1 U4340 ( .A1(n3544), .A2(n3224), .ZN(n3502) );
  NAND2_X1 U4341 ( .A1(n3502), .A2(n3207), .ZN(n3512) );
  INV_X1 U4342 ( .A(n3512), .ZN(n3520) );
  XNOR2_X1 U4343 ( .A(n3503), .B(n3506), .ZN(n3563) );
  AND2_X1 U4344 ( .A1(n3563), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3511) );
  INV_X1 U4345 ( .A(n3511), .ZN(n3519) );
  NAND2_X1 U4346 ( .A1(n3505), .A2(n3504), .ZN(n3551) );
  OAI21_X1 U4347 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4955), .A(n3506), 
        .ZN(n3507) );
  INV_X1 U4348 ( .A(n3507), .ZN(n3514) );
  AOI21_X1 U4349 ( .B1(n3508), .B2(n3514), .A(n4269), .ZN(n3510) );
  OAI22_X1 U4350 ( .A1(n3512), .A2(n3511), .B1(n3510), .B2(n3509), .ZN(n3513)
         );
  OAI21_X1 U4351 ( .B1(n3563), .B2(n3551), .A(n3513), .ZN(n3517) );
  NAND2_X1 U4352 ( .A1(n3544), .A2(n3514), .ZN(n3515) );
  NAND2_X1 U4353 ( .A1(n3515), .A2(n3551), .ZN(n3516) );
  NAND2_X1 U4354 ( .A1(n3517), .A2(n3516), .ZN(n3518) );
  OAI21_X1 U4355 ( .B1(n3520), .B2(n3519), .A(n3518), .ZN(n3522) );
  OAI211_X1 U4356 ( .C1(n3564), .C2(n3539), .A(n3524), .B(n3525), .ZN(n3521)
         );
  NAND2_X1 U4357 ( .A1(n3522), .A2(n3521), .ZN(n3523) );
  OAI21_X1 U4358 ( .B1(n3525), .B2(n3524), .A(n3523), .ZN(n3549) );
  INV_X1 U4359 ( .A(n3526), .ZN(n3527) );
  NAND2_X1 U4360 ( .A1(n3528), .A2(n3527), .ZN(n3530) );
  NAND2_X1 U4361 ( .A1(n6351), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U4362 ( .A1(n3530), .A2(n3529), .ZN(n3535) );
  XNOR2_X1 U4363 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U4364 ( .A1(n3535), .A2(n3533), .ZN(n3532) );
  NAND2_X1 U4365 ( .A1(n6358), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U4366 ( .A1(n3532), .A2(n3531), .ZN(n3541) );
  INV_X1 U4367 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U4368 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6646), .ZN(n3542) );
  OR2_X1 U4369 ( .A1(n3541), .A2(n3542), .ZN(n3537) );
  INV_X1 U4370 ( .A(n3533), .ZN(n3534) );
  XNOR2_X1 U4371 ( .A(n3535), .B(n3534), .ZN(n3536) );
  INV_X1 U4372 ( .A(n3565), .ZN(n3538) );
  NAND2_X1 U4373 ( .A1(n3539), .A2(n3538), .ZN(n3548) );
  INV_X1 U4374 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6355) );
  AND2_X1 U4375 ( .A1(n6355), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3540)
         );
  OR2_X1 U4376 ( .A1(n3541), .A2(n3540), .ZN(n3543) );
  NAND2_X1 U4377 ( .A1(n3544), .A2(n3550), .ZN(n3546) );
  NAND2_X1 U4378 ( .A1(n6379), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3545) );
  OAI211_X1 U4379 ( .C1(n3551), .C2(n3565), .A(n3546), .B(n3545), .ZN(n3547)
         );
  AOI21_X1 U4380 ( .B1(n3549), .B2(n3548), .A(n3547), .ZN(n3553) );
  NOR2_X1 U4381 ( .A1(n3551), .A2(n3566), .ZN(n3552) );
  NAND2_X1 U4382 ( .A1(n3554), .A2(n3207), .ZN(n4419) );
  NOR2_X1 U4383 ( .A1(n4419), .A2(n3222), .ZN(n3593) );
  INV_X1 U4384 ( .A(n3593), .ZN(n3569) );
  INV_X1 U4385 ( .A(n3555), .ZN(n4335) );
  INV_X1 U4386 ( .A(n3582), .ZN(n3557) );
  NAND2_X1 U4387 ( .A1(n4419), .A2(n4269), .ZN(n3556) );
  AND3_X1 U4388 ( .A1(n3557), .A2(n3347), .A3(n3556), .ZN(n3578) );
  NAND2_X1 U4389 ( .A1(n3558), .A2(n4590), .ZN(n3560) );
  INV_X1 U4390 ( .A(n3212), .ZN(n3559) );
  MUX2_X1 U4391 ( .A(n3560), .B(n6488), .S(n3559), .Z(n4416) );
  NAND2_X1 U4392 ( .A1(n3578), .A2(n4416), .ZN(n3561) );
  NAND2_X1 U4393 ( .A1(n4335), .A2(n3561), .ZN(n4401) );
  INV_X1 U4394 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6403) );
  NAND2_X1 U4395 ( .A1(n3562), .A2(n6403), .ZN(n6398) );
  INV_X1 U4396 ( .A(n6398), .ZN(n4327) );
  NAND3_X1 U4397 ( .A1(n3565), .A2(n3564), .A3(n3563), .ZN(n3567) );
  NAND2_X1 U4398 ( .A1(n3567), .A2(n3566), .ZN(n4234) );
  NOR2_X1 U4399 ( .A1(READY_N), .A2(n4234), .ZN(n4405) );
  OAI211_X1 U4400 ( .C1(n3222), .C2(n4327), .A(n3155), .B(n4405), .ZN(n3568)
         );
  OAI211_X1 U4401 ( .C1(n4404), .C2(n3569), .A(n4401), .B(n3568), .ZN(n3571)
         );
  NAND2_X1 U4402 ( .A1(n3570), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6384) );
  INV_X1 U4403 ( .A(n6384), .ZN(n4494) );
  NAND2_X1 U4404 ( .A1(n3571), .A2(n4494), .ZN(n3575) );
  INV_X1 U4405 ( .A(READY_N), .ZN(n6485) );
  AND2_X1 U4406 ( .A1(n4415), .A2(n6485), .ZN(n4394) );
  NAND2_X1 U4407 ( .A1(n3222), .A2(n6398), .ZN(n4270) );
  NAND2_X1 U4408 ( .A1(n4590), .A2(n4500), .ZN(n3572) );
  AOI21_X1 U4409 ( .B1(n4394), .B2(n4270), .A(n3572), .ZN(n3573) );
  AND2_X1 U4410 ( .A1(n3578), .A2(n5082), .ZN(n4403) );
  INV_X1 U4411 ( .A(n4403), .ZN(n4519) );
  NAND2_X1 U4412 ( .A1(n3678), .A2(n4585), .ZN(n3576) );
  NAND2_X1 U4413 ( .A1(n4415), .A2(n4422), .ZN(n4395) );
  AND2_X1 U4414 ( .A1(n3576), .A2(n4395), .ZN(n3579) );
  NAND2_X1 U4415 ( .A1(n3578), .A2(n3577), .ZN(n6360) );
  NAND4_X1 U4416 ( .A1(n4519), .A2(n3579), .A3(n4557), .A4(n6360), .ZN(n3580)
         );
  NAND2_X1 U4417 ( .A1(n3682), .A2(n3580), .ZN(n5805) );
  NAND2_X1 U4418 ( .A1(n3699), .A2(n6129), .ZN(n3698) );
  NOR2_X1 U4419 ( .A1(n6074), .A2(n6066), .ZN(n6061) );
  NAND3_X1 U4420 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6061), .ZN(n3595) );
  NAND2_X1 U4421 ( .A1(n3582), .A2(n5373), .ZN(n3590) );
  NAND2_X1 U4422 ( .A1(n3155), .A2(n4500), .ZN(n3583) );
  AND2_X1 U4423 ( .A1(n3584), .A2(n3583), .ZN(n3588) );
  INV_X4 U4424 ( .A(n5373), .ZN(n5317) );
  OR2_X1 U4425 ( .A1(n5085), .A2(n3155), .ZN(n4400) );
  NAND2_X1 U4426 ( .A1(n2973), .A2(n4400), .ZN(n3586) );
  INV_X1 U4427 ( .A(n3347), .ZN(n3585) );
  NAND2_X1 U4428 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  NAND4_X1 U4429 ( .A1(n3590), .A2(n3589), .A3(n3588), .A4(n3587), .ZN(n4411)
         );
  OAI21_X1 U4430 ( .B1(n4412), .B2(n4590), .A(n4542), .ZN(n3591) );
  NOR2_X1 U4431 ( .A1(n4411), .A2(n3591), .ZN(n3592) );
  AND2_X1 U4432 ( .A1(n3592), .A2(n4416), .ZN(n3596) );
  NAND2_X1 U4433 ( .A1(n3596), .A2(n3593), .ZN(n4520) );
  INV_X1 U4434 ( .A(n4520), .ZN(n4332) );
  NAND2_X1 U4435 ( .A1(n3682), .A2(n4332), .ZN(n6116) );
  INV_X1 U4436 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U4437 ( .B1(n6127), .B2(n6117), .A(n3355), .ZN(n6118) );
  NAND3_X1 U4438 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6118), .ZN(n5120) );
  NOR2_X1 U4439 ( .A1(n6116), .A2(n5120), .ZN(n6086) );
  NAND3_X1 U4440 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6086), .ZN(n5117) );
  NOR2_X1 U4441 ( .A1(n3595), .A2(n5117), .ZN(n3683) );
  NOR2_X1 U4442 ( .A1(n3355), .A2(n6127), .ZN(n6098) );
  NAND3_X1 U4443 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6098), .ZN(n6088) );
  NAND2_X1 U4444 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3594) );
  OR2_X1 U4445 ( .A1(n6088), .A2(n3594), .ZN(n5118) );
  OR2_X1 U4446 ( .A1(n5118), .A2(n3595), .ZN(n3684) );
  INV_X1 U4447 ( .A(n3596), .ZN(n3597) );
  NAND2_X1 U4448 ( .A1(n3682), .A2(n3597), .ZN(n5223) );
  AND2_X1 U4449 ( .A1(n3555), .A2(n3224), .ZN(n4536) );
  NAND2_X1 U4450 ( .A1(n3682), .A2(n4536), .ZN(n5228) );
  NAND2_X1 U4451 ( .A1(n5223), .A2(n5228), .ZN(n6078) );
  NAND2_X1 U4452 ( .A1(n5228), .A2(n6117), .ZN(n4425) );
  NAND2_X1 U4453 ( .A1(n6078), .A2(n4425), .ZN(n6126) );
  NOR2_X1 U4454 ( .A1(n3684), .A2(n6126), .ZN(n6041) );
  NOR2_X1 U4455 ( .A1(n3683), .A2(n6041), .ZN(n5817) );
  INV_X1 U4456 ( .A(n5817), .ZN(n6043) );
  NAND2_X1 U4457 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6042) );
  NOR2_X1 U4458 ( .A1(n3645), .A2(n6042), .ZN(n5229) );
  INV_X1 U4459 ( .A(n5229), .ZN(n5231) );
  NOR2_X1 U4460 ( .A1(n6548), .A2(n5231), .ZN(n3685) );
  NAND3_X1 U4461 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5708), .ZN(n5811) );
  INV_X1 U4462 ( .A(n5811), .ZN(n3598) );
  AND2_X1 U4463 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n3598), .ZN(n5799)
         );
  NAND2_X1 U4464 ( .A1(n5799), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5685) );
  AND2_X1 U4465 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U4466 ( .A1(n5676), .A2(n5655), .ZN(n3599) );
  NOR2_X1 U4467 ( .A1(n5685), .A2(n3599), .ZN(n5643) );
  INV_X1 U4468 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5524) );
  OR2_X1 U4469 ( .A1(n4038), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6123) );
  INV_X1 U4470 ( .A(REIP_REG_23__SCAN_IN), .ZN(n3600) );
  NOR2_X1 U4471 ( .A1(n6123), .A2(n3600), .ZN(n4045) );
  AND2_X1 U4472 ( .A1(n5373), .A2(EBX_REG_1__SCAN_IN), .ZN(n3602) );
  NAND2_X1 U4473 ( .A1(n3605), .A2(n3604), .ZN(n3608) );
  INV_X1 U4474 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U4475 ( .A1(n5373), .A2(n5088), .ZN(n3607) );
  OAI21_X1 U4476 ( .B1(n3606), .B2(n5088), .A(n3607), .ZN(n4365) );
  XNOR2_X1 U4477 ( .A(n3608), .B(n4365), .ZN(n5094) );
  AOI21_X1 U4478 ( .B1(n5094), .B2(n4422), .A(n3608), .ZN(n4437) );
  MUX2_X1 U4479 ( .A(n3609), .B(n5373), .S(EBX_REG_2__SCAN_IN), .Z(n3611) );
  NOR2_X1 U4480 ( .A1(n4304), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3610)
         );
  NOR2_X1 U4481 ( .A1(n3611), .A2(n3610), .ZN(n4436) );
  NAND2_X1 U4482 ( .A1(n4437), .A2(n4436), .ZN(n4509) );
  OR2_X1 U4483 ( .A1(n4300), .A2(EBX_REG_3__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U4484 ( .A1(n3606), .A2(n6099), .ZN(n3613) );
  OAI211_X1 U4485 ( .C1(n3612), .C2(EBX_REG_3__SCAN_IN), .A(n5317), .B(n3613), 
        .ZN(n3614) );
  NAND2_X1 U4486 ( .A1(n5317), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3617)
         );
  OAI211_X1 U4487 ( .C1(n3612), .C2(EBX_REG_4__SCAN_IN), .A(n3606), .B(n3617), 
        .ZN(n3618) );
  OAI21_X1 U4488 ( .B1(n3601), .B2(EBX_REG_4__SCAN_IN), .A(n3618), .ZN(n5920)
         );
  OR2_X1 U4489 ( .A1(n4300), .A2(EBX_REG_5__SCAN_IN), .ZN(n3621) );
  OAI21_X1 U4490 ( .B1(n5373), .B2(n5121), .A(n3606), .ZN(n3619) );
  OAI21_X1 U4491 ( .B1(n3612), .B2(EBX_REG_5__SCAN_IN), .A(n3619), .ZN(n3620)
         );
  NAND2_X1 U4492 ( .A1(n3621), .A2(n3620), .ZN(n4573) );
  INV_X1 U4493 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U4494 ( .A1(n3609), .A2(n5954), .ZN(n3624) );
  NAND2_X1 U4495 ( .A1(n5317), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3622)
         );
  OAI211_X1 U4496 ( .C1(n3612), .C2(EBX_REG_6__SCAN_IN), .A(n3606), .B(n3622), 
        .ZN(n3623) );
  MUX2_X1 U4497 ( .A(n3609), .B(n5373), .S(EBX_REG_8__SCAN_IN), .Z(n3625) );
  INV_X1 U4498 ( .A(n3625), .ZN(n3626) );
  NAND2_X1 U4499 ( .A1(n3626), .A2(n3065), .ZN(n4909) );
  OR2_X1 U4500 ( .A1(n4300), .A2(EBX_REG_7__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U4501 ( .A1(n3606), .A2(n6074), .ZN(n3627) );
  OAI211_X1 U4502 ( .C1(n3612), .C2(EBX_REG_7__SCAN_IN), .A(n5317), .B(n3627), 
        .ZN(n3628) );
  OR2_X1 U4503 ( .A1(n4300), .A2(EBX_REG_9__SCAN_IN), .ZN(n3634) );
  NAND2_X1 U4504 ( .A1(n3606), .A2(n6050), .ZN(n3632) );
  OAI211_X1 U4505 ( .C1(n3612), .C2(EBX_REG_9__SCAN_IN), .A(n5317), .B(n3632), 
        .ZN(n3633) );
  AND2_X1 U4506 ( .A1(n3634), .A2(n3633), .ZN(n5048) );
  MUX2_X1 U4507 ( .A(n3609), .B(n5373), .S(EBX_REG_10__SCAN_IN), .Z(n3636) );
  NOR2_X1 U4508 ( .A1(n4304), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3635)
         );
  NOR2_X1 U4509 ( .A1(n3636), .A2(n3635), .ZN(n5109) );
  OR2_X1 U4510 ( .A1(n4300), .A2(EBX_REG_11__SCAN_IN), .ZN(n3639) );
  INV_X1 U4511 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U4512 ( .A1(n3606), .A2(n5184), .ZN(n3637) );
  OAI211_X1 U4513 ( .C1(n3612), .C2(EBX_REG_11__SCAN_IN), .A(n5317), .B(n3637), 
        .ZN(n3638) );
  AND2_X1 U4514 ( .A1(n3639), .A2(n3638), .ZN(n5168) );
  MUX2_X1 U4515 ( .A(n3609), .B(n5373), .S(EBX_REG_12__SCAN_IN), .Z(n3640) );
  INV_X1 U4516 ( .A(n3640), .ZN(n3641) );
  NAND2_X1 U4517 ( .A1(n3641), .A2(n3066), .ZN(n5176) );
  MUX2_X1 U4518 ( .A(n3609), .B(n5373), .S(EBX_REG_14__SCAN_IN), .Z(n3642) );
  INV_X1 U4519 ( .A(n3642), .ZN(n3644) );
  NAND2_X1 U4520 ( .A1(n2973), .A2(n6548), .ZN(n3643) );
  NAND2_X1 U4521 ( .A1(n3644), .A2(n3643), .ZN(n5206) );
  OR2_X1 U4522 ( .A1(n4300), .A2(EBX_REG_13__SCAN_IN), .ZN(n3648) );
  OAI21_X1 U4523 ( .B1(n5373), .B2(n3645), .A(n3606), .ZN(n3646) );
  OAI21_X1 U4524 ( .B1(n3612), .B2(EBX_REG_13__SCAN_IN), .A(n3646), .ZN(n3647)
         );
  AND2_X1 U4525 ( .A1(n3648), .A2(n3647), .ZN(n5205) );
  NOR2_X1 U4526 ( .A1(n5206), .A2(n5205), .ZN(n3649) );
  OR2_X1 U4527 ( .A1(n4300), .A2(EBX_REG_15__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U4528 ( .A1(n3606), .A2(n5707), .ZN(n3650) );
  OAI211_X1 U4529 ( .C1(n3612), .C2(EBX_REG_15__SCAN_IN), .A(n5317), .B(n3650), 
        .ZN(n3651) );
  NAND2_X1 U4530 ( .A1(n3652), .A2(n3651), .ZN(n5242) );
  NAND2_X1 U4531 ( .A1(n5243), .A2(n5242), .ZN(n5391) );
  NAND2_X1 U4532 ( .A1(n5317), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3653) );
  OAI211_X1 U4533 ( .C1(n3612), .C2(EBX_REG_16__SCAN_IN), .A(n3606), .B(n3653), 
        .ZN(n3654) );
  OAI21_X1 U4534 ( .B1(n3601), .B2(EBX_REG_16__SCAN_IN), .A(n3654), .ZN(n5392)
         );
  OR2_X1 U4535 ( .A1(n4300), .A2(EBX_REG_17__SCAN_IN), .ZN(n3657) );
  INV_X1 U4536 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U4537 ( .A1(n3606), .A2(n6529), .ZN(n3655) );
  OAI211_X1 U4538 ( .C1(n3612), .C2(EBX_REG_17__SCAN_IN), .A(n5317), .B(n3655), 
        .ZN(n3656) );
  AND2_X1 U4539 ( .A1(n3657), .A2(n3656), .ZN(n5445) );
  NAND2_X1 U4540 ( .A1(n5317), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3658) );
  OAI211_X1 U4541 ( .C1(n3612), .C2(EBX_REG_19__SCAN_IN), .A(n3606), .B(n3658), 
        .ZN(n3659) );
  OAI21_X1 U4542 ( .B1(n3601), .B2(EBX_REG_19__SCAN_IN), .A(n3659), .ZN(n5376)
         );
  INV_X1 U4543 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U4544 ( .A1(n2973), .A2(n5803), .ZN(n3660) );
  OR2_X1 U4545 ( .A1(n3612), .A2(EBX_REG_18__SCAN_IN), .ZN(n5372) );
  AND2_X1 U4546 ( .A1(n3660), .A2(n5372), .ZN(n5375) );
  OAI22_X1 U4547 ( .A1(n4304), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n3612), .B2(EBX_REG_20__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U4548 ( .A1(n5375), .A2(n5358), .ZN(n3662) );
  NAND2_X1 U4549 ( .A1(n5373), .A2(EBX_REG_20__SCAN_IN), .ZN(n3661) );
  OAI211_X1 U4550 ( .C1(n5375), .C2(n5373), .A(n3662), .B(n3661), .ZN(n3663)
         );
  INV_X1 U4551 ( .A(n3663), .ZN(n3664) );
  MUX2_X1 U4552 ( .A(n3609), .B(n5373), .S(EBX_REG_21__SCAN_IN), .Z(n3666) );
  NOR2_X1 U4553 ( .A1(n4304), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3665)
         );
  NOR2_X1 U4554 ( .A1(n3666), .A2(n3665), .ZN(n5424) );
  OR2_X1 U4555 ( .A1(n4300), .A2(EBX_REG_22__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4556 ( .A1(n3606), .A2(n5661), .ZN(n3667) );
  OAI211_X1 U4557 ( .C1(n3612), .C2(EBX_REG_22__SCAN_IN), .A(n5317), .B(n3667), 
        .ZN(n3668) );
  NAND2_X1 U4558 ( .A1(n3669), .A2(n3668), .ZN(n5652) );
  INV_X1 U4559 ( .A(n5652), .ZN(n3674) );
  INV_X1 U4560 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U4561 ( .A1(n3609), .A2(n5729), .ZN(n3672) );
  NAND2_X1 U4562 ( .A1(n5317), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3670) );
  OAI211_X1 U4563 ( .C1(n3612), .C2(EBX_REG_23__SCAN_IN), .A(n3606), .B(n3670), 
        .ZN(n3671) );
  AND2_X1 U4564 ( .A1(n3672), .A2(n3671), .ZN(n3675) );
  INV_X1 U4565 ( .A(n3675), .ZN(n3673) );
  OAI21_X1 U4566 ( .B1(n5653), .B2(n3674), .A(n3673), .ZN(n3677) );
  NAND2_X1 U4567 ( .A1(n3675), .A2(n5652), .ZN(n3676) );
  NAND2_X1 U4568 ( .A1(n3677), .A2(n5413), .ZN(n5737) );
  NAND2_X1 U4569 ( .A1(n3678), .A2(n4370), .ZN(n3679) );
  NAND2_X1 U4570 ( .A1(n4415), .A2(n4351), .ZN(n6370) );
  NAND2_X1 U4571 ( .A1(n3679), .A2(n6370), .ZN(n3680) );
  INV_X1 U4572 ( .A(n6121), .ZN(n6089) );
  NOR2_X1 U4573 ( .A1(n5737), .A2(n6089), .ZN(n3681) );
  AOI211_X1 U4574 ( .C1(n5643), .C2(n5524), .A(n4045), .B(n3681), .ZN(n3696)
         );
  NAND2_X1 U4575 ( .A1(n6116), .A2(n5223), .ZN(n5225) );
  AND2_X1 U4576 ( .A1(n6117), .A2(n5225), .ZN(n4377) );
  INV_X2 U4577 ( .A(n6123), .ZN(n6101) );
  NOR2_X1 U4578 ( .A1(n6101), .A2(n3682), .ZN(n4380) );
  NOR2_X1 U4579 ( .A1(n4377), .A2(n4380), .ZN(n4424) );
  NAND2_X1 U4580 ( .A1(n4424), .A2(n6116), .ZN(n5669) );
  INV_X1 U4581 ( .A(n3683), .ZN(n5224) );
  AOI22_X1 U4582 ( .A1(n6078), .A2(n3684), .B1(n5669), .B2(n5224), .ZN(n5227)
         );
  INV_X1 U4583 ( .A(n5228), .ZN(n4381) );
  INV_X1 U4584 ( .A(n3685), .ZN(n3686) );
  NAND2_X1 U4585 ( .A1(n5674), .A2(n3686), .ZN(n3687) );
  NAND2_X1 U4586 ( .A1(n5227), .A2(n3687), .ZN(n5693) );
  NOR2_X1 U4587 ( .A1(n5707), .A2(n5775), .ZN(n5695) );
  INV_X1 U4588 ( .A(n5695), .ZN(n3688) );
  AND2_X1 U4589 ( .A1(n5674), .A2(n3688), .ZN(n3689) );
  OR2_X1 U4590 ( .A1(n5693), .A2(n3689), .ZN(n5808) );
  INV_X1 U4591 ( .A(n3690), .ZN(n3691) );
  NAND2_X1 U4592 ( .A1(n3691), .A2(n5676), .ZN(n5654) );
  AND2_X1 U4593 ( .A1(n5674), .A2(n5654), .ZN(n3692) );
  NOR2_X1 U4594 ( .A1(n5808), .A2(n3692), .ZN(n5668) );
  INV_X1 U4595 ( .A(n5655), .ZN(n3693) );
  NAND2_X1 U4596 ( .A1(n5674), .A2(n3693), .ZN(n3694) );
  AND2_X1 U4597 ( .A1(n5668), .A2(n3694), .ZN(n4293) );
  OR2_X1 U4598 ( .A1(n4293), .A2(n5524), .ZN(n3695) );
  NAND2_X1 U4599 ( .A1(n3698), .A2(n3697), .ZN(U2995) );
  INV_X1 U4600 ( .A(n6011), .ZN(n6035) );
  NAND2_X1 U4601 ( .A1(n3699), .A2(n6035), .ZN(n4050) );
  NAND2_X1 U4602 ( .A1(n3231), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3880) );
  INV_X2 U4603 ( .A(n2980), .ZN(n4227) );
  AOI22_X1 U4604 ( .A1(n4227), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6285), .ZN(n3701) );
  INV_X1 U4605 ( .A(n4500), .ZN(n4503) );
  NAND2_X1 U4606 ( .A1(n4503), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3730) );
  INV_X1 U4607 ( .A(n3730), .ZN(n3707) );
  NAND2_X1 U4608 ( .A1(n3707), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3700) );
  AND2_X1 U4609 ( .A1(n3701), .A2(n3700), .ZN(n3702) );
  INV_X1 U4610 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5829) );
  NAND2_X1 U4611 ( .A1(n6285), .A2(n5829), .ZN(n3731) );
  NAND2_X1 U4612 ( .A1(n4227), .A2(EAX_REG_0__SCAN_IN), .ZN(n3705) );
  NAND2_X1 U4613 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3704)
         );
  OAI211_X1 U4614 ( .C1(n3730), .C2(n3070), .A(n3705), .B(n3704), .ZN(n3706)
         );
  NAND2_X1 U4615 ( .A1(n3707), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3711) );
  OAI21_X1 U4616 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3719), .ZN(n6038) );
  INV_X1 U4617 ( .A(n6038), .ZN(n3708) );
  NAND2_X1 U4618 ( .A1(n6285), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4075) );
  INV_X1 U4619 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5940) );
  OAI22_X1 U4620 ( .A1(n3731), .A2(n3708), .B1(n4075), .B2(n5940), .ZN(n3709)
         );
  AOI21_X1 U4621 ( .B1(n4227), .B2(EAX_REG_2__SCAN_IN), .A(n3709), .ZN(n3710)
         );
  AND2_X1 U4622 ( .A1(n3711), .A2(n3710), .ZN(n4433) );
  INV_X1 U4623 ( .A(n4433), .ZN(n3712) );
  NAND2_X1 U4624 ( .A1(n3713), .A2(n3712), .ZN(n3714) );
  INV_X1 U4625 ( .A(n4575), .ZN(n4734) );
  NAND2_X1 U4626 ( .A1(n3714), .A2(n4434), .ZN(n3716) );
  NAND2_X1 U4627 ( .A1(n4387), .A2(n4433), .ZN(n3715) );
  NAND2_X1 U4628 ( .A1(n3716), .A2(n3715), .ZN(n4432) );
  INV_X1 U4629 ( .A(n4432), .ZN(n3727) );
  INV_X1 U4630 ( .A(n3719), .ZN(n3718) );
  INV_X1 U4631 ( .A(n3733), .ZN(n3722) );
  INV_X1 U4632 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3720) );
  NAND2_X1 U4633 ( .A1(n3720), .A2(n3719), .ZN(n3721) );
  NAND2_X1 U4634 ( .A1(n3722), .A2(n3721), .ZN(n5147) );
  INV_X1 U4635 ( .A(n4075), .ZN(n4226) );
  AOI22_X1 U4636 ( .A1(n5147), .A2(n4212), .B1(n4226), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3724) );
  NAND2_X1 U4637 ( .A1(n4227), .A2(EAX_REG_3__SCAN_IN), .ZN(n3723) );
  OAI211_X1 U4638 ( .C1(n3730), .C2(n4539), .A(n3724), .B(n3723), .ZN(n3725)
         );
  NAND2_X1 U4639 ( .A1(n3727), .A2(n3726), .ZN(n4506) );
  NAND2_X1 U4640 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3729)
         );
  NAND2_X1 U4641 ( .A1(n4227), .A2(EAX_REG_4__SCAN_IN), .ZN(n3728) );
  OAI211_X1 U4642 ( .C1(n3730), .C2(n6646), .A(n3729), .B(n3728), .ZN(n3732)
         );
  NAND2_X1 U4643 ( .A1(n3732), .A2(n3731), .ZN(n3735) );
  OAI21_X1 U4644 ( .B1(n3733), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3742), 
        .ZN(n6029) );
  NAND2_X1 U4645 ( .A1(n6029), .A2(n4212), .ZN(n3734) );
  NAND2_X1 U4646 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  AOI21_X1 U4647 ( .B1(n3737), .B2(n3814), .A(n3736), .ZN(n4662) );
  NAND2_X1 U4648 ( .A1(n3738), .A2(n3814), .ZN(n3741) );
  XNOR2_X1 U4649 ( .A(n3742), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5913) );
  INV_X1 U4650 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4852) );
  OAI22_X1 U4651 ( .A1(n5913), .A2(n3731), .B1(n4075), .B2(n4852), .ZN(n3739)
         );
  AOI21_X1 U4652 ( .B1(n4227), .B2(EAX_REG_5__SCAN_IN), .A(n3739), .ZN(n3740)
         );
  NAND2_X1 U4653 ( .A1(n3741), .A2(n3740), .ZN(n4569) );
  NOR2_X1 U4654 ( .A1(n3743), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3744)
         );
  OR2_X1 U4655 ( .A1(n3753), .A2(n3744), .ZN(n6020) );
  INV_X1 U4656 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4862) );
  INV_X1 U4657 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5902) );
  OAI22_X1 U4658 ( .A1(n2980), .A2(n4862), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5902), .ZN(n3745) );
  MUX2_X1 U4659 ( .A(n6020), .B(n3745), .S(n3731), .Z(n3746) );
  INV_X1 U4660 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4946) );
  XNOR2_X1 U4661 ( .A(n3753), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U4662 ( .A1(n5081), .A2(n4212), .ZN(n3750) );
  NAND2_X1 U4663 ( .A1(n4226), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3749)
         );
  OAI211_X1 U4664 ( .C1(n2980), .C2(n4946), .A(n3750), .B(n3749), .ZN(n3751)
         );
  NAND2_X1 U4665 ( .A1(n4227), .A2(EAX_REG_8__SCAN_IN), .ZN(n3768) );
  XNOR2_X1 U4666 ( .A(n3769), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U4667 ( .A1(n5065), .A2(n4212), .ZN(n3767) );
  AOI22_X1 U4668 ( .A1(n3436), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4669 ( .A1(n3366), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4670 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4188), .B1(n4187), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4671 ( .A1(n4194), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4672 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3763)
         );
  AOI22_X1 U4673 ( .A1(n4168), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4674 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n3371), .B1(n4186), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4675 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n2964), .B1(n4195), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4676 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n4196), .B1(n4169), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3758) );
  NAND4_X1 U4677 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3762)
         );
  NOR2_X1 U4678 ( .A1(n3763), .A2(n3762), .ZN(n3764) );
  OR2_X1 U4679 ( .A1(n3880), .A2(n3764), .ZN(n3766) );
  NAND2_X1 U4680 ( .A1(n4226), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3765)
         );
  NAND4_X1 U4681 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n4908)
         );
  NAND2_X1 U4682 ( .A1(n4905), .A2(n4908), .ZN(n4906) );
  INV_X1 U4683 ( .A(n4906), .ZN(n3785) );
  XNOR2_X1 U4684 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3787), .ZN(n5054) );
  INV_X1 U4685 ( .A(n5054), .ZN(n5128) );
  AOI22_X1 U4686 ( .A1(n4168), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4687 ( .A1(n4187), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4688 ( .A1(n4188), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4689 ( .A1(n3435), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3770) );
  NAND4_X1 U4690 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3779)
         );
  AOI22_X1 U4691 ( .A1(n3366), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4692 ( .A1(n3390), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4693 ( .A1(n2964), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4694 ( .A1(n4196), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3774) );
  NAND4_X1 U4695 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3778)
         );
  NOR2_X1 U4696 ( .A1(n3779), .A2(n3778), .ZN(n3782) );
  NAND2_X1 U4697 ( .A1(n4227), .A2(EAX_REG_9__SCAN_IN), .ZN(n3781) );
  NAND2_X1 U4698 ( .A1(n4226), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3780)
         );
  OAI211_X1 U4699 ( .C1(n3782), .C2(n3880), .A(n3781), .B(n3780), .ZN(n3783)
         );
  AOI21_X1 U4700 ( .B1(n5128), .B2(n4212), .A(n3783), .ZN(n5046) );
  INV_X1 U4701 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3786) );
  XNOR2_X1 U4702 ( .A(n3802), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5162)
         );
  AOI22_X1 U4703 ( .A1(n3436), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4704 ( .A1(n4196), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4705 ( .A1(n2964), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4706 ( .A1(n4168), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3788) );
  NAND4_X1 U4707 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3797)
         );
  AOI22_X1 U4708 ( .A1(n3366), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4709 ( .A1(n4187), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4710 ( .A1(n3435), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4711 ( .A1(n4195), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4712 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3796)
         );
  NOR2_X1 U4713 ( .A1(n3797), .A2(n3796), .ZN(n3800) );
  NAND2_X1 U4714 ( .A1(n4227), .A2(EAX_REG_10__SCAN_IN), .ZN(n3799) );
  NAND2_X1 U4715 ( .A1(n4226), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3798)
         );
  OAI211_X1 U4716 ( .C1(n3800), .C2(n3880), .A(n3799), .B(n3798), .ZN(n3801)
         );
  AOI21_X1 U4717 ( .B1(n5162), .B2(n4212), .A(n3801), .ZN(n5105) );
  NAND2_X1 U4718 ( .A1(n3802), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3817)
         );
  XNOR2_X1 U4719 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3817), .ZN(n6006)
         );
  AOI22_X1 U4720 ( .A1(n3366), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4721 ( .A1(n4187), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4722 ( .A1(n4196), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4723 ( .A1(n3390), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4724 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3812)
         );
  AOI22_X1 U4725 ( .A1(n4168), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4726 ( .A1(n4541), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4727 ( .A1(n3435), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4728 ( .A1(n4188), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4729 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3811)
         );
  OR2_X1 U4730 ( .A1(n3812), .A2(n3811), .ZN(n3813) );
  AOI22_X1 U4731 ( .A1(n3814), .A2(n3813), .B1(n4226), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3816) );
  NAND2_X1 U4732 ( .A1(n4227), .A2(EAX_REG_11__SCAN_IN), .ZN(n3815) );
  OAI211_X1 U4733 ( .C1(n6006), .C2(n3731), .A(n3816), .B(n3815), .ZN(n5145)
         );
  INV_X1 U4734 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5888) );
  XNOR2_X1 U4735 ( .A(n3834), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5879)
         );
  INV_X1 U4736 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5877) );
  NOR2_X1 U4737 ( .A1(n5877), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3818) );
  AOI21_X1 U4738 ( .B1(n4227), .B2(EAX_REG_12__SCAN_IN), .A(n3818), .ZN(n3830)
         );
  AOI22_X1 U4739 ( .A1(n3390), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4740 ( .A1(n2964), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4741 ( .A1(n3436), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4742 ( .A1(n4188), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4743 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3828)
         );
  AOI22_X1 U4744 ( .A1(n4168), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3366), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4745 ( .A1(n4187), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4746 ( .A1(n4196), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4747 ( .A1(n3435), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4748 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3827)
         );
  NOR2_X1 U4749 ( .A1(n3828), .A2(n3827), .ZN(n3829) );
  OAI22_X1 U4750 ( .A1(n3830), .A2(n4212), .B1(n3829), .B2(n3880), .ZN(n3831)
         );
  AOI21_X1 U4751 ( .B1(n5879), .B2(n4212), .A(n3831), .ZN(n5173) );
  INV_X1 U4752 ( .A(n5173), .ZN(n3832) );
  NAND2_X1 U4753 ( .A1(n3833), .A2(n3832), .ZN(n3839) );
  NAND2_X1 U4754 ( .A1(n4227), .A2(EAX_REG_13__SCAN_IN), .ZN(n3837) );
  OAI21_X1 U4755 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3835), .A(n3866), 
        .ZN(n5875) );
  AOI22_X1 U4756 ( .A1(n4212), .A2(n5875), .B1(n4226), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3836) );
  AND2_X1 U4757 ( .A1(n3837), .A2(n3836), .ZN(n3838) );
  OR2_X2 U4758 ( .A1(n3839), .A2(n3838), .ZN(n3852) );
  NAND2_X1 U4759 ( .A1(n3839), .A2(n3838), .ZN(n3840) );
  AOI22_X1 U4760 ( .A1(n3366), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4761 ( .A1(n4196), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4762 ( .A1(n4187), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4763 ( .A1(n4168), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4764 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3850)
         );
  AOI22_X1 U4765 ( .A1(n3436), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4766 ( .A1(n4186), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4767 ( .A1(n3435), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4768 ( .A1(n4195), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3845) );
  NAND4_X1 U4769 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3849)
         );
  NOR2_X1 U4770 ( .A1(n3850), .A2(n3849), .ZN(n3851) );
  NOR2_X1 U4771 ( .A1(n3880), .A2(n3851), .ZN(n5195) );
  AOI22_X1 U4772 ( .A1(n4168), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4773 ( .A1(n4196), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4774 ( .A1(n3435), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4775 ( .A1(n3366), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4776 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3862)
         );
  AOI22_X1 U4777 ( .A1(n4541), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4778 ( .A1(n4187), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4779 ( .A1(n3390), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4780 ( .A1(n2964), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4781 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  NOR2_X1 U4782 ( .A1(n3862), .A2(n3861), .ZN(n3865) );
  NAND2_X1 U4783 ( .A1(n4227), .A2(EAX_REG_14__SCAN_IN), .ZN(n3864) );
  XNOR2_X1 U4784 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3866), .ZN(n5211)
         );
  INV_X1 U4785 ( .A(n5211), .ZN(n5590) );
  AOI22_X1 U4786 ( .A1(n4212), .A2(n5590), .B1(n4226), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3863) );
  OAI211_X1 U4787 ( .C1(n3880), .C2(n3865), .A(n3864), .B(n3863), .ZN(n5199)
         );
  INV_X1 U4788 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5204) );
  INV_X1 U4789 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3867) );
  XNOR2_X1 U4790 ( .A(n3883), .B(n3867), .ZN(n5584) );
  AOI22_X1 U4791 ( .A1(n4196), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4792 ( .A1(n4541), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4793 ( .A1(n3390), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4794 ( .A1(n3969), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3868) );
  NAND4_X1 U4795 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3877)
         );
  AOI22_X1 U4796 ( .A1(n4168), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4797 ( .A1(n3366), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4798 ( .A1(n2964), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4799 ( .A1(n3435), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3872) );
  NAND4_X1 U4800 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3876)
         );
  NOR2_X1 U4801 ( .A1(n3877), .A2(n3876), .ZN(n3881) );
  NAND2_X1 U4802 ( .A1(n4227), .A2(EAX_REG_15__SCAN_IN), .ZN(n3879) );
  NAND2_X1 U4803 ( .A1(n4226), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3878)
         );
  OAI211_X1 U4804 ( .C1(n3881), .C2(n3880), .A(n3879), .B(n3878), .ZN(n3882)
         );
  AOI21_X1 U4805 ( .B1(n5584), .B2(n4212), .A(n3882), .ZN(n5237) );
  XOR2_X1 U4806 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3896), .Z(n5576) );
  AOI22_X1 U4807 ( .A1(n4227), .A2(EAX_REG_16__SCAN_IN), .B1(n4226), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4808 ( .A1(n3366), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4809 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n4196), .B1(n4188), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4810 ( .A1(n4168), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4811 ( .A1(n4187), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3884) );
  NAND4_X1 U4812 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3893)
         );
  AOI22_X1 U4813 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3436), .B1(n3390), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4814 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n3969), .B1(n4186), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4815 ( .A1(n2964), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4816 ( .A1(n3435), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3888) );
  NAND4_X1 U4817 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3892)
         );
  NOR2_X1 U4818 ( .A1(n4419), .A2(n6379), .ZN(n4180) );
  OAI21_X1 U4819 ( .B1(n3893), .B2(n3892), .A(n4180), .ZN(n3894) );
  OAI211_X1 U4820 ( .C1(n5576), .C2(n3731), .A(n3895), .B(n3894), .ZN(n5384)
         );
  NAND2_X1 U4821 ( .A1(n3896), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3914)
         );
  INV_X1 U4822 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5854) );
  OR2_X1 U4823 ( .A1(n3897), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3898)
         );
  NAND2_X1 U4824 ( .A1(n3898), .A2(n3947), .ZN(n5848) );
  INV_X1 U4825 ( .A(n4180), .ZN(n4207) );
  AOI22_X1 U4826 ( .A1(n3435), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4827 ( .A1(n4196), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4828 ( .A1(n3366), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4829 ( .A1(n2964), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4830 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3908)
         );
  AOI22_X1 U4831 ( .A1(n4168), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4832 ( .A1(n3390), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4833 ( .A1(n3969), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4834 ( .A1(n4194), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4835 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3907)
         );
  NOR2_X1 U4836 ( .A1(n3908), .A2(n3907), .ZN(n3909) );
  NOR2_X1 U4837 ( .A1(n4207), .A2(n3909), .ZN(n3913) );
  INV_X1 U4838 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U4839 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3910)
         );
  OAI211_X1 U4840 ( .C1(n2980), .C2(n3911), .A(n3731), .B(n3910), .ZN(n3912)
         );
  OAI22_X1 U4841 ( .A1(n5848), .A2(n3731), .B1(n3913), .B2(n3912), .ZN(n5432)
         );
  XNOR2_X1 U4842 ( .A(n3914), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5856)
         );
  NAND2_X1 U4843 ( .A1(n5856), .A2(n4212), .ZN(n3929) );
  AOI22_X1 U4844 ( .A1(n4168), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4845 ( .A1(n4187), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4846 ( .A1(n4196), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4847 ( .A1(n2964), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3915) );
  NAND4_X1 U4848 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(n3924)
         );
  AOI22_X1 U4849 ( .A1(n3436), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4850 ( .A1(n3366), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4851 ( .A1(n4194), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4852 ( .A1(n4195), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3919) );
  NAND4_X1 U4853 ( .A1(n3922), .A2(n3921), .A3(n3920), .A4(n3919), .ZN(n3923)
         );
  NOR2_X1 U4854 ( .A1(n3924), .A2(n3923), .ZN(n3927) );
  AOI21_X1 U4855 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5854), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3925) );
  AOI21_X1 U4856 ( .B1(n4227), .B2(EAX_REG_17__SCAN_IN), .A(n3925), .ZN(n3926)
         );
  OAI21_X1 U4857 ( .B1(n4207), .B2(n3927), .A(n3926), .ZN(n3928) );
  NAND2_X1 U4858 ( .A1(n3929), .A2(n3928), .ZN(n5444) );
  OR2_X1 U4859 ( .A1(n5432), .A2(n5444), .ZN(n5366) );
  AOI22_X1 U4860 ( .A1(n4168), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3436), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4861 ( .A1(n3366), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4862 ( .A1(n4196), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4863 ( .A1(n3435), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U4864 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3939)
         );
  AOI22_X1 U4865 ( .A1(n4187), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4866 ( .A1(n4541), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4867 ( .A1(n2964), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4868 ( .A1(n4188), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3934) );
  NAND4_X1 U4869 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(n3938)
         );
  NOR2_X1 U4870 ( .A1(n3939), .A2(n3938), .ZN(n3943) );
  NAND2_X1 U4871 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3940)
         );
  NAND2_X1 U4872 ( .A1(n3731), .A2(n3940), .ZN(n3941) );
  AOI21_X1 U4873 ( .B1(n4227), .B2(EAX_REG_19__SCAN_IN), .A(n3941), .ZN(n3942)
         );
  OAI21_X1 U4874 ( .B1(n4207), .B2(n3943), .A(n3942), .ZN(n3945) );
  XNOR2_X1 U4875 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3947), .ZN(n5562)
         );
  NAND2_X1 U4876 ( .A1(n4212), .A2(n5562), .ZN(n3944) );
  NAND2_X1 U4877 ( .A1(n3945), .A2(n3944), .ZN(n5369) );
  INV_X1 U4878 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3946) );
  OR2_X1 U4879 ( .A1(n3948), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3949)
         );
  NAND2_X1 U4880 ( .A1(n3948), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3979)
         );
  NAND2_X1 U4881 ( .A1(n3949), .A2(n3979), .ZN(n5555) );
  INV_X1 U4882 ( .A(n5555), .ZN(n5360) );
  AOI22_X1 U4883 ( .A1(n3366), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4884 ( .A1(n4196), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4885 ( .A1(n3436), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4886 ( .A1(n4186), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3950) );
  NAND4_X1 U4887 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3959)
         );
  AOI22_X1 U4888 ( .A1(n4168), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4889 ( .A1(n4187), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4890 ( .A1(n3435), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4891 ( .A1(n2964), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U4892 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3958)
         );
  OR2_X1 U4893 ( .A1(n3959), .A2(n3958), .ZN(n3963) );
  INV_X1 U4894 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3961) );
  NAND2_X1 U4895 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3960)
         );
  OAI211_X1 U4896 ( .C1(n2980), .C2(n3961), .A(n3731), .B(n3960), .ZN(n3962)
         );
  AOI21_X1 U4897 ( .B1(n4180), .B2(n3963), .A(n3962), .ZN(n3964) );
  AOI21_X1 U4898 ( .B1(n5360), .B2(n4212), .A(n3964), .ZN(n5356) );
  AOI22_X1 U4899 ( .A1(n3186), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3366), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4900 ( .A1(n4196), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4901 ( .A1(n3435), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4902 ( .A1(n2964), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3965) );
  NAND4_X1 U4903 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3975)
         );
  AOI22_X1 U4904 ( .A1(n3390), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4905 ( .A1(n4187), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4906 ( .A1(n3969), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4907 ( .A1(n3436), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4908 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3974)
         );
  NOR2_X1 U4909 ( .A1(n3975), .A2(n3974), .ZN(n3978) );
  INV_X1 U4910 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6571) );
  OAI21_X1 U4911 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6571), .A(n3731), .ZN(
        n3976) );
  AOI21_X1 U4912 ( .B1(n4227), .B2(EAX_REG_21__SCAN_IN), .A(n3976), .ZN(n3977)
         );
  OAI21_X1 U4913 ( .B1(n4207), .B2(n3978), .A(n3977), .ZN(n3983) );
  NOR2_X1 U4914 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3980), .ZN(n3981)
         );
  NOR2_X1 U4915 ( .A1(n3998), .A2(n3981), .ZN(n5748) );
  NAND2_X1 U4916 ( .A1(n5748), .A2(n4212), .ZN(n3982) );
  NAND2_X1 U4917 ( .A1(n3983), .A2(n3982), .ZN(n5537) );
  AOI22_X1 U4918 ( .A1(n4168), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4919 ( .A1(n4187), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4920 ( .A1(n3194), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4921 ( .A1(n4196), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3984) );
  NAND4_X1 U4922 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(n3993)
         );
  AOI22_X1 U4923 ( .A1(n3390), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4924 ( .A1(n3366), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4925 ( .A1(n4188), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4926 ( .A1(n3436), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3988) );
  NAND4_X1 U4927 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n3988), .ZN(n3992)
         );
  NOR2_X1 U4928 ( .A1(n3993), .A2(n3992), .ZN(n3997) );
  OAI21_X1 U4929 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5829), .A(n6285), 
        .ZN(n3994) );
  INV_X1 U4930 ( .A(n3994), .ZN(n3995) );
  AOI21_X1 U4931 ( .B1(n4227), .B2(EAX_REG_22__SCAN_IN), .A(n3995), .ZN(n3996)
         );
  OAI21_X1 U4932 ( .B1(n4207), .B2(n3997), .A(n3996), .ZN(n4004) );
  INV_X1 U4933 ( .A(n4057), .ZN(n4002) );
  INV_X1 U4934 ( .A(n3998), .ZN(n4000) );
  INV_X1 U4935 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3999) );
  NAND2_X1 U4936 ( .A1(n4000), .A2(n3999), .ZN(n4001) );
  NAND2_X1 U4937 ( .A1(n4002), .A2(n4001), .ZN(n5738) );
  OR2_X1 U4938 ( .A1(n5738), .A2(n3731), .ZN(n4003) );
  NAND2_X1 U4939 ( .A1(n4004), .A2(n4003), .ZN(n5536) );
  AOI22_X1 U4940 ( .A1(n3366), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4941 ( .A1(n2964), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4942 ( .A1(n4168), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4943 ( .A1(n4196), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U4944 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4015)
         );
  AOI22_X1 U4945 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3436), .B1(n3390), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4946 ( .A1(n4541), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4947 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4188), .B1(n4195), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4948 ( .A1(n3435), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4949 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4014)
         );
  NOR2_X1 U4950 ( .A1(n4015), .A2(n4014), .ZN(n4060) );
  AOI22_X1 U4951 ( .A1(n3436), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4952 ( .A1(n2964), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3969), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4953 ( .A1(n4168), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4954 ( .A1(n4195), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U4955 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4025)
         );
  AOI22_X1 U4956 ( .A1(n3390), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4957 ( .A1(n4196), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4958 ( .A1(n3366), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4959 ( .A1(n3435), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U4960 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4024)
         );
  NOR2_X1 U4961 ( .A1(n4025), .A2(n4024), .ZN(n4059) );
  XOR2_X1 U4962 ( .A(n4060), .B(n4059), .Z(n4026) );
  NAND2_X1 U4963 ( .A1(n4180), .A2(n4026), .ZN(n4030) );
  NAND2_X1 U4964 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4027)
         );
  NAND2_X1 U4965 ( .A1(n3731), .A2(n4027), .ZN(n4028) );
  AOI21_X1 U4966 ( .B1(n4227), .B2(EAX_REG_23__SCAN_IN), .A(n4028), .ZN(n4029)
         );
  NAND2_X1 U4967 ( .A1(n4030), .A2(n4029), .ZN(n4033) );
  INV_X1 U4968 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4031) );
  XNOR2_X1 U4969 ( .A(n4057), .B(n4031), .ZN(n5735) );
  NAND2_X1 U4970 ( .A1(n5735), .A2(n4212), .ZN(n4032) );
  NAND2_X1 U4971 ( .A1(n4033), .A2(n4032), .ZN(n4034) );
  AND2_X1 U4972 ( .A1(n4035), .A2(n4034), .ZN(n4036) );
  OR2_X1 U4973 ( .A1(n4036), .A2(n4079), .ZN(n5732) );
  NAND3_X1 U4974 ( .A1(n6379), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6391) );
  INV_X1 U4975 ( .A(n6391), .ZN(n4037) );
  NOR2_X2 U4976 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6284) );
  NAND2_X1 U4977 ( .A1(n4037), .A2(n6284), .ZN(n5579) );
  INV_X1 U4978 ( .A(n6284), .ZN(n6235) );
  NAND2_X1 U4979 ( .A1(n6235), .A2(n4038), .ZN(n6484) );
  NAND2_X1 U4980 ( .A1(n6484), .A2(n6379), .ZN(n4039) );
  NAND2_X1 U4981 ( .A1(n6011), .A2(n4039), .ZN(n5574) );
  NAND2_X1 U4982 ( .A1(n6379), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U4983 ( .A1(n5829), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4040) );
  AND2_X1 U4984 ( .A1(n4041), .A2(n4040), .ZN(n4344) );
  INV_X1 U4985 ( .A(n4344), .ZN(n4042) );
  NAND2_X1 U4986 ( .A1(n5574), .A2(n4042), .ZN(n6039) );
  INV_X1 U4987 ( .A(n5735), .ZN(n4043) );
  NOR2_X1 U4988 ( .A1(n6039), .A2(n4043), .ZN(n4044) );
  AOI211_X1 U4989 ( .C1(n6030), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4045), 
        .B(n4044), .ZN(n4046) );
  INV_X1 U4990 ( .A(n4046), .ZN(n4047) );
  NAND2_X1 U4991 ( .A1(n4050), .A2(n4049), .ZN(U2963) );
  AND2_X1 U4992 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4296) );
  NAND3_X1 U4993 ( .A1(n5676), .A2(n4296), .A3(n5655), .ZN(n4051) );
  NAND2_X1 U4994 ( .A1(n5581), .A2(n4051), .ZN(n4053) );
  NOR2_X1 U4995 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5677) );
  NOR2_X1 U4996 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5656) );
  INV_X1 U4997 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5529) );
  AND4_X1 U4998 ( .A1(n5677), .A2(n5656), .A3(n5524), .A4(n5529), .ZN(n4052)
         );
  XNOR2_X1 U4999 ( .A(n5581), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5519)
         );
  INV_X1 U5000 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U5001 ( .A1(n5581), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5509) );
  AND2_X1 U5002 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U5003 ( .A1(n5616), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5595) );
  NOR2_X1 U5004 ( .A1(n5581), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5508)
         );
  NOR2_X1 U5005 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U5006 ( .A1(n5508), .A2(n5615), .ZN(n5482) );
  NOR2_X1 U5007 ( .A1(n5482), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4054)
         );
  AND2_X1 U5008 ( .A1(n5481), .A2(n4054), .ZN(n4055) );
  OR2_X1 U5009 ( .A1(n4216), .A2(n4055), .ZN(n4056) );
  XNOR2_X1 U5010 ( .A(n4056), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5602)
         );
  INV_X1 U5011 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6634) );
  INV_X1 U5012 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U5013 ( .A1(n4159), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4165)
         );
  INV_X1 U5014 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5326) );
  XNOR2_X1 U5015 ( .A(n4222), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4262)
         );
  INV_X1 U5016 ( .A(n6039), .ZN(n6007) );
  INV_X1 U5017 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U5018 ( .A1(n6101), .A2(REIP_REG_30__SCAN_IN), .ZN(n5597) );
  OAI21_X1 U5019 ( .B1(n5574), .B2(n6586), .A(n5597), .ZN(n4058) );
  AOI21_X1 U5020 ( .B1(n4262), .B2(n6007), .A(n4058), .ZN(n4215) );
  OR2_X1 U5021 ( .A1(n4060), .A2(n4059), .ZN(n4093) );
  AOI22_X1 U5022 ( .A1(n3366), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4196), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5023 ( .A1(n4188), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5024 ( .A1(n4168), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5025 ( .A1(n4187), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4061) );
  NAND4_X1 U5026 ( .A1(n4064), .A2(n4063), .A3(n4062), .A4(n4061), .ZN(n4070)
         );
  AOI22_X1 U5027 ( .A1(n3390), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5028 ( .A1(n3436), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5029 ( .A1(n3435), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5030 ( .A1(n3969), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4065) );
  NAND4_X1 U5031 ( .A1(n4068), .A2(n4067), .A3(n4066), .A4(n4065), .ZN(n4069)
         );
  NOR2_X1 U5032 ( .A1(n4070), .A2(n4069), .ZN(n4092) );
  XNOR2_X1 U5033 ( .A(n4093), .B(n4092), .ZN(n4078) );
  NAND2_X1 U5034 ( .A1(n4071), .A2(n6634), .ZN(n4073) );
  INV_X1 U5035 ( .A(n4072), .ZN(n4080) );
  NAND2_X1 U5036 ( .A1(n4073), .A2(n4080), .ZN(n5532) );
  NAND2_X1 U5037 ( .A1(n5532), .A2(n4212), .ZN(n4074) );
  OAI21_X1 U5038 ( .B1(n6634), .B2(n4075), .A(n4074), .ZN(n4076) );
  AOI21_X1 U5039 ( .B1(n4227), .B2(EAX_REG_24__SCAN_IN), .A(n4076), .ZN(n4077)
         );
  OAI21_X1 U5040 ( .B1(n4078), .B2(n4207), .A(n4077), .ZN(n5347) );
  XNOR2_X1 U5041 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4080), .ZN(n5721)
         );
  AOI22_X1 U5042 ( .A1(n4168), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5043 ( .A1(n3436), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5044 ( .A1(n3366), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5045 ( .A1(n4194), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4082) );
  NAND4_X1 U5046 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4091)
         );
  AOI22_X1 U5047 ( .A1(n4187), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5048 ( .A1(n4196), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5049 ( .A1(n2964), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3969), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5050 ( .A1(n4195), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4086) );
  NAND4_X1 U5051 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4090)
         );
  NOR2_X1 U5052 ( .A1(n4091), .A2(n4090), .ZN(n4100) );
  OR2_X1 U5053 ( .A1(n4093), .A2(n4092), .ZN(n4099) );
  XOR2_X1 U5054 ( .A(n4100), .B(n4099), .Z(n4094) );
  NAND2_X1 U5055 ( .A1(n4094), .A2(n4180), .ZN(n4096) );
  AOI22_X1 U5056 ( .A1(n4227), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6285), .ZN(n4095) );
  NAND2_X1 U5057 ( .A1(n4096), .A2(n4095), .ZN(n4097) );
  NAND2_X1 U5058 ( .A1(n4097), .A2(n3731), .ZN(n4098) );
  OAI21_X1 U5059 ( .B1(n5721), .B2(n3731), .A(n4098), .ZN(n5412) );
  NOR2_X1 U5060 ( .A1(n4100), .A2(n4099), .ZN(n4124) );
  AOI22_X1 U5061 ( .A1(n3186), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5062 ( .A1(n3436), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5063 ( .A1(n3366), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5064 ( .A1(n4194), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U5065 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4110)
         );
  AOI22_X1 U5066 ( .A1(n4187), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5067 ( .A1(n4196), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5068 ( .A1(n2964), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5069 ( .A1(n4195), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4105) );
  NAND4_X1 U5070 ( .A1(n4108), .A2(n4107), .A3(n4106), .A4(n4105), .ZN(n4109)
         );
  OR2_X1 U5071 ( .A1(n4110), .A2(n4109), .ZN(n4123) );
  INV_X1 U5072 ( .A(n4123), .ZN(n4111) );
  XNOR2_X1 U5073 ( .A(n4124), .B(n4111), .ZN(n4115) );
  INV_X1 U5074 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4113) );
  NAND2_X1 U5075 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4112)
         );
  OAI211_X1 U5076 ( .C1(n2980), .C2(n4113), .A(n3731), .B(n4112), .ZN(n4114)
         );
  AOI21_X1 U5077 ( .B1(n4115), .B2(n4180), .A(n4114), .ZN(n4121) );
  INV_X1 U5078 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4118) );
  INV_X1 U5079 ( .A(n4116), .ZN(n4117) );
  NAND2_X1 U5080 ( .A1(n4118), .A2(n4117), .ZN(n4119) );
  NAND2_X1 U5081 ( .A1(n4140), .A2(n4119), .ZN(n5711) );
  NOR2_X1 U5082 ( .A1(n5711), .A2(n3731), .ZN(n4120) );
  NAND2_X1 U5083 ( .A1(n4124), .A2(n4123), .ZN(n4143) );
  AOI22_X1 U5084 ( .A1(n3366), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5085 ( .A1(n4186), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n2964), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5086 ( .A1(n4196), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5087 ( .A1(n3436), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4125) );
  NAND4_X1 U5088 ( .A1(n4128), .A2(n4127), .A3(n4126), .A4(n4125), .ZN(n4134)
         );
  AOI22_X1 U5089 ( .A1(n4168), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5090 ( .A1(n4187), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5091 ( .A1(n3194), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5092 ( .A1(n4188), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4129) );
  NAND4_X1 U5093 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4133)
         );
  NOR2_X1 U5094 ( .A1(n4134), .A2(n4133), .ZN(n4144) );
  XOR2_X1 U5095 ( .A(n4143), .B(n4144), .Z(n4135) );
  NAND2_X1 U5096 ( .A1(n4135), .A2(n4180), .ZN(n4139) );
  NAND2_X1 U5097 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4136)
         );
  NAND2_X1 U5098 ( .A1(n3731), .A2(n4136), .ZN(n4137) );
  AOI21_X1 U5099 ( .B1(n4227), .B2(EAX_REG_27__SCAN_IN), .A(n4137), .ZN(n4138)
         );
  NAND2_X1 U5100 ( .A1(n4139), .A2(n4138), .ZN(n4142) );
  XNOR2_X1 U5101 ( .A(n4140), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5502)
         );
  NAND2_X1 U5102 ( .A1(n5502), .A2(n4212), .ZN(n4141) );
  NAND2_X1 U5103 ( .A1(n4142), .A2(n4141), .ZN(n4312) );
  NOR2_X1 U5104 ( .A1(n4144), .A2(n4143), .ZN(n4167) );
  AOI22_X1 U5105 ( .A1(n3186), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5106 ( .A1(n3436), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5107 ( .A1(n3366), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5108 ( .A1(n4194), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4145) );
  NAND4_X1 U5109 ( .A1(n4148), .A2(n4147), .A3(n4146), .A4(n4145), .ZN(n4154)
         );
  AOI22_X1 U5110 ( .A1(n4187), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5111 ( .A1(n4196), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5112 ( .A1(n2964), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3969), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5113 ( .A1(n4195), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4149) );
  NAND4_X1 U5114 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4153)
         );
  OR2_X1 U5115 ( .A1(n4154), .A2(n4153), .ZN(n4166) );
  INV_X1 U5116 ( .A(n4166), .ZN(n4155) );
  XNOR2_X1 U5117 ( .A(n4167), .B(n4155), .ZN(n4156) );
  NAND2_X1 U5118 ( .A1(n4156), .A2(n4180), .ZN(n4164) );
  NAND2_X1 U5119 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4157)
         );
  NAND2_X1 U5120 ( .A1(n3731), .A2(n4157), .ZN(n4158) );
  AOI21_X1 U5121 ( .B1(n4227), .B2(EAX_REG_28__SCAN_IN), .A(n4158), .ZN(n4163)
         );
  INV_X1 U5122 ( .A(n4159), .ZN(n4160) );
  INV_X1 U5123 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U5124 ( .A1(n4160), .A2(n5338), .ZN(n4161) );
  NAND2_X1 U5125 ( .A1(n4165), .A2(n4161), .ZN(n5491) );
  NOR2_X1 U5126 ( .A1(n5491), .A2(n3731), .ZN(n4162) );
  AOI21_X1 U5127 ( .B1(n4164), .B2(n4163), .A(n4162), .ZN(n5333) );
  XOR2_X1 U5128 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .B(n4165), .Z(n5486) );
  INV_X1 U5129 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4184) );
  NAND2_X1 U5130 ( .A1(n4167), .A2(n4166), .ZN(n4203) );
  AOI22_X1 U5131 ( .A1(n3436), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5132 ( .A1(n3366), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4187), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5133 ( .A1(n4168), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4194), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5134 ( .A1(n4188), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4170) );
  NAND4_X1 U5135 ( .A1(n4173), .A2(n4172), .A3(n4171), .A4(n4170), .ZN(n4179)
         );
  AOI22_X1 U5136 ( .A1(n3390), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5137 ( .A1(n2964), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5138 ( .A1(n4196), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5139 ( .A1(n3435), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4174) );
  NAND4_X1 U5140 ( .A1(n4177), .A2(n4176), .A3(n4175), .A4(n4174), .ZN(n4178)
         );
  NOR2_X1 U5141 ( .A1(n4179), .A2(n4178), .ZN(n4204) );
  XOR2_X1 U5142 ( .A(n4203), .B(n4204), .Z(n4181) );
  NAND2_X1 U5143 ( .A1(n4181), .A2(n4180), .ZN(n4183) );
  AOI21_X1 U5144 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6285), .A(n4212), 
        .ZN(n4182) );
  OAI211_X1 U5145 ( .C1(n2980), .C2(n4184), .A(n4183), .B(n4182), .ZN(n4185)
         );
  OAI21_X1 U5146 ( .B1(n3028), .B2(n5486), .A(n4185), .ZN(n5316) );
  NOR2_X2 U5147 ( .A1(n5314), .A2(n5316), .ZN(n4213) );
  OAI21_X1 U5148 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6586), .A(n3731), .ZN(
        n4210) );
  AOI22_X1 U5149 ( .A1(n3366), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5150 ( .A1(n4187), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4186), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5151 ( .A1(n2964), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3371), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U5152 ( .A1(n4188), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4169), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4189) );
  NAND4_X1 U5153 ( .A1(n4192), .A2(n4191), .A3(n4190), .A4(n4189), .ZN(n4202)
         );
  AOI22_X1 U5154 ( .A1(n3186), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5155 ( .A1(n3436), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4541), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U5156 ( .A1(n4194), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4193), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5157 ( .A1(n4196), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4195), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4197) );
  NAND4_X1 U5158 ( .A1(n4200), .A2(n4199), .A3(n4198), .A4(n4197), .ZN(n4201)
         );
  NOR2_X1 U5159 ( .A1(n4202), .A2(n4201), .ZN(n4206) );
  NOR2_X1 U5160 ( .A1(n4204), .A2(n4203), .ZN(n4205) );
  XOR2_X1 U5161 ( .A(n4206), .B(n4205), .Z(n4208) );
  NOR2_X1 U5162 ( .A1(n4208), .A2(n4207), .ZN(n4209) );
  AOI211_X1 U5163 ( .C1(n4227), .C2(EAX_REG_30__SCAN_IN), .A(n4210), .B(n4209), 
        .ZN(n4211) );
  AOI21_X1 U5164 ( .B1(n4212), .B2(n4262), .A(n4211), .ZN(n4214) );
  NAND2_X1 U5165 ( .A1(n4216), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4220) );
  NOR4_X1 U5166 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A3(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4218) );
  NOR2_X1 U5167 ( .A1(n4222), .A2(n6586), .ZN(n4223) );
  XNOR2_X1 U5168 ( .A(n4223), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4260)
         );
  INV_X1 U5169 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6454) );
  NOR2_X1 U5170 ( .A1(n6123), .A2(n6454), .ZN(n4299) );
  AOI21_X1 U5171 ( .B1(n6030), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4299), 
        .ZN(n4224) );
  OAI21_X1 U5172 ( .B1(n6039), .B2(n4260), .A(n4224), .ZN(n4225) );
  INV_X1 U5173 ( .A(n4225), .ZN(n4232) );
  AOI22_X1 U5174 ( .A1(n4227), .A2(EAX_REG_31__SCAN_IN), .B1(n4226), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4228) );
  INV_X1 U5175 ( .A(n4228), .ZN(n4229) );
  XNOR2_X2 U5176 ( .A(n4230), .B(n4229), .ZN(n5460) );
  NAND2_X1 U5177 ( .A1(n5460), .A2(n2963), .ZN(n4231) );
  INV_X1 U5178 ( .A(n4326), .ZN(n4329) );
  INV_X1 U5179 ( .A(n4234), .ZN(n4336) );
  NAND2_X1 U5180 ( .A1(n3555), .A2(n4336), .ZN(n4324) );
  INV_X1 U5181 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U5182 ( .A1(n6374), .A2(n6285), .ZN(n6390) );
  NOR3_X1 U5183 ( .A1(n6379), .A2(n6464), .A3(n6390), .ZN(n6375) );
  NOR3_X1 U5184 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6374), .A3(n3731), .ZN(
        n6386) );
  NOR2_X1 U5185 ( .A1(n4260), .A2(n6374), .ZN(n4235) );
  MUX2_X1 U5186 ( .A(n3609), .B(n5373), .S(EBX_REG_25__SCAN_IN), .Z(n4237) );
  NOR2_X1 U5187 ( .A1(n4304), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4236)
         );
  NOR2_X1 U5188 ( .A1(n4237), .A2(n4236), .ZN(n5414) );
  OR2_X1 U5189 ( .A1(n4300), .A2(EBX_REG_24__SCAN_IN), .ZN(n4240) );
  OAI21_X1 U5190 ( .B1(n5373), .B2(n5529), .A(n3606), .ZN(n4238) );
  OAI21_X1 U5191 ( .B1(n3612), .B2(EBX_REG_24__SCAN_IN), .A(n4238), .ZN(n4239)
         );
  NAND2_X1 U5192 ( .A1(n4240), .A2(n4239), .ZN(n5415) );
  NAND2_X1 U5193 ( .A1(n5414), .A2(n5415), .ZN(n4241) );
  NOR2_X2 U5194 ( .A1(n5413), .A2(n4241), .ZN(n5417) );
  OR2_X1 U5195 ( .A1(n4300), .A2(EBX_REG_26__SCAN_IN), .ZN(n4244) );
  INV_X1 U5196 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U5197 ( .A1(n3606), .A2(n5635), .ZN(n4242) );
  OAI211_X1 U5198 ( .C1(n3612), .C2(EBX_REG_26__SCAN_IN), .A(n5317), .B(n4242), 
        .ZN(n4243) );
  NAND2_X1 U5199 ( .A1(n4244), .A2(n4243), .ZN(n5407) );
  NAND2_X1 U5200 ( .A1(n5317), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4245) );
  OAI211_X1 U5201 ( .C1(n3612), .C2(EBX_REG_27__SCAN_IN), .A(n3606), .B(n4245), 
        .ZN(n4246) );
  OAI21_X1 U5202 ( .B1(n3601), .B2(EBX_REG_27__SCAN_IN), .A(n4246), .ZN(n4314)
         );
  OR2_X1 U5203 ( .A1(n4300), .A2(EBX_REG_28__SCAN_IN), .ZN(n4249) );
  INV_X1 U5204 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5622) );
  OAI21_X1 U5205 ( .B1(n5373), .B2(n5622), .A(n3606), .ZN(n4247) );
  OAI21_X1 U5206 ( .B1(n3612), .B2(EBX_REG_28__SCAN_IN), .A(n4247), .ZN(n4248)
         );
  AND2_X1 U5207 ( .A1(n4249), .A2(n4248), .ZN(n5335) );
  INV_X1 U5208 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5606) );
  INV_X1 U5209 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U5210 ( .A1(n2973), .A2(n5606), .B1(n4422), .B2(n4250), .ZN(n5318)
         );
  INV_X1 U5211 ( .A(n4301), .ZN(n4251) );
  NAND2_X1 U5212 ( .A1(n4251), .A2(n5317), .ZN(n4302) );
  NAND2_X1 U5213 ( .A1(n4304), .A2(EBX_REG_30__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U5214 ( .A1(n3612), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4252) );
  NAND2_X1 U5215 ( .A1(n4253), .A2(n4252), .ZN(n4303) );
  OAI211_X1 U5216 ( .C1(n4301), .C2(n3000), .A(n4302), .B(n4303), .ZN(n4257)
         );
  INV_X1 U5217 ( .A(n4303), .ZN(n4254) );
  OAI21_X1 U5218 ( .B1(n5323), .B2(n5317), .A(n4254), .ZN(n4255) );
  OR2_X1 U5219 ( .A1(n4301), .A2(n4255), .ZN(n4256) );
  NAND2_X1 U5220 ( .A1(n4257), .A2(n4256), .ZN(n5598) );
  AND2_X1 U5221 ( .A1(n5087), .A2(EBX_REG_31__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U5222 ( .A1(n6485), .A2(n5829), .ZN(n4268) );
  INV_X1 U5223 ( .A(n4268), .ZN(n4258) );
  NOR2_X1 U5224 ( .A1(n3612), .A2(n4258), .ZN(n4259) );
  AND2_X1 U5225 ( .A1(n4260), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4261) );
  AOI22_X1 U5226 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5927), .B1(n5928), 
        .B2(n4262), .ZN(n4267) );
  INV_X1 U5227 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U5228 ( .A1(n4268), .A2(n5398), .ZN(n4264) );
  OR2_X1 U5229 ( .A1(n6398), .A2(n4268), .ZN(n6369) );
  AND2_X1 U5230 ( .A1(n4351), .A2(n6369), .ZN(n5304) );
  INV_X1 U5231 ( .A(n5304), .ZN(n4263) );
  OAI21_X1 U5232 ( .B1(n4269), .B2(n4264), .A(n4263), .ZN(n4265) );
  NAND2_X1 U5233 ( .A1(n5943), .A2(EBX_REG_30__SCAN_IN), .ZN(n4266) );
  OAI211_X1 U5234 ( .C1(n5598), .C2(n5910), .A(n4267), .B(n4266), .ZN(n4289)
         );
  INV_X1 U5235 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6431) );
  INV_X1 U5236 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6427) );
  INV_X1 U5237 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6425) );
  NAND3_X1 U5238 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U5239 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5869) );
  NOR3_X1 U5240 ( .A1(n6425), .A2(n5201), .A3(n5869), .ZN(n4276) );
  NAND3_X1 U5241 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_8__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .ZN(n4275) );
  NOR2_X1 U5242 ( .A1(n4269), .A2(n4268), .ZN(n4271) );
  AND2_X1 U5243 ( .A1(n4271), .A2(n4270), .ZN(n4272) );
  INV_X1 U5244 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6414) );
  NAND3_X1 U5245 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n5930) );
  NOR2_X1 U5246 ( .A1(n6414), .A2(n5930), .ZN(n4274) );
  NAND2_X1 U5247 ( .A1(n4276), .A2(n5886), .ZN(n5247) );
  NOR2_X1 U5248 ( .A1(n6427), .A2(n5247), .ZN(n5388) );
  NAND2_X1 U5249 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5388), .ZN(n5857) );
  NAND4_X1 U5250 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5371), .ZN(n5742) );
  NAND3_X1 U5251 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4280) );
  NOR2_X1 U5252 ( .A1(n5742), .A2(n4280), .ZN(n5714) );
  AND3_X1 U5253 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4283) );
  NAND2_X1 U5254 ( .A1(n5714), .A2(n4283), .ZN(n5343) );
  NAND2_X1 U5255 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4273) );
  NOR3_X1 U5256 ( .A1(n5343), .A2(REIP_REG_29__SCAN_IN), .A3(n4273), .ZN(n5330) );
  INV_X1 U5257 ( .A(n4273), .ZN(n4285) );
  INV_X1 U5258 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6574) );
  INV_X1 U5259 ( .A(n5100), .ZN(n5936) );
  NAND2_X1 U5260 ( .A1(REIP_REG_5__SCAN_IN), .A2(n4274), .ZN(n5070) );
  NOR3_X1 U5261 ( .A1(n5936), .A2(n5070), .A3(n4275), .ZN(n5865) );
  NAND2_X1 U5262 ( .A1(n5865), .A2(n4276), .ZN(n5202) );
  NOR4_X1 U5263 ( .A1(n6574), .A2(n6431), .A3(n6427), .A4(n5202), .ZN(n4277)
         );
  AND2_X1 U5264 ( .A1(n5931), .A2(n5100), .ZN(n5863) );
  OR2_X1 U5265 ( .A1(n4277), .A2(n5863), .ZN(n5378) );
  NAND2_X1 U5266 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5370) );
  NOR2_X1 U5267 ( .A1(n5554), .A2(n5370), .ZN(n4278) );
  OR2_X1 U5268 ( .A1(n5863), .A2(n4278), .ZN(n4279) );
  NAND2_X1 U5269 ( .A1(n5378), .A2(n4279), .ZN(n5752) );
  INV_X1 U5270 ( .A(n4280), .ZN(n4281) );
  NOR2_X1 U5271 ( .A1(n5931), .A2(n4281), .ZN(n4282) );
  NOR2_X1 U5272 ( .A1(n5752), .A2(n4282), .ZN(n5731) );
  OR2_X1 U5273 ( .A1(n5863), .A2(n4283), .ZN(n4284) );
  AND2_X1 U5274 ( .A1(n5731), .A2(n4284), .ZN(n5715) );
  OAI21_X1 U5275 ( .B1(n4285), .B2(n5931), .A(n5715), .ZN(n5342) );
  NOR2_X1 U5276 ( .A1(n5330), .A2(n5342), .ZN(n5302) );
  INV_X1 U5277 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6452) );
  NOR2_X1 U5278 ( .A1(n5302), .A2(n6452), .ZN(n4288) );
  NAND2_X1 U5279 ( .A1(REIP_REG_29__SCAN_IN), .A2(n4285), .ZN(n4286) );
  NOR2_X1 U5280 ( .A1(n5343), .A2(n4286), .ZN(n5303) );
  INV_X1 U5281 ( .A(n5674), .ZN(n6080) );
  AND2_X1 U5282 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4295) );
  INV_X1 U5283 ( .A(n5616), .ZN(n5483) );
  NAND2_X1 U5284 ( .A1(n6126), .A2(n6116), .ZN(n6096) );
  INV_X1 U5285 ( .A(n4296), .ZN(n4291) );
  NAND2_X1 U5286 ( .A1(n6096), .A2(n4291), .ZN(n4292) );
  NAND2_X1 U5287 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U5288 ( .A1(n5674), .A2(n5633), .ZN(n4294) );
  NAND2_X1 U5289 ( .A1(n5645), .A2(n4294), .ZN(n5629) );
  AOI21_X1 U5290 ( .B1(n5483), .B2(n5674), .A(n5629), .ZN(n5607) );
  OAI21_X1 U5291 ( .B1(n6080), .B2(n4295), .A(n5607), .ZN(n5600) );
  NAND2_X1 U5292 ( .A1(n5643), .A2(n4296), .ZN(n5798) );
  OR2_X1 U5293 ( .A1(n5798), .A2(n5633), .ZN(n5626) );
  INV_X1 U5294 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4297) );
  NOR4_X1 U5295 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5595), 
        .A4(n4297), .ZN(n4298) );
  AOI211_X1 U5296 ( .C1(n5600), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n4299), .B(n4298), .ZN(n4307) );
  NOR2_X1 U5297 ( .A1(n4300), .A2(EBX_REG_29__SCAN_IN), .ZN(n5319) );
  AOI22_X1 U5298 ( .A1(n4301), .A2(n5317), .B1(n5319), .B2(n5323), .ZN(n5325)
         );
  OAI21_X1 U5299 ( .B1(n5325), .B2(n4303), .A(n4302), .ZN(n4306) );
  OAI22_X1 U5300 ( .A1(n4304), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n3612), .B2(EBX_REG_31__SCAN_IN), .ZN(n4305) );
  XNOR2_X1 U5301 ( .A(n4306), .B(n4305), .ZN(n5399) );
  BUF_X1 U5302 ( .A(n4310), .Z(n4311) );
  AOI21_X1 U5303 ( .B1(n4312), .B2(n4309), .A(n4311), .ZN(n5506) );
  INV_X1 U5304 ( .A(n5506), .ZN(n5470) );
  NOR2_X1 U5305 ( .A1(n5470), .A2(n5880), .ZN(n4321) );
  NOR2_X1 U5306 ( .A1(n5343), .A2(REIP_REG_27__SCAN_IN), .ZN(n4320) );
  INV_X1 U5307 ( .A(REIP_REG_27__SCAN_IN), .ZN(n4313) );
  NOR2_X1 U5308 ( .A1(n5715), .A2(n4313), .ZN(n4319) );
  NAND2_X1 U5309 ( .A1(n5409), .A2(n4314), .ZN(n4315) );
  NAND2_X1 U5310 ( .A1(n5334), .A2(n4315), .ZN(n5624) );
  AOI22_X1 U5311 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n5927), .B1(n5928), 
        .B2(n5502), .ZN(n4317) );
  NAND2_X1 U5312 ( .A1(n5943), .A2(EBX_REG_27__SCAN_IN), .ZN(n4316) );
  OAI211_X1 U5313 ( .C1(n5624), .C2(n5910), .A(n4317), .B(n4316), .ZN(n4318)
         );
  OR4_X1 U5314 ( .A1(n4321), .A2(n4320), .A3(n4319), .A4(n4318), .ZN(U2800) );
  AND2_X1 U5315 ( .A1(n6284), .A2(n6374), .ZN(n4339) );
  NOR2_X1 U5316 ( .A1(n4339), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4323) );
  OAI21_X1 U5317 ( .B1(n5082), .B2(n4422), .A(n6483), .ZN(n4322) );
  OAI21_X1 U5318 ( .B1(n4323), .B2(n6483), .A(n4322), .ZN(U3474) );
  INV_X1 U5319 ( .A(n4324), .ZN(n4325) );
  OAI22_X1 U5320 ( .A1(n4404), .A2(n5082), .B1(n4326), .B2(n4325), .ZN(n5824)
         );
  NOR3_X1 U5321 ( .A1(n4422), .A2(n5082), .A3(n4327), .ZN(n4328) );
  NOR2_X1 U5322 ( .A1(n4328), .A2(READY_N), .ZN(n6487) );
  NOR2_X1 U5323 ( .A1(n5824), .A2(n6487), .ZN(n6364) );
  NOR2_X1 U5324 ( .A1(n6364), .A2(n6384), .ZN(n5831) );
  INV_X1 U5325 ( .A(MORE_REG_SCAN_IN), .ZN(n4338) );
  NAND2_X1 U5326 ( .A1(n6360), .A2(n4329), .ZN(n4330) );
  NOR2_X1 U5327 ( .A1(n4330), .A2(n4403), .ZN(n4331) );
  OR2_X1 U5328 ( .A1(n4404), .A2(n4331), .ZN(n4334) );
  NAND2_X1 U5329 ( .A1(n4404), .A2(n4332), .ZN(n4333) );
  OAI211_X1 U5330 ( .C1(n4336), .C2(n4335), .A(n4334), .B(n4333), .ZN(n6361)
         );
  NAND2_X1 U5331 ( .A1(n5831), .A2(n6361), .ZN(n4337) );
  OAI21_X1 U5332 ( .B1(n5831), .B2(n4338), .A(n4337), .ZN(U3471) );
  INV_X1 U5333 ( .A(n4349), .ZN(n4350) );
  AOI211_X1 U5334 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4340), .A(n4339), .B(
        n4350), .ZN(n4341) );
  INV_X1 U5335 ( .A(n4341), .ZN(U2788) );
  XOR2_X1 U5336 ( .A(n4342), .B(n2991), .Z(n5093) );
  INV_X1 U5337 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4343) );
  AOI21_X1 U5338 ( .B1(n4344), .B2(n5574), .A(n4343), .ZN(n4345) );
  INV_X1 U5339 ( .A(n4345), .ZN(n4348) );
  XOR2_X1 U5340 ( .A(n4346), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n4376) );
  INV_X1 U5341 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6478) );
  NOR2_X1 U5342 ( .A1(n6123), .A2(n6478), .ZN(n4378) );
  AOI21_X1 U5343 ( .B1(n4376), .B2(n6035), .A(n4378), .ZN(n4347) );
  OAI211_X1 U5344 ( .C1(n5093), .C2(n5579), .A(n4348), .B(n4347), .ZN(U2986)
         );
  NOR2_X1 U5345 ( .A1(n4349), .A2(n3224), .ZN(n4443) );
  INV_X2 U5346 ( .A(n4443), .ZN(n4484) );
  INV_X1 U5347 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6636) );
  OR3_X1 U5348 ( .A1(n4349), .A2(n3222), .A3(READY_N), .ZN(n4497) );
  NAND2_X1 U5349 ( .A1(n4475), .A2(DATAI_5_), .ZN(n4482) );
  OAI21_X1 U5350 ( .B1(n4351), .B2(n6485), .A(n4350), .ZN(n4362) );
  NAND2_X1 U5351 ( .A1(n4362), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4352) );
  OAI211_X1 U5352 ( .C1(n4484), .C2(n6636), .A(n4482), .B(n4352), .ZN(U2929)
         );
  NAND2_X1 U5353 ( .A1(n4475), .A2(DATAI_4_), .ZN(n4479) );
  NAND2_X1 U5354 ( .A1(n4362), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4353) );
  OAI211_X1 U5355 ( .C1(n4484), .C2(n3961), .A(n4479), .B(n4353), .ZN(U2928)
         );
  INV_X1 U5356 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4678) );
  NAND2_X1 U5357 ( .A1(n4475), .A2(DATAI_9_), .ZN(n4457) );
  NAND2_X1 U5358 ( .A1(n4362), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4354) );
  OAI211_X1 U5359 ( .C1(n4484), .C2(n4678), .A(n4457), .B(n4354), .ZN(U2933)
         );
  INV_X1 U5360 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U5361 ( .A1(n4475), .A2(DATAI_3_), .ZN(n4467) );
  NAND2_X1 U5362 ( .A1(n4362), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4355) );
  OAI211_X1 U5363 ( .C1(n4484), .C2(n4673), .A(n4467), .B(n4355), .ZN(U2927)
         );
  INV_X1 U5364 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4489) );
  NAND2_X1 U5365 ( .A1(n4475), .A2(DATAI_8_), .ZN(n4459) );
  NAND2_X1 U5366 ( .A1(n4362), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4356) );
  OAI211_X1 U5367 ( .C1(n4484), .C2(n4489), .A(n4459), .B(n4356), .ZN(U2932)
         );
  INV_X1 U5368 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4487) );
  NAND2_X1 U5369 ( .A1(n4475), .A2(DATAI_7_), .ZN(n4472) );
  NAND2_X1 U5370 ( .A1(n4362), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4357) );
  OAI211_X1 U5371 ( .C1(n4484), .C2(n4487), .A(n4472), .B(n4357), .ZN(U2931)
         );
  INV_X1 U5372 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U5373 ( .A1(n4475), .A2(DATAI_12_), .ZN(n4451) );
  NAND2_X1 U5374 ( .A1(n4362), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4358) );
  OAI211_X1 U5375 ( .C1(n4484), .C2(n6583), .A(n4451), .B(n4358), .ZN(U2936)
         );
  INV_X1 U5376 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4447) );
  NAND2_X1 U5377 ( .A1(n4475), .A2(DATAI_11_), .ZN(n4453) );
  NAND2_X1 U5378 ( .A1(n4362), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4359) );
  OAI211_X1 U5379 ( .C1(n4484), .C2(n4447), .A(n4453), .B(n4359), .ZN(U2935)
         );
  NAND2_X1 U5380 ( .A1(n4475), .A2(DATAI_10_), .ZN(n4455) );
  NAND2_X1 U5381 ( .A1(n4362), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4360) );
  OAI211_X1 U5382 ( .C1(n4484), .C2(n4113), .A(n4455), .B(n4360), .ZN(U2934)
         );
  INV_X1 U5383 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U5384 ( .A1(n4475), .A2(DATAI_1_), .ZN(n4449) );
  NAND2_X1 U5385 ( .A1(n4362), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4361) );
  OAI211_X1 U5386 ( .C1(n4484), .C2(n4669), .A(n4449), .B(n4361), .ZN(U2925)
         );
  INV_X1 U5387 ( .A(DATAI_15_), .ZN(n4364) );
  INV_X1 U5388 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4363) );
  INV_X1 U5389 ( .A(n4362), .ZN(n4440) );
  INV_X1 U5390 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5976) );
  OAI222_X1 U5391 ( .A1(n4364), .A2(n4497), .B1(n4363), .B2(n4440), .C1(n4484), 
        .C2(n5976), .ZN(U2954) );
  INV_X1 U5392 ( .A(n4365), .ZN(n4367) );
  NAND2_X1 U5393 ( .A1(n2973), .A2(n6117), .ZN(n4366) );
  NAND2_X1 U5394 ( .A1(n4367), .A2(n4366), .ZN(n5084) );
  OR2_X1 U5395 ( .A1(n4404), .A2(n4520), .ZN(n4402) );
  NAND4_X1 U5396 ( .A1(n4370), .A2(n4369), .A3(n5459), .A4(n4368), .ZN(n4372)
         );
  OR2_X1 U5397 ( .A1(n4372), .A2(n4371), .ZN(n4493) );
  INV_X1 U5398 ( .A(n4493), .ZN(n4373) );
  NAND2_X1 U5399 ( .A1(n4373), .A2(n4422), .ZN(n4374) );
  NAND2_X1 U5400 ( .A1(n4402), .A2(n4374), .ZN(n4375) );
  NAND2_X1 U5401 ( .A1(n5959), .A2(n5459), .ZN(n5455) );
  NAND2_X1 U5402 ( .A1(n5959), .A2(n3232), .ZN(n5441) );
  OAI222_X1 U5403 ( .A1(n5084), .A2(n5455), .B1(n5088), .B2(n5959), .C1(n5441), 
        .C2(n5093), .ZN(U2859) );
  INV_X1 U5404 ( .A(n4376), .ZN(n4384) );
  INV_X1 U5405 ( .A(n5084), .ZN(n4379) );
  AOI211_X1 U5406 ( .C1(n6121), .C2(n4379), .A(n4378), .B(n4377), .ZN(n4383)
         );
  OAI21_X1 U5407 ( .B1(n4381), .B2(n4380), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4382) );
  OAI211_X1 U5408 ( .C1(n4384), .C2(n5805), .A(n4383), .B(n4382), .ZN(U3018)
         );
  XNOR2_X1 U5409 ( .A(n4386), .B(n4385), .ZN(n4431) );
  OAI21_X1 U5410 ( .B1(n4389), .B2(n4388), .A(n4387), .ZN(n5104) );
  INV_X1 U5411 ( .A(n5104), .ZN(n4390) );
  NAND2_X1 U5412 ( .A1(n4390), .A2(n2963), .ZN(n4393) );
  NOR2_X1 U5413 ( .A1(n6123), .A2(n6573), .ZN(n4427) );
  AND2_X1 U5414 ( .A1(n6030), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4391)
         );
  AOI211_X1 U5415 ( .C1(n6007), .C2(n5097), .A(n4427), .B(n4391), .ZN(n4392)
         );
  OAI211_X1 U5416 ( .C1(n4431), .C2(n6011), .A(n4393), .B(n4392), .ZN(U2985)
         );
  NAND2_X1 U5417 ( .A1(n4536), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6340) );
  INV_X1 U5418 ( .A(n5818), .ZN(n6469) );
  INV_X1 U5419 ( .A(n5287), .ZN(n6467) );
  NAND2_X1 U5420 ( .A1(n4536), .A2(n6485), .ZN(n4397) );
  INV_X1 U5421 ( .A(n4394), .ZN(n4396) );
  AOI22_X1 U5422 ( .A1(n4397), .A2(n4396), .B1(n6398), .B2(n4395), .ZN(n4398)
         );
  NAND2_X1 U5423 ( .A1(n4404), .A2(n4398), .ZN(n4399) );
  NAND4_X1 U5424 ( .A1(n4402), .A2(n4401), .A3(n4400), .A4(n4399), .ZN(n4409)
         );
  NAND2_X1 U5425 ( .A1(n4404), .A2(n4403), .ZN(n4408) );
  INV_X1 U5426 ( .A(n4405), .ZN(n4406) );
  OR2_X1 U5427 ( .A1(n4557), .A2(n4406), .ZN(n4407) );
  NAND2_X1 U5428 ( .A1(n4408), .A2(n4407), .ZN(n4496) );
  OR2_X1 U5429 ( .A1(n4409), .A2(n4496), .ZN(n6343) );
  INV_X1 U5430 ( .A(n6343), .ZN(n4558) );
  NAND2_X1 U5431 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4562) );
  OR2_X1 U5432 ( .A1(n6379), .A2(n4562), .ZN(n6462) );
  INV_X1 U5433 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5830) );
  OAI22_X1 U5434 ( .A1(n4558), .A2(n6384), .B1(n6462), .B2(n5830), .ZN(n5820)
         );
  NAND2_X1 U5435 ( .A1(n6379), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6463) );
  INV_X1 U5436 ( .A(n6463), .ZN(n4410) );
  NOR2_X1 U5437 ( .A1(n5820), .A2(n4410), .ZN(n6471) );
  INV_X1 U5438 ( .A(n6471), .ZN(n5822) );
  OAI21_X1 U5439 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6467), .A(n5822), 
        .ZN(n5273) );
  INV_X1 U5440 ( .A(n4411), .ZN(n4418) );
  NAND2_X1 U5441 ( .A1(n4413), .A2(n4412), .ZN(n4414) );
  NOR2_X1 U5442 ( .A1(n4415), .A2(n4414), .ZN(n4417) );
  NAND4_X1 U5443 ( .A1(n4418), .A2(n4417), .A3(n4557), .A4(n4416), .ZN(n4534)
         );
  INV_X1 U5444 ( .A(n4419), .ZN(n5275) );
  AOI22_X1 U5445 ( .A1(n6278), .A2(n4534), .B1(n5275), .B2(n3070), .ZN(n6341)
         );
  OAI22_X1 U5446 ( .A1(n6341), .A2(n6469), .B1(n6374), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4420) );
  OAI22_X1 U5447 ( .A1(n5273), .A2(n4420), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5822), .ZN(n4421) );
  OAI21_X1 U5448 ( .B1(n6340), .B2(n6469), .A(n4421), .ZN(U3461) );
  XNOR2_X1 U5449 ( .A(n5094), .B(n4422), .ZN(n4428) );
  INV_X1 U5450 ( .A(n5959), .ZN(n5451) );
  AOI22_X1 U5451 ( .A1(n5955), .A2(n4428), .B1(EBX_REG_1__SCAN_IN), .B2(n5451), 
        .ZN(n4423) );
  OAI21_X1 U5452 ( .B1(n5104), .B2(n5441), .A(n4423), .ZN(U2858) );
  INV_X1 U5453 ( .A(n4424), .ZN(n6077) );
  NAND2_X1 U5454 ( .A1(n6077), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4430)
         );
  AND3_X1 U5455 ( .A1(n5674), .A2(n4425), .A3(n6127), .ZN(n4426) );
  AOI211_X1 U5456 ( .C1(n6121), .C2(n4428), .A(n4427), .B(n4426), .ZN(n4429)
         );
  OAI211_X1 U5457 ( .C1(n4431), .C2(n5805), .A(n4430), .B(n4429), .ZN(U3017)
         );
  NAND3_X1 U5458 ( .A1(n4434), .A2(n4433), .A3(n4387), .ZN(n4435) );
  AND2_X1 U5459 ( .A1(n4432), .A2(n4435), .ZN(n6034) );
  INV_X1 U5460 ( .A(n6034), .ZN(n4505) );
  OR2_X1 U5461 ( .A1(n4437), .A2(n4436), .ZN(n4438) );
  AND2_X1 U5462 ( .A1(n4509), .A2(n4438), .ZN(n6120) );
  AOI22_X1 U5463 ( .A1(n5955), .A2(n6120), .B1(EBX_REG_2__SCAN_IN), .B2(n5451), 
        .ZN(n4439) );
  OAI21_X1 U5464 ( .B1(n4505), .B2(n5441), .A(n4439), .ZN(U2857) );
  AOI22_X1 U5465 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n4481), .B1(n4443), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n4441) );
  NAND2_X1 U5466 ( .A1(n4475), .A2(DATAI_6_), .ZN(n4462) );
  NAND2_X1 U5467 ( .A1(n4441), .A2(n4462), .ZN(U2930) );
  INV_X1 U5468 ( .A(n4442), .ZN(n4444) );
  AOI21_X1 U5469 ( .B1(n4536), .B2(n4444), .A(n4443), .ZN(n4445) );
  NOR2_X1 U5470 ( .A1(n4445), .A2(n6398), .ZN(n5974) );
  NAND2_X1 U5471 ( .A1(n5974), .A2(n4590), .ZN(n4682) );
  NOR2_X1 U5472 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4562), .ZN(n6001) );
  AOI22_X1 U5473 ( .A1(DATAO_REG_27__SCAN_IN), .A2(n5993), .B1(n6001), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n4446) );
  OAI21_X1 U5474 ( .B1(n4447), .B2(n4682), .A(n4446), .ZN(U2896) );
  INV_X1 U5475 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U5476 ( .A1(n4481), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4448) );
  OAI211_X1 U5477 ( .C1(n4484), .C2(n6542), .A(n4449), .B(n4448), .ZN(U2940)
         );
  INV_X1 U5478 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U5479 ( .A1(n4481), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4450) );
  OAI211_X1 U5480 ( .C1(n4484), .C2(n5982), .A(n4451), .B(n4450), .ZN(U2951)
         );
  INV_X1 U5481 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U5482 ( .A1(n4481), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4452) );
  OAI211_X1 U5483 ( .C1(n4484), .C2(n5984), .A(n4453), .B(n4452), .ZN(U2950)
         );
  INV_X1 U5484 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U5485 ( .A1(n4481), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4454) );
  OAI211_X1 U5486 ( .C1(n4484), .C2(n6579), .A(n4455), .B(n4454), .ZN(U2949)
         );
  INV_X1 U5487 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U5488 ( .A1(n4481), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4456) );
  OAI211_X1 U5489 ( .C1(n4484), .C2(n6526), .A(n4457), .B(n4456), .ZN(U2948)
         );
  INV_X1 U5490 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U5491 ( .A1(n4481), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4458) );
  OAI211_X1 U5492 ( .C1(n4484), .C2(n5988), .A(n4459), .B(n4458), .ZN(U2947)
         );
  INV_X1 U5493 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U5494 ( .A1(n4475), .A2(DATAI_14_), .ZN(n4465) );
  NAND2_X1 U5495 ( .A1(n4481), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4460) );
  OAI211_X1 U5496 ( .C1(n4484), .C2(n5978), .A(n4465), .B(n4460), .ZN(U2953)
         );
  NAND2_X1 U5497 ( .A1(n4481), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4461) );
  OAI211_X1 U5498 ( .C1(n4484), .C2(n4862), .A(n4462), .B(n4461), .ZN(U2945)
         );
  INV_X1 U5499 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U5500 ( .A1(n4475), .A2(DATAI_0_), .ZN(n4474) );
  NAND2_X1 U5501 ( .A1(n4481), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4463) );
  OAI211_X1 U5502 ( .C1(n4484), .C2(n6005), .A(n4474), .B(n4463), .ZN(U2939)
         );
  INV_X1 U5503 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U5504 ( .A1(n4481), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4464) );
  OAI211_X1 U5505 ( .C1(n4484), .C2(n6591), .A(n4465), .B(n4464), .ZN(U2938)
         );
  INV_X1 U5506 ( .A(EAX_REG_3__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U5507 ( .A1(n4481), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4466) );
  OAI211_X1 U5508 ( .C1(n4484), .C2(n5997), .A(n4467), .B(n4466), .ZN(U2942)
         );
  INV_X1 U5509 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U5510 ( .A1(n4475), .A2(DATAI_2_), .ZN(n4470) );
  NAND2_X1 U5511 ( .A1(n4481), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4468) );
  OAI211_X1 U5512 ( .C1(n4484), .C2(n5999), .A(n4470), .B(n4468), .ZN(U2941)
         );
  NAND2_X1 U5513 ( .A1(n4481), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4469) );
  OAI211_X1 U5514 ( .C1(n4484), .C2(n3911), .A(n4470), .B(n4469), .ZN(U2926)
         );
  NAND2_X1 U5515 ( .A1(n4481), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4471) );
  OAI211_X1 U5516 ( .C1(n4484), .C2(n4946), .A(n4472), .B(n4471), .ZN(U2946)
         );
  INV_X1 U5517 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4675) );
  NAND2_X1 U5518 ( .A1(n4481), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4473) );
  OAI211_X1 U5519 ( .C1(n4484), .C2(n4675), .A(n4474), .B(n4473), .ZN(U2924)
         );
  NAND2_X1 U5520 ( .A1(n4475), .A2(DATAI_13_), .ZN(n4478) );
  NAND2_X1 U5521 ( .A1(n4481), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4476) );
  OAI211_X1 U5522 ( .C1(n4484), .C2(n4184), .A(n4478), .B(n4476), .ZN(U2937)
         );
  INV_X1 U5523 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U5524 ( .A1(n4481), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4477) );
  OAI211_X1 U5525 ( .C1(n4484), .C2(n5980), .A(n4478), .B(n4477), .ZN(U2952)
         );
  INV_X1 U5526 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U5527 ( .A1(n4481), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4480) );
  OAI211_X1 U5528 ( .C1(n4484), .C2(n5995), .A(n4480), .B(n4479), .ZN(U2943)
         );
  INV_X1 U5529 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U5530 ( .A1(n4481), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4483) );
  OAI211_X1 U5531 ( .C1(n4484), .C2(n5992), .A(n4483), .B(n4482), .ZN(U2944)
         );
  AOI22_X1 U5532 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6001), .B1(n5993), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4485) );
  OAI21_X1 U5533 ( .B1(n6591), .B2(n4682), .A(n4485), .ZN(U2893) );
  AOI22_X1 U5534 ( .A1(n6486), .A2(UWORD_REG_7__SCAN_IN), .B1(n5993), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4486) );
  OAI21_X1 U5535 ( .B1(n4487), .B2(n4682), .A(n4486), .ZN(U2900) );
  AOI22_X1 U5536 ( .A1(n6001), .A2(UWORD_REG_8__SCAN_IN), .B1(n5993), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4488) );
  OAI21_X1 U5537 ( .B1(n4489), .B2(n4682), .A(n4488), .ZN(U2899) );
  AOI22_X1 U5538 ( .A1(n6001), .A2(UWORD_REG_12__SCAN_IN), .B1(n5993), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4490) );
  OAI21_X1 U5539 ( .B1(n6583), .B2(n4682), .A(n4490), .ZN(U2895) );
  AOI22_X1 U5540 ( .A1(n6001), .A2(UWORD_REG_10__SCAN_IN), .B1(n5993), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4491) );
  OAI21_X1 U5541 ( .B1(n4113), .B2(n4682), .A(n4491), .ZN(U2897) );
  NOR2_X1 U5542 ( .A1(n4493), .A2(n4492), .ZN(n4495) );
  OAI21_X1 U5543 ( .B1(n4496), .B2(n4495), .A(n4494), .ZN(n4498) );
  AND2_X1 U5544 ( .A1(n4499), .A2(n3232), .ZN(n4504) );
  INV_X1 U5545 ( .A(n4504), .ZN(n4501) );
  AND2_X1 U5546 ( .A1(n4501), .A2(n4500), .ZN(n4502) );
  INV_X1 U5547 ( .A(DATAI_2_), .ZN(n4608) );
  OAI222_X1 U5548 ( .A1(n4505), .A2(n5760), .B1(n4944), .B2(n4608), .C1(n5458), 
        .C2(n5999), .ZN(U2889) );
  INV_X1 U5549 ( .A(DATAI_1_), .ZN(n4599) );
  OAI222_X1 U5550 ( .A1(n5104), .A2(n5760), .B1(n4944), .B2(n4599), .C1(n5458), 
        .C2(n6542), .ZN(U2890) );
  AOI21_X1 U5551 ( .B1(n4507), .B2(n4432), .A(n3014), .ZN(n4517) );
  INV_X1 U5552 ( .A(n4517), .ZN(n5159) );
  NAND2_X1 U5553 ( .A1(n4509), .A2(n4508), .ZN(n4510) );
  AND2_X1 U5554 ( .A1(n5919), .A2(n4510), .ZN(n6109) );
  AOI22_X1 U5555 ( .A1(n5955), .A2(n6109), .B1(EBX_REG_3__SCAN_IN), .B2(n5451), 
        .ZN(n4511) );
  OAI21_X1 U5556 ( .B1(n5159), .B2(n5441), .A(n4511), .ZN(U2856) );
  OAI21_X1 U5557 ( .B1(n4512), .B2(n4514), .A(n4513), .ZN(n6110) );
  NAND2_X1 U5558 ( .A1(n6101), .A2(REIP_REG_3__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U5559 ( .A1(n6030), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4515)
         );
  OAI211_X1 U5560 ( .C1(n6039), .C2(n5147), .A(n6107), .B(n4515), .ZN(n4516)
         );
  AOI21_X1 U5561 ( .B1(n4517), .B2(n2963), .A(n4516), .ZN(n4518) );
  OAI21_X1 U5562 ( .B1(n6011), .B2(n6110), .A(n4518), .ZN(U2983) );
  INV_X1 U5563 ( .A(n4542), .ZN(n4524) );
  NAND2_X1 U5564 ( .A1(n4520), .A2(n4519), .ZN(n4548) );
  INV_X1 U5565 ( .A(n4521), .ZN(n5285) );
  MUX2_X1 U5566 ( .A(n4524), .B(n4548), .S(n5285), .Z(n4523) );
  AND2_X1 U5567 ( .A1(n4536), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4522)
         );
  NOR2_X1 U5568 ( .A1(n4523), .A2(n4522), .ZN(n4528) );
  MUX2_X1 U5569 ( .A(n4524), .B(n4548), .S(n4521), .Z(n4526) );
  NAND2_X1 U5570 ( .A1(n4536), .A2(n3075), .ZN(n5278) );
  INV_X1 U5571 ( .A(n5278), .ZN(n4525) );
  NOR2_X1 U5572 ( .A1(n4526), .A2(n4525), .ZN(n4527) );
  MUX2_X1 U5573 ( .A(n4528), .B(n4527), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4531) );
  INV_X1 U5574 ( .A(n4529), .ZN(n4625) );
  NAND2_X1 U5575 ( .A1(n4625), .A2(n4534), .ZN(n4530) );
  NAND2_X1 U5576 ( .A1(n4531), .A2(n4530), .ZN(n5290) );
  INV_X1 U5577 ( .A(n5290), .ZN(n4532) );
  MUX2_X1 U5578 ( .A(n5292), .B(n4532), .S(n6343), .Z(n6348) );
  NOR2_X1 U5579 ( .A1(n6348), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4552) );
  INV_X1 U5580 ( .A(n2969), .ZN(n6230) );
  INV_X1 U5581 ( .A(n4534), .ZN(n5279) );
  NOR2_X1 U5582 ( .A1(n4521), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4535)
         );
  XNOR2_X1 U5583 ( .A(n4535), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4547)
         );
  NOR2_X1 U5584 ( .A1(n5278), .A2(n4539), .ZN(n4546) );
  INV_X1 U5585 ( .A(n4536), .ZN(n4544) );
  AOI21_X1 U5586 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n4538), .A(n4537), 
        .ZN(n4543) );
  AOI21_X1 U5587 ( .B1(n4521), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4539), 
        .ZN(n4540) );
  NOR2_X1 U5588 ( .A1(n4541), .A2(n4540), .ZN(n6468) );
  OAI22_X1 U5589 ( .A1(n4544), .A2(n4543), .B1(n6468), .B2(n4542), .ZN(n4545)
         );
  AOI211_X1 U5590 ( .C1(n4548), .C2(n4547), .A(n4546), .B(n4545), .ZN(n4549)
         );
  OAI21_X1 U5591 ( .B1(n6230), .B2(n5279), .A(n4549), .ZN(n6466) );
  MUX2_X1 U5592 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6466), .S(n6343), 
        .Z(n6357) );
  NAND2_X1 U5593 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5830), .ZN(n4559) );
  INV_X1 U5594 ( .A(n4559), .ZN(n4550) );
  AOI22_X1 U5595 ( .A1(n4552), .A2(n6357), .B1(n4551), .B2(n4550), .ZN(n6366)
         );
  NOR2_X1 U5596 ( .A1(n6366), .A2(n4553), .ZN(n4563) );
  INV_X1 U5597 ( .A(n4555), .ZN(n4915) );
  NOR2_X1 U5598 ( .A1(n4554), .A2(n4915), .ZN(n4556) );
  XNOR2_X1 U5599 ( .A(n4556), .B(n6646), .ZN(n5921) );
  INV_X1 U5600 ( .A(n4557), .ZN(n5819) );
  AOI22_X1 U5601 ( .A1(n5921), .A2(n5819), .B1(n4558), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4560) );
  OAI22_X1 U5602 ( .A1(n4560), .A2(STATE2_REG_1__SCAN_IN), .B1(n4559), .B2(
        n6646), .ZN(n6359) );
  NOR3_X1 U5603 ( .A1(n4563), .A2(n6359), .A3(FLUSH_REG_SCAN_IN), .ZN(n4561)
         );
  OAI21_X1 U5604 ( .B1(n4561), .B2(n6462), .A(n4628), .ZN(n6134) );
  NOR3_X1 U5605 ( .A1(n4563), .A2(n4562), .A3(n6359), .ZN(n6376) );
  NAND2_X1 U5606 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6464), .ZN(n4658) );
  INV_X1 U5607 ( .A(n4658), .ZN(n4565) );
  OAI22_X1 U5608 ( .A1(n4564), .A2(n6235), .B1(n3703), .B2(n4565), .ZN(n4566)
         );
  OAI21_X1 U5609 ( .B1(n6376), .B2(n4566), .A(n6134), .ZN(n4567) );
  OAI21_X1 U5610 ( .B1(n6134), .B2(n4955), .A(n4567), .ZN(U3465) );
  INV_X1 U5611 ( .A(DATAI_0_), .ZN(n4591) );
  OAI222_X1 U5612 ( .A1(n5760), .A2(n5093), .B1(n5458), .B2(n6005), .C1(n4591), 
        .C2(n4944), .ZN(U2891) );
  INV_X1 U5613 ( .A(DATAI_3_), .ZN(n4604) );
  OAI222_X1 U5614 ( .A1(n5159), .A2(n5760), .B1(n4944), .B2(n4604), .C1(n5458), 
        .C2(n5997), .ZN(U2888) );
  OR2_X1 U5615 ( .A1(n4570), .A2(n4569), .ZN(n4571) );
  NAND2_X1 U5616 ( .A1(n4568), .A2(n4571), .ZN(n5912) );
  INV_X1 U5617 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4574) );
  INV_X1 U5618 ( .A(n4572), .ZN(n5900) );
  OAI21_X1 U5619 ( .B1(n2989), .B2(n4573), .A(n5900), .ZN(n6090) );
  OAI222_X1 U5620 ( .A1(n5912), .A2(n5441), .B1(n5959), .B2(n4574), .C1(n6090), 
        .C2(n5455), .ZN(U2854) );
  NAND2_X1 U5621 ( .A1(n3717), .A2(n4575), .ZN(n6277) );
  NAND2_X1 U5622 ( .A1(n4577), .A2(n4914), .ZN(n6189) );
  NAND2_X1 U5623 ( .A1(n2963), .A2(DATAI_28_), .ZN(n6258) );
  NAND3_X1 U5624 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6345), .ZN(n4804) );
  NOR2_X1 U5625 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4804), .ZN(n4620)
         );
  INV_X1 U5626 ( .A(n4620), .ZN(n4579) );
  AND2_X1 U5627 ( .A1(n4586), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4919) );
  INV_X1 U5628 ( .A(n4736), .ZN(n4578) );
  NOR2_X1 U5629 ( .A1(n4578), .A2(n4989), .ZN(n6231) );
  OAI21_X1 U5630 ( .B1(n6231), .B2(n6285), .A(n4737), .ZN(n6239) );
  AOI211_X1 U5631 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4579), .A(n4919), .B(
        n6239), .ZN(n4583) );
  INV_X1 U5632 ( .A(n4580), .ZN(n5280) );
  NAND2_X1 U5633 ( .A1(n4625), .A2(n5280), .ZN(n4799) );
  INV_X1 U5634 ( .A(n6192), .ZN(n4659) );
  OR2_X1 U5635 ( .A1(n4575), .A2(n4659), .ZN(n4630) );
  OAI21_X1 U5636 ( .B1(n6318), .B2(n5267), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4581) );
  OAI211_X1 U5637 ( .C1(n6230), .C2(n4799), .A(n4581), .B(n6284), .ZN(n4582)
         );
  NAND2_X1 U5638 ( .A1(n4583), .A2(n4582), .ZN(n4621) );
  NAND2_X1 U5639 ( .A1(n4621), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4589)
         );
  NAND2_X1 U5640 ( .A1(n4616), .A2(n4585), .ZN(n4993) );
  INV_X1 U5641 ( .A(n4993), .ZN(n6312) );
  INV_X1 U5642 ( .A(n5267), .ZN(n4617) );
  NAND2_X1 U5643 ( .A1(n2963), .A2(DATAI_20_), .ZN(n6316) );
  NOR2_X1 U5644 ( .A1(n4799), .A2(n6235), .ZN(n4923) );
  NOR2_X1 U5645 ( .A1(n4586), .A2(n6285), .ZN(n6240) );
  AOI22_X1 U5646 ( .A1(n4923), .A2(n2969), .B1(n6231), .B2(n6240), .ZN(n4618)
         );
  INV_X1 U5647 ( .A(DATAI_4_), .ZN(n4663) );
  NOR2_X1 U5648 ( .A1(n4663), .A2(n4628), .ZN(n6313) );
  INV_X1 U5649 ( .A(n6313), .ZN(n5032) );
  OAI22_X1 U5650 ( .A1(n4617), .A2(n6316), .B1(n4618), .B2(n5032), .ZN(n4587)
         );
  AOI21_X1 U5651 ( .B1(n6312), .B2(n4620), .A(n4587), .ZN(n4588) );
  OAI211_X1 U5652 ( .C1(n6339), .C2(n6258), .A(n4589), .B(n4588), .ZN(U3120)
         );
  NAND2_X1 U5653 ( .A1(n2963), .A2(DATAI_24_), .ZN(n6292) );
  NAND2_X1 U5654 ( .A1(n4621), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4594)
         );
  NAND2_X1 U5655 ( .A1(n4616), .A2(n4590), .ZN(n5008) );
  NAND2_X1 U5656 ( .A1(n2963), .A2(DATAI_16_), .ZN(n6178) );
  NOR2_X1 U5657 ( .A1(n4591), .A2(n4628), .ZN(n6289) );
  INV_X1 U5658 ( .A(n6289), .ZN(n5007) );
  OAI22_X1 U5659 ( .A1(n4617), .A2(n6178), .B1(n4618), .B2(n5007), .ZN(n4592)
         );
  AOI21_X1 U5660 ( .B1(n6275), .B2(n4620), .A(n4592), .ZN(n4593) );
  OAI211_X1 U5661 ( .C1(n6339), .C2(n6292), .A(n4594), .B(n4593), .ZN(U3116)
         );
  NAND2_X1 U5662 ( .A1(n2963), .A2(DATAI_29_), .ZN(n6324) );
  NAND2_X1 U5663 ( .A1(n4621), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4597)
         );
  NAND2_X1 U5664 ( .A1(n4616), .A2(n3207), .ZN(n5272) );
  INV_X1 U5665 ( .A(n5272), .ZN(n6319) );
  NAND2_X1 U5666 ( .A1(n2963), .A2(DATAI_21_), .ZN(n5260) );
  INV_X1 U5667 ( .A(DATAI_5_), .ZN(n4665) );
  NOR2_X1 U5668 ( .A1(n4665), .A2(n4628), .ZN(n6320) );
  INV_X1 U5669 ( .A(n6320), .ZN(n5258) );
  OAI22_X1 U5670 ( .A1(n4617), .A2(n5260), .B1(n4618), .B2(n5258), .ZN(n4595)
         );
  AOI21_X1 U5671 ( .B1(n6319), .B2(n4620), .A(n4595), .ZN(n4596) );
  OAI211_X1 U5672 ( .C1(n6339), .C2(n6324), .A(n4597), .B(n4596), .ZN(U3121)
         );
  NAND2_X1 U5673 ( .A1(n2963), .A2(DATAI_25_), .ZN(n6298) );
  NAND2_X1 U5674 ( .A1(n4621), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4602)
         );
  NAND2_X1 U5675 ( .A1(n4616), .A2(n3224), .ZN(n5003) );
  INV_X1 U5676 ( .A(n5003), .ZN(n6294) );
  NAND2_X1 U5677 ( .A1(n2963), .A2(DATAI_17_), .ZN(n6208) );
  NOR2_X1 U5678 ( .A1(n4599), .A2(n4628), .ZN(n6295) );
  INV_X1 U5679 ( .A(n6295), .ZN(n5002) );
  OAI22_X1 U5680 ( .A1(n4617), .A2(n6208), .B1(n4618), .B2(n5002), .ZN(n4600)
         );
  AOI21_X1 U5681 ( .B1(n6294), .B2(n4620), .A(n4600), .ZN(n4601) );
  OAI211_X1 U5682 ( .C1(n6339), .C2(n6298), .A(n4602), .B(n4601), .ZN(U3117)
         );
  NAND2_X1 U5683 ( .A1(n2963), .A2(DATAI_27_), .ZN(n6254) );
  NAND2_X1 U5684 ( .A1(n4621), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4607)
         );
  NAND2_X1 U5685 ( .A1(n4616), .A2(n4603), .ZN(n5024) );
  INV_X1 U5686 ( .A(n5024), .ZN(n6306) );
  NAND2_X1 U5687 ( .A1(n2963), .A2(DATAI_19_), .ZN(n6310) );
  NOR2_X1 U5688 ( .A1(n4604), .A2(n4628), .ZN(n6307) );
  INV_X1 U5689 ( .A(n6307), .ZN(n5021) );
  OAI22_X1 U5690 ( .A1(n4617), .A2(n6310), .B1(n4618), .B2(n5021), .ZN(n4605)
         );
  AOI21_X1 U5691 ( .B1(n6306), .B2(n4620), .A(n4605), .ZN(n4606) );
  OAI211_X1 U5692 ( .C1(n6339), .C2(n6254), .A(n4607), .B(n4606), .ZN(U3119)
         );
  NAND2_X1 U5693 ( .A1(n2963), .A2(DATAI_26_), .ZN(n6304) );
  NAND2_X1 U5694 ( .A1(n4621), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4611)
         );
  NAND2_X1 U5695 ( .A1(n4616), .A2(n3155), .ZN(n4998) );
  INV_X1 U5696 ( .A(n4998), .ZN(n6300) );
  NAND2_X1 U5697 ( .A1(n2963), .A2(DATAI_18_), .ZN(n6213) );
  NOR2_X1 U5698 ( .A1(n4608), .A2(n4628), .ZN(n6301) );
  INV_X1 U5699 ( .A(n6301), .ZN(n4997) );
  OAI22_X1 U5700 ( .A1(n4617), .A2(n6213), .B1(n4618), .B2(n4997), .ZN(n4609)
         );
  AOI21_X1 U5701 ( .B1(n6300), .B2(n4620), .A(n4609), .ZN(n4610) );
  OAI211_X1 U5702 ( .C1(n6339), .C2(n6304), .A(n4611), .B(n4610), .ZN(U3118)
         );
  NAND2_X1 U5703 ( .A1(n2963), .A2(DATAI_30_), .ZN(n6264) );
  NAND2_X1 U5704 ( .A1(n4616), .A2(n4612), .ZN(n5016) );
  INV_X1 U5705 ( .A(n5016), .ZN(n6326) );
  AND2_X1 U5706 ( .A1(DATAI_6_), .A2(n4737), .ZN(n6327) );
  INV_X1 U5707 ( .A(n6327), .ZN(n5042) );
  NAND2_X1 U5708 ( .A1(n2963), .A2(DATAI_22_), .ZN(n6330) );
  OAI22_X1 U5709 ( .A1(n4618), .A2(n5042), .B1(n4617), .B2(n6330), .ZN(n4613)
         );
  AOI21_X1 U5710 ( .B1(n6326), .B2(n4620), .A(n4613), .ZN(n4615) );
  NAND2_X1 U5711 ( .A1(n4621), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4614)
         );
  OAI211_X1 U5712 ( .C1(n6339), .C2(n6264), .A(n4615), .B(n4614), .ZN(U3122)
         );
  NAND2_X1 U5713 ( .A1(n2963), .A2(DATAI_31_), .ZN(n6498) );
  NAND2_X1 U5714 ( .A1(n4616), .A2(n3232), .ZN(n6506) );
  INV_X1 U5715 ( .A(n6506), .ZN(n6334) );
  AND2_X1 U5716 ( .A1(DATAI_7_), .A2(n4737), .ZN(n6502) );
  INV_X1 U5717 ( .A(n6502), .ZN(n5012) );
  NAND2_X1 U5718 ( .A1(n2963), .A2(DATAI_23_), .ZN(n6497) );
  OAI22_X1 U5719 ( .A1(n4618), .A2(n5012), .B1(n4617), .B2(n6497), .ZN(n4619)
         );
  AOI21_X1 U5720 ( .B1(n6334), .B2(n4620), .A(n4619), .ZN(n4623) );
  NAND2_X1 U5721 ( .A1(n4621), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4622)
         );
  OAI211_X1 U5722 ( .C1(n6339), .C2(n6498), .A(n4623), .B(n4622), .ZN(U3123)
         );
  INV_X1 U5723 ( .A(n4630), .ZN(n4624) );
  AOI21_X1 U5724 ( .B1(n4624), .B2(n4577), .A(n5579), .ZN(n4627) );
  NOR2_X1 U5725 ( .A1(n6235), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6237) );
  NAND2_X1 U5726 ( .A1(n4625), .A2(n4580), .ZN(n4772) );
  INV_X1 U5727 ( .A(n4772), .ZN(n6194) );
  AND2_X1 U5728 ( .A1(n2969), .A2(n6278), .ZN(n4801) );
  INV_X1 U5729 ( .A(n5257), .ZN(n4626) );
  AOI21_X1 U5730 ( .B1(n6194), .B2(n4801), .A(n4626), .ZN(n4631) );
  OAI21_X1 U5731 ( .B1(n4627), .B2(n6237), .A(n4631), .ZN(n4629) );
  AOI21_X1 U5732 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4955), .A(n4628), .ZN(
        n6281) );
  OAI211_X1 U5733 ( .C1(n6284), .C2(n4633), .A(n4629), .B(n6281), .ZN(n5251)
         );
  NAND2_X1 U5734 ( .A1(n5251), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4638)
         );
  INV_X1 U5735 ( .A(n6316), .ZN(n6255) );
  OR2_X1 U5736 ( .A1(n4630), .A2(n6189), .ZN(n4767) );
  NAND2_X1 U5737 ( .A1(n4577), .A2(n4564), .ZN(n4980) );
  INV_X1 U5738 ( .A(n4631), .ZN(n4632) );
  NAND2_X1 U5739 ( .A1(n4632), .A2(n6284), .ZN(n4635) );
  NAND2_X1 U5740 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4633), .ZN(n4634) );
  AND2_X1 U5741 ( .A1(n4635), .A2(n4634), .ZN(n5252) );
  OAI22_X1 U5742 ( .A1(n6496), .A2(n6258), .B1(n5252), .B2(n5032), .ZN(n4636)
         );
  AOI21_X1 U5743 ( .B1(n6255), .B2(n5254), .A(n4636), .ZN(n4637) );
  OAI211_X1 U5744 ( .C1(n4993), .C2(n5257), .A(n4638), .B(n4637), .ZN(U3144)
         );
  NAND2_X1 U5745 ( .A1(n5251), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4641)
         );
  INV_X1 U5746 ( .A(n5252), .ZN(n4643) );
  OAI22_X1 U5747 ( .A1(n6498), .A2(n6496), .B1(n4767), .B2(n6497), .ZN(n4639)
         );
  AOI21_X1 U5748 ( .B1(n6502), .B2(n4643), .A(n4639), .ZN(n4640) );
  OAI211_X1 U5749 ( .C1(n6506), .C2(n5257), .A(n4641), .B(n4640), .ZN(U3147)
         );
  NAND2_X1 U5750 ( .A1(n5251), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4645)
         );
  OAI22_X1 U5751 ( .A1(n6264), .A2(n6496), .B1(n4767), .B2(n6330), .ZN(n4642)
         );
  AOI21_X1 U5752 ( .B1(n6327), .B2(n4643), .A(n4642), .ZN(n4644) );
  OAI211_X1 U5753 ( .C1(n5016), .C2(n5257), .A(n4645), .B(n4644), .ZN(U3146)
         );
  NAND2_X1 U5754 ( .A1(n5251), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4648)
         );
  INV_X1 U5755 ( .A(n6208), .ZN(n6293) );
  OAI22_X1 U5756 ( .A1(n6496), .A2(n6298), .B1(n5252), .B2(n5002), .ZN(n4646)
         );
  AOI21_X1 U5757 ( .B1(n6293), .B2(n5254), .A(n4646), .ZN(n4647) );
  OAI211_X1 U5758 ( .C1(n5003), .C2(n5257), .A(n4648), .B(n4647), .ZN(U3141)
         );
  NAND2_X1 U5759 ( .A1(n5251), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4651)
         );
  INV_X1 U5760 ( .A(n6310), .ZN(n6251) );
  OAI22_X1 U5761 ( .A1(n6496), .A2(n6254), .B1(n5252), .B2(n5021), .ZN(n4649)
         );
  AOI21_X1 U5762 ( .B1(n6251), .B2(n5254), .A(n4649), .ZN(n4650) );
  OAI211_X1 U5763 ( .C1(n5024), .C2(n5257), .A(n4651), .B(n4650), .ZN(U3143)
         );
  NAND2_X1 U5764 ( .A1(n5251), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4654)
         );
  INV_X1 U5765 ( .A(n6178), .ZN(n6274) );
  OAI22_X1 U5766 ( .A1(n6496), .A2(n6292), .B1(n5252), .B2(n5007), .ZN(n4652)
         );
  AOI21_X1 U5767 ( .B1(n6274), .B2(n5254), .A(n4652), .ZN(n4653) );
  OAI211_X1 U5768 ( .C1(n5008), .C2(n5257), .A(n4654), .B(n4653), .ZN(U3140)
         );
  NAND2_X1 U5769 ( .A1(n5251), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4657)
         );
  INV_X1 U5770 ( .A(n6213), .ZN(n6299) );
  OAI22_X1 U5771 ( .A1(n6496), .A2(n6304), .B1(n5252), .B2(n4997), .ZN(n4655)
         );
  AOI21_X1 U5772 ( .B1(n6299), .B2(n5254), .A(n4655), .ZN(n4656) );
  OAI211_X1 U5773 ( .C1(n4998), .C2(n5257), .A(n4657), .B(n4656), .ZN(U3142)
         );
  NAND2_X1 U5774 ( .A1(n6134), .A2(n4658), .ZN(n5298) );
  INV_X1 U5775 ( .A(n6134), .ZN(n5294) );
  NOR2_X1 U5776 ( .A1(n5294), .A2(n6235), .ZN(n5296) );
  NAND2_X1 U5777 ( .A1(n4577), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6276) );
  NOR2_X1 U5778 ( .A1(n4575), .A2(n6276), .ZN(n6191) );
  MUX2_X1 U5779 ( .A(n3717), .B(n4659), .S(n6191), .Z(n4660) );
  AOI22_X1 U5780 ( .A1(n5296), .A2(n4660), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n5294), .ZN(n4661) );
  OAI21_X1 U5781 ( .B1(n6230), .B2(n5298), .A(n4661), .ZN(U3462) );
  XOR2_X1 U5782 ( .A(n4506), .B(n4662), .Z(n6026) );
  INV_X1 U5783 ( .A(n6026), .ZN(n4664) );
  OAI222_X1 U5784 ( .A1(n5760), .A2(n4664), .B1(n5458), .B2(n5995), .C1(n4663), 
        .C2(n4944), .ZN(U2887) );
  OAI222_X1 U5785 ( .A1(n5912), .A2(n5760), .B1(n4944), .B2(n4665), .C1(n5458), 
        .C2(n5992), .ZN(U2886) );
  OAI211_X1 U5786 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4577), .A(n5296), .B(
        n6276), .ZN(n4667) );
  NAND2_X1 U5787 ( .A1(n5294), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4666) );
  OAI211_X1 U5788 ( .C1(n5298), .C2(n5280), .A(n4667), .B(n4666), .ZN(U3464)
         );
  AOI22_X1 U5789 ( .A1(n6486), .A2(UWORD_REG_1__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4668) );
  OAI21_X1 U5790 ( .B1(n4669), .B2(n4682), .A(n4668), .ZN(U2906) );
  AOI22_X1 U5791 ( .A1(n6486), .A2(UWORD_REG_2__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4670) );
  OAI21_X1 U5792 ( .B1(n3911), .B2(n4682), .A(n4670), .ZN(U2905) );
  AOI22_X1 U5793 ( .A1(n6486), .A2(UWORD_REG_5__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4671) );
  OAI21_X1 U5794 ( .B1(n6636), .B2(n4682), .A(n4671), .ZN(U2902) );
  AOI22_X1 U5795 ( .A1(n6486), .A2(UWORD_REG_3__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4672) );
  OAI21_X1 U5796 ( .B1(n4673), .B2(n4682), .A(n4672), .ZN(U2904) );
  AOI22_X1 U5797 ( .A1(n6486), .A2(UWORD_REG_0__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4674) );
  OAI21_X1 U5798 ( .B1(n4675), .B2(n4682), .A(n4674), .ZN(U2907) );
  AOI22_X1 U5799 ( .A1(n6486), .A2(UWORD_REG_4__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4676) );
  OAI21_X1 U5800 ( .B1(n3961), .B2(n4682), .A(n4676), .ZN(U2903) );
  AOI22_X1 U5801 ( .A1(n6486), .A2(UWORD_REG_9__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4677) );
  OAI21_X1 U5802 ( .B1(n4678), .B2(n4682), .A(n4677), .ZN(U2898) );
  INV_X1 U5803 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U5804 ( .A1(n6486), .A2(UWORD_REG_6__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4679) );
  OAI21_X1 U5805 ( .B1(n4680), .B2(n4682), .A(n4679), .ZN(U2901) );
  AOI22_X1 U5806 ( .A1(n6001), .A2(UWORD_REG_13__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4681) );
  OAI21_X1 U5807 ( .B1(n4184), .B2(n4682), .A(n4681), .ZN(U2894) );
  OR2_X1 U5808 ( .A1(n4689), .A2(n5829), .ZN(n4683) );
  NAND2_X1 U5809 ( .A1(n5280), .A2(n4529), .ZN(n6229) );
  INV_X1 U5810 ( .A(n6229), .ZN(n4684) );
  NAND3_X1 U5811 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6351), .A3(n6345), .ZN(n6228) );
  NOR2_X1 U5812 ( .A1(n4955), .A2(n6228), .ZN(n4706) );
  AOI21_X1 U5813 ( .B1(n4801), .B2(n4684), .A(n4706), .ZN(n4688) );
  AOI22_X1 U5814 ( .A1(n4686), .A2(n4688), .B1(n6235), .B2(n6228), .ZN(n4685)
         );
  NAND2_X1 U5815 ( .A1(n6281), .A2(n4685), .ZN(n4705) );
  INV_X1 U5816 ( .A(n4686), .ZN(n4687) );
  OAI22_X1 U5817 ( .A1(n4688), .A2(n4687), .B1(n6285), .B2(n6228), .ZN(n4704)
         );
  AOI22_X1 U5818 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4705), .B1(n6327), 
        .B2(n4704), .ZN(n4691) );
  NOR2_X2 U5819 ( .A1(n4689), .A2(n4914), .ZN(n6267) );
  INV_X1 U5820 ( .A(n6264), .ZN(n6325) );
  AOI22_X1 U5821 ( .A1(n6267), .A2(n6325), .B1(n6326), .B2(n4706), .ZN(n4690)
         );
  OAI211_X1 U5822 ( .C1(n4876), .C2(n6330), .A(n4691), .B(n4690), .ZN(U3098)
         );
  AOI22_X1 U5823 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4705), .B1(n6307), 
        .B2(n4704), .ZN(n4693) );
  INV_X1 U5824 ( .A(n6254), .ZN(n6305) );
  AOI22_X1 U5825 ( .A1(n6267), .A2(n6305), .B1(n6306), .B2(n4706), .ZN(n4692)
         );
  OAI211_X1 U5826 ( .C1(n4876), .C2(n6310), .A(n4693), .B(n4692), .ZN(U3095)
         );
  AOI22_X1 U5827 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4705), .B1(n6295), 
        .B2(n4704), .ZN(n4695) );
  INV_X1 U5828 ( .A(n6298), .ZN(n6205) );
  AOI22_X1 U5829 ( .A1(n6267), .A2(n6205), .B1(n6294), .B2(n4706), .ZN(n4694)
         );
  OAI211_X1 U5830 ( .C1(n4876), .C2(n6208), .A(n4695), .B(n4694), .ZN(U3093)
         );
  AOI22_X1 U5831 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4705), .B1(n6320), 
        .B2(n4704), .ZN(n4697) );
  INV_X1 U5832 ( .A(n6324), .ZN(n5268) );
  AOI22_X1 U5833 ( .A1(n6267), .A2(n5268), .B1(n6319), .B2(n4706), .ZN(n4696)
         );
  OAI211_X1 U5834 ( .C1(n4876), .C2(n5260), .A(n4697), .B(n4696), .ZN(U3097)
         );
  AOI22_X1 U5835 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4705), .B1(n6289), 
        .B2(n4704), .ZN(n4699) );
  INV_X1 U5836 ( .A(n6292), .ZN(n6175) );
  AOI22_X1 U5837 ( .A1(n6267), .A2(n6175), .B1(n6275), .B2(n4706), .ZN(n4698)
         );
  OAI211_X1 U5838 ( .C1(n4876), .C2(n6178), .A(n4699), .B(n4698), .ZN(U3092)
         );
  AOI22_X1 U5839 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4705), .B1(n6313), 
        .B2(n4704), .ZN(n4701) );
  INV_X1 U5840 ( .A(n6258), .ZN(n6311) );
  AOI22_X1 U5841 ( .A1(n6267), .A2(n6311), .B1(n6312), .B2(n4706), .ZN(n4700)
         );
  OAI211_X1 U5842 ( .C1(n4876), .C2(n6316), .A(n4701), .B(n4700), .ZN(U3096)
         );
  AOI22_X1 U5843 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4705), .B1(n6301), 
        .B2(n4704), .ZN(n4703) );
  INV_X1 U5844 ( .A(n6304), .ZN(n6210) );
  AOI22_X1 U5845 ( .A1(n6267), .A2(n6210), .B1(n6300), .B2(n4706), .ZN(n4702)
         );
  OAI211_X1 U5846 ( .C1(n4876), .C2(n6213), .A(n4703), .B(n4702), .ZN(U3094)
         );
  AOI22_X1 U5847 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4705), .B1(n6502), 
        .B2(n4704), .ZN(n4708) );
  INV_X1 U5848 ( .A(n6498), .ZN(n6331) );
  AOI22_X1 U5849 ( .A1(n6267), .A2(n6331), .B1(n6334), .B2(n4706), .ZN(n4707)
         );
  OAI211_X1 U5850 ( .C1(n4876), .C2(n6497), .A(n4708), .B(n4707), .ZN(U3099)
         );
  NOR2_X1 U5851 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4709), .ZN(n4714)
         );
  INV_X1 U5852 ( .A(n4714), .ZN(n6505) );
  OAI21_X1 U5853 ( .B1(n4989), .B2(n6285), .A(n4737), .ZN(n4872) );
  NOR3_X1 U5854 ( .A1(n4872), .A2(n6358), .A3(n4919), .ZN(n4713) );
  NOR2_X2 U5855 ( .A1(n4797), .A2(n4564), .ZN(n5266) );
  INV_X1 U5856 ( .A(n6496), .ZN(n4710) );
  OAI21_X1 U5857 ( .B1(n5266), .B2(n4710), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4711) );
  NAND3_X1 U5858 ( .A1(n4772), .A2(n6284), .A3(n4711), .ZN(n4712) );
  OAI211_X1 U5859 ( .C1(n4714), .C2(n6464), .A(n4713), .B(n4712), .ZN(n6495)
         );
  NAND2_X1 U5860 ( .A1(n6495), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4718)
         );
  OR2_X1 U5861 ( .A1(n4772), .A2(n6235), .ZN(n4778) );
  NAND3_X1 U5862 ( .A1(n6240), .A2(n4989), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4715) );
  OAI21_X1 U5863 ( .B1(n4778), .B2(n6230), .A(n4715), .ZN(n6501) );
  INV_X1 U5864 ( .A(n5266), .ZN(n6499) );
  OAI22_X1 U5865 ( .A1(n6499), .A2(n6264), .B1(n6330), .B2(n6496), .ZN(n4716)
         );
  AOI21_X1 U5866 ( .B1(n6327), .B2(n6501), .A(n4716), .ZN(n4717) );
  OAI211_X1 U5867 ( .C1(n6505), .C2(n5016), .A(n4718), .B(n4717), .ZN(U3138)
         );
  NAND2_X1 U5868 ( .A1(n6495), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4721)
         );
  INV_X1 U5869 ( .A(n6501), .ZN(n5259) );
  OAI22_X1 U5870 ( .A1(n6496), .A2(n6213), .B1(n5259), .B2(n4997), .ZN(n4719)
         );
  AOI21_X1 U5871 ( .B1(n5266), .B2(n6210), .A(n4719), .ZN(n4720) );
  OAI211_X1 U5872 ( .C1(n6505), .C2(n4998), .A(n4721), .B(n4720), .ZN(U3134)
         );
  NAND2_X1 U5873 ( .A1(n6495), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4724)
         );
  OAI22_X1 U5874 ( .A1(n6496), .A2(n6178), .B1(n5259), .B2(n5007), .ZN(n4722)
         );
  AOI21_X1 U5875 ( .B1(n5266), .B2(n6175), .A(n4722), .ZN(n4723) );
  OAI211_X1 U5876 ( .C1(n6505), .C2(n5008), .A(n4724), .B(n4723), .ZN(U3132)
         );
  NAND2_X1 U5877 ( .A1(n6495), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4727)
         );
  OAI22_X1 U5878 ( .A1(n6496), .A2(n6316), .B1(n5259), .B2(n5032), .ZN(n4725)
         );
  AOI21_X1 U5879 ( .B1(n5266), .B2(n6311), .A(n4725), .ZN(n4726) );
  OAI211_X1 U5880 ( .C1(n6505), .C2(n4993), .A(n4727), .B(n4726), .ZN(U3136)
         );
  NAND2_X1 U5881 ( .A1(n6495), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4730)
         );
  OAI22_X1 U5882 ( .A1(n6496), .A2(n6208), .B1(n5259), .B2(n5002), .ZN(n4728)
         );
  AOI21_X1 U5883 ( .B1(n5266), .B2(n6205), .A(n4728), .ZN(n4729) );
  OAI211_X1 U5884 ( .C1(n6505), .C2(n5003), .A(n4730), .B(n4729), .ZN(U3133)
         );
  NAND2_X1 U5885 ( .A1(n6495), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4733)
         );
  OAI22_X1 U5886 ( .A1(n6496), .A2(n6310), .B1(n5259), .B2(n5021), .ZN(n4731)
         );
  AOI21_X1 U5887 ( .B1(n5266), .B2(n6305), .A(n4731), .ZN(n4732) );
  OAI211_X1 U5888 ( .C1(n6505), .C2(n5024), .A(n4733), .B(n4732), .ZN(U3135)
         );
  NAND2_X1 U5889 ( .A1(n4827), .A2(n4564), .ZN(n4847) );
  NOR2_X1 U5890 ( .A1(n5254), .A2(n6235), .ZN(n4735) );
  AOI21_X1 U5891 ( .B1(n4847), .B2(n4735), .A(n6237), .ZN(n4740) );
  NOR2_X1 U5892 ( .A1(n2969), .A2(n6229), .ZN(n4821) );
  NAND3_X1 U5893 ( .A1(n6358), .A2(n6351), .A3(n6345), .ZN(n4824) );
  NOR2_X1 U5894 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4824), .ZN(n4769)
         );
  INV_X1 U5895 ( .A(n4769), .ZN(n4738) );
  NOR2_X1 U5896 ( .A1(n4989), .A2(n4736), .ZN(n4922) );
  OAI21_X1 U5897 ( .B1(n4922), .B2(n6285), .A(n4737), .ZN(n4918) );
  AOI211_X1 U5898 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4738), .A(n6240), .B(
        n4918), .ZN(n4739) );
  OAI21_X1 U5899 ( .B1(n4740), .B2(n4821), .A(n4739), .ZN(n4765) );
  NAND2_X1 U5900 ( .A1(n4765), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4746) );
  INV_X1 U5901 ( .A(n4821), .ZN(n4741) );
  OR2_X1 U5902 ( .A1(n4741), .A2(n6235), .ZN(n4743) );
  NAND2_X1 U5903 ( .A1(n4922), .A2(n4919), .ZN(n4742) );
  AND2_X1 U5904 ( .A1(n4743), .A2(n4742), .ZN(n4766) );
  OAI22_X1 U5905 ( .A1(n4767), .A2(n6292), .B1(n4766), .B2(n5007), .ZN(n4744)
         );
  AOI21_X1 U5906 ( .B1(n6275), .B2(n4769), .A(n4744), .ZN(n4745) );
  OAI211_X1 U5907 ( .C1(n4847), .C2(n6178), .A(n4746), .B(n4745), .ZN(U3020)
         );
  NAND2_X1 U5908 ( .A1(n4765), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4749) );
  OAI22_X1 U5909 ( .A1(n4767), .A2(n6304), .B1(n4766), .B2(n4997), .ZN(n4747)
         );
  AOI21_X1 U5910 ( .B1(n6300), .B2(n4769), .A(n4747), .ZN(n4748) );
  OAI211_X1 U5911 ( .C1(n4847), .C2(n6213), .A(n4749), .B(n4748), .ZN(U3022)
         );
  NAND2_X1 U5912 ( .A1(n4765), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4752) );
  OAI22_X1 U5913 ( .A1(n4767), .A2(n6258), .B1(n4766), .B2(n5032), .ZN(n4750)
         );
  AOI21_X1 U5914 ( .B1(n6312), .B2(n4769), .A(n4750), .ZN(n4751) );
  OAI211_X1 U5915 ( .C1(n4847), .C2(n6316), .A(n4752), .B(n4751), .ZN(U3024)
         );
  NAND2_X1 U5916 ( .A1(n4765), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4755) );
  OAI22_X1 U5917 ( .A1(n4767), .A2(n6254), .B1(n4766), .B2(n5021), .ZN(n4753)
         );
  AOI21_X1 U5918 ( .B1(n6306), .B2(n4769), .A(n4753), .ZN(n4754) );
  OAI211_X1 U5919 ( .C1(n4847), .C2(n6310), .A(n4755), .B(n4754), .ZN(U3023)
         );
  NAND2_X1 U5920 ( .A1(n4765), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4758) );
  OAI22_X1 U5921 ( .A1(n5042), .A2(n4766), .B1(n6264), .B2(n4767), .ZN(n4756)
         );
  AOI21_X1 U5922 ( .B1(n6326), .B2(n4769), .A(n4756), .ZN(n4757) );
  OAI211_X1 U5923 ( .C1(n4847), .C2(n6330), .A(n4758), .B(n4757), .ZN(U3026)
         );
  NAND2_X1 U5924 ( .A1(n4765), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4761) );
  OAI22_X1 U5925 ( .A1(n5012), .A2(n4766), .B1(n6498), .B2(n4767), .ZN(n4759)
         );
  AOI21_X1 U5926 ( .B1(n6334), .B2(n4769), .A(n4759), .ZN(n4760) );
  OAI211_X1 U5927 ( .C1(n4847), .C2(n6497), .A(n4761), .B(n4760), .ZN(U3027)
         );
  NAND2_X1 U5928 ( .A1(n4765), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4764) );
  OAI22_X1 U5929 ( .A1(n4767), .A2(n6324), .B1(n4766), .B2(n5258), .ZN(n4762)
         );
  AOI21_X1 U5930 ( .B1(n6319), .B2(n4769), .A(n4762), .ZN(n4763) );
  OAI211_X1 U5931 ( .C1(n4847), .C2(n5260), .A(n4764), .B(n4763), .ZN(U3025)
         );
  NAND2_X1 U5932 ( .A1(n4765), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4771) );
  OAI22_X1 U5933 ( .A1(n4767), .A2(n6298), .B1(n4766), .B2(n5002), .ZN(n4768)
         );
  AOI21_X1 U5934 ( .B1(n6294), .B2(n4769), .A(n4768), .ZN(n4770) );
  OAI211_X1 U5935 ( .C1(n4847), .C2(n6208), .A(n4771), .B(n4770), .ZN(U3021)
         );
  OR2_X1 U5936 ( .A1(n4575), .A2(n6192), .ZN(n6190) );
  NOR3_X1 U5937 ( .A1(n6185), .A2(n6209), .A3(n6235), .ZN(n4773) );
  OAI21_X1 U5938 ( .B1(n4773), .B2(n6237), .A(n4772), .ZN(n4776) );
  INV_X1 U5939 ( .A(n6199), .ZN(n6200) );
  NOR2_X1 U5940 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6200), .ZN(n6184)
         );
  INV_X1 U5941 ( .A(n6184), .ZN(n4774) );
  AOI211_X1 U5942 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4774), .A(n4919), .B(
        n4872), .ZN(n4775) );
  NAND3_X1 U5943 ( .A1(n4776), .A2(n4775), .A3(n6358), .ZN(n6186) );
  INV_X1 U5944 ( .A(n6186), .ZN(n4796) );
  INV_X1 U5945 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4782) );
  NAND3_X1 U5946 ( .A1(n6240), .A2(n4989), .A3(n6358), .ZN(n4777) );
  OAI21_X1 U5947 ( .B1(n4778), .B2(n2969), .A(n4777), .ZN(n6183) );
  INV_X1 U5948 ( .A(n6183), .ZN(n4788) );
  INV_X1 U5949 ( .A(n6497), .ZN(n6268) );
  AOI22_X1 U5950 ( .A1(n6185), .A2(n6331), .B1(n6268), .B2(n6209), .ZN(n4779)
         );
  OAI21_X1 U5951 ( .B1(n5012), .B2(n4788), .A(n4779), .ZN(n4780) );
  AOI21_X1 U5952 ( .B1(n6334), .B2(n6184), .A(n4780), .ZN(n4781) );
  OAI21_X1 U5953 ( .B1(n4796), .B2(n4782), .A(n4781), .ZN(U3075) );
  INV_X1 U5954 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4786) );
  INV_X1 U5955 ( .A(n5260), .ZN(n6317) );
  AOI22_X1 U5956 ( .A1(n6209), .A2(n6317), .B1(n6320), .B2(n6183), .ZN(n4783)
         );
  OAI21_X1 U5957 ( .B1(n5038), .B2(n6324), .A(n4783), .ZN(n4784) );
  AOI21_X1 U5958 ( .B1(n6319), .B2(n6184), .A(n4784), .ZN(n4785) );
  OAI21_X1 U5959 ( .B1(n4796), .B2(n4786), .A(n4785), .ZN(U3073) );
  INV_X1 U5960 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4791) );
  INV_X1 U5961 ( .A(n6330), .ZN(n6261) );
  AOI22_X1 U5962 ( .A1(n6185), .A2(n6325), .B1(n6261), .B2(n6209), .ZN(n4787)
         );
  OAI21_X1 U5963 ( .B1(n5042), .B2(n4788), .A(n4787), .ZN(n4789) );
  AOI21_X1 U5964 ( .B1(n6326), .B2(n6184), .A(n4789), .ZN(n4790) );
  OAI21_X1 U5965 ( .B1(n4796), .B2(n4791), .A(n4790), .ZN(U3074) );
  INV_X1 U5966 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U5967 ( .A1(n6209), .A2(n6255), .B1(n6313), .B2(n6183), .ZN(n4792)
         );
  OAI21_X1 U5968 ( .B1(n5038), .B2(n6258), .A(n4792), .ZN(n4793) );
  AOI21_X1 U5969 ( .B1(n6312), .B2(n6184), .A(n4793), .ZN(n4794) );
  OAI21_X1 U5970 ( .B1(n4796), .B2(n4795), .A(n4794), .ZN(U3072) );
  NOR2_X1 U5971 ( .A1(n4955), .A2(n4804), .ZN(n4800) );
  INV_X1 U5972 ( .A(n4800), .ZN(n5271) );
  INV_X1 U5973 ( .A(n4797), .ZN(n4798) );
  AOI21_X1 U5974 ( .B1(n4798), .B2(STATEBS16_REG_SCAN_IN), .A(n6235), .ZN(
        n4803) );
  INV_X1 U5975 ( .A(n4799), .ZN(n4916) );
  AOI21_X1 U5976 ( .B1(n4916), .B2(n4801), .A(n4800), .ZN(n4806) );
  AOI22_X1 U5977 ( .A1(n4803), .A2(n4806), .B1(n6235), .B2(n4804), .ZN(n4802)
         );
  NAND2_X1 U5978 ( .A1(n6281), .A2(n4802), .ZN(n5265) );
  INV_X1 U5979 ( .A(n4803), .ZN(n4805) );
  OAI22_X1 U5980 ( .A1(n4806), .A2(n4805), .B1(n6285), .B2(n4804), .ZN(n5264)
         );
  AOI22_X1 U5981 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5265), .B1(n6502), 
        .B2(n5264), .ZN(n4808) );
  AOI22_X1 U5982 ( .A1(n6331), .A2(n5267), .B1(n5266), .B2(n6268), .ZN(n4807)
         );
  OAI211_X1 U5983 ( .C1(n6506), .C2(n5271), .A(n4808), .B(n4807), .ZN(U3131)
         );
  AOI22_X1 U5984 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5265), .B1(n6327), 
        .B2(n5264), .ZN(n4810) );
  AOI22_X1 U5985 ( .A1(n6325), .A2(n5267), .B1(n5266), .B2(n6261), .ZN(n4809)
         );
  OAI211_X1 U5986 ( .C1(n5016), .C2(n5271), .A(n4810), .B(n4809), .ZN(U3130)
         );
  AOI22_X1 U5987 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5265), .B1(n6295), 
        .B2(n5264), .ZN(n4812) );
  AOI22_X1 U5988 ( .A1(n6205), .A2(n5267), .B1(n5266), .B2(n6293), .ZN(n4811)
         );
  OAI211_X1 U5989 ( .C1(n5003), .C2(n5271), .A(n4812), .B(n4811), .ZN(U3125)
         );
  AOI22_X1 U5990 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5265), .B1(n6313), 
        .B2(n5264), .ZN(n4814) );
  AOI22_X1 U5991 ( .A1(n6311), .A2(n5267), .B1(n5266), .B2(n6255), .ZN(n4813)
         );
  OAI211_X1 U5992 ( .C1(n4993), .C2(n5271), .A(n4814), .B(n4813), .ZN(U3128)
         );
  AOI22_X1 U5993 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5265), .B1(n6307), 
        .B2(n5264), .ZN(n4816) );
  AOI22_X1 U5994 ( .A1(n6305), .A2(n5267), .B1(n5266), .B2(n6251), .ZN(n4815)
         );
  OAI211_X1 U5995 ( .C1(n5024), .C2(n5271), .A(n4816), .B(n4815), .ZN(U3127)
         );
  AOI22_X1 U5996 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5265), .B1(n6289), 
        .B2(n5264), .ZN(n4818) );
  AOI22_X1 U5997 ( .A1(n6175), .A2(n5267), .B1(n5266), .B2(n6274), .ZN(n4817)
         );
  OAI211_X1 U5998 ( .C1(n5008), .C2(n5271), .A(n4818), .B(n4817), .ZN(U3124)
         );
  AOI22_X1 U5999 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5265), .B1(n6301), 
        .B2(n5264), .ZN(n4820) );
  AOI22_X1 U6000 ( .A1(n6210), .A2(n5267), .B1(n5266), .B2(n6299), .ZN(n4819)
         );
  OAI211_X1 U6001 ( .C1(n4998), .C2(n5271), .A(n4820), .B(n4819), .ZN(U3126)
         );
  NOR2_X1 U6002 ( .A1(n4955), .A2(n4824), .ZN(n4844) );
  AOI21_X1 U6003 ( .B1(n4821), .B2(n6278), .A(n4844), .ZN(n4825) );
  AOI21_X1 U6004 ( .B1(n4827), .B2(STATEBS16_REG_SCAN_IN), .A(n6235), .ZN(
        n4823) );
  AOI22_X1 U6005 ( .A1(n4825), .A2(n4823), .B1(n6235), .B2(n4824), .ZN(n4822)
         );
  NAND2_X1 U6006 ( .A1(n6281), .A2(n4822), .ZN(n4843) );
  INV_X1 U6007 ( .A(n4823), .ZN(n4826) );
  OAI22_X1 U6008 ( .A1(n4826), .A2(n4825), .B1(n6285), .B2(n4824), .ZN(n4842)
         );
  AOI22_X1 U6009 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4843), .B1(n6320), 
        .B2(n4842), .ZN(n4829) );
  NAND2_X1 U6010 ( .A1(n4827), .A2(n4914), .ZN(n5028) );
  AOI22_X1 U6011 ( .A1(n4981), .A2(n6317), .B1(n6319), .B2(n4844), .ZN(n4828)
         );
  OAI211_X1 U6012 ( .C1(n6324), .C2(n4847), .A(n4829), .B(n4828), .ZN(U3033)
         );
  AOI22_X1 U6013 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4843), .B1(n6295), 
        .B2(n4842), .ZN(n4831) );
  AOI22_X1 U6014 ( .A1(n4981), .A2(n6293), .B1(n6294), .B2(n4844), .ZN(n4830)
         );
  OAI211_X1 U6015 ( .C1(n6298), .C2(n4847), .A(n4831), .B(n4830), .ZN(U3029)
         );
  AOI22_X1 U6016 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4843), .B1(n6289), 
        .B2(n4842), .ZN(n4833) );
  AOI22_X1 U6017 ( .A1(n4981), .A2(n6274), .B1(n6275), .B2(n4844), .ZN(n4832)
         );
  OAI211_X1 U6018 ( .C1(n6292), .C2(n4847), .A(n4833), .B(n4832), .ZN(U3028)
         );
  AOI22_X1 U6019 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4843), .B1(n6307), 
        .B2(n4842), .ZN(n4835) );
  AOI22_X1 U6020 ( .A1(n4981), .A2(n6251), .B1(n6306), .B2(n4844), .ZN(n4834)
         );
  OAI211_X1 U6021 ( .C1(n6254), .C2(n4847), .A(n4835), .B(n4834), .ZN(U3031)
         );
  AOI22_X1 U6022 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4843), .B1(n6313), 
        .B2(n4842), .ZN(n4837) );
  AOI22_X1 U6023 ( .A1(n4981), .A2(n6255), .B1(n6312), .B2(n4844), .ZN(n4836)
         );
  OAI211_X1 U6024 ( .C1(n6258), .C2(n4847), .A(n4837), .B(n4836), .ZN(U3032)
         );
  AOI22_X1 U6025 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4843), .B1(n6301), 
        .B2(n4842), .ZN(n4839) );
  AOI22_X1 U6026 ( .A1(n4981), .A2(n6299), .B1(n6300), .B2(n4844), .ZN(n4838)
         );
  OAI211_X1 U6027 ( .C1(n6304), .C2(n4847), .A(n4839), .B(n4838), .ZN(U3030)
         );
  AOI22_X1 U6028 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4843), .B1(n6327), 
        .B2(n4842), .ZN(n4841) );
  AOI22_X1 U6029 ( .A1(n4981), .A2(n6261), .B1(n6326), .B2(n4844), .ZN(n4840)
         );
  OAI211_X1 U6030 ( .C1(n6264), .C2(n4847), .A(n4841), .B(n4840), .ZN(U3034)
         );
  AOI22_X1 U6031 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4843), .B1(n6502), 
        .B2(n4842), .ZN(n4846) );
  AOI22_X1 U6032 ( .A1(n4981), .A2(n6268), .B1(n6334), .B2(n4844), .ZN(n4845)
         );
  OAI211_X1 U6033 ( .C1(n6498), .C2(n4847), .A(n4846), .B(n4845), .ZN(U3035)
         );
  OAI21_X1 U6034 ( .B1(n4850), .B2(n4849), .A(n4848), .ZN(n6087) );
  INV_X1 U6035 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4851) );
  OAI22_X1 U6036 ( .A1(n5574), .A2(n4852), .B1(n6123), .B2(n4851), .ZN(n4854)
         );
  NOR2_X1 U6037 ( .A1(n5912), .A2(n5579), .ZN(n4853) );
  AOI211_X1 U6038 ( .C1(n6007), .C2(n5913), .A(n4854), .B(n4853), .ZN(n4855)
         );
  OAI21_X1 U6039 ( .B1(n6011), .B2(n6087), .A(n4855), .ZN(U2981) );
  XOR2_X1 U6040 ( .A(n4856), .B(n4857), .Z(n5078) );
  INV_X1 U6041 ( .A(n5078), .ZN(n4943) );
  XOR2_X1 U6042 ( .A(n4910), .B(n5899), .Z(n6068) );
  AOI22_X1 U6043 ( .A1(n6068), .A2(n5955), .B1(EBX_REG_7__SCAN_IN), .B2(n5451), 
        .ZN(n4858) );
  OAI21_X1 U6044 ( .B1(n4943), .B2(n5441), .A(n4858), .ZN(U2852) );
  INV_X1 U6045 ( .A(DATAI_6_), .ZN(n4861) );
  XOR2_X1 U6046 ( .A(n4568), .B(n4859), .Z(n6017) );
  INV_X1 U6047 ( .A(n6017), .ZN(n4860) );
  OAI222_X1 U6048 ( .A1(n5458), .A2(n4862), .B1(n4861), .B2(n4944), .C1(n5760), 
        .C2(n4860), .ZN(U2885) );
  OAI21_X1 U6049 ( .B1(n4865), .B2(n4864), .A(n4863), .ZN(n6069) );
  INV_X1 U6050 ( .A(REIP_REG_7__SCAN_IN), .ZN(n4866) );
  NOR2_X1 U6051 ( .A1(n6123), .A2(n4866), .ZN(n6067) );
  AOI21_X1 U6052 ( .B1(n6030), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6067), 
        .ZN(n4867) );
  OAI21_X1 U6053 ( .B1(n5081), .B2(n6039), .A(n4867), .ZN(n4868) );
  AOI21_X1 U6054 ( .B1(n5078), .B2(n2963), .A(n4868), .ZN(n4869) );
  OAI21_X1 U6055 ( .B1(n6069), .B2(n6011), .A(n4869), .ZN(U2979) );
  AOI21_X1 U6056 ( .B1(n4876), .B2(n6323), .A(n5829), .ZN(n4870) );
  NOR2_X1 U6057 ( .A1(n4870), .A2(n6235), .ZN(n4874) );
  AND2_X1 U6058 ( .A1(n4580), .A2(n4529), .ZN(n4982) );
  AND2_X1 U6059 ( .A1(n4982), .A2(n2969), .ZN(n6279) );
  INV_X1 U6060 ( .A(n4919), .ZN(n6233) );
  NOR2_X1 U6061 ( .A1(n6233), .A2(n6358), .ZN(n4871) );
  AOI22_X1 U6062 ( .A1(n4874), .A2(n6279), .B1(n4989), .B2(n4871), .ZN(n4904)
         );
  NOR2_X1 U6063 ( .A1(n6240), .A2(n4872), .ZN(n4985) );
  INV_X1 U6064 ( .A(n6279), .ZN(n4873) );
  NAND2_X1 U6065 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4979), .ZN(n6286) );
  OR2_X1 U6066 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6286), .ZN(n4899)
         );
  AOI22_X1 U6067 ( .A1(n4874), .A2(n4873), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4899), .ZN(n4875) );
  OAI211_X1 U6068 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6285), .A(n4985), .B(n4875), .ZN(n4898) );
  NAND2_X1 U6069 ( .A1(n4898), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4879)
         );
  INV_X1 U6070 ( .A(n4876), .ZN(n4901) );
  OAI22_X1 U6071 ( .A1(n5008), .A2(n4899), .B1(n6323), .B2(n6178), .ZN(n4877)
         );
  AOI21_X1 U6072 ( .B1(n4901), .B2(n6175), .A(n4877), .ZN(n4878) );
  OAI211_X1 U6073 ( .C1(n4904), .C2(n5007), .A(n4879), .B(n4878), .ZN(U3100)
         );
  NAND2_X1 U6074 ( .A1(n4898), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4882)
         );
  OAI22_X1 U6075 ( .A1(n4899), .A2(n5003), .B1(n6323), .B2(n6208), .ZN(n4880)
         );
  AOI21_X1 U6076 ( .B1(n4901), .B2(n6205), .A(n4880), .ZN(n4881) );
  OAI211_X1 U6077 ( .C1(n4904), .C2(n5002), .A(n4882), .B(n4881), .ZN(U3101)
         );
  NAND2_X1 U6078 ( .A1(n4898), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4885)
         );
  OAI22_X1 U6079 ( .A1(n4899), .A2(n4993), .B1(n6323), .B2(n6316), .ZN(n4883)
         );
  AOI21_X1 U6080 ( .B1(n4901), .B2(n6311), .A(n4883), .ZN(n4884) );
  OAI211_X1 U6081 ( .C1(n4904), .C2(n5032), .A(n4885), .B(n4884), .ZN(U3104)
         );
  NAND2_X1 U6082 ( .A1(n4898), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4888)
         );
  OAI22_X1 U6083 ( .A1(n4899), .A2(n5272), .B1(n6323), .B2(n5260), .ZN(n4886)
         );
  AOI21_X1 U6084 ( .B1(n4901), .B2(n5268), .A(n4886), .ZN(n4887) );
  OAI211_X1 U6085 ( .C1(n4904), .C2(n5258), .A(n4888), .B(n4887), .ZN(U3105)
         );
  NAND2_X1 U6086 ( .A1(n4898), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4891)
         );
  OAI22_X1 U6087 ( .A1(n4899), .A2(n5024), .B1(n6323), .B2(n6310), .ZN(n4889)
         );
  AOI21_X1 U6088 ( .B1(n4901), .B2(n6305), .A(n4889), .ZN(n4890) );
  OAI211_X1 U6089 ( .C1(n4904), .C2(n5021), .A(n4891), .B(n4890), .ZN(U3103)
         );
  NAND2_X1 U6090 ( .A1(n4898), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4894)
         );
  OAI22_X1 U6091 ( .A1(n4899), .A2(n5016), .B1(n6323), .B2(n6330), .ZN(n4892)
         );
  AOI21_X1 U6092 ( .B1(n4901), .B2(n6325), .A(n4892), .ZN(n4893) );
  OAI211_X1 U6093 ( .C1(n4904), .C2(n5042), .A(n4894), .B(n4893), .ZN(U3106)
         );
  NAND2_X1 U6094 ( .A1(n4898), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4897)
         );
  OAI22_X1 U6095 ( .A1(n4899), .A2(n6506), .B1(n6323), .B2(n6497), .ZN(n4895)
         );
  AOI21_X1 U6096 ( .B1(n4901), .B2(n6331), .A(n4895), .ZN(n4896) );
  OAI211_X1 U6097 ( .C1(n4904), .C2(n5012), .A(n4897), .B(n4896), .ZN(U3107)
         );
  NAND2_X1 U6098 ( .A1(n4898), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4903)
         );
  OAI22_X1 U6099 ( .A1(n4899), .A2(n4998), .B1(n6323), .B2(n6213), .ZN(n4900)
         );
  AOI21_X1 U6100 ( .B1(n4901), .B2(n6210), .A(n4900), .ZN(n4902) );
  OAI211_X1 U6101 ( .C1(n4904), .C2(n4997), .A(n4903), .B(n4902), .ZN(U3102)
         );
  OAI21_X1 U6102 ( .B1(n4905), .B2(n4908), .A(n4907), .ZN(n5069) );
  OAI21_X1 U6103 ( .B1(n5899), .B2(n4910), .A(n4909), .ZN(n4911) );
  AND2_X1 U6104 ( .A1(n4911), .A2(n5049), .ZN(n6060) );
  AOI22_X1 U6105 ( .A1(n6060), .A2(n5955), .B1(EBX_REG_8__SCAN_IN), .B2(n5451), 
        .ZN(n4912) );
  OAI21_X1 U6106 ( .B1(n5069), .B2(n5441), .A(n4912), .ZN(U2851) );
  AOI22_X1 U6107 ( .A1(n5240), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n5970), .ZN(n4913) );
  OAI21_X1 U6108 ( .B1(n5069), .B2(n5760), .A(n4913), .ZN(U2883) );
  NAND3_X1 U6109 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6358), .A3(n6345), .ZN(n4960) );
  NOR2_X1 U6110 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4960), .ZN(n6169)
         );
  OAI21_X1 U6111 ( .B1(n6159), .B2(n6170), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4917) );
  NAND2_X1 U6112 ( .A1(n4916), .A2(n4915), .ZN(n4957) );
  AND2_X1 U6113 ( .A1(n4917), .A2(n4957), .ZN(n4920) );
  AOI211_X1 U6114 ( .C1(n6284), .C2(n4920), .A(n4919), .B(n4918), .ZN(n4921)
         );
  NAND2_X1 U6115 ( .A1(n6171), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4926) );
  INV_X1 U6116 ( .A(n6170), .ZN(n4939) );
  AOI22_X1 U6117 ( .A1(n4923), .A2(n6230), .B1(n6240), .B2(n4922), .ZN(n6165)
         );
  OAI22_X1 U6118 ( .A1(n4939), .A2(n6178), .B1(n6165), .B2(n5007), .ZN(n4924)
         );
  AOI21_X1 U6119 ( .B1(n6275), .B2(n6169), .A(n4924), .ZN(n4925) );
  OAI211_X1 U6120 ( .C1(n6292), .C2(n6174), .A(n4926), .B(n4925), .ZN(U3052)
         );
  NAND2_X1 U6121 ( .A1(n6171), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4929) );
  OAI22_X1 U6122 ( .A1(n4939), .A2(n6310), .B1(n6165), .B2(n5021), .ZN(n4927)
         );
  AOI21_X1 U6123 ( .B1(n6306), .B2(n6169), .A(n4927), .ZN(n4928) );
  OAI211_X1 U6124 ( .C1(n6174), .C2(n6254), .A(n4929), .B(n4928), .ZN(U3055)
         );
  NAND2_X1 U6125 ( .A1(n6171), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4932) );
  OAI22_X1 U6126 ( .A1(n4939), .A2(n6208), .B1(n6165), .B2(n5002), .ZN(n4930)
         );
  AOI21_X1 U6127 ( .B1(n6294), .B2(n6169), .A(n4930), .ZN(n4931) );
  OAI211_X1 U6128 ( .C1(n6174), .C2(n6298), .A(n4932), .B(n4931), .ZN(U3053)
         );
  NAND2_X1 U6129 ( .A1(n6171), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4935) );
  OAI22_X1 U6130 ( .A1(n4939), .A2(n5260), .B1(n6165), .B2(n5258), .ZN(n4933)
         );
  AOI21_X1 U6131 ( .B1(n6319), .B2(n6169), .A(n4933), .ZN(n4934) );
  OAI211_X1 U6132 ( .C1(n6174), .C2(n6324), .A(n4935), .B(n4934), .ZN(U3057)
         );
  NAND2_X1 U6133 ( .A1(n6171), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4938) );
  OAI22_X1 U6134 ( .A1(n6165), .A2(n5012), .B1(n4939), .B2(n6497), .ZN(n4936)
         );
  AOI21_X1 U6135 ( .B1(n6334), .B2(n6169), .A(n4936), .ZN(n4937) );
  OAI211_X1 U6136 ( .C1(n6174), .C2(n6498), .A(n4938), .B(n4937), .ZN(U3059)
         );
  NAND2_X1 U6137 ( .A1(n6171), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4942) );
  OAI22_X1 U6138 ( .A1(n4939), .A2(n6213), .B1(n6165), .B2(n4997), .ZN(n4940)
         );
  AOI21_X1 U6139 ( .B1(n6300), .B2(n6169), .A(n4940), .ZN(n4941) );
  OAI211_X1 U6140 ( .C1(n6174), .C2(n6304), .A(n4942), .B(n4941), .ZN(U3054)
         );
  INV_X1 U6141 ( .A(DATAI_7_), .ZN(n4945) );
  OAI222_X1 U6142 ( .A1(n5458), .A2(n4946), .B1(n4945), .B2(n4944), .C1(n5760), 
        .C2(n4943), .ZN(U2884) );
  INV_X1 U6143 ( .A(n5065), .ZN(n4950) );
  INV_X1 U6144 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4948) );
  AOI22_X1 U6145 ( .A1(EBX_REG_8__SCAN_IN), .A2(n5943), .B1(n5944), .B2(n6060), 
        .ZN(n4947) );
  NOR3_X2 U6146 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5936), .A3(n6235), .ZN(
        n5926) );
  INV_X1 U6147 ( .A(n5926), .ZN(n5887) );
  OAI211_X1 U6148 ( .C1(n5939), .C2(n4948), .A(n4947), .B(n5887), .ZN(n4949)
         );
  AOI21_X1 U6149 ( .B1(n5928), .B2(n4950), .A(n4949), .ZN(n4952) );
  INV_X1 U6150 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6635) );
  NOR2_X1 U6151 ( .A1(n6635), .A2(n5897), .ZN(n5077) );
  NOR2_X1 U6152 ( .A1(n5863), .A2(n5865), .ZN(n5134) );
  OAI221_X1 U6153 ( .B1(REIP_REG_8__SCAN_IN), .B2(REIP_REG_7__SCAN_IN), .C1(
        REIP_REG_8__SCAN_IN), .C2(n5077), .A(n5134), .ZN(n4951) );
  OAI211_X1 U6154 ( .C1(n5069), .C2(n5880), .A(n4952), .B(n4951), .ZN(U2819)
         );
  INV_X1 U6155 ( .A(n4953), .ZN(n4954) );
  AOI21_X1 U6156 ( .B1(n4954), .B2(STATEBS16_REG_SCAN_IN), .A(n6235), .ZN(
        n4962) );
  NOR2_X1 U6157 ( .A1(n4955), .A2(n4960), .ZN(n5040) );
  INV_X1 U6158 ( .A(n5040), .ZN(n4956) );
  OAI21_X1 U6159 ( .B1(n4957), .B2(n3703), .A(n4956), .ZN(n4959) );
  INV_X1 U6160 ( .A(n4960), .ZN(n4958) );
  AOI22_X1 U6161 ( .A1(n4962), .A2(n4959), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4958), .ZN(n5043) );
  INV_X1 U6162 ( .A(n4959), .ZN(n4961) );
  AOI22_X1 U6163 ( .A1(n4962), .A2(n4961), .B1(n4960), .B2(n6235), .ZN(n4963)
         );
  NAND2_X1 U6164 ( .A1(n6281), .A2(n4963), .ZN(n5036) );
  AOI22_X1 U6165 ( .A1(n6170), .A2(n6175), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n5036), .ZN(n4964) );
  OAI21_X1 U6166 ( .B1(n6178), .B2(n5038), .A(n4964), .ZN(n4965) );
  AOI21_X1 U6167 ( .B1(n6275), .B2(n5040), .A(n4965), .ZN(n4966) );
  OAI21_X1 U6168 ( .B1(n5043), .B2(n5007), .A(n4966), .ZN(U3060) );
  AOI22_X1 U6169 ( .A1(n6170), .A2(n6305), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n5036), .ZN(n4967) );
  OAI21_X1 U6170 ( .B1(n6310), .B2(n5038), .A(n4967), .ZN(n4968) );
  AOI21_X1 U6171 ( .B1(n6306), .B2(n5040), .A(n4968), .ZN(n4969) );
  OAI21_X1 U6172 ( .B1(n5043), .B2(n5021), .A(n4969), .ZN(U3063) );
  AOI22_X1 U6173 ( .A1(n6170), .A2(n6331), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n5036), .ZN(n4970) );
  OAI21_X1 U6174 ( .B1(n6497), .B2(n5038), .A(n4970), .ZN(n4971) );
  AOI21_X1 U6175 ( .B1(n6334), .B2(n5040), .A(n4971), .ZN(n4972) );
  OAI21_X1 U6176 ( .B1(n5043), .B2(n5012), .A(n4972), .ZN(U3067) );
  AOI22_X1 U6177 ( .A1(n6170), .A2(n6210), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n5036), .ZN(n4973) );
  OAI21_X1 U6178 ( .B1(n6213), .B2(n5038), .A(n4973), .ZN(n4974) );
  AOI21_X1 U6179 ( .B1(n6300), .B2(n5040), .A(n4974), .ZN(n4975) );
  OAI21_X1 U6180 ( .B1(n5043), .B2(n4997), .A(n4975), .ZN(U3062) );
  AOI22_X1 U6181 ( .A1(n6170), .A2(n6205), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n5036), .ZN(n4976) );
  OAI21_X1 U6182 ( .B1(n6208), .B2(n5038), .A(n4976), .ZN(n4977) );
  AOI21_X1 U6183 ( .B1(n6294), .B2(n5040), .A(n4977), .ZN(n4978) );
  OAI21_X1 U6184 ( .B1(n5043), .B2(n5002), .A(n4978), .ZN(U3061) );
  NAND2_X1 U6185 ( .A1(n4979), .A2(n6358), .ZN(n6141) );
  NOR2_X1 U6186 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6141), .ZN(n4987)
         );
  NOR2_X1 U6187 ( .A1(n4981), .A2(n6135), .ZN(n4984) );
  AND2_X1 U6188 ( .A1(n6230), .A2(n4982), .ZN(n6137) );
  INV_X1 U6189 ( .A(n6137), .ZN(n4983) );
  OAI21_X1 U6190 ( .B1(n4984), .B2(n6237), .A(n4983), .ZN(n4986) );
  OAI221_X1 U6191 ( .B1(n4987), .B2(n6464), .C1(n4987), .C2(n4986), .A(n4985), 
        .ZN(n5020) );
  NAND2_X1 U6192 ( .A1(n5020), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4992) );
  INV_X1 U6193 ( .A(n4987), .ZN(n5023) );
  NOR2_X1 U6194 ( .A1(n6233), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4988)
         );
  AOI22_X1 U6195 ( .A1(n6137), .A2(n6284), .B1(n4989), .B2(n4988), .ZN(n5022)
         );
  OAI22_X1 U6196 ( .A1(n5272), .A2(n5023), .B1(n5022), .B2(n5258), .ZN(n4990)
         );
  AOI21_X1 U6197 ( .B1(n6317), .B2(n6135), .A(n4990), .ZN(n4991) );
  OAI211_X1 U6198 ( .C1(n5028), .C2(n6324), .A(n4992), .B(n4991), .ZN(U3041)
         );
  NAND2_X1 U6199 ( .A1(n5020), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4996) );
  OAI22_X1 U6200 ( .A1(n4993), .A2(n5023), .B1(n5022), .B2(n5032), .ZN(n4994)
         );
  AOI21_X1 U6201 ( .B1(n6255), .B2(n6135), .A(n4994), .ZN(n4995) );
  OAI211_X1 U6202 ( .C1(n5028), .C2(n6258), .A(n4996), .B(n4995), .ZN(U3040)
         );
  NAND2_X1 U6203 ( .A1(n5020), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5001) );
  OAI22_X1 U6204 ( .A1(n4998), .A2(n5023), .B1(n5022), .B2(n4997), .ZN(n4999)
         );
  AOI21_X1 U6205 ( .B1(n6299), .B2(n6135), .A(n4999), .ZN(n5000) );
  OAI211_X1 U6206 ( .C1(n5028), .C2(n6304), .A(n5001), .B(n5000), .ZN(U3038)
         );
  NAND2_X1 U6207 ( .A1(n5020), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5006) );
  OAI22_X1 U6208 ( .A1(n5003), .A2(n5023), .B1(n5022), .B2(n5002), .ZN(n5004)
         );
  AOI21_X1 U6209 ( .B1(n6293), .B2(n6135), .A(n5004), .ZN(n5005) );
  OAI211_X1 U6210 ( .C1(n5028), .C2(n6298), .A(n5006), .B(n5005), .ZN(U3037)
         );
  NAND2_X1 U6211 ( .A1(n5020), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5011) );
  OAI22_X1 U6212 ( .A1(n5008), .A2(n5023), .B1(n5022), .B2(n5007), .ZN(n5009)
         );
  AOI21_X1 U6213 ( .B1(n6274), .B2(n6135), .A(n5009), .ZN(n5010) );
  OAI211_X1 U6214 ( .C1(n6292), .C2(n5028), .A(n5011), .B(n5010), .ZN(U3036)
         );
  NAND2_X1 U6215 ( .A1(n5020), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5015) );
  OAI22_X1 U6216 ( .A1(n5012), .A2(n5022), .B1(n6506), .B2(n5023), .ZN(n5013)
         );
  AOI21_X1 U6217 ( .B1(n6268), .B2(n6135), .A(n5013), .ZN(n5014) );
  OAI211_X1 U6218 ( .C1(n5028), .C2(n6498), .A(n5015), .B(n5014), .ZN(U3043)
         );
  NAND2_X1 U6219 ( .A1(n5020), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5019) );
  OAI22_X1 U6220 ( .A1(n5042), .A2(n5022), .B1(n5016), .B2(n5023), .ZN(n5017)
         );
  AOI21_X1 U6221 ( .B1(n6261), .B2(n6135), .A(n5017), .ZN(n5018) );
  OAI211_X1 U6222 ( .C1(n5028), .C2(n6264), .A(n5019), .B(n5018), .ZN(U3042)
         );
  NAND2_X1 U6223 ( .A1(n5020), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5027) );
  OAI22_X1 U6224 ( .A1(n5024), .A2(n5023), .B1(n5022), .B2(n5021), .ZN(n5025)
         );
  AOI21_X1 U6225 ( .B1(n6251), .B2(n6135), .A(n5025), .ZN(n5026) );
  OAI211_X1 U6226 ( .C1(n5028), .C2(n6254), .A(n5027), .B(n5026), .ZN(U3039)
         );
  AOI22_X1 U6227 ( .A1(n6170), .A2(n6311), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n5036), .ZN(n5029) );
  OAI21_X1 U6228 ( .B1(n6316), .B2(n5038), .A(n5029), .ZN(n5030) );
  AOI21_X1 U6229 ( .B1(n6312), .B2(n5040), .A(n5030), .ZN(n5031) );
  OAI21_X1 U6230 ( .B1(n5043), .B2(n5032), .A(n5031), .ZN(U3064) );
  AOI22_X1 U6231 ( .A1(n6170), .A2(n5268), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n5036), .ZN(n5033) );
  OAI21_X1 U6232 ( .B1(n5260), .B2(n5038), .A(n5033), .ZN(n5034) );
  AOI21_X1 U6233 ( .B1(n6319), .B2(n5040), .A(n5034), .ZN(n5035) );
  OAI21_X1 U6234 ( .B1(n5043), .B2(n5258), .A(n5035), .ZN(U3065) );
  AOI22_X1 U6235 ( .A1(n6170), .A2(n6325), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n5036), .ZN(n5037) );
  OAI21_X1 U6236 ( .B1(n6330), .B2(n5038), .A(n5037), .ZN(n5039) );
  AOI21_X1 U6237 ( .B1(n6326), .B2(n5040), .A(n5039), .ZN(n5041) );
  OAI21_X1 U6238 ( .B1(n5043), .B2(n5042), .A(n5041), .ZN(U3066) );
  INV_X1 U6239 ( .A(n5044), .ZN(n5045) );
  AOI21_X1 U6240 ( .B1(n5046), .B2(n4907), .A(n5045), .ZN(n5130) );
  INV_X1 U6241 ( .A(n5130), .ZN(n5056) );
  AOI22_X1 U6242 ( .A1(n5240), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5970), .ZN(n5047) );
  OAI21_X1 U6243 ( .B1(n5056), .B2(n5760), .A(n5047), .ZN(U2882) );
  AND2_X1 U6244 ( .A1(n5049), .A2(n5048), .ZN(n5050) );
  OR2_X1 U6245 ( .A1(n5050), .A2(n5110), .ZN(n5119) );
  AOI21_X1 U6246 ( .B1(n5927), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5926), 
        .ZN(n5052) );
  AOI22_X1 U6247 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5943), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5134), .ZN(n5051) );
  OAI211_X1 U6248 ( .C1(n5910), .C2(n5119), .A(n5052), .B(n5051), .ZN(n5053)
         );
  INV_X1 U6249 ( .A(n5886), .ZN(n5140) );
  NOR2_X1 U6250 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5140), .ZN(n5133) );
  AOI211_X1 U6251 ( .C1(n5054), .C2(n5928), .A(n5053), .B(n5133), .ZN(n5055)
         );
  OAI21_X1 U6252 ( .B1(n5880), .B2(n5056), .A(n5055), .ZN(U2818) );
  INV_X1 U6253 ( .A(n5441), .ZN(n5956) );
  INV_X1 U6254 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5057) );
  OAI22_X1 U6255 ( .A1(n5119), .A2(n5455), .B1(n5057), .B2(n5959), .ZN(n5058)
         );
  AOI21_X1 U6256 ( .B1(n5130), .B2(n5956), .A(n5058), .ZN(n5059) );
  INV_X1 U6257 ( .A(n5059), .ZN(U2850) );
  OAI21_X1 U6258 ( .B1(n5062), .B2(n5061), .A(n5060), .ZN(n5063) );
  INV_X1 U6259 ( .A(n5063), .ZN(n6063) );
  NAND2_X1 U6260 ( .A1(n6063), .A2(n6035), .ZN(n5068) );
  INV_X1 U6261 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5064) );
  NOR2_X1 U6262 ( .A1(n6123), .A2(n5064), .ZN(n6059) );
  NOR2_X1 U6263 ( .A1(n6039), .A2(n5065), .ZN(n5066) );
  AOI211_X1 U6264 ( .C1(n6030), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6059), 
        .B(n5066), .ZN(n5067) );
  OAI211_X1 U6265 ( .C1(n5579), .C2(n5069), .A(n5068), .B(n5067), .ZN(U2978)
         );
  INV_X1 U6266 ( .A(n5070), .ZN(n5071) );
  AND2_X1 U6267 ( .A1(n5100), .A2(n5071), .ZN(n5072) );
  OR2_X1 U6268 ( .A1(n5863), .A2(n5072), .ZN(n5918) );
  OAI21_X1 U6269 ( .B1(REIP_REG_6__SCAN_IN), .B2(n5897), .A(n5918), .ZN(n5076)
         );
  INV_X1 U6270 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5074) );
  AOI22_X1 U6271 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5943), .B1(n5944), .B2(n6068), 
        .ZN(n5073) );
  OAI211_X1 U6272 ( .C1(n5939), .C2(n5074), .A(n5073), .B(n5887), .ZN(n5075)
         );
  AOI221_X1 U6273 ( .B1(n5077), .B2(n4866), .C1(n5076), .C2(
        REIP_REG_7__SCAN_IN), .A(n5075), .ZN(n5080) );
  NAND2_X1 U6274 ( .A1(n5078), .A2(n5907), .ZN(n5079) );
  OAI211_X1 U6275 ( .C1(n5952), .C2(n5081), .A(n5080), .B(n5079), .ZN(U2820)
         );
  NAND2_X1 U6276 ( .A1(n5087), .A2(n5082), .ZN(n5083) );
  NAND2_X1 U6277 ( .A1(n5083), .A2(n5880), .ZN(n5950) );
  INV_X1 U6278 ( .A(n5950), .ZN(n5158) );
  NAND2_X1 U6279 ( .A1(n5939), .A2(n5952), .ZN(n5091) );
  OAI22_X1 U6280 ( .A1(n5863), .A2(n6478), .B1(n5910), .B2(n5084), .ZN(n5090)
         );
  INV_X1 U6281 ( .A(n5085), .ZN(n5086) );
  AND2_X1 U6282 ( .A1(n5087), .A2(n5086), .ZN(n5922) );
  INV_X1 U6283 ( .A(n5922), .ZN(n5941) );
  OAI22_X1 U6284 ( .A1(n5088), .A2(n5924), .B1(n5941), .B2(n3703), .ZN(n5089)
         );
  AOI211_X1 U6285 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n5091), .A(n5090), 
        .B(n5089), .ZN(n5092) );
  OAI21_X1 U6286 ( .B1(n5158), .B2(n5093), .A(n5092), .ZN(U2827) );
  INV_X1 U6287 ( .A(n5094), .ZN(n5096) );
  AOI22_X1 U6288 ( .A1(n5943), .A2(EBX_REG_1__SCAN_IN), .B1(n5922), .B2(n4580), 
        .ZN(n5095) );
  OAI21_X1 U6289 ( .B1(n5910), .B2(n5096), .A(n5095), .ZN(n5102) );
  NOR2_X1 U6290 ( .A1(n5931), .A2(REIP_REG_1__SCAN_IN), .ZN(n5937) );
  INV_X1 U6291 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6292 ( .A1(n5928), .A2(n5097), .ZN(n5099) );
  NAND2_X1 U6293 ( .A1(n5927), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5098)
         );
  OAI211_X1 U6294 ( .C1(n6573), .C2(n5100), .A(n5099), .B(n5098), .ZN(n5101)
         );
  NOR3_X1 U6295 ( .A1(n5102), .A2(n5937), .A3(n5101), .ZN(n5103) );
  OAI21_X1 U6296 ( .B1(n5158), .B2(n5104), .A(n5103), .ZN(U2826) );
  AND2_X1 U6297 ( .A1(n5044), .A2(n5105), .ZN(n5107) );
  OR2_X1 U6298 ( .A1(n5107), .A2(n5106), .ZN(n5166) );
  AOI22_X1 U6299 ( .A1(n5240), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5970), .ZN(n5108) );
  OAI21_X1 U6300 ( .B1(n5166), .B2(n5760), .A(n5108), .ZN(U2881) );
  OR2_X1 U6301 ( .A1(n5110), .A2(n5109), .ZN(n5111) );
  AND2_X1 U6302 ( .A1(n5169), .A2(n5111), .ZN(n6052) );
  AOI22_X1 U6303 ( .A1(n6052), .A2(n5955), .B1(EBX_REG_10__SCAN_IN), .B2(n5451), .ZN(n5112) );
  OAI21_X1 U6304 ( .B1(n5166), .B2(n5441), .A(n5112), .ZN(U2849) );
  NAND2_X1 U6305 ( .A1(n5114), .A2(n5113), .ZN(n5116) );
  XOR2_X1 U6306 ( .A(n5116), .B(n5115), .Z(n5132) );
  AOI22_X1 U6307 ( .A1(n6078), .A2(n5118), .B1(n5669), .B2(n5117), .ZN(n6075)
         );
  OAI21_X1 U6308 ( .B1(n6080), .B2(n6061), .A(n6075), .ZN(n6053) );
  NOR2_X1 U6309 ( .A1(n5119), .A2(n6089), .ZN(n5124) );
  INV_X1 U6310 ( .A(n6116), .ZN(n6097) );
  NOR2_X1 U6311 ( .A1(n5121), .A2(n5120), .ZN(n6079) );
  OAI211_X1 U6312 ( .C1(n6098), .C2(n6097), .A(n6079), .B(n6096), .ZN(n6084)
         );
  NOR2_X1 U6313 ( .A1(n5122), .A2(n6084), .ZN(n6070) );
  NAND2_X1 U6314 ( .A1(n6061), .A2(n6070), .ZN(n6058) );
  NAND2_X1 U6315 ( .A1(n6101), .A2(REIP_REG_9__SCAN_IN), .ZN(n5127) );
  OAI21_X1 U6316 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6058), .A(n5127), 
        .ZN(n5123) );
  AOI211_X1 U6317 ( .C1(n6053), .C2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5124), 
        .B(n5123), .ZN(n5125) );
  OAI21_X1 U6318 ( .B1(n5132), .B2(n5805), .A(n5125), .ZN(U3009) );
  NAND2_X1 U6319 ( .A1(n6030), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5126)
         );
  OAI211_X1 U6320 ( .C1(n6039), .C2(n5128), .A(n5127), .B(n5126), .ZN(n5129)
         );
  AOI21_X1 U6321 ( .B1(n5130), .B2(n2963), .A(n5129), .ZN(n5131) );
  OAI21_X1 U6322 ( .B1(n5132), .B2(n6011), .A(n5131), .ZN(U2977) );
  OAI21_X1 U6323 ( .B1(n5134), .B2(n5133), .A(REIP_REG_10__SCAN_IN), .ZN(n5139) );
  INV_X1 U6324 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5136) );
  AOI22_X1 U6325 ( .A1(EBX_REG_10__SCAN_IN), .A2(n5943), .B1(n5944), .B2(n6052), .ZN(n5135) );
  OAI211_X1 U6326 ( .C1(n5939), .C2(n5136), .A(n5135), .B(n5887), .ZN(n5137)
         );
  INV_X1 U6327 ( .A(n5137), .ZN(n5138) );
  OAI211_X1 U6328 ( .C1(n5952), .C2(n5162), .A(n5139), .B(n5138), .ZN(n5142)
         );
  INV_X1 U6329 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6420) );
  NOR3_X1 U6330 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6420), .A3(n5140), .ZN(n5141) );
  NOR2_X1 U6331 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  OAI21_X1 U6332 ( .B1(n5880), .B2(n5166), .A(n5143), .ZN(U2817) );
  OAI21_X1 U6333 ( .B1(n5106), .B2(n5145), .A(n5174), .ZN(n5167) );
  AOI22_X1 U6334 ( .A1(n5240), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n5970), .ZN(n5146) );
  OAI21_X1 U6335 ( .B1(n5167), .B2(n5760), .A(n5146), .ZN(U2880) );
  NAND4_X1 U6336 ( .A1(n5938), .A2(n5930), .A3(REIP_REG_2__SCAN_IN), .A4(
        REIP_REG_1__SCAN_IN), .ZN(n5152) );
  INV_X1 U6337 ( .A(n5147), .ZN(n5148) );
  AOI22_X1 U6338 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n5927), .B1(n5928), 
        .B2(n5148), .ZN(n5151) );
  NAND2_X1 U6339 ( .A1(n5922), .A2(n2969), .ZN(n5150) );
  NAND2_X1 U6340 ( .A1(n5943), .A2(EBX_REG_3__SCAN_IN), .ZN(n5149) );
  NAND4_X1 U6341 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .ZN(n5156)
         );
  INV_X1 U6342 ( .A(n5863), .ZN(n5153) );
  OAI21_X1 U6343 ( .B1(n5936), .B2(n5930), .A(n5153), .ZN(n5923) );
  INV_X1 U6344 ( .A(REIP_REG_3__SCAN_IN), .ZN(n5154) );
  NOR2_X1 U6345 ( .A1(n5923), .A2(n5154), .ZN(n5155) );
  AOI211_X1 U6346 ( .C1(n6109), .C2(n5944), .A(n5156), .B(n5155), .ZN(n5157)
         );
  OAI21_X1 U6347 ( .B1(n5159), .B2(n5158), .A(n5157), .ZN(U2824) );
  XNOR2_X1 U6348 ( .A(n5776), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5160)
         );
  XNOR2_X1 U6349 ( .A(n3482), .B(n5160), .ZN(n6054) );
  NAND2_X1 U6350 ( .A1(n6054), .A2(n6035), .ZN(n5165) );
  INV_X1 U6351 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5161) );
  NOR2_X1 U6352 ( .A1(n6123), .A2(n5161), .ZN(n6051) );
  NOR2_X1 U6353 ( .A1(n6039), .A2(n5162), .ZN(n5163) );
  AOI211_X1 U6354 ( .C1(n6030), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6051), 
        .B(n5163), .ZN(n5164) );
  OAI211_X1 U6355 ( .C1(n5579), .C2(n5166), .A(n5165), .B(n5164), .ZN(U2976)
         );
  INV_X1 U6356 ( .A(n5167), .ZN(n6008) );
  NAND2_X1 U6357 ( .A1(n5169), .A2(n5168), .ZN(n5170) );
  NAND2_X1 U6358 ( .A1(n5175), .A2(n5170), .ZN(n5889) );
  INV_X1 U6359 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5890) );
  OAI22_X1 U6360 ( .A1(n5889), .A2(n5455), .B1(n5890), .B2(n5959), .ZN(n5171)
         );
  AOI21_X1 U6361 ( .B1(n6008), .B2(n5956), .A(n5171), .ZN(n5172) );
  INV_X1 U6362 ( .A(n5172), .ZN(U2848) );
  XNOR2_X1 U6363 ( .A(n5174), .B(n5173), .ZN(n5881) );
  AOI21_X1 U6364 ( .B1(n5176), .B2(n5175), .A(n5209), .ZN(n6044) );
  AOI22_X1 U6365 ( .A1(n6044), .A2(n5955), .B1(EBX_REG_12__SCAN_IN), .B2(n5451), .ZN(n5177) );
  OAI21_X1 U6366 ( .B1(n5881), .B2(n5441), .A(n5177), .ZN(U2847) );
  AOI22_X1 U6367 ( .A1(n5240), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n5970), .ZN(n5178) );
  OAI21_X1 U6368 ( .B1(n5881), .B2(n5760), .A(n5178), .ZN(U2879) );
  AOI22_X1 U6369 ( .A1(n5179), .A2(n5776), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n3482), .ZN(n5181) );
  XNOR2_X1 U6370 ( .A(n5581), .B(n5184), .ZN(n5180) );
  XNOR2_X1 U6371 ( .A(n5181), .B(n5180), .ZN(n6012) );
  INV_X1 U6372 ( .A(n5227), .ZN(n6040) );
  AOI22_X1 U6373 ( .A1(n6101), .A2(REIP_REG_11__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6040), .ZN(n5182) );
  OAI21_X1 U6374 ( .B1(n5889), .B2(n6089), .A(n5182), .ZN(n5183) );
  AOI21_X1 U6375 ( .B1(n6043), .B2(n5184), .A(n5183), .ZN(n5185) );
  OAI21_X1 U6376 ( .B1(n6012), .B2(n5805), .A(n5185), .ZN(U3007) );
  NAND2_X1 U6377 ( .A1(n2990), .A2(n5186), .ZN(n5187) );
  XNOR2_X1 U6378 ( .A(n5188), .B(n5187), .ZN(n6045) );
  NAND2_X1 U6379 ( .A1(n6045), .A2(n6035), .ZN(n5193) );
  INV_X1 U6380 ( .A(n5879), .ZN(n5191) );
  INV_X1 U6381 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5189) );
  OAI22_X1 U6382 ( .A1(n5574), .A2(n5877), .B1(n6123), .B2(n5189), .ZN(n5190)
         );
  AOI21_X1 U6383 ( .B1(n6007), .B2(n5191), .A(n5190), .ZN(n5192) );
  OAI211_X1 U6384 ( .C1(n5881), .C2(n5579), .A(n5193), .B(n5192), .ZN(U2974)
         );
  OAI21_X1 U6385 ( .B1(n2988), .B2(n5195), .A(n5194), .ZN(n5871) );
  XNOR2_X1 U6386 ( .A(n5209), .B(n5205), .ZN(n5866) );
  AOI22_X1 U6387 ( .A1(n5866), .A2(n5955), .B1(EBX_REG_13__SCAN_IN), .B2(n5451), .ZN(n5196) );
  OAI21_X1 U6388 ( .B1(n5871), .B2(n5441), .A(n5196), .ZN(U2846) );
  AOI22_X1 U6389 ( .A1(n5240), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n5970), .ZN(n5197) );
  OAI21_X1 U6390 ( .B1(n5871), .B2(n5760), .A(n5197), .ZN(U2878) );
  OAI21_X1 U6391 ( .B1(n5200), .B2(n5199), .A(n5198), .ZN(n5588) );
  INV_X1 U6392 ( .A(n5201), .ZN(n5864) );
  NAND2_X1 U6393 ( .A1(n5864), .A2(n5886), .ZN(n5885) );
  OAI21_X1 U6394 ( .B1(n5869), .B2(n5885), .A(n6425), .ZN(n5215) );
  INV_X1 U6395 ( .A(n5202), .ZN(n5203) );
  NOR2_X1 U6396 ( .A1(n5863), .A2(n5203), .ZN(n5387) );
  INV_X1 U6397 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6653) );
  OAI22_X1 U6398 ( .A1(n6653), .A2(n5924), .B1(n5204), .B2(n5939), .ZN(n5214)
         );
  INV_X1 U6399 ( .A(n5205), .ZN(n5208) );
  INV_X1 U6400 ( .A(n5206), .ZN(n5207) );
  AOI21_X1 U6401 ( .B1(n5209), .B2(n5208), .A(n5207), .ZN(n5210) );
  OR2_X1 U6402 ( .A1(n5243), .A2(n5210), .ZN(n5236) );
  AOI21_X1 U6403 ( .B1(n5928), .B2(n5211), .A(n5926), .ZN(n5212) );
  OAI21_X1 U6404 ( .B1(n5236), .B2(n5910), .A(n5212), .ZN(n5213) );
  AOI211_X1 U6405 ( .C1(n5215), .C2(n5387), .A(n5214), .B(n5213), .ZN(n5216)
         );
  OAI21_X1 U6406 ( .B1(n5588), .B2(n5880), .A(n5216), .ZN(U2813) );
  AOI22_X1 U6407 ( .A1(n5240), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n5970), .ZN(n5217) );
  OAI21_X1 U6408 ( .B1(n5588), .B2(n5760), .A(n5217), .ZN(U2877) );
  INV_X1 U6409 ( .A(n5219), .ZN(n5221) );
  NAND2_X1 U6410 ( .A1(n5221), .A2(n5220), .ZN(n5222) );
  XNOR2_X1 U6411 ( .A(n5218), .B(n5222), .ZN(n5594) );
  AOI21_X1 U6412 ( .B1(n5224), .B2(n5223), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5230) );
  NAND2_X1 U6413 ( .A1(n5225), .A2(n6042), .ZN(n5226) );
  OAI211_X1 U6414 ( .C1(n5229), .C2(n5228), .A(n5227), .B(n5226), .ZN(n5812)
         );
  OAI21_X1 U6415 ( .B1(n5230), .B2(n5812), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5235) );
  NOR3_X1 U6416 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5817), .A3(n5231), 
        .ZN(n5233) );
  OAI22_X1 U6417 ( .A1(n5236), .A2(n6089), .B1(n6425), .B2(n6123), .ZN(n5232)
         );
  NOR2_X1 U6418 ( .A1(n5233), .A2(n5232), .ZN(n5234) );
  OAI211_X1 U6419 ( .C1(n5594), .C2(n5805), .A(n5235), .B(n5234), .ZN(U3004)
         );
  OAI222_X1 U6420 ( .A1(n5236), .A2(n5455), .B1(n5959), .B2(n6653), .C1(n5588), 
        .C2(n5441), .ZN(U2845) );
  AND2_X1 U6421 ( .A1(n5198), .A2(n5237), .ZN(n5239) );
  OR2_X1 U6422 ( .A1(n5239), .A2(n5238), .ZN(n5453) );
  AOI22_X1 U6423 ( .A1(n5240), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5970), .ZN(n5241) );
  OAI21_X1 U6424 ( .B1(n5453), .B2(n5760), .A(n5241), .ZN(U2876) );
  INV_X1 U6425 ( .A(n5584), .ZN(n5249) );
  OR2_X1 U6426 ( .A1(n5243), .A2(n5242), .ZN(n5244) );
  NAND2_X1 U6427 ( .A1(n5391), .A2(n5244), .ZN(n5703) );
  AOI21_X1 U6428 ( .B1(n5927), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5926), 
        .ZN(n5246) );
  AOI22_X1 U6429 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5943), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5387), .ZN(n5245) );
  OAI211_X1 U6430 ( .C1(n5910), .C2(n5703), .A(n5246), .B(n5245), .ZN(n5248)
         );
  NOR2_X1 U6431 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5247), .ZN(n5386) );
  AOI211_X1 U6432 ( .C1(n5928), .C2(n5249), .A(n5248), .B(n5386), .ZN(n5250)
         );
  OAI21_X1 U6433 ( .B1(n5453), .B2(n5880), .A(n5250), .ZN(U2812) );
  NAND2_X1 U6434 ( .A1(n5251), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5256)
         );
  OAI22_X1 U6435 ( .A1(n6496), .A2(n6324), .B1(n5252), .B2(n5258), .ZN(n5253)
         );
  AOI21_X1 U6436 ( .B1(n6317), .B2(n5254), .A(n5253), .ZN(n5255) );
  OAI211_X1 U6437 ( .C1(n5272), .C2(n5257), .A(n5256), .B(n5255), .ZN(U3145)
         );
  NAND2_X1 U6438 ( .A1(n6495), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5263)
         );
  OAI22_X1 U6439 ( .A1(n6496), .A2(n5260), .B1(n5259), .B2(n5258), .ZN(n5261)
         );
  AOI21_X1 U6440 ( .B1(n5266), .B2(n5268), .A(n5261), .ZN(n5262) );
  OAI211_X1 U6441 ( .C1(n6505), .C2(n5272), .A(n5263), .B(n5262), .ZN(U3137)
         );
  AOI22_X1 U6442 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5265), .B1(n6320), 
        .B2(n5264), .ZN(n5270) );
  AOI22_X1 U6443 ( .A1(n5268), .A2(n5267), .B1(n5266), .B2(n6317), .ZN(n5269)
         );
  OAI211_X1 U6444 ( .C1(n5272), .C2(n5271), .A(n5270), .B(n5269), .ZN(U3129)
         );
  INV_X1 U6445 ( .A(n5273), .ZN(n5284) );
  OAI21_X1 U6446 ( .B1(n5276), .B2(n5274), .A(n5275), .ZN(n5277) );
  OAI211_X1 U6447 ( .C1(n5280), .C2(n5279), .A(n5278), .B(n5277), .ZN(n6342)
         );
  INV_X1 U6448 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5281) );
  AOI22_X1 U6449 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5281), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6127), .ZN(n5286) );
  NOR2_X1 U6450 ( .A1(n6374), .A2(n6117), .ZN(n5282) );
  AOI222_X1 U6451 ( .A1(n6342), .A2(n5818), .B1(n5286), .B2(n5282), .C1(n5274), 
        .C2(n5287), .ZN(n5283) );
  OAI22_X1 U6452 ( .A1(n5284), .A2(n3075), .B1(n6471), .B2(n5283), .ZN(U3460)
         );
  AOI21_X1 U6453 ( .B1(n5287), .B2(n5285), .A(n6471), .ZN(n5293) );
  NOR3_X1 U6454 ( .A1(n6374), .A2(n6117), .A3(n5286), .ZN(n5289) );
  AND3_X1 U6455 ( .A1(n5287), .A2(n4521), .A3(n5292), .ZN(n5288) );
  AOI211_X1 U6456 ( .C1(n5290), .C2(n5818), .A(n5289), .B(n5288), .ZN(n5291)
         );
  OAI22_X1 U6457 ( .A1(n5293), .A2(n5292), .B1(n6471), .B2(n5291), .ZN(U3459)
         );
  AOI21_X1 U6458 ( .B1(n4575), .B2(n6276), .A(n6191), .ZN(n5295) );
  AOI22_X1 U6459 ( .A1(n5296), .A2(n5295), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n5294), .ZN(n5297) );
  OAI21_X1 U6460 ( .B1(n4529), .B2(n5298), .A(n5297), .ZN(U3463) );
  AOI22_X1 U6461 ( .A1(n5967), .A2(DATAI_30_), .B1(n5970), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6462 ( .A1(n5971), .A2(DATAI_14_), .ZN(n5299) );
  OAI211_X1 U6463 ( .C1(n4233), .C2(n5760), .A(n5300), .B(n5299), .ZN(U2861)
         );
  INV_X1 U6464 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5301) );
  OAI222_X1 U6465 ( .A1(n5441), .A2(n4233), .B1(n5301), .B2(n5959), .C1(n5598), 
        .C2(n5455), .ZN(U2829) );
  INV_X1 U6466 ( .A(n5460), .ZN(n5313) );
  OAI21_X1 U6467 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5931), .A(n5302), .ZN(n5309) );
  NAND3_X1 U6468 ( .A1(n5303), .A2(REIP_REG_30__SCAN_IN), .A3(n6454), .ZN(
        n5307) );
  AOI22_X1 U6469 ( .A1(n5305), .A2(n5304), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n5927), .ZN(n5306) );
  OAI21_X1 U6470 ( .B1(n5313), .B2(n5880), .A(n5312), .ZN(U2796) );
  AOI21_X1 U6471 ( .B1(n5316), .B2(n5314), .A(n5315), .ZN(n5488) );
  INV_X1 U6472 ( .A(n5488), .ZN(n5465) );
  NAND2_X1 U6473 ( .A1(n5318), .A2(n5317), .ZN(n5321) );
  INV_X1 U6474 ( .A(n5319), .ZN(n5320) );
  NAND2_X1 U6475 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  OR2_X1 U6476 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  INV_X1 U6477 ( .A(n5342), .ZN(n5329) );
  INV_X1 U6478 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6447) );
  OAI22_X1 U6479 ( .A1(n5326), .A2(n5939), .B1(n5952), .B2(n5486), .ZN(n5327)
         );
  AOI21_X1 U6480 ( .B1(n5943), .B2(EBX_REG_29__SCAN_IN), .A(n5327), .ZN(n5328)
         );
  OAI21_X1 U6481 ( .B1(n5329), .B2(n6447), .A(n5328), .ZN(n5331) );
  AOI211_X1 U6482 ( .C1(n5610), .C2(n5944), .A(n5331), .B(n5330), .ZN(n5332)
         );
  OAI21_X1 U6483 ( .B1(n5465), .B2(n5880), .A(n5332), .ZN(U2798) );
  OAI21_X1 U6484 ( .B1(n4311), .B2(n5333), .A(n5314), .ZN(n5498) );
  INV_X1 U6485 ( .A(n5334), .ZN(n5337) );
  INV_X1 U6486 ( .A(n5335), .ZN(n5336) );
  OAI21_X1 U6487 ( .B1(n5337), .B2(n5336), .A(n3000), .ZN(n5614) );
  OAI22_X1 U6488 ( .A1(n5338), .A2(n5939), .B1(n5952), .B2(n5491), .ZN(n5339)
         );
  AOI21_X1 U6489 ( .B1(n5943), .B2(EBX_REG_28__SCAN_IN), .A(n5339), .ZN(n5340)
         );
  OAI21_X1 U6490 ( .B1(n5614), .B2(n5910), .A(n5340), .ZN(n5341) );
  AOI21_X1 U6491 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5342), .A(n5341), .ZN(n5346) );
  INV_X1 U6492 ( .A(n5343), .ZN(n5344) );
  INV_X1 U6493 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5490) );
  NAND3_X1 U6494 ( .A1(n5344), .A2(REIP_REG_27__SCAN_IN), .A3(n5490), .ZN(
        n5345) );
  OAI211_X1 U6495 ( .C1(n5498), .C2(n5880), .A(n5346), .B(n5345), .ZN(U2799)
         );
  INV_X1 U6496 ( .A(n5347), .ZN(n5350) );
  INV_X1 U6497 ( .A(n4079), .ZN(n5349) );
  AOI21_X1 U6498 ( .B1(n5350), .B2(n5349), .A(n5348), .ZN(n5534) );
  INV_X1 U6499 ( .A(n5534), .ZN(n5475) );
  XNOR2_X1 U6500 ( .A(n5413), .B(n5415), .ZN(n5648) );
  INV_X1 U6501 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6439) );
  OAI22_X1 U6502 ( .A1(n5731), .A2(n6439), .B1(n5532), .B2(n5952), .ZN(n5352)
         );
  INV_X1 U6503 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5421) );
  OAI22_X1 U6504 ( .A1(n5421), .A2(n5924), .B1(n6634), .B2(n5939), .ZN(n5351)
         );
  AOI211_X1 U6505 ( .C1(n5648), .C2(n5944), .A(n5352), .B(n5351), .ZN(n5353)
         );
  NAND2_X1 U6506 ( .A1(n5714), .A2(n6439), .ZN(n5728) );
  OAI211_X1 U6507 ( .C1(n5475), .C2(n5880), .A(n5353), .B(n5728), .ZN(U2803)
         );
  OAI21_X1 U6508 ( .B1(n5354), .B2(n5356), .A(n5538), .ZN(n5771) );
  INV_X1 U6509 ( .A(n5371), .ZN(n5853) );
  OAI21_X1 U6510 ( .B1(n5370), .B2(n5853), .A(n5554), .ZN(n5364) );
  INV_X1 U6511 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5429) );
  MUX2_X1 U6512 ( .A(n5373), .B(n5375), .S(n5357), .Z(n5359) );
  XNOR2_X1 U6513 ( .A(n5359), .B(n5358), .ZN(n5680) );
  NAND2_X1 U6514 ( .A1(n5680), .A2(n5944), .ZN(n5362) );
  AOI22_X1 U6515 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n5927), .B1(n5360), 
        .B2(n5928), .ZN(n5361) );
  OAI211_X1 U6516 ( .C1(n5924), .C2(n5429), .A(n5362), .B(n5361), .ZN(n5363)
         );
  AOI21_X1 U6517 ( .B1(n5364), .B2(n5752), .A(n5363), .ZN(n5365) );
  OAI21_X1 U6518 ( .B1(n5771), .B2(n5880), .A(n5365), .ZN(U2807) );
  INV_X1 U6519 ( .A(n5443), .ZN(n5368) );
  INV_X1 U6520 ( .A(n5366), .ZN(n5367) );
  NAND2_X1 U6521 ( .A1(n5368), .A2(n5367), .ZN(n5435) );
  AOI21_X1 U6522 ( .B1(n5369), .B2(n5435), .A(n5354), .ZN(n5566) );
  INV_X1 U6523 ( .A(n5566), .ZN(n5480) );
  OAI211_X1 U6524 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5371), .B(n5370), .ZN(n5383) );
  INV_X1 U6525 ( .A(n5372), .ZN(n5374) );
  MUX2_X1 U6526 ( .A(n5375), .B(n5374), .S(n5373), .Z(n5436) );
  NAND2_X1 U6527 ( .A1(n3004), .A2(n5436), .ZN(n5439) );
  INV_X1 U6528 ( .A(n5376), .ZN(n5377) );
  XNOR2_X1 U6529 ( .A(n5439), .B(n5377), .ZN(n5690) );
  INV_X1 U6530 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6651) );
  AOI21_X1 U6531 ( .B1(n5927), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5926), 
        .ZN(n5380) );
  INV_X1 U6532 ( .A(n5378), .ZN(n5859) );
  AOI22_X1 U6533 ( .A1(n5562), .A2(n5928), .B1(REIP_REG_19__SCAN_IN), .B2(
        n5859), .ZN(n5379) );
  OAI211_X1 U6534 ( .C1(n6651), .C2(n5924), .A(n5380), .B(n5379), .ZN(n5381)
         );
  AOI21_X1 U6535 ( .B1(n5944), .B2(n5690), .A(n5381), .ZN(n5382) );
  OAI211_X1 U6536 ( .C1(n5480), .C2(n5880), .A(n5383), .B(n5382), .ZN(U2808)
         );
  OR2_X1 U6537 ( .A1(n5238), .A2(n5384), .ZN(n5385) );
  NAND2_X1 U6538 ( .A1(n5443), .A2(n5385), .ZN(n5966) );
  OAI33_X1 U6540 ( .A1(1'b0), .A2(n5388), .A3(REIP_REG_16__SCAN_IN), .B1(n6574), .B2(n5387), .B3(n5386), .ZN(n5397) );
  INV_X1 U6541 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5394) );
  INV_X1 U6542 ( .A(n5446), .ZN(n5390) );
  AOI21_X1 U6543 ( .B1(n5392), .B2(n5391), .A(n5390), .ZN(n5696) );
  AOI22_X1 U6544 ( .A1(n5576), .A2(n5928), .B1(n5944), .B2(n5696), .ZN(n5393)
         );
  OAI21_X1 U6545 ( .B1(n5394), .B2(n5924), .A(n5393), .ZN(n5395) );
  AOI211_X1 U6546 ( .C1(n5927), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5926), 
        .B(n5395), .ZN(n5396) );
  OAI211_X1 U6547 ( .C1(n5966), .C2(n5880), .A(n5397), .B(n5396), .ZN(U2811)
         );
  OAI22_X1 U6548 ( .A1(n5399), .A2(n5455), .B1(n5959), .B2(n5398), .ZN(U2828)
         );
  AOI22_X1 U6549 ( .A1(n5610), .A2(n5955), .B1(EBX_REG_29__SCAN_IN), .B2(n5451), .ZN(n5400) );
  OAI21_X1 U6550 ( .B1(n5465), .B2(n5441), .A(n5400), .ZN(U2830) );
  INV_X1 U6551 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5401) );
  OAI222_X1 U6552 ( .A1(n5441), .A2(n5498), .B1(n5401), .B2(n5959), .C1(n5614), 
        .C2(n5455), .ZN(U2831) );
  INV_X1 U6553 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6560) );
  OAI22_X1 U6554 ( .A1(n5624), .A2(n5455), .B1(n6560), .B2(n5959), .ZN(n5402)
         );
  AOI21_X1 U6555 ( .B1(n5506), .B2(n5956), .A(n5402), .ZN(n5403) );
  INV_X1 U6556 ( .A(n5403), .ZN(U2832) );
  NAND2_X1 U6557 ( .A1(n5404), .A2(n5405), .ZN(n5406) );
  AND2_X1 U6558 ( .A1(n4309), .A2(n5406), .ZN(n5761) );
  OR2_X1 U6559 ( .A1(n5417), .A2(n5407), .ZN(n5408) );
  NAND2_X1 U6560 ( .A1(n5409), .A2(n5408), .ZN(n5720) );
  INV_X1 U6561 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5712) );
  OAI22_X1 U6562 ( .A1(n5720), .A2(n5455), .B1(n5712), .B2(n5959), .ZN(n5410)
         );
  AOI21_X1 U6563 ( .B1(n5761), .B2(n5956), .A(n5410), .ZN(n5411) );
  INV_X1 U6564 ( .A(n5411), .ZN(U2833) );
  OAI21_X1 U6565 ( .B1(n5348), .B2(n5412), .A(n5404), .ZN(n5724) );
  INV_X1 U6566 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5419) );
  INV_X1 U6567 ( .A(n5413), .ZN(n5416) );
  AOI21_X1 U6568 ( .B1(n5416), .B2(n5415), .A(n5414), .ZN(n5418) );
  OR2_X1 U6569 ( .A1(n5418), .A2(n5417), .ZN(n5793) );
  OAI222_X1 U6570 ( .A1(n5441), .A2(n5724), .B1(n5959), .B2(n5419), .C1(n5793), 
        .C2(n5455), .ZN(U2834) );
  INV_X1 U6571 ( .A(n5648), .ZN(n5420) );
  OAI222_X1 U6572 ( .A1(n5475), .A2(n5441), .B1(n5959), .B2(n5421), .C1(n5455), 
        .C2(n5420), .ZN(U2835) );
  OAI22_X1 U6573 ( .A1(n5737), .A2(n5455), .B1(n5729), .B2(n5959), .ZN(n5422)
         );
  INV_X1 U6574 ( .A(n5422), .ZN(n5423) );
  OAI21_X1 U6575 ( .B1(n5732), .B2(n5441), .A(n5423), .ZN(U2836) );
  XNOR2_X1 U6576 ( .A(n5538), .B(n5537), .ZN(n5767) );
  OR2_X1 U6577 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  AND2_X1 U6578 ( .A1(n5426), .A2(n5653), .ZN(n5753) );
  AOI22_X1 U6579 ( .A1(n5753), .A2(n5955), .B1(EBX_REG_21__SCAN_IN), .B2(n5451), .ZN(n5427) );
  OAI21_X1 U6580 ( .B1(n5767), .B2(n5441), .A(n5427), .ZN(U2838) );
  INV_X1 U6581 ( .A(n5680), .ZN(n5428) );
  OAI222_X1 U6582 ( .A1(n5441), .A2(n5771), .B1(n5429), .B2(n5959), .C1(n5428), 
        .C2(n5455), .ZN(U2839) );
  NOR2_X1 U6583 ( .A1(n5959), .A2(n6651), .ZN(n5430) );
  AOI21_X1 U6584 ( .B1(n5690), .B2(n5955), .A(n5430), .ZN(n5431) );
  OAI21_X1 U6585 ( .B1(n5480), .B2(n5441), .A(n5431), .ZN(U2840) );
  OR2_X1 U6586 ( .A1(n5443), .A2(n5444), .ZN(n5433) );
  NAND2_X1 U6587 ( .A1(n5433), .A2(n5432), .ZN(n5434) );
  INV_X1 U6588 ( .A(n5960), .ZN(n5442) );
  INV_X1 U6589 ( .A(n5436), .ZN(n5437) );
  NAND2_X1 U6590 ( .A1(n5448), .A2(n5437), .ZN(n5438) );
  AND2_X1 U6591 ( .A1(n5439), .A2(n5438), .ZN(n5850) );
  AOI22_X1 U6592 ( .A1(n5850), .A2(n5955), .B1(EBX_REG_18__SCAN_IN), .B2(n5451), .ZN(n5440) );
  OAI21_X1 U6593 ( .B1(n5442), .B2(n5441), .A(n5440), .ZN(U2841) );
  XOR2_X1 U6594 ( .A(n5444), .B(n5443), .Z(n5963) );
  NAND2_X1 U6595 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  NAND2_X1 U6596 ( .A1(n5448), .A2(n5447), .ZN(n5862) );
  INV_X1 U6597 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6654) );
  OAI22_X1 U6598 ( .A1(n5862), .A2(n5455), .B1(n6654), .B2(n5959), .ZN(n5449)
         );
  AOI21_X1 U6599 ( .B1(n5963), .B2(n5956), .A(n5449), .ZN(n5450) );
  INV_X1 U6600 ( .A(n5450), .ZN(U2842) );
  AOI22_X1 U6601 ( .A1(n5696), .A2(n5955), .B1(EBX_REG_16__SCAN_IN), .B2(n5451), .ZN(n5452) );
  OAI21_X1 U6602 ( .B1(n5966), .B2(n5441), .A(n5452), .ZN(U2843) );
  INV_X1 U6603 ( .A(n5453), .ZN(n5586) );
  INV_X1 U6604 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5454) );
  OAI22_X1 U6605 ( .A1(n5703), .A2(n5455), .B1(n5454), .B2(n5959), .ZN(n5456)
         );
  AOI21_X1 U6606 ( .B1(n5586), .B2(n5956), .A(n5456), .ZN(n5457) );
  INV_X1 U6607 ( .A(n5457), .ZN(U2844) );
  NAND3_X1 U6608 ( .A1(n5460), .A2(n5459), .A3(n5458), .ZN(n5462) );
  AOI22_X1 U6609 ( .A1(n5967), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5970), .ZN(n5461) );
  NAND2_X1 U6610 ( .A1(n5462), .A2(n5461), .ZN(U2860) );
  AOI22_X1 U6611 ( .A1(n5967), .A2(DATAI_29_), .B1(n5970), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6612 ( .A1(n5971), .A2(DATAI_13_), .ZN(n5463) );
  OAI211_X1 U6613 ( .C1(n5465), .C2(n5760), .A(n5464), .B(n5463), .ZN(U2862)
         );
  AOI22_X1 U6614 ( .A1(n5967), .A2(DATAI_28_), .B1(n5970), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U6615 ( .A1(n5971), .A2(DATAI_12_), .ZN(n5466) );
  OAI211_X1 U6616 ( .C1(n5498), .C2(n5760), .A(n5467), .B(n5466), .ZN(U2863)
         );
  AOI22_X1 U6617 ( .A1(n5967), .A2(DATAI_27_), .B1(n5970), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6618 ( .A1(n5971), .A2(DATAI_11_), .ZN(n5468) );
  OAI211_X1 U6619 ( .C1(n5470), .C2(n5760), .A(n5469), .B(n5468), .ZN(U2864)
         );
  AOI22_X1 U6620 ( .A1(n5971), .A2(DATAI_9_), .B1(n5970), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6621 ( .A1(n5967), .A2(DATAI_25_), .ZN(n5471) );
  OAI211_X1 U6622 ( .C1(n5724), .C2(n5760), .A(n5472), .B(n5471), .ZN(U2866)
         );
  AOI22_X1 U6623 ( .A1(n5967), .A2(DATAI_24_), .B1(n5970), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6624 ( .A1(n5971), .A2(DATAI_8_), .ZN(n5473) );
  OAI211_X1 U6625 ( .C1(n5475), .C2(n5760), .A(n5474), .B(n5473), .ZN(U2867)
         );
  AOI22_X1 U6626 ( .A1(n5971), .A2(DATAI_7_), .B1(n5970), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6627 ( .A1(n5967), .A2(DATAI_23_), .ZN(n5476) );
  OAI211_X1 U6628 ( .C1(n5732), .C2(n5760), .A(n5477), .B(n5476), .ZN(U2868)
         );
  AOI22_X1 U6629 ( .A1(n5967), .A2(DATAI_19_), .B1(n5970), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6630 ( .A1(n5971), .A2(DATAI_3_), .ZN(n5478) );
  OAI211_X1 U6631 ( .C1(n5480), .C2(n5760), .A(n5479), .B(n5478), .ZN(U2872)
         );
  INV_X1 U6632 ( .A(n5481), .ZN(n5512) );
  OAI22_X1 U6633 ( .A1(n5483), .A2(n5493), .B1(n5512), .B2(n5482), .ZN(n5484)
         );
  XNOR2_X1 U6634 ( .A(n5484), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5612)
         );
  NOR2_X1 U6635 ( .A1(n6123), .A2(n6447), .ZN(n5603) );
  AOI21_X1 U6636 ( .B1(n6030), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5603), 
        .ZN(n5485) );
  OAI21_X1 U6637 ( .B1(n5486), .B2(n6039), .A(n5485), .ZN(n5487) );
  AOI21_X1 U6638 ( .B1(n5488), .B2(n2963), .A(n5487), .ZN(n5489) );
  OAI21_X1 U6639 ( .B1(n5612), .B2(n6011), .A(n5489), .ZN(U2957) );
  NOR2_X1 U6640 ( .A1(n6123), .A2(n5490), .ZN(n5618) );
  NOR2_X1 U6641 ( .A1(n6039), .A2(n5491), .ZN(n5492) );
  AOI211_X1 U6642 ( .C1(n6030), .C2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5618), 
        .B(n5492), .ZN(n5497) );
  INV_X1 U6643 ( .A(n5493), .ZN(n5499) );
  OAI22_X1 U6644 ( .A1(n5494), .A2(n5499), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5635), .ZN(n5495) );
  NAND2_X1 U6645 ( .A1(n5613), .A2(n6035), .ZN(n5496) );
  OAI211_X1 U6646 ( .C1(n5498), .C2(n5579), .A(n5497), .B(n5496), .ZN(U2958)
         );
  INV_X1 U6647 ( .A(n4217), .ZN(n5500) );
  AOI21_X1 U6648 ( .B1(n5500), .B2(n5508), .A(n5499), .ZN(n5501) );
  XOR2_X1 U6649 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(n5501), .Z(n5632) );
  NAND2_X1 U6650 ( .A1(n6007), .A2(n5502), .ZN(n5503) );
  NAND2_X1 U6651 ( .A1(n6101), .A2(REIP_REG_27__SCAN_IN), .ZN(n5625) );
  OAI211_X1 U6652 ( .C1(n5574), .C2(n5504), .A(n5503), .B(n5625), .ZN(n5505)
         );
  AOI21_X1 U6653 ( .B1(n5506), .B2(n2963), .A(n5505), .ZN(n5507) );
  OAI21_X1 U6654 ( .B1(n5632), .B2(n6011), .A(n5507), .ZN(U2959) );
  INV_X1 U6655 ( .A(n5508), .ZN(n5510) );
  NAND2_X1 U6656 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  XNOR2_X1 U6657 ( .A(n5512), .B(n5511), .ZN(n5642) );
  INV_X1 U6658 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6443) );
  NOR2_X1 U6659 ( .A1(n6123), .A2(n6443), .ZN(n5638) );
  AOI21_X1 U6660 ( .B1(n6030), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5638), 
        .ZN(n5513) );
  OAI21_X1 U6661 ( .B1(n5711), .B2(n6039), .A(n5513), .ZN(n5514) );
  AOI21_X1 U6662 ( .B1(n5761), .B2(n2963), .A(n5514), .ZN(n5515) );
  OAI21_X1 U6663 ( .B1(n5642), .B2(n6011), .A(n5515), .ZN(U2960) );
  INV_X1 U6664 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5517) );
  INV_X1 U6665 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5516) );
  OAI22_X1 U6666 ( .A1(n5574), .A2(n5517), .B1(n6123), .B2(n5516), .ZN(n5518)
         );
  AOI21_X1 U6667 ( .B1(n6007), .B2(n5721), .A(n5518), .ZN(n5522) );
  OAI21_X1 U6668 ( .B1(n5520), .B2(n5519), .A(n4217), .ZN(n5795) );
  NAND2_X1 U6669 ( .A1(n5795), .A2(n6035), .ZN(n5521) );
  OAI211_X1 U6670 ( .C1(n5724), .C2(n5579), .A(n5522), .B(n5521), .ZN(U2961)
         );
  NAND2_X1 U6671 ( .A1(n5523), .A2(n5524), .ZN(n5528) );
  NAND2_X1 U6672 ( .A1(n5547), .A2(n3069), .ZN(n5542) );
  INV_X1 U6673 ( .A(n5542), .ZN(n5526) );
  NAND2_X1 U6674 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  NAND2_X1 U6675 ( .A1(n5528), .A2(n5527), .ZN(n5530) );
  XNOR2_X1 U6676 ( .A(n5530), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5650)
         );
  NOR2_X1 U6677 ( .A1(n6123), .A2(n6439), .ZN(n5647) );
  AOI21_X1 U6678 ( .B1(n6030), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5647), 
        .ZN(n5531) );
  OAI21_X1 U6679 ( .B1(n5532), .B2(n6039), .A(n5531), .ZN(n5533) );
  AOI21_X1 U6680 ( .B1(n5534), .B2(n2963), .A(n5533), .ZN(n5535) );
  OAI21_X1 U6681 ( .B1(n5650), .B2(n6011), .A(n5535), .ZN(U2962) );
  OAI21_X1 U6682 ( .B1(n5538), .B2(n5537), .A(n5536), .ZN(n5539) );
  NAND2_X1 U6683 ( .A1(n5539), .A2(n4035), .ZN(n5740) );
  OAI21_X1 U6684 ( .B1(n5776), .B2(n5661), .A(n5540), .ZN(n5541) );
  XNOR2_X1 U6685 ( .A(n5542), .B(n5541), .ZN(n5651) );
  NAND2_X1 U6686 ( .A1(n5651), .A2(n6035), .ZN(n5546) );
  INV_X1 U6687 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5543) );
  NOR2_X1 U6688 ( .A1(n6123), .A2(n5543), .ZN(n5658) );
  NOR2_X1 U6689 ( .A1(n6039), .A2(n5738), .ZN(n5544) );
  AOI211_X1 U6690 ( .C1(n6030), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5658), 
        .B(n5544), .ZN(n5545) );
  OAI211_X1 U6691 ( .C1(n5579), .C2(n5740), .A(n5546), .B(n5545), .ZN(U2964)
         );
  OAI21_X1 U6692 ( .B1(n5549), .B2(n5548), .A(n5547), .ZN(n5662) );
  NAND2_X1 U6693 ( .A1(n5662), .A2(n6035), .ZN(n5552) );
  NAND2_X1 U6694 ( .A1(n6101), .A2(REIP_REG_21__SCAN_IN), .ZN(n5663) );
  OAI21_X1 U6695 ( .B1(n5574), .B2(n6571), .A(n5663), .ZN(n5550) );
  AOI21_X1 U6696 ( .B1(n6007), .B2(n5748), .A(n5550), .ZN(n5551) );
  OAI211_X1 U6697 ( .C1(n5579), .C2(n5767), .A(n5552), .B(n5551), .ZN(U2965)
         );
  XOR2_X1 U6698 ( .A(n5553), .B(n3495), .Z(n5675) );
  NAND2_X1 U6699 ( .A1(n5675), .A2(n6035), .ZN(n5558) );
  INV_X1 U6700 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5554) );
  NOR2_X1 U6701 ( .A1(n6123), .A2(n5554), .ZN(n5679) );
  NOR2_X1 U6702 ( .A1(n5555), .A2(n6039), .ZN(n5556) );
  AOI211_X1 U6703 ( .C1(n6030), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5679), 
        .B(n5556), .ZN(n5557) );
  OAI211_X1 U6704 ( .C1(n5579), .C2(n5771), .A(n5558), .B(n5557), .ZN(U2966)
         );
  AOI21_X1 U6705 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5559), .A(n5560), 
        .ZN(n5561) );
  XNOR2_X1 U6706 ( .A(n5561), .B(n5776), .ZN(n5692) );
  INV_X1 U6707 ( .A(n5562), .ZN(n5564) );
  NAND2_X1 U6708 ( .A1(n6030), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5563)
         );
  NAND2_X1 U6709 ( .A1(n6101), .A2(REIP_REG_19__SCAN_IN), .ZN(n5684) );
  OAI211_X1 U6710 ( .C1(n6039), .C2(n5564), .A(n5563), .B(n5684), .ZN(n5565)
         );
  AOI21_X1 U6711 ( .B1(n5566), .B2(n2963), .A(n5565), .ZN(n5567) );
  OAI21_X1 U6712 ( .B1(n5692), .B2(n6011), .A(n5567), .ZN(U2967) );
  INV_X1 U6713 ( .A(n5569), .ZN(n5571) );
  NOR2_X1 U6714 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  XNOR2_X1 U6715 ( .A(n5568), .B(n5572), .ZN(n5694) );
  NAND2_X1 U6716 ( .A1(n5694), .A2(n6035), .ZN(n5578) );
  NOR2_X1 U6717 ( .A1(n6123), .A2(n6574), .ZN(n5699) );
  INV_X1 U6718 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5573) );
  NOR2_X1 U6719 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  AOI211_X1 U6720 ( .C1(n6007), .C2(n5576), .A(n5699), .B(n5575), .ZN(n5577)
         );
  OAI211_X1 U6721 ( .C1(n5579), .C2(n5966), .A(n5578), .B(n5577), .ZN(U2970)
         );
  XNOR2_X1 U6722 ( .A(n5581), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5582)
         );
  XNOR2_X1 U6723 ( .A(n5580), .B(n5582), .ZN(n5710) );
  AOI22_X1 U6724 ( .A1(n6030), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6101), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5583) );
  OAI21_X1 U6725 ( .B1(n5584), .B2(n6039), .A(n5583), .ZN(n5585) );
  AOI21_X1 U6726 ( .B1(n5586), .B2(n2963), .A(n5585), .ZN(n5587) );
  OAI21_X1 U6727 ( .B1(n5710), .B2(n6011), .A(n5587), .ZN(U2971) );
  INV_X1 U6728 ( .A(n5588), .ZN(n5592) );
  AOI22_X1 U6729 ( .A1(n6030), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6101), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5589) );
  OAI21_X1 U6730 ( .B1(n6039), .B2(n5590), .A(n5589), .ZN(n5591) );
  AOI21_X1 U6731 ( .B1(n5592), .B2(n2963), .A(n5591), .ZN(n5593) );
  OAI21_X1 U6732 ( .B1(n5594), .B2(n6011), .A(n5593), .ZN(U2972) );
  OR3_X1 U6733 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5595), 
        .ZN(n5596) );
  OAI211_X1 U6734 ( .C1(n5598), .C2(n6089), .A(n5597), .B(n5596), .ZN(n5599)
         );
  AOI21_X1 U6735 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5600), .A(n5599), 
        .ZN(n5601) );
  OAI21_X1 U6736 ( .B1(n5602), .B2(n5805), .A(n5601), .ZN(U2988) );
  NAND2_X1 U6737 ( .A1(n5616), .A2(n5606), .ZN(n5605) );
  INV_X1 U6738 ( .A(n5603), .ZN(n5604) );
  OAI21_X1 U6739 ( .B1(n5626), .B2(n5605), .A(n5604), .ZN(n5609) );
  NOR2_X1 U6740 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  AOI211_X1 U6741 ( .C1(n6121), .C2(n5610), .A(n5609), .B(n5608), .ZN(n5611)
         );
  OAI21_X1 U6742 ( .B1(n5612), .B2(n5805), .A(n5611), .ZN(U2989) );
  INV_X1 U6743 ( .A(n5629), .ZN(n5623) );
  NAND2_X1 U6744 ( .A1(n5613), .A2(n6129), .ZN(n5621) );
  INV_X1 U6745 ( .A(n5614), .ZN(n5619) );
  NOR3_X1 U6746 ( .A1(n5626), .A2(n5616), .A3(n5615), .ZN(n5617) );
  AOI211_X1 U6747 ( .C1(n5619), .C2(n6121), .A(n5618), .B(n5617), .ZN(n5620)
         );
  OAI211_X1 U6748 ( .C1(n5623), .C2(n5622), .A(n5621), .B(n5620), .ZN(U2990)
         );
  INV_X1 U6749 ( .A(n5624), .ZN(n5628) );
  OAI21_X1 U6750 ( .B1(n5626), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5625), 
        .ZN(n5627) );
  AOI21_X1 U6751 ( .B1(n5628), .B2(n6121), .A(n5627), .ZN(n5631) );
  NAND2_X1 U6752 ( .A1(n5629), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5630) );
  OAI211_X1 U6753 ( .C1(n5632), .C2(n5805), .A(n5631), .B(n5630), .ZN(U2991)
         );
  INV_X1 U6754 ( .A(n5720), .ZN(n5639) );
  INV_X1 U6755 ( .A(n5633), .ZN(n5634) );
  AOI211_X1 U6756 ( .C1(n5636), .C2(n5635), .A(n5634), .B(n5798), .ZN(n5637)
         );
  AOI211_X1 U6757 ( .C1(n5639), .C2(n6121), .A(n5638), .B(n5637), .ZN(n5641)
         );
  INV_X1 U6758 ( .A(n5645), .ZN(n5792) );
  NAND2_X1 U6759 ( .A1(n5792), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5640) );
  OAI211_X1 U6760 ( .C1(n5642), .C2(n5805), .A(n5641), .B(n5640), .ZN(U2992)
         );
  AOI21_X1 U6761 ( .B1(n5643), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5644) );
  NOR2_X1 U6762 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  AOI211_X1 U6763 ( .C1(n6121), .C2(n5648), .A(n5647), .B(n5646), .ZN(n5649)
         );
  OAI21_X1 U6764 ( .B1(n5650), .B2(n5805), .A(n5649), .ZN(U2994) );
  NAND2_X1 U6765 ( .A1(n5651), .A2(n6129), .ZN(n5660) );
  XNOR2_X1 U6766 ( .A(n5653), .B(n5652), .ZN(n5758) );
  OR2_X1 U6767 ( .A1(n5654), .A2(n5811), .ZN(n5664) );
  NOR3_X1 U6768 ( .A1(n5664), .A2(n5656), .A3(n5655), .ZN(n5657) );
  AOI211_X1 U6769 ( .C1(n5758), .C2(n6121), .A(n5658), .B(n5657), .ZN(n5659)
         );
  OAI211_X1 U6770 ( .C1(n5668), .C2(n5661), .A(n5660), .B(n5659), .ZN(U2996)
         );
  INV_X1 U6771 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U6772 ( .A1(n5662), .A2(n6129), .ZN(n5667) );
  OAI21_X1 U6773 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5664), .A(n5663), 
        .ZN(n5665) );
  AOI21_X1 U6774 ( .B1(n5753), .B2(n6121), .A(n5665), .ZN(n5666) );
  OAI211_X1 U6775 ( .C1(n5668), .C2(n6551), .A(n5667), .B(n5666), .ZN(U2997)
         );
  INV_X1 U6776 ( .A(n5669), .ZN(n5671) );
  INV_X1 U6777 ( .A(n6041), .ZN(n5670) );
  NAND2_X1 U6778 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  AOI21_X1 U6779 ( .B1(n6529), .B2(n5672), .A(n5808), .ZN(n5804) );
  INV_X1 U6780 ( .A(n5804), .ZN(n5673) );
  AOI21_X1 U6781 ( .B1(n5803), .B2(n5674), .A(n5673), .ZN(n5687) );
  INV_X1 U6782 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U6783 ( .A1(n5675), .A2(n6129), .ZN(n5682) );
  NOR3_X1 U6784 ( .A1(n5685), .A2(n5677), .A3(n5676), .ZN(n5678) );
  AOI211_X1 U6785 ( .C1(n5680), .C2(n6121), .A(n5679), .B(n5678), .ZN(n5681)
         );
  OAI211_X1 U6786 ( .C1(n5687), .C2(n5683), .A(n5682), .B(n5681), .ZN(U2998)
         );
  OAI21_X1 U6787 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5685), .A(n5684), 
        .ZN(n5689) );
  INV_X1 U6788 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5686) );
  NOR2_X1 U6789 ( .A1(n5687), .A2(n5686), .ZN(n5688) );
  AOI211_X1 U6790 ( .C1(n6121), .C2(n5690), .A(n5689), .B(n5688), .ZN(n5691)
         );
  OAI21_X1 U6791 ( .B1(n5692), .B2(n5805), .A(n5691), .ZN(U2999) );
  INV_X1 U6792 ( .A(n5693), .ZN(n5704) );
  NAND2_X1 U6793 ( .A1(n5694), .A2(n6129), .ZN(n5702) );
  AOI21_X1 U6794 ( .B1(n5707), .B2(n5775), .A(n5695), .ZN(n5700) );
  INV_X1 U6795 ( .A(n5696), .ZN(n5697) );
  NOR2_X1 U6796 ( .A1(n5697), .A2(n6089), .ZN(n5698) );
  AOI211_X1 U6797 ( .C1(n5700), .C2(n5708), .A(n5699), .B(n5698), .ZN(n5701)
         );
  OAI211_X1 U6798 ( .C1(n5704), .C2(n5775), .A(n5702), .B(n5701), .ZN(U3002)
         );
  OAI22_X1 U6799 ( .A1(n5703), .A2(n6089), .B1(n6427), .B2(n6123), .ZN(n5706)
         );
  NOR2_X1 U6800 ( .A1(n5704), .A2(n5707), .ZN(n5705) );
  AOI211_X1 U6801 ( .C1(n5708), .C2(n5707), .A(n5706), .B(n5705), .ZN(n5709)
         );
  OAI21_X1 U6802 ( .B1(n5710), .B2(n5805), .A(n5709), .ZN(U3003) );
  AND2_X1 U6803 ( .A1(n5993), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OAI22_X1 U6804 ( .A1(n5712), .A2(n5924), .B1(n5711), .B2(n5952), .ZN(n5713)
         );
  AOI21_X1 U6805 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5927), .A(n5713), 
        .ZN(n5719) );
  NAND2_X1 U6806 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5714), .ZN(n5723) );
  OAI21_X1 U6807 ( .B1(n5516), .B2(n5723), .A(n6443), .ZN(n5717) );
  INV_X1 U6808 ( .A(n5715), .ZN(n5716) );
  AOI22_X1 U6809 ( .A1(n5761), .A2(n5907), .B1(n5717), .B2(n5716), .ZN(n5718)
         );
  OAI211_X1 U6810 ( .C1(n5720), .C2(n5910), .A(n5719), .B(n5718), .ZN(U2801)
         );
  AOI22_X1 U6811 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n5927), .B1(n5721), 
        .B2(n5928), .ZN(n5722) );
  OAI21_X1 U6812 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5723), .A(n5722), .ZN(n5726) );
  OAI22_X1 U6813 ( .A1(n5724), .A2(n5880), .B1(n5910), .B2(n5793), .ZN(n5725)
         );
  AOI211_X1 U6814 ( .C1(EBX_REG_25__SCAN_IN), .C2(n5943), .A(n5726), .B(n5725), 
        .ZN(n5727) );
  OAI221_X1 U6815 ( .B1(n5516), .B2(n5731), .C1(n5516), .C2(n5728), .A(n5727), 
        .ZN(U2802) );
  OAI22_X1 U6816 ( .A1(n5729), .A2(n5924), .B1(n4031), .B2(n5939), .ZN(n5734)
         );
  INV_X1 U6817 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6561) );
  NOR2_X1 U6818 ( .A1(n5543), .A2(n6561), .ZN(n5741) );
  INV_X1 U6819 ( .A(n5742), .ZN(n5751) );
  AOI21_X1 U6820 ( .B1(n5741), .B2(n5751), .A(REIP_REG_23__SCAN_IN), .ZN(n5730) );
  OAI22_X1 U6821 ( .A1(n5732), .A2(n5880), .B1(n5731), .B2(n5730), .ZN(n5733)
         );
  AOI211_X1 U6822 ( .C1(n5735), .C2(n5928), .A(n5734), .B(n5733), .ZN(n5736)
         );
  OAI21_X1 U6823 ( .B1(n5737), .B2(n5910), .A(n5736), .ZN(U2804) );
  AOI22_X1 U6824 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5943), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5927), .ZN(n5747) );
  INV_X1 U6825 ( .A(n5738), .ZN(n5739) );
  AOI22_X1 U6826 ( .A1(n5739), .A2(n5928), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5752), .ZN(n5746) );
  AOI22_X1 U6827 ( .A1(n5764), .A2(n5907), .B1(n5944), .B2(n5758), .ZN(n5745)
         );
  AOI211_X1 U6828 ( .C1(n5543), .C2(n6561), .A(n5742), .B(n5741), .ZN(n5743)
         );
  INV_X1 U6829 ( .A(n5743), .ZN(n5744) );
  NAND4_X1 U6830 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(U2805)
         );
  AOI22_X1 U6831 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5943), .B1(n5748), .B2(n5928), .ZN(n5749) );
  OAI21_X1 U6832 ( .B1(n6571), .B2(n5939), .A(n5749), .ZN(n5750) );
  AOI221_X1 U6833 ( .B1(n5752), .B2(REIP_REG_21__SCAN_IN), .C1(n5751), .C2(
        n6561), .A(n5750), .ZN(n5757) );
  OR2_X1 U6834 ( .A1(n5767), .A2(n5880), .ZN(n5755) );
  NAND2_X1 U6835 ( .A1(n5753), .A2(n5944), .ZN(n5754) );
  AND2_X1 U6836 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  NAND2_X1 U6837 ( .A1(n5757), .A2(n5756), .ZN(U2806) );
  INV_X1 U6838 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6517) );
  AOI22_X1 U6839 ( .A1(n5764), .A2(n5956), .B1(n5955), .B2(n5758), .ZN(n5759)
         );
  OAI21_X1 U6840 ( .B1(n5959), .B2(n6517), .A(n5759), .ZN(U2837) );
  INV_X1 U6841 ( .A(n5760), .ZN(n5968) );
  AOI22_X1 U6842 ( .A1(n5761), .A2(n5968), .B1(n5967), .B2(DATAI_26_), .ZN(
        n5763) );
  AOI22_X1 U6843 ( .A1(n5971), .A2(DATAI_10_), .B1(n5970), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U6844 ( .A1(n5763), .A2(n5762), .ZN(U2865) );
  AOI22_X1 U6845 ( .A1(n5764), .A2(n5968), .B1(n5967), .B2(DATAI_22_), .ZN(
        n5766) );
  AOI22_X1 U6846 ( .A1(n5971), .A2(DATAI_6_), .B1(n5970), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U6847 ( .A1(n5766), .A2(n5765), .ZN(U2869) );
  INV_X1 U6848 ( .A(n5767), .ZN(n5768) );
  AOI22_X1 U6849 ( .A1(n5768), .A2(n5968), .B1(n5967), .B2(DATAI_21_), .ZN(
        n5770) );
  AOI22_X1 U6850 ( .A1(n5971), .A2(DATAI_5_), .B1(n5970), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U6851 ( .A1(n5770), .A2(n5769), .ZN(U2870) );
  INV_X1 U6852 ( .A(n5771), .ZN(n5772) );
  AOI22_X1 U6853 ( .A1(n5772), .A2(n5968), .B1(n5967), .B2(DATAI_20_), .ZN(
        n5774) );
  AOI22_X1 U6854 ( .A1(n5971), .A2(DATAI_4_), .B1(n5970), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U6855 ( .A1(n5774), .A2(n5773), .ZN(U2871) );
  AOI22_X1 U6856 ( .A1(n6101), .A2(REIP_REG_18__SCAN_IN), .B1(n6030), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5780) );
  NAND3_X1 U6857 ( .A1(n5568), .A2(n5776), .A3(n5775), .ZN(n5781) );
  NOR3_X1 U6858 ( .A1(n5568), .A2(n5776), .A3(n5775), .ZN(n5783) );
  NAND2_X1 U6859 ( .A1(n5783), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5777) );
  OAI21_X1 U6860 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5781), .A(n5777), 
        .ZN(n5778) );
  XNOR2_X1 U6861 ( .A(n5778), .B(n5803), .ZN(n5800) );
  AOI22_X1 U6862 ( .A1(n5800), .A2(n6035), .B1(n2963), .B2(n5960), .ZN(n5779)
         );
  OAI211_X1 U6863 ( .C1(n6039), .C2(n5848), .A(n5780), .B(n5779), .ZN(U2968)
         );
  INV_X1 U6864 ( .A(n5781), .ZN(n5782) );
  NOR2_X1 U6865 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  XNOR2_X1 U6866 ( .A(n5784), .B(n6529), .ZN(n5806) );
  AOI22_X1 U6867 ( .A1(n6101), .A2(REIP_REG_17__SCAN_IN), .B1(n6030), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5786) );
  AOI22_X1 U6868 ( .A1(n5963), .A2(n2963), .B1(n6007), .B2(n5856), .ZN(n5785)
         );
  OAI211_X1 U6869 ( .C1(n5806), .C2(n6011), .A(n5786), .B(n5785), .ZN(U2969)
         );
  AOI22_X1 U6870 ( .A1(n6101), .A2(REIP_REG_13__SCAN_IN), .B1(n6030), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5791) );
  XNOR2_X1 U6871 ( .A(n5788), .B(n5787), .ZN(n5813) );
  INV_X1 U6872 ( .A(n5871), .ZN(n5789) );
  AOI22_X1 U6873 ( .A1(n5813), .A2(n6035), .B1(n2963), .B2(n5789), .ZN(n5790)
         );
  OAI211_X1 U6874 ( .C1(n6039), .C2(n5875), .A(n5791), .B(n5790), .ZN(U2973)
         );
  AOI22_X1 U6875 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n5792), .B1(n6101), .B2(REIP_REG_25__SCAN_IN), .ZN(n5797) );
  INV_X1 U6876 ( .A(n5793), .ZN(n5794) );
  AOI22_X1 U6877 ( .A1(n5795), .A2(n6129), .B1(n6121), .B2(n5794), .ZN(n5796)
         );
  OAI211_X1 U6878 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5798), .A(n5797), .B(n5796), .ZN(U2993) );
  AOI22_X1 U6879 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6101), .B1(n5799), .B2(
        n5803), .ZN(n5802) );
  AOI22_X1 U6880 ( .A1(n5800), .A2(n6129), .B1(n6121), .B2(n5850), .ZN(n5801)
         );
  OAI211_X1 U6881 ( .C1(n5804), .C2(n5803), .A(n5802), .B(n5801), .ZN(U3000)
         );
  OAI22_X1 U6882 ( .A1(n5806), .A2(n5805), .B1(n6089), .B2(n5862), .ZN(n5807)
         );
  AOI21_X1 U6883 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5808), .A(n5807), 
        .ZN(n5810) );
  NAND2_X1 U6884 ( .A1(n6101), .A2(REIP_REG_17__SCAN_IN), .ZN(n5809) );
  OAI211_X1 U6885 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5811), .A(n5810), .B(n5809), .ZN(U3001) );
  OR2_X1 U6886 ( .A1(n6042), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5816)
         );
  AOI22_X1 U6887 ( .A1(n5866), .A2(n6121), .B1(n6101), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5815) );
  AOI22_X1 U6888 ( .A1(n5813), .A2(n6129), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5812), .ZN(n5814) );
  OAI211_X1 U6889 ( .C1(n5817), .C2(n5816), .A(n5815), .B(n5814), .ZN(U3005)
         );
  NAND4_X1 U6890 ( .A1(n5820), .A2(n5819), .A3(n5818), .A4(n5921), .ZN(n5821)
         );
  OAI21_X1 U6891 ( .B1(n5822), .B2(n6646), .A(n5821), .ZN(U3455) );
  INV_X1 U6892 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6409) );
  AOI21_X1 U6893 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6409), .A(n6403), .ZN(n5827) );
  INV_X1 U6894 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5823) );
  NOR2_X1 U6895 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6399), .ZN(n6494) );
  AOI21_X1 U6896 ( .B1(n5827), .B2(n5823), .A(n6494), .ZN(U2789) );
  OAI21_X1 U6897 ( .B1(n5824), .B2(n6384), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5825) );
  OAI21_X1 U6898 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6385), .A(n5825), .ZN(
        U2790) );
  INV_X1 U6899 ( .A(n6494), .ZN(n6482) );
  NOR2_X1 U6900 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5828) );
  OAI21_X1 U6901 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5828), .A(n6448), .ZN(n5826)
         );
  OAI21_X1 U6902 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6482), .A(n5826), .ZN(
        U2791) );
  NOR2_X1 U6903 ( .A1(n6494), .A2(n5827), .ZN(n6461) );
  OAI21_X1 U6904 ( .B1(n5828), .B2(BS16_N), .A(n6461), .ZN(n6459) );
  OAI21_X1 U6905 ( .B1(n6461), .B2(n5829), .A(n6459), .ZN(U2792) );
  OAI21_X1 U6906 ( .B1(n5831), .B2(n5830), .A(n6011), .ZN(U2793) );
  NOR4_X1 U6907 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5835) );
  NOR4_X1 U6908 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5834) );
  NOR4_X1 U6909 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5833) );
  NOR4_X1 U6910 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5832) );
  NAND4_X1 U6911 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n5841)
         );
  NOR4_X1 U6912 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5839) );
  AOI211_X1 U6913 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_7__SCAN_IN), .B(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n5838) );
  NOR4_X1 U6914 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n5837)
         );
  NOR4_X1 U6915 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5836) );
  NAND4_X1 U6916 ( .A1(n5839), .A2(n5838), .A3(n5837), .A4(n5836), .ZN(n5840)
         );
  NOR2_X1 U6917 ( .A1(n5841), .A2(n5840), .ZN(n6476) );
  INV_X1 U6918 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5843) );
  NOR3_X1 U6919 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5844) );
  OAI21_X1 U6920 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5844), .A(n6476), .ZN(n5842)
         );
  OAI21_X1 U6921 ( .B1(n6476), .B2(n5843), .A(n5842), .ZN(U2794) );
  INV_X1 U6922 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6573) );
  INV_X1 U6923 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6460) );
  AOI21_X1 U6924 ( .B1(n6573), .B2(n6460), .A(n5844), .ZN(n5846) );
  INV_X1 U6925 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5845) );
  INV_X1 U6926 ( .A(n6476), .ZN(n6479) );
  AOI22_X1 U6927 ( .A1(n6476), .A2(n5846), .B1(n5845), .B2(n6479), .ZN(U2795)
         );
  AOI22_X1 U6928 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5943), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5859), .ZN(n5847) );
  OAI21_X1 U6929 ( .B1(n5848), .B2(n5952), .A(n5847), .ZN(n5849) );
  AOI211_X1 U6930 ( .C1(n5927), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5926), 
        .B(n5849), .ZN(n5852) );
  AOI22_X1 U6931 ( .A1(n5960), .A2(n5907), .B1(n5944), .B2(n5850), .ZN(n5851)
         );
  OAI211_X1 U6932 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5853), .A(n5852), .B(n5851), .ZN(U2809) );
  OAI22_X1 U6933 ( .A1(n6654), .A2(n5924), .B1(n5854), .B2(n5939), .ZN(n5855)
         );
  AOI211_X1 U6934 ( .C1(n5928), .C2(n5856), .A(n5926), .B(n5855), .ZN(n5861)
         );
  NAND2_X1 U6935 ( .A1(n6431), .A2(n5857), .ZN(n5858) );
  AOI22_X1 U6936 ( .A1(n5963), .A2(n5907), .B1(n5859), .B2(n5858), .ZN(n5860)
         );
  OAI211_X1 U6937 ( .C1(n5910), .C2(n5862), .A(n5861), .B(n5860), .ZN(U2810)
         );
  INV_X1 U6938 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5868) );
  AOI21_X1 U6939 ( .B1(n5865), .B2(n5864), .A(n5863), .ZN(n5893) );
  AOI22_X1 U6940 ( .A1(n5944), .A2(n5866), .B1(REIP_REG_13__SCAN_IN), .B2(
        n5893), .ZN(n5867) );
  OAI211_X1 U6941 ( .C1(n5939), .C2(n5868), .A(n5867), .B(n5887), .ZN(n5873)
         );
  OAI21_X1 U6942 ( .B1(REIP_REG_13__SCAN_IN), .B2(REIP_REG_12__SCAN_IN), .A(
        n5869), .ZN(n5870) );
  OAI22_X1 U6943 ( .A1(n5871), .A2(n5880), .B1(n5870), .B2(n5885), .ZN(n5872)
         );
  AOI211_X1 U6944 ( .C1(EBX_REG_13__SCAN_IN), .C2(n5943), .A(n5873), .B(n5872), 
        .ZN(n5874) );
  OAI21_X1 U6945 ( .B1(n5875), .B2(n5952), .A(n5874), .ZN(U2814) );
  AOI22_X1 U6946 ( .A1(EBX_REG_12__SCAN_IN), .A2(n5943), .B1(n5944), .B2(n6044), .ZN(n5876) );
  OAI211_X1 U6947 ( .C1(n5939), .C2(n5877), .A(n5876), .B(n5887), .ZN(n5878)
         );
  AOI21_X1 U6948 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5893), .A(n5878), .ZN(n5884) );
  OAI22_X1 U6949 ( .A1(n5881), .A2(n5880), .B1(n5879), .B2(n5952), .ZN(n5882)
         );
  INV_X1 U6950 ( .A(n5882), .ZN(n5883) );
  OAI211_X1 U6951 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5885), .A(n5884), .B(n5883), .ZN(U2815) );
  NAND3_X1 U6952 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n5886), .ZN(n5896) );
  OAI21_X1 U6953 ( .B1(n5939), .B2(n5888), .A(n5887), .ZN(n5892) );
  OAI22_X1 U6954 ( .A1(n5890), .A2(n5924), .B1(n5910), .B2(n5889), .ZN(n5891)
         );
  AOI211_X1 U6955 ( .C1(REIP_REG_11__SCAN_IN), .C2(n5893), .A(n5892), .B(n5891), .ZN(n5895) );
  AOI22_X1 U6956 ( .A1(n6008), .A2(n5907), .B1(n5928), .B2(n6006), .ZN(n5894)
         );
  OAI211_X1 U6957 ( .C1(REIP_REG_11__SCAN_IN), .C2(n5896), .A(n5895), .B(n5894), .ZN(U2816) );
  OAI22_X1 U6958 ( .A1(n5918), .A2(n6635), .B1(n5897), .B2(REIP_REG_6__SCAN_IN), .ZN(n5906) );
  INV_X1 U6959 ( .A(n5898), .ZN(n5901) );
  AOI21_X1 U6960 ( .B1(n5901), .B2(n5900), .A(n3631), .ZN(n6076) );
  OAI22_X1 U6961 ( .A1(n5954), .A2(n5924), .B1(n5902), .B2(n5939), .ZN(n5903)
         );
  AOI211_X1 U6962 ( .C1(n5944), .C2(n6076), .A(n5926), .B(n5903), .ZN(n5904)
         );
  INV_X1 U6963 ( .A(n5904), .ZN(n5905) );
  AOI211_X1 U6964 ( .C1(n5907), .C2(n6017), .A(n5906), .B(n5905), .ZN(n5908)
         );
  OAI21_X1 U6965 ( .B1(n6020), .B2(n5952), .A(n5908), .ZN(U2821) );
  NOR2_X1 U6966 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5909), .ZN(n5917) );
  OAI22_X1 U6967 ( .A1(n4852), .A2(n5939), .B1(n5910), .B2(n6090), .ZN(n5911)
         );
  AOI211_X1 U6968 ( .C1(n5943), .C2(EBX_REG_5__SCAN_IN), .A(n5926), .B(n5911), 
        .ZN(n5916) );
  INV_X1 U6969 ( .A(n5912), .ZN(n5914) );
  AOI22_X1 U6970 ( .A1(n5914), .A2(n5950), .B1(n5913), .B2(n5928), .ZN(n5915)
         );
  OAI211_X1 U6971 ( .C1(n5918), .C2(n5917), .A(n5916), .B(n5915), .ZN(U2822)
         );
  AOI21_X1 U6972 ( .B1(n5920), .B2(n5919), .A(n2989), .ZN(n6102) );
  AOI22_X1 U6973 ( .A1(n5944), .A2(n6102), .B1(n5922), .B2(n5921), .ZN(n5935)
         );
  INV_X1 U6974 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5958) );
  OAI22_X1 U6975 ( .A1(n5958), .A2(n5924), .B1(n6414), .B2(n5923), .ZN(n5925)
         );
  AOI211_X1 U6976 ( .C1(n5927), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5926), 
        .B(n5925), .ZN(n5934) );
  INV_X1 U6977 ( .A(n6029), .ZN(n5929) );
  AOI22_X1 U6978 ( .A1(n6026), .A2(n5950), .B1(n5929), .B2(n5928), .ZN(n5933)
         );
  OR3_X1 U6979 ( .A1(n5931), .A2(n5930), .A3(REIP_REG_4__SCAN_IN), .ZN(n5932)
         );
  NAND4_X1 U6980 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(U2823)
         );
  INV_X1 U6981 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6532) );
  NOR3_X1 U6982 ( .A1(n5937), .A2(n5936), .A3(n6532), .ZN(n5948) );
  AOI21_X1 U6983 ( .B1(n5938), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5947) );
  OAI22_X1 U6984 ( .A1(n5941), .A2(n4529), .B1(n5940), .B2(n5939), .ZN(n5942)
         );
  AOI21_X1 U6985 ( .B1(n5943), .B2(EBX_REG_2__SCAN_IN), .A(n5942), .ZN(n5946)
         );
  NAND2_X1 U6986 ( .A1(n5944), .A2(n6120), .ZN(n5945) );
  OAI211_X1 U6987 ( .C1(n5948), .C2(n5947), .A(n5946), .B(n5945), .ZN(n5949)
         );
  AOI21_X1 U6988 ( .B1(n6034), .B2(n5950), .A(n5949), .ZN(n5951) );
  OAI21_X1 U6989 ( .B1(n6038), .B2(n5952), .A(n5951), .ZN(U2825) );
  AOI22_X1 U6990 ( .A1(n6017), .A2(n5956), .B1(n5955), .B2(n6076), .ZN(n5953)
         );
  OAI21_X1 U6991 ( .B1(n5959), .B2(n5954), .A(n5953), .ZN(U2853) );
  AOI22_X1 U6992 ( .A1(n6026), .A2(n5956), .B1(n5955), .B2(n6102), .ZN(n5957)
         );
  OAI21_X1 U6993 ( .B1(n5959), .B2(n5958), .A(n5957), .ZN(U2855) );
  AOI22_X1 U6994 ( .A1(n5960), .A2(n5968), .B1(n5967), .B2(DATAI_18_), .ZN(
        n5962) );
  AOI22_X1 U6995 ( .A1(n5971), .A2(DATAI_2_), .B1(n5970), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U6996 ( .A1(n5962), .A2(n5961), .ZN(U2873) );
  AOI22_X1 U6997 ( .A1(n5963), .A2(n5968), .B1(n5967), .B2(DATAI_17_), .ZN(
        n5965) );
  AOI22_X1 U6998 ( .A1(n5971), .A2(DATAI_1_), .B1(n5970), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U6999 ( .A1(n5965), .A2(n5964), .ZN(U2874) );
  INV_X1 U7000 ( .A(n5966), .ZN(n5969) );
  AOI22_X1 U7001 ( .A1(n5969), .A2(n5968), .B1(n5967), .B2(DATAI_16_), .ZN(
        n5973) );
  AOI22_X1 U7002 ( .A1(n5971), .A2(DATAI_0_), .B1(n5970), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7003 ( .A1(n5973), .A2(n5972), .ZN(U2875) );
  AOI22_X1 U7004 ( .A1(n6486), .A2(LWORD_REG_15__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5975) );
  OAI21_X1 U7005 ( .B1(n5976), .B2(n6004), .A(n5975), .ZN(U2908) );
  AOI22_X1 U7006 ( .A1(n6486), .A2(LWORD_REG_14__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5977) );
  OAI21_X1 U7007 ( .B1(n5978), .B2(n6004), .A(n5977), .ZN(U2909) );
  AOI22_X1 U7008 ( .A1(n6486), .A2(LWORD_REG_13__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5979) );
  OAI21_X1 U7009 ( .B1(n5980), .B2(n6004), .A(n5979), .ZN(U2910) );
  AOI22_X1 U7010 ( .A1(n6486), .A2(LWORD_REG_12__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5981) );
  OAI21_X1 U7011 ( .B1(n5982), .B2(n6004), .A(n5981), .ZN(U2911) );
  AOI22_X1 U7012 ( .A1(DATAO_REG_11__SCAN_IN), .A2(n6002), .B1(
        LWORD_REG_11__SCAN_IN), .B2(n6001), .ZN(n5983) );
  OAI21_X1 U7013 ( .B1(n5984), .B2(n6004), .A(n5983), .ZN(U2912) );
  AOI22_X1 U7014 ( .A1(n6486), .A2(LWORD_REG_10__SCAN_IN), .B1(n5993), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5985) );
  OAI21_X1 U7015 ( .B1(n6579), .B2(n6004), .A(n5985), .ZN(U2913) );
  AOI22_X1 U7016 ( .A1(n6486), .A2(LWORD_REG_9__SCAN_IN), .B1(n5993), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5986) );
  OAI21_X1 U7017 ( .B1(n6526), .B2(n6004), .A(n5986), .ZN(U2914) );
  AOI22_X1 U7018 ( .A1(n6486), .A2(LWORD_REG_8__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5987) );
  OAI21_X1 U7019 ( .B1(n5988), .B2(n6004), .A(n5987), .ZN(U2915) );
  AOI22_X1 U7020 ( .A1(DATAO_REG_7__SCAN_IN), .A2(n6002), .B1(n6001), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n5989) );
  OAI21_X1 U7021 ( .B1(n4946), .B2(n6004), .A(n5989), .ZN(U2916) );
  AOI22_X1 U7022 ( .A1(n6486), .A2(LWORD_REG_6__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5990) );
  OAI21_X1 U7023 ( .B1(n4862), .B2(n6004), .A(n5990), .ZN(U2917) );
  AOI22_X1 U7024 ( .A1(n6486), .A2(LWORD_REG_5__SCAN_IN), .B1(n5993), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5991) );
  OAI21_X1 U7025 ( .B1(n5992), .B2(n6004), .A(n5991), .ZN(U2918) );
  AOI22_X1 U7026 ( .A1(n6486), .A2(LWORD_REG_4__SCAN_IN), .B1(n5993), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5994) );
  OAI21_X1 U7027 ( .B1(n5995), .B2(n6004), .A(n5994), .ZN(U2919) );
  AOI22_X1 U7028 ( .A1(DATAO_REG_3__SCAN_IN), .A2(n6002), .B1(n6001), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n5996) );
  OAI21_X1 U7029 ( .B1(n5997), .B2(n6004), .A(n5996), .ZN(U2920) );
  AOI22_X1 U7030 ( .A1(n6486), .A2(LWORD_REG_2__SCAN_IN), .B1(n6002), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5998) );
  OAI21_X1 U7031 ( .B1(n5999), .B2(n6004), .A(n5998), .ZN(U2921) );
  AOI22_X1 U7032 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6001), .B1(n6002), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6000) );
  OAI21_X1 U7033 ( .B1(n6542), .B2(n6004), .A(n6000), .ZN(U2922) );
  AOI22_X1 U7034 ( .A1(DATAO_REG_0__SCAN_IN), .A2(n6002), .B1(n6001), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n6003) );
  OAI21_X1 U7035 ( .B1(n6005), .B2(n6004), .A(n6003), .ZN(U2923) );
  AOI22_X1 U7036 ( .A1(n6101), .A2(REIP_REG_11__SCAN_IN), .B1(n6030), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6010) );
  AOI22_X1 U7037 ( .A1(n6008), .A2(n2963), .B1(n6007), .B2(n6006), .ZN(n6009)
         );
  OAI211_X1 U7038 ( .C1(n6012), .C2(n6011), .A(n6010), .B(n6009), .ZN(U2975)
         );
  AOI22_X1 U7039 ( .A1(n6101), .A2(REIP_REG_6__SCAN_IN), .B1(n6030), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6019) );
  OAI21_X1 U7040 ( .B1(n6015), .B2(n6014), .A(n6013), .ZN(n6016) );
  INV_X1 U7041 ( .A(n6016), .ZN(n6081) );
  AOI22_X1 U7042 ( .A1(n6081), .A2(n6035), .B1(n2963), .B2(n6017), .ZN(n6018)
         );
  OAI211_X1 U7043 ( .C1(n6039), .C2(n6020), .A(n6019), .B(n6018), .ZN(U2980)
         );
  AOI22_X1 U7044 ( .A1(n6101), .A2(REIP_REG_4__SCAN_IN), .B1(n6030), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7045 ( .B1(n6021), .B2(n6022), .A(n6023), .ZN(n6025) );
  INV_X1 U7046 ( .A(n6025), .ZN(n6103) );
  AOI22_X1 U7047 ( .A1(n6103), .A2(n6035), .B1(n6026), .B2(n2963), .ZN(n6027)
         );
  OAI211_X1 U7048 ( .C1(n6039), .C2(n6029), .A(n6028), .B(n6027), .ZN(U2982)
         );
  AOI22_X1 U7049 ( .A1(n6101), .A2(REIP_REG_2__SCAN_IN), .B1(n6030), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6037) );
  XOR2_X1 U7050 ( .A(n6031), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6033) );
  XNOR2_X1 U7051 ( .A(n6033), .B(n6032), .ZN(n6130) );
  AOI22_X1 U7052 ( .A1(n6130), .A2(n6035), .B1(n2963), .B2(n6034), .ZN(n6036)
         );
  OAI211_X1 U7053 ( .C1(n6039), .C2(n6038), .A(n6037), .B(n6036), .ZN(U2984)
         );
  AOI221_X1 U7054 ( .B1(n6097), .B2(n6042), .C1(n6041), .C2(n6042), .A(n6040), 
        .ZN(n6049) );
  AOI21_X1 U7055 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6043), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6048) );
  AOI22_X1 U7056 ( .A1(n6045), .A2(n6129), .B1(n6121), .B2(n6044), .ZN(n6047)
         );
  NAND2_X1 U7057 ( .A1(n6101), .A2(REIP_REG_12__SCAN_IN), .ZN(n6046) );
  OAI211_X1 U7058 ( .C1(n6049), .C2(n6048), .A(n6047), .B(n6046), .ZN(U3006)
         );
  AOI22_X1 U7059 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n3481), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6050), .ZN(n6057) );
  AOI21_X1 U7060 ( .B1(n6052), .B2(n6121), .A(n6051), .ZN(n6056) );
  AOI22_X1 U7061 ( .A1(n6054), .A2(n6129), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6053), .ZN(n6055) );
  OAI211_X1 U7062 ( .C1(n6058), .C2(n6057), .A(n6056), .B(n6055), .ZN(U3008)
         );
  AOI21_X1 U7063 ( .B1(n6060), .B2(n6121), .A(n6059), .ZN(n6065) );
  AOI21_X1 U7064 ( .B1(n6074), .B2(n6066), .A(n6061), .ZN(n6062) );
  AOI22_X1 U7065 ( .A1(n6063), .A2(n6129), .B1(n6070), .B2(n6062), .ZN(n6064)
         );
  OAI211_X1 U7066 ( .C1(n6075), .C2(n6066), .A(n6065), .B(n6064), .ZN(U3010)
         );
  AOI21_X1 U7067 ( .B1(n6068), .B2(n6121), .A(n6067), .ZN(n6073) );
  INV_X1 U7068 ( .A(n6069), .ZN(n6071) );
  AOI22_X1 U7069 ( .A1(n6071), .A2(n6129), .B1(n6070), .B2(n6074), .ZN(n6072)
         );
  OAI211_X1 U7070 ( .C1(n6075), .C2(n6074), .A(n6073), .B(n6072), .ZN(U3011)
         );
  AOI22_X1 U7071 ( .A1(n6076), .A2(n6121), .B1(n6101), .B2(REIP_REG_6__SCAN_IN), .ZN(n6083) );
  INV_X1 U7072 ( .A(n6098), .ZN(n6119) );
  AOI22_X1 U7073 ( .A1(n6078), .A2(n6119), .B1(n6116), .B2(n6077), .ZN(n6133)
         );
  OAI21_X1 U7074 ( .B1(n6080), .B2(n6079), .A(n6133), .ZN(n6085) );
  AOI22_X1 U7075 ( .A1(n6085), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .B1(n6081), 
        .B2(n6129), .ZN(n6082) );
  OAI211_X1 U7076 ( .C1(INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n6084), .A(n6083), 
        .B(n6082), .ZN(U3012) );
  OAI21_X1 U7077 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n6086), .A(n6085), 
        .ZN(n6095) );
  INV_X1 U7078 ( .A(n6087), .ZN(n6093) );
  NOR3_X1 U7079 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6088), .A3(n6126), 
        .ZN(n6092) );
  OAI22_X1 U7080 ( .A1(n6090), .A2(n6089), .B1(n4851), .B2(n6123), .ZN(n6091)
         );
  AOI211_X1 U7081 ( .C1(n6093), .C2(n6129), .A(n6092), .B(n6091), .ZN(n6094)
         );
  NAND2_X1 U7082 ( .A1(n6095), .A2(n6094), .ZN(U3013) );
  OAI211_X1 U7083 ( .C1(n6098), .C2(n6097), .A(n6096), .B(n6118), .ZN(n6115)
         );
  AOI22_X1 U7084 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n6100), .B1(
        INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n6099), .ZN(n6106) );
  AOI22_X1 U7085 ( .A1(n6102), .A2(n6121), .B1(n6101), .B2(REIP_REG_4__SCAN_IN), .ZN(n6105) );
  OAI21_X1 U7086 ( .B1(n6116), .B2(n6118), .A(n6133), .ZN(n6112) );
  AOI22_X1 U7087 ( .A1(n6112), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n6129), 
        .B2(n6103), .ZN(n6104) );
  OAI211_X1 U7088 ( .C1(n6115), .C2(n6106), .A(n6105), .B(n6104), .ZN(U3014)
         );
  INV_X1 U7089 ( .A(n6107), .ZN(n6108) );
  AOI21_X1 U7090 ( .B1(n6121), .B2(n6109), .A(n6108), .ZN(n6114) );
  INV_X1 U7091 ( .A(n6110), .ZN(n6111) );
  AOI22_X1 U7092 ( .A1(n6112), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6129), 
        .B2(n6111), .ZN(n6113) );
  OAI211_X1 U7093 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6115), .A(n6114), 
        .B(n6113), .ZN(U3015) );
  AOI221_X1 U7094 ( .B1(n6119), .B2(n6118), .C1(n6117), .C2(n6118), .A(n6116), 
        .ZN(n6125) );
  NAND2_X1 U7095 ( .A1(n6121), .A2(n6120), .ZN(n6122) );
  OAI21_X1 U7096 ( .B1(n6532), .B2(n6123), .A(n6122), .ZN(n6124) );
  NOR2_X1 U7097 ( .A1(n6125), .A2(n6124), .ZN(n6132) );
  NOR3_X1 U7098 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6127), .A3(n6126), 
        .ZN(n6128) );
  AOI21_X1 U7099 ( .B1(n6130), .B2(n6129), .A(n6128), .ZN(n6131) );
  OAI211_X1 U7100 ( .C1(n6133), .C2(n3355), .A(n6132), .B(n6131), .ZN(U3016)
         );
  NOR2_X1 U7101 ( .A1(n6355), .A2(n6134), .ZN(U3019) );
  NOR2_X1 U7102 ( .A1(n6273), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6158)
         );
  AOI22_X1 U7103 ( .A1(n6175), .A2(n6135), .B1(n6275), .B2(n6158), .ZN(n6145)
         );
  INV_X1 U7104 ( .A(n6141), .ZN(n6140) );
  OAI21_X1 U7105 ( .B1(n6136), .B2(n6276), .A(n6284), .ZN(n6143) );
  INV_X1 U7106 ( .A(n6143), .ZN(n6138) );
  AOI21_X1 U7107 ( .B1(n6137), .B2(n6278), .A(n6158), .ZN(n6142) );
  NAND2_X1 U7108 ( .A1(n6138), .A2(n6142), .ZN(n6139) );
  OAI211_X1 U7109 ( .C1(n6284), .C2(n6140), .A(n6139), .B(n6281), .ZN(n6161)
         );
  OAI22_X1 U7110 ( .A1(n6143), .A2(n6142), .B1(n6141), .B2(n6285), .ZN(n6160)
         );
  AOI22_X1 U7111 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6161), .B1(n6289), 
        .B2(n6160), .ZN(n6144) );
  OAI211_X1 U7112 ( .C1(n6178), .C2(n6174), .A(n6145), .B(n6144), .ZN(U3044)
         );
  AOI22_X1 U7113 ( .A1(n6293), .A2(n6159), .B1(n6294), .B2(n6158), .ZN(n6147)
         );
  AOI22_X1 U7114 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6161), .B1(n6295), 
        .B2(n6160), .ZN(n6146) );
  OAI211_X1 U7115 ( .C1(n6164), .C2(n6298), .A(n6147), .B(n6146), .ZN(U3045)
         );
  AOI22_X1 U7116 ( .A1(n6299), .A2(n6159), .B1(n6300), .B2(n6158), .ZN(n6149)
         );
  AOI22_X1 U7117 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6161), .B1(n6301), 
        .B2(n6160), .ZN(n6148) );
  OAI211_X1 U7118 ( .C1(n6164), .C2(n6304), .A(n6149), .B(n6148), .ZN(U3046)
         );
  AOI22_X1 U7119 ( .A1(n6251), .A2(n6159), .B1(n6306), .B2(n6158), .ZN(n6151)
         );
  AOI22_X1 U7120 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6161), .B1(n6307), 
        .B2(n6160), .ZN(n6150) );
  OAI211_X1 U7121 ( .C1(n6164), .C2(n6254), .A(n6151), .B(n6150), .ZN(U3047)
         );
  AOI22_X1 U7122 ( .A1(n6255), .A2(n6159), .B1(n6312), .B2(n6158), .ZN(n6153)
         );
  AOI22_X1 U7123 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6161), .B1(n6313), 
        .B2(n6160), .ZN(n6152) );
  OAI211_X1 U7124 ( .C1(n6164), .C2(n6258), .A(n6153), .B(n6152), .ZN(U3048)
         );
  AOI22_X1 U7125 ( .A1(n6317), .A2(n6159), .B1(n6319), .B2(n6158), .ZN(n6155)
         );
  AOI22_X1 U7126 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6161), .B1(n6320), 
        .B2(n6160), .ZN(n6154) );
  OAI211_X1 U7127 ( .C1(n6164), .C2(n6324), .A(n6155), .B(n6154), .ZN(U3049)
         );
  AOI22_X1 U7128 ( .A1(n6261), .A2(n6159), .B1(n6326), .B2(n6158), .ZN(n6157)
         );
  AOI22_X1 U7129 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6161), .B1(n6327), 
        .B2(n6160), .ZN(n6156) );
  OAI211_X1 U7130 ( .C1(n6164), .C2(n6264), .A(n6157), .B(n6156), .ZN(U3050)
         );
  AOI22_X1 U7131 ( .A1(n6268), .A2(n6159), .B1(n6334), .B2(n6158), .ZN(n6163)
         );
  AOI22_X1 U7132 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6161), .B1(n6502), 
        .B2(n6160), .ZN(n6162) );
  OAI211_X1 U7133 ( .C1(n6164), .C2(n6498), .A(n6163), .B(n6162), .ZN(U3051)
         );
  INV_X1 U7134 ( .A(n6165), .ZN(n6168) );
  AOI22_X1 U7135 ( .A1(n6312), .A2(n6169), .B1(n6313), .B2(n6168), .ZN(n6167)
         );
  AOI22_X1 U7136 ( .A1(n6171), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6255), 
        .B2(n6170), .ZN(n6166) );
  OAI211_X1 U7137 ( .C1(n6258), .C2(n6174), .A(n6167), .B(n6166), .ZN(U3056)
         );
  AOI22_X1 U7138 ( .A1(n6326), .A2(n6169), .B1(n6327), .B2(n6168), .ZN(n6173)
         );
  AOI22_X1 U7139 ( .A1(n6171), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6261), 
        .B2(n6170), .ZN(n6172) );
  OAI211_X1 U7140 ( .C1(n6264), .C2(n6174), .A(n6173), .B(n6172), .ZN(U3058)
         );
  AOI22_X1 U7141 ( .A1(n6275), .A2(n6184), .B1(n6289), .B2(n6183), .ZN(n6177)
         );
  AOI22_X1 U7142 ( .A1(n6186), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6175), 
        .B2(n6185), .ZN(n6176) );
  OAI211_X1 U7143 ( .C1(n6178), .C2(n6227), .A(n6177), .B(n6176), .ZN(U3068)
         );
  AOI22_X1 U7144 ( .A1(n6294), .A2(n6184), .B1(n6295), .B2(n6183), .ZN(n6180)
         );
  AOI22_X1 U7145 ( .A1(n6186), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6205), 
        .B2(n6185), .ZN(n6179) );
  OAI211_X1 U7146 ( .C1(n6208), .C2(n6227), .A(n6180), .B(n6179), .ZN(U3069)
         );
  AOI22_X1 U7147 ( .A1(n6300), .A2(n6184), .B1(n6301), .B2(n6183), .ZN(n6182)
         );
  AOI22_X1 U7148 ( .A1(n6186), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6210), 
        .B2(n6185), .ZN(n6181) );
  OAI211_X1 U7149 ( .C1(n6213), .C2(n6227), .A(n6182), .B(n6181), .ZN(U3070)
         );
  AOI22_X1 U7150 ( .A1(n6306), .A2(n6184), .B1(n6307), .B2(n6183), .ZN(n6188)
         );
  AOI22_X1 U7151 ( .A1(n6186), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6305), 
        .B2(n6185), .ZN(n6187) );
  OAI211_X1 U7152 ( .C1(n6310), .C2(n6227), .A(n6188), .B(n6187), .ZN(U3071)
         );
  INV_X1 U7153 ( .A(n6195), .ZN(n6222) );
  AOI22_X1 U7154 ( .A1(n6275), .A2(n6222), .B1(n6274), .B2(n6236), .ZN(n6204)
         );
  INV_X1 U7155 ( .A(n6191), .ZN(n6193) );
  OAI21_X1 U7156 ( .B1(n6193), .B2(n6192), .A(n6284), .ZN(n6201) );
  INV_X1 U7157 ( .A(n6201), .ZN(n6197) );
  NAND3_X1 U7158 ( .A1(n6194), .A2(n6230), .A3(n6278), .ZN(n6196) );
  AND2_X1 U7159 ( .A1(n6196), .A2(n6195), .ZN(n6202) );
  NAND2_X1 U7160 ( .A1(n6197), .A2(n6202), .ZN(n6198) );
  OAI211_X1 U7161 ( .C1(n6199), .C2(n6284), .A(n6281), .B(n6198), .ZN(n6224)
         );
  OAI22_X1 U7162 ( .A1(n6202), .A2(n6201), .B1(n6285), .B2(n6200), .ZN(n6223)
         );
  AOI22_X1 U7163 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6224), .B1(n6289), 
        .B2(n6223), .ZN(n6203) );
  OAI211_X1 U7164 ( .C1(n6292), .C2(n6227), .A(n6204), .B(n6203), .ZN(U3076)
         );
  AOI22_X1 U7165 ( .A1(n6294), .A2(n6222), .B1(n6205), .B2(n6209), .ZN(n6207)
         );
  AOI22_X1 U7166 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6224), .B1(n6295), 
        .B2(n6223), .ZN(n6206) );
  OAI211_X1 U7167 ( .C1(n6208), .C2(n6272), .A(n6207), .B(n6206), .ZN(U3077)
         );
  AOI22_X1 U7168 ( .A1(n6300), .A2(n6222), .B1(n6210), .B2(n6209), .ZN(n6212)
         );
  AOI22_X1 U7169 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6224), .B1(n6301), 
        .B2(n6223), .ZN(n6211) );
  OAI211_X1 U7170 ( .C1(n6213), .C2(n6272), .A(n6212), .B(n6211), .ZN(U3078)
         );
  AOI22_X1 U7171 ( .A1(n6306), .A2(n6222), .B1(n6251), .B2(n6236), .ZN(n6215)
         );
  AOI22_X1 U7172 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6224), .B1(n6307), 
        .B2(n6223), .ZN(n6214) );
  OAI211_X1 U7173 ( .C1(n6254), .C2(n6227), .A(n6215), .B(n6214), .ZN(U3079)
         );
  AOI22_X1 U7174 ( .A1(n6312), .A2(n6222), .B1(n6255), .B2(n6236), .ZN(n6217)
         );
  AOI22_X1 U7175 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6224), .B1(n6313), 
        .B2(n6223), .ZN(n6216) );
  OAI211_X1 U7176 ( .C1(n6258), .C2(n6227), .A(n6217), .B(n6216), .ZN(U3080)
         );
  AOI22_X1 U7177 ( .A1(n6319), .A2(n6222), .B1(n6317), .B2(n6236), .ZN(n6219)
         );
  AOI22_X1 U7178 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6224), .B1(n6320), 
        .B2(n6223), .ZN(n6218) );
  OAI211_X1 U7179 ( .C1(n6324), .C2(n6227), .A(n6219), .B(n6218), .ZN(U3081)
         );
  AOI22_X1 U7180 ( .A1(n6326), .A2(n6222), .B1(n6261), .B2(n6236), .ZN(n6221)
         );
  AOI22_X1 U7181 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6224), .B1(n6327), 
        .B2(n6223), .ZN(n6220) );
  OAI211_X1 U7182 ( .C1(n6264), .C2(n6227), .A(n6221), .B(n6220), .ZN(U3082)
         );
  AOI22_X1 U7183 ( .A1(n6334), .A2(n6222), .B1(n6268), .B2(n6236), .ZN(n6226)
         );
  AOI22_X1 U7184 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6224), .B1(n6502), 
        .B2(n6223), .ZN(n6225) );
  OAI211_X1 U7185 ( .C1(n6498), .C2(n6227), .A(n6226), .B(n6225), .ZN(U3083)
         );
  NOR2_X1 U7186 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6228), .ZN(n6266)
         );
  NOR2_X1 U7187 ( .A1(n6230), .A2(n6229), .ZN(n6243) );
  INV_X1 U7188 ( .A(n6243), .ZN(n6234) );
  INV_X1 U7189 ( .A(n6231), .ZN(n6232) );
  OAI22_X1 U7190 ( .A1(n6234), .A2(n6235), .B1(n6233), .B2(n6232), .ZN(n6265)
         );
  AOI22_X1 U7191 ( .A1(n6275), .A2(n6266), .B1(n6289), .B2(n6265), .ZN(n6246)
         );
  NOR3_X1 U7192 ( .A1(n6267), .A2(n6236), .A3(n6235), .ZN(n6238) );
  NOR2_X1 U7193 ( .A1(n6238), .A2(n6237), .ZN(n6244) );
  INV_X1 U7194 ( .A(n6266), .ZN(n6241) );
  AOI211_X1 U7195 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6241), .A(n6240), .B(
        n6239), .ZN(n6242) );
  OAI21_X1 U7196 ( .B1(n6244), .B2(n6243), .A(n6242), .ZN(n6269) );
  AOI22_X1 U7197 ( .A1(n6269), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6274), 
        .B2(n6267), .ZN(n6245) );
  OAI211_X1 U7198 ( .C1(n6292), .C2(n6272), .A(n6246), .B(n6245), .ZN(U3084)
         );
  AOI22_X1 U7199 ( .A1(n6294), .A2(n6266), .B1(n6295), .B2(n6265), .ZN(n6248)
         );
  AOI22_X1 U7200 ( .A1(n6269), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6293), 
        .B2(n6267), .ZN(n6247) );
  OAI211_X1 U7201 ( .C1(n6298), .C2(n6272), .A(n6248), .B(n6247), .ZN(U3085)
         );
  AOI22_X1 U7202 ( .A1(n6300), .A2(n6266), .B1(n6301), .B2(n6265), .ZN(n6250)
         );
  AOI22_X1 U7203 ( .A1(n6269), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6299), 
        .B2(n6267), .ZN(n6249) );
  OAI211_X1 U7204 ( .C1(n6304), .C2(n6272), .A(n6250), .B(n6249), .ZN(U3086)
         );
  AOI22_X1 U7205 ( .A1(n6306), .A2(n6266), .B1(n6307), .B2(n6265), .ZN(n6253)
         );
  AOI22_X1 U7206 ( .A1(n6269), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6251), 
        .B2(n6267), .ZN(n6252) );
  OAI211_X1 U7207 ( .C1(n6254), .C2(n6272), .A(n6253), .B(n6252), .ZN(U3087)
         );
  AOI22_X1 U7208 ( .A1(n6312), .A2(n6266), .B1(n6313), .B2(n6265), .ZN(n6257)
         );
  AOI22_X1 U7209 ( .A1(n6269), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6255), 
        .B2(n6267), .ZN(n6256) );
  OAI211_X1 U7210 ( .C1(n6258), .C2(n6272), .A(n6257), .B(n6256), .ZN(U3088)
         );
  AOI22_X1 U7211 ( .A1(n6319), .A2(n6266), .B1(n6320), .B2(n6265), .ZN(n6260)
         );
  AOI22_X1 U7212 ( .A1(n6269), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6317), 
        .B2(n6267), .ZN(n6259) );
  OAI211_X1 U7213 ( .C1(n6324), .C2(n6272), .A(n6260), .B(n6259), .ZN(U3089)
         );
  AOI22_X1 U7214 ( .A1(n6326), .A2(n6266), .B1(n6327), .B2(n6265), .ZN(n6263)
         );
  AOI22_X1 U7215 ( .A1(n6269), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6261), 
        .B2(n6267), .ZN(n6262) );
  OAI211_X1 U7216 ( .C1(n6264), .C2(n6272), .A(n6263), .B(n6262), .ZN(U3090)
         );
  AOI22_X1 U7217 ( .A1(n6334), .A2(n6266), .B1(n6502), .B2(n6265), .ZN(n6271)
         );
  AOI22_X1 U7218 ( .A1(n6269), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6268), 
        .B2(n6267), .ZN(n6270) );
  OAI211_X1 U7219 ( .C1(n6498), .C2(n6272), .A(n6271), .B(n6270), .ZN(U3091)
         );
  NOR2_X1 U7220 ( .A1(n6358), .A2(n6273), .ZN(n6333) );
  AOI22_X1 U7221 ( .A1(n6275), .A2(n6333), .B1(n6318), .B2(n6274), .ZN(n6291)
         );
  INV_X1 U7222 ( .A(n6286), .ZN(n6283) );
  OAI21_X1 U7223 ( .B1(n6277), .B2(n6276), .A(n6284), .ZN(n6288) );
  INV_X1 U7224 ( .A(n6288), .ZN(n6280) );
  AOI21_X1 U7225 ( .B1(n6279), .B2(n6278), .A(n6333), .ZN(n6287) );
  NAND2_X1 U7226 ( .A1(n6280), .A2(n6287), .ZN(n6282) );
  OAI211_X1 U7227 ( .C1(n6284), .C2(n6283), .A(n6282), .B(n6281), .ZN(n6336)
         );
  OAI22_X1 U7228 ( .A1(n6288), .A2(n6287), .B1(n6286), .B2(n6285), .ZN(n6335)
         );
  AOI22_X1 U7229 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6336), .B1(n6289), 
        .B2(n6335), .ZN(n6290) );
  OAI211_X1 U7230 ( .C1(n6292), .C2(n6323), .A(n6291), .B(n6290), .ZN(U3108)
         );
  AOI22_X1 U7231 ( .A1(n6294), .A2(n6333), .B1(n6318), .B2(n6293), .ZN(n6297)
         );
  AOI22_X1 U7232 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6336), .B1(n6295), 
        .B2(n6335), .ZN(n6296) );
  OAI211_X1 U7233 ( .C1(n6298), .C2(n6323), .A(n6297), .B(n6296), .ZN(U3109)
         );
  AOI22_X1 U7234 ( .A1(n6300), .A2(n6333), .B1(n6318), .B2(n6299), .ZN(n6303)
         );
  AOI22_X1 U7235 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6336), .B1(n6301), 
        .B2(n6335), .ZN(n6302) );
  OAI211_X1 U7236 ( .C1(n6304), .C2(n6323), .A(n6303), .B(n6302), .ZN(U3110)
         );
  INV_X1 U7237 ( .A(n6323), .ZN(n6332) );
  AOI22_X1 U7238 ( .A1(n6306), .A2(n6333), .B1(n6332), .B2(n6305), .ZN(n6309)
         );
  AOI22_X1 U7239 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6336), .B1(n6307), 
        .B2(n6335), .ZN(n6308) );
  OAI211_X1 U7240 ( .C1(n6310), .C2(n6339), .A(n6309), .B(n6308), .ZN(U3111)
         );
  AOI22_X1 U7241 ( .A1(n6312), .A2(n6333), .B1(n6332), .B2(n6311), .ZN(n6315)
         );
  AOI22_X1 U7242 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6336), .B1(n6313), 
        .B2(n6335), .ZN(n6314) );
  OAI211_X1 U7243 ( .C1(n6316), .C2(n6339), .A(n6315), .B(n6314), .ZN(U3112)
         );
  AOI22_X1 U7244 ( .A1(n6319), .A2(n6333), .B1(n6318), .B2(n6317), .ZN(n6322)
         );
  AOI22_X1 U7245 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6336), .B1(n6320), 
        .B2(n6335), .ZN(n6321) );
  OAI211_X1 U7246 ( .C1(n6324), .C2(n6323), .A(n6322), .B(n6321), .ZN(U3113)
         );
  AOI22_X1 U7247 ( .A1(n6326), .A2(n6333), .B1(n6332), .B2(n6325), .ZN(n6329)
         );
  AOI22_X1 U7248 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6336), .B1(n6327), 
        .B2(n6335), .ZN(n6328) );
  OAI211_X1 U7249 ( .C1(n6330), .C2(n6339), .A(n6329), .B(n6328), .ZN(U3114)
         );
  AOI22_X1 U7250 ( .A1(n6334), .A2(n6333), .B1(n6332), .B2(n6331), .ZN(n6338)
         );
  AOI22_X1 U7251 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6336), .B1(n6502), 
        .B2(n6335), .ZN(n6337) );
  OAI211_X1 U7252 ( .C1(n6497), .C2(n6339), .A(n6338), .B(n6337), .ZN(U3115)
         );
  INV_X1 U7253 ( .A(n6357), .ZN(n6354) );
  AND3_X1 U7254 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6341), .A3(n6340), 
        .ZN(n6347) );
  INV_X1 U7255 ( .A(n6347), .ZN(n6344) );
  OAI211_X1 U7256 ( .C1(n6345), .C2(n6344), .A(n6343), .B(n6342), .ZN(n6346)
         );
  OAI21_X1 U7257 ( .B1(n6347), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6346), 
        .ZN(n6352) );
  INV_X1 U7258 ( .A(n6352), .ZN(n6349) );
  OAI21_X1 U7259 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6349), .A(n6348), 
        .ZN(n6350) );
  OAI21_X1 U7260 ( .B1(n6352), .B2(n6351), .A(n6350), .ZN(n6353) );
  OAI21_X1 U7261 ( .B1(n6354), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6353), 
        .ZN(n6356) );
  OAI211_X1 U7262 ( .C1(n6358), .C2(n6357), .A(n6356), .B(n6355), .ZN(n6368)
         );
  INV_X1 U7263 ( .A(n6359), .ZN(n6367) );
  OR2_X1 U7264 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6363) );
  INV_X1 U7265 ( .A(n6360), .ZN(n6362) );
  AOI211_X1 U7266 ( .C1(n6364), .C2(n6363), .A(n6362), .B(n6361), .ZN(n6365)
         );
  AND4_X1 U7267 ( .A1(n6368), .A2(n6367), .A3(n6366), .A4(n6365), .ZN(n6382)
         );
  OR2_X1 U7268 ( .A1(n6370), .A2(n6369), .ZN(n6373) );
  AOI21_X1 U7269 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6371) );
  INV_X1 U7270 ( .A(n6371), .ZN(n6372) );
  AND3_X1 U7271 ( .A1(n6373), .A2(STATE2_REG_2__SCAN_IN), .A3(n6372), .ZN(
        n6377) );
  OAI221_X1 U7272 ( .B1(n6379), .B2(n6382), .C1(n6379), .C2(n6374), .A(n6377), 
        .ZN(n6465) );
  OAI21_X1 U7273 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6485), .A(n6465), .ZN(
        n6383) );
  AOI221_X1 U7274 ( .B1(n6376), .B2(STATE2_REG_0__SCAN_IN), .C1(n6383), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6375), .ZN(n6381) );
  INV_X1 U7275 ( .A(n6377), .ZN(n6378) );
  OAI211_X1 U7276 ( .C1(n6390), .C2(n6467), .A(n6379), .B(n6378), .ZN(n6380)
         );
  OAI211_X1 U7277 ( .C1(n6382), .C2(n6384), .A(n6381), .B(n6380), .ZN(U3148)
         );
  OAI211_X1 U7278 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6383), .ZN(n6389) );
  OAI21_X1 U7279 ( .B1(READY_N), .B2(n6385), .A(n6384), .ZN(n6387) );
  AOI21_X1 U7280 ( .B1(n6387), .B2(n6465), .A(n6386), .ZN(n6388) );
  NAND2_X1 U7281 ( .A1(n6389), .A2(n6388), .ZN(U3149) );
  INV_X1 U7282 ( .A(n6390), .ZN(n6489) );
  OAI221_X1 U7283 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6485), .A(n6462), .ZN(n6392) );
  OAI21_X1 U7284 ( .B1(n6489), .B2(n6392), .A(n6391), .ZN(U3150) );
  INV_X1 U7285 ( .A(n6461), .ZN(n6457) );
  AND2_X1 U7286 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6457), .ZN(U3151) );
  AND2_X1 U7287 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6457), .ZN(U3152) );
  AND2_X1 U7288 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6457), .ZN(U3153) );
  AND2_X1 U7289 ( .A1(n6457), .A2(DATAWIDTH_REG_28__SCAN_IN), .ZN(U3154) );
  INV_X1 U7290 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6577) );
  NOR2_X1 U7291 ( .A1(n6461), .A2(n6577), .ZN(U3155) );
  AND2_X1 U7292 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6457), .ZN(U3156) );
  AND2_X1 U7293 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6457), .ZN(U3157) );
  AND2_X1 U7294 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6457), .ZN(U3158) );
  AND2_X1 U7295 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6457), .ZN(U3159) );
  AND2_X1 U7296 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6457), .ZN(U3160) );
  AND2_X1 U7297 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6457), .ZN(U3161) );
  AND2_X1 U7298 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6457), .ZN(U3162) );
  AND2_X1 U7299 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6457), .ZN(U3163) );
  AND2_X1 U7300 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6457), .ZN(U3164) );
  AND2_X1 U7301 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6457), .ZN(U3165) );
  AND2_X1 U7302 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6457), .ZN(U3166) );
  AND2_X1 U7303 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6457), .ZN(U3167) );
  AND2_X1 U7304 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6457), .ZN(U3168) );
  AND2_X1 U7305 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6457), .ZN(U3169) );
  AND2_X1 U7306 ( .A1(n6457), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U7307 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6457), .ZN(U3171) );
  AND2_X1 U7308 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6457), .ZN(U3172) );
  AND2_X1 U7309 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6457), .ZN(U3173) );
  AND2_X1 U7310 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6457), .ZN(U3174) );
  AND2_X1 U7311 ( .A1(n6457), .A2(DATAWIDTH_REG_7__SCAN_IN), .ZN(U3175) );
  AND2_X1 U7312 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6457), .ZN(U3176) );
  AND2_X1 U7313 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6457), .ZN(U3177) );
  AND2_X1 U7314 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6457), .ZN(U3178) );
  AND2_X1 U7315 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6457), .ZN(U3179) );
  AND2_X1 U7316 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6457), .ZN(U3180) );
  NOR2_X1 U7317 ( .A1(n6409), .A2(n6399), .ZN(n6400) );
  AOI22_X1 U7318 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6408) );
  AND2_X1 U7319 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6396) );
  INV_X1 U7320 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6394) );
  INV_X1 U7321 ( .A(NA_N), .ZN(n6401) );
  AOI221_X1 U7322 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6401), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6405) );
  AOI221_X1 U7323 ( .B1(n6396), .B2(n6448), .C1(n6394), .C2(n6448), .A(n6405), 
        .ZN(n6393) );
  OAI21_X1 U7324 ( .B1(n6400), .B2(n6408), .A(n6393), .ZN(U3181) );
  NOR2_X1 U7325 ( .A1(n6403), .A2(n6394), .ZN(n6402) );
  NAND2_X1 U7326 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6395) );
  OAI21_X1 U7327 ( .B1(n6402), .B2(n6396), .A(n6395), .ZN(n6397) );
  OAI211_X1 U7328 ( .C1(n6399), .C2(n6485), .A(n6398), .B(n6397), .ZN(U3182)
         );
  AOI21_X1 U7329 ( .B1(n6402), .B2(n6401), .A(n6400), .ZN(n6407) );
  AOI221_X1 U7330 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6485), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6404) );
  AOI221_X1 U7331 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6404), .C2(HOLD), .A(n6403), .ZN(n6406) );
  OAI22_X1 U7332 ( .A1(n6408), .A2(n6407), .B1(n6406), .B2(n6405), .ZN(U3183)
         );
  NAND2_X1 U7333 ( .A1(n6494), .A2(n6409), .ZN(n6455) );
  NOR2_X2 U7334 ( .A1(n6409), .A2(n6448), .ZN(n6449) );
  AOI22_X1 U7335 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6482), .ZN(n6410) );
  OAI21_X1 U7336 ( .B1(n6532), .B2(n6455), .A(n6410), .ZN(U3184) );
  INV_X1 U7337 ( .A(n6449), .ZN(n6451) );
  INV_X1 U7338 ( .A(n6455), .ZN(n6444) );
  AOI22_X1 U7339 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6482), .ZN(n6411) );
  OAI21_X1 U7340 ( .B1(n6532), .B2(n6451), .A(n6411), .ZN(U3185) );
  AOI22_X1 U7341 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6482), .ZN(n6412) );
  OAI21_X1 U7342 ( .B1(n6414), .B2(n6455), .A(n6412), .ZN(U3186) );
  AOI22_X1 U7343 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6482), .ZN(n6413) );
  OAI21_X1 U7344 ( .B1(n6414), .B2(n6451), .A(n6413), .ZN(U3187) );
  AOI22_X1 U7345 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6482), .ZN(n6415) );
  OAI21_X1 U7346 ( .B1(n6635), .B2(n6455), .A(n6415), .ZN(U3188) );
  INV_X1 U7347 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6416) );
  OAI222_X1 U7348 ( .A1(n6455), .A2(n4866), .B1(n6416), .B2(n6494), .C1(n6635), 
        .C2(n6451), .ZN(U3189) );
  AOI22_X1 U7349 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6482), .ZN(n6417) );
  OAI21_X1 U7350 ( .B1(n4866), .B2(n6451), .A(n6417), .ZN(U3190) );
  AOI22_X1 U7351 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6482), .ZN(n6418) );
  OAI21_X1 U7352 ( .B1(n6420), .B2(n6455), .A(n6418), .ZN(U3191) );
  AOI22_X1 U7353 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6448), .ZN(n6419) );
  OAI21_X1 U7354 ( .B1(n6420), .B2(n6451), .A(n6419), .ZN(U3192) );
  AOI22_X1 U7355 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6482), .ZN(n6421) );
  OAI21_X1 U7356 ( .B1(n5161), .B2(n6451), .A(n6421), .ZN(U3193) );
  AOI22_X1 U7357 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6482), .ZN(n6422) );
  OAI21_X1 U7358 ( .B1(n5189), .B2(n6455), .A(n6422), .ZN(U3194) );
  AOI22_X1 U7359 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6482), .ZN(n6423) );
  OAI21_X1 U7360 ( .B1(n5189), .B2(n6451), .A(n6423), .ZN(U3195) );
  AOI22_X1 U7361 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6482), .ZN(n6424) );
  OAI21_X1 U7362 ( .B1(n6425), .B2(n6455), .A(n6424), .ZN(U3196) );
  AOI22_X1 U7363 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6482), .ZN(n6426) );
  OAI21_X1 U7364 ( .B1(n6427), .B2(n6455), .A(n6426), .ZN(U3197) );
  AOI22_X1 U7365 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6482), .ZN(n6428) );
  OAI21_X1 U7366 ( .B1(n6574), .B2(n6455), .A(n6428), .ZN(U3198) );
  AOI22_X1 U7367 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6482), .ZN(n6429) );
  OAI21_X1 U7368 ( .B1(n6431), .B2(n6455), .A(n6429), .ZN(U3199) );
  AOI22_X1 U7369 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6482), .ZN(n6430) );
  OAI21_X1 U7370 ( .B1(n6431), .B2(n6451), .A(n6430), .ZN(U3200) );
  INV_X1 U7371 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6433) );
  AOI22_X1 U7372 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6482), .ZN(n6432) );
  OAI21_X1 U7373 ( .B1(n6433), .B2(n6451), .A(n6432), .ZN(U3201) );
  AOI22_X1 U7374 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6482), .ZN(n6434) );
  OAI21_X1 U7375 ( .B1(n5554), .B2(n6455), .A(n6434), .ZN(U3202) );
  AOI22_X1 U7376 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6448), .ZN(n6435) );
  OAI21_X1 U7377 ( .B1(n6561), .B2(n6455), .A(n6435), .ZN(U3203) );
  AOI22_X1 U7378 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6448), .ZN(n6436) );
  OAI21_X1 U7379 ( .B1(n5543), .B2(n6455), .A(n6436), .ZN(U3204) );
  AOI22_X1 U7380 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6448), .ZN(n6437) );
  OAI21_X1 U7381 ( .B1(n5543), .B2(n6451), .A(n6437), .ZN(U3205) );
  AOI22_X1 U7382 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6482), .ZN(n6438) );
  OAI21_X1 U7383 ( .B1(n6439), .B2(n6455), .A(n6438), .ZN(U3206) );
  AOI22_X1 U7384 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6448), .ZN(n6440) );
  OAI21_X1 U7385 ( .B1(n5516), .B2(n6455), .A(n6440), .ZN(U3207) );
  AOI22_X1 U7386 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6448), .ZN(n6441) );
  OAI21_X1 U7387 ( .B1(n6443), .B2(n6455), .A(n6441), .ZN(U3208) );
  AOI22_X1 U7388 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6448), .ZN(n6442) );
  OAI21_X1 U7389 ( .B1(n6443), .B2(n6451), .A(n6442), .ZN(U3209) );
  AOI22_X1 U7390 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6444), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6448), .ZN(n6445) );
  OAI21_X1 U7391 ( .B1(n4313), .B2(n6451), .A(n6445), .ZN(U3210) );
  AOI22_X1 U7392 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6448), .ZN(n6446) );
  OAI21_X1 U7393 ( .B1(n6447), .B2(n6455), .A(n6446), .ZN(U3211) );
  AOI22_X1 U7394 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6449), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6448), .ZN(n6450) );
  OAI21_X1 U7395 ( .B1(n6452), .B2(n6455), .A(n6450), .ZN(U3212) );
  INV_X1 U7396 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6453) );
  OAI222_X1 U7397 ( .A1(n6455), .A2(n6454), .B1(n6453), .B2(n6494), .C1(n6452), 
        .C2(n6451), .ZN(U3213) );
  MUX2_X1 U7398 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6494), .Z(U3445) );
  MUX2_X1 U7399 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6494), .Z(U3446) );
  MUX2_X1 U7400 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6494), .Z(U3447) );
  MUX2_X1 U7401 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6494), .Z(U3448) );
  INV_X1 U7402 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6458) );
  INV_X1 U7403 ( .A(n6459), .ZN(n6456) );
  AOI21_X1 U7404 ( .B1(n6458), .B2(n6457), .A(n6456), .ZN(U3451) );
  OAI21_X1 U7405 ( .B1(n6461), .B2(n6460), .A(n6459), .ZN(U3452) );
  OAI211_X1 U7406 ( .C1(n6465), .C2(n6464), .A(n6463), .B(n6462), .ZN(U3453)
         );
  INV_X1 U7407 ( .A(n6466), .ZN(n6470) );
  OAI22_X1 U7408 ( .A1(n6470), .A2(n6469), .B1(n6468), .B2(n6467), .ZN(n6472)
         );
  MUX2_X1 U7409 ( .A(n6472), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6471), 
        .Z(U3456) );
  AOI21_X1 U7410 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6473) );
  AOI22_X1 U7411 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6473), .B2(n6573), .ZN(n6475) );
  INV_X1 U7412 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6474) );
  AOI22_X1 U7413 ( .A1(n6476), .A2(n6475), .B1(n6474), .B2(n6479), .ZN(U3468)
         );
  INV_X1 U7414 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6480) );
  NOR2_X1 U7415 ( .A1(n6479), .A2(REIP_REG_1__SCAN_IN), .ZN(n6477) );
  AOI22_X1 U7416 ( .A1(n6480), .A2(n6479), .B1(n6478), .B2(n6477), .ZN(U3469)
         );
  NAND2_X1 U7417 ( .A1(n6482), .A2(W_R_N_REG_SCAN_IN), .ZN(n6481) );
  OAI21_X1 U7418 ( .B1(n6482), .B2(READREQUEST_REG_SCAN_IN), .A(n6481), .ZN(
        U3470) );
  AOI211_X1 U7419 ( .C1(n6486), .C2(n6485), .A(n6484), .B(n6483), .ZN(n6493)
         );
  OAI211_X1 U7420 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6488), .A(n6487), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6490) );
  AOI21_X1 U7421 ( .B1(n6490), .B2(STATE2_REG_0__SCAN_IN), .A(n6489), .ZN(
        n6492) );
  NAND2_X1 U7422 ( .A1(n6493), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6491) );
  OAI21_X1 U7423 ( .B1(n6493), .B2(n6492), .A(n6491), .ZN(U3472) );
  MUX2_X1 U7424 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6494), .Z(U3473) );
  NAND2_X1 U7425 ( .A1(n6495), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6504)
         );
  OAI22_X1 U7426 ( .A1(n6499), .A2(n6498), .B1(n6497), .B2(n6496), .ZN(n6500)
         );
  AOI21_X1 U7427 ( .B1(n6502), .B2(n6501), .A(n6500), .ZN(n6503) );
  OAI211_X1 U7428 ( .C1(n6506), .C2(n6505), .A(n6504), .B(n6503), .ZN(n6671)
         );
  INV_X1 U7429 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6509) );
  INV_X1 U7430 ( .A(keyinput34), .ZN(n6508) );
  AOI22_X1 U7431 ( .A1(n6509), .A2(keyinput61), .B1(ADDRESS_REG_18__SCAN_IN), 
        .B2(n6508), .ZN(n6507) );
  OAI221_X1 U7432 ( .B1(n6509), .B2(keyinput61), .C1(n6508), .C2(
        ADDRESS_REG_18__SCAN_IN), .A(n6507), .ZN(n6521) );
  INV_X1 U7433 ( .A(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n6512) );
  INV_X1 U7434 ( .A(keyinput3), .ZN(n6511) );
  AOI22_X1 U7435 ( .A1(n6512), .A2(keyinput35), .B1(LWORD_REG_1__SCAN_IN), 
        .B2(n6511), .ZN(n6510) );
  OAI221_X1 U7436 ( .B1(n6512), .B2(keyinput35), .C1(n6511), .C2(
        LWORD_REG_1__SCAN_IN), .A(n6510), .ZN(n6520) );
  INV_X1 U7437 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6515) );
  INV_X1 U7438 ( .A(keyinput55), .ZN(n6514) );
  AOI22_X1 U7439 ( .A1(n6515), .A2(keyinput17), .B1(DATAWIDTH_REG_0__SCAN_IN), 
        .B2(n6514), .ZN(n6513) );
  OAI221_X1 U7440 ( .B1(n6515), .B2(keyinput17), .C1(n6514), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(n6513), .ZN(n6519) );
  AOI22_X1 U7441 ( .A1(n5398), .A2(keyinput26), .B1(n6517), .B2(keyinput10), 
        .ZN(n6516) );
  OAI221_X1 U7442 ( .B1(n5398), .B2(keyinput26), .C1(n6517), .C2(keyinput10), 
        .A(n6516), .ZN(n6518) );
  NOR4_X1 U7443 ( .A1(n6521), .A2(n6520), .A3(n6519), .A4(n6518), .ZN(n6669)
         );
  INV_X1 U7444 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6523) );
  AOI22_X1 U7445 ( .A1(n6524), .A2(keyinput57), .B1(keyinput5), .B2(n6523), 
        .ZN(n6522) );
  OAI221_X1 U7446 ( .B1(n6524), .B2(keyinput57), .C1(n6523), .C2(keyinput5), 
        .A(n6522), .ZN(n6536) );
  AOI22_X1 U7447 ( .A1(n4782), .A2(keyinput56), .B1(keyinput40), .B2(n6526), 
        .ZN(n6525) );
  OAI221_X1 U7448 ( .B1(n4782), .B2(keyinput56), .C1(n6526), .C2(keyinput40), 
        .A(n6525), .ZN(n6535) );
  INV_X1 U7449 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U7450 ( .A1(n6529), .A2(keyinput39), .B1(keyinput53), .B2(n6528), 
        .ZN(n6527) );
  OAI221_X1 U7451 ( .B1(n6529), .B2(keyinput39), .C1(n6528), .C2(keyinput53), 
        .A(n6527), .ZN(n6534) );
  INV_X1 U7452 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6531) );
  AOI22_X1 U7453 ( .A1(n6532), .A2(keyinput23), .B1(n6531), .B2(keyinput16), 
        .ZN(n6530) );
  OAI221_X1 U7454 ( .B1(n6532), .B2(keyinput23), .C1(n6531), .C2(keyinput16), 
        .A(n6530), .ZN(n6533) );
  NOR4_X1 U7455 ( .A1(n6536), .A2(n6535), .A3(n6534), .A4(n6533), .ZN(n6668)
         );
  INV_X1 U7456 ( .A(keyinput21), .ZN(n6539) );
  INV_X1 U7457 ( .A(keyinput18), .ZN(n6538) );
  OAI22_X1 U7458 ( .A1(n6539), .A2(ADDRESS_REG_8__SCAN_IN), .B1(n6538), .B2(
        ADDRESS_REG_29__SCAN_IN), .ZN(n6537) );
  AOI221_X1 U7459 ( .B1(n6539), .B2(ADDRESS_REG_8__SCAN_IN), .C1(
        ADDRESS_REG_29__SCAN_IN), .C2(n6538), .A(n6537), .ZN(n6541) );
  XNOR2_X1 U7460 ( .A(keyinput58), .B(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6540) );
  OAI211_X1 U7461 ( .C1(keyinput11), .C2(n6542), .A(n6541), .B(n6540), .ZN(
        n6568) );
  INV_X1 U7462 ( .A(keyinput4), .ZN(n6545) );
  INV_X1 U7463 ( .A(keyinput13), .ZN(n6544) );
  OAI22_X1 U7464 ( .A1(n6545), .A2(DATAO_REG_0__SCAN_IN), .B1(n6544), .B2(
        ADDRESS_REG_6__SCAN_IN), .ZN(n6543) );
  AOI221_X1 U7465 ( .B1(n6545), .B2(DATAO_REG_0__SCAN_IN), .C1(
        ADDRESS_REG_6__SCAN_IN), .C2(n6544), .A(n6543), .ZN(n6558) );
  INV_X1 U7466 ( .A(keyinput19), .ZN(n6547) );
  OAI22_X1 U7467 ( .A1(n6548), .A2(keyinput8), .B1(n6547), .B2(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n6546) );
  AOI221_X1 U7468 ( .B1(n6548), .B2(keyinput8), .C1(DATAWIDTH_REG_12__SCAN_IN), 
        .C2(n6547), .A(n6546), .ZN(n6557) );
  INV_X1 U7469 ( .A(keyinput59), .ZN(n6550) );
  OAI22_X1 U7470 ( .A1(n6551), .A2(keyinput15), .B1(n6550), .B2(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n6549) );
  AOI221_X1 U7471 ( .B1(n6551), .B2(keyinput15), .C1(DATAWIDTH_REG_28__SCAN_IN), .C2(n6550), .A(n6549), .ZN(n6556) );
  INV_X1 U7472 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6554) );
  INV_X1 U7473 ( .A(keyinput52), .ZN(n6553) );
  OAI22_X1 U7474 ( .A1(n6554), .A2(keyinput31), .B1(n6553), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n6552) );
  AOI221_X1 U7475 ( .B1(n6554), .B2(keyinput31), .C1(DATAO_REG_27__SCAN_IN), 
        .C2(n6553), .A(n6552), .ZN(n6555) );
  NAND4_X1 U7476 ( .A1(n6558), .A2(n6557), .A3(n6556), .A4(n6555), .ZN(n6567)
         );
  AOI22_X1 U7477 ( .A1(n6561), .A2(keyinput0), .B1(n6560), .B2(keyinput33), 
        .ZN(n6559) );
  OAI221_X1 U7478 ( .B1(n6561), .B2(keyinput0), .C1(n6560), .C2(keyinput33), 
        .A(n6559), .ZN(n6566) );
  INV_X1 U7479 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6562) );
  XOR2_X1 U7480 ( .A(n6562), .B(keyinput22), .Z(n6564) );
  XNOR2_X1 U7481 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput9), .ZN(n6563)
         );
  NAND2_X1 U7482 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  NOR4_X1 U7483 ( .A1(n6568), .A2(n6567), .A3(n6566), .A4(n6565), .ZN(n6667)
         );
  INV_X1 U7484 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6570) );
  AOI22_X1 U7485 ( .A1(n6571), .A2(keyinput50), .B1(n6570), .B2(keyinput44), 
        .ZN(n6569) );
  OAI221_X1 U7486 ( .B1(n6571), .B2(keyinput50), .C1(n6570), .C2(keyinput44), 
        .A(n6569), .ZN(n6665) );
  AOI22_X1 U7487 ( .A1(n6574), .A2(keyinput49), .B1(keyinput14), .B2(n6573), 
        .ZN(n6572) );
  OAI221_X1 U7488 ( .B1(n6574), .B2(keyinput49), .C1(n6573), .C2(keyinput14), 
        .A(n6572), .ZN(n6664) );
  INV_X1 U7489 ( .A(keyinput41), .ZN(n6576) );
  OAI22_X1 U7490 ( .A1(keyinput2), .A2(n6577), .B1(n6576), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6575) );
  AOI221_X1 U7491 ( .B1(n6577), .B2(keyinput2), .C1(n6576), .C2(
        LWORD_REG_11__SCAN_IN), .A(n6575), .ZN(n6599) );
  INV_X1 U7492 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6580) );
  OAI22_X1 U7493 ( .A1(n6580), .A2(keyinput27), .B1(n6579), .B2(keyinput24), 
        .ZN(n6578) );
  AOI221_X1 U7494 ( .B1(n6580), .B2(keyinput27), .C1(keyinput24), .C2(n6579), 
        .A(n6578), .ZN(n6598) );
  INV_X1 U7495 ( .A(keyinput32), .ZN(n6582) );
  AOI22_X1 U7496 ( .A1(n6583), .A2(keyinput43), .B1(DATAO_REG_3__SCAN_IN), 
        .B2(n6582), .ZN(n6581) );
  OAI221_X1 U7497 ( .B1(n6583), .B2(keyinput43), .C1(n6582), .C2(
        DATAO_REG_3__SCAN_IN), .A(n6581), .ZN(n6596) );
  INV_X1 U7498 ( .A(keyinput46), .ZN(n6585) );
  AOI22_X1 U7499 ( .A1(n6586), .A2(keyinput38), .B1(ADDRESS_REG_2__SCAN_IN), 
        .B2(n6585), .ZN(n6584) );
  OAI221_X1 U7500 ( .B1(n6586), .B2(keyinput38), .C1(n6585), .C2(
        ADDRESS_REG_2__SCAN_IN), .A(n6584), .ZN(n6595) );
  INV_X1 U7501 ( .A(keyinput54), .ZN(n6589) );
  INV_X1 U7502 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6588) );
  AOI22_X1 U7503 ( .A1(n6589), .A2(UWORD_REG_14__SCAN_IN), .B1(keyinput28), 
        .B2(n6588), .ZN(n6587) );
  OAI221_X1 U7504 ( .B1(n6589), .B2(UWORD_REG_14__SCAN_IN), .C1(n6588), .C2(
        keyinput28), .A(n6587), .ZN(n6594) );
  INV_X1 U7505 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6592) );
  AOI22_X1 U7506 ( .A1(n6592), .A2(keyinput12), .B1(keyinput36), .B2(n6591), 
        .ZN(n6590) );
  OAI221_X1 U7507 ( .B1(n6592), .B2(keyinput12), .C1(n6591), .C2(keyinput36), 
        .A(n6590), .ZN(n6593) );
  NOR4_X1 U7508 ( .A1(n6596), .A2(n6595), .A3(n6594), .A4(n6593), .ZN(n6597)
         );
  NAND3_X1 U7509 ( .A1(n6599), .A2(n6598), .A3(n6597), .ZN(n6663) );
  NAND2_X1 U7510 ( .A1(keyinput58), .A2(keyinput22), .ZN(n6605) );
  INV_X1 U7511 ( .A(keyinput17), .ZN(n6600) );
  NAND4_X1 U7512 ( .A1(keyinput55), .A2(keyinput35), .A3(keyinput26), .A4(
        n6600), .ZN(n6604) );
  NOR3_X1 U7513 ( .A1(keyinput9), .A2(keyinput0), .A3(keyinput21), .ZN(n6602)
         );
  NOR3_X1 U7514 ( .A1(keyinput34), .A2(keyinput61), .A3(keyinput3), .ZN(n6601)
         );
  NAND4_X1 U7515 ( .A1(keyinput33), .A2(n6602), .A3(keyinput18), .A4(n6601), 
        .ZN(n6603) );
  NOR4_X1 U7516 ( .A1(keyinput54), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(
        n6629) );
  NAND3_X1 U7517 ( .A1(keyinput31), .A2(keyinput57), .A3(keyinput56), .ZN(
        n6627) );
  NAND2_X1 U7518 ( .A1(keyinput19), .A2(keyinput10), .ZN(n6606) );
  NOR3_X1 U7519 ( .A1(keyinput13), .A2(keyinput4), .A3(n6606), .ZN(n6610) );
  NAND2_X1 U7520 ( .A1(keyinput52), .A2(keyinput59), .ZN(n6607) );
  NOR3_X1 U7521 ( .A1(keyinput8), .A2(keyinput15), .A3(n6607), .ZN(n6609) );
  NOR3_X1 U7522 ( .A1(keyinput39), .A2(keyinput53), .A3(keyinput23), .ZN(n6608) );
  NAND4_X1 U7523 ( .A1(n6610), .A2(n6609), .A3(keyinput40), .A4(n6608), .ZN(
        n6626) );
  NOR4_X1 U7524 ( .A1(keyinput63), .A2(keyinput30), .A3(keyinput1), .A4(
        keyinput48), .ZN(n6624) );
  NAND3_X1 U7525 ( .A1(keyinput16), .A2(keyinput45), .A3(keyinput20), .ZN(
        n6615) );
  INV_X1 U7526 ( .A(keyinput6), .ZN(n6611) );
  NAND4_X1 U7527 ( .A1(keyinput29), .A2(keyinput62), .A3(keyinput51), .A4(
        n6611), .ZN(n6614) );
  INV_X1 U7528 ( .A(keyinput60), .ZN(n6612) );
  NAND4_X1 U7529 ( .A1(keyinput7), .A2(keyinput25), .A3(keyinput37), .A4(n6612), .ZN(n6613) );
  NOR4_X1 U7530 ( .A1(keyinput47), .A2(n6615), .A3(n6614), .A4(n6613), .ZN(
        n6623) );
  NAND2_X1 U7531 ( .A1(keyinput2), .A2(keyinput27), .ZN(n6616) );
  NOR3_X1 U7532 ( .A1(keyinput32), .A2(keyinput24), .A3(n6616), .ZN(n6622) );
  NAND2_X1 U7533 ( .A1(keyinput41), .A2(keyinput36), .ZN(n6620) );
  NOR3_X1 U7534 ( .A1(keyinput42), .A2(keyinput14), .A3(keyinput50), .ZN(n6618) );
  NOR3_X1 U7535 ( .A1(keyinput44), .A2(keyinput38), .A3(keyinput43), .ZN(n6617) );
  NAND4_X1 U7536 ( .A1(keyinput49), .A2(n6618), .A3(keyinput46), .A4(n6617), 
        .ZN(n6619) );
  NOR4_X1 U7537 ( .A1(keyinput12), .A2(keyinput28), .A3(n6620), .A4(n6619), 
        .ZN(n6621) );
  NAND4_X1 U7538 ( .A1(n6624), .A2(n6623), .A3(n6622), .A4(n6621), .ZN(n6625)
         );
  NOR4_X1 U7539 ( .A1(keyinput5), .A2(n6627), .A3(n6626), .A4(n6625), .ZN(
        n6628) );
  AOI21_X1 U7540 ( .B1(n6629), .B2(n6628), .A(keyinput11), .ZN(n6661) );
  INV_X1 U7541 ( .A(keyinput37), .ZN(n6632) );
  INV_X1 U7542 ( .A(keyinput42), .ZN(n6631) );
  AOI22_X1 U7543 ( .A1(n6632), .A2(DATAO_REG_7__SCAN_IN), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6631), .ZN(n6630) );
  OAI221_X1 U7544 ( .B1(n6632), .B2(DATAO_REG_7__SCAN_IN), .C1(n6631), .C2(
        ADDRESS_REG_5__SCAN_IN), .A(n6630), .ZN(n6643) );
  AOI22_X1 U7545 ( .A1(n6635), .A2(keyinput51), .B1(n6634), .B2(keyinput7), 
        .ZN(n6633) );
  OAI221_X1 U7546 ( .B1(n6635), .B2(keyinput51), .C1(n6634), .C2(keyinput7), 
        .A(n6633), .ZN(n6642) );
  XOR2_X1 U7547 ( .A(n6636), .B(keyinput29), .Z(n6640) );
  XNOR2_X1 U7548 ( .A(keyinput60), .B(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6639) );
  XNOR2_X1 U7549 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .B(keyinput6), .ZN(n6638)
         );
  XNOR2_X1 U7550 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput25), .ZN(
        n6637) );
  NAND4_X1 U7551 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n6641)
         );
  NOR3_X1 U7552 ( .A1(n6643), .A2(n6642), .A3(n6641), .ZN(n6660) );
  INV_X1 U7553 ( .A(keyinput63), .ZN(n6645) );
  AOI22_X1 U7554 ( .A1(n6646), .A2(keyinput47), .B1(DATAO_REG_11__SCAN_IN), 
        .B2(n6645), .ZN(n6644) );
  OAI221_X1 U7555 ( .B1(n6646), .B2(keyinput47), .C1(n6645), .C2(
        DATAO_REG_11__SCAN_IN), .A(n6644), .ZN(n6658) );
  AOI22_X1 U7556 ( .A1(n6648), .A2(keyinput45), .B1(keyinput20), .B2(n4113), 
        .ZN(n6647) );
  OAI221_X1 U7557 ( .B1(n6648), .B2(keyinput45), .C1(n4113), .C2(keyinput20), 
        .A(n6647), .ZN(n6657) );
  INV_X1 U7558 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6650) );
  AOI22_X1 U7559 ( .A1(n6651), .A2(keyinput48), .B1(n6650), .B2(keyinput62), 
        .ZN(n6649) );
  OAI221_X1 U7560 ( .B1(n6651), .B2(keyinput48), .C1(n6650), .C2(keyinput62), 
        .A(n6649), .ZN(n6656) );
  AOI22_X1 U7561 ( .A1(n6654), .A2(keyinput30), .B1(n6653), .B2(keyinput1), 
        .ZN(n6652) );
  OAI221_X1 U7562 ( .B1(n6654), .B2(keyinput30), .C1(n6653), .C2(keyinput1), 
        .A(n6652), .ZN(n6655) );
  NOR4_X1 U7563 ( .A1(n6658), .A2(n6657), .A3(n6656), .A4(n6655), .ZN(n6659)
         );
  OAI211_X1 U7564 ( .C1(EAX_REG_1__SCAN_IN), .C2(n6661), .A(n6660), .B(n6659), 
        .ZN(n6662) );
  NOR4_X1 U7565 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6666)
         );
  NAND4_X1 U7566 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6670)
         );
  XNOR2_X1 U7567 ( .A(n6671), .B(n6670), .ZN(U3139) );
  CLKBUF_X1 U3417 ( .A(n3194), .Z(n3435) );
  CLKBUF_X1 U34460 ( .A(n5993), .Z(n6002) );
  CLKBUF_X1 U3480 ( .A(n4533), .Z(n2969) );
endmodule

