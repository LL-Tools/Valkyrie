

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915;

  NAND2_X2 U2250 ( .A1(n2023), .A2(n2127), .ZN(n4309) );
  CLKBUF_X2 U2252 ( .A(n3260), .Z(n4253) );
  AND4_X2 U2253 ( .A1(n2544), .A2(n2543), .A3(n2542), .A4(n2541), .ZN(n3165)
         );
  CLKBUF_X1 U2254 ( .A(n2576), .Z(n2012) );
  INV_X1 U2255 ( .A(IR_REG_31__SCAN_IN), .ZN(n2472) );
  INV_X1 U2256 ( .A(n3267), .ZN(n3383) );
  CLKBUF_X2 U2257 ( .A(n3264), .Z(n4043) );
  NAND2_X1 U2258 ( .A1(n2140), .A2(n2137), .ZN(n3764) );
  NAND2_X1 U2259 ( .A1(n2900), .A2(n2862), .ZN(n3256) );
  OR2_X1 U2260 ( .A1(n4390), .A2(n3929), .ZN(n2170) );
  INV_X1 U2261 ( .A(n3261), .ZN(n3164) );
  NAND2_X1 U2262 ( .A1(n2014), .A2(REG3_REG_1__SCAN_IN), .ZN(n2337) );
  INV_X2 U2263 ( .A(n3652), .ZN(n4078) );
  INV_X1 U2264 ( .A(n4311), .ZN(n3361) );
  NAND4_X1 U2265 ( .A1(n2336), .A2(n2337), .A3(n2335), .A4(n2334), .ZN(n3260)
         );
  NAND2_X1 U2266 ( .A1(n2530), .A2(n2531), .ZN(n2805) );
  INV_X1 U2267 ( .A(n4426), .ZN(n4396) );
  AOI211_X1 U2268 ( .C1(n2333), .C2(n4823), .A(n3229), .B(n3228), .ZN(n3298)
         );
  INV_X1 U2269 ( .A(n4915), .ZN(n4912) );
  NAND2_X1 U2270 ( .A1(n3111), .A2(n3191), .ZN(n4870) );
  INV_X2 U2271 ( .A(n2376), .ZN(n2377) );
  NAND3_X2 U2272 ( .A1(n2356), .A2(n2333), .A3(n2332), .ZN(n2376) );
  INV_X2 U2273 ( .A(n2390), .ZN(n2164) );
  NAND2_X2 U2274 ( .A1(n2377), .A2(n2347), .ZN(n2390) );
  INV_X4 U2275 ( .A(IR_REG_0__SCAN_IN), .ZN(n2333) );
  CLKBUF_X1 U2276 ( .A(n2914), .Z(n2008) );
  BUF_X4 U2277 ( .A(n2914), .Z(n2009) );
  INV_X2 U2278 ( .A(n2805), .ZN(n2914) );
  AND2_X4 U2279 ( .A1(n3256), .A2(n3245), .ZN(n4079) );
  NAND4_X2 U2280 ( .A1(n2463), .A2(n3105), .A3(n3101), .A4(n2462), .ZN(n3245)
         );
  NAND2_X2 U2281 ( .A1(n3161), .A2(n3162), .ZN(n3160) );
  XNOR2_X2 U2282 ( .A(n2464), .B(IR_REG_22__SCAN_IN), .ZN(n2807) );
  NOR2_X2 U2283 ( .A1(n4829), .A2(n2257), .ZN(n2439) );
  OAI21_X2 U2284 ( .B1(n4327), .B2(n2432), .A(n2433), .ZN(n2135) );
  NAND2_X2 U2285 ( .A1(n2428), .A2(n2427), .ZN(n4327) );
  NAND2_X2 U2286 ( .A1(n3425), .A2(n2827), .ZN(n2829) );
  NAND2_X2 U2287 ( .A1(n2826), .A2(n2825), .ZN(n3425) );
  NAND2_X2 U2288 ( .A1(n4609), .A2(n2839), .ZN(n2343) );
  NAND2_X2 U2289 ( .A1(n3092), .A2(IR_REG_31__SCAN_IN), .ZN(n2132) );
  CLKBUF_X1 U2290 ( .A(n3194), .Z(n4597) );
  INV_X2 U2291 ( .A(n3264), .ZN(n4087) );
  AND4_X1 U2292 ( .A1(n2596), .A2(n2595), .A3(n2594), .A4(n2593), .ZN(n3539)
         );
  BUF_X2 U2293 ( .A(n2012), .Z(n2913) );
  NOR2_X1 U2294 ( .A1(n2459), .A2(n2458), .ZN(n3105) );
  CLKBUF_X2 U2296 ( .A(IR_REG_0__SCAN_IN), .Z(n2379) );
  AND2_X1 U2297 ( .A1(n2207), .A2(n2168), .ZN(n2167) );
  MUX2_X1 U2298 ( .A(n3969), .B(n3968), .S(n4811), .Z(n3970) );
  NAND2_X1 U2299 ( .A1(n2131), .A2(n2130), .ZN(n2282) );
  NAND2_X1 U2300 ( .A1(n2700), .A2(n3940), .ZN(n4485) );
  NOR2_X1 U2301 ( .A1(n2910), .A2(n4386), .ZN(n4385) );
  AND2_X1 U2302 ( .A1(n4470), .A2(n4474), .ZN(n4472) );
  NAND2_X1 U2303 ( .A1(n2273), .A2(n2272), .ZN(n3417) );
  NAND2_X1 U2304 ( .A1(n2575), .A2(n3835), .ZN(n3571) );
  NAND2_X1 U2305 ( .A1(n2728), .A2(n2727), .ZN(n4665) );
  NAND2_X1 U2306 ( .A1(n2214), .A2(n2211), .ZN(n3301) );
  NOR2_X1 U2307 ( .A1(n3647), .A2(n2276), .ZN(n2275) );
  OR2_X1 U2308 ( .A1(n2045), .A2(n2302), .ZN(n2300) );
  NOR2_X1 U2309 ( .A1(n3481), .A2(n3480), .ZN(n2302) );
  NAND2_X1 U2310 ( .A1(n3572), .A2(n3599), .ZN(n3839) );
  AND2_X1 U2311 ( .A1(n3829), .A2(n3826), .ZN(n3912) );
  BUF_X2 U2312 ( .A(n3383), .Z(n3652) );
  NAND2_X1 U2313 ( .A1(n3211), .A2(n3261), .ZN(n3824) );
  AND2_X2 U2314 ( .A1(n3207), .A2(n4896), .ZN(n4859) );
  INV_X1 U2315 ( .A(n3539), .ZN(n4307) );
  NAND4_X1 U2316 ( .A1(n2632), .A2(n2631), .A3(n2630), .A4(n2629), .ZN(n4736)
         );
  INV_X1 U2317 ( .A(n4079), .ZN(n4089) );
  INV_X1 U2318 ( .A(n3256), .ZN(n3462) );
  NAND4_X2 U2319 ( .A1(n2551), .A2(n2550), .A3(n2549), .A4(n2548), .ZN(n4311)
         );
  NAND2_X1 U2320 ( .A1(n2012), .A2(REG2_REG_3__SCAN_IN), .ZN(n2548) );
  OR2_X1 U2321 ( .A1(n2636), .A2(n2635), .ZN(n2641) );
  OAI21_X1 U2322 ( .B1(n2798), .B2(n2792), .A(n2348), .ZN(n2900) );
  INV_X1 U2323 ( .A(n3340), .ZN(n3349) );
  OAI21_X1 U2324 ( .B1(n2011), .B2(n2554), .A(n2553), .ZN(n3340) );
  XNOR2_X1 U2325 ( .A(n2388), .B(n3295), .ZN(n3290) );
  INV_X1 U2326 ( .A(n3570), .ZN(n3572) );
  NAND2_X1 U2327 ( .A1(n2240), .A2(n2384), .ZN(n2388) );
  OAI21_X1 U2328 ( .B1(n2533), .B2(n3295), .A(n2171), .ZN(n3470) );
  INV_X2 U2329 ( .A(n2533), .ZN(n2909) );
  OR2_X1 U2330 ( .A1(n2465), .A2(n2472), .ZN(n2464) );
  AND2_X1 U2331 ( .A1(n2466), .A2(n2467), .ZN(n2465) );
  XNOR2_X1 U2332 ( .A(n2471), .B(IR_REG_26__SCAN_IN), .ZN(n3101) );
  MUX2_X1 U2333 ( .A(n2456), .B(n2472), .S(n2518), .Z(n2459) );
  NOR2_X1 U2334 ( .A1(n2447), .A2(n2452), .ZN(n2466) );
  NAND2_X1 U2335 ( .A1(n2457), .A2(n2518), .ZN(n2477) );
  AND4_X1 U2336 ( .A1(n2113), .A2(n2112), .A3(n2111), .A4(n2114), .ZN(n2454)
         );
  AND2_X1 U2337 ( .A1(n2929), .A2(n2357), .ZN(n2347) );
  INV_X1 U2338 ( .A(IR_REG_26__SCAN_IN), .ZN(n2519) );
  INV_X1 U2339 ( .A(IR_REG_24__SCAN_IN), .ZN(n2871) );
  NOR2_X1 U2340 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2111)
         );
  NOR2_X1 U2341 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2112)
         );
  NOR2_X1 U2342 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2113)
         );
  INV_X1 U2343 ( .A(IR_REG_22__SCAN_IN), .ZN(n2925) );
  INV_X1 U2344 ( .A(IR_REG_21__SCAN_IN), .ZN(n2467) );
  INV_X1 U2345 ( .A(IR_REG_13__SCAN_IN), .ZN(n2455) );
  NOR2_X1 U2346 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2360)
         );
  NOR2_X1 U2347 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2361)
         );
  INV_X1 U2348 ( .A(IR_REG_2__SCAN_IN), .ZN(n2356) );
  NOR2_X1 U2349 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2359)
         );
  AND3_X1 U2350 ( .A1(n2166), .A2(n2162), .A3(n2164), .ZN(n2457) );
  OAI21_X1 U2351 ( .B1(n4468), .B2(n2854), .A(n2330), .ZN(n4453) );
  NAND2_X1 U2352 ( .A1(n4468), .A2(n2327), .ZN(n2324) );
  INV_X4 U2353 ( .A(n2533), .ZN(n2011) );
  AND2_X2 U2354 ( .A1(n2164), .A2(n2163), .ZN(n2524) );
  OAI21_X4 U2355 ( .B1(n4115), .B2(n2308), .A(n2305), .ZN(n4134) );
  NAND2_X2 U2356 ( .A1(n3990), .A2(n3989), .ZN(n4115) );
  INV_X1 U2357 ( .A(n3354), .ZN(n3913) );
  NAND2_X2 U2358 ( .A1(n4634), .A2(n2838), .ZN(n4609) );
  INV_X1 U2359 ( .A(n3165), .ZN(n4313) );
  NOR2_X1 U2360 ( .A1(n2378), .A2(n2377), .ZN(n2485) );
  MUX2_X2 U2361 ( .A(n3088), .B(n3087), .S(n4905), .Z(n3090) );
  MUX2_X2 U2362 ( .A(n3088), .B(n3083), .S(n4912), .Z(n3086) );
  AND2_X1 U2363 ( .A1(n4809), .A2(n3097), .ZN(n2014) );
  AND2_X4 U2364 ( .A1(n4809), .A2(n3097), .ZN(n2581) );
  NAND3_X1 U2365 ( .A1(n2455), .A2(n2925), .A3(n2467), .ZN(n2517) );
  NAND2_X1 U2366 ( .A1(n4134), .A2(n2050), .ZN(n2131) );
  INV_X1 U2367 ( .A(n2581), .ZN(n2782) );
  NAND2_X1 U2368 ( .A1(n3256), .A2(n3255), .ZN(n3264) );
  INV_X1 U2369 ( .A(n2159), .ZN(n2158) );
  OAI21_X1 U2370 ( .B1(n2342), .B2(n2160), .A(n2843), .ZN(n2159) );
  AND2_X1 U2371 ( .A1(n2317), .A2(n2016), .ZN(n2314) );
  AND2_X1 U2372 ( .A1(n2020), .A2(n3911), .ZN(n2340) );
  AND2_X1 U2373 ( .A1(n2807), .A2(n2862), .ZN(n3185) );
  NAND2_X1 U2374 ( .A1(n4077), .A2(n2031), .ZN(n2116) );
  INV_X1 U2375 ( .A(n4273), .ZN(n2117) );
  NOR2_X1 U2376 ( .A1(n2286), .A2(n4030), .ZN(n2130) );
  INV_X1 U2377 ( .A(n2287), .ZN(n2286) );
  NOR2_X1 U2378 ( .A1(n2082), .A2(n3330), .ZN(n2081) );
  INV_X1 U2379 ( .A(n2349), .ZN(n2082) );
  NAND2_X1 U2380 ( .A1(n2042), .A2(n2074), .ZN(n2221) );
  NAND2_X1 U2381 ( .A1(n2498), .A2(n2497), .ZN(n3683) );
  INV_X1 U2382 ( .A(n3685), .ZN(n2497) );
  AND2_X1 U2383 ( .A1(n2435), .A2(n2258), .ZN(n4829) );
  INV_X1 U2384 ( .A(n4830), .ZN(n2258) );
  NAND2_X1 U2385 ( .A1(n2271), .A2(n2665), .ZN(n2270) );
  NAND2_X1 U2386 ( .A1(n2073), .A2(n2057), .ZN(n2072) );
  INV_X1 U2387 ( .A(n4848), .ZN(n2073) );
  NAND2_X1 U2388 ( .A1(n2070), .A2(n2072), .ZN(n4367) );
  AND2_X1 U2389 ( .A1(n2237), .A2(n2071), .ZN(n2070) );
  AND2_X1 U2390 ( .A1(n2509), .A2(n2056), .ZN(n2071) );
  AND2_X1 U2391 ( .A1(n2278), .A2(n2344), .ZN(n2161) );
  AND2_X1 U2392 ( .A1(n2769), .A2(n2768), .ZN(n4438) );
  OR2_X1 U2393 ( .A1(n4421), .A2(n2782), .ZN(n2769) );
  NAND2_X1 U2394 ( .A1(n4515), .A2(n2850), .ZN(n4484) );
  NAND2_X1 U2395 ( .A1(n2343), .A2(n2342), .ZN(n4587) );
  NAND2_X1 U2396 ( .A1(n3775), .A2(n2836), .ZN(n2153) );
  INV_X1 U2397 ( .A(n4678), .ZN(n4900) );
  INV_X1 U2398 ( .A(n3403), .ZN(n2147) );
  NOR2_X1 U2399 ( .A1(n2147), .A2(n2148), .ZN(n2145) );
  INV_X1 U2400 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2148) );
  NOR2_X1 U2401 ( .A1(n4328), .A2(n2235), .ZN(n2234) );
  NOR2_X1 U2402 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2358)
         );
  NOR2_X1 U2403 ( .A1(n2641), .A2(n3041), .ZN(n2654) );
  NAND2_X1 U2404 ( .A1(n2061), .A2(REG3_REG_13__SCAN_IN), .ZN(n2636) );
  INV_X1 U2405 ( .A(n2627), .ZN(n2061) );
  XNOR2_X1 U2406 ( .A(n3265), .B(n4087), .ZN(n3271) );
  AND2_X1 U2407 ( .A1(n3888), .A2(n4464), .ZN(n3948) );
  AND2_X1 U2408 ( .A1(n2010), .A2(REG1_REG_2__SCAN_IN), .ZN(n2487) );
  AND2_X1 U2409 ( .A1(n4821), .A2(REG1_REG_1__SCAN_IN), .ZN(n2091) );
  INV_X1 U2410 ( .A(n2487), .ZN(n2084) );
  INV_X1 U2411 ( .A(n2246), .ZN(n2244) );
  INV_X1 U2412 ( .A(n2228), .ZN(n2227) );
  AOI22_X1 U2413 ( .A1(n3767), .A2(n2234), .B1(n4814), .B2(n2233), .ZN(n2228)
         );
  INV_X1 U2414 ( .A(n2234), .ZN(n2229) );
  INV_X1 U2415 ( .A(n3945), .ZN(n2198) );
  NAND2_X1 U2416 ( .A1(n4683), .A2(n4549), .ZN(n3905) );
  INV_X1 U2417 ( .A(n2319), .ZN(n2315) );
  INV_X1 U2418 ( .A(n3306), .ZN(n2817) );
  OAI21_X1 U2419 ( .B1(n3161), .B2(n3819), .A(n3824), .ZN(n3357) );
  NAND2_X1 U2420 ( .A1(n3164), .A2(n3260), .ZN(n3820) );
  NOR2_X1 U2421 ( .A1(n4557), .A2(n4682), .ZN(n4517) );
  NOR2_X1 U2422 ( .A1(n2188), .A2(n4143), .ZN(n2187) );
  NAND2_X1 U2423 ( .A1(n4620), .A2(n4598), .ZN(n2188) );
  NAND2_X1 U2424 ( .A1(n3991), .A2(n3677), .ZN(n2175) );
  NAND2_X1 U2425 ( .A1(n2184), .A2(n2183), .ZN(n2182) );
  NAND2_X1 U2426 ( .A1(n3182), .A2(n2808), .ZN(n2899) );
  INV_X1 U2427 ( .A(n3456), .ZN(n3458) );
  NOR2_X1 U2428 ( .A1(n2165), .A2(n2517), .ZN(n2162) );
  NAND2_X1 U2429 ( .A1(n2346), .A2(n2363), .ZN(n2364) );
  INV_X1 U2430 ( .A(IR_REG_16__SCAN_IN), .ZN(n2362) );
  INV_X1 U2431 ( .A(IR_REG_17__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U2432 ( .A1(n4057), .A2(n4056), .ZN(n4125) );
  INV_X1 U2433 ( .A(n4127), .ZN(n4056) );
  INV_X1 U2434 ( .A(n4126), .ZN(n4057) );
  NAND2_X1 U2435 ( .A1(n2701), .A2(REG3_REG_22__SCAN_IN), .ZN(n2721) );
  INV_X1 U2436 ( .A(n2713), .ZN(n2701) );
  OR2_X1 U2437 ( .A1(n2721), .A2(n4129), .ZN(n2733) );
  NAND2_X1 U2438 ( .A1(n2666), .A2(REG3_REG_18__SCAN_IN), .ZN(n2679) );
  INV_X1 U2439 ( .A(n2677), .ZN(n2666) );
  OR2_X1 U2440 ( .A1(n2711), .A2(n2710), .ZN(n2713) );
  NAND2_X1 U2441 ( .A1(n2297), .A2(n2296), .ZN(n2295) );
  NAND2_X1 U2442 ( .A1(n4175), .A2(n4174), .ZN(n2296) );
  NAND2_X1 U2443 ( .A1(n4171), .A2(n4073), .ZN(n2297) );
  INV_X1 U2444 ( .A(n2295), .ZN(n2293) );
  NAND2_X1 U2445 ( .A1(n4209), .A2(n4173), .ZN(n2298) );
  NOR2_X1 U2446 ( .A1(n2295), .A2(n2298), .ZN(n2291) );
  INV_X1 U2447 ( .A(n2654), .ZN(n2657) );
  NAND2_X1 U2448 ( .A1(n3392), .A2(n2128), .ZN(n3393) );
  NAND2_X1 U2449 ( .A1(n2129), .A2(n4309), .ZN(n2128) );
  INV_X1 U2450 ( .A(n4011), .ZN(n2311) );
  OR2_X1 U2451 ( .A1(n3542), .A2(n3541), .ZN(n3648) );
  OAI21_X1 U2452 ( .B1(n3282), .B2(n3196), .A(n3195), .ZN(n3204) );
  NAND2_X1 U2453 ( .A1(n2605), .A2(REG3_REG_10__SCAN_IN), .ZN(n2620) );
  INV_X1 U2454 ( .A(n2607), .ZN(n2605) );
  OR2_X1 U2455 ( .A1(n2311), .A2(n4198), .ZN(n2307) );
  OAI22_X1 U2456 ( .A1(n4010), .A2(n4190), .B1(n2310), .B2(n4011), .ZN(n2309)
         );
  INV_X1 U2457 ( .A(n4117), .ZN(n2310) );
  NAND2_X1 U2458 ( .A1(n2563), .A2(REG3_REG_5__SCAN_IN), .ZN(n2569) );
  INV_X1 U2459 ( .A(n4314), .ZN(n2089) );
  INV_X1 U2460 ( .A(n3237), .ZN(n2087) );
  INV_X1 U2461 ( .A(n2393), .ZN(n2250) );
  NAND2_X1 U2462 ( .A1(n2224), .A2(n2068), .ZN(n2067) );
  NOR2_X1 U2463 ( .A1(n2069), .A2(n2054), .ZN(n2068) );
  INV_X1 U2464 ( .A(n2222), .ZN(n2069) );
  NAND2_X1 U2465 ( .A1(n3683), .A2(n2351), .ZN(n2066) );
  INV_X1 U2466 ( .A(n4328), .ZN(n2233) );
  NOR2_X1 U2467 ( .A1(n3767), .A2(n2139), .ZN(n2138) );
  NOR2_X1 U2468 ( .A1(n2267), .A2(n4356), .ZN(n2265) );
  OR2_X1 U2469 ( .A1(n2263), .A2(n2265), .ZN(n2262) );
  INV_X1 U2470 ( .A(n2264), .ZN(n2263) );
  OAI21_X1 U2471 ( .B1(n2484), .B2(n2441), .A(n2268), .ZN(n2264) );
  OR2_X1 U2472 ( .A1(n2773), .A2(n2772), .ZN(n4397) );
  NAND2_X1 U2473 ( .A1(n4434), .A2(n3952), .ZN(n2210) );
  OAI21_X1 U2474 ( .B1(n2856), .B2(n2326), .A(n2855), .ZN(n2325) );
  NAND2_X1 U2475 ( .A1(n2854), .A2(n2330), .ZN(n2326) );
  NOR2_X1 U2476 ( .A1(n2856), .A2(n2328), .ZN(n2327) );
  INV_X1 U2477 ( .A(n2330), .ZN(n2328) );
  NAND2_X1 U2478 ( .A1(n4485), .A2(n3944), .ZN(n2195) );
  NAND2_X1 U2479 ( .A1(n4528), .A2(n2846), .ZN(n2848) );
  AOI21_X1 U2480 ( .B1(n2158), .B2(n2160), .A(n2040), .ZN(n2156) );
  INV_X1 U2481 ( .A(n2063), .ZN(n2691) );
  NAND2_X1 U2482 ( .A1(n2063), .A2(REG3_REG_20__SCAN_IN), .ZN(n2711) );
  INV_X1 U2483 ( .A(n4507), .ZN(n4551) );
  AOI21_X1 U2484 ( .B1(n2202), .B2(n2204), .A(n2037), .ZN(n2200) );
  AOI21_X1 U2485 ( .B1(n2340), .B2(n2835), .A(n2035), .ZN(n2338) );
  NOR2_X1 U2486 ( .A1(n2830), .A2(n2318), .ZN(n2317) );
  INV_X1 U2487 ( .A(n2828), .ZN(n2318) );
  INV_X1 U2488 ( .A(n3566), .ZN(n3567) );
  INV_X1 U2489 ( .A(n2212), .ZN(n2211) );
  NAND2_X1 U2490 ( .A1(n3467), .A2(n2215), .ZN(n2214) );
  OAI21_X1 U2491 ( .B1(n3833), .B2(n2213), .A(n3844), .ZN(n2212) );
  NAND2_X1 U2492 ( .A1(n2561), .A2(n4310), .ZN(n3832) );
  AND2_X1 U2493 ( .A1(n3178), .A2(n3177), .ZN(n3452) );
  INV_X1 U2494 ( .A(n4590), .ZN(n4631) );
  AND2_X1 U2495 ( .A1(n2891), .A2(n2890), .ZN(n3180) );
  AND2_X1 U2496 ( .A1(n4517), .A2(n2896), .ZN(n4516) );
  NOR2_X1 U2497 ( .A1(n4618), .A2(n2188), .ZN(n4599) );
  AND3_X1 U2498 ( .A1(n2889), .A2(n2888), .A3(n3178), .ZN(n2922) );
  NOR2_X1 U2499 ( .A1(n2523), .A2(n2522), .ZN(n2525) );
  NAND2_X1 U2500 ( .A1(n2420), .A2(IR_REG_31__SCAN_IN), .ZN(n2424) );
  INV_X1 U2501 ( .A(IR_REG_6__SCAN_IN), .ZN(n2399) );
  INV_X1 U2502 ( .A(IR_REG_4__SCAN_IN), .ZN(n2357) );
  NAND2_X1 U2503 ( .A1(n2356), .A2(n2472), .ZN(n2374) );
  NAND2_X1 U2504 ( .A1(n3395), .A2(n2110), .ZN(n2109) );
  NAND2_X1 U2505 ( .A1(n2116), .A2(n2115), .ZN(n4106) );
  NOR2_X1 U2506 ( .A1(n2119), .A2(n4107), .ZN(n2115) );
  NAND2_X1 U2507 ( .A1(n2034), .A2(n2122), .ZN(n2121) );
  INV_X1 U2508 ( .A(n3470), .ZN(n2561) );
  INV_X1 U2509 ( .A(n4238), .ZN(n2281) );
  OAI21_X1 U2510 ( .B1(n2011), .B2(n2546), .A(n2545), .ZN(n4252) );
  NAND2_X1 U2511 ( .A1(n2909), .A2(n2010), .ZN(n2545) );
  INV_X1 U2512 ( .A(n4296), .ZN(n4250) );
  OR2_X1 U2513 ( .A1(n3251), .A2(n4822), .ZN(n4267) );
  INV_X1 U2514 ( .A(n4276), .ZN(n4294) );
  NAND2_X1 U2515 ( .A1(n2758), .A2(n2757), .ZN(n4424) );
  OR2_X1 U2516 ( .A1(n4446), .A2(n2782), .ZN(n2758) );
  INV_X1 U2517 ( .A(n4718), .ZN(n4611) );
  NAND2_X1 U2518 ( .A1(n3142), .A2(n2491), .ZN(n3214) );
  NAND2_X1 U2519 ( .A1(n2067), .A2(n2251), .ZN(n2491) );
  NAND2_X1 U2520 ( .A1(n3214), .A2(n2492), .ZN(n2493) );
  OR2_X1 U2521 ( .A1(n4818), .A2(REG1_REG_7__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U2522 ( .A1(n2493), .A2(n2081), .ZN(n2076) );
  NAND2_X1 U2523 ( .A1(n3328), .A2(REG2_REG_8__SCAN_IN), .ZN(n2146) );
  INV_X1 U2524 ( .A(n2221), .ZN(n3406) );
  INV_X1 U2525 ( .A(n3405), .ZN(n2220) );
  INV_X1 U2526 ( .A(n4840), .ZN(n4342) );
  INV_X1 U2527 ( .A(n2435), .ZN(n4831) );
  NAND2_X1 U2528 ( .A1(n2096), .A2(n2502), .ZN(n4835) );
  OR2_X1 U2529 ( .A1(n4338), .A2(n4731), .ZN(n2096) );
  OR2_X1 U2530 ( .A1(n4828), .A2(n4810), .ZN(n4360) );
  NAND2_X1 U2531 ( .A1(n2483), .A2(n2484), .ZN(n2151) );
  NAND2_X1 U2532 ( .A1(n2270), .A2(n2269), .ZN(n2483) );
  AOI21_X1 U2533 ( .B1(n2036), .B2(n2270), .A(n4840), .ZN(n2152) );
  AND2_X1 U2534 ( .A1(n2072), .A2(n2017), .ZN(n2508) );
  OR2_X1 U2535 ( .A1(n4828), .A2(n3971), .ZN(n4840) );
  NAND2_X1 U2536 ( .A1(n2343), .A2(n2840), .ZN(n4585) );
  NAND2_X1 U2537 ( .A1(n2167), .A2(n2169), .ZN(n3071) );
  AND2_X1 U2538 ( .A1(n2208), .A2(n2806), .ZN(n2168) );
  NAND2_X1 U2539 ( .A1(n4416), .A2(n3081), .ZN(n3082) );
  AND2_X1 U2540 ( .A1(n3080), .A2(n2352), .ZN(n3081) );
  XNOR2_X1 U2541 ( .A(n2410), .B(IR_REG_9__SCAN_IN), .ZN(n4817) );
  INV_X1 U2542 ( .A(IR_REG_8__SCAN_IN), .ZN(n2405) );
  NOR2_X1 U2543 ( .A1(n3895), .A2(n2218), .ZN(n2217) );
  INV_X1 U2544 ( .A(n3938), .ZN(n2218) );
  NOR2_X1 U2545 ( .A1(n3794), .A2(n3795), .ZN(n2125) );
  NOR2_X1 U2546 ( .A1(n4157), .A2(n2288), .ZN(n2287) );
  INV_X1 U2547 ( .A(n3789), .ZN(n3745) );
  NOR2_X1 U2548 ( .A1(n4115), .A2(n4117), .ZN(n4185) );
  NAND2_X1 U2549 ( .A1(n3128), .A2(n2393), .ZN(n2396) );
  NOR2_X1 U2550 ( .A1(n2081), .A2(n2080), .ZN(n2077) );
  NAND2_X1 U2551 ( .A1(n2079), .A2(n2494), .ZN(n2078) );
  NOR2_X1 U2552 ( .A1(n2053), .A2(n2100), .ZN(n2099) );
  INV_X1 U2553 ( .A(n2107), .ZN(n2103) );
  NOR2_X1 U2554 ( .A1(n2350), .A2(n3524), .ZN(n2098) );
  NAND2_X1 U2555 ( .A1(n2144), .A2(n2142), .ZN(n2416) );
  INV_X1 U2556 ( .A(n2143), .ZN(n2142) );
  OAI21_X1 U2557 ( .B1(n2408), .B2(n2147), .A(n2411), .ZN(n2143) );
  INV_X1 U2558 ( .A(n3688), .ZN(n2255) );
  INV_X1 U2559 ( .A(n4836), .ZN(n2095) );
  INV_X1 U2560 ( .A(n4349), .ZN(n2239) );
  AND2_X1 U2561 ( .A1(n2645), .A2(REG2_REG_15__SCAN_IN), .ZN(n2257) );
  NOR2_X1 U2562 ( .A1(n2476), .A2(IR_REG_25__SCAN_IN), .ZN(n2278) );
  XNOR2_X1 U2563 ( .A(IR_REG_28__SCAN_IN), .B(IR_REG_27__SCAN_IN), .ZN(n2474)
         );
  AND2_X1 U2564 ( .A1(n2481), .A2(IR_REG_31__SCAN_IN), .ZN(n2277) );
  NOR2_X1 U2565 ( .A1(n2752), .A2(n2751), .ZN(n2060) );
  INV_X1 U2566 ( .A(n2842), .ZN(n2160) );
  NOR2_X1 U2567 ( .A1(n2679), .A2(n2667), .ZN(n2063) );
  AND2_X1 U2568 ( .A1(n2841), .A2(n2840), .ZN(n2342) );
  INV_X1 U2569 ( .A(n4588), .ZN(n2841) );
  NAND2_X1 U2570 ( .A1(n2654), .A2(n2653), .ZN(n2677) );
  NOR2_X1 U2571 ( .A1(n3854), .A2(n2206), .ZN(n2205) );
  INV_X1 U2572 ( .A(n3851), .ZN(n2206) );
  AOI21_X1 U2573 ( .B1(n3816), .B2(n2203), .A(n3911), .ZN(n2202) );
  INV_X1 U2574 ( .A(n2205), .ZN(n2203) );
  INV_X1 U2575 ( .A(n3816), .ZN(n2204) );
  NOR2_X1 U2576 ( .A1(n2569), .A2(n2059), .ZN(n2577) );
  NAND2_X1 U2577 ( .A1(n2562), .A2(n3832), .ZN(n2213) );
  NOR2_X1 U2578 ( .A1(n3833), .A2(n2216), .ZN(n2215) );
  INV_X1 U2579 ( .A(n3894), .ZN(n2155) );
  INV_X1 U2580 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3041) );
  AND2_X1 U2581 ( .A1(n4472), .A2(n2018), .ZN(n2897) );
  NOR2_X1 U2582 ( .A1(n2190), .A2(n4109), .ZN(n2189) );
  INV_X1 U2583 ( .A(n2191), .ZN(n2190) );
  NOR2_X1 U2584 ( .A1(n4655), .A2(n4442), .ZN(n2191) );
  NAND2_X1 U2585 ( .A1(n2583), .A2(n2582), .ZN(n2585) );
  NAND2_X1 U2586 ( .A1(n3554), .A2(n2561), .ZN(n2179) );
  INV_X1 U2587 ( .A(n2899), .ZN(n3457) );
  INV_X1 U2588 ( .A(IR_REG_23__SCAN_IN), .ZN(n2453) );
  INV_X1 U2589 ( .A(IR_REG_15__SCAN_IN), .ZN(n2363) );
  INV_X1 U2590 ( .A(IR_REG_10__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U2591 ( .A1(n3481), .A2(n3480), .ZN(n2303) );
  INV_X1 U2592 ( .A(n2302), .ZN(n2301) );
  NAND2_X1 U2593 ( .A1(n2060), .A2(REG3_REG_27__SCAN_IN), .ZN(n2773) );
  AND2_X1 U2594 ( .A1(n4003), .A2(n4004), .ZN(n4117) );
  NAND2_X1 U2595 ( .A1(n2062), .A2(n2052), .ZN(n2627) );
  INV_X1 U2596 ( .A(n2620), .ZN(n2062) );
  NAND2_X1 U2597 ( .A1(n3794), .A2(n3795), .ZN(n2126) );
  NOR2_X1 U2598 ( .A1(n2280), .A2(n2125), .ZN(n2124) );
  INV_X1 U2599 ( .A(n2125), .ZN(n2122) );
  AND2_X1 U2600 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2563) );
  NAND2_X1 U2601 ( .A1(n2533), .A2(DATAI_4_), .ZN(n2171) );
  NAND2_X1 U2602 ( .A1(n3376), .A2(n3375), .ZN(n2273) );
  INV_X1 U2603 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2597) );
  OR2_X1 U2604 ( .A1(n2598), .A2(n2597), .ZN(n2607) );
  AOI21_X1 U2605 ( .B1(n2287), .B2(n2285), .A(n2284), .ZN(n2283) );
  INV_X1 U2606 ( .A(n4158), .ZN(n2284) );
  OR2_X1 U2607 ( .A1(n3182), .A2(n3181), .ZN(n3255) );
  NAND2_X1 U2608 ( .A1(n2584), .A2(REG1_REG_1__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U2609 ( .A1(n2914), .A2(REG0_REG_1__SCAN_IN), .ZN(n2336) );
  INV_X1 U2610 ( .A(n2091), .ZN(n2088) );
  NAND2_X1 U2611 ( .A1(n2085), .A2(n2083), .ZN(n2488) );
  NAND2_X1 U2612 ( .A1(n2089), .A2(n2086), .ZN(n2085) );
  NOR2_X1 U2613 ( .A1(n2091), .A2(n2487), .ZN(n2086) );
  NAND2_X1 U2614 ( .A1(n2490), .A2(n2223), .ZN(n2222) );
  INV_X1 U2615 ( .A(n3127), .ZN(n2223) );
  OR2_X1 U2616 ( .A1(n3292), .A2(n2047), .ZN(n2224) );
  NOR2_X1 U2617 ( .A1(n2251), .A2(n2247), .ZN(n2246) );
  INV_X1 U2618 ( .A(n3130), .ZN(n2247) );
  XNOR2_X1 U2619 ( .A(n2067), .B(n2251), .ZN(n3138) );
  NOR2_X1 U2620 ( .A1(n2108), .A2(n3524), .ZN(n2107) );
  INV_X1 U2621 ( .A(n2350), .ZN(n2108) );
  OAI21_X1 U2622 ( .B1(n3410), .B2(n2101), .A(n2097), .ZN(n2498) );
  AOI21_X1 U2623 ( .B1(n2104), .B2(REG1_REG_10__SCAN_IN), .A(n4816), .ZN(n2101) );
  AOI21_X1 U2624 ( .B1(n3410), .B2(n2099), .A(n2098), .ZN(n2097) );
  NAND2_X1 U2625 ( .A1(n2105), .A2(n4816), .ZN(n2104) );
  OAI211_X1 U2626 ( .C1(n2066), .C2(n2051), .A(n2500), .B(n2065), .ZN(n2501)
         );
  NAND2_X1 U2627 ( .A1(n2066), .A2(n2227), .ZN(n2065) );
  NAND2_X1 U2628 ( .A1(n2134), .A2(n4812), .ZN(n2133) );
  NAND2_X1 U2629 ( .A1(n2093), .A2(n2092), .ZN(n2505) );
  INV_X1 U2630 ( .A(n2094), .ZN(n2093) );
  OR2_X1 U2631 ( .A1(n4338), .A2(n2055), .ZN(n2092) );
  OAI21_X1 U2632 ( .B1(n2502), .B2(n2095), .A(n2504), .ZN(n2094) );
  XNOR2_X1 U2633 ( .A(n2439), .B(n2652), .ZN(n4843) );
  NOR2_X1 U2634 ( .A1(n2505), .A2(n2652), .ZN(n2506) );
  AND2_X1 U2635 ( .A1(n2770), .A2(n3954), .ZN(n2209) );
  NOR2_X1 U2636 ( .A1(n2325), .A2(n2329), .ZN(n2323) );
  INV_X1 U2637 ( .A(n2354), .ZN(n2329) );
  NAND2_X1 U2638 ( .A1(n2732), .A2(REG3_REG_24__SCAN_IN), .ZN(n2752) );
  INV_X1 U2639 ( .A(n2733), .ZN(n2732) );
  INV_X1 U2640 ( .A(n2060), .ZN(n2762) );
  AOI21_X1 U2641 ( .B1(n2025), .B2(n2198), .A(n2193), .ZN(n2192) );
  INV_X1 U2642 ( .A(n3887), .ZN(n2193) );
  NAND2_X1 U2643 ( .A1(n2331), .A2(n4474), .ZN(n2330) );
  NOR2_X1 U2644 ( .A1(n4513), .A2(n2321), .ZN(n2320) );
  INV_X1 U2645 ( .A(n2847), .ZN(n2321) );
  AND2_X1 U2646 ( .A1(n2684), .A2(n2683), .ZN(n4572) );
  AND2_X1 U2647 ( .A1(n4568), .A2(n4569), .ZN(n4588) );
  NAND2_X1 U2648 ( .A1(n2201), .A2(n3816), .ZN(n3931) );
  NAND2_X1 U2649 ( .A1(n3634), .A2(n2205), .ZN(n2201) );
  OAI21_X1 U2650 ( .B1(n3634), .B2(n2204), .A(n2202), .ZN(n3772) );
  NAND2_X1 U2651 ( .A1(n3634), .A2(n3851), .ZN(n3667) );
  NAND2_X1 U2652 ( .A1(n2154), .A2(n2313), .ZN(n3637) );
  NAND2_X1 U2653 ( .A1(n2043), .A2(n2016), .ZN(n2313) );
  NAND2_X1 U2654 ( .A1(n2829), .A2(n2314), .ZN(n2154) );
  NAND2_X1 U2655 ( .A1(n3637), .A2(n3636), .ZN(n3635) );
  NAND2_X1 U2656 ( .A1(n3194), .A2(n4373), .ZN(n3494) );
  OAI21_X1 U2657 ( .B1(n3571), .B2(n2588), .A(n3839), .ZN(n3424) );
  NAND2_X1 U2658 ( .A1(n2577), .A2(REG3_REG_7__SCAN_IN), .ZN(n2591) );
  CLKBUF_X1 U2659 ( .A(n3302), .Z(n3303) );
  INV_X1 U2660 ( .A(n4419), .ZN(n4109) );
  NAND2_X1 U2661 ( .A1(n4472), .A2(n2191), .ZN(n4444) );
  NAND2_X1 U2662 ( .A1(n4472), .A2(n4456), .ZN(n4455) );
  INV_X1 U2663 ( .A(n4424), .ZN(n4659) );
  AND2_X1 U2664 ( .A1(n2708), .A2(n2707), .ZN(n4686) );
  AND2_X1 U2665 ( .A1(n2187), .A2(n4558), .ZN(n2185) );
  NAND2_X1 U2666 ( .A1(n2186), .A2(n2187), .ZN(n4578) );
  NOR2_X1 U2667 ( .A1(n2175), .A2(n4715), .ZN(n2174) );
  INV_X1 U2668 ( .A(n4723), .ZN(n3991) );
  NAND2_X1 U2669 ( .A1(n2341), .A2(n2340), .ZN(n3695) );
  AND2_X1 U2670 ( .A1(n2341), .A2(n2020), .ZN(n3696) );
  OR2_X1 U2671 ( .A1(n3673), .A2(n2835), .ZN(n2341) );
  NAND2_X1 U2672 ( .A1(n2181), .A2(n3640), .ZN(n2180) );
  INV_X1 U2673 ( .A(n2182), .ZN(n2181) );
  INV_X1 U2674 ( .A(n3756), .ZN(n3640) );
  OR2_X1 U2675 ( .A1(n3506), .A2(n3656), .ZN(n3515) );
  INV_X1 U2676 ( .A(n4306), .ZN(n3653) );
  NOR2_X1 U2677 ( .A1(n3347), .A2(n2177), .ZN(n3565) );
  NAND2_X1 U2678 ( .A1(n2178), .A2(n3595), .ZN(n2177) );
  INV_X1 U2679 ( .A(n2179), .ZN(n2178) );
  INV_X1 U2680 ( .A(n4738), .ZN(n4707) );
  AND2_X1 U2681 ( .A1(n3185), .A2(n3226), .ZN(n4738) );
  OR2_X1 U2682 ( .A1(n3455), .A2(n2807), .ZN(n3363) );
  INV_X1 U2683 ( .A(n2523), .ZN(n2166) );
  INV_X1 U2684 ( .A(IR_REG_18__SCAN_IN), .ZN(n2367) );
  INV_X1 U2685 ( .A(IR_REG_9__SCAN_IN), .ZN(n2413) );
  OR3_X1 U2686 ( .A1(n2409), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2412) );
  NOR2_X1 U2687 ( .A1(n2390), .A2(IR_REG_5__SCAN_IN), .ZN(n2400) );
  INV_X1 U2688 ( .A(IR_REG_3__SCAN_IN), .ZN(n2929) );
  NAND2_X1 U2689 ( .A1(n2379), .A2(IR_REG_31__SCAN_IN), .ZN(n2241) );
  NAND2_X1 U2690 ( .A1(n2116), .A2(n2118), .ZN(n4108) );
  AND2_X1 U2691 ( .A1(n2733), .A2(n2722), .ZN(n4501) );
  OR2_X1 U2692 ( .A1(n3257), .A2(n4043), .ZN(n3258) );
  NAND2_X1 U2693 ( .A1(n4218), .A2(n4161), .ZN(n4164) );
  AND2_X1 U2694 ( .A1(n3806), .A2(n3805), .ZN(n3978) );
  OR2_X1 U2695 ( .A1(n4180), .A2(n2291), .ZN(n2290) );
  AND2_X1 U2696 ( .A1(n4180), .A2(n2298), .ZN(n2294) );
  NAND2_X1 U2697 ( .A1(n4180), .A2(n2293), .ZN(n2292) );
  NAND2_X1 U2698 ( .A1(n3395), .A2(n3394), .ZN(n3437) );
  INV_X1 U2699 ( .A(n2304), .ZN(n4201) );
  AOI21_X1 U2700 ( .B1(n4115), .B2(n2311), .A(n2309), .ZN(n2304) );
  INV_X1 U2701 ( .A(n3534), .ZN(n2276) );
  INV_X1 U2702 ( .A(n4305), .ZN(n3743) );
  NAND2_X1 U2703 ( .A1(n2533), .A2(DATAI_0_), .ZN(n2176) );
  NAND2_X1 U2704 ( .A1(n4160), .A2(n4216), .ZN(n4218) );
  AND3_X1 U2705 ( .A1(n2640), .A2(n2639), .A3(n2638), .ZN(n4231) );
  INV_X1 U2706 ( .A(n4288), .ZN(n4241) );
  NAND2_X1 U2707 ( .A1(n2282), .A2(n2283), .ZN(n4237) );
  INV_X1 U2708 ( .A(n4304), .ZN(n3797) );
  NAND2_X1 U2709 ( .A1(n3208), .A2(n4560), .ZN(n4288) );
  INV_X1 U2710 ( .A(n4291), .ZN(n4262) );
  OR2_X1 U2711 ( .A1(n2309), .A2(n4198), .ZN(n2308) );
  AND2_X1 U2712 ( .A1(n2306), .A2(n4197), .ZN(n2305) );
  OR2_X1 U2713 ( .A1(n2309), .A2(n2307), .ZN(n2306) );
  NAND2_X1 U2714 ( .A1(n3437), .A2(n3436), .ZN(n3482) );
  NOR2_X1 U2715 ( .A1(n2033), .A2(n4076), .ZN(n4275) );
  AND2_X1 U2716 ( .A1(n2651), .A2(n2650), .ZN(n4718) );
  INV_X1 U2717 ( .A(n4438), .ZN(n4301) );
  INV_X1 U2718 ( .A(n4686), .ZN(n4496) );
  NAND2_X1 U2719 ( .A1(n2719), .A2(n2718), .ZN(n4507) );
  NAND2_X1 U2720 ( .A1(n2697), .A2(n2696), .ZN(n4683) );
  OR2_X1 U2721 ( .A1(n4561), .A2(n2782), .ZN(n2697) );
  NAND2_X1 U2722 ( .A1(n2674), .A2(n2673), .ZN(n4593) );
  INV_X1 U2723 ( .A(n4627), .ZN(n4302) );
  OAI211_X1 U2724 ( .C1(n3776), .C2(n2782), .A(n2644), .B(n2643), .ZN(n4303)
         );
  INV_X1 U2725 ( .A(n4231), .ZN(n4716) );
  AOI21_X1 U2726 ( .B1(REG0_REG_5__SCAN_IN), .B2(n2009), .A(n2032), .ZN(n2127)
         );
  NAND2_X1 U2727 ( .A1(n2581), .A2(n4853), .ZN(n2550) );
  NAND2_X1 U2728 ( .A1(n4320), .A2(n2380), .ZN(n4319) );
  AND2_X1 U2729 ( .A1(n2090), .A2(n2087), .ZN(n3236) );
  NAND2_X1 U2730 ( .A1(n2089), .A2(n2088), .ZN(n2090) );
  NAND2_X1 U2731 ( .A1(n3122), .A2(REG1_REG_3__SCAN_IN), .ZN(n3121) );
  OR2_X1 U2732 ( .A1(n3292), .A2(n4910), .ZN(n2226) );
  INV_X1 U2733 ( .A(n2490), .ZN(n2225) );
  NAND2_X1 U2734 ( .A1(n2224), .A2(n2222), .ZN(n3126) );
  NAND2_X1 U2735 ( .A1(n3290), .A2(REG2_REG_4__SCAN_IN), .ZN(n2149) );
  NOR2_X1 U2736 ( .A1(n2024), .A2(n2249), .ZN(n2248) );
  NOR2_X1 U2737 ( .A1(n2019), .A2(n3130), .ZN(n2249) );
  OR2_X1 U2738 ( .A1(n3138), .A2(n3137), .ZN(n3142) );
  AOI21_X1 U2739 ( .B1(n3410), .B2(n2107), .A(n2106), .ZN(n2102) );
  OR2_X1 U2740 ( .A1(n2232), .A2(n2231), .ZN(n4334) );
  OAI21_X1 U2741 ( .B1(n2236), .B2(REG1_REG_12__SCAN_IN), .A(n2233), .ZN(n2232) );
  NOR2_X1 U2742 ( .A1(n3763), .A2(n2236), .ZN(n2231) );
  AND2_X1 U2743 ( .A1(n2064), .A2(n2230), .ZN(n4329) );
  NAND2_X1 U2744 ( .A1(n3763), .A2(REG1_REG_12__SCAN_IN), .ZN(n2230) );
  XNOR2_X1 U2745 ( .A(n2135), .B(n4812), .ZN(n4344) );
  NAND2_X1 U2746 ( .A1(n4344), .A2(REG2_REG_14__SCAN_IN), .ZN(n4343) );
  XNOR2_X1 U2747 ( .A(n2505), .B(n2652), .ZN(n4848) );
  NOR2_X1 U2748 ( .A1(n4848), .A2(REG1_REG_16__SCAN_IN), .ZN(n4849) );
  NAND2_X1 U2749 ( .A1(n2072), .A2(n2237), .ZN(n4348) );
  NAND2_X1 U2750 ( .A1(n2261), .A2(n2259), .ZN(n4363) );
  AOI21_X1 U2751 ( .B1(n2263), .B2(n2484), .A(n2260), .ZN(n2259) );
  AND2_X1 U2752 ( .A1(n2265), .A2(n2441), .ZN(n2260) );
  XNOR2_X1 U2753 ( .A(n4370), .B(n4369), .ZN(n4375) );
  NAND2_X1 U2754 ( .A1(n4367), .A2(n4366), .ZN(n4370) );
  NAND2_X1 U2755 ( .A1(n2210), .A2(n3954), .ZN(n3057) );
  AND2_X1 U2756 ( .A1(n2779), .A2(n2778), .ZN(n4426) );
  OR2_X1 U2757 ( .A1(n4408), .A2(n2782), .ZN(n2779) );
  NAND2_X1 U2758 ( .A1(n2324), .A2(n2322), .ZN(n4432) );
  INV_X1 U2759 ( .A(n2325), .ZN(n2322) );
  NAND2_X1 U2760 ( .A1(n2195), .A2(n3945), .ZN(n4465) );
  NAND2_X1 U2761 ( .A1(n2219), .A2(n3938), .ZN(n4607) );
  CLKBUF_X1 U2762 ( .A(n4634), .Z(n4635) );
  AND4_X1 U2763 ( .A1(n2617), .A2(n2616), .A3(n2615), .A4(n2614), .ZN(n3751)
         );
  NAND2_X1 U2764 ( .A1(n2829), .A2(n2317), .ZN(n2316) );
  INV_X1 U2765 ( .A(n4605), .ZN(n4644) );
  OR2_X1 U2766 ( .A1(n4624), .A2(n4707), .ZN(n4535) );
  OR2_X1 U2767 ( .A1(n4624), .A2(n4741), .ZN(n4617) );
  OAI21_X1 U2768 ( .B1(n3467), .B2(n2562), .A(n3832), .ZN(n3320) );
  INV_X1 U2769 ( .A(n4642), .ZN(n4862) );
  OR2_X1 U2770 ( .A1(n4646), .A2(n3551), .ZN(n4566) );
  INV_X1 U2771 ( .A(n4566), .ZN(n4861) );
  OR2_X1 U2772 ( .A1(n4703), .A2(n4702), .ZN(n4783) );
  INV_X1 U2773 ( .A(IR_REG_29__SCAN_IN), .ZN(n2526) );
  INV_X1 U2774 ( .A(IR_REG_30__SCAN_IN), .ZN(n3093) );
  AND2_X1 U2775 ( .A1(n3246), .A2(STATE_REG_SCAN_IN), .ZN(n4873) );
  MUX2_X1 U2776 ( .A(n2468), .B(IR_REG_31__SCAN_IN), .S(n2467), .Z(n2469) );
  XNOR2_X1 U2777 ( .A(n2424), .B(IR_REG_11__SCAN_IN), .ZN(n4815) );
  XNOR2_X1 U2778 ( .A(n2403), .B(IR_REG_7__SCAN_IN), .ZN(n4818) );
  XNOR2_X1 U2779 ( .A(n2391), .B(IR_REG_5__SCAN_IN), .ZN(n4819) );
  INV_X1 U2780 ( .A(n2552), .ZN(n3119) );
  OAI21_X1 U2781 ( .B1(n2373), .B2(n2375), .A(n2374), .ZN(n2378) );
  NAND2_X1 U2782 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2375)
         );
  BUF_X1 U2783 ( .A(n2486), .Z(n4821) );
  NAND2_X1 U2784 ( .A1(n4106), .A2(n2021), .ZN(n4104) );
  OAI211_X1 U2785 ( .C1(n2493), .C2(n2494), .A(n2076), .B(n2079), .ZN(n3327)
         );
  NAND2_X1 U2786 ( .A1(n2146), .A2(n2408), .ZN(n3404) );
  NAND2_X1 U2787 ( .A1(n4835), .A2(n4836), .ZN(n4834) );
  NAND2_X1 U2788 ( .A1(n2038), .A2(n2150), .ZN(U3258) );
  NAND2_X1 U2789 ( .A1(n2152), .A2(n2151), .ZN(n2150) );
  OR2_X1 U2790 ( .A1(n4746), .A2(n4405), .ZN(n3085) );
  NOR2_X1 U2791 ( .A1(n4907), .A2(n3072), .ZN(n3073) );
  OR2_X1 U2792 ( .A1(n4405), .A2(n4807), .ZN(n3089) );
  INV_X1 U2793 ( .A(n3656), .ZN(n2183) );
  NAND4_X1 U2794 ( .A1(n2162), .A2(n2164), .A3(n2161), .A4(n2454), .ZN(n2015)
         );
  NAND2_X1 U2795 ( .A1(n3741), .A2(n4305), .ZN(n2016) );
  NAND2_X1 U2796 ( .A1(n3738), .A2(n3737), .ZN(n3786) );
  AND2_X1 U2797 ( .A1(n2237), .A2(n2056), .ZN(n2017) );
  NAND2_X1 U2798 ( .A1(n2739), .A2(n2738), .ZN(n4656) );
  OR2_X1 U2799 ( .A1(n3506), .A2(n2180), .ZN(n3633) );
  AND2_X1 U2800 ( .A1(n2189), .A2(n4406), .ZN(n2018) );
  INV_X1 U2801 ( .A(n2484), .ZN(n2266) );
  INV_X1 U2802 ( .A(n3140), .ZN(n2251) );
  OR2_X1 U2803 ( .A1(n4236), .A2(n4125), .ZN(n4077) );
  OR2_X1 U2804 ( .A1(n2250), .A2(n3140), .ZN(n2019) );
  NAND2_X1 U2805 ( .A1(n4736), .A2(n4228), .ZN(n2020) );
  NAND2_X1 U2806 ( .A1(n2131), .A2(n4031), .ZN(n4160) );
  AND3_X1 U2807 ( .A1(n4099), .A2(n4098), .A3(n4250), .ZN(n2021) );
  AND2_X1 U2808 ( .A1(n2470), .A2(n2469), .ZN(n2862) );
  NOR2_X1 U2809 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2373)
         );
  AND2_X1 U2810 ( .A1(n4472), .A2(n2189), .ZN(n2022) );
  AND2_X1 U2811 ( .A1(n2567), .A2(n2568), .ZN(n2023) );
  NAND2_X1 U2812 ( .A1(n2524), .A2(n2455), .ZN(n2447) );
  AND2_X1 U2813 ( .A1(n2250), .A2(n3140), .ZN(n2024) );
  NAND2_X1 U2814 ( .A1(n4587), .A2(n2842), .ZN(n4576) );
  AND2_X1 U2815 ( .A1(n3948), .A2(n2196), .ZN(n2025) );
  AND4_X1 U2816 ( .A1(n3554), .A2(n2561), .A3(n3572), .A4(n3595), .ZN(n2026)
         );
  OR2_X1 U2817 ( .A1(n4176), .A2(n4171), .ZN(n2027) );
  OR3_X1 U2818 ( .A1(n4176), .A2(n4180), .A3(n2295), .ZN(n2028) );
  NOR2_X1 U2819 ( .A1(n3741), .A2(n4305), .ZN(n2029) );
  NAND2_X1 U2820 ( .A1(n2848), .A2(n2847), .ZN(n4512) );
  NOR2_X1 U2821 ( .A1(n4849), .A2(n2506), .ZN(n2030) );
  NAND2_X1 U2822 ( .A1(n3494), .A2(n4079), .ZN(n3282) );
  AND2_X1 U2823 ( .A1(n2345), .A2(n2117), .ZN(n2031) );
  AND2_X1 U2824 ( .A1(n2912), .A2(REG1_REG_5__SCAN_IN), .ZN(n2032) );
  INV_X1 U2825 ( .A(n2119), .ZN(n2118) );
  OAI21_X1 U2826 ( .B1(n2120), .B2(n4273), .A(n4271), .ZN(n2119) );
  AND2_X1 U2827 ( .A1(n4077), .A2(n2345), .ZN(n2033) );
  OAI21_X1 U2828 ( .B1(n4029), .B2(n4028), .A(n4138), .ZN(n4030) );
  NAND2_X1 U2829 ( .A1(n3748), .A2(n2126), .ZN(n2034) );
  AND2_X1 U2830 ( .A1(n3933), .A2(n3938), .ZN(n4637) );
  INV_X1 U2831 ( .A(n2280), .ZN(n2279) );
  NAND2_X1 U2832 ( .A1(n3745), .A2(n3737), .ZN(n2280) );
  AND2_X1 U2833 ( .A1(n4231), .A2(n3991), .ZN(n2035) );
  AND2_X1 U2834 ( .A1(n2269), .A2(n2266), .ZN(n2036) );
  OR2_X1 U2835 ( .A1(n3909), .A2(n3930), .ZN(n2037) );
  AND2_X1 U2836 ( .A1(n2516), .A2(n2515), .ZN(n2038) );
  INV_X1 U2837 ( .A(IR_REG_25__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U2838 ( .A1(n2219), .A2(n2217), .ZN(n2039) );
  AND2_X1 U2839 ( .A1(n2844), .A2(n4579), .ZN(n2040) );
  NAND3_X1 U2840 ( .A1(n2475), .A2(n2474), .A3(n2473), .ZN(n2041) );
  INV_X1 U2841 ( .A(n3944), .ZN(n2197) );
  NAND2_X1 U2842 ( .A1(n2495), .A2(n2494), .ZN(n2042) );
  OR2_X1 U2843 ( .A1(n2029), .A2(n2315), .ZN(n2043) );
  AND2_X1 U2844 ( .A1(n2248), .A2(n2244), .ZN(n2044) );
  AND2_X1 U2845 ( .A1(n3436), .A2(n2303), .ZN(n2045) );
  AND2_X1 U2846 ( .A1(n2281), .A2(n2283), .ZN(n2046) );
  OR2_X1 U2847 ( .A1(n3127), .A2(n4910), .ZN(n2047) );
  AND2_X1 U2848 ( .A1(n2686), .A2(n2217), .ZN(n2048) );
  INV_X1 U2849 ( .A(IR_REG_27__SCAN_IN), .ZN(n2481) );
  INV_X1 U2850 ( .A(IR_REG_14__SCAN_IN), .ZN(n2114) );
  INV_X1 U2851 ( .A(n3741), .ZN(n2184) );
  INV_X1 U2852 ( .A(n4161), .ZN(n2288) );
  XNOR2_X1 U2853 ( .A(n2406), .B(n2405), .ZN(n3330) );
  NOR2_X1 U2854 ( .A1(n4618), .A2(n4704), .ZN(n4596) );
  NOR2_X1 U2855 ( .A1(n3674), .A2(n4228), .ZN(n3675) );
  NOR2_X1 U2856 ( .A1(n3674), .A2(n2175), .ZN(n3700) );
  AND2_X1 U2857 ( .A1(n4516), .A2(n4499), .ZN(n4470) );
  NAND2_X1 U2858 ( .A1(n2555), .A2(n3829), .ZN(n3467) );
  OAI21_X1 U2859 ( .B1(n3410), .B2(n4816), .A(n2102), .ZN(n3520) );
  NAND2_X1 U2860 ( .A1(n2123), .A2(n2121), .ZN(n3979) );
  NAND2_X1 U2861 ( .A1(n2109), .A2(n2300), .ZN(n3530) );
  NAND2_X1 U2862 ( .A1(n3787), .A2(n3748), .ZN(n3796) );
  NAND2_X1 U2863 ( .A1(n3535), .A2(n3534), .ZN(n3646) );
  NAND2_X1 U2864 ( .A1(n2274), .A2(n3648), .ZN(n3733) );
  NAND2_X1 U2865 ( .A1(n2316), .A2(n2319), .ZN(n3511) );
  INV_X1 U2866 ( .A(n4216), .ZN(n2285) );
  NOR2_X1 U2867 ( .A1(n2447), .A2(n2364), .ZN(n2442) );
  INV_X1 U2868 ( .A(n3832), .ZN(n2216) );
  NOR2_X1 U2869 ( .A1(n3506), .A2(n2182), .ZN(n2049) );
  INV_X1 U2870 ( .A(n4143), .ZN(n4579) );
  INV_X1 U2871 ( .A(n4715), .ZN(n3779) );
  INV_X1 U2872 ( .A(n4620), .ZN(n4704) );
  AND2_X1 U2873 ( .A1(n4139), .A2(n4023), .ZN(n2050) );
  OR2_X1 U2874 ( .A1(n3767), .A2(n2229), .ZN(n2051) );
  INV_X1 U2875 ( .A(n4618), .ZN(n2186) );
  INV_X1 U2876 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2059) );
  AND2_X1 U2877 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .ZN(
        n2052) );
  NAND2_X1 U2878 ( .A1(n3738), .A2(n2279), .ZN(n3787) );
  XNOR2_X1 U2879 ( .A(n2501), .B(n4812), .ZN(n4338) );
  AND2_X1 U2880 ( .A1(n2103), .A2(n2105), .ZN(n2053) );
  INV_X1 U2881 ( .A(n2080), .ZN(n2079) );
  NOR2_X1 U2882 ( .A1(n2349), .A2(n2494), .ZN(n2080) );
  AND2_X1 U2883 ( .A1(n4819), .A2(REG1_REG_5__SCAN_IN), .ZN(n2054) );
  AOI21_X1 U2884 ( .B1(n3424), .B2(n3841), .A(n3423), .ZN(n3503) );
  XNOR2_X1 U2885 ( .A(n2426), .B(IR_REG_12__SCAN_IN), .ZN(n4814) );
  OR2_X1 U2886 ( .A1(n2095), .A2(n4731), .ZN(n2055) );
  INV_X1 U2887 ( .A(n2064), .ZN(n2236) );
  AND2_X2 U2888 ( .A1(n2922), .A2(n3180), .ZN(n4915) );
  NAND2_X1 U2889 ( .A1(n3259), .A2(n3258), .ZN(n4151) );
  NOR2_X1 U2890 ( .A1(n3347), .A2(n2179), .ZN(n3311) );
  NOR2_X1 U2891 ( .A1(n3173), .A2(n2013), .ZN(n3348) );
  OR2_X1 U2892 ( .A1(n4356), .A2(REG1_REG_17__SCAN_IN), .ZN(n2056) );
  NAND2_X1 U2893 ( .A1(n2273), .A2(n3380), .ZN(n3416) );
  AND2_X1 U2894 ( .A1(n2239), .A2(n2238), .ZN(n2057) );
  INV_X1 U2895 ( .A(n2106), .ZN(n2105) );
  NOR2_X1 U2896 ( .A1(n2350), .A2(n4816), .ZN(n2106) );
  INV_X1 U2897 ( .A(n2268), .ZN(n2267) );
  NAND2_X1 U2898 ( .A1(n4362), .A2(REG2_REG_18__SCAN_IN), .ZN(n2268) );
  AND2_X1 U2899 ( .A1(n2226), .A2(n2225), .ZN(n2058) );
  INV_X1 U2900 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2100) );
  INV_X1 U2901 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2238) );
  INV_X1 U2902 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2235) );
  NAND2_X2 U2903 ( .A1(n2613), .A2(n3849), .ZN(n3634) );
  NAND2_X1 U2904 ( .A1(n2219), .A2(n2048), .ZN(n4546) );
  NAND2_X1 U2905 ( .A1(n2590), .A2(REG3_REG_8__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U2906 ( .A1(n2194), .A2(n2192), .ZN(n4451) );
  OAI22_X1 U2907 ( .A1(n3959), .A2(n3958), .B1(n3961), .B2(n3960), .ZN(n3966)
         );
  NAND2_X1 U2908 ( .A1(n3880), .A2(n3951), .ZN(n3958) );
  NAND2_X1 U2909 ( .A1(n3945), .A2(n2197), .ZN(n2196) );
  NAND2_X1 U2910 ( .A1(n2339), .A2(n2338), .ZN(n3775) );
  NAND2_X1 U2911 ( .A1(n2153), .A2(n2837), .ZN(n4633) );
  NAND2_X2 U2912 ( .A1(n2853), .A2(n2852), .ZN(n4468) );
  NAND2_X1 U2913 ( .A1(n2525), .A2(n2524), .ZN(n2528) );
  NAND2_X1 U2914 ( .A1(n2157), .A2(n2156), .ZN(n4543) );
  NAND2_X1 U2915 ( .A1(n2815), .A2(n2155), .ZN(n3302) );
  NAND2_X1 U2916 ( .A1(n2066), .A2(n4814), .ZN(n2064) );
  XNOR2_X1 U2917 ( .A(n2066), .B(n3767), .ZN(n3763) );
  NAND2_X1 U2918 ( .A1(n2493), .A2(n2349), .ZN(n2495) );
  OAI211_X1 U2919 ( .C1(n2493), .C2(n2078), .A(n2075), .B(REG1_REG_8__SCAN_IN), 
        .ZN(n2074) );
  NAND2_X1 U2920 ( .A1(n2493), .A2(n2077), .ZN(n2075) );
  NAND2_X1 U2921 ( .A1(n2084), .A2(n3237), .ZN(n2083) );
  INV_X1 U2922 ( .A(n2090), .ZN(n3238) );
  NOR2_X1 U2923 ( .A1(n4315), .A2(n4316), .ZN(n4314) );
  INV_X1 U2924 ( .A(n2498), .ZN(n3686) );
  AND2_X1 U2925 ( .A1(n2301), .A2(n3394), .ZN(n2110) );
  NAND2_X1 U2926 ( .A1(n2454), .A2(n2344), .ZN(n2523) );
  INV_X1 U2927 ( .A(n2454), .ZN(n2452) );
  INV_X1 U2928 ( .A(n4076), .ZN(n2120) );
  NAND2_X1 U2929 ( .A1(n3738), .A2(n2124), .ZN(n2123) );
  INV_X1 U2930 ( .A(n3383), .ZN(n2129) );
  INV_X2 U2931 ( .A(n4309), .ZN(n3596) );
  AND2_X2 U2932 ( .A1(n2282), .A2(n2046), .ZN(n4236) );
  XNOR2_X2 U2933 ( .A(n2132), .B(n3093), .ZN(n2531) );
  NAND2_X1 U2934 ( .A1(n4343), .A2(n2133), .ZN(n2435) );
  INV_X1 U2935 ( .A(n2135), .ZN(n2134) );
  NAND2_X2 U2936 ( .A1(n4842), .A2(n2440), .ZN(n4351) );
  NAND2_X1 U2937 ( .A1(n4843), .A2(n4841), .ZN(n4842) );
  NAND2_X1 U2938 ( .A1(n3687), .A2(n2422), .ZN(n2136) );
  NAND2_X1 U2939 ( .A1(n2136), .A2(n3767), .ZN(n2140) );
  NAND2_X1 U2940 ( .A1(n3687), .A2(n2422), .ZN(n2141) );
  NAND2_X1 U2941 ( .A1(n3687), .A2(n2138), .ZN(n2137) );
  INV_X1 U2942 ( .A(n2422), .ZN(n2139) );
  NAND2_X1 U2943 ( .A1(n2141), .A2(n4814), .ZN(n2427) );
  NAND2_X1 U2944 ( .A1(n3328), .A2(n2145), .ZN(n2144) );
  NAND2_X2 U2945 ( .A1(n2149), .A2(n2389), .ZN(n3129) );
  OR2_X2 U2946 ( .A1(n4633), .A2(n4637), .ZN(n4634) );
  AND2_X2 U2947 ( .A1(n3832), .A2(n3830), .ZN(n3894) );
  NAND2_X1 U2948 ( .A1(n2343), .A2(n2158), .ZN(n2157) );
  NAND4_X1 U2949 ( .A1(n2358), .A2(n2359), .A3(n2361), .A4(n2360), .ZN(n2165)
         );
  INV_X1 U2950 ( .A(n2165), .ZN(n2163) );
  NAND3_X1 U2951 ( .A1(n2868), .A2(n2869), .A3(n2170), .ZN(n2169) );
  NAND2_X2 U2952 ( .A1(n2015), .A2(n2172), .ZN(n2533) );
  AOI21_X2 U2953 ( .B1(n2477), .B2(n2277), .A(n2041), .ZN(n2172) );
  INV_X1 U2954 ( .A(n3674), .ZN(n2173) );
  NAND2_X1 U2955 ( .A1(n2173), .A2(n2174), .ZN(n4638) );
  INV_X1 U2956 ( .A(n4638), .ZN(n2895) );
  OAI21_X1 U2957 ( .B1(n2533), .B2(n2333), .A(n2176), .ZN(n3456) );
  NAND2_X1 U2958 ( .A1(n2892), .A2(n2026), .ZN(n3566) );
  NAND2_X1 U2959 ( .A1(n2892), .A2(n2561), .ZN(n3466) );
  INV_X1 U2960 ( .A(n3633), .ZN(n2894) );
  NAND2_X1 U2961 ( .A1(n2186), .A2(n2185), .ZN(n4557) );
  NAND2_X1 U2962 ( .A1(n4485), .A2(n2025), .ZN(n2194) );
  NAND2_X1 U2963 ( .A1(n3634), .A2(n2202), .ZN(n2199) );
  NAND2_X1 U2964 ( .A1(n2199), .A2(n2200), .ZN(n2646) );
  NAND2_X1 U2965 ( .A1(n2801), .A2(n4590), .ZN(n2207) );
  NAND2_X1 U2966 ( .A1(n2207), .A2(n2806), .ZN(n4400) );
  INV_X1 U2967 ( .A(n2810), .ZN(n2208) );
  NAND2_X1 U2968 ( .A1(n2210), .A2(n2209), .ZN(n2771) );
  NAND2_X1 U2969 ( .A1(n4626), .A2(n4637), .ZN(n2219) );
  INV_X1 U2970 ( .A(n4149), .ZN(n3196) );
  NAND2_X1 U2971 ( .A1(n2646), .A2(n3818), .ZN(n4626) );
  NAND2_X1 U2972 ( .A1(n2221), .A2(n2220), .ZN(n3410) );
  INV_X1 U2973 ( .A(n2226), .ZN(n3291) );
  NAND2_X1 U2974 ( .A1(n2506), .A2(n2239), .ZN(n2237) );
  XNOR2_X2 U2975 ( .A(n2407), .B(n3330), .ZN(n3328) );
  NAND2_X2 U2976 ( .A1(n3216), .A2(n2401), .ZN(n2407) );
  NAND2_X1 U2977 ( .A1(n3218), .A2(n3217), .ZN(n3216) );
  NAND2_X1 U2978 ( .A1(n3118), .A2(REG2_REG_3__SCAN_IN), .ZN(n2240) );
  MUX2_X1 U2979 ( .A(REG2_REG_1__SCAN_IN), .B(n3496), .S(n2486), .Z(n4320) );
  XNOR2_X2 U2980 ( .A(n2241), .B(IR_REG_1__SCAN_IN), .ZN(n2486) );
  OAI211_X1 U2981 ( .C1(n3129), .C2(n2245), .A(n2242), .B(REG2_REG_6__SCAN_IN), 
        .ZN(n2398) );
  NAND2_X1 U2982 ( .A1(n2044), .A2(n3129), .ZN(n2242) );
  NAND2_X1 U2983 ( .A1(n3129), .A2(n3130), .ZN(n3128) );
  OAI211_X1 U2984 ( .C1(n3129), .C2(n2019), .A(n2248), .B(n2243), .ZN(n3136)
         );
  NAND2_X1 U2985 ( .A1(n3129), .A2(n2246), .ZN(n2243) );
  NAND2_X1 U2986 ( .A1(n2248), .A2(n2019), .ZN(n2245) );
  OAI21_X2 U2987 ( .B1(n3521), .B2(n2253), .A(n2252), .ZN(n3687) );
  AOI21_X2 U2988 ( .B1(n2417), .B2(n2256), .A(n2255), .ZN(n2252) );
  INV_X1 U2989 ( .A(n2417), .ZN(n2253) );
  NAND2_X1 U2990 ( .A1(n2254), .A2(n2417), .ZN(n3689) );
  NAND2_X1 U2991 ( .A1(n3521), .A2(REG2_REG_10__SCAN_IN), .ZN(n2254) );
  INV_X1 U2992 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2256) );
  OR2_X1 U2993 ( .A1(n4351), .A2(n2441), .ZN(n2271) );
  NAND2_X1 U2994 ( .A1(n4351), .A2(n2262), .ZN(n2261) );
  NAND2_X1 U2995 ( .A1(n4351), .A2(n2441), .ZN(n2269) );
  AND2_X1 U2996 ( .A1(n3386), .A2(n3380), .ZN(n2272) );
  NAND2_X1 U2997 ( .A1(n3535), .A2(n2275), .ZN(n2274) );
  NAND2_X1 U2998 ( .A1(n2477), .A2(IR_REG_31__SCAN_IN), .ZN(n2471) );
  OAI21_X1 U2999 ( .B1(n4176), .B2(n4175), .A(n4174), .ZN(n4208) );
  NAND2_X1 U3000 ( .A1(n2028), .A2(n2289), .ZN(n2299) );
  AOI22_X1 U3001 ( .A1(n4176), .A2(n2294), .B1(n2292), .B2(n2290), .ZN(n2289)
         );
  OAI21_X1 U3002 ( .B1(n2299), .B2(n4296), .A(n4183), .ZN(U3222) );
  OR2_X1 U3003 ( .A1(n2312), .A2(n2867), .ZN(n2868) );
  NAND2_X1 U3004 ( .A1(n2312), .A2(n3077), .ZN(n4390) );
  XNOR2_X2 U3005 ( .A(n2312), .B(n3076), .ZN(n4404) );
  NAND2_X2 U3006 ( .A1(n2861), .A2(n2860), .ZN(n2312) );
  NAND2_X1 U3007 ( .A1(n2829), .A2(n2828), .ZN(n3501) );
  OR2_X1 U3008 ( .A1(n4306), .A2(n3656), .ZN(n2319) );
  NAND2_X1 U3009 ( .A1(n2848), .A2(n2320), .ZN(n4515) );
  NAND2_X1 U3010 ( .A1(n2324), .A2(n2323), .ZN(n3055) );
  INV_X1 U3011 ( .A(n4656), .ZN(n2331) );
  INV_X1 U3012 ( .A(IR_REG_1__SCAN_IN), .ZN(n2332) );
  NOR2_X2 U3013 ( .A1(n2531), .A2(n3097), .ZN(n2576) );
  AND2_X2 U3014 ( .A1(n2531), .A2(n3097), .ZN(n2584) );
  NAND2_X1 U3015 ( .A1(n2576), .A2(REG2_REG_1__SCAN_IN), .ZN(n2335) );
  NAND2_X1 U3016 ( .A1(n3673), .A2(n2340), .ZN(n2339) );
  NAND2_X1 U3017 ( .A1(n2897), .A2(n4394), .ZN(n2910) );
  NAND2_X1 U3018 ( .A1(n2895), .A2(n4639), .ZN(n4618) );
  INV_X1 U3019 ( .A(n2466), .ZN(n2797) );
  NAND2_X1 U3020 ( .A1(n2894), .A2(n2893), .ZN(n3674) );
  NOR2_X1 U3021 ( .A1(n4236), .A2(n4125), .ZN(n4176) );
  NAND2_X1 U3022 ( .A1(n3567), .A2(n3623), .ZN(n3506) );
  INV_X1 U3023 ( .A(n3347), .ZN(n2892) );
  NOR2_X1 U3024 ( .A1(n3272), .A2(n3271), .ZN(n3273) );
  CLKBUF_X1 U3025 ( .A(n4150), .Z(n4153) );
  INV_X1 U3026 ( .A(n4517), .ZN(n4530) );
  OR2_X1 U3027 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  INV_X1 U3028 ( .A(n3260), .ZN(n3211) );
  AND2_X1 U3029 ( .A1(n2900), .A2(n3457), .ZN(n3194) );
  INV_X1 U3030 ( .A(n2900), .ZN(n4811) );
  AND2_X1 U3031 ( .A1(n3055), .A2(n3886), .ZN(n3056) );
  INV_X1 U3032 ( .A(n3097), .ZN(n2530) );
  AND2_X1 U3033 ( .A1(n2871), .A2(n2453), .ZN(n2344) );
  AND2_X1 U3034 ( .A1(n4071), .A2(n4070), .ZN(n2345) );
  AND2_X1 U3035 ( .A1(n2114), .A2(n2362), .ZN(n2346) );
  AND2_X1 U3036 ( .A1(n2797), .A2(n2796), .ZN(n2348) );
  OAI21_X1 U3037 ( .B1(n3979), .B2(n3978), .A(n3977), .ZN(n4224) );
  OR2_X1 U3038 ( .A1(n3221), .A2(n4913), .ZN(n2349) );
  OR2_X1 U3039 ( .A1(n3408), .A2(n2496), .ZN(n2350) );
  OR2_X1 U3040 ( .A1(n3692), .A2(n2991), .ZN(n2351) );
  OR2_X1 U3041 ( .A1(n4409), .A2(n4726), .ZN(n2352) );
  INV_X1 U3042 ( .A(DATAI_0_), .ZN(n2540) );
  INV_X1 U3043 ( .A(DATAI_3_), .ZN(n2554) );
  AND4_X1 U3044 ( .A1(n3076), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n2353)
         );
  NAND2_X1 U3045 ( .A1(n4424), .A2(n4442), .ZN(n2354) );
  AND2_X1 U3046 ( .A1(n4473), .A2(n4456), .ZN(n3925) );
  INV_X1 U3047 ( .A(n3925), .ZN(n2748) );
  INV_X1 U3048 ( .A(n4398), .ZN(n2902) );
  INV_X1 U3049 ( .A(n3077), .ZN(n3076) );
  AND2_X1 U3050 ( .A1(n2584), .A2(REG1_REG_7__SCAN_IN), .ZN(n2355) );
  AND2_X2 U3051 ( .A1(n2922), .A2(n3453), .ZN(n4907) );
  INV_X1 U3052 ( .A(n4746), .ZN(n2901) );
  INV_X1 U3053 ( .A(n3304), .ZN(n2816) );
  OR2_X1 U3054 ( .A1(n4259), .A2(n4258), .ZN(n4023) );
  INV_X1 U3055 ( .A(n3936), .ZN(n2686) );
  INV_X1 U3056 ( .A(n4030), .ZN(n4031) );
  OAI21_X1 U3057 ( .B1(n3165), .B2(n3383), .A(n3276), .ZN(n3277) );
  INV_X1 U3058 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2635) );
  AND2_X1 U3059 ( .A1(n2760), .A2(n4433), .ZN(n3952) );
  NAND2_X1 U3060 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2792) );
  INV_X1 U3061 ( .A(n2591), .ZN(n2590) );
  OR2_X1 U3062 ( .A1(n3805), .A2(n3806), .ZN(n3977) );
  INV_X1 U3063 ( .A(n3419), .ZN(n3386) );
  INV_X1 U3064 ( .A(n2913), .ZN(n2785) );
  AOI21_X1 U3065 ( .B1(n4846), .B2(ADDR_REG_18__SCAN_IN), .A(n4263), .ZN(n2513) );
  OR2_X1 U3066 ( .A1(n4239), .A2(n2782), .ZN(n2708) );
  INV_X1 U3067 ( .A(n4518), .ZN(n2896) );
  INV_X1 U3068 ( .A(n3801), .ZN(n2893) );
  INV_X1 U3069 ( .A(n3623), .ZN(n3536) );
  NAND2_X1 U3070 ( .A1(n2011), .A2(n2552), .ZN(n2553) );
  AND2_X1 U3071 ( .A1(n2489), .A2(n4820), .ZN(n2490) );
  OAI21_X1 U3072 ( .B1(n4852), .B2(n4875), .A(n2513), .ZN(n2514) );
  INV_X1 U3073 ( .A(n4382), .ZN(n2911) );
  OR2_X1 U3074 ( .A1(n3926), .A2(n3925), .ZN(n4454) );
  AND2_X1 U3075 ( .A1(n4489), .A2(n2849), .ZN(n4513) );
  NAND2_X1 U3076 ( .A1(n3823), .A2(n3827), .ZN(n3354) );
  OAI21_X1 U3077 ( .B1(n4382), .B2(n4741), .A(n4383), .ZN(n2919) );
  AND2_X1 U3078 ( .A1(n4555), .A2(n3363), .ZN(n4678) );
  XNOR2_X1 U3079 ( .A(n4063), .B(n4087), .ZN(n4209) );
  INV_X1 U3080 ( .A(n4267), .ZN(n4287) );
  OR2_X1 U3081 ( .A1(n4476), .A2(n2782), .ZN(n2739) );
  AND2_X1 U3082 ( .A1(n2663), .A2(n2662), .ZN(n4627) );
  INV_X1 U3083 ( .A(n3751), .ZN(n4739) );
  OR2_X1 U3084 ( .A1(n2899), .A2(n2900), .ZN(n4741) );
  INV_X1 U3085 ( .A(n4859), .ZN(n4560) );
  INV_X1 U3086 ( .A(n4535), .ZN(n4612) );
  INV_X1 U3087 ( .A(n4624), .ZN(n4556) );
  INV_X1 U3088 ( .A(n2919), .ZN(n2920) );
  INV_X1 U3089 ( .A(n4741), .ZN(n4724) );
  NAND2_X1 U3090 ( .A1(n2800), .A2(n2799), .ZN(n4590) );
  INV_X1 U3091 ( .A(n3363), .ZN(n4896) );
  INV_X1 U3092 ( .A(n3180), .ZN(n3453) );
  OR2_X1 U3093 ( .A1(n2431), .A2(n2430), .ZN(n4332) );
  XNOR2_X1 U3094 ( .A(n2395), .B(n2399), .ZN(n3140) );
  AND2_X1 U3095 ( .A1(n2512), .A2(n2511), .ZN(n4846) );
  AND2_X1 U3096 ( .A1(n3250), .A2(n3249), .ZN(n4276) );
  OR2_X1 U3097 ( .A1(n3251), .A2(n3226), .ZN(n4291) );
  OR3_X1 U3098 ( .A1(n3206), .A2(n3449), .A3(n3193), .ZN(n4296) );
  NAND2_X1 U3099 ( .A1(n2746), .A2(n2745), .ZN(n4473) );
  INV_X1 U3100 ( .A(n4572), .ZN(n4705) );
  OR2_X1 U3101 ( .A1(n4828), .A2(n3226), .ZN(n4852) );
  AND2_X1 U3102 ( .A1(n3454), .A2(n4560), .ZN(n4624) );
  OR2_X1 U3103 ( .A1(n4624), .A2(n3552), .ZN(n4605) );
  AND2_X1 U3104 ( .A1(n2905), .A2(n2904), .ZN(n2906) );
  NAND2_X1 U3105 ( .A1(n4915), .A2(n4597), .ZN(n4746) );
  AOI21_X1 U3106 ( .B1(n2902), .B2(n4889), .A(n3073), .ZN(n3074) );
  NAND2_X1 U3107 ( .A1(n4907), .A2(n4597), .ZN(n4807) );
  INV_X1 U3108 ( .A(n4907), .ZN(n4905) );
  XNOR2_X1 U3109 ( .A(n2872), .B(n2871), .ZN(n3113) );
  INV_X1 U3110 ( .A(n2531), .ZN(n4809) );
  INV_X1 U3111 ( .A(n4332), .ZN(n4813) );
  INV_X2 U3112 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U3113 ( .A1(n2442), .A2(n2444), .ZN(n2366) );
  NAND2_X1 U3114 ( .A1(n2366), .A2(IR_REG_31__SCAN_IN), .ZN(n2365) );
  MUX2_X1 U3115 ( .A(IR_REG_31__SCAN_IN), .B(n2365), .S(IR_REG_18__SCAN_IN), 
        .Z(n2369) );
  INV_X1 U3116 ( .A(n2366), .ZN(n2368) );
  NAND2_X1 U3117 ( .A1(n2368), .A2(n2367), .ZN(n2791) );
  NAND2_X1 U3118 ( .A1(n2369), .A2(n2791), .ZN(n4875) );
  INV_X1 U3119 ( .A(n4875), .ZN(n4362) );
  INV_X1 U3120 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2370) );
  AOI22_X1 U3121 ( .A1(n4362), .A2(n2370), .B1(REG2_REG_18__SCAN_IN), .B2(
        n4875), .ZN(n2484) );
  OR2_X1 U3122 ( .A1(n2447), .A2(IR_REG_14__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3123 ( .A1(n2371), .A2(IR_REG_31__SCAN_IN), .ZN(n2436) );
  XNOR2_X1 U3124 ( .A(n2436), .B(IR_REG_15__SCAN_IN), .ZN(n2645) );
  INV_X1 U3125 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2372) );
  MUX2_X1 U3126 ( .A(REG2_REG_2__SCAN_IN), .B(n2372), .S(n2010), .Z(n3231) );
  INV_X1 U3127 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3496) );
  AND2_X1 U3128 ( .A1(n2379), .A2(REG2_REG_0__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U3129 ( .A1(n4821), .A2(REG2_REG_1__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3130 ( .A1(n4319), .A2(n2381), .ZN(n3230) );
  NAND2_X1 U3131 ( .A1(n3231), .A2(n3230), .ZN(n3232) );
  NAND2_X1 U3132 ( .A1(n2010), .A2(REG2_REG_2__SCAN_IN), .ZN(n2382) );
  NAND2_X1 U3133 ( .A1(n3232), .A2(n2382), .ZN(n2383) );
  NAND2_X1 U3134 ( .A1(n2376), .A2(IR_REG_31__SCAN_IN), .ZN(n2385) );
  XNOR2_X1 U3135 ( .A(n2385), .B(IR_REG_3__SCAN_IN), .ZN(n2552) );
  XNOR2_X2 U3136 ( .A(n2383), .B(n3119), .ZN(n3118) );
  NAND2_X1 U3137 ( .A1(n2383), .A2(n2552), .ZN(n2384) );
  NAND2_X1 U3138 ( .A1(n2385), .A2(n2929), .ZN(n2386) );
  NAND2_X1 U3139 ( .A1(n2386), .A2(IR_REG_31__SCAN_IN), .ZN(n2387) );
  XNOR2_X1 U3140 ( .A(n2387), .B(IR_REG_4__SCAN_IN), .ZN(n4820) );
  INV_X1 U3141 ( .A(n4820), .ZN(n3295) );
  NAND2_X1 U3142 ( .A1(n2388), .A2(n4820), .ZN(n2389) );
  INV_X1 U3143 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2392) );
  NAND2_X1 U3144 ( .A1(n2390), .A2(IR_REG_31__SCAN_IN), .ZN(n2391) );
  MUX2_X1 U3145 ( .A(REG2_REG_5__SCAN_IN), .B(n2392), .S(n4819), .Z(n3130) );
  NAND2_X1 U3146 ( .A1(n4819), .A2(REG2_REG_5__SCAN_IN), .ZN(n2393) );
  INV_X1 U3147 ( .A(n2400), .ZN(n2394) );
  NAND2_X1 U31480 ( .A1(n2394), .A2(IR_REG_31__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U31490 ( .A1(n2396), .A2(n2251), .ZN(n2397) );
  NAND2_X1 U3150 ( .A1(n2398), .A2(n2397), .ZN(n3218) );
  INV_X1 U3151 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2955) );
  NAND2_X1 U3152 ( .A1(n2400), .A2(n2399), .ZN(n2409) );
  NAND2_X1 U3153 ( .A1(n2409), .A2(IR_REG_31__SCAN_IN), .ZN(n2403) );
  MUX2_X1 U3154 ( .A(REG2_REG_7__SCAN_IN), .B(n2955), .S(n4818), .Z(n3217) );
  NAND2_X1 U3155 ( .A1(n4818), .A2(REG2_REG_7__SCAN_IN), .ZN(n2401) );
  INV_X1 U3156 ( .A(IR_REG_7__SCAN_IN), .ZN(n2402) );
  NAND2_X1 U3157 ( .A1(n2403), .A2(n2402), .ZN(n2404) );
  NAND2_X1 U3158 ( .A1(n2404), .A2(IR_REG_31__SCAN_IN), .ZN(n2406) );
  INV_X1 U3159 ( .A(n3330), .ZN(n2494) );
  NAND2_X1 U3160 ( .A1(n2407), .A2(n2494), .ZN(n2408) );
  NAND2_X1 U3161 ( .A1(n2412), .A2(IR_REG_31__SCAN_IN), .ZN(n2410) );
  INV_X1 U3162 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3005) );
  XNOR2_X1 U3163 ( .A(n4817), .B(n3005), .ZN(n3403) );
  NAND2_X1 U3164 ( .A1(n4817), .A2(REG2_REG_9__SCAN_IN), .ZN(n2411) );
  INV_X1 U3165 ( .A(n2412), .ZN(n2414) );
  NAND2_X1 U3166 ( .A1(n2414), .A2(n2413), .ZN(n2418) );
  NAND2_X1 U3167 ( .A1(n2418), .A2(IR_REG_31__SCAN_IN), .ZN(n2415) );
  XNOR2_X1 U3168 ( .A(n2415), .B(IR_REG_10__SCAN_IN), .ZN(n4816) );
  INV_X1 U3169 ( .A(n4816), .ZN(n3524) );
  XNOR2_X1 U3170 ( .A(n2416), .B(n3524), .ZN(n3521) );
  NAND2_X1 U3171 ( .A1(n2416), .A2(n4816), .ZN(n2417) );
  INV_X1 U3172 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2421) );
  INV_X1 U3173 ( .A(n2418), .ZN(n2419) );
  NAND2_X1 U3174 ( .A1(n2419), .A2(n2971), .ZN(n2420) );
  MUX2_X1 U3175 ( .A(REG2_REG_11__SCAN_IN), .B(n2421), .S(n4815), .Z(n3688) );
  NAND2_X1 U3176 ( .A1(n4815), .A2(REG2_REG_11__SCAN_IN), .ZN(n2422) );
  INV_X1 U3177 ( .A(IR_REG_11__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3178 ( .A1(n2424), .A2(n2423), .ZN(n2425) );
  NAND2_X1 U3179 ( .A1(n2425), .A2(IR_REG_31__SCAN_IN), .ZN(n2426) );
  INV_X1 U3180 ( .A(n4814), .ZN(n3767) );
  NAND2_X1 U3181 ( .A1(n3764), .A2(REG2_REG_12__SCAN_IN), .ZN(n2428) );
  NOR2_X1 U3182 ( .A1(n2524), .A2(n2472), .ZN(n2429) );
  MUX2_X1 U3183 ( .A(n2472), .B(n2429), .S(IR_REG_13__SCAN_IN), .Z(n2431) );
  INV_X1 U3184 ( .A(n2447), .ZN(n2430) );
  INV_X1 U3185 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4325) );
  NOR2_X1 U3186 ( .A1(n4332), .A2(n4325), .ZN(n2432) );
  NAND2_X1 U3187 ( .A1(n4332), .A2(n4325), .ZN(n2433) );
  NAND2_X1 U3188 ( .A1(n2447), .A2(IR_REG_31__SCAN_IN), .ZN(n2434) );
  XNOR2_X1 U3189 ( .A(n2434), .B(IR_REG_14__SCAN_IN), .ZN(n4812) );
  INV_X1 U3190 ( .A(n4812), .ZN(n4339) );
  INV_X1 U3191 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2954) );
  INV_X1 U3192 ( .A(n2645), .ZN(n4879) );
  AOI22_X1 U3193 ( .A1(n2645), .A2(n2954), .B1(REG2_REG_15__SCAN_IN), .B2(
        n4879), .ZN(n4830) );
  NAND2_X1 U3194 ( .A1(n2436), .A2(n2363), .ZN(n2437) );
  NAND2_X1 U3195 ( .A1(n2437), .A2(IR_REG_31__SCAN_IN), .ZN(n2438) );
  XNOR2_X1 U3196 ( .A(n2438), .B(IR_REG_16__SCAN_IN), .ZN(n2652) );
  INV_X1 U3197 ( .A(n2652), .ZN(n4877) );
  INV_X1 U3198 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4841) );
  NAND2_X1 U3199 ( .A1(n2439), .A2(n4877), .ZN(n2440) );
  INV_X1 U3200 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2441) );
  INV_X1 U3201 ( .A(n2442), .ZN(n2443) );
  NAND2_X1 U3202 ( .A1(n2443), .A2(IR_REG_31__SCAN_IN), .ZN(n2445) );
  MUX2_X1 U3203 ( .A(n2445), .B(IR_REG_31__SCAN_IN), .S(n2444), .Z(n2446) );
  NAND2_X1 U3204 ( .A1(n2446), .A2(n2366), .ZN(n2665) );
  INV_X1 U3205 ( .A(n2665), .ZN(n4356) );
  NAND2_X1 U3206 ( .A1(n2465), .A2(n2925), .ZN(n2450) );
  NAND2_X1 U3207 ( .A1(n2450), .A2(IR_REG_31__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U3208 ( .A1(n2448), .A2(n2453), .ZN(n2870) );
  OR2_X1 U3209 ( .A1(n2448), .A2(n2453), .ZN(n2449) );
  NAND2_X1 U32100 ( .A1(n2870), .A2(n2449), .ZN(n3246) );
  INV_X1 U32110 ( .A(n2450), .ZN(n2451) );
  NAND2_X1 U32120 ( .A1(n2451), .A2(n2871), .ZN(n2463) );
  NOR2_X1 U32130 ( .A1(n2457), .A2(n2472), .ZN(n2456) );
  INV_X1 U32140 ( .A(n2477), .ZN(n2458) );
  NAND2_X1 U32150 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(
        n2460) );
  NAND2_X1 U32160 ( .A1(n2460), .A2(IR_REG_31__SCAN_IN), .ZN(n2461) );
  OAI21_X1 U32170 ( .B1(n2871), .B2(IR_REG_31__SCAN_IN), .A(n2461), .ZN(n2462)
         );
  NAND2_X1 U32180 ( .A1(n4873), .A2(n3245), .ZN(n3449) );
  OR2_X1 U32190 ( .A1(n3246), .A2(U3149), .ZN(n3975) );
  NAND2_X1 U32200 ( .A1(n3449), .A2(n3975), .ZN(n2511) );
  INV_X1 U32210 ( .A(n2465), .ZN(n2470) );
  NAND2_X1 U32220 ( .A1(n2797), .A2(IR_REG_31__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U32230 ( .A1(n2519), .A2(IR_REG_27__SCAN_IN), .ZN(n2476) );
  NAND3_X1 U32240 ( .A1(n2481), .A2(IR_REG_31__SCAN_IN), .A3(
        IR_REG_26__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U32250 ( .A1(n2472), .A2(IR_REG_27__SCAN_IN), .ZN(n2473) );
  AOI21_X1 U32260 ( .B1(n3185), .B2(n3246), .A(n2011), .ZN(n2510) );
  NAND2_X1 U32270 ( .A1(n2511), .A2(n2510), .ZN(n4828) );
  NAND2_X1 U32280 ( .A1(n2481), .A2(n2519), .ZN(n2478) );
  OAI21_X1 U32290 ( .B1(n2477), .B2(n2478), .A(IR_REG_31__SCAN_IN), .ZN(n2480)
         );
  INV_X1 U32300 ( .A(IR_REG_28__SCAN_IN), .ZN(n2479) );
  XNOR2_X1 U32310 ( .A(n2480), .B(n2479), .ZN(n4822) );
  OAI21_X1 U32320 ( .B1(n2477), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2482) );
  XNOR2_X1 U32330 ( .A(n2482), .B(n2481), .ZN(n4824) );
  OR2_X1 U32340 ( .A1(n4822), .A2(n4824), .ZN(n3971) );
  INV_X1 U32350 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4365) );
  AOI22_X1 U32360 ( .A1(n4362), .A2(REG1_REG_18__SCAN_IN), .B1(n4365), .B2(
        n4875), .ZN(n2509) );
  XNOR2_X1 U32370 ( .A(n2010), .B(REG1_REG_2__SCAN_IN), .ZN(n3237) );
  XNOR2_X1 U32380 ( .A(n2486), .B(REG1_REG_1__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U32390 ( .A1(n2379), .A2(REG1_REG_0__SCAN_IN), .ZN(n4316) );
  XNOR2_X1 U32400 ( .A(n2488), .B(n2552), .ZN(n3122) );
  INV_X1 U32410 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3016) );
  OAI21_X1 U32420 ( .B1(n2488), .B2(n3119), .A(n3121), .ZN(n2489) );
  XNOR2_X1 U32430 ( .A(n2489), .B(n4820), .ZN(n3292) );
  INV_X1 U32440 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4910) );
  INV_X1 U32450 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3373) );
  MUX2_X1 U32460 ( .A(n3373), .B(REG1_REG_5__SCAN_IN), .S(n4819), .Z(n3127) );
  INV_X1 U32470 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3137) );
  INV_X1 U32480 ( .A(n4818), .ZN(n3221) );
  INV_X1 U32490 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4913) );
  INV_X1 U32500 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2496) );
  MUX2_X1 U32510 ( .A(n2496), .B(REG1_REG_9__SCAN_IN), .S(n4817), .Z(n3405) );
  INV_X1 U32520 ( .A(n4817), .ZN(n3408) );
  INV_X1 U32530 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2991) );
  MUX2_X1 U32540 ( .A(n2991), .B(REG1_REG_11__SCAN_IN), .S(n4815), .Z(n3685)
         );
  INV_X1 U32550 ( .A(n4815), .ZN(n3692) );
  INV_X1 U32560 ( .A(REG1_REG_13__SCAN_IN), .ZN(n2499) );
  MUX2_X1 U32570 ( .A(REG1_REG_13__SCAN_IN), .B(n2499), .S(n4332), .Z(n4328)
         );
  NAND2_X1 U32580 ( .A1(n4813), .A2(REG1_REG_13__SCAN_IN), .ZN(n2500) );
  INV_X1 U32590 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U32600 ( .A1(n2501), .A2(n4812), .ZN(n2502) );
  INV_X1 U32610 ( .A(REG1_REG_15__SCAN_IN), .ZN(n2503) );
  AOI22_X1 U32620 ( .A1(n2645), .A2(REG1_REG_15__SCAN_IN), .B1(n2503), .B2(
        n4879), .ZN(n4836) );
  NAND2_X1 U32630 ( .A1(n2645), .A2(REG1_REG_15__SCAN_IN), .ZN(n2504) );
  INV_X1 U32640 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2507) );
  OAI21_X1 U32650 ( .B1(n2507), .B2(n2665), .A(n2056), .ZN(n4349) );
  INV_X1 U32660 ( .A(n4824), .ZN(n4810) );
  INV_X1 U32670 ( .A(n4360), .ZN(n4847) );
  OAI211_X1 U32680 ( .C1(n2509), .C2(n2508), .A(n4847), .B(n4367), .ZN(n2516)
         );
  INV_X1 U32690 ( .A(n4822), .ZN(n3226) );
  INV_X1 U32700 ( .A(n2510), .ZN(n2512) );
  AND2_X1 U32710 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4263) );
  INV_X1 U32720 ( .A(n2514), .ZN(n2515) );
  INV_X1 U32730 ( .A(n2517), .ZN(n2521) );
  NOR2_X1 U32740 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2520) );
  NAND4_X1 U32750 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(n2522)
         );
  INV_X1 U32760 ( .A(n2528), .ZN(n2527) );
  NAND2_X1 U32770 ( .A1(n2527), .A2(n2526), .ZN(n3092) );
  NAND2_X1 U32780 ( .A1(n2528), .A2(IR_REG_31__SCAN_IN), .ZN(n2529) );
  XNOR2_X2 U32790 ( .A(n2529), .B(IR_REG_29__SCAN_IN), .ZN(n3097) );
  INV_X1 U32800 ( .A(DATAI_1_), .ZN(n2535) );
  INV_X1 U32810 ( .A(n4821), .ZN(n2532) );
  OAI21_X2 U32820 ( .B1(n2909), .B2(n2535), .A(n2534), .ZN(n3261) );
  NAND2_X2 U32830 ( .A1(n3824), .A2(n3820), .ZN(n3161) );
  NAND2_X1 U32840 ( .A1(n2581), .A2(REG3_REG_0__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U32850 ( .A1(n2914), .A2(REG0_REG_0__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U32860 ( .A1(n2584), .A2(REG1_REG_0__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U32870 ( .A1(n2576), .A2(REG2_REG_0__SCAN_IN), .ZN(n2536) );
  NAND4_X2 U32880 ( .A1(n2539), .A2(n2538), .A3(n2537), .A4(n2536), .ZN(n4149)
         );
  NAND2_X1 U32890 ( .A1(n3196), .A2(n3456), .ZN(n3819) );
  NAND2_X1 U32900 ( .A1(n2581), .A2(REG3_REG_2__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U32910 ( .A1(n2914), .A2(REG0_REG_2__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U32920 ( .A1(n2584), .A2(REG1_REG_2__SCAN_IN), .ZN(n2542) );
  NAND2_X1 U32930 ( .A1(n2576), .A2(REG2_REG_2__SCAN_IN), .ZN(n2541) );
  INV_X1 U32940 ( .A(DATAI_2_), .ZN(n2546) );
  NAND2_X1 U32950 ( .A1(n3165), .A2(n2013), .ZN(n3823) );
  INV_X1 U32960 ( .A(n4252), .ZN(n2547) );
  NAND2_X1 U32970 ( .A1(n2547), .A2(n4313), .ZN(n3827) );
  NAND2_X1 U32980 ( .A1(n3357), .A2(n3913), .ZN(n3356) );
  NAND2_X1 U32990 ( .A1(n3356), .A2(n3823), .ZN(n3339) );
  NAND2_X1 U33000 ( .A1(n2914), .A2(REG0_REG_3__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U33010 ( .A1(n2584), .A2(REG1_REG_3__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U33020 ( .A1(n3361), .A2(n3340), .ZN(n3829) );
  NAND2_X1 U33030 ( .A1(n3349), .A2(n4311), .ZN(n3826) );
  NAND2_X1 U33040 ( .A1(n3339), .A2(n3912), .ZN(n2555) );
  NAND2_X1 U33050 ( .A1(n2576), .A2(REG2_REG_4__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U33060 ( .A1(n2008), .A2(REG0_REG_4__SCAN_IN), .ZN(n2559) );
  INV_X1 U33070 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2556) );
  XNOR2_X1 U33080 ( .A(n2556), .B(REG3_REG_3__SCAN_IN), .ZN(n3477) );
  NAND2_X1 U33090 ( .A1(n2581), .A2(n3477), .ZN(n2558) );
  NAND2_X1 U33100 ( .A1(n2584), .A2(REG1_REG_4__SCAN_IN), .ZN(n2557) );
  AND4_X2 U33110 ( .A1(n2560), .A2(n2559), .A3(n2558), .A4(n2557), .ZN(n3555)
         );
  NAND2_X1 U33120 ( .A1(n3555), .A2(n3470), .ZN(n3830) );
  INV_X1 U33130 ( .A(n3830), .ZN(n2562) );
  INV_X2 U33140 ( .A(n3555), .ZN(n4310) );
  MUX2_X1 U33150 ( .A(DATAI_5_), .B(n4819), .S(n2909), .Z(n3397) );
  INV_X1 U33160 ( .A(n3397), .ZN(n3554) );
  BUF_X4 U33170 ( .A(n2584), .Z(n2912) );
  INV_X1 U33180 ( .A(n2563), .ZN(n2565) );
  INV_X1 U33190 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U33200 ( .A1(n2565), .A2(n2564), .ZN(n2566) );
  AND2_X1 U33210 ( .A1(n2569), .A2(n2566), .ZN(n3556) );
  NAND2_X1 U33220 ( .A1(n2581), .A2(n3556), .ZN(n2568) );
  NAND2_X1 U33230 ( .A1(n2012), .A2(REG2_REG_5__SCAN_IN), .ZN(n2567) );
  AND2_X1 U33240 ( .A1(n3554), .A2(n4309), .ZN(n3833) );
  NAND2_X1 U33250 ( .A1(n3596), .A2(n3397), .ZN(n3844) );
  INV_X1 U33260 ( .A(DATAI_6_), .ZN(n3099) );
  MUX2_X1 U33270 ( .A(n3099), .B(n3140), .S(n2011), .Z(n3595) );
  NAND2_X1 U33280 ( .A1(n2012), .A2(REG2_REG_6__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U33290 ( .A1(n2009), .A2(REG0_REG_6__SCAN_IN), .ZN(n2573) );
  INV_X1 U33300 ( .A(n2577), .ZN(n2579) );
  NAND2_X1 U33310 ( .A1(n2569), .A2(n2059), .ZN(n2570) );
  AND2_X1 U33320 ( .A1(n2579), .A2(n2570), .ZN(n3592) );
  NAND2_X1 U33330 ( .A1(n2581), .A2(n3592), .ZN(n2572) );
  NAND2_X1 U33340 ( .A1(n2912), .A2(REG1_REG_6__SCAN_IN), .ZN(n2571) );
  AND4_X2 U33350 ( .A1(n2574), .A2(n2573), .A3(n2572), .A4(n2571), .ZN(n3579)
         );
  INV_X1 U33360 ( .A(n3579), .ZN(n4308) );
  NAND2_X1 U33370 ( .A1(n3595), .A2(n4308), .ZN(n3845) );
  NAND2_X1 U33380 ( .A1(n3301), .A2(n3845), .ZN(n2575) );
  INV_X1 U33390 ( .A(n3595), .ZN(n3443) );
  NAND2_X1 U33400 ( .A1(n3579), .A2(n3443), .ZN(n3835) );
  NAND2_X1 U33410 ( .A1(n2576), .A2(REG2_REG_7__SCAN_IN), .ZN(n2583) );
  INV_X1 U33420 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U33430 ( .A1(n2579), .A2(n2578), .ZN(n2580) );
  AND2_X1 U33440 ( .A1(n2591), .A2(n2580), .ZN(n3576) );
  NAND2_X1 U33450 ( .A1(n2581), .A2(n3576), .ZN(n2582) );
  NOR2_X1 U33460 ( .A1(n2585), .A2(n2355), .ZN(n2587) );
  NAND2_X1 U33470 ( .A1(n2914), .A2(REG0_REG_7__SCAN_IN), .ZN(n2586) );
  AND2_X2 U33480 ( .A1(n2587), .A2(n2586), .ZN(n2589) );
  MUX2_X1 U33490 ( .A(DATAI_7_), .B(n4818), .S(n2011), .Z(n3570) );
  NAND2_X1 U33500 ( .A1(n2589), .A2(n3570), .ZN(n2819) );
  INV_X1 U33510 ( .A(n2819), .ZN(n2588) );
  INV_X2 U33520 ( .A(n2589), .ZN(n3599) );
  NAND2_X1 U3353 ( .A1(n2009), .A2(REG0_REG_8__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U33540 ( .A1(n2912), .A2(REG1_REG_8__SCAN_IN), .ZN(n2595) );
  INV_X1 U3355 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2972) );
  NAND2_X1 U3356 ( .A1(n2591), .A2(n2972), .ZN(n2592) );
  AND2_X1 U3357 ( .A1(n2598), .A2(n2592), .ZN(n3625) );
  NAND2_X1 U3358 ( .A1(n2581), .A2(n3625), .ZN(n2594) );
  NAND2_X1 U3359 ( .A1(n2913), .A2(REG2_REG_8__SCAN_IN), .ZN(n2593) );
  INV_X1 U3360 ( .A(DATAI_8_), .ZN(n3103) );
  MUX2_X1 U3361 ( .A(n3103), .B(n3330), .S(n2909), .Z(n3623) );
  NAND2_X1 U3362 ( .A1(n3539), .A2(n3536), .ZN(n3841) );
  AND2_X1 U3363 ( .A1(n3623), .A2(n4307), .ZN(n3423) );
  MUX2_X1 U3364 ( .A(DATAI_9_), .B(n4817), .S(n2011), .Z(n3656) );
  NAND2_X1 U3365 ( .A1(n2913), .A2(REG2_REG_9__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U3366 ( .A1(n2009), .A2(REG0_REG_9__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U3367 ( .A1(n2598), .A2(n2597), .ZN(n2599) );
  AND2_X1 U3368 ( .A1(n2607), .A2(n2599), .ZN(n3660) );
  NAND2_X1 U3369 ( .A1(n2581), .A2(n3660), .ZN(n2601) );
  NAND2_X1 U3370 ( .A1(n2912), .A2(REG1_REG_9__SCAN_IN), .ZN(n2600) );
  NAND4_X1 U3371 ( .A1(n2603), .A2(n2602), .A3(n2601), .A4(n2600), .ZN(n4306)
         );
  NAND2_X1 U3372 ( .A1(n2183), .A2(n4306), .ZN(n3852) );
  NAND2_X1 U3373 ( .A1(n3503), .A2(n3852), .ZN(n2604) );
  NAND2_X1 U3374 ( .A1(n3653), .A2(n3656), .ZN(n3842) );
  NAND2_X1 U3375 ( .A1(n2604), .A2(n3842), .ZN(n3510) );
  MUX2_X1 U3376 ( .A(DATAI_10_), .B(n4816), .S(n2011), .Z(n3741) );
  NAND2_X1 U3377 ( .A1(n2009), .A2(REG0_REG_10__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U3378 ( .A1(n2912), .A2(REG1_REG_10__SCAN_IN), .ZN(n2611) );
  INV_X1 U3379 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U3380 ( .A1(n2607), .A2(n2606), .ZN(n2608) );
  AND2_X1 U3381 ( .A1(n2620), .A2(n2608), .ZN(n3792) );
  NAND2_X1 U3382 ( .A1(n2581), .A2(n3792), .ZN(n2610) );
  NAND2_X1 U3383 ( .A1(n2913), .A2(REG2_REG_10__SCAN_IN), .ZN(n2609) );
  NAND4_X1 U3384 ( .A1(n2612), .A2(n2611), .A3(n2610), .A4(n2609), .ZN(n4305)
         );
  NAND2_X1 U3385 ( .A1(n2184), .A2(n4305), .ZN(n3850) );
  NAND2_X1 U3386 ( .A1(n3510), .A2(n3850), .ZN(n2613) );
  NAND2_X1 U3387 ( .A1(n3743), .A2(n3741), .ZN(n3849) );
  MUX2_X1 U3388 ( .A(DATAI_11_), .B(n4815), .S(n2909), .Z(n3756) );
  NAND2_X1 U3389 ( .A1(n2009), .A2(REG0_REG_11__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U3390 ( .A1(n2912), .A2(REG1_REG_11__SCAN_IN), .ZN(n2616) );
  XNOR2_X1 U3391 ( .A(n2620), .B(REG3_REG_11__SCAN_IN), .ZN(n3760) );
  NAND2_X1 U3392 ( .A1(n2581), .A2(n3760), .ZN(n2615) );
  NAND2_X1 U3393 ( .A1(n2913), .A2(REG2_REG_11__SCAN_IN), .ZN(n2614) );
  NAND2_X1 U3394 ( .A1(n3640), .A2(n4739), .ZN(n3851) );
  MUX2_X1 U3395 ( .A(DATAI_12_), .B(n4814), .S(n2011), .Z(n3801) );
  NAND2_X1 U3396 ( .A1(n2913), .A2(REG2_REG_12__SCAN_IN), .ZN(n2625) );
  INV_X1 U3397 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2619) );
  INV_X1 U3398 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2618) );
  OAI21_X1 U3399 ( .B1(n2620), .B2(n2619), .A(n2618), .ZN(n2621) );
  AND2_X1 U3400 ( .A1(n2621), .A2(n2627), .ZN(n3812) );
  NAND2_X1 U3401 ( .A1(n2581), .A2(n3812), .ZN(n2624) );
  NAND2_X1 U3402 ( .A1(n2009), .A2(REG0_REG_12__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U3403 ( .A1(n2912), .A2(REG1_REG_12__SCAN_IN), .ZN(n2622) );
  NAND4_X1 U3404 ( .A1(n2625), .A2(n2624), .A3(n2623), .A4(n2622), .ZN(n4304)
         );
  NAND2_X1 U3405 ( .A1(n2893), .A2(n4304), .ZN(n3722) );
  INV_X1 U3406 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2626) );
  NAND2_X1 U3407 ( .A1(n2627), .A2(n2626), .ZN(n2628) );
  NAND2_X1 U3408 ( .A1(n2636), .A2(n2628), .ZN(n3678) );
  OR2_X1 U3409 ( .A1(n3678), .A2(n2782), .ZN(n2632) );
  NAND2_X1 U3410 ( .A1(n2913), .A2(REG2_REG_13__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3411 ( .A1(n2009), .A2(REG0_REG_13__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U3412 ( .A1(n2912), .A2(REG1_REG_13__SCAN_IN), .ZN(n2629) );
  MUX2_X1 U3413 ( .A(DATAI_13_), .B(n4813), .S(n2011), .Z(n4228) );
  INV_X1 U3414 ( .A(n4228), .ZN(n3677) );
  NAND2_X1 U3415 ( .A1(n4736), .A2(n3677), .ZN(n3663) );
  NAND2_X1 U3416 ( .A1(n3722), .A2(n3663), .ZN(n3854) );
  INV_X1 U3417 ( .A(n3854), .ZN(n2634) );
  NAND2_X1 U3418 ( .A1(n3801), .A2(n3797), .ZN(n3721) );
  NAND2_X1 U3419 ( .A1(n3751), .A2(n3756), .ZN(n3666) );
  NAND2_X1 U3420 ( .A1(n3721), .A2(n3666), .ZN(n2633) );
  NOR2_X1 U3421 ( .A1(n4736), .A2(n3677), .ZN(n3664) );
  AOI21_X1 U3422 ( .B1(n2634), .B2(n2633), .A(n3664), .ZN(n3816) );
  NAND2_X1 U3423 ( .A1(n2636), .A2(n2635), .ZN(n2637) );
  NAND2_X1 U3424 ( .A1(n2641), .A2(n2637), .ZN(n3702) );
  OR2_X1 U3425 ( .A1(n3702), .A2(n2782), .ZN(n2640) );
  AOI22_X1 U3426 ( .A1(n2009), .A2(REG0_REG_14__SCAN_IN), .B1(n2912), .B2(
        REG1_REG_14__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U3427 ( .A1(n2913), .A2(REG2_REG_14__SCAN_IN), .ZN(n2638) );
  MUX2_X1 U3428 ( .A(DATAI_14_), .B(n4812), .S(n2011), .Z(n4723) );
  NAND2_X1 U3429 ( .A1(n4231), .A2(n4723), .ZN(n3815) );
  NAND2_X1 U3430 ( .A1(n4716), .A2(n3991), .ZN(n3817) );
  NAND2_X1 U3431 ( .A1(n3815), .A2(n3817), .ZN(n3911) );
  NAND2_X1 U3432 ( .A1(n2641), .A2(n3041), .ZN(n2642) );
  NAND2_X1 U3433 ( .A1(n2657), .A2(n2642), .ZN(n3776) );
  AOI22_X1 U3434 ( .A1(n2913), .A2(REG2_REG_15__SCAN_IN), .B1(n2009), .B2(
        REG0_REG_15__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U3435 ( .A1(n2912), .A2(REG1_REG_15__SCAN_IN), .ZN(n2643) );
  MUX2_X1 U3436 ( .A(DATAI_15_), .B(n2645), .S(n2011), .Z(n4715) );
  OR2_X1 U3437 ( .A1(n4303), .A2(n3779), .ZN(n3932) );
  NAND2_X1 U3438 ( .A1(n4303), .A2(n3779), .ZN(n3818) );
  NAND2_X1 U3439 ( .A1(n3932), .A2(n3818), .ZN(n3909) );
  INV_X1 U3440 ( .A(n3815), .ZN(n3930) );
  XNOR2_X1 U3441 ( .A(n2657), .B(REG3_REG_16__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U3442 ( .A1(n4640), .A2(n2581), .ZN(n2651) );
  NAND2_X1 U3443 ( .A1(n2912), .A2(REG1_REG_16__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3444 ( .A1(n2009), .A2(REG0_REG_16__SCAN_IN), .ZN(n2647) );
  OAI211_X1 U3445 ( .C1(n2785), .C2(n4841), .A(n2648), .B(n2647), .ZN(n2649)
         );
  INV_X1 U3446 ( .A(n2649), .ZN(n2650) );
  MUX2_X1 U3447 ( .A(DATAI_16_), .B(n2652), .S(n2909), .Z(n4629) );
  NAND2_X1 U3448 ( .A1(n4718), .A2(n4629), .ZN(n3933) );
  INV_X1 U3449 ( .A(n4629), .ZN(n4639) );
  NAND2_X1 U3450 ( .A1(n4611), .A2(n4639), .ZN(n3938) );
  AND2_X1 U3451 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2653) );
  INV_X1 U3452 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2656) );
  INV_X1 U3453 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2655) );
  OAI21_X1 U3454 ( .B1(n2657), .B2(n2656), .A(n2655), .ZN(n2658) );
  NAND2_X1 U3455 ( .A1(n2677), .A2(n2658), .ZN(n4202) );
  OR2_X1 U3456 ( .A1(n4202), .A2(n2782), .ZN(n2663) );
  INV_X1 U3457 ( .A(n2912), .ZN(n2766) );
  NAND2_X1 U34580 ( .A1(n2009), .A2(REG0_REG_17__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U34590 ( .A1(n2913), .A2(REG2_REG_17__SCAN_IN), .ZN(n2659) );
  OAI211_X1 U3460 ( .C1(n2766), .C2(n2507), .A(n2660), .B(n2659), .ZN(n2661)
         );
  INV_X1 U3461 ( .A(n2661), .ZN(n2662) );
  INV_X1 U3462 ( .A(DATAI_17_), .ZN(n2664) );
  MUX2_X1 U3463 ( .A(n2665), .B(n2664), .S(n2533), .Z(n4620) );
  AND2_X1 U3464 ( .A1(n4302), .A2(n4620), .ZN(n3895) );
  INV_X1 U3465 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3466 ( .A1(n2679), .A2(n2667), .ZN(n2668) );
  AND2_X1 U34670 ( .A1(n2691), .A2(n2668), .ZN(n4580) );
  NAND2_X1 U3468 ( .A1(n4580), .A2(n2581), .ZN(n2674) );
  INV_X1 U34690 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U3470 ( .A1(n2912), .A2(REG1_REG_19__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U34710 ( .A1(n2009), .A2(REG0_REG_19__SCAN_IN), .ZN(n2669) );
  OAI211_X1 U3472 ( .C1(n2785), .C2(n2671), .A(n2670), .B(n2669), .ZN(n2672)
         );
  INV_X1 U34730 ( .A(n2672), .ZN(n2673) );
  NAND2_X1 U3474 ( .A1(n2791), .A2(IR_REG_31__SCAN_IN), .ZN(n2675) );
  XNOR2_X2 U34750 ( .A(n2675), .B(IR_REG_19__SCAN_IN), .ZN(n3181) );
  MUX2_X1 U3476 ( .A(DATAI_19_), .B(n3181), .S(n2909), .Z(n4143) );
  NAND2_X1 U34770 ( .A1(n4593), .A2(n4579), .ZN(n2685) );
  INV_X1 U3478 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2676) );
  NAND2_X1 U34790 ( .A1(n2677), .A2(n2676), .ZN(n2678) );
  NAND2_X1 U3480 ( .A1(n2679), .A2(n2678), .ZN(n4261) );
  OR2_X1 U34810 ( .A1(n4261), .A2(n2782), .ZN(n2684) );
  NAND2_X1 U3482 ( .A1(n2009), .A2(REG0_REG_18__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U34830 ( .A1(n2913), .A2(REG2_REG_18__SCAN_IN), .ZN(n2680) );
  OAI211_X1 U3484 ( .C1(n2766), .C2(n4365), .A(n2681), .B(n2680), .ZN(n2682)
         );
  INV_X1 U34850 ( .A(n2682), .ZN(n2683) );
  INV_X1 U3486 ( .A(DATAI_18_), .ZN(n4874) );
  MUX2_X1 U34870 ( .A(n4874), .B(n4875), .S(n2011), .Z(n4598) );
  NAND2_X1 U3488 ( .A1(n4705), .A2(n4598), .ZN(n4569) );
  NAND2_X1 U34890 ( .A1(n2685), .A2(n4569), .ZN(n3936) );
  INV_X1 U3490 ( .A(n4598), .ZN(n4264) );
  NAND2_X1 U34910 ( .A1(n4572), .A2(n4264), .ZN(n4568) );
  NAND2_X1 U3492 ( .A1(n4627), .A2(n4704), .ZN(n4567) );
  AND2_X1 U34930 ( .A1(n4568), .A2(n4567), .ZN(n2687) );
  OR2_X1 U3494 ( .A1(n2687), .A2(n3936), .ZN(n2689) );
  INV_X1 U34950 ( .A(n4593), .ZN(n2844) );
  NAND2_X1 U3496 ( .A1(n2844), .A2(n4143), .ZN(n2688) );
  NAND2_X1 U34970 ( .A1(n2689), .A2(n2688), .ZN(n4544) );
  INV_X1 U3498 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U34990 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  NAND2_X1 U3500 ( .A1(n2711), .A2(n2692), .ZN(n4561) );
  INV_X1 U35010 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4776) );
  NAND2_X1 U3502 ( .A1(n2913), .A2(REG2_REG_20__SCAN_IN), .ZN(n2694) );
  NAND2_X1 U35030 ( .A1(n2912), .A2(REG1_REG_20__SCAN_IN), .ZN(n2693) );
  OAI211_X1 U3504 ( .C1(n2805), .C2(n4776), .A(n2694), .B(n2693), .ZN(n2695)
         );
  INV_X1 U35050 ( .A(n2695), .ZN(n2696) );
  INV_X1 U35060 ( .A(DATAI_20_), .ZN(n2698) );
  NOR2_X1 U35070 ( .A1(n2909), .A2(n2698), .ZN(n4549) );
  INV_X1 U35080 ( .A(n4549), .ZN(n4558) );
  NOR2_X1 U35090 ( .A1(n4683), .A2(n4558), .ZN(n2699) );
  NOR2_X1 U35100 ( .A1(n4544), .A2(n2699), .ZN(n3942) );
  NAND2_X1 U35110 ( .A1(n4546), .A2(n3942), .ZN(n2700) );
  NAND2_X1 U35120 ( .A1(n4683), .A2(n4558), .ZN(n3940) );
  INV_X1 U35130 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2710) );
  INV_X1 U35140 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4240) );
  NAND2_X1 U35150 ( .A1(n2713), .A2(n4240), .ZN(n2702) );
  NAND2_X1 U35160 ( .A1(n2721), .A2(n2702), .ZN(n4239) );
  INV_X1 U35170 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U35180 ( .A1(n2009), .A2(REG0_REG_22__SCAN_IN), .ZN(n2704) );
  NAND2_X1 U35190 ( .A1(n2912), .A2(REG1_REG_22__SCAN_IN), .ZN(n2703) );
  OAI211_X1 U35200 ( .C1(n2705), .C2(n2785), .A(n2704), .B(n2703), .ZN(n2706)
         );
  INV_X1 U35210 ( .A(n2706), .ZN(n2707) );
  INV_X1 U35220 ( .A(DATAI_22_), .ZN(n2709) );
  NOR2_X1 U35230 ( .A1(n2011), .A2(n2709), .ZN(n4518) );
  NAND2_X1 U35240 ( .A1(n4686), .A2(n4518), .ZN(n4489) );
  NAND2_X1 U35250 ( .A1(n2711), .A2(n2710), .ZN(n2712) );
  AND2_X1 U35260 ( .A1(n2713), .A2(n2712), .ZN(n4532) );
  NAND2_X1 U35270 ( .A1(n4532), .A2(n2581), .ZN(n2719) );
  INV_X1 U35280 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U35290 ( .A1(n2912), .A2(REG1_REG_21__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U35300 ( .A1(n2009), .A2(REG0_REG_21__SCAN_IN), .ZN(n2714) );
  OAI211_X1 U35310 ( .C1(n2785), .C2(n2716), .A(n2715), .B(n2714), .ZN(n2717)
         );
  INV_X1 U35320 ( .A(n2717), .ZN(n2718) );
  INV_X1 U35330 ( .A(DATAI_21_), .ZN(n2720) );
  NOR2_X1 U35340 ( .A1(n2011), .A2(n2720), .ZN(n4682) );
  NAND2_X1 U35350 ( .A1(n4551), .A2(n4682), .ZN(n4487) );
  AND2_X1 U35360 ( .A1(n4489), .A2(n4487), .ZN(n3944) );
  INV_X1 U35370 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4129) );
  NAND2_X1 U35380 ( .A1(n2721), .A2(n4129), .ZN(n2722) );
  NAND2_X1 U35390 ( .A1(n4501), .A2(n2014), .ZN(n2728) );
  INV_X1 U35400 ( .A(REG2_REG_23__SCAN_IN), .ZN(n2725) );
  NAND2_X1 U35410 ( .A1(n2912), .A2(REG1_REG_23__SCAN_IN), .ZN(n2724) );
  NAND2_X1 U35420 ( .A1(n2009), .A2(REG0_REG_23__SCAN_IN), .ZN(n2723) );
  OAI211_X1 U35430 ( .C1(n2785), .C2(n2725), .A(n2724), .B(n2723), .ZN(n2726)
         );
  INV_X1 U35440 ( .A(n2726), .ZN(n2727) );
  INV_X1 U35450 ( .A(DATAI_23_), .ZN(n2729) );
  NOR2_X1 U35460 ( .A1(n2011), .A2(n2729), .ZN(n4495) );
  INV_X1 U35470 ( .A(n4495), .ZN(n4499) );
  NAND2_X1 U35480 ( .A1(n4665), .A2(n4499), .ZN(n2730) );
  NAND2_X1 U35490 ( .A1(n4496), .A2(n2896), .ZN(n2849) );
  NAND2_X1 U35500 ( .A1(n2730), .A2(n2849), .ZN(n3866) );
  INV_X1 U35510 ( .A(n4682), .ZN(n4534) );
  AND2_X1 U35520 ( .A1(n4507), .A2(n4534), .ZN(n4486) );
  AND2_X1 U35530 ( .A1(n4489), .A2(n4486), .ZN(n2731) );
  NOR2_X1 U35540 ( .A1(n3866), .A2(n2731), .ZN(n3945) );
  INV_X1 U35550 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3031) );
  NAND2_X1 U35560 ( .A1(n2733), .A2(n3031), .ZN(n2734) );
  NAND2_X1 U35570 ( .A1(n2752), .A2(n2734), .ZN(n4476) );
  INV_X1 U35580 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U35590 ( .A1(n2913), .A2(REG2_REG_24__SCAN_IN), .ZN(n2736) );
  NAND2_X1 U35600 ( .A1(n2009), .A2(REG0_REG_24__SCAN_IN), .ZN(n2735) );
  OAI211_X1 U35610 ( .C1(n4671), .C2(n2766), .A(n2736), .B(n2735), .ZN(n2737)
         );
  INV_X1 U35620 ( .A(n2737), .ZN(n2738) );
  INV_X1 U35630 ( .A(DATAI_24_), .ZN(n2740) );
  NOR2_X1 U35640 ( .A1(n2011), .A2(n2740), .ZN(n4664) );
  INV_X1 U35650 ( .A(n4664), .ZN(n4474) );
  OR2_X1 U35660 ( .A1(n4656), .A2(n4474), .ZN(n3888) );
  OR2_X1 U35670 ( .A1(n4665), .A2(n4499), .ZN(n4464) );
  NAND2_X1 U35680 ( .A1(n4656), .A2(n4474), .ZN(n3887) );
  INV_X1 U35690 ( .A(n4451), .ZN(n2749) );
  XNOR2_X1 U35700 ( .A(n2752), .B(REG3_REG_25__SCAN_IN), .ZN(n4457) );
  NAND2_X1 U35710 ( .A1(n4457), .A2(n2581), .ZN(n2746) );
  INV_X1 U35720 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2743) );
  NAND2_X1 U35730 ( .A1(n2912), .A2(REG1_REG_25__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U35740 ( .A1(n2009), .A2(REG0_REG_25__SCAN_IN), .ZN(n2741) );
  OAI211_X1 U35750 ( .C1(n2785), .C2(n2743), .A(n2742), .B(n2741), .ZN(n2744)
         );
  INV_X1 U35760 ( .A(n2744), .ZN(n2745) );
  INV_X1 U35770 ( .A(DATAI_25_), .ZN(n2747) );
  NOR2_X1 U35780 ( .A1(n2011), .A2(n2747), .ZN(n4655) );
  INV_X1 U35790 ( .A(n4655), .ZN(n4456) );
  NAND2_X1 U35800 ( .A1(n2749), .A2(n2748), .ZN(n4434) );
  INV_X1 U35810 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2750) );
  OAI21_X1 U3582 ( .B1(n2752), .B2(n3003), .A(n2750), .ZN(n2753) );
  NAND2_X1 U3583 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2751) );
  NAND2_X1 U3584 ( .A1(n2753), .A2(n2762), .ZN(n4446) );
  INV_X1 U3585 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4445) );
  NAND2_X1 U3586 ( .A1(n2912), .A2(REG1_REG_26__SCAN_IN), .ZN(n2755) );
  NAND2_X1 U3587 ( .A1(n2009), .A2(REG0_REG_26__SCAN_IN), .ZN(n2754) );
  OAI211_X1 U3588 ( .C1(n2785), .C2(n4445), .A(n2755), .B(n2754), .ZN(n2756)
         );
  INV_X1 U3589 ( .A(n2756), .ZN(n2757) );
  INV_X1 U3590 ( .A(DATAI_26_), .ZN(n2759) );
  NOR2_X1 U3591 ( .A1(n2909), .A2(n2759), .ZN(n4442) );
  NAND2_X1 U3592 ( .A1(n4659), .A2(n4442), .ZN(n2760) );
  OR2_X1 U3593 ( .A1(n4473), .A2(n4456), .ZN(n4433) );
  INV_X1 U3594 ( .A(n4442), .ZN(n4437) );
  NAND2_X1 U3595 ( .A1(n4424), .A2(n4437), .ZN(n3954) );
  INV_X1 U3596 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U3597 ( .A1(n2762), .A2(n2761), .ZN(n2763) );
  NAND2_X1 U3598 ( .A1(n2773), .A2(n2763), .ZN(n4421) );
  INV_X1 U3599 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3062) );
  NAND2_X1 U3600 ( .A1(n2913), .A2(REG2_REG_27__SCAN_IN), .ZN(n2765) );
  NAND2_X1 U3601 ( .A1(n2009), .A2(REG0_REG_27__SCAN_IN), .ZN(n2764) );
  OAI211_X1 U3602 ( .C1(n2766), .C2(n3062), .A(n2765), .B(n2764), .ZN(n2767)
         );
  INV_X1 U3603 ( .A(n2767), .ZN(n2768) );
  NAND2_X1 U3604 ( .A1(n2533), .A2(DATAI_27_), .ZN(n4419) );
  NAND2_X1 U3605 ( .A1(n4438), .A2(n4109), .ZN(n3950) );
  NAND2_X1 U3606 ( .A1(n4301), .A2(n4419), .ZN(n3874) );
  NAND2_X1 U3607 ( .A1(n3950), .A2(n3874), .ZN(n3956) );
  INV_X1 U3608 ( .A(n3956), .ZN(n2770) );
  NAND2_X1 U3609 ( .A1(n2771), .A2(n3950), .ZN(n3078) );
  INV_X1 U3610 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U3611 ( .A1(n2773), .A2(n2772), .ZN(n2774) );
  NAND2_X1 U3612 ( .A1(n4397), .A2(n2774), .ZN(n4408) );
  INV_X1 U3613 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4407) );
  NAND2_X1 U3614 ( .A1(n2912), .A2(REG1_REG_28__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U3615 ( .A1(n2009), .A2(REG0_REG_28__SCAN_IN), .ZN(n2775) );
  OAI211_X1 U3616 ( .C1(n2785), .C2(n4407), .A(n2776), .B(n2775), .ZN(n2777)
         );
  INV_X1 U3617 ( .A(n2777), .ZN(n2778) );
  INV_X1 U3618 ( .A(DATAI_28_), .ZN(n2780) );
  NOR2_X1 U3619 ( .A1(n2011), .A2(n2780), .ZN(n4095) );
  INV_X1 U3620 ( .A(n4095), .ZN(n4406) );
  NAND2_X1 U3621 ( .A1(n4396), .A2(n4406), .ZN(n3873) );
  NAND2_X1 U3622 ( .A1(n3078), .A2(n3873), .ZN(n2781) );
  NAND2_X1 U3623 ( .A1(n4426), .A2(n4095), .ZN(n3953) );
  NAND2_X1 U3624 ( .A1(n2781), .A2(n3953), .ZN(n2790) );
  OR2_X1 U3625 ( .A1(n4397), .A2(n2782), .ZN(n2788) );
  INV_X1 U3626 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U3627 ( .A1(n2912), .A2(REG1_REG_29__SCAN_IN), .ZN(n2784) );
  NAND2_X1 U3628 ( .A1(n2009), .A2(REG0_REG_29__SCAN_IN), .ZN(n2783) );
  OAI211_X1 U3629 ( .C1(n2785), .C2(n4393), .A(n2784), .B(n2783), .ZN(n2786)
         );
  INV_X1 U3630 ( .A(n2786), .ZN(n2787) );
  NAND2_X1 U3631 ( .A1(n2788), .A2(n2787), .ZN(n4300) );
  INV_X1 U3632 ( .A(DATAI_29_), .ZN(n2789) );
  NOR2_X1 U3633 ( .A1(n2909), .A2(n2789), .ZN(n3879) );
  XNOR2_X1 U3634 ( .A(n4300), .B(n3879), .ZN(n3929) );
  XNOR2_X1 U3635 ( .A(n2790), .B(n3929), .ZN(n2801) );
  NAND2_X1 U3636 ( .A1(n3181), .A2(n2807), .ZN(n2800) );
  INV_X1 U3637 ( .A(n2791), .ZN(n2798) );
  INV_X1 U3638 ( .A(IR_REG_20__SCAN_IN), .ZN(n2795) );
  NAND2_X1 U3639 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2793) );
  NAND2_X1 U3640 ( .A1(n2793), .A2(IR_REG_31__SCAN_IN), .ZN(n2794) );
  OAI21_X1 U3641 ( .B1(n2795), .B2(IR_REG_31__SCAN_IN), .A(n2794), .ZN(n2796)
         );
  NAND2_X1 U3642 ( .A1(n4811), .A2(n2862), .ZN(n2799) );
  NAND2_X1 U3643 ( .A1(n3185), .A2(n4822), .ZN(n4726) );
  INV_X1 U3644 ( .A(B_REG_SCAN_IN), .ZN(n2873) );
  NOR2_X1 U3645 ( .A1(n4824), .A2(n2873), .ZN(n2802) );
  NOR2_X1 U3646 ( .A1(n4726), .A2(n2802), .ZN(n2918) );
  INV_X1 U3647 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2994) );
  NAND2_X1 U3648 ( .A1(n2913), .A2(REG2_REG_30__SCAN_IN), .ZN(n2804) );
  NAND2_X1 U3649 ( .A1(n2912), .A2(REG1_REG_30__SCAN_IN), .ZN(n2803) );
  OAI211_X1 U3650 ( .C1(n2805), .C2(n2994), .A(n2804), .B(n2803), .ZN(n4299)
         );
  NAND2_X1 U3651 ( .A1(n2918), .A2(n4299), .ZN(n2806) );
  INV_X1 U3652 ( .A(n3879), .ZN(n4394) );
  INV_X1 U3653 ( .A(n2807), .ZN(n3182) );
  INV_X1 U3654 ( .A(n2862), .ZN(n2808) );
  NAND2_X1 U3655 ( .A1(n4396), .A2(n4738), .ZN(n2809) );
  OAI21_X1 U3656 ( .B1(n4394), .B2(n4741), .A(n2809), .ZN(n2810) );
  AND2_X1 U3657 ( .A1(n3456), .A2(n4149), .ZN(n3162) );
  NAND2_X1 U3658 ( .A1(n3340), .A2(n4311), .ZN(n2812) );
  NAND2_X1 U3659 ( .A1(n3261), .A2(n4253), .ZN(n3335) );
  AND2_X1 U3660 ( .A1(n2812), .A2(n3335), .ZN(n2811) );
  NAND3_X1 U3661 ( .A1(n3160), .A2(n2811), .A3(n3354), .ZN(n2814) );
  NOR2_X1 U3662 ( .A1(n2013), .A2(n4313), .ZN(n3336) );
  AOI22_X1 U3663 ( .A1(n3336), .A2(n2812), .B1(n3361), .B2(n3349), .ZN(n2813)
         );
  NAND2_X1 U3664 ( .A1(n2814), .A2(n2813), .ZN(n3468) );
  INV_X1 U3665 ( .A(n3468), .ZN(n2815) );
  NAND2_X1 U3666 ( .A1(n3397), .A2(n4309), .ZN(n3306) );
  NAND2_X1 U3667 ( .A1(n3470), .A2(n4310), .ZN(n3304) );
  NOR2_X1 U3668 ( .A1(n2817), .A2(n2816), .ZN(n2818) );
  NAND2_X1 U3669 ( .A1(n3302), .A2(n2818), .ZN(n2823) );
  NAND2_X2 U3670 ( .A1(n2819), .A2(n3839), .ZN(n3890) );
  INV_X1 U3671 ( .A(n3890), .ZN(n3584) );
  NAND2_X1 U3672 ( .A1(n3596), .A2(n3554), .ZN(n3305) );
  NAND2_X1 U3673 ( .A1(n3579), .A2(n3595), .ZN(n2820) );
  NAND2_X1 U3674 ( .A1(n3305), .A2(n2820), .ZN(n2821) );
  NOR2_X1 U3675 ( .A1(n3584), .A2(n2821), .ZN(n2822) );
  NAND2_X1 U3676 ( .A1(n2823), .A2(n2822), .ZN(n2826) );
  AND2_X1 U3677 ( .A1(n3443), .A2(n4308), .ZN(n2824) );
  AOI22_X1 U3678 ( .A1(n3890), .A2(n2824), .B1(n3570), .B2(n3599), .ZN(n2825)
         );
  NAND2_X1 U3679 ( .A1(n3539), .A2(n3623), .ZN(n2827) );
  NAND2_X1 U3680 ( .A1(n3536), .A2(n4307), .ZN(n2828) );
  AND2_X1 U3681 ( .A1(n3656), .A2(n4306), .ZN(n2830) );
  NAND2_X1 U3682 ( .A1(n3666), .A2(n3851), .ZN(n3636) );
  NAND2_X1 U3683 ( .A1(n3751), .A2(n3640), .ZN(n2831) );
  NAND2_X1 U3684 ( .A1(n3635), .A2(n2831), .ZN(n3725) );
  NAND2_X1 U3685 ( .A1(n3801), .A2(n4304), .ZN(n2832) );
  NAND2_X1 U3686 ( .A1(n3725), .A2(n2832), .ZN(n2834) );
  NAND2_X1 U3687 ( .A1(n2893), .A2(n3797), .ZN(n2833) );
  NAND2_X1 U3688 ( .A1(n2834), .A2(n2833), .ZN(n3673) );
  NOR2_X1 U3689 ( .A1(n4736), .A2(n4228), .ZN(n2835) );
  NAND2_X1 U3690 ( .A1(n4303), .A2(n4715), .ZN(n2836) );
  OR2_X1 U3691 ( .A1(n4303), .A2(n4715), .ZN(n2837) );
  NAND2_X1 U3692 ( .A1(n4611), .A2(n4629), .ZN(n2838) );
  NAND2_X1 U3693 ( .A1(n4627), .A2(n4620), .ZN(n2839) );
  NAND2_X1 U3694 ( .A1(n4302), .A2(n4704), .ZN(n2840) );
  NAND2_X1 U3695 ( .A1(n4572), .A2(n4598), .ZN(n2842) );
  NAND2_X1 U3696 ( .A1(n4593), .A2(n4143), .ZN(n2843) );
  NAND2_X1 U3697 ( .A1(n4543), .A2(n3905), .ZN(n2845) );
  INV_X1 U3698 ( .A(n4683), .ZN(n4536) );
  NAND2_X1 U3699 ( .A1(n4536), .A2(n4558), .ZN(n3906) );
  NAND2_X1 U3700 ( .A1(n2845), .A2(n3906), .ZN(n4528) );
  NAND2_X1 U3701 ( .A1(n4507), .A2(n4682), .ZN(n2846) );
  NAND2_X1 U3702 ( .A1(n4551), .A2(n4534), .ZN(n2847) );
  NAND2_X1 U3703 ( .A1(n4496), .A2(n4518), .ZN(n2850) );
  OR2_X1 U3704 ( .A1(n4665), .A2(n4495), .ZN(n2851) );
  NAND2_X1 U3705 ( .A1(n4484), .A2(n2851), .ZN(n2853) );
  NAND2_X1 U3706 ( .A1(n4665), .A2(n4495), .ZN(n2852) );
  AND2_X1 U3707 ( .A1(n4656), .A2(n4664), .ZN(n2854) );
  NOR2_X1 U3708 ( .A1(n4473), .A2(n4655), .ZN(n2856) );
  NAND2_X1 U3709 ( .A1(n4473), .A2(n4655), .ZN(n2855) );
  NAND2_X1 U3710 ( .A1(n4659), .A2(n4437), .ZN(n3886) );
  INV_X1 U3711 ( .A(n3886), .ZN(n2858) );
  AND2_X1 U3712 ( .A1(n4438), .A2(n4419), .ZN(n2857) );
  NOR2_X1 U3713 ( .A1(n2858), .A2(n2857), .ZN(n2859) );
  NAND2_X1 U3714 ( .A1(n3055), .A2(n2859), .ZN(n2861) );
  NAND2_X1 U3715 ( .A1(n4301), .A2(n4109), .ZN(n2860) );
  NAND2_X1 U3716 ( .A1(n3953), .A2(n3873), .ZN(n3077) );
  NAND2_X1 U3717 ( .A1(n4396), .A2(n4095), .ZN(n4389) );
  NAND2_X1 U3718 ( .A1(n3929), .A2(n4389), .ZN(n2867) );
  INV_X1 U3719 ( .A(n4389), .ZN(n2864) );
  INV_X1 U3720 ( .A(n3929), .ZN(n4391) );
  XNOR2_X1 U3721 ( .A(n3256), .B(n2807), .ZN(n2863) );
  INV_X1 U3722 ( .A(n3181), .ZN(n4373) );
  NAND2_X1 U3723 ( .A1(n2863), .A2(n4373), .ZN(n4555) );
  NAND2_X1 U3724 ( .A1(n3181), .A2(n2900), .ZN(n3455) );
  AOI21_X1 U3725 ( .B1(n2864), .B2(n4391), .A(n4678), .ZN(n2865) );
  OAI21_X1 U3726 ( .B1(n3077), .B2(n2867), .A(n2865), .ZN(n2866) );
  INV_X1 U3727 ( .A(n2866), .ZN(n2869) );
  NAND2_X1 U3728 ( .A1(n2870), .A2(IR_REG_31__SCAN_IN), .ZN(n2872) );
  INV_X1 U3729 ( .A(n3113), .ZN(n3109) );
  NAND2_X1 U3730 ( .A1(n3109), .A2(n2873), .ZN(n2876) );
  INV_X1 U3731 ( .A(n3105), .ZN(n2874) );
  NAND3_X1 U3732 ( .A1(n3113), .A2(B_REG_SCAN_IN), .A3(n2874), .ZN(n2875) );
  NAND3_X1 U3733 ( .A1(n2876), .A2(n2875), .A3(n3101), .ZN(n3111) );
  OR2_X1 U3734 ( .A1(n3111), .A2(D_REG_1__SCAN_IN), .ZN(n3179) );
  OR2_X1 U3735 ( .A1(n3105), .A2(n3101), .ZN(n3177) );
  NAND2_X1 U3736 ( .A1(n3179), .A2(n3177), .ZN(n2889) );
  INV_X1 U3737 ( .A(n3449), .ZN(n3191) );
  OR2_X1 U3738 ( .A1(n4811), .A2(n3181), .ZN(n3184) );
  NAND2_X1 U3739 ( .A1(n3184), .A2(n3185), .ZN(n3451) );
  OAI211_X1 U3740 ( .C1(n2862), .C2(n3363), .A(n3191), .B(n3451), .ZN(n2877)
         );
  INV_X1 U3741 ( .A(n2877), .ZN(n2888) );
  NOR4_X1 U3742 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2950) );
  NOR2_X1 U3743 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_31__SCAN_IN), .ZN(n2880)
         );
  NOR4_X1 U3744 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2879) );
  NOR4_X1 U3745 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2878) );
  NAND4_X1 U3746 ( .A1(n2950), .A2(n2880), .A3(n2879), .A4(n2878), .ZN(n2886)
         );
  NOR4_X1 U3747 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2884) );
  NOR4_X1 U3748 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2883) );
  NOR4_X1 U3749 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2882) );
  NOR4_X1 U3750 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2881) );
  NAND4_X1 U3751 ( .A1(n2884), .A2(n2883), .A3(n2882), .A4(n2881), .ZN(n2885)
         );
  NOR2_X1 U3752 ( .A1(n2886), .A2(n2885), .ZN(n2887) );
  OR2_X1 U3753 ( .A1(n3111), .A2(n2887), .ZN(n3178) );
  OR2_X1 U3754 ( .A1(n3111), .A2(D_REG_0__SCAN_IN), .ZN(n2891) );
  INV_X1 U3755 ( .A(n3101), .ZN(n3112) );
  NAND2_X1 U3756 ( .A1(n3113), .A2(n3112), .ZN(n2890) );
  NAND2_X1 U3757 ( .A1(n3071), .A2(n4915), .ZN(n2907) );
  NAND2_X1 U3758 ( .A1(n3164), .A2(n3458), .ZN(n3173) );
  NAND2_X1 U3759 ( .A1(n3348), .A2(n3349), .ZN(n3347) );
  INV_X1 U3760 ( .A(n2897), .ZN(n3084) );
  NAND2_X1 U3761 ( .A1(n3084), .A2(n3879), .ZN(n2898) );
  NAND2_X1 U3762 ( .A1(n2910), .A2(n2898), .ZN(n4398) );
  NAND2_X1 U3763 ( .A1(n2902), .A2(n2901), .ZN(n2905) );
  INV_X1 U3764 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2903) );
  OR2_X1 U3765 ( .A1(n4915), .A2(n2903), .ZN(n2904) );
  NAND2_X1 U3766 ( .A1(n2907), .A2(n2906), .ZN(U3547) );
  INV_X1 U3767 ( .A(DATAI_30_), .ZN(n2908) );
  NOR2_X1 U3768 ( .A1(n2909), .A2(n2908), .ZN(n4386) );
  NAND2_X1 U3769 ( .A1(n2533), .A2(DATAI_31_), .ZN(n4382) );
  XNOR2_X1 U3770 ( .A(n4385), .B(n2911), .ZN(n4378) );
  NAND2_X1 U3771 ( .A1(n4378), .A2(n4597), .ZN(n2921) );
  NAND2_X1 U3772 ( .A1(n2912), .A2(REG1_REG_31__SCAN_IN), .ZN(n2917) );
  NAND2_X1 U3773 ( .A1(n2913), .A2(REG2_REG_31__SCAN_IN), .ZN(n2916) );
  NAND2_X1 U3774 ( .A1(n2009), .A2(REG0_REG_31__SCAN_IN), .ZN(n2915) );
  NAND3_X1 U3775 ( .A1(n2917), .A2(n2916), .A3(n2915), .ZN(n4298) );
  NAND2_X1 U3776 ( .A1(n2918), .A2(n4298), .ZN(n4383) );
  NAND2_X1 U3777 ( .A1(n2921), .A2(n2920), .ZN(n4648) );
  NAND2_X1 U3778 ( .A1(n4648), .A2(n4907), .ZN(n2924) );
  OR2_X1 U3779 ( .A1(n4907), .A2(n3017), .ZN(n2923) );
  NAND2_X1 U3780 ( .A1(n2924), .A2(n2923), .ZN(n3054) );
  NAND4_X1 U3781 ( .A1(n3003), .A2(n2925), .A3(REG2_REG_20__SCAN_IN), .A4(
        REG1_REG_16__SCAN_IN), .ZN(n2933) );
  INV_X1 U3782 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2926) );
  NAND4_X1 U3783 ( .A1(n2926), .A2(n3103), .A3(REG2_REG_0__SCAN_IN), .A4(
        DATAI_7_), .ZN(n2932) );
  NOR3_X1 U3784 ( .A1(IR_REG_6__SCAN_IN), .A2(REG1_REG_3__SCAN_IN), .A3(
        REG0_REG_31__SCAN_IN), .ZN(n2928) );
  AND4_X1 U3785 ( .A1(REG2_REG_25__SCAN_IN), .A2(REG2_REG_17__SCAN_IN), .A3(
        REG1_REG_24__SCAN_IN), .A4(n3031), .ZN(n2927) );
  NAND4_X1 U3786 ( .A1(n2929), .A2(D_REG_30__SCAN_IN), .A3(n2928), .A4(n2927), 
        .ZN(n2931) );
  NAND4_X1 U3787 ( .A1(REG2_REG_9__SCAN_IN), .A2(ADDR_REG_12__SCAN_IN), .A3(
        DATAO_REG_11__SCAN_IN), .A4(DATAO_REG_14__SCAN_IN), .ZN(n2930) );
  NOR4_X1 U3788 ( .A1(n2933), .A2(n2932), .A3(n2931), .A4(n2930), .ZN(n2937)
         );
  INV_X1 U3789 ( .A(DATAI_5_), .ZN(n3038) );
  NAND4_X1 U3790 ( .A1(IR_REG_30__SCAN_IN), .A2(REG1_REG_5__SCAN_IN), .A3(
        DATAO_REG_7__SCAN_IN), .A4(n3038), .ZN(n2935) );
  NAND4_X1 U3791 ( .A1(REG3_REG_15__SCAN_IN), .A2(D_REG_1__SCAN_IN), .A3(
        DATAI_23_), .A4(n3062), .ZN(n2934) );
  NOR2_X1 U3792 ( .A1(n2935), .A2(n2934), .ZN(n2936) );
  INV_X1 U3793 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n3157) );
  NAND4_X1 U3794 ( .A1(n2937), .A2(n2936), .A3(n3157), .A4(
        DATAO_REG_12__SCAN_IN), .ZN(n2948) );
  INV_X1 U3795 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4797) );
  NOR4_X1 U3796 ( .A1(REG3_REG_22__SCAN_IN), .A2(REG1_REG_11__SCAN_IN), .A3(
        n4797), .A4(n4913), .ZN(n2942) );
  NOR3_X1 U3797 ( .A1(IR_REG_19__SCAN_IN), .A2(DATAI_18_), .A3(
        DATAO_REG_19__SCAN_IN), .ZN(n2941) );
  NAND3_X1 U3798 ( .A1(DATAI_11_), .A2(REG2_REG_7__SCAN_IN), .A3(
        ADDR_REG_8__SCAN_IN), .ZN(n2939) );
  INV_X1 U3799 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4898) );
  NAND3_X1 U3800 ( .A1(REG0_REG_2__SCAN_IN), .A2(REG0_REG_30__SCAN_IN), .A3(
        n4898), .ZN(n2938) );
  NOR4_X1 U3801 ( .A1(DATAI_15_), .A2(DATAO_REG_0__SCAN_IN), .A3(n2939), .A4(
        n2938), .ZN(n2940) );
  NAND4_X1 U3802 ( .A1(REG3_REG_8__SCAN_IN), .A2(n2942), .A3(n2941), .A4(n2940), .ZN(n2947) );
  NOR4_X1 U3803 ( .A1(REG0_REG_0__SCAN_IN), .A2(REG1_REG_10__SCAN_IN), .A3(
        ADDR_REG_15__SCAN_IN), .A4(n4776), .ZN(n2945) );
  INV_X1 U3804 ( .A(DATAI_14_), .ZN(n2998) );
  NOR4_X1 U3805 ( .A1(IR_REG_27__SCAN_IN), .A2(DATAO_REG_1__SCAN_IN), .A3(
        n2954), .A4(n2998), .ZN(n2944) );
  NOR3_X1 U3806 ( .A1(IR_REG_24__SCAN_IN), .A2(DATAI_0_), .A3(
        DATAO_REG_22__SCAN_IN), .ZN(n2943) );
  NAND4_X1 U3807 ( .A1(DATAI_19_), .A2(n2945), .A3(n2944), .A4(n2943), .ZN(
        n2946) );
  NOR3_X1 U3808 ( .A1(n2948), .A2(n2947), .A3(n2946), .ZN(n2949) );
  AOI21_X1 U3809 ( .B1(n2950), .B2(n2949), .A(IR_REG_10__SCAN_IN), .ZN(n3052)
         );
  INV_X1 U3810 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n3149) );
  INV_X1 U3811 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n2952) );
  AOI22_X1 U3812 ( .A1(n3149), .A2(keyinput16), .B1(keyinput21), .B2(n2952), 
        .ZN(n2951) );
  OAI221_X1 U3813 ( .B1(n3149), .B2(keyinput16), .C1(n2952), .C2(keyinput21), 
        .A(n2951), .ZN(n2967) );
  INV_X1 U3814 ( .A(D_REG_30__SCAN_IN), .ZN(n4866) );
  AOI22_X1 U3815 ( .A1(n3157), .A2(keyinput40), .B1(n4866), .B2(keyinput37), 
        .ZN(n2953) );
  OAI221_X1 U3816 ( .B1(n3157), .B2(keyinput40), .C1(n4866), .C2(keyinput37), 
        .A(n2953), .ZN(n2966) );
  XOR2_X1 U3817 ( .A(n2954), .B(keyinput35), .Z(n2959) );
  XOR2_X1 U3818 ( .A(n2540), .B(keyinput27), .Z(n2958) );
  XOR2_X1 U3819 ( .A(n2955), .B(keyinput17), .Z(n2957) );
  XNOR2_X1 U3820 ( .A(IR_REG_3__SCAN_IN), .B(keyinput47), .ZN(n2956) );
  NAND4_X1 U3821 ( .A1(n2959), .A2(n2958), .A3(n2957), .A4(n2956), .ZN(n2965)
         );
  XNOR2_X1 U3822 ( .A(IR_REG_6__SCAN_IN), .B(keyinput38), .ZN(n2963) );
  XNOR2_X1 U3823 ( .A(IR_REG_19__SCAN_IN), .B(keyinput42), .ZN(n2962) );
  XNOR2_X1 U3824 ( .A(IR_REG_27__SCAN_IN), .B(keyinput20), .ZN(n2961) );
  XNOR2_X1 U3825 ( .A(IR_REG_22__SCAN_IN), .B(keyinput33), .ZN(n2960) );
  NAND4_X1 U3826 ( .A1(n2963), .A2(n2962), .A3(n2961), .A4(n2960), .ZN(n2964)
         );
  NOR4_X1 U3827 ( .A1(n2967), .A2(n2966), .A3(n2965), .A4(n2964), .ZN(n2980)
         );
  INV_X1 U3828 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n2968) );
  XOR2_X1 U3829 ( .A(keyinput54), .B(n2968), .Z(n2979) );
  XNOR2_X1 U3830 ( .A(keyinput41), .B(n2926), .ZN(n2970) );
  XOR2_X1 U3831 ( .A(REG1_REG_16__SCAN_IN), .B(keyinput14), .Z(n2969) );
  AOI211_X1 U3832 ( .C1(keyinput56), .C2(n2971), .A(n2970), .B(n2969), .ZN(
        n2978) );
  XOR2_X1 U3833 ( .A(REG2_REG_0__SCAN_IN), .B(keyinput13), .Z(n2976) );
  XNOR2_X1 U3834 ( .A(n2972), .B(keyinput61), .ZN(n2975) );
  XNOR2_X1 U3835 ( .A(n4874), .B(keyinput46), .ZN(n2974) );
  XNOR2_X1 U3836 ( .A(n3103), .B(keyinput12), .ZN(n2973) );
  NOR4_X1 U3837 ( .A1(n2976), .A2(n2975), .A3(n2974), .A4(n2973), .ZN(n2977)
         );
  AND4_X1 U3838 ( .A1(n2980), .A2(n2979), .A3(n2978), .A4(n2977), .ZN(n2985)
         );
  OAI22_X1 U3839 ( .A1(n4240), .A2(keyinput58), .B1(n4913), .B2(keyinput49), 
        .ZN(n2981) );
  AOI221_X1 U3840 ( .B1(n4240), .B2(keyinput58), .C1(keyinput49), .C2(n4913), 
        .A(n2981), .ZN(n2984) );
  INV_X1 U3841 ( .A(D_REG_12__SCAN_IN), .ZN(n4868) );
  INV_X1 U3842 ( .A(D_REG_10__SCAN_IN), .ZN(n4869) );
  OAI22_X1 U3843 ( .A1(n4868), .A2(keyinput62), .B1(n4869), .B2(keyinput52), 
        .ZN(n2982) );
  AOI221_X1 U3844 ( .B1(n4868), .B2(keyinput62), .C1(keyinput52), .C2(n4869), 
        .A(n2982), .ZN(n2983) );
  NAND3_X1 U3845 ( .A1(n2985), .A2(n2984), .A3(n2983), .ZN(n3014) );
  INV_X1 U3846 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4892) );
  OAI22_X1 U3847 ( .A1(n4898), .A2(keyinput45), .B1(n4892), .B2(keyinput48), 
        .ZN(n2986) );
  AOI221_X1 U3848 ( .B1(n4898), .B2(keyinput45), .C1(keyinput48), .C2(n4892), 
        .A(n2986), .ZN(n2989) );
  INV_X1 U3849 ( .A(DATAI_15_), .ZN(n4878) );
  INV_X1 U3850 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n3159) );
  OAI22_X1 U3851 ( .A1(n4878), .A2(keyinput50), .B1(n3159), .B2(keyinput44), 
        .ZN(n2987) );
  AOI221_X1 U3852 ( .B1(n4878), .B2(keyinput50), .C1(keyinput44), .C2(n3159), 
        .A(n2987), .ZN(n2988) );
  NAND2_X1 U3853 ( .A1(n2989), .A2(n2988), .ZN(n3013) );
  INV_X1 U3854 ( .A(DATAI_11_), .ZN(n2992) );
  OAI22_X1 U3855 ( .A1(n2992), .A2(keyinput18), .B1(n2991), .B2(keyinput57), 
        .ZN(n2990) );
  AOI221_X1 U3856 ( .B1(n2992), .B2(keyinput18), .C1(keyinput57), .C2(n2991), 
        .A(n2990), .ZN(n3011) );
  OAI22_X1 U3857 ( .A1(n4797), .A2(keyinput60), .B1(n2994), .B2(keyinput53), 
        .ZN(n2993) );
  AOI221_X1 U3858 ( .B1(n4797), .B2(keyinput60), .C1(keyinput53), .C2(n2994), 
        .A(n2993), .ZN(n3010) );
  INV_X1 U3859 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U3860 ( .A1(n3062), .A2(keyinput8), .B1(keyinput10), .B2(n3155), 
        .ZN(n2995) );
  OAI221_X1 U3861 ( .B1(n3062), .B2(keyinput8), .C1(n3155), .C2(keyinput10), 
        .A(n2995), .ZN(n3000) );
  INV_X1 U3862 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n2997) );
  AOI22_X1 U3863 ( .A1(n2998), .A2(keyinput55), .B1(keyinput59), .B2(n2997), 
        .ZN(n2996) );
  OAI221_X1 U3864 ( .B1(n2998), .B2(keyinput55), .C1(n2997), .C2(keyinput59), 
        .A(n2996), .ZN(n2999) );
  NOR2_X1 U3865 ( .A1(n3000), .A2(n2999), .ZN(n3009) );
  INV_X1 U3866 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3003) );
  INV_X1 U3867 ( .A(DATAI_7_), .ZN(n3002) );
  AOI22_X1 U3868 ( .A1(n3003), .A2(keyinput32), .B1(keyinput34), .B2(n3002), 
        .ZN(n3001) );
  OAI221_X1 U3869 ( .B1(n3003), .B2(keyinput32), .C1(n3002), .C2(keyinput34), 
        .A(n3001), .ZN(n3007) );
  INV_X1 U3870 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U3871 ( .A1(n3005), .A2(keyinput51), .B1(keyinput39), .B2(n3151), 
        .ZN(n3004) );
  OAI221_X1 U3872 ( .B1(n3005), .B2(keyinput51), .C1(n3151), .C2(keyinput39), 
        .A(n3004), .ZN(n3006) );
  NOR2_X1 U3873 ( .A1(n3007), .A2(n3006), .ZN(n3008) );
  NAND4_X1 U3874 ( .A1(n3011), .A2(n3010), .A3(n3009), .A4(n3008), .ZN(n3012)
         );
  NOR3_X1 U3875 ( .A1(n3014), .A2(n3013), .A3(n3012), .ZN(n3050) );
  INV_X1 U3876 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3017) );
  AOI22_X1 U3877 ( .A1(n3017), .A2(keyinput36), .B1(n3016), .B2(keyinput22), 
        .ZN(n3015) );
  OAI221_X1 U3878 ( .B1(n3017), .B2(keyinput36), .C1(n3016), .C2(keyinput22), 
        .A(n3015), .ZN(n3026) );
  INV_X1 U3879 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3020) );
  INV_X1 U3880 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n3019) );
  AOI22_X1 U3881 ( .A1(n3020), .A2(keyinput24), .B1(keyinput28), .B2(n3019), 
        .ZN(n3018) );
  OAI221_X1 U3882 ( .B1(n3020), .B2(keyinput24), .C1(n3019), .C2(keyinput28), 
        .A(n3018), .ZN(n3025) );
  INV_X1 U3883 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4885) );
  AOI22_X1 U3884 ( .A1(n2100), .A2(keyinput30), .B1(keyinput29), .B2(n4885), 
        .ZN(n3021) );
  OAI221_X1 U3885 ( .B1(n2100), .B2(keyinput30), .C1(n4885), .C2(keyinput29), 
        .A(n3021), .ZN(n3024) );
  INV_X1 U3886 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U3887 ( .A1(n4776), .A2(keyinput25), .B1(keyinput26), .B2(n3153), 
        .ZN(n3022) );
  OAI221_X1 U3888 ( .B1(n4776), .B2(keyinput25), .C1(n3153), .C2(keyinput26), 
        .A(n3022), .ZN(n3023) );
  NOR4_X1 U3889 ( .A1(n3026), .A2(n3025), .A3(n3024), .A4(n3023), .ZN(n3049)
         );
  INV_X1 U3890 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U3891 ( .A1(n2871), .A2(keyinput19), .B1(keyinput23), .B2(n3213), 
        .ZN(n3027) );
  OAI221_X1 U3892 ( .B1(n2871), .B2(keyinput19), .C1(n3213), .C2(keyinput23), 
        .A(n3027), .ZN(n3036) );
  INV_X1 U3893 ( .A(DATAI_19_), .ZN(n3029) );
  AOI22_X1 U3894 ( .A1(n3029), .A2(keyinput11), .B1(n2743), .B2(keyinput3), 
        .ZN(n3028) );
  OAI221_X1 U3895 ( .B1(n3029), .B2(keyinput11), .C1(n2743), .C2(keyinput3), 
        .A(n3028), .ZN(n3035) );
  AOI22_X1 U3896 ( .A1(n3031), .A2(keyinput7), .B1(keyinput31), .B2(n2441), 
        .ZN(n3030) );
  OAI221_X1 U3897 ( .B1(n3031), .B2(keyinput7), .C1(n2441), .C2(keyinput31), 
        .A(n3030), .ZN(n3034) );
  INV_X1 U3898 ( .A(D_REG_2__SCAN_IN), .ZN(n4871) );
  AOI22_X1 U3899 ( .A1(n4671), .A2(keyinput15), .B1(n4871), .B2(keyinput63), 
        .ZN(n3032) );
  OAI221_X1 U3900 ( .B1(n4671), .B2(keyinput15), .C1(n4871), .C2(keyinput63), 
        .A(n3032), .ZN(n3033) );
  NOR4_X1 U3901 ( .A1(n3036), .A2(n3035), .A3(n3034), .A4(n3033), .ZN(n3048)
         );
  INV_X1 U3902 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U3903 ( .A1(n3038), .A2(keyinput1), .B1(keyinput2), .B2(n3147), 
        .ZN(n3037) );
  OAI221_X1 U3904 ( .B1(n3038), .B2(keyinput1), .C1(n3147), .C2(keyinput2), 
        .A(n3037), .ZN(n3046) );
  INV_X1 U3905 ( .A(D_REG_25__SCAN_IN), .ZN(n4867) );
  AOI22_X1 U3906 ( .A1(n4867), .A2(keyinput43), .B1(keyinput0), .B2(n3373), 
        .ZN(n3039) );
  OAI221_X1 U3907 ( .B1(n4867), .B2(keyinput43), .C1(n3373), .C2(keyinput0), 
        .A(n3039), .ZN(n3045) );
  INV_X1 U3908 ( .A(D_REG_1__SCAN_IN), .ZN(n3117) );
  AOI22_X1 U3909 ( .A1(n3117), .A2(keyinput4), .B1(keyinput9), .B2(n3041), 
        .ZN(n3040) );
  OAI221_X1 U3910 ( .B1(n3117), .B2(keyinput4), .C1(n3041), .C2(keyinput9), 
        .A(n3040), .ZN(n3044) );
  AOI22_X1 U3911 ( .A1(n3093), .A2(keyinput5), .B1(keyinput6), .B2(n2729), 
        .ZN(n3042) );
  OAI221_X1 U3912 ( .B1(n3093), .B2(keyinput5), .C1(n2729), .C2(keyinput6), 
        .A(n3042), .ZN(n3043) );
  NOR4_X1 U3913 ( .A1(n3046), .A2(n3045), .A3(n3044), .A4(n3043), .ZN(n3047)
         );
  AND4_X1 U3914 ( .A1(n3050), .A2(n3049), .A3(n3048), .A4(n3047), .ZN(n3051)
         );
  OAI21_X1 U3915 ( .B1(n3052), .B2(keyinput56), .A(n3051), .ZN(n3053) );
  XNOR2_X1 U3916 ( .A(n3054), .B(n3053), .ZN(U3517) );
  XOR2_X1 U3917 ( .A(n3956), .B(n3056), .Z(n4417) );
  XNOR2_X1 U3918 ( .A(n3057), .B(n3956), .ZN(n3058) );
  NAND2_X1 U3919 ( .A1(n3058), .A2(n4590), .ZN(n4431) );
  AOI22_X1 U3920 ( .A1(n4424), .A2(n4738), .B1(n4109), .B2(n4724), .ZN(n3059)
         );
  OAI211_X1 U3921 ( .C1(n4426), .C2(n4726), .A(n4431), .B(n3059), .ZN(n3060)
         );
  AOI21_X1 U3922 ( .B1(n4417), .B2(n4900), .A(n3060), .ZN(n3066) );
  OR2_X1 U3923 ( .A1(n3066), .A2(n4912), .ZN(n3065) );
  AND2_X1 U3924 ( .A1(n4444), .A2(n4109), .ZN(n3061) );
  OR2_X1 U3925 ( .A1(n3061), .A2(n2022), .ZN(n4418) );
  OAI22_X1 U3926 ( .A1(n4418), .A2(n4746), .B1(n3062), .B2(n4915), .ZN(n3063)
         );
  INV_X1 U3927 ( .A(n3063), .ZN(n3064) );
  NAND2_X1 U3928 ( .A1(n3065), .A2(n3064), .ZN(U3545) );
  OR2_X1 U3929 ( .A1(n3066), .A2(n4905), .ZN(n3070) );
  INV_X1 U3930 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3067) );
  OAI22_X1 U3931 ( .A1(n4418), .A2(n4807), .B1(n3067), .B2(n4907), .ZN(n3068)
         );
  INV_X1 U3932 ( .A(n3068), .ZN(n3069) );
  NAND2_X1 U3933 ( .A1(n3070), .A2(n3069), .ZN(U3513) );
  NAND2_X1 U3934 ( .A1(n3071), .A2(n4907), .ZN(n3075) );
  INV_X1 U3935 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3072) );
  NAND2_X1 U3936 ( .A1(n3075), .A2(n3074), .ZN(U3515) );
  XNOR2_X1 U3937 ( .A(n3078), .B(n3076), .ZN(n3079) );
  NAND2_X1 U3938 ( .A1(n3079), .A2(n4590), .ZN(n4416) );
  AOI22_X1 U3939 ( .A1(n4301), .A2(n4738), .B1(n4095), .B2(n4724), .ZN(n3080)
         );
  INV_X1 U3940 ( .A(n4300), .ZN(n4409) );
  AOI21_X1 U3941 ( .B1(n4404), .B2(n4900), .A(n3082), .ZN(n3088) );
  INV_X1 U3942 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3083) );
  OAI21_X1 U3943 ( .B1(n2022), .B2(n4406), .A(n3084), .ZN(n4405) );
  NAND2_X1 U3944 ( .A1(n3086), .A2(n3085), .ZN(U3546) );
  INV_X1 U3945 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U3946 ( .A1(n3090), .A2(n3089), .ZN(U3514) );
  INV_X1 U3947 ( .A(n3245), .ZN(n3091) );
  AND2_X2 U3948 ( .A1(n4873), .A2(n3091), .ZN(U4043) );
  NAND3_X1 U3949 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n3093), 
        .ZN(n3095) );
  INV_X1 U3950 ( .A(DATAI_31_), .ZN(n3094) );
  OAI22_X1 U3951 ( .A1(n3092), .A2(n3095), .B1(STATE_REG_SCAN_IN), .B2(n3094), 
        .ZN(U3321) );
  MUX2_X1 U3952 ( .A(n2554), .B(n3119), .S(STATE_REG_SCAN_IN), .Z(n3096) );
  INV_X1 U3953 ( .A(n3096), .ZN(U3349) );
  NAND2_X1 U3954 ( .A1(n3097), .A2(STATE_REG_SCAN_IN), .ZN(n3098) );
  OAI21_X1 U3955 ( .B1(STATE_REG_SCAN_IN), .B2(n2789), .A(n3098), .ZN(U3323)
         );
  MUX2_X1 U3956 ( .A(n3099), .B(n3140), .S(STATE_REG_SCAN_IN), .Z(n3100) );
  INV_X1 U3957 ( .A(n3100), .ZN(U3346) );
  NAND2_X1 U3958 ( .A1(n3101), .A2(STATE_REG_SCAN_IN), .ZN(n3102) );
  OAI21_X1 U3959 ( .B1(STATE_REG_SCAN_IN), .B2(n2759), .A(n3102), .ZN(U3326)
         );
  MUX2_X1 U3960 ( .A(n3103), .B(n3330), .S(STATE_REG_SCAN_IN), .Z(n3104) );
  INV_X1 U3961 ( .A(n3104), .ZN(U3344) );
  NAND2_X1 U3962 ( .A1(n3105), .A2(STATE_REG_SCAN_IN), .ZN(n3106) );
  OAI21_X1 U3963 ( .B1(STATE_REG_SCAN_IN), .B2(n2747), .A(n3106), .ZN(U3327)
         );
  NAND2_X1 U3964 ( .A1(n4356), .A2(STATE_REG_SCAN_IN), .ZN(n3107) );
  OAI21_X1 U3965 ( .B1(STATE_REG_SCAN_IN), .B2(n2664), .A(n3107), .ZN(U3335)
         );
  NAND2_X1 U3966 ( .A1(n2807), .A2(STATE_REG_SCAN_IN), .ZN(n3108) );
  OAI21_X1 U3967 ( .B1(STATE_REG_SCAN_IN), .B2(n2709), .A(n3108), .ZN(U3330)
         );
  NAND2_X1 U3968 ( .A1(n3109), .A2(STATE_REG_SCAN_IN), .ZN(n3110) );
  OAI21_X1 U3969 ( .B1(STATE_REG_SCAN_IN), .B2(n2740), .A(n3110), .ZN(U3328)
         );
  INV_X1 U3970 ( .A(D_REG_0__SCAN_IN), .ZN(n3115) );
  AND2_X1 U3971 ( .A1(n4873), .A2(n3112), .ZN(n3114) );
  AOI22_X1 U3972 ( .A1(n4870), .A2(n3115), .B1(n3114), .B2(n3113), .ZN(U3458)
         );
  INV_X1 U3973 ( .A(n3177), .ZN(n3116) );
  AOI22_X1 U3974 ( .A1(n4870), .A2(n3117), .B1(n3116), .B2(n4873), .ZN(U3459)
         );
  XNOR2_X1 U3975 ( .A(n3118), .B(REG2_REG_3__SCAN_IN), .ZN(n3125) );
  INV_X1 U3976 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4853) );
  NOR2_X1 U3977 ( .A1(STATE_REG_SCAN_IN), .A2(n4853), .ZN(n3253) );
  NOR2_X1 U3978 ( .A1(n4852), .A2(n3119), .ZN(n3120) );
  AOI211_X1 U3979 ( .C1(n4846), .C2(ADDR_REG_3__SCAN_IN), .A(n3253), .B(n3120), 
        .ZN(n3124) );
  OAI211_X1 U3980 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3122), .A(n4847), .B(n3121), 
        .ZN(n3123) );
  OAI211_X1 U3981 ( .C1(n3125), .C2(n4840), .A(n3124), .B(n3123), .ZN(U3243)
         );
  AOI211_X1 U3982 ( .C1(n2058), .C2(n3127), .A(n4360), .B(n3126), .ZN(n3135)
         );
  INV_X1 U3983 ( .A(n4819), .ZN(n3133) );
  OAI211_X1 U3984 ( .C1(n3130), .C2(n3129), .A(n4342), .B(n3128), .ZN(n3132)
         );
  AND2_X1 U3985 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3396) );
  AOI21_X1 U3986 ( .B1(n4846), .B2(ADDR_REG_5__SCAN_IN), .A(n3396), .ZN(n3131)
         );
  OAI211_X1 U3987 ( .C1(n4852), .C2(n3133), .A(n3132), .B(n3131), .ZN(n3134)
         );
  OR2_X1 U3988 ( .A1(n3135), .A2(n3134), .ZN(U3245) );
  NOR2_X1 U3989 ( .A1(n4846), .A2(U4043), .ZN(U3148) );
  XNOR2_X1 U3990 ( .A(n3136), .B(REG2_REG_6__SCAN_IN), .ZN(n3145) );
  AOI21_X1 U3991 ( .B1(n3138), .B2(n3137), .A(n4360), .ZN(n3143) );
  AND2_X1 U3992 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3442) );
  AOI21_X1 U3993 ( .B1(n4846), .B2(ADDR_REG_6__SCAN_IN), .A(n3442), .ZN(n3139)
         );
  OAI21_X1 U3994 ( .B1(n4852), .B2(n3140), .A(n3139), .ZN(n3141) );
  AOI21_X1 U3995 ( .B1(n3143), .B2(n3142), .A(n3141), .ZN(n3144) );
  OAI21_X1 U3996 ( .B1(n3145), .B2(n4840), .A(n3144), .ZN(U3246) );
  NAND2_X1 U3997 ( .A1(U4043), .A2(n3599), .ZN(n3146) );
  OAI21_X1 U3998 ( .B1(U4043), .B2(n3147), .A(n3146), .ZN(U3557) );
  NAND2_X1 U3999 ( .A1(U4043), .A2(n4149), .ZN(n3148) );
  OAI21_X1 U4000 ( .B1(U4043), .B2(n3149), .A(n3148), .ZN(U3550) );
  NAND2_X1 U4001 ( .A1(U4043), .A2(n4739), .ZN(n3150) );
  OAI21_X1 U4002 ( .B1(U4043), .B2(n3151), .A(n3150), .ZN(U3561) );
  NAND2_X1 U4003 ( .A1(U4043), .A2(n4253), .ZN(n3152) );
  OAI21_X1 U4004 ( .B1(U4043), .B2(n3153), .A(n3152), .ZN(U3551) );
  NAND2_X1 U4005 ( .A1(n4716), .A2(U4043), .ZN(n3154) );
  OAI21_X1 U4006 ( .B1(U4043), .B2(n3155), .A(n3154), .ZN(U3564) );
  NAND2_X1 U4007 ( .A1(n4507), .A2(U4043), .ZN(n3156) );
  OAI21_X1 U4008 ( .B1(n3157), .B2(U4043), .A(n3156), .ZN(U3571) );
  NAND2_X1 U4009 ( .A1(n4593), .A2(U4043), .ZN(n3158) );
  OAI21_X1 U4010 ( .B1(U4043), .B2(n3159), .A(n3158), .ZN(U3569) );
  OR2_X1 U4011 ( .A1(n3162), .A2(n3161), .ZN(n3163) );
  AND2_X1 U4012 ( .A1(n3160), .A2(n3163), .ZN(n3493) );
  INV_X1 U4013 ( .A(n4555), .ZN(n3473) );
  NAND2_X1 U4014 ( .A1(n3493), .A2(n3473), .ZN(n3172) );
  OR2_X1 U4015 ( .A1(n4726), .A2(n3165), .ZN(n3167) );
  NAND2_X1 U4016 ( .A1(n4738), .A2(n4149), .ZN(n3166) );
  OAI211_X1 U4017 ( .C1(n4741), .C2(n3164), .A(n3167), .B(n3166), .ZN(n3168)
         );
  INV_X1 U4018 ( .A(n3168), .ZN(n3171) );
  XNOR2_X1 U4019 ( .A(n3161), .B(n3819), .ZN(n3169) );
  NAND2_X1 U4020 ( .A1(n3169), .A2(n4590), .ZN(n3170) );
  AND3_X1 U4021 ( .A1(n3172), .A2(n3171), .A3(n3170), .ZN(n3497) );
  INV_X1 U4022 ( .A(n3173), .ZN(n3174) );
  AOI21_X1 U4023 ( .B1(n3456), .B2(n3261), .A(n3174), .ZN(n3495) );
  AOI22_X1 U4024 ( .A1(n3493), .A2(n4896), .B1(n3495), .B2(n4597), .ZN(n3175)
         );
  AND2_X1 U4025 ( .A1(n3497), .A2(n3175), .ZN(n4887) );
  NAND2_X1 U4026 ( .A1(n4912), .A2(REG1_REG_1__SCAN_IN), .ZN(n3176) );
  OAI21_X1 U4027 ( .B1(n4887), .B2(n4912), .A(n3176), .ZN(U3519) );
  NAND3_X1 U4028 ( .A1(n3452), .A2(n3180), .A3(n3179), .ZN(n3206) );
  AND2_X2 U4029 ( .A1(n3462), .A2(n3245), .ZN(n3267) );
  INV_X1 U4030 ( .A(n3255), .ZN(n3183) );
  NAND3_X1 U4031 ( .A1(n4078), .A2(n4873), .A3(n3183), .ZN(n3972) );
  OR2_X1 U4032 ( .A1(n3206), .A2(n3972), .ZN(n3251) );
  NAND2_X1 U4033 ( .A1(n3457), .A2(n3184), .ZN(n3187) );
  INV_X1 U4034 ( .A(n3185), .ZN(n3186) );
  NAND2_X1 U4035 ( .A1(n3187), .A2(n3186), .ZN(n3193) );
  NAND2_X1 U4036 ( .A1(n3193), .A2(n4741), .ZN(n3188) );
  NAND2_X1 U4037 ( .A1(n3206), .A2(n3188), .ZN(n3189) );
  NAND2_X1 U4038 ( .A1(n3189), .A2(n3451), .ZN(n3248) );
  INV_X1 U4039 ( .A(n3248), .ZN(n3192) );
  INV_X1 U4040 ( .A(n3972), .ZN(n3190) );
  NAND2_X1 U4041 ( .A1(n3206), .A2(n3190), .ZN(n3249) );
  NAND3_X1 U4042 ( .A1(n3192), .A2(n3191), .A3(n3249), .ZN(n4254) );
  NAND2_X1 U40430 ( .A1(n4254), .A2(REG3_REG_0__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4044 ( .A1(n3267), .A2(n3456), .ZN(n3195) );
  NAND2_X1 U4045 ( .A1(n3267), .A2(n4149), .ZN(n3198) );
  NAND2_X1 U4046 ( .A1(n4079), .A2(n3456), .ZN(n3197) );
  NAND2_X1 U4047 ( .A1(n3198), .A2(n3197), .ZN(n3257) );
  NAND2_X1 U4048 ( .A1(n3204), .A2(n3257), .ZN(n3200) );
  OR2_X1 U4049 ( .A1(n3245), .A2(n4316), .ZN(n3199) );
  NAND2_X1 U4050 ( .A1(n3200), .A2(n3199), .ZN(n3254) );
  NOR2_X1 U4051 ( .A1(n2379), .A2(REG1_REG_0__SCAN_IN), .ZN(n3201) );
  NOR2_X1 U4052 ( .A1(n3245), .A2(n3201), .ZN(n3202) );
  OR2_X1 U4053 ( .A1(n3257), .A2(n3202), .ZN(n3203) );
  NOR2_X1 U4054 ( .A1(n3204), .A2(n3203), .ZN(n3205) );
  NOR2_X1 U4055 ( .A1(n3254), .A2(n3205), .ZN(n3227) );
  OR3_X1 U4056 ( .A1(n3206), .A2(n3449), .A3(n4741), .ZN(n3208) );
  NOR2_X1 U4057 ( .A1(n3449), .A2(n2862), .ZN(n3207) );
  AOI22_X1 U4058 ( .A1(n4250), .A2(n3227), .B1(n4288), .B2(n3456), .ZN(n3209)
         );
  OAI211_X1 U4059 ( .C1(n3211), .C2(n4291), .A(n3210), .B(n3209), .ZN(U3229)
         );
  NAND2_X1 U4060 ( .A1(n4496), .A2(U4043), .ZN(n3212) );
  OAI21_X1 U4061 ( .B1(U4043), .B2(n3213), .A(n3212), .ZN(U3572) );
  MUX2_X1 U4062 ( .A(REG1_REG_7__SCAN_IN), .B(n4913), .S(n4818), .Z(n3215) );
  XOR2_X1 U4063 ( .A(n3215), .B(n3214), .Z(n3223) );
  OAI211_X1 U4064 ( .C1(n3218), .C2(n3217), .A(n3216), .B(n4342), .ZN(n3220)
         );
  AND2_X1 U4065 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3487) );
  AOI21_X1 U4066 ( .B1(n4846), .B2(ADDR_REG_7__SCAN_IN), .A(n3487), .ZN(n3219)
         );
  OAI211_X1 U4067 ( .C1(n4852), .C2(n3221), .A(n3220), .B(n3219), .ZN(n3222)
         );
  AOI21_X1 U4068 ( .B1(n3223), .B2(n4847), .A(n3222), .ZN(n3224) );
  INV_X1 U4069 ( .A(n3224), .ZN(U3247) );
  OR2_X1 U4070 ( .A1(n4824), .A2(REG2_REG_0__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4071 ( .A1(n3226), .A2(n3225), .ZN(n4823) );
  NAND2_X1 U4072 ( .A1(n2379), .A2(REG2_REG_0__SCAN_IN), .ZN(n4318) );
  OAI21_X1 U4073 ( .B1(n4318), .B2(n3971), .A(U4043), .ZN(n3229) );
  NOR3_X1 U4074 ( .A1(n3227), .A2(n4810), .A3(n4822), .ZN(n3228) );
  INV_X1 U4075 ( .A(n2010), .ZN(n3243) );
  INV_X1 U4076 ( .A(n3230), .ZN(n3235) );
  INV_X1 U4077 ( .A(n3231), .ZN(n3234) );
  INV_X1 U4078 ( .A(n3232), .ZN(n3233) );
  AOI211_X1 U4079 ( .C1(n3235), .C2(n3234), .A(n3233), .B(n4840), .ZN(n3240)
         );
  AOI211_X1 U4080 ( .C1(n3238), .C2(n3237), .A(n3236), .B(n4360), .ZN(n3239)
         );
  NOR2_X1 U4081 ( .A1(n3240), .A2(n3239), .ZN(n3242) );
  AOI22_X1 U4082 ( .A1(n4846), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3241) );
  OAI211_X1 U4083 ( .C1(n3243), .C2(n4852), .A(n3242), .B(n3241), .ZN(n3244)
         );
  OR2_X1 U4084 ( .A1(n3298), .A2(n3244), .ZN(U3242) );
  NAND2_X1 U4085 ( .A1(n3246), .A2(n3245), .ZN(n3247) );
  OAI21_X1 U4086 ( .B1(n3248), .B2(n3247), .A(STATE_REG_SCAN_IN), .ZN(n3250)
         );
  OAI22_X1 U4087 ( .A1(n3165), .A2(n4267), .B1(n4291), .B2(n3555), .ZN(n3252)
         );
  AOI211_X1 U4088 ( .C1(n3340), .C2(n4288), .A(n3253), .B(n3252), .ZN(n3289)
         );
  INV_X1 U4089 ( .A(n3254), .ZN(n3259) );
  NAND2_X1 U4090 ( .A1(n3267), .A2(n4253), .ZN(n3263) );
  NAND2_X1 U4091 ( .A1(n4079), .A2(n3261), .ZN(n3262) );
  NAND2_X1 U4092 ( .A1(n3263), .A2(n3262), .ZN(n3265) );
  INV_X1 U4093 ( .A(n3282), .ZN(n3266) );
  NAND2_X1 U4094 ( .A1(n3266), .A2(n4253), .ZN(n3269) );
  NAND2_X1 U4095 ( .A1(n3267), .A2(n3261), .ZN(n3268) );
  NAND2_X1 U4096 ( .A1(n3269), .A2(n3268), .ZN(n3270) );
  XNOR2_X1 U4097 ( .A(n3271), .B(n3270), .ZN(n4150) );
  INV_X1 U4098 ( .A(n3270), .ZN(n3272) );
  AOI21_X1 U4099 ( .B1(n4151), .B2(n4150), .A(n3273), .ZN(n4249) );
  OR2_X1 U4100 ( .A1(n3282), .A2(n3165), .ZN(n3275) );
  NAND2_X1 U4101 ( .A1(n2129), .A2(n2013), .ZN(n3274) );
  NAND2_X1 U4102 ( .A1(n3275), .A2(n3274), .ZN(n3280) );
  NAND2_X1 U4103 ( .A1(n4079), .A2(n2013), .ZN(n3276) );
  XNOR2_X1 U4104 ( .A(n3277), .B(n4087), .ZN(n3278) );
  XNOR2_X1 U4105 ( .A(n3280), .B(n3278), .ZN(n4248) );
  NAND2_X1 U4106 ( .A1(n4249), .A2(n4248), .ZN(n4247) );
  INV_X1 U4107 ( .A(n3278), .ZN(n3279) );
  OR2_X1 U4108 ( .A1(n3280), .A2(n3279), .ZN(n3281) );
  NAND2_X1 U4109 ( .A1(n4247), .A2(n3281), .ZN(n3376) );
  INV_X2 U4110 ( .A(n3266), .ZN(n3798) );
  OR2_X1 U4111 ( .A1(n3798), .A2(n3361), .ZN(n3284) );
  NAND2_X1 U4112 ( .A1(n3267), .A2(n3340), .ZN(n3283) );
  NAND2_X1 U4113 ( .A1(n3284), .A2(n3283), .ZN(n3379) );
  NAND2_X1 U4114 ( .A1(n4079), .A2(n3340), .ZN(n3285) );
  OAI21_X1 U4115 ( .B1(n3361), .B2(n3383), .A(n3285), .ZN(n3286) );
  XNOR2_X1 U4116 ( .A(n3286), .B(n4087), .ZN(n3377) );
  XNOR2_X1 U4117 ( .A(n3379), .B(n3377), .ZN(n3375) );
  XNOR2_X1 U4118 ( .A(n3376), .B(n3375), .ZN(n3287) );
  NAND2_X1 U4119 ( .A1(n3287), .A2(n4250), .ZN(n3288) );
  OAI211_X1 U4120 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4276), .A(n3289), .B(n3288), 
        .ZN(U3215) );
  XNOR2_X1 U4121 ( .A(n3290), .B(REG2_REG_4__SCAN_IN), .ZN(n3300) );
  AOI211_X1 U4122 ( .C1(n4910), .C2(n3292), .A(n4360), .B(n3291), .ZN(n3297)
         );
  NAND2_X1 U4123 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3414) );
  INV_X1 U4124 ( .A(n3414), .ZN(n3293) );
  AOI21_X1 U4125 ( .B1(n4846), .B2(ADDR_REG_4__SCAN_IN), .A(n3293), .ZN(n3294)
         );
  OAI21_X1 U4126 ( .B1(n4852), .B2(n3295), .A(n3294), .ZN(n3296) );
  NOR3_X1 U4127 ( .A1(n3298), .A2(n3297), .A3(n3296), .ZN(n3299) );
  OAI21_X1 U4128 ( .B1(n3300), .B2(n4840), .A(n3299), .ZN(U3244) );
  NAND2_X1 U4129 ( .A1(n3835), .A2(n3845), .ZN(n3910) );
  XOR2_X1 U4130 ( .A(n3301), .B(n3910), .Z(n3591) );
  NAND2_X1 U4131 ( .A1(n3303), .A2(n3304), .ZN(n3318) );
  NAND2_X1 U4132 ( .A1(n3318), .A2(n3305), .ZN(n3307) );
  NAND2_X1 U4133 ( .A1(n3307), .A2(n3306), .ZN(n3578) );
  XNOR2_X1 U4134 ( .A(n3578), .B(n3910), .ZN(n3602) );
  INV_X1 U4135 ( .A(n4726), .ZN(n4737) );
  OAI22_X1 U4136 ( .A1(n4707), .A2(n3596), .B1(n4741), .B2(n3595), .ZN(n3308)
         );
  AOI21_X1 U4137 ( .B1(n4737), .B2(n3599), .A(n3308), .ZN(n3309) );
  OAI21_X1 U4138 ( .B1(n3602), .B2(n4678), .A(n3309), .ZN(n3310) );
  AOI21_X1 U4139 ( .B1(n3591), .B2(n4590), .A(n3310), .ZN(n3371) );
  NOR2_X1 U4140 ( .A1(n3311), .A2(n3595), .ZN(n3312) );
  OR2_X1 U4141 ( .A1(n3565), .A2(n3312), .ZN(n3594) );
  INV_X1 U4142 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3313) );
  OAI22_X1 U4143 ( .A1(n3594), .A2(n4807), .B1(n4907), .B2(n3313), .ZN(n3314)
         );
  INV_X1 U4144 ( .A(n3314), .ZN(n3315) );
  OAI21_X1 U4145 ( .B1(n3371), .B2(n4905), .A(n3315), .ZN(U3479) );
  INV_X1 U4146 ( .A(n3833), .ZN(n3316) );
  NAND2_X1 U4147 ( .A1(n3316), .A2(n3844), .ZN(n3891) );
  INV_X1 U4148 ( .A(n3891), .ZN(n3317) );
  XNOR2_X1 U4149 ( .A(n3318), .B(n3317), .ZN(n3550) );
  AOI22_X1 U4150 ( .A1(n4724), .A2(n3397), .B1(n4310), .B2(n4738), .ZN(n3319)
         );
  OAI21_X1 U4151 ( .B1(n3579), .B2(n4726), .A(n3319), .ZN(n3322) );
  XOR2_X1 U4152 ( .A(n3320), .B(n3891), .Z(n3321) );
  NOR2_X1 U4153 ( .A1(n3321), .A2(n4631), .ZN(n3553) );
  AOI211_X1 U4154 ( .C1(n3550), .C2(n4900), .A(n3322), .B(n3553), .ZN(n3372)
         );
  AND2_X1 U4155 ( .A1(n3466), .A2(n3397), .ZN(n3323) );
  OR2_X1 U4156 ( .A1(n3323), .A2(n3311), .ZN(n3559) );
  INV_X1 U4157 ( .A(REG0_REG_5__SCAN_IN), .ZN(n3324) );
  OAI22_X1 U4158 ( .A1(n4807), .A2(n3559), .B1(n4907), .B2(n3324), .ZN(n3325)
         );
  INV_X1 U4159 ( .A(n3325), .ZN(n3326) );
  OAI21_X1 U4160 ( .B1(n3372), .B2(n4905), .A(n3326), .ZN(U3477) );
  XNOR2_X1 U4161 ( .A(n3327), .B(REG1_REG_8__SCAN_IN), .ZN(n3334) );
  XOR2_X1 U4162 ( .A(n3328), .B(REG2_REG_8__SCAN_IN), .Z(n3332) );
  NAND2_X1 U4163 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n3545) );
  NAND2_X1 U4164 ( .A1(n4846), .A2(ADDR_REG_8__SCAN_IN), .ZN(n3329) );
  OAI211_X1 U4165 ( .C1(n4852), .C2(n3330), .A(n3545), .B(n3329), .ZN(n3331)
         );
  AOI21_X1 U4166 ( .B1(n3332), .B2(n4342), .A(n3331), .ZN(n3333) );
  OAI21_X1 U4167 ( .B1(n3334), .B2(n4360), .A(n3333), .ZN(U3248) );
  NAND2_X1 U4168 ( .A1(n3160), .A2(n3335), .ZN(n3352) );
  OR2_X1 U4169 ( .A1(n3352), .A2(n3913), .ZN(n3353) );
  INV_X1 U4170 ( .A(n3336), .ZN(n3337) );
  NAND2_X1 U4171 ( .A1(n3353), .A2(n3337), .ZN(n3338) );
  XNOR2_X1 U4172 ( .A(n3338), .B(n3912), .ZN(n3342) );
  INV_X1 U4173 ( .A(n3342), .ZN(n4854) );
  XNOR2_X1 U4174 ( .A(n3339), .B(n3912), .ZN(n3345) );
  AOI22_X1 U4175 ( .A1(n4724), .A2(n3340), .B1(n4310), .B2(n4737), .ZN(n3341)
         );
  OAI21_X1 U4176 ( .B1(n3165), .B2(n4707), .A(n3341), .ZN(n3344) );
  NOR2_X1 U4177 ( .A1(n3342), .A2(n4555), .ZN(n3343) );
  AOI211_X1 U4178 ( .C1(n3345), .C2(n4590), .A(n3344), .B(n3343), .ZN(n4858)
         );
  INV_X1 U4179 ( .A(n4858), .ZN(n3346) );
  AOI21_X1 U4180 ( .B1(n4896), .B2(n4854), .A(n3346), .ZN(n3368) );
  INV_X1 U4181 ( .A(n4807), .ZN(n4889) );
  OR2_X1 U4182 ( .A1(n3348), .A2(n3349), .ZN(n3350) );
  AND2_X1 U4183 ( .A1(n3347), .A2(n3350), .ZN(n4855) );
  AOI22_X1 U4184 ( .A1(n4889), .A2(n4855), .B1(REG0_REG_3__SCAN_IN), .B2(n4905), .ZN(n3351) );
  OAI21_X1 U4185 ( .B1(n3368), .B2(n4905), .A(n3351), .ZN(U3473) );
  INV_X1 U4186 ( .A(n3352), .ZN(n3355) );
  OAI21_X1 U4187 ( .B1(n3355), .B2(n3354), .A(n3353), .ZN(n4860) );
  INV_X1 U4188 ( .A(n4860), .ZN(n3364) );
  OAI21_X1 U4189 ( .B1(n3913), .B2(n3357), .A(n3356), .ZN(n3358) );
  NAND2_X1 U4190 ( .A1(n3358), .A2(n4590), .ZN(n3360) );
  AOI22_X1 U4191 ( .A1(n2013), .A2(n4724), .B1(n4253), .B2(n4738), .ZN(n3359)
         );
  OAI211_X1 U4192 ( .C1(n3361), .C2(n4726), .A(n3360), .B(n3359), .ZN(n3362)
         );
  AOI21_X1 U4193 ( .B1(n3473), .B2(n4860), .A(n3362), .ZN(n4865) );
  OAI21_X1 U4194 ( .B1(n3364), .B2(n3363), .A(n4865), .ZN(n4890) );
  INV_X1 U4195 ( .A(n4890), .ZN(n3366) );
  AOI21_X1 U4196 ( .B1(n2013), .B2(n3173), .A(n3348), .ZN(n4888) );
  AOI22_X1 U4197 ( .A1(n2901), .A2(n4888), .B1(REG1_REG_2__SCAN_IN), .B2(n4912), .ZN(n3365) );
  OAI21_X1 U4198 ( .B1(n3366), .B2(n4912), .A(n3365), .ZN(U3520) );
  AOI22_X1 U4199 ( .A1(n2901), .A2(n4855), .B1(REG1_REG_3__SCAN_IN), .B2(n4912), .ZN(n3367) );
  OAI21_X1 U4200 ( .B1(n3368), .B2(n4912), .A(n3367), .ZN(U3521) );
  INV_X1 U4201 ( .A(n3594), .ZN(n3369) );
  AOI22_X1 U4202 ( .A1(n3369), .A2(n2901), .B1(n4912), .B2(REG1_REG_6__SCAN_IN), .ZN(n3370) );
  OAI21_X1 U4203 ( .B1(n3371), .B2(n4912), .A(n3370), .ZN(U3524) );
  MUX2_X1 U4204 ( .A(n3373), .B(n3372), .S(n4915), .Z(n3374) );
  OAI21_X1 U4205 ( .B1(n4746), .B2(n3559), .A(n3374), .ZN(U3523) );
  INV_X1 U4206 ( .A(n3377), .ZN(n3378) );
  OR2_X1 U4207 ( .A1(n3379), .A2(n3378), .ZN(n3380) );
  OR2_X1 U4208 ( .A1(n3798), .A2(n3555), .ZN(n3382) );
  NAND2_X1 U4209 ( .A1(n2129), .A2(n3470), .ZN(n3381) );
  NAND2_X1 U4210 ( .A1(n3382), .A2(n3381), .ZN(n3388) );
  NAND2_X1 U4211 ( .A1(n4079), .A2(n3470), .ZN(n3384) );
  OAI21_X1 U4212 ( .B1(n3555), .B2(n3383), .A(n3384), .ZN(n3385) );
  XNOR2_X1 U4213 ( .A(n3385), .B(n4043), .ZN(n3387) );
  XNOR2_X1 U4214 ( .A(n3388), .B(n3387), .ZN(n3419) );
  NAND2_X1 U4215 ( .A1(n3388), .A2(n3387), .ZN(n3389) );
  NAND2_X1 U4216 ( .A1(n3417), .A2(n3389), .ZN(n3395) );
  INV_X1 U4217 ( .A(n3798), .ZN(n4018) );
  OR2_X1 U4218 ( .A1(n3798), .A2(n3596), .ZN(n3391) );
  NAND2_X1 U4219 ( .A1(n4078), .A2(n3397), .ZN(n3390) );
  NAND2_X1 U4220 ( .A1(n3391), .A2(n3390), .ZN(n3435) );
  NAND2_X1 U4221 ( .A1(n4079), .A2(n3397), .ZN(n3392) );
  XNOR2_X1 U4222 ( .A(n3393), .B(n4087), .ZN(n3433) );
  XNOR2_X1 U4223 ( .A(n3435), .B(n3433), .ZN(n3394) );
  OAI211_X1 U4224 ( .C1(n3395), .C2(n3394), .A(n3437), .B(n4250), .ZN(n3402)
         );
  NAND2_X1 U4225 ( .A1(n4287), .A2(n4310), .ZN(n3399) );
  AOI21_X1 U4226 ( .B1(n4288), .B2(n3397), .A(n3396), .ZN(n3398) );
  OAI211_X1 U4227 ( .C1(n3579), .C2(n4291), .A(n3399), .B(n3398), .ZN(n3400)
         );
  AOI21_X1 U4228 ( .B1(n4294), .B2(n3556), .A(n3400), .ZN(n3401) );
  NAND2_X1 U4229 ( .A1(n3402), .A2(n3401), .ZN(U3224) );
  XNOR2_X1 U4230 ( .A(n3404), .B(n3403), .ZN(n3413) );
  AOI21_X1 U4231 ( .B1(n3406), .B2(n3405), .A(n4360), .ZN(n3411) );
  AND2_X1 U4232 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3655) );
  AOI21_X1 U4233 ( .B1(n4846), .B2(ADDR_REG_9__SCAN_IN), .A(n3655), .ZN(n3407)
         );
  OAI21_X1 U4234 ( .B1(n4852), .B2(n3408), .A(n3407), .ZN(n3409) );
  AOI21_X1 U4235 ( .B1(n3411), .B2(n3410), .A(n3409), .ZN(n3412) );
  OAI21_X1 U4236 ( .B1(n3413), .B2(n4840), .A(n3412), .ZN(U3249) );
  AOI22_X1 U4237 ( .A1(n4262), .A2(n4309), .B1(n4287), .B2(n4311), .ZN(n3415)
         );
  OAI211_X1 U4238 ( .C1(n4241), .C2(n2561), .A(n3415), .B(n3414), .ZN(n3421)
         );
  INV_X1 U4239 ( .A(n3417), .ZN(n3418) );
  AOI211_X1 U4240 ( .C1(n3419), .C2(n3416), .A(n4296), .B(n3418), .ZN(n3420)
         );
  AOI211_X1 U4241 ( .C1(n3477), .C2(n4294), .A(n3421), .B(n3420), .ZN(n3422)
         );
  INV_X1 U4242 ( .A(n3422), .ZN(U3227) );
  INV_X1 U4243 ( .A(n3423), .ZN(n3840) );
  AND2_X1 U4244 ( .A1(n3840), .A2(n3841), .ZN(n3902) );
  XOR2_X1 U4245 ( .A(n3424), .B(n3902), .Z(n3621) );
  XOR2_X1 U4246 ( .A(n3425), .B(n3902), .Z(n3622) );
  OAI22_X1 U4247 ( .A1(n4707), .A2(n2589), .B1(n3653), .B2(n4726), .ZN(n3426)
         );
  AOI21_X1 U4248 ( .B1(n3536), .B2(n4724), .A(n3426), .ZN(n3427) );
  OAI21_X1 U4249 ( .B1(n3622), .B2(n4678), .A(n3427), .ZN(n3428) );
  AOI21_X1 U4250 ( .B1(n3621), .B2(n4590), .A(n3428), .ZN(n3432) );
  NAND2_X1 U4251 ( .A1(n3566), .A2(n3536), .ZN(n3429) );
  AND2_X1 U4252 ( .A1(n3506), .A2(n3429), .ZN(n3624) );
  AOI22_X1 U4253 ( .A1(n3624), .A2(n2901), .B1(REG1_REG_8__SCAN_IN), .B2(n4912), .ZN(n3430) );
  OAI21_X1 U4254 ( .B1(n3432), .B2(n4912), .A(n3430), .ZN(U3526) );
  AOI22_X1 U4255 ( .A1(n3624), .A2(n4889), .B1(REG0_REG_8__SCAN_IN), .B2(n4905), .ZN(n3431) );
  OAI21_X1 U4256 ( .B1(n3432), .B2(n4905), .A(n3431), .ZN(U3483) );
  INV_X1 U4257 ( .A(n3433), .ZN(n3434) );
  NAND2_X1 U4258 ( .A1(n3435), .A2(n3434), .ZN(n3436) );
  OAI22_X1 U4259 ( .A1(n3579), .A2(n3652), .B1(n3595), .B2(n4089), .ZN(n3438)
         );
  XNOR2_X1 U4260 ( .A(n3438), .B(n4043), .ZN(n3480) );
  OR2_X1 U4261 ( .A1(n3798), .A2(n3579), .ZN(n3440) );
  NAND2_X1 U4262 ( .A1(n4078), .A2(n3443), .ZN(n3439) );
  NAND2_X1 U4263 ( .A1(n3440), .A2(n3439), .ZN(n3481) );
  XOR2_X1 U4264 ( .A(n3480), .B(n3481), .Z(n3441) );
  XNOR2_X1 U4265 ( .A(n3482), .B(n3441), .ZN(n3448) );
  NAND2_X1 U4266 ( .A1(n4262), .A2(n3599), .ZN(n3445) );
  AOI21_X1 U4267 ( .B1(n4288), .B2(n3443), .A(n3442), .ZN(n3444) );
  OAI211_X1 U4268 ( .C1(n3596), .C2(n4267), .A(n3445), .B(n3444), .ZN(n3446)
         );
  AOI21_X1 U4269 ( .B1(n4294), .B2(n3592), .A(n3446), .ZN(n3447) );
  OAI21_X1 U4270 ( .B1(n3448), .B2(n4296), .A(n3447), .ZN(U3236) );
  OAI21_X1 U4271 ( .B1(n3449), .B2(n3117), .A(n4870), .ZN(n3450) );
  NAND4_X1 U4272 ( .A1(n3453), .A2(n3452), .A3(n3451), .A4(n3450), .ZN(n3454)
         );
  INV_X1 U4273 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3465) );
  INV_X1 U4274 ( .A(n3455), .ZN(n3460) );
  NAND2_X1 U4275 ( .A1(n3457), .A2(n3456), .ZN(n4880) );
  NAND2_X1 U4276 ( .A1(n3458), .A2(n4149), .ZN(n3821) );
  NAND2_X1 U4277 ( .A1(n3821), .A2(n3819), .ZN(n4884) );
  NAND2_X1 U4278 ( .A1(n4555), .A2(n4631), .ZN(n3459) );
  AOI22_X1 U4279 ( .A1(n4884), .A2(n3459), .B1(n4737), .B2(n4253), .ZN(n4881)
         );
  OAI21_X1 U4280 ( .B1(n3460), .B2(n4880), .A(n4881), .ZN(n3461) );
  AOI22_X1 U4281 ( .A1(n4556), .A2(n3461), .B1(REG3_REG_0__SCAN_IN), .B2(n4859), .ZN(n3464) );
  NAND2_X1 U4282 ( .A1(n3462), .A2(n3181), .ZN(n3551) );
  NAND2_X1 U4283 ( .A1(n4861), .A2(n4884), .ZN(n3463) );
  OAI211_X1 U4284 ( .C1(n4556), .C2(n3465), .A(n3464), .B(n3463), .ZN(U3290)
         );
  OAI211_X1 U4285 ( .C1(n2892), .C2(n2561), .A(n4597), .B(n3466), .ZN(n4893)
         );
  NOR2_X1 U4286 ( .A1(n4893), .A2(n3181), .ZN(n3476) );
  XOR2_X1 U4287 ( .A(n3467), .B(n3894), .Z(n3475) );
  INV_X1 U4288 ( .A(n3303), .ZN(n3469) );
  AOI21_X1 U4289 ( .B1(n3894), .B2(n3468), .A(n3469), .ZN(n4897) );
  AOI22_X1 U4290 ( .A1(n4724), .A2(n3470), .B1(n4738), .B2(n4311), .ZN(n3471)
         );
  OAI21_X1 U4291 ( .B1(n3596), .B2(n4726), .A(n3471), .ZN(n3472) );
  AOI21_X1 U4292 ( .B1(n4897), .B2(n3473), .A(n3472), .ZN(n3474) );
  OAI21_X1 U4293 ( .B1(n3475), .B2(n4631), .A(n3474), .ZN(n4894) );
  AOI211_X1 U4294 ( .C1(n4859), .C2(n3477), .A(n3476), .B(n4894), .ZN(n3479)
         );
  INV_X2 U4295 ( .A(n4556), .ZN(n4646) );
  AOI22_X1 U4296 ( .A1(n4861), .A2(n4897), .B1(REG2_REG_4__SCAN_IN), .B2(n4624), .ZN(n3478) );
  OAI21_X1 U4297 ( .B1(n3479), .B2(n4646), .A(n3478), .ZN(U3286) );
  OR2_X1 U4298 ( .A1(n3798), .A2(n2589), .ZN(n3484) );
  NAND2_X1 U4299 ( .A1(n4078), .A2(n3570), .ZN(n3483) );
  NAND2_X1 U4300 ( .A1(n3484), .A2(n3483), .ZN(n3533) );
  NAND2_X1 U4301 ( .A1(n4079), .A2(n3570), .ZN(n3485) );
  OAI21_X1 U4302 ( .B1(n2589), .B2(n3652), .A(n3485), .ZN(n3486) );
  XNOR2_X1 U4303 ( .A(n3486), .B(n4087), .ZN(n3531) );
  XNOR2_X1 U4304 ( .A(n3533), .B(n3531), .ZN(n3529) );
  XNOR2_X1 U4305 ( .A(n3530), .B(n3529), .ZN(n3492) );
  NAND2_X1 U4306 ( .A1(n4287), .A2(n4308), .ZN(n3489) );
  AOI21_X1 U4307 ( .B1(n4288), .B2(n3570), .A(n3487), .ZN(n3488) );
  OAI211_X1 U4308 ( .C1(n3539), .C2(n4291), .A(n3489), .B(n3488), .ZN(n3490)
         );
  AOI21_X1 U4309 ( .B1(n4294), .B2(n3576), .A(n3490), .ZN(n3491) );
  OAI21_X1 U4310 ( .B1(n3492), .B2(n4296), .A(n3491), .ZN(U3210) );
  INV_X1 U4311 ( .A(n3493), .ZN(n3500) );
  OR2_X1 U4312 ( .A1(n4624), .A2(n3494), .ZN(n4642) );
  AOI22_X1 U4313 ( .A1(n4862), .A2(n3495), .B1(REG3_REG_1__SCAN_IN), .B2(n4859), .ZN(n3499) );
  MUX2_X1 U4314 ( .A(n3497), .B(n3496), .S(n4646), .Z(n3498) );
  OAI211_X1 U4315 ( .C1(n3500), .C2(n4566), .A(n3499), .B(n3498), .ZN(U3289)
         );
  NAND2_X1 U4316 ( .A1(n3842), .A2(n3852), .ZN(n3898) );
  XOR2_X1 U4317 ( .A(n3501), .B(n3898), .Z(n3612) );
  AOI22_X1 U4318 ( .A1(n4307), .A2(n4738), .B1(n4737), .B2(n4305), .ZN(n3502)
         );
  OAI21_X1 U4319 ( .B1(n2183), .B2(n4741), .A(n3502), .ZN(n3505) );
  XNOR2_X1 U4320 ( .A(n3503), .B(n3898), .ZN(n3504) );
  NOR2_X1 U4321 ( .A1(n3504), .A2(n4631), .ZN(n3613) );
  AOI211_X1 U4322 ( .C1(n3612), .C2(n4900), .A(n3505), .B(n3613), .ZN(n3589)
         );
  INV_X1 U4323 ( .A(n3506), .ZN(n3507) );
  OAI21_X1 U4324 ( .B1(n3507), .B2(n2183), .A(n3515), .ZN(n3615) );
  INV_X1 U4325 ( .A(n3615), .ZN(n3508) );
  AOI22_X1 U4326 ( .A1(n3508), .A2(n4889), .B1(REG0_REG_9__SCAN_IN), .B2(n4905), .ZN(n3509) );
  OAI21_X1 U4327 ( .B1(n3589), .B2(n4905), .A(n3509), .ZN(U3485) );
  NAND2_X1 U4328 ( .A1(n3849), .A2(n3850), .ZN(n3908) );
  XOR2_X1 U4329 ( .A(n3510), .B(n3908), .Z(n3604) );
  XOR2_X1 U4330 ( .A(n3511), .B(n3908), .Z(n3611) );
  OAI22_X1 U4331 ( .A1(n4707), .A2(n3653), .B1(n3751), .B2(n4726), .ZN(n3512)
         );
  AOI21_X1 U4332 ( .B1(n3741), .B2(n4724), .A(n3512), .ZN(n3513) );
  OAI21_X1 U4333 ( .B1(n3611), .B2(n4678), .A(n3513), .ZN(n3514) );
  AOI21_X1 U4334 ( .B1(n3604), .B2(n4590), .A(n3514), .ZN(n3519) );
  AND2_X1 U4335 ( .A1(n3515), .A2(n3741), .ZN(n3516) );
  NOR2_X1 U4336 ( .A1(n2049), .A2(n3516), .ZN(n3608) );
  AOI22_X1 U4337 ( .A1(n3608), .A2(n4889), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4905), .ZN(n3517) );
  OAI21_X1 U4338 ( .B1(n3519), .B2(n4905), .A(n3517), .ZN(U3487) );
  AOI22_X1 U4339 ( .A1(n3608), .A2(n2901), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4912), .ZN(n3518) );
  OAI21_X1 U4340 ( .B1(n3519), .B2(n4912), .A(n3518), .ZN(U3528) );
  XNOR2_X1 U4341 ( .A(n3520), .B(REG1_REG_10__SCAN_IN), .ZN(n3528) );
  XOR2_X1 U4342 ( .A(REG2_REG_10__SCAN_IN), .B(n3521), .Z(n3522) );
  NAND2_X1 U4343 ( .A1(n4342), .A2(n3522), .ZN(n3523) );
  NAND2_X1 U4344 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4345 ( .A1(n3523), .A2(n3784), .ZN(n3526) );
  NOR2_X1 U4346 ( .A1(n4852), .A2(n3524), .ZN(n3525) );
  AOI211_X1 U4347 ( .C1(n4846), .C2(ADDR_REG_10__SCAN_IN), .A(n3526), .B(n3525), .ZN(n3527) );
  OAI21_X1 U4348 ( .B1(n3528), .B2(n4360), .A(n3527), .ZN(U3250) );
  NAND2_X1 U4349 ( .A1(n3530), .A2(n3529), .ZN(n3535) );
  INV_X1 U4350 ( .A(n3531), .ZN(n3532) );
  NAND2_X1 U4351 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  OR2_X1 U4352 ( .A1(n3798), .A2(n3539), .ZN(n3538) );
  NAND2_X1 U4353 ( .A1(n4078), .A2(n3536), .ZN(n3537) );
  NAND2_X1 U4354 ( .A1(n3538), .A2(n3537), .ZN(n3542) );
  OAI22_X1 U4355 ( .A1(n3539), .A2(n3652), .B1(n3623), .B2(n4089), .ZN(n3540)
         );
  XNOR2_X1 U4356 ( .A(n3540), .B(n4043), .ZN(n3541) );
  INV_X1 U4357 ( .A(n3648), .ZN(n3543) );
  AND2_X1 U4358 ( .A1(n3542), .A2(n3541), .ZN(n3647) );
  NOR2_X1 U4359 ( .A1(n3543), .A2(n3647), .ZN(n3544) );
  XNOR2_X1 U4360 ( .A(n3646), .B(n3544), .ZN(n3549) );
  AOI22_X1 U4361 ( .A1(n4262), .A2(n4306), .B1(n4287), .B2(n3599), .ZN(n3546)
         );
  OAI211_X1 U4362 ( .C1(n4241), .C2(n3623), .A(n3546), .B(n3545), .ZN(n3547)
         );
  AOI21_X1 U4363 ( .B1(n3625), .B2(n4294), .A(n3547), .ZN(n3548) );
  OAI21_X1 U4364 ( .B1(n3549), .B2(n4296), .A(n3548), .ZN(U3218) );
  INV_X1 U4365 ( .A(n3550), .ZN(n3564) );
  AND2_X1 U4366 ( .A1(n4555), .A2(n3551), .ZN(n3552) );
  NAND2_X1 U4367 ( .A1(n3553), .A2(n4556), .ZN(n3563) );
  OR2_X1 U4368 ( .A1(n4624), .A2(n4726), .ZN(n4537) );
  OAI22_X1 U4369 ( .A1(n3579), .A2(n4537), .B1(n4617), .B2(n3554), .ZN(n3561)
         );
  OR2_X1 U4370 ( .A1(n4535), .A2(n3555), .ZN(n3558) );
  AOI22_X1 U4371 ( .A1(n4646), .A2(REG2_REG_5__SCAN_IN), .B1(n3556), .B2(n4859), .ZN(n3557) );
  OAI211_X1 U4372 ( .C1(n4642), .C2(n3559), .A(n3558), .B(n3557), .ZN(n3560)
         );
  NOR2_X1 U4373 ( .A1(n3561), .A2(n3560), .ZN(n3562) );
  OAI211_X1 U4374 ( .C1(n3564), .C2(n4605), .A(n3563), .B(n3562), .ZN(U3285)
         );
  INV_X1 U4375 ( .A(n3565), .ZN(n3569) );
  INV_X1 U4376 ( .A(n4597), .ZN(n3568) );
  AOI211_X1 U4377 ( .C1(n3570), .C2(n3569), .A(n3568), .B(n3567), .ZN(n4903)
         );
  XNOR2_X1 U4378 ( .A(n3571), .B(n3890), .ZN(n3575) );
  OAI22_X1 U4379 ( .A1(n4707), .A2(n3579), .B1(n4741), .B2(n3572), .ZN(n3573)
         );
  AOI21_X1 U4380 ( .B1(n4737), .B2(n4307), .A(n3573), .ZN(n3574) );
  OAI21_X1 U4381 ( .B1(n3575), .B2(n4631), .A(n3574), .ZN(n4904) );
  AOI21_X1 U4382 ( .B1(n4903), .B2(n4373), .A(n4904), .ZN(n3588) );
  AOI22_X1 U4383 ( .A1(n4646), .A2(REG2_REG_7__SCAN_IN), .B1(n3576), .B2(n4859), .ZN(n3587) );
  NAND2_X1 U4384 ( .A1(n3578), .A2(n4308), .ZN(n3577) );
  NAND2_X1 U4385 ( .A1(n3577), .A2(n3595), .ZN(n3582) );
  INV_X1 U4386 ( .A(n3578), .ZN(n3580) );
  NAND2_X1 U4387 ( .A1(n3580), .A2(n3579), .ZN(n3581) );
  AND2_X1 U4388 ( .A1(n3582), .A2(n3581), .ZN(n3583) );
  NAND2_X1 U4389 ( .A1(n3583), .A2(n3890), .ZN(n4901) );
  INV_X1 U4390 ( .A(n3583), .ZN(n3585) );
  NAND2_X1 U4391 ( .A1(n3585), .A2(n3584), .ZN(n4899) );
  NAND3_X1 U4392 ( .A1(n4901), .A2(n4644), .A3(n4899), .ZN(n3586) );
  OAI211_X1 U4393 ( .C1(n3588), .C2(n4646), .A(n3587), .B(n3586), .ZN(U3283)
         );
  MUX2_X1 U4394 ( .A(n2496), .B(n3589), .S(n4915), .Z(n3590) );
  OAI21_X1 U4395 ( .B1(n4746), .B2(n3615), .A(n3590), .ZN(U3527) );
  NAND2_X1 U4396 ( .A1(n4556), .A2(n4590), .ZN(n3719) );
  INV_X1 U4397 ( .A(n3719), .ZN(n3603) );
  NAND2_X1 U4398 ( .A1(n3591), .A2(n3603), .ZN(n3601) );
  INV_X1 U4399 ( .A(n4537), .ZN(n4613) );
  AOI22_X1 U4400 ( .A1(n4646), .A2(REG2_REG_6__SCAN_IN), .B1(n3592), .B2(n4859), .ZN(n3593) );
  OAI21_X1 U4401 ( .B1(n4642), .B2(n3594), .A(n3593), .ZN(n3598) );
  OAI22_X1 U4402 ( .A1(n3596), .A2(n4535), .B1(n4617), .B2(n3595), .ZN(n3597)
         );
  AOI211_X1 U4403 ( .C1(n4613), .C2(n3599), .A(n3598), .B(n3597), .ZN(n3600)
         );
  OAI211_X1 U4404 ( .C1(n4605), .C2(n3602), .A(n3601), .B(n3600), .ZN(U3284)
         );
  NAND2_X1 U4405 ( .A1(n3604), .A2(n3603), .ZN(n3610) );
  AOI22_X1 U4406 ( .A1(n4646), .A2(REG2_REG_10__SCAN_IN), .B1(n3792), .B2(
        n4859), .ZN(n3605) );
  OAI21_X1 U4407 ( .B1(n4535), .B2(n3653), .A(n3605), .ZN(n3607) );
  OAI22_X1 U4408 ( .A1(n3751), .A2(n4537), .B1(n4617), .B2(n2184), .ZN(n3606)
         );
  AOI211_X1 U4409 ( .C1(n3608), .C2(n4862), .A(n3607), .B(n3606), .ZN(n3609)
         );
  OAI211_X1 U4410 ( .C1(n4605), .C2(n3611), .A(n3610), .B(n3609), .ZN(U3280)
         );
  INV_X1 U4411 ( .A(n3612), .ZN(n3620) );
  NAND2_X1 U4412 ( .A1(n3613), .A2(n4556), .ZN(n3619) );
  AOI22_X1 U4413 ( .A1(n4646), .A2(REG2_REG_9__SCAN_IN), .B1(n3660), .B2(n4859), .ZN(n3614) );
  OAI21_X1 U4414 ( .B1(n4617), .B2(n2183), .A(n3614), .ZN(n3617) );
  OAI22_X1 U4415 ( .A1(n3615), .A2(n4642), .B1(n3743), .B2(n4537), .ZN(n3616)
         );
  AOI211_X1 U4416 ( .C1(n4612), .C2(n4307), .A(n3617), .B(n3616), .ZN(n3618)
         );
  OAI211_X1 U4417 ( .C1(n3620), .C2(n4605), .A(n3619), .B(n3618), .ZN(U3281)
         );
  INV_X1 U4418 ( .A(n3621), .ZN(n3632) );
  INV_X1 U4419 ( .A(n3622), .ZN(n3630) );
  OAI22_X1 U4420 ( .A1(n2589), .A2(n4535), .B1(n4617), .B2(n3623), .ZN(n3629)
         );
  NAND2_X1 U4421 ( .A1(n3624), .A2(n4862), .ZN(n3627) );
  AOI22_X1 U4422 ( .A1(n4624), .A2(REG2_REG_8__SCAN_IN), .B1(n3625), .B2(n4859), .ZN(n3626) );
  OAI211_X1 U4423 ( .C1(n3653), .C2(n4537), .A(n3627), .B(n3626), .ZN(n3628)
         );
  AOI211_X1 U4424 ( .C1(n3630), .C2(n4644), .A(n3629), .B(n3628), .ZN(n3631)
         );
  OAI21_X1 U4425 ( .B1(n3632), .B2(n3719), .A(n3631), .ZN(U3282) );
  OAI21_X1 U4426 ( .B1(n2049), .B2(n3640), .A(n3633), .ZN(n3714) );
  INV_X1 U4427 ( .A(n3636), .ZN(n3914) );
  XNOR2_X1 U4428 ( .A(n3634), .B(n3914), .ZN(n3710) );
  OAI21_X1 U4429 ( .B1(n3637), .B2(n3636), .A(n3635), .ZN(n3717) );
  NAND2_X1 U4430 ( .A1(n3717), .A2(n4900), .ZN(n3639) );
  AOI22_X1 U4431 ( .A1(n4737), .A2(n4304), .B1(n4738), .B2(n4305), .ZN(n3638)
         );
  OAI211_X1 U4432 ( .C1(n4741), .C2(n3640), .A(n3639), .B(n3638), .ZN(n3641)
         );
  AOI21_X1 U4433 ( .B1(n3710), .B2(n4590), .A(n3641), .ZN(n3643) );
  MUX2_X1 U4434 ( .A(n2991), .B(n3643), .S(n4915), .Z(n3642) );
  OAI21_X1 U4435 ( .B1(n4746), .B2(n3714), .A(n3642), .ZN(U3529) );
  INV_X1 U4436 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3644) );
  MUX2_X1 U4437 ( .A(n3644), .B(n3643), .S(n4907), .Z(n3645) );
  OAI21_X1 U4438 ( .B1(n3714), .B2(n4807), .A(n3645), .ZN(U3489) );
  OR2_X1 U4439 ( .A1(n3798), .A2(n3653), .ZN(n3650) );
  NAND2_X1 U4440 ( .A1(n4078), .A2(n3656), .ZN(n3649) );
  NAND2_X1 U4441 ( .A1(n3650), .A2(n3649), .ZN(n3736) );
  NAND2_X1 U4442 ( .A1(n4079), .A2(n3656), .ZN(n3651) );
  OAI21_X1 U4443 ( .B1(n3653), .B2(n3652), .A(n3651), .ZN(n3654) );
  XNOR2_X1 U4444 ( .A(n3654), .B(n4087), .ZN(n3734) );
  XNOR2_X1 U4445 ( .A(n3736), .B(n3734), .ZN(n3732) );
  XOR2_X1 U4446 ( .A(n3733), .B(n3732), .Z(n3662) );
  NAND2_X1 U4447 ( .A1(n4287), .A2(n4307), .ZN(n3658) );
  AOI21_X1 U4448 ( .B1(n4288), .B2(n3656), .A(n3655), .ZN(n3657) );
  OAI211_X1 U4449 ( .C1(n3743), .C2(n4291), .A(n3658), .B(n3657), .ZN(n3659)
         );
  AOI21_X1 U4450 ( .B1(n4294), .B2(n3660), .A(n3659), .ZN(n3661) );
  OAI21_X1 U4451 ( .B1(n3662), .B2(n4296), .A(n3661), .ZN(U3228) );
  INV_X1 U4452 ( .A(n3663), .ZN(n3665) );
  OR2_X1 U4453 ( .A1(n3665), .A2(n3664), .ZN(n3899) );
  NAND2_X1 U4454 ( .A1(n3667), .A2(n3666), .ZN(n3723) );
  INV_X1 U4455 ( .A(n3721), .ZN(n3668) );
  OAI21_X1 U4456 ( .B1(n3723), .B2(n3668), .A(n3722), .ZN(n3669) );
  XOR2_X1 U4457 ( .A(n3899), .B(n3669), .Z(n3672) );
  OAI22_X1 U4458 ( .A1(n4707), .A2(n3797), .B1(n4741), .B2(n3677), .ZN(n3670)
         );
  AOI21_X1 U4459 ( .B1(n4737), .B2(n4716), .A(n3670), .ZN(n3671) );
  OAI21_X1 U4460 ( .B1(n3672), .B2(n4631), .A(n3671), .ZN(n4733) );
  INV_X1 U4461 ( .A(n4733), .ZN(n3682) );
  XNOR2_X1 U4462 ( .A(n3673), .B(n3899), .ZN(n4734) );
  INV_X1 U4463 ( .A(n3675), .ZN(n3676) );
  OAI21_X1 U4464 ( .B1(n2173), .B2(n3677), .A(n3676), .ZN(n4803) );
  INV_X1 U4465 ( .A(n3678), .ZN(n4233) );
  AOI22_X1 U4466 ( .A1(n4646), .A2(REG2_REG_13__SCAN_IN), .B1(n4233), .B2(
        n4859), .ZN(n3679) );
  OAI21_X1 U4467 ( .B1(n4803), .B2(n4642), .A(n3679), .ZN(n3680) );
  AOI21_X1 U4468 ( .B1(n4734), .B2(n4644), .A(n3680), .ZN(n3681) );
  OAI21_X1 U4469 ( .B1(n3682), .B2(n4646), .A(n3681), .ZN(U3277) );
  INV_X1 U4470 ( .A(n3683), .ZN(n3684) );
  AOI211_X1 U4471 ( .C1(n3686), .C2(n3685), .A(n4360), .B(n3684), .ZN(n3694)
         );
  OAI211_X1 U4472 ( .C1(n3689), .C2(n3688), .A(n3687), .B(n4342), .ZN(n3691)
         );
  AND2_X1 U4473 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3755) );
  AOI21_X1 U4474 ( .B1(n4846), .B2(ADDR_REG_11__SCAN_IN), .A(n3755), .ZN(n3690) );
  OAI211_X1 U4475 ( .C1(n4852), .C2(n3692), .A(n3691), .B(n3690), .ZN(n3693)
         );
  OR2_X1 U4476 ( .A1(n3694), .A2(n3693), .ZN(U3251) );
  OAI21_X1 U4477 ( .B1(n3696), .B2(n3911), .A(n3695), .ZN(n4730) );
  INV_X1 U4478 ( .A(n4730), .ZN(n3709) );
  INV_X1 U4479 ( .A(n3931), .ZN(n3698) );
  INV_X1 U4480 ( .A(n3772), .ZN(n3697) );
  AOI21_X1 U4481 ( .B1(n3698), .B2(n3911), .A(n3697), .ZN(n3699) );
  OAI22_X1 U4482 ( .A1(n3699), .A2(n4631), .B1(n3709), .B2(n4555), .ZN(n4728)
         );
  NAND2_X1 U4483 ( .A1(n4728), .A2(n4556), .ZN(n3708) );
  INV_X1 U4484 ( .A(n3700), .ZN(n3701) );
  OAI21_X1 U4485 ( .B1(n3675), .B2(n3991), .A(n3701), .ZN(n4799) );
  INV_X1 U4486 ( .A(n4799), .ZN(n3706) );
  AOI22_X1 U4487 ( .A1(n4612), .A2(n4736), .B1(n4613), .B2(n4303), .ZN(n3704)
         );
  INV_X1 U4488 ( .A(n3702), .ZN(n4122) );
  AOI22_X1 U4489 ( .A1(n4646), .A2(REG2_REG_14__SCAN_IN), .B1(n4122), .B2(
        n4859), .ZN(n3703) );
  OAI211_X1 U4490 ( .C1(n3991), .C2(n4617), .A(n3704), .B(n3703), .ZN(n3705)
         );
  AOI21_X1 U4491 ( .B1(n3706), .B2(n4862), .A(n3705), .ZN(n3707) );
  OAI211_X1 U4492 ( .C1(n3709), .C2(n4566), .A(n3708), .B(n3707), .ZN(U3276)
         );
  INV_X1 U4493 ( .A(n3710), .ZN(n3720) );
  INV_X1 U4494 ( .A(n4617), .ZN(n3711) );
  AOI22_X1 U4495 ( .A1(n3711), .A2(n3756), .B1(n4613), .B2(n4304), .ZN(n3713)
         );
  AOI22_X1 U4496 ( .A1(n4624), .A2(REG2_REG_11__SCAN_IN), .B1(n3760), .B2(
        n4859), .ZN(n3712) );
  OAI211_X1 U4497 ( .C1(n3743), .C2(n4535), .A(n3713), .B(n3712), .ZN(n3716)
         );
  NOR2_X1 U4498 ( .A1(n3714), .A2(n4642), .ZN(n3715) );
  AOI211_X1 U4499 ( .C1(n3717), .C2(n4644), .A(n3716), .B(n3715), .ZN(n3718)
         );
  OAI21_X1 U4500 ( .B1(n3720), .B2(n3719), .A(n3718), .ZN(U3279) );
  AND2_X1 U4501 ( .A1(n3722), .A2(n3721), .ZN(n3916) );
  XOR2_X1 U4502 ( .A(n3916), .B(n3723), .Z(n3724) );
  NOR2_X1 U4503 ( .A1(n3724), .A2(n4631), .ZN(n4742) );
  INV_X1 U4504 ( .A(n4742), .ZN(n3731) );
  XOR2_X1 U4505 ( .A(n3725), .B(n3916), .Z(n4744) );
  AOI22_X1 U4506 ( .A1(n4612), .A2(n4739), .B1(n4613), .B2(n4736), .ZN(n3727)
         );
  AOI22_X1 U4507 ( .A1(n4624), .A2(REG2_REG_12__SCAN_IN), .B1(n3812), .B2(
        n4859), .ZN(n3726) );
  OAI211_X1 U4508 ( .C1(n2893), .C2(n4617), .A(n3727), .B(n3726), .ZN(n3729)
         );
  OAI21_X1 U4509 ( .B1(n2894), .B2(n2893), .A(n3674), .ZN(n4808) );
  NOR2_X1 U4510 ( .A1(n4808), .A2(n4642), .ZN(n3728) );
  AOI211_X1 U4511 ( .C1(n4744), .C2(n4644), .A(n3729), .B(n3728), .ZN(n3730)
         );
  OAI21_X1 U4512 ( .B1(n3731), .B2(n4646), .A(n3730), .ZN(U3278) );
  NAND2_X1 U4513 ( .A1(n3733), .A2(n3732), .ZN(n3738) );
  INV_X1 U4514 ( .A(n3734), .ZN(n3735) );
  OR2_X1 U4515 ( .A1(n3736), .A2(n3735), .ZN(n3737) );
  OR2_X1 U4516 ( .A1(n3798), .A2(n3743), .ZN(n3740) );
  NAND2_X1 U4517 ( .A1(n4078), .A2(n3741), .ZN(n3739) );
  NAND2_X1 U4518 ( .A1(n3740), .A2(n3739), .ZN(n3747) );
  NAND2_X1 U4519 ( .A1(n4079), .A2(n3741), .ZN(n3742) );
  OAI21_X1 U4520 ( .B1(n3743), .B2(n3652), .A(n3742), .ZN(n3744) );
  XNOR2_X1 U4521 ( .A(n3744), .B(n4043), .ZN(n3746) );
  XNOR2_X1 U4522 ( .A(n3747), .B(n3746), .ZN(n3789) );
  NAND2_X1 U4523 ( .A1(n3747), .A2(n3746), .ZN(n3748) );
  NAND2_X1 U4524 ( .A1(n3756), .A2(n4079), .ZN(n3749) );
  OAI21_X1 U4525 ( .B1(n3751), .B2(n3652), .A(n3749), .ZN(n3750) );
  XNOR2_X1 U4526 ( .A(n3750), .B(n4043), .ZN(n3794) );
  OR2_X1 U4527 ( .A1(n3798), .A2(n3751), .ZN(n3753) );
  NAND2_X1 U4528 ( .A1(n4078), .A2(n3756), .ZN(n3752) );
  NAND2_X1 U4529 ( .A1(n3753), .A2(n3752), .ZN(n3795) );
  XOR2_X1 U4530 ( .A(n3794), .B(n3795), .Z(n3754) );
  XNOR2_X1 U4531 ( .A(n3796), .B(n3754), .ZN(n3762) );
  NAND2_X1 U4532 ( .A1(n4287), .A2(n4305), .ZN(n3758) );
  AOI21_X1 U4533 ( .B1(n4288), .B2(n3756), .A(n3755), .ZN(n3757) );
  OAI211_X1 U4534 ( .C1(n3797), .C2(n4291), .A(n3758), .B(n3757), .ZN(n3759)
         );
  AOI21_X1 U4535 ( .B1(n4294), .B2(n3760), .A(n3759), .ZN(n3761) );
  OAI21_X1 U4536 ( .B1(n3762), .B2(n4296), .A(n3761), .ZN(U3233) );
  XNOR2_X1 U4537 ( .A(n3763), .B(REG1_REG_12__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4538 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3809) );
  XOR2_X1 U4539 ( .A(REG2_REG_12__SCAN_IN), .B(n3764), .Z(n3765) );
  NAND2_X1 U4540 ( .A1(n4342), .A2(n3765), .ZN(n3766) );
  NAND2_X1 U4541 ( .A1(n3809), .A2(n3766), .ZN(n3769) );
  NOR2_X1 U4542 ( .A1(n4852), .A2(n3767), .ZN(n3768) );
  AOI211_X1 U4543 ( .C1(n4846), .C2(ADDR_REG_12__SCAN_IN), .A(n3769), .B(n3768), .ZN(n3770) );
  OAI21_X1 U4544 ( .B1(n3771), .B2(n4360), .A(n3770), .ZN(U3252) );
  NAND2_X1 U4545 ( .A1(n3772), .A2(n3815), .ZN(n3773) );
  XNOR2_X1 U4546 ( .A(n3773), .B(n3909), .ZN(n3774) );
  NOR2_X1 U4547 ( .A1(n3774), .A2(n4631), .ZN(n4719) );
  INV_X1 U4548 ( .A(n4719), .ZN(n3783) );
  XNOR2_X1 U4549 ( .A(n3775), .B(n3909), .ZN(n4721) );
  OAI21_X1 U4550 ( .B1(n3700), .B2(n3779), .A(n4638), .ZN(n4795) );
  NOR2_X1 U4551 ( .A1(n4795), .A2(n4642), .ZN(n3781) );
  AOI22_X1 U4552 ( .A1(n4612), .A2(n4716), .B1(n4613), .B2(n4611), .ZN(n3778)
         );
  INV_X1 U4553 ( .A(n3776), .ZN(n4293) );
  AOI22_X1 U4554 ( .A1(n4646), .A2(REG2_REG_15__SCAN_IN), .B1(n4293), .B2(
        n4859), .ZN(n3777) );
  OAI211_X1 U4555 ( .C1(n3779), .C2(n4617), .A(n3778), .B(n3777), .ZN(n3780)
         );
  AOI211_X1 U4556 ( .C1(n4721), .C2(n4644), .A(n3781), .B(n3780), .ZN(n3782)
         );
  OAI21_X1 U4557 ( .B1(n3783), .B2(n4624), .A(n3782), .ZN(U3275) );
  AOI22_X1 U4558 ( .A1(n4287), .A2(n4306), .B1(n4262), .B2(n4739), .ZN(n3785)
         );
  OAI211_X1 U4559 ( .C1(n4241), .C2(n2184), .A(n3785), .B(n3784), .ZN(n3791)
         );
  INV_X1 U4560 ( .A(n3787), .ZN(n3788) );
  AOI211_X1 U4561 ( .C1(n3789), .C2(n3786), .A(n4296), .B(n3788), .ZN(n3790)
         );
  AOI211_X1 U4562 ( .C1(n3792), .C2(n4294), .A(n3791), .B(n3790), .ZN(n3793)
         );
  INV_X1 U4563 ( .A(n3793), .ZN(U3214) );
  OR2_X1 U4564 ( .A1(n3798), .A2(n3797), .ZN(n3800) );
  NAND2_X1 U4565 ( .A1(n3801), .A2(n4078), .ZN(n3799) );
  NAND2_X1 U4566 ( .A1(n3800), .A2(n3799), .ZN(n3805) );
  NAND2_X1 U4567 ( .A1(n3801), .A2(n4079), .ZN(n3803) );
  NAND2_X1 U4568 ( .A1(n4078), .A2(n4304), .ZN(n3802) );
  NAND2_X1 U4569 ( .A1(n3803), .A2(n3802), .ZN(n3804) );
  XNOR2_X1 U4570 ( .A(n3804), .B(n4043), .ZN(n3806) );
  INV_X1 U4571 ( .A(n3977), .ZN(n3807) );
  NOR2_X1 U4572 ( .A1(n3807), .A2(n3978), .ZN(n3808) );
  XNOR2_X1 U4573 ( .A(n3979), .B(n3808), .ZN(n3814) );
  AOI22_X1 U4574 ( .A1(n4287), .A2(n4739), .B1(n4262), .B2(n4736), .ZN(n3810)
         );
  OAI211_X1 U4575 ( .C1(n4241), .C2(n2893), .A(n3810), .B(n3809), .ZN(n3811)
         );
  AOI21_X1 U4576 ( .B1(n3812), .B2(n4294), .A(n3811), .ZN(n3813) );
  OAI21_X1 U4577 ( .B1(n3814), .B2(n4296), .A(n3813), .ZN(U3221) );
  AND2_X1 U4578 ( .A1(n3816), .A2(n3815), .ZN(n3861) );
  NAND2_X1 U4579 ( .A1(n3818), .A2(n3817), .ZN(n3934) );
  INV_X1 U4580 ( .A(n3819), .ZN(n3822) );
  OAI211_X1 U4581 ( .C1(n3822), .C2(n2862), .A(n3821), .B(n3820), .ZN(n3825)
         );
  NAND3_X1 U4582 ( .A1(n3825), .A2(n3824), .A3(n3823), .ZN(n3828) );
  NAND3_X1 U4583 ( .A1(n3828), .A2(n3827), .A3(n3826), .ZN(n3831) );
  NAND3_X1 U4584 ( .A1(n3831), .A2(n3830), .A3(n3829), .ZN(n3838) );
  INV_X1 U4585 ( .A(n3845), .ZN(n3834) );
  NOR3_X1 U4586 ( .A1(n3834), .A2(n2216), .A3(n3833), .ZN(n3837) );
  INV_X1 U4587 ( .A(n3835), .ZN(n3836) );
  AOI211_X1 U4588 ( .C1(n3838), .C2(n3837), .A(n3836), .B(n3890), .ZN(n3843)
         );
  NAND2_X1 U4589 ( .A1(n3840), .A2(n3839), .ZN(n3847) );
  OAI211_X1 U4590 ( .C1(n3843), .C2(n3847), .A(n3842), .B(n3841), .ZN(n3859)
         );
  INV_X1 U4591 ( .A(n3844), .ZN(n3846) );
  NAND2_X1 U4592 ( .A1(n3846), .A2(n3845), .ZN(n3848) );
  OAI21_X1 U4593 ( .B1(n3848), .B2(n3847), .A(n3849), .ZN(n3858) );
  INV_X1 U4594 ( .A(n3934), .ZN(n3857) );
  INV_X1 U4595 ( .A(n3849), .ZN(n3853) );
  OAI211_X1 U4596 ( .C1(n3853), .C2(n3852), .A(n3851), .B(n3850), .ZN(n3855)
         );
  NOR2_X1 U4597 ( .A1(n3855), .A2(n3854), .ZN(n3856) );
  OAI211_X1 U4598 ( .C1(n3859), .C2(n3858), .A(n3857), .B(n3856), .ZN(n3860)
         );
  OAI211_X1 U4599 ( .C1(n3861), .C2(n3934), .A(n3860), .B(n3932), .ZN(n3862)
         );
  NAND2_X1 U4600 ( .A1(n3862), .A2(n3938), .ZN(n3863) );
  AOI211_X1 U4601 ( .C1(n3863), .C2(n3933), .A(n3895), .B(n3936), .ZN(n3865)
         );
  INV_X1 U4602 ( .A(n3942), .ZN(n3864) );
  INV_X1 U4603 ( .A(n4486), .ZN(n3889) );
  OAI211_X1 U4604 ( .C1(n3865), .C2(n3864), .A(n3940), .B(n3889), .ZN(n3867)
         );
  AOI21_X1 U4605 ( .B1(n3867), .B2(n3944), .A(n3866), .ZN(n3870) );
  INV_X1 U4606 ( .A(n3948), .ZN(n3869) );
  NAND2_X1 U4607 ( .A1(n2748), .A2(n3887), .ZN(n3947) );
  INV_X1 U4608 ( .A(n3947), .ZN(n3868) );
  OAI21_X1 U4609 ( .B1(n3870), .B2(n3869), .A(n3868), .ZN(n3871) );
  NAND2_X1 U4610 ( .A1(n3871), .A2(n3952), .ZN(n3875) );
  NAND2_X1 U4611 ( .A1(n4300), .A2(n4394), .ZN(n3872) );
  NAND2_X1 U4612 ( .A1(n3873), .A2(n3872), .ZN(n3957) );
  INV_X1 U4613 ( .A(n3957), .ZN(n3877) );
  NAND4_X1 U4614 ( .A1(n3875), .A2(n3877), .A3(n3954), .A4(n3874), .ZN(n3885)
         );
  NAND2_X1 U4615 ( .A1(n3953), .A2(n3950), .ZN(n3876) );
  NAND2_X1 U4616 ( .A1(n3877), .A2(n3876), .ZN(n3880) );
  INV_X1 U4617 ( .A(n4386), .ZN(n3881) );
  OR2_X1 U4618 ( .A1(n4299), .A2(n3881), .ZN(n3878) );
  NAND2_X1 U4619 ( .A1(n4298), .A2(n4382), .ZN(n3883) );
  NAND2_X1 U4620 ( .A1(n3878), .A2(n3883), .ZN(n3897) );
  AOI21_X1 U4621 ( .B1(n4409), .B2(n3879), .A(n3897), .ZN(n3951) );
  INV_X1 U4622 ( .A(n3958), .ZN(n3884) );
  NAND2_X1 U4623 ( .A1(n3881), .A2(n4299), .ZN(n3963) );
  OR2_X1 U4624 ( .A1(n4298), .A2(n4382), .ZN(n3882) );
  NAND2_X1 U4625 ( .A1(n3963), .A2(n3882), .ZN(n3896) );
  AOI22_X1 U4626 ( .A1(n3885), .A2(n3884), .B1(n3883), .B2(n3896), .ZN(n3969)
         );
  NAND2_X1 U4627 ( .A1(n2354), .A2(n3886), .ZN(n4436) );
  XNOR2_X1 U4628 ( .A(n4665), .B(n4495), .ZN(n4491) );
  NAND2_X1 U4629 ( .A1(n3888), .A2(n3887), .ZN(n4469) );
  AND2_X1 U4630 ( .A1(n3889), .A2(n4487), .ZN(n4529) );
  INV_X1 U4631 ( .A(n3161), .ZN(n3893) );
  NOR2_X1 U4632 ( .A1(n3891), .A2(n3890), .ZN(n3892) );
  NAND4_X1 U4633 ( .A1(n4588), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3904)
         );
  INV_X1 U4634 ( .A(n3895), .ZN(n3937) );
  AND2_X1 U4635 ( .A1(n3937), .A2(n4567), .ZN(n4610) );
  NOR2_X1 U4636 ( .A1(n3897), .A2(n3896), .ZN(n3901) );
  NOR2_X1 U4637 ( .A1(n3899), .A2(n3898), .ZN(n3900) );
  NAND4_X1 U4638 ( .A1(n4610), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3903)
         );
  NOR2_X1 U4639 ( .A1(n3904), .A2(n3903), .ZN(n3907) );
  NAND2_X1 U4640 ( .A1(n3906), .A2(n3905), .ZN(n4547) );
  AND2_X1 U4641 ( .A1(n3907), .A2(n4547), .ZN(n3921) );
  XNOR2_X1 U4642 ( .A(n4593), .B(n4579), .ZN(n4577) );
  NOR3_X1 U4643 ( .A1(n3909), .A2(n3908), .A3(n4884), .ZN(n3918) );
  NOR2_X1 U4644 ( .A1(n3911), .A2(n3910), .ZN(n3915) );
  AND4_X1 U4645 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(n3917)
         );
  NAND4_X1 U4646 ( .A1(n3918), .A2(n3917), .A3(n4637), .A4(n3916), .ZN(n3919)
         );
  NOR2_X1 U4647 ( .A1(n4577), .A2(n3919), .ZN(n3920) );
  NAND4_X1 U4648 ( .A1(n4513), .A2(n4529), .A3(n3921), .A4(n3920), .ZN(n3922)
         );
  NOR2_X1 U4649 ( .A1(n4469), .A2(n3922), .ZN(n3923) );
  NAND3_X1 U4650 ( .A1(n4436), .A2(n4491), .A3(n3923), .ZN(n3924) );
  NOR2_X1 U4651 ( .A1(n3924), .A2(n3956), .ZN(n3928) );
  INV_X1 U4652 ( .A(n4433), .ZN(n3926) );
  INV_X1 U4653 ( .A(n4454), .ZN(n3927) );
  NOR2_X1 U4654 ( .A1(n3931), .A2(n3930), .ZN(n3935) );
  OAI211_X1 U4655 ( .C1(n3935), .C2(n3934), .A(n3933), .B(n3932), .ZN(n3939)
         );
  NAND4_X1 U4656 ( .A1(n3939), .A2(n2686), .A3(n3938), .A4(n3937), .ZN(n3943)
         );
  INV_X1 U4657 ( .A(n3940), .ZN(n3941) );
  AOI21_X1 U4658 ( .B1(n3943), .B2(n3942), .A(n3941), .ZN(n3946) );
  OAI21_X1 U4659 ( .B1(n3946), .B2(n2197), .A(n3945), .ZN(n3949) );
  AOI21_X1 U4660 ( .B1(n3949), .B2(n3948), .A(n3947), .ZN(n3961) );
  NAND4_X1 U4661 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3960)
         );
  INV_X1 U4662 ( .A(n3954), .ZN(n3955) );
  NOR3_X1 U4663 ( .A1(n3957), .A2(n3956), .A3(n3955), .ZN(n3959) );
  INV_X1 U4664 ( .A(n4298), .ZN(n3962) );
  NAND2_X1 U4665 ( .A1(n3962), .A2(n4386), .ZN(n3965) );
  AOI21_X1 U4666 ( .B1(n3963), .B2(n4298), .A(n4382), .ZN(n3964) );
  AOI21_X1 U4667 ( .B1(n3966), .B2(n3965), .A(n3964), .ZN(n3967) );
  MUX2_X1 U4668 ( .A(n2353), .B(n3967), .S(n2862), .Z(n3968) );
  XNOR2_X1 U4669 ( .A(n3970), .B(n3181), .ZN(n3976) );
  NOR2_X1 U4670 ( .A1(n3972), .A2(n3971), .ZN(n3974) );
  OAI21_X1 U4671 ( .B1(n3975), .B2(n2807), .A(B_REG_SCAN_IN), .ZN(n3973) );
  OAI22_X1 U4672 ( .A1(n3976), .A2(n3975), .B1(n3974), .B2(n3973), .ZN(U3239)
         );
  NAND2_X1 U4673 ( .A1(n4078), .A2(n4736), .ZN(n3981) );
  NAND2_X1 U4674 ( .A1(n4079), .A2(n4228), .ZN(n3980) );
  NAND2_X1 U4675 ( .A1(n3981), .A2(n3980), .ZN(n3982) );
  XNOR2_X1 U4676 ( .A(n3982), .B(n4087), .ZN(n4226) );
  NAND2_X1 U4677 ( .A1(n4224), .A2(n4226), .ZN(n3986) );
  INV_X1 U4678 ( .A(n4736), .ZN(n3983) );
  OR2_X1 U4679 ( .A1(n3798), .A2(n3983), .ZN(n3985) );
  NAND2_X1 U4680 ( .A1(n4078), .A2(n4228), .ZN(n3984) );
  NAND2_X1 U4681 ( .A1(n3985), .A2(n3984), .ZN(n4225) );
  NAND2_X1 U4682 ( .A1(n3986), .A2(n4225), .ZN(n3990) );
  INV_X1 U4683 ( .A(n4224), .ZN(n3988) );
  INV_X1 U4684 ( .A(n4226), .ZN(n3987) );
  NAND2_X1 U4685 ( .A1(n3988), .A2(n3987), .ZN(n3989) );
  OAI22_X1 U4686 ( .A1(n4231), .A2(n3652), .B1(n4089), .B2(n3991), .ZN(n3992)
         );
  XNOR2_X1 U4687 ( .A(n3992), .B(n4043), .ZN(n4003) );
  OR2_X1 U4688 ( .A1(n3798), .A2(n4231), .ZN(n3994) );
  NAND2_X1 U4689 ( .A1(n4078), .A2(n4723), .ZN(n3993) );
  NAND2_X1 U4690 ( .A1(n3994), .A2(n3993), .ZN(n4004) );
  INV_X1 U4691 ( .A(n4303), .ZN(n4727) );
  OR2_X1 U4692 ( .A1(n4727), .A2(n3798), .ZN(n3996) );
  NAND2_X1 U4693 ( .A1(n4078), .A2(n4715), .ZN(n3995) );
  NAND2_X1 U4694 ( .A1(n3996), .A2(n3995), .ZN(n4184) );
  NAND2_X1 U4695 ( .A1(n4303), .A2(n4078), .ZN(n3998) );
  NAND2_X1 U4696 ( .A1(n4079), .A2(n4715), .ZN(n3997) );
  NAND2_X1 U4697 ( .A1(n3998), .A2(n3997), .ZN(n3999) );
  XNOR2_X1 U4698 ( .A(n3999), .B(n4043), .ZN(n4187) );
  OAI22_X1 U4699 ( .A1(n4718), .A2(n3652), .B1(n4089), .B2(n4639), .ZN(n4000)
         );
  XNOR2_X1 U4700 ( .A(n4000), .B(n4043), .ZN(n4009) );
  INV_X1 U4701 ( .A(n4009), .ZN(n4002) );
  OAI22_X1 U4702 ( .A1(n4718), .A2(n3798), .B1(n3652), .B2(n4639), .ZN(n4008)
         );
  INV_X1 U4703 ( .A(n4008), .ZN(n4001) );
  NAND2_X1 U4704 ( .A1(n4002), .A2(n4001), .ZN(n4007) );
  INV_X1 U4705 ( .A(n4003), .ZN(n4006) );
  INV_X1 U4706 ( .A(n4004), .ZN(n4005) );
  NAND2_X1 U4707 ( .A1(n4006), .A2(n4005), .ZN(n4116) );
  OAI211_X1 U4708 ( .C1(n4184), .C2(n4187), .A(n4007), .B(n4116), .ZN(n4011)
         );
  INV_X1 U4709 ( .A(n4007), .ZN(n4190) );
  AND2_X1 U4710 ( .A1(n4009), .A2(n4008), .ZN(n4189) );
  AOI21_X1 U4711 ( .B1(n4184), .B2(n4187), .A(n4189), .ZN(n4010) );
  OAI22_X1 U4712 ( .A1(n4627), .A2(n3652), .B1(n4089), .B2(n4620), .ZN(n4012)
         );
  XNOR2_X1 U4713 ( .A(n4012), .B(n4043), .ZN(n4014) );
  OAI22_X1 U4714 ( .A1(n4627), .A2(n3798), .B1(n3652), .B2(n4620), .ZN(n4013)
         );
  AND2_X1 U4715 ( .A1(n4014), .A2(n4013), .ZN(n4198) );
  OR2_X1 U4716 ( .A1(n4014), .A2(n4013), .ZN(n4197) );
  NAND2_X1 U4717 ( .A1(n4593), .A2(n4078), .ZN(n4016) );
  NAND2_X1 U4718 ( .A1(n4143), .A2(n4079), .ZN(n4015) );
  NAND2_X1 U4719 ( .A1(n4016), .A2(n4015), .ZN(n4017) );
  XNOR2_X1 U4720 ( .A(n4017), .B(n4043), .ZN(n4024) );
  NAND2_X1 U4721 ( .A1(n4593), .A2(n4018), .ZN(n4020) );
  NAND2_X1 U4722 ( .A1(n4078), .A2(n4143), .ZN(n4019) );
  NAND2_X1 U4723 ( .A1(n4020), .A2(n4019), .ZN(n4025) );
  NAND2_X1 U4724 ( .A1(n4024), .A2(n4025), .ZN(n4139) );
  OAI22_X1 U4725 ( .A1(n4572), .A2(n3652), .B1(n4089), .B2(n4598), .ZN(n4021)
         );
  XNOR2_X1 U4726 ( .A(n4021), .B(n4087), .ZN(n4259) );
  NOR2_X1 U4727 ( .A1(n4598), .A2(n3652), .ZN(n4022) );
  AOI21_X1 U4728 ( .B1(n4705), .B2(n3266), .A(n4022), .ZN(n4258) );
  INV_X1 U4729 ( .A(n4139), .ZN(n4029) );
  NAND2_X1 U4730 ( .A1(n4259), .A2(n4258), .ZN(n4028) );
  INV_X1 U4731 ( .A(n4024), .ZN(n4027) );
  INV_X1 U4732 ( .A(n4025), .ZN(n4026) );
  NAND2_X1 U4733 ( .A1(n4027), .A2(n4026), .ZN(n4138) );
  NAND2_X1 U4734 ( .A1(n4683), .A2(n4078), .ZN(n4033) );
  NAND2_X1 U4735 ( .A1(n4079), .A2(n4549), .ZN(n4032) );
  NAND2_X1 U4736 ( .A1(n4033), .A2(n4032), .ZN(n4034) );
  XNOR2_X1 U4737 ( .A(n4034), .B(n4043), .ZN(n4037) );
  NAND2_X1 U4738 ( .A1(n4683), .A2(n4018), .ZN(n4036) );
  NAND2_X1 U4739 ( .A1(n4078), .A2(n4549), .ZN(n4035) );
  NAND2_X1 U4740 ( .A1(n4036), .A2(n4035), .ZN(n4038) );
  NAND2_X1 U4741 ( .A1(n4037), .A2(n4038), .ZN(n4216) );
  INV_X1 U4742 ( .A(n4037), .ZN(n4040) );
  INV_X1 U4743 ( .A(n4038), .ZN(n4039) );
  NAND2_X1 U4744 ( .A1(n4040), .A2(n4039), .ZN(n4161) );
  NAND2_X1 U4745 ( .A1(n4507), .A2(n4078), .ZN(n4042) );
  NAND2_X1 U4746 ( .A1(n4079), .A2(n4682), .ZN(n4041) );
  NAND2_X1 U4747 ( .A1(n4042), .A2(n4041), .ZN(n4044) );
  XNOR2_X1 U4748 ( .A(n4044), .B(n4043), .ZN(n4048) );
  NAND2_X1 U4749 ( .A1(n4507), .A2(n4018), .ZN(n4046) );
  NAND2_X1 U4750 ( .A1(n4078), .A2(n4682), .ZN(n4045) );
  NAND2_X1 U4751 ( .A1(n4046), .A2(n4045), .ZN(n4047) );
  NOR2_X1 U4752 ( .A1(n4048), .A2(n4047), .ZN(n4157) );
  NAND2_X1 U4753 ( .A1(n4048), .A2(n4047), .ZN(n4158) );
  OAI22_X1 U4754 ( .A1(n4686), .A2(n3652), .B1(n4089), .B2(n2896), .ZN(n4049)
         );
  XNOR2_X1 U4755 ( .A(n4049), .B(n4043), .ZN(n4055) );
  OAI22_X1 U4756 ( .A1(n4686), .A2(n3798), .B1(n3652), .B2(n2896), .ZN(n4054)
         );
  XNOR2_X1 U4757 ( .A(n4055), .B(n4054), .ZN(n4238) );
  NAND2_X1 U4758 ( .A1(n4665), .A2(n4078), .ZN(n4051) );
  NAND2_X1 U4759 ( .A1(n4079), .A2(n4495), .ZN(n4050) );
  NAND2_X1 U4760 ( .A1(n4051), .A2(n4050), .ZN(n4052) );
  XNOR2_X1 U4761 ( .A(n4052), .B(n4087), .ZN(n4064) );
  NOR2_X1 U4762 ( .A1(n3652), .A2(n4499), .ZN(n4053) );
  AOI21_X1 U4763 ( .B1(n4665), .B2(n4018), .A(n4053), .ZN(n4065) );
  XNOR2_X1 U4764 ( .A(n4064), .B(n4065), .ZN(n4126) );
  NOR2_X1 U4765 ( .A1(n4055), .A2(n4054), .ZN(n4127) );
  NAND2_X1 U4766 ( .A1(n4473), .A2(n4078), .ZN(n4059) );
  NAND2_X1 U4767 ( .A1(n4079), .A2(n4655), .ZN(n4058) );
  NAND2_X1 U4768 ( .A1(n4059), .A2(n4058), .ZN(n4060) );
  XNOR2_X1 U4769 ( .A(n4060), .B(n4087), .ZN(n4179) );
  AOI22_X1 U4770 ( .A1(n4473), .A2(n4018), .B1(n4078), .B2(n4655), .ZN(n4178)
         );
  NOR2_X1 U4771 ( .A1(n4179), .A2(n4178), .ZN(n4177) );
  INV_X1 U4772 ( .A(n4177), .ZN(n4071) );
  NAND2_X1 U4773 ( .A1(n4656), .A2(n4078), .ZN(n4062) );
  NAND2_X1 U4774 ( .A1(n4079), .A2(n4664), .ZN(n4061) );
  NAND2_X1 U4775 ( .A1(n4062), .A2(n4061), .ZN(n4063) );
  INV_X1 U4776 ( .A(n4064), .ZN(n4067) );
  INV_X1 U4777 ( .A(n4065), .ZN(n4066) );
  NAND2_X1 U4778 ( .A1(n4067), .A2(n4066), .ZN(n4172) );
  NAND2_X1 U4779 ( .A1(n4209), .A2(n4172), .ZN(n4069) );
  NOR2_X1 U4780 ( .A1(n3652), .A2(n4474), .ZN(n4068) );
  AOI21_X1 U4781 ( .B1(n4656), .B2(n4018), .A(n4068), .ZN(n4173) );
  NAND2_X1 U4782 ( .A1(n4172), .A2(n4173), .ZN(n4171) );
  NAND2_X1 U4783 ( .A1(n4069), .A2(n4171), .ZN(n4070) );
  AOI21_X1 U4784 ( .B1(n4209), .B2(n4173), .A(n4178), .ZN(n4075) );
  INV_X1 U4785 ( .A(n4179), .ZN(n4074) );
  INV_X1 U4786 ( .A(n4209), .ZN(n4073) );
  NAND2_X1 U4787 ( .A1(n4178), .A2(n4173), .ZN(n4072) );
  OAI22_X1 U4788 ( .A1(n4075), .A2(n4074), .B1(n4073), .B2(n4072), .ZN(n4076)
         );
  NAND2_X1 U4789 ( .A1(n4424), .A2(n4078), .ZN(n4081) );
  NAND2_X1 U4790 ( .A1(n4079), .A2(n4442), .ZN(n4080) );
  NAND2_X1 U4791 ( .A1(n4081), .A2(n4080), .ZN(n4082) );
  XNOR2_X1 U4792 ( .A(n4082), .B(n4087), .ZN(n4085) );
  NOR2_X1 U4793 ( .A1(n3652), .A2(n4437), .ZN(n4083) );
  AOI21_X1 U4794 ( .B1(n4424), .B2(n4018), .A(n4083), .ZN(n4084) );
  NOR2_X1 U4795 ( .A1(n4085), .A2(n4084), .ZN(n4273) );
  NAND2_X1 U4796 ( .A1(n4085), .A2(n4084), .ZN(n4271) );
  OAI22_X1 U4797 ( .A1(n4438), .A2(n3652), .B1(n4419), .B2(n4089), .ZN(n4086)
         );
  XNOR2_X1 U4798 ( .A(n4086), .B(n4043), .ZN(n4094) );
  OAI22_X1 U4799 ( .A1(n4438), .A2(n3798), .B1(n4419), .B2(n3383), .ZN(n4093)
         );
  XNOR2_X1 U4800 ( .A(n4094), .B(n4093), .ZN(n4107) );
  OAI22_X1 U4801 ( .A1(n4426), .A2(n3798), .B1(n3652), .B2(n4406), .ZN(n4088)
         );
  XNOR2_X1 U4802 ( .A(n4088), .B(n4087), .ZN(n4091) );
  OAI22_X1 U4803 ( .A1(n4426), .A2(n3383), .B1(n4089), .B2(n4406), .ZN(n4090)
         );
  XNOR2_X1 U4804 ( .A(n4091), .B(n4090), .ZN(n4099) );
  INV_X1 U4805 ( .A(n4099), .ZN(n4092) );
  NAND2_X1 U4806 ( .A1(n4092), .A2(n4250), .ZN(n4105) );
  NAND2_X1 U4807 ( .A1(n4094), .A2(n4093), .ZN(n4098) );
  INV_X1 U4808 ( .A(n4408), .ZN(n4102) );
  AOI22_X1 U4809 ( .A1(n4288), .A2(n4095), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n4097) );
  NAND2_X1 U4810 ( .A1(n4300), .A2(n4262), .ZN(n4096) );
  OAI211_X1 U4811 ( .C1(n4438), .C2(n4267), .A(n4097), .B(n4096), .ZN(n4101)
         );
  NOR3_X1 U4812 ( .A1(n4099), .A2(n4296), .A3(n4098), .ZN(n4100) );
  AOI211_X1 U4813 ( .C1(n4102), .C2(n4294), .A(n4101), .B(n4100), .ZN(n4103)
         );
  OAI211_X1 U4814 ( .C1(n4106), .C2(n4105), .A(n4104), .B(n4103), .ZN(U3217)
         );
  XNOR2_X1 U4815 ( .A(n4108), .B(n4107), .ZN(n4114) );
  NOR2_X1 U4816 ( .A1(n4421), .A2(n4276), .ZN(n4112) );
  AOI22_X1 U4817 ( .A1(n4288), .A2(n4109), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n4110) );
  OAI21_X1 U4818 ( .B1(n4659), .B2(n4267), .A(n4110), .ZN(n4111) );
  AOI211_X1 U4819 ( .C1(n4396), .C2(n4262), .A(n4112), .B(n4111), .ZN(n4113)
         );
  OAI21_X1 U4820 ( .B1(n4114), .B2(n4296), .A(n4113), .ZN(U3211) );
  INV_X1 U4821 ( .A(n4116), .ZN(n4186) );
  NOR2_X1 U4822 ( .A1(n4186), .A2(n4117), .ZN(n4118) );
  XNOR2_X1 U4823 ( .A(n4115), .B(n4118), .ZN(n4124) );
  NAND2_X1 U4824 ( .A1(n4287), .A2(n4736), .ZN(n4120) );
  AND2_X1 U4825 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4341) );
  AOI21_X1 U4826 ( .B1(n4288), .B2(n4723), .A(n4341), .ZN(n4119) );
  OAI211_X1 U4827 ( .C1(n4727), .C2(n4291), .A(n4120), .B(n4119), .ZN(n4121)
         );
  AOI21_X1 U4828 ( .B1(n4294), .B2(n4122), .A(n4121), .ZN(n4123) );
  OAI21_X1 U4829 ( .B1(n4124), .B2(n4296), .A(n4123), .ZN(U3212) );
  OAI21_X1 U4830 ( .B1(n4236), .B2(n4127), .A(n4126), .ZN(n4128) );
  NAND3_X1 U4831 ( .A1(n4077), .A2(n4250), .A3(n4128), .ZN(n4133) );
  OAI22_X1 U4832 ( .A1(n4241), .A2(n4499), .B1(STATE_REG_SCAN_IN), .B2(n4129), 
        .ZN(n4131) );
  OAI22_X1 U4833 ( .A1(n2331), .A2(n4291), .B1(n4686), .B2(n4267), .ZN(n4130)
         );
  AOI211_X1 U4834 ( .C1(n4501), .C2(n4294), .A(n4131), .B(n4130), .ZN(n4132)
         );
  NAND2_X1 U4835 ( .A1(n4133), .A2(n4132), .ZN(U3213) );
  INV_X1 U4836 ( .A(n4134), .ZN(n4137) );
  INV_X1 U4837 ( .A(n4258), .ZN(n4136) );
  AOI21_X1 U4838 ( .B1(n4134), .B2(n4258), .A(n4259), .ZN(n4135) );
  AOI21_X1 U4839 ( .B1(n4137), .B2(n4136), .A(n4135), .ZN(n4141) );
  NAND2_X1 U4840 ( .A1(n4139), .A2(n4138), .ZN(n4140) );
  XNOR2_X1 U4841 ( .A(n4141), .B(n4140), .ZN(n4148) );
  NAND2_X1 U4842 ( .A1(n4287), .A2(n4705), .ZN(n4145) );
  NAND2_X1 U4843 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4372) );
  INV_X1 U4844 ( .A(n4372), .ZN(n4142) );
  AOI21_X1 U4845 ( .B1(n4288), .B2(n4143), .A(n4142), .ZN(n4144) );
  OAI211_X1 U4846 ( .C1(n4536), .C2(n4291), .A(n4145), .B(n4144), .ZN(n4146)
         );
  AOI21_X1 U4847 ( .B1(n4294), .B2(n4580), .A(n4146), .ZN(n4147) );
  OAI21_X1 U4848 ( .B1(n4148), .B2(n4296), .A(n4147), .ZN(U3216) );
  AOI22_X1 U4849 ( .A1(n4254), .A2(REG3_REG_1__SCAN_IN), .B1(n4262), .B2(n4313), .ZN(n4156) );
  AOI22_X1 U4850 ( .A1(n4287), .A2(n4149), .B1(n3261), .B2(n4288), .ZN(n4155)
         );
  NAND2_X1 U4851 ( .A1(n4151), .A2(n4153), .ZN(n4152) );
  OAI211_X1 U4852 ( .C1(n4153), .C2(n4151), .A(n4250), .B(n4152), .ZN(n4154)
         );
  NAND3_X1 U4853 ( .A1(n4156), .A2(n4155), .A3(n4154), .ZN(U3219) );
  INV_X1 U4854 ( .A(n4532), .ZN(n4170) );
  INV_X1 U4855 ( .A(n4157), .ZN(n4159) );
  NAND2_X1 U4856 ( .A1(n4159), .A2(n4158), .ZN(n4163) );
  OAI211_X1 U4857 ( .C1(n4160), .C2(n2288), .A(n4216), .B(n4163), .ZN(n4162)
         );
  OAI211_X1 U4858 ( .C1(n4164), .C2(n4163), .A(n4250), .B(n4162), .ZN(n4169)
         );
  AOI22_X1 U4859 ( .A1(n4288), .A2(n4682), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n4166) );
  NAND2_X1 U4860 ( .A1(n4287), .A2(n4683), .ZN(n4165) );
  OAI211_X1 U4861 ( .C1(n4686), .C2(n4291), .A(n4166), .B(n4165), .ZN(n4167)
         );
  INV_X1 U4862 ( .A(n4167), .ZN(n4168) );
  OAI211_X1 U4863 ( .C1(n4276), .C2(n4170), .A(n4169), .B(n4168), .ZN(U3220)
         );
  INV_X1 U4864 ( .A(n4172), .ZN(n4175) );
  INV_X1 U4865 ( .A(n4173), .ZN(n4174) );
  AOI21_X1 U4866 ( .B1(n4179), .B2(n4178), .A(n4177), .ZN(n4180) );
  OAI22_X1 U4867 ( .A1(n4241), .A2(n4456), .B1(STATE_REG_SCAN_IN), .B2(n3003), 
        .ZN(n4182) );
  OAI22_X1 U4868 ( .A1(n4659), .A2(n4291), .B1(n2331), .B2(n4267), .ZN(n4181)
         );
  AOI211_X1 U4869 ( .C1(n4457), .C2(n4294), .A(n4182), .B(n4181), .ZN(n4183)
         );
  INV_X1 U4870 ( .A(n4184), .ZN(n4285) );
  NOR2_X1 U4871 ( .A1(n4185), .A2(n4186), .ZN(n4188) );
  NAND2_X1 U4872 ( .A1(n4188), .A2(n4187), .ZN(n4283) );
  NOR2_X1 U4873 ( .A1(n4188), .A2(n4187), .ZN(n4282) );
  AOI21_X1 U4874 ( .B1(n4285), .B2(n4283), .A(n4282), .ZN(n4192) );
  NOR2_X1 U4875 ( .A1(n4190), .A2(n4189), .ZN(n4191) );
  XNOR2_X1 U4876 ( .A(n4192), .B(n4191), .ZN(n4196) );
  AOI22_X1 U4877 ( .A1(n4287), .A2(n4303), .B1(n4262), .B2(n4302), .ZN(n4193)
         );
  NAND2_X1 U4878 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4839) );
  OAI211_X1 U4879 ( .C1(n4241), .C2(n4639), .A(n4193), .B(n4839), .ZN(n4194)
         );
  AOI21_X1 U4880 ( .B1(n4640), .B2(n4294), .A(n4194), .ZN(n4195) );
  OAI21_X1 U4881 ( .B1(n4196), .B2(n4296), .A(n4195), .ZN(U3223) );
  INV_X1 U4882 ( .A(n4197), .ZN(n4199) );
  NOR2_X1 U4883 ( .A1(n4199), .A2(n4198), .ZN(n4200) );
  XNOR2_X1 U4884 ( .A(n4201), .B(n4200), .ZN(n4207) );
  INV_X1 U4885 ( .A(n4202), .ZN(n4614) );
  NAND2_X1 U4886 ( .A1(n4262), .A2(n4705), .ZN(n4204) );
  AND2_X1 U4887 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4355) );
  AOI21_X1 U4888 ( .B1(n4288), .B2(n4704), .A(n4355), .ZN(n4203) );
  OAI211_X1 U4889 ( .C1(n4718), .C2(n4267), .A(n4204), .B(n4203), .ZN(n4205)
         );
  AOI21_X1 U4890 ( .B1(n4294), .B2(n4614), .A(n4205), .ZN(n4206) );
  OAI21_X1 U4891 ( .B1(n4207), .B2(n4296), .A(n4206), .ZN(U3225) );
  NAND2_X1 U4892 ( .A1(n2027), .A2(n4208), .ZN(n4210) );
  XNOR2_X1 U4893 ( .A(n4210), .B(n4209), .ZN(n4215) );
  NOR2_X1 U4894 ( .A1(n4476), .A2(n4276), .ZN(n4213) );
  INV_X1 U4895 ( .A(n4665), .ZN(n4242) );
  AOI22_X1 U4896 ( .A1(n4288), .A2(n4664), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n4211) );
  OAI21_X1 U4897 ( .B1(n4242), .B2(n4267), .A(n4211), .ZN(n4212) );
  AOI211_X1 U4898 ( .C1(n4262), .C2(n4473), .A(n4213), .B(n4212), .ZN(n4214)
         );
  OAI21_X1 U4899 ( .B1(n4215), .B2(n4296), .A(n4214), .ZN(U3226) );
  NOR2_X1 U4900 ( .A1(n2288), .A2(n2285), .ZN(n4217) );
  OAI22_X1 U4901 ( .A1(n4218), .A2(n2288), .B1(n4217), .B2(n4160), .ZN(n4222)
         );
  AOI22_X1 U4902 ( .A1(n4287), .A2(n4593), .B1(n4262), .B2(n4507), .ZN(n4220)
         );
  AOI22_X1 U4903 ( .A1(n4288), .A2(n4549), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n4219) );
  OAI211_X1 U4904 ( .C1(n4276), .C2(n4561), .A(n4220), .B(n4219), .ZN(n4221)
         );
  AOI21_X1 U4905 ( .B1(n4222), .B2(n4250), .A(n4221), .ZN(n4223) );
  INV_X1 U4906 ( .A(n4223), .ZN(U3230) );
  XOR2_X1 U4907 ( .A(n4226), .B(n4225), .Z(n4227) );
  XNOR2_X1 U4908 ( .A(n4224), .B(n4227), .ZN(n4235) );
  NAND2_X1 U4909 ( .A1(n4287), .A2(n4304), .ZN(n4230) );
  AND2_X1 U4910 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4330) );
  AOI21_X1 U4911 ( .B1(n4288), .B2(n4228), .A(n4330), .ZN(n4229) );
  OAI211_X1 U4912 ( .C1(n4231), .C2(n4291), .A(n4230), .B(n4229), .ZN(n4232)
         );
  AOI21_X1 U4913 ( .B1(n4294), .B2(n4233), .A(n4232), .ZN(n4234) );
  OAI21_X1 U4914 ( .B1(n4235), .B2(n4296), .A(n4234), .ZN(U3231) );
  AOI21_X1 U4915 ( .B1(n4238), .B2(n4237), .A(n4236), .ZN(n4246) );
  INV_X1 U4916 ( .A(n4239), .ZN(n4521) );
  OAI22_X1 U4917 ( .A1(n4241), .A2(n2896), .B1(STATE_REG_SCAN_IN), .B2(n4240), 
        .ZN(n4244) );
  OAI22_X1 U4918 ( .A1(n4242), .A2(n4291), .B1(n4551), .B2(n4267), .ZN(n4243)
         );
  AOI211_X1 U4919 ( .C1(n4521), .C2(n4294), .A(n4244), .B(n4243), .ZN(n4245)
         );
  OAI21_X1 U4920 ( .B1(n4246), .B2(n4296), .A(n4245), .ZN(U3232) );
  OAI21_X1 U4921 ( .B1(n4249), .B2(n4248), .A(n4247), .ZN(n4251) );
  NAND2_X1 U4922 ( .A1(n4251), .A2(n4250), .ZN(n4257) );
  AOI22_X1 U4923 ( .A1(n4287), .A2(n4253), .B1(n2013), .B2(n4288), .ZN(n4256)
         );
  AOI22_X1 U4924 ( .A1(n4254), .A2(REG3_REG_2__SCAN_IN), .B1(n4262), .B2(n4311), .ZN(n4255) );
  NAND3_X1 U4925 ( .A1(n4257), .A2(n4256), .A3(n4255), .ZN(U3234) );
  XNOR2_X1 U4926 ( .A(n4259), .B(n4258), .ZN(n4260) );
  XNOR2_X1 U4927 ( .A(n4134), .B(n4260), .ZN(n4270) );
  INV_X1 U4928 ( .A(n4261), .ZN(n4602) );
  NAND2_X1 U4929 ( .A1(n4262), .A2(n4593), .ZN(n4266) );
  AOI21_X1 U4930 ( .B1(n4288), .B2(n4264), .A(n4263), .ZN(n4265) );
  OAI211_X1 U4931 ( .C1(n4627), .C2(n4267), .A(n4266), .B(n4265), .ZN(n4268)
         );
  AOI21_X1 U4932 ( .B1(n4294), .B2(n4602), .A(n4268), .ZN(n4269) );
  OAI21_X1 U4933 ( .B1(n4270), .B2(n4296), .A(n4269), .ZN(U3235) );
  INV_X1 U4934 ( .A(n4271), .ZN(n4272) );
  NOR2_X1 U4935 ( .A1(n4273), .A2(n4272), .ZN(n4274) );
  XNOR2_X1 U4936 ( .A(n4275), .B(n4274), .ZN(n4281) );
  NOR2_X1 U4937 ( .A1(n4446), .A2(n4276), .ZN(n4279) );
  AOI22_X1 U4938 ( .A1(n4288), .A2(n4442), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4277) );
  OAI21_X1 U4939 ( .B1(n4438), .B2(n4291), .A(n4277), .ZN(n4278) );
  AOI211_X1 U4940 ( .C1(n4287), .C2(n4473), .A(n4279), .B(n4278), .ZN(n4280)
         );
  OAI21_X1 U4941 ( .B1(n4281), .B2(n4296), .A(n4280), .ZN(U3237) );
  INV_X1 U4942 ( .A(n4282), .ZN(n4284) );
  NAND2_X1 U4943 ( .A1(n4284), .A2(n4283), .ZN(n4286) );
  XNOR2_X1 U4944 ( .A(n4286), .B(n4285), .ZN(n4297) );
  NAND2_X1 U4945 ( .A1(n4287), .A2(n4716), .ZN(n4290) );
  AND2_X1 U4946 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4833) );
  AOI21_X1 U4947 ( .B1(n4288), .B2(n4715), .A(n4833), .ZN(n4289) );
  OAI211_X1 U4948 ( .C1(n4718), .C2(n4291), .A(n4290), .B(n4289), .ZN(n4292)
         );
  AOI21_X1 U4949 ( .B1(n4294), .B2(n4293), .A(n4292), .ZN(n4295) );
  OAI21_X1 U4950 ( .B1(n4297), .B2(n4296), .A(n4295), .ZN(U3238) );
  MUX2_X1 U4951 ( .A(DATAO_REG_31__SCAN_IN), .B(n4298), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4952 ( .A(DATAO_REG_30__SCAN_IN), .B(n4299), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4953 ( .A(DATAO_REG_29__SCAN_IN), .B(n4300), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4954 ( .A(DATAO_REG_28__SCAN_IN), .B(n4396), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4955 ( .A(DATAO_REG_27__SCAN_IN), .B(n4301), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4956 ( .A(DATAO_REG_26__SCAN_IN), .B(n4424), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4957 ( .A(DATAO_REG_25__SCAN_IN), .B(n4473), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4958 ( .A(DATAO_REG_24__SCAN_IN), .B(n4656), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4959 ( .A(DATAO_REG_23__SCAN_IN), .B(n4665), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4960 ( .A(DATAO_REG_20__SCAN_IN), .B(n4683), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4961 ( .A(DATAO_REG_18__SCAN_IN), .B(n4705), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4962 ( .A(DATAO_REG_17__SCAN_IN), .B(n4302), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4963 ( .A(DATAO_REG_16__SCAN_IN), .B(n4611), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4964 ( .A(DATAO_REG_15__SCAN_IN), .B(n4303), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4965 ( .A(DATAO_REG_13__SCAN_IN), .B(n4736), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4966 ( .A(DATAO_REG_12__SCAN_IN), .B(n4304), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4967 ( .A(DATAO_REG_10__SCAN_IN), .B(n4305), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4968 ( .A(DATAO_REG_9__SCAN_IN), .B(n4306), .S(U4043), .Z(U3559) );
  MUX2_X1 U4969 ( .A(DATAO_REG_8__SCAN_IN), .B(n4307), .S(U4043), .Z(U3558) );
  MUX2_X1 U4970 ( .A(DATAO_REG_6__SCAN_IN), .B(n4308), .S(U4043), .Z(U3556) );
  MUX2_X1 U4971 ( .A(DATAO_REG_5__SCAN_IN), .B(n4309), .S(U4043), .Z(U3555) );
  MUX2_X1 U4972 ( .A(DATAO_REG_4__SCAN_IN), .B(n4310), .S(U4043), .Z(U3554) );
  MUX2_X1 U4973 ( .A(DATAO_REG_3__SCAN_IN), .B(n4311), .S(U4043), .Z(U3553) );
  MUX2_X1 U4974 ( .A(DATAO_REG_2__SCAN_IN), .B(n4313), .S(U4043), .Z(U3552) );
  AOI211_X1 U4975 ( .C1(n4316), .C2(n4315), .A(n4314), .B(n4360), .ZN(n4317)
         );
  INV_X1 U4976 ( .A(n4317), .ZN(n4324) );
  AOI22_X1 U4977 ( .A1(n4846), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4323) );
  INV_X1 U4978 ( .A(n4852), .ZN(n4357) );
  NAND2_X1 U4979 ( .A1(n4357), .A2(n4821), .ZN(n4322) );
  OAI211_X1 U4980 ( .C1(n2380), .C2(n4320), .A(n4342), .B(n4319), .ZN(n4321)
         );
  NAND4_X1 U4981 ( .A1(n4324), .A2(n4323), .A3(n4322), .A4(n4321), .ZN(U3241)
         );
  XNOR2_X1 U4982 ( .A(n4813), .B(n4325), .ZN(n4326) );
  XNOR2_X1 U4983 ( .A(n4327), .B(n4326), .ZN(n4337) );
  AOI21_X1 U4984 ( .B1(n4329), .B2(n4328), .A(n4360), .ZN(n4335) );
  AOI21_X1 U4985 ( .B1(n4846), .B2(ADDR_REG_13__SCAN_IN), .A(n4330), .ZN(n4331) );
  OAI21_X1 U4986 ( .B1(n4852), .B2(n4332), .A(n4331), .ZN(n4333) );
  AOI21_X1 U4987 ( .B1(n4335), .B2(n4334), .A(n4333), .ZN(n4336) );
  OAI21_X1 U4988 ( .B1(n4840), .B2(n4337), .A(n4336), .ZN(U3253) );
  XOR2_X1 U4989 ( .A(REG1_REG_14__SCAN_IN), .B(n4338), .Z(n4347) );
  NOR2_X1 U4990 ( .A1(n4852), .A2(n4339), .ZN(n4340) );
  AOI211_X1 U4991 ( .C1(n4846), .C2(ADDR_REG_14__SCAN_IN), .A(n4341), .B(n4340), .ZN(n4346) );
  OAI211_X1 U4992 ( .C1(n4344), .C2(REG2_REG_14__SCAN_IN), .A(n4343), .B(n4342), .ZN(n4345) );
  OAI211_X1 U4993 ( .C1(n4347), .C2(n4360), .A(n4346), .B(n4345), .ZN(U3254)
         );
  AOI21_X1 U4994 ( .B1(n2030), .B2(n4349), .A(n4348), .ZN(n4361) );
  NOR2_X1 U4995 ( .A1(n4356), .A2(REG2_REG_17__SCAN_IN), .ZN(n4350) );
  AOI21_X1 U4996 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4356), .A(n4350), .ZN(n4353) );
  NAND2_X1 U4997 ( .A1(n4351), .A2(n4353), .ZN(n4352) );
  AOI221_X1 U4998 ( .B1(n4353), .B2(n4352), .C1(n4351), .C2(n4352), .A(n4840), 
        .ZN(n4354) );
  AOI211_X1 U4999 ( .C1(n4846), .C2(ADDR_REG_17__SCAN_IN), .A(n4355), .B(n4354), .ZN(n4359) );
  NAND2_X1 U5000 ( .A1(n4357), .A2(n4356), .ZN(n4358) );
  OAI211_X1 U5001 ( .C1(n4361), .C2(n4360), .A(n4359), .B(n4358), .ZN(U3257)
         );
  MUX2_X1 U5002 ( .A(REG2_REG_19__SCAN_IN), .B(n2671), .S(n3181), .Z(n4364) );
  XOR2_X1 U5003 ( .A(n4364), .B(n4363), .Z(n4377) );
  NAND2_X1 U5004 ( .A1(n4362), .A2(REG1_REG_18__SCAN_IN), .ZN(n4366) );
  INV_X1 U5005 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4368) );
  MUX2_X1 U5006 ( .A(n4368), .B(REG1_REG_19__SCAN_IN), .S(n3181), .Z(n4369) );
  NAND2_X1 U5007 ( .A1(n4846), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4371) );
  OAI211_X1 U5008 ( .C1(n4852), .C2(n4373), .A(n4372), .B(n4371), .ZN(n4374)
         );
  AOI21_X1 U5009 ( .B1(n4375), .B2(n4847), .A(n4374), .ZN(n4376) );
  OAI21_X1 U5010 ( .B1(n4377), .B2(n4840), .A(n4376), .ZN(U3259) );
  NAND2_X1 U5011 ( .A1(n4378), .A2(n4862), .ZN(n4381) );
  NOR2_X1 U5012 ( .A1(n4646), .A2(n4383), .ZN(n4379) );
  AOI21_X1 U5013 ( .B1(REG2_REG_31__SCAN_IN), .B2(n4646), .A(n4379), .ZN(n4380) );
  OAI211_X1 U5014 ( .C1(n4382), .C2(n4617), .A(n4381), .B(n4380), .ZN(U3260)
         );
  INV_X1 U5015 ( .A(n4383), .ZN(n4384) );
  AOI21_X1 U5016 ( .B1(n4386), .B2(n4724), .A(n4384), .ZN(n4750) );
  AOI21_X1 U5017 ( .B1(n4386), .B2(n2910), .A(n4385), .ZN(n4747) );
  NAND2_X1 U5018 ( .A1(n4747), .A2(n4862), .ZN(n4388) );
  NAND2_X1 U5019 ( .A1(n4624), .A2(REG2_REG_30__SCAN_IN), .ZN(n4387) );
  OAI211_X1 U5020 ( .C1(n4624), .C2(n4750), .A(n4388), .B(n4387), .ZN(U3261)
         );
  NAND2_X1 U5021 ( .A1(n4390), .A2(n4389), .ZN(n4392) );
  XNOR2_X1 U5022 ( .A(n4392), .B(n4391), .ZN(n4403) );
  OAI22_X1 U5023 ( .A1(n4394), .A2(n4617), .B1(n4556), .B2(n4393), .ZN(n4395)
         );
  AOI21_X1 U5024 ( .B1(n4396), .B2(n4612), .A(n4395), .ZN(n4402) );
  OAI22_X1 U5025 ( .A1(n4398), .A2(n4642), .B1(n4397), .B2(n4560), .ZN(n4399)
         );
  OAI21_X1 U5026 ( .B1(n4400), .B2(n4399), .A(n4556), .ZN(n4401) );
  OAI211_X1 U5027 ( .C1(n4403), .C2(n4605), .A(n4402), .B(n4401), .ZN(U3354)
         );
  NAND2_X1 U5028 ( .A1(n4404), .A2(n4644), .ZN(n4415) );
  NOR2_X1 U5029 ( .A1(n4405), .A2(n4642), .ZN(n4413) );
  NOR2_X1 U5030 ( .A1(n4617), .A2(n4406), .ZN(n4412) );
  OAI22_X1 U5031 ( .A1(n4408), .A2(n4560), .B1(n4407), .B2(n4556), .ZN(n4411)
         );
  OAI22_X1 U5032 ( .A1(n4409), .A2(n4537), .B1(n4438), .B2(n4535), .ZN(n4410)
         );
  NOR4_X1 U5033 ( .A1(n4413), .A2(n4412), .A3(n4411), .A4(n4410), .ZN(n4414)
         );
  OAI211_X1 U5034 ( .C1(n4624), .C2(n4416), .A(n4415), .B(n4414), .ZN(U3262)
         );
  NAND2_X1 U5035 ( .A1(n4417), .A2(n4644), .ZN(n4430) );
  INV_X1 U5036 ( .A(n4418), .ZN(n4428) );
  NOR2_X1 U5037 ( .A1(n4617), .A2(n4419), .ZN(n4423) );
  INV_X1 U5038 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4420) );
  OAI22_X1 U5039 ( .A1(n4421), .A2(n4560), .B1(n4420), .B2(n4556), .ZN(n4422)
         );
  AOI211_X1 U5040 ( .C1(n4612), .C2(n4424), .A(n4423), .B(n4422), .ZN(n4425)
         );
  OAI21_X1 U5041 ( .B1(n4426), .B2(n4537), .A(n4425), .ZN(n4427) );
  AOI21_X1 U5042 ( .B1(n4428), .B2(n4862), .A(n4427), .ZN(n4429) );
  OAI211_X1 U5043 ( .C1(n4624), .C2(n4431), .A(n4430), .B(n4429), .ZN(U3263)
         );
  XNOR2_X1 U5044 ( .A(n4432), .B(n4436), .ZN(n4652) );
  INV_X1 U5045 ( .A(n4652), .ZN(n4450) );
  NAND2_X1 U5046 ( .A1(n4434), .A2(n4433), .ZN(n4435) );
  XOR2_X1 U5047 ( .A(n4436), .B(n4435), .Z(n4441) );
  OAI22_X1 U5048 ( .A1(n4438), .A2(n4726), .B1(n4741), .B2(n4437), .ZN(n4439)
         );
  AOI21_X1 U5049 ( .B1(n4738), .B2(n4473), .A(n4439), .ZN(n4440) );
  OAI21_X1 U5050 ( .B1(n4441), .B2(n4631), .A(n4440), .ZN(n4651) );
  NAND2_X1 U5051 ( .A1(n4455), .A2(n4442), .ZN(n4443) );
  NAND2_X1 U5052 ( .A1(n4444), .A2(n4443), .ZN(n4754) );
  NOR2_X1 U5053 ( .A1(n4754), .A2(n4642), .ZN(n4448) );
  OAI22_X1 U5054 ( .A1(n4446), .A2(n4560), .B1(n4445), .B2(n4556), .ZN(n4447)
         );
  AOI211_X1 U5055 ( .C1(n4651), .C2(n4556), .A(n4448), .B(n4447), .ZN(n4449)
         );
  OAI21_X1 U5056 ( .B1(n4450), .B2(n4605), .A(n4449), .ZN(U3264) );
  XNOR2_X1 U5057 ( .A(n4451), .B(n4454), .ZN(n4452) );
  NAND2_X1 U5058 ( .A1(n4452), .A2(n4590), .ZN(n4658) );
  XNOR2_X1 U5059 ( .A(n4453), .B(n4454), .ZN(n4661) );
  NAND2_X1 U5060 ( .A1(n4661), .A2(n4644), .ZN(n4463) );
  OAI21_X1 U5061 ( .B1(n4472), .B2(n4456), .A(n4455), .ZN(n4758) );
  INV_X1 U5062 ( .A(n4758), .ZN(n4461) );
  OAI22_X1 U5063 ( .A1(n2331), .A2(n4535), .B1(n4617), .B2(n4456), .ZN(n4460)
         );
  AOI22_X1 U5064 ( .A1(n4457), .A2(n4859), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4646), .ZN(n4458) );
  OAI21_X1 U5065 ( .B1(n4659), .B2(n4537), .A(n4458), .ZN(n4459) );
  AOI211_X1 U5066 ( .C1(n4461), .C2(n4862), .A(n4460), .B(n4459), .ZN(n4462)
         );
  OAI211_X1 U5067 ( .C1(n4624), .C2(n4658), .A(n4463), .B(n4462), .ZN(U3265)
         );
  NAND2_X1 U5068 ( .A1(n4465), .A2(n4464), .ZN(n4466) );
  XOR2_X1 U5069 ( .A(n4469), .B(n4466), .Z(n4467) );
  NAND2_X1 U5070 ( .A1(n4467), .A2(n4590), .ZN(n4667) );
  XOR2_X1 U5071 ( .A(n4469), .B(n4468), .Z(n4670) );
  NAND2_X1 U5072 ( .A1(n4670), .A2(n4644), .ZN(n4483) );
  NOR2_X1 U5073 ( .A1(n4470), .A2(n4474), .ZN(n4471) );
  OR2_X1 U5074 ( .A1(n4472), .A2(n4471), .ZN(n4762) );
  INV_X1 U5075 ( .A(n4762), .ZN(n4481) );
  INV_X1 U5076 ( .A(n4473), .ZN(n4668) );
  NOR2_X1 U5077 ( .A1(n4617), .A2(n4474), .ZN(n4478) );
  INV_X1 U5078 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4475) );
  OAI22_X1 U5079 ( .A1(n4476), .A2(n4560), .B1(n4475), .B2(n4556), .ZN(n4477)
         );
  AOI211_X1 U5080 ( .C1(n4612), .C2(n4665), .A(n4478), .B(n4477), .ZN(n4479)
         );
  OAI21_X1 U5081 ( .B1(n4668), .B2(n4537), .A(n4479), .ZN(n4480) );
  AOI21_X1 U5082 ( .B1(n4481), .B2(n4862), .A(n4480), .ZN(n4482) );
  OAI211_X1 U5083 ( .C1(n4624), .C2(n4667), .A(n4483), .B(n4482), .ZN(U3266)
         );
  XNOR2_X1 U5084 ( .A(n4484), .B(n4491), .ZN(n4674) );
  INV_X1 U5085 ( .A(n4674), .ZN(n4505) );
  OR2_X1 U5086 ( .A1(n4485), .A2(n4486), .ZN(n4488) );
  NAND2_X1 U5087 ( .A1(n4488), .A2(n4487), .ZN(n4506) );
  INV_X1 U5088 ( .A(n4489), .ZN(n4490) );
  AOI21_X1 U5089 ( .B1(n4506), .B2(n4513), .A(n4490), .ZN(n4493) );
  INV_X1 U5090 ( .A(n4491), .ZN(n4492) );
  XNOR2_X1 U5091 ( .A(n4493), .B(n4492), .ZN(n4494) );
  NAND2_X1 U5092 ( .A1(n4494), .A2(n4590), .ZN(n4498) );
  AOI22_X1 U5093 ( .A1(n4496), .A2(n4738), .B1(n4724), .B2(n4495), .ZN(n4497)
         );
  OAI211_X1 U5094 ( .C1(n2331), .C2(n4726), .A(n4498), .B(n4497), .ZN(n4673)
         );
  NOR2_X1 U5095 ( .A1(n4516), .A2(n4499), .ZN(n4500) );
  OR2_X1 U5096 ( .A1(n4470), .A2(n4500), .ZN(n4766) );
  AOI22_X1 U5097 ( .A1(n4501), .A2(n4859), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4624), .ZN(n4502) );
  OAI21_X1 U5098 ( .B1(n4766), .B2(n4642), .A(n4502), .ZN(n4503) );
  AOI21_X1 U5099 ( .B1(n4673), .B2(n4556), .A(n4503), .ZN(n4504) );
  OAI21_X1 U5100 ( .B1(n4505), .B2(n4605), .A(n4504), .ZN(U3267) );
  XNOR2_X1 U5101 ( .A(n4506), .B(n4513), .ZN(n4511) );
  NAND2_X1 U5102 ( .A1(n4665), .A2(n4737), .ZN(n4509) );
  AOI22_X1 U5103 ( .A1(n4507), .A2(n4738), .B1(n4518), .B2(n4724), .ZN(n4508)
         );
  NAND2_X1 U5104 ( .A1(n4509), .A2(n4508), .ZN(n4510) );
  AOI21_X1 U5105 ( .B1(n4511), .B2(n4590), .A(n4510), .ZN(n4677) );
  NAND2_X1 U5106 ( .A1(n4512), .A2(n4513), .ZN(n4514) );
  NAND2_X1 U5107 ( .A1(n4515), .A2(n4514), .ZN(n4679) );
  INV_X1 U5108 ( .A(n4679), .ZN(n4524) );
  INV_X1 U5109 ( .A(n4516), .ZN(n4520) );
  NAND2_X1 U5110 ( .A1(n4530), .A2(n4518), .ZN(n4519) );
  NAND2_X1 U5111 ( .A1(n4520), .A2(n4519), .ZN(n4770) );
  AOI22_X1 U5112 ( .A1(n4521), .A2(n4859), .B1(REG2_REG_22__SCAN_IN), .B2(
        n4624), .ZN(n4522) );
  OAI21_X1 U5113 ( .B1(n4770), .B2(n4642), .A(n4522), .ZN(n4523) );
  AOI21_X1 U5114 ( .B1(n4524), .B2(n4644), .A(n4523), .ZN(n4525) );
  OAI21_X1 U5115 ( .B1(n4624), .B2(n4677), .A(n4525), .ZN(U3268) );
  INV_X1 U5116 ( .A(n4529), .ZN(n4526) );
  XNOR2_X1 U5117 ( .A(n4485), .B(n4526), .ZN(n4527) );
  NAND2_X1 U5118 ( .A1(n4527), .A2(n4590), .ZN(n4685) );
  XOR2_X1 U5119 ( .A(n4529), .B(n4528), .Z(n4688) );
  NAND2_X1 U5120 ( .A1(n4688), .A2(n4644), .ZN(n4542) );
  INV_X1 U5121 ( .A(n4557), .ZN(n4531) );
  OAI21_X1 U5122 ( .B1(n4531), .B2(n4534), .A(n4530), .ZN(n4774) );
  INV_X1 U5123 ( .A(n4774), .ZN(n4540) );
  AOI22_X1 U5124 ( .A1(n4624), .A2(REG2_REG_21__SCAN_IN), .B1(n4532), .B2(
        n4859), .ZN(n4533) );
  OAI21_X1 U5125 ( .B1(n4617), .B2(n4534), .A(n4533), .ZN(n4539) );
  OAI22_X1 U5126 ( .A1(n4686), .A2(n4537), .B1(n4536), .B2(n4535), .ZN(n4538)
         );
  AOI211_X1 U5127 ( .C1(n4540), .C2(n4862), .A(n4539), .B(n4538), .ZN(n4541)
         );
  OAI211_X1 U5128 ( .C1(n4624), .C2(n4685), .A(n4542), .B(n4541), .ZN(U3269)
         );
  XNOR2_X1 U5129 ( .A(n4543), .B(n4547), .ZN(n4691) );
  INV_X1 U5130 ( .A(n4544), .ZN(n4545) );
  NAND2_X1 U5131 ( .A1(n4546), .A2(n4545), .ZN(n4548) );
  XNOR2_X1 U5132 ( .A(n4548), .B(n4547), .ZN(n4553) );
  AOI22_X1 U5133 ( .A1(n4593), .A2(n4738), .B1(n4549), .B2(n4724), .ZN(n4550)
         );
  OAI21_X1 U5134 ( .B1(n4551), .B2(n4726), .A(n4550), .ZN(n4552) );
  AOI21_X1 U5135 ( .B1(n4553), .B2(n4590), .A(n4552), .ZN(n4554) );
  OAI21_X1 U5136 ( .B1(n4691), .B2(n4555), .A(n4554), .ZN(n4692) );
  NAND2_X1 U5137 ( .A1(n4692), .A2(n4556), .ZN(n4565) );
  INV_X1 U5138 ( .A(n4578), .ZN(n4559) );
  OAI21_X1 U5139 ( .B1(n4559), .B2(n4558), .A(n4557), .ZN(n4778) );
  INV_X1 U5140 ( .A(n4778), .ZN(n4563) );
  OAI22_X1 U5141 ( .A1(n4556), .A2(n3020), .B1(n4561), .B2(n4560), .ZN(n4562)
         );
  AOI21_X1 U5142 ( .B1(n4563), .B2(n4862), .A(n4562), .ZN(n4564) );
  OAI211_X1 U5143 ( .C1(n4691), .C2(n4566), .A(n4565), .B(n4564), .ZN(U3270)
         );
  NAND2_X1 U5144 ( .A1(n2039), .A2(n4567), .ZN(n4589) );
  INV_X1 U5145 ( .A(n4568), .ZN(n4570) );
  OAI21_X1 U5146 ( .B1(n4589), .B2(n4570), .A(n4569), .ZN(n4571) );
  XOR2_X1 U5147 ( .A(n4577), .B(n4571), .Z(n4575) );
  OAI22_X1 U5148 ( .A1(n4572), .A2(n4707), .B1(n4579), .B2(n4741), .ZN(n4573)
         );
  AOI21_X1 U5149 ( .B1(n4683), .B2(n4737), .A(n4573), .ZN(n4574) );
  OAI21_X1 U5150 ( .B1(n4575), .B2(n4631), .A(n4574), .ZN(n4696) );
  INV_X1 U5151 ( .A(n4696), .ZN(n4584) );
  XNOR2_X1 U5152 ( .A(n4576), .B(n4577), .ZN(n4697) );
  OAI21_X1 U5153 ( .B1(n4599), .B2(n4579), .A(n4578), .ZN(n4782) );
  AOI22_X1 U5154 ( .A1(n4646), .A2(REG2_REG_19__SCAN_IN), .B1(n4580), .B2(
        n4859), .ZN(n4581) );
  OAI21_X1 U5155 ( .B1(n4782), .B2(n4642), .A(n4581), .ZN(n4582) );
  AOI21_X1 U5156 ( .B1(n4697), .B2(n4644), .A(n4582), .ZN(n4583) );
  OAI21_X1 U5157 ( .B1(n4584), .B2(n4646), .A(n4583), .ZN(U3271) );
  NAND2_X1 U5158 ( .A1(n4585), .A2(n4588), .ZN(n4586) );
  NAND2_X1 U5159 ( .A1(n4587), .A2(n4586), .ZN(n4699) );
  INV_X1 U5160 ( .A(n4699), .ZN(n4606) );
  XNOR2_X1 U5161 ( .A(n4589), .B(n4588), .ZN(n4591) );
  NAND2_X1 U5162 ( .A1(n4591), .A2(n4590), .ZN(n4595) );
  OAI22_X1 U5163 ( .A1(n4627), .A2(n4707), .B1(n4741), .B2(n4598), .ZN(n4592)
         );
  AOI21_X1 U5164 ( .B1(n4737), .B2(n4593), .A(n4592), .ZN(n4594) );
  NAND2_X1 U5165 ( .A1(n4595), .A2(n4594), .ZN(n4703) );
  OAI21_X1 U5166 ( .B1(n4596), .B2(n4598), .A(n4597), .ZN(n4600) );
  OR2_X1 U5167 ( .A1(n4600), .A2(n4599), .ZN(n4700) );
  NOR2_X1 U5168 ( .A1(n4700), .A2(n3181), .ZN(n4601) );
  OAI21_X1 U5169 ( .B1(n4703), .B2(n4601), .A(n4556), .ZN(n4604) );
  AOI22_X1 U5170 ( .A1(n4624), .A2(REG2_REG_18__SCAN_IN), .B1(n4602), .B2(
        n4859), .ZN(n4603) );
  OAI211_X1 U5171 ( .C1(n4606), .C2(n4605), .A(n4604), .B(n4603), .ZN(U3272)
         );
  XNOR2_X1 U5172 ( .A(n4607), .B(n4610), .ZN(n4608) );
  NOR2_X1 U5173 ( .A1(n4608), .A2(n4631), .ZN(n4708) );
  INV_X1 U5174 ( .A(n4708), .ZN(n4625) );
  XNOR2_X1 U5175 ( .A(n4609), .B(n4610), .ZN(n4710) );
  AOI22_X1 U5176 ( .A1(n4613), .A2(n4705), .B1(n4612), .B2(n4611), .ZN(n4616)
         );
  AOI22_X1 U5177 ( .A1(n4624), .A2(REG2_REG_17__SCAN_IN), .B1(n4614), .B2(
        n4859), .ZN(n4615) );
  OAI211_X1 U5178 ( .C1(n4620), .C2(n4617), .A(n4616), .B(n4615), .ZN(n4622)
         );
  INV_X1 U5179 ( .A(n4596), .ZN(n4619) );
  OAI21_X1 U5180 ( .B1(n2186), .B2(n4620), .A(n4619), .ZN(n4787) );
  NOR2_X1 U5181 ( .A1(n4787), .A2(n4642), .ZN(n4621) );
  AOI211_X1 U5182 ( .C1(n4710), .C2(n4644), .A(n4622), .B(n4621), .ZN(n4623)
         );
  OAI21_X1 U5183 ( .B1(n4625), .B2(n4624), .A(n4623), .ZN(U3273) );
  XNOR2_X1 U5184 ( .A(n4626), .B(n4637), .ZN(n4632) );
  OAI22_X1 U5185 ( .A1(n4627), .A2(n4726), .B1(n4727), .B2(n4707), .ZN(n4628)
         );
  AOI21_X1 U5186 ( .B1(n4629), .B2(n4724), .A(n4628), .ZN(n4630) );
  OAI21_X1 U5187 ( .B1(n4632), .B2(n4631), .A(n4630), .ZN(n4712) );
  INV_X1 U5188 ( .A(n4712), .ZN(n4647) );
  INV_X1 U5189 ( .A(n4635), .ZN(n4636) );
  AOI21_X1 U5190 ( .B1(n4637), .B2(n4633), .A(n4636), .ZN(n4713) );
  OAI21_X1 U5191 ( .B1(n2895), .B2(n4639), .A(n4618), .ZN(n4791) );
  AOI22_X1 U5192 ( .A1(n4646), .A2(REG2_REG_16__SCAN_IN), .B1(n4640), .B2(
        n4859), .ZN(n4641) );
  OAI21_X1 U5193 ( .B1(n4791), .B2(n4642), .A(n4641), .ZN(n4643) );
  AOI21_X1 U5194 ( .B1(n4713), .B2(n4644), .A(n4643), .ZN(n4645) );
  OAI21_X1 U5195 ( .B1(n4647), .B2(n4646), .A(n4645), .ZN(U3274) );
  MUX2_X1 U5196 ( .A(REG1_REG_31__SCAN_IN), .B(n4648), .S(n4915), .Z(U3549) );
  NAND2_X1 U5197 ( .A1(n4747), .A2(n2901), .ZN(n4650) );
  NAND2_X1 U5198 ( .A1(n4912), .A2(REG1_REG_30__SCAN_IN), .ZN(n4649) );
  OAI211_X1 U5199 ( .C1(n4750), .C2(n4912), .A(n4650), .B(n4649), .ZN(U3548)
         );
  INV_X1 U5200 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4653) );
  AOI21_X1 U5201 ( .B1(n4652), .B2(n4900), .A(n4651), .ZN(n4751) );
  MUX2_X1 U5202 ( .A(n4653), .B(n4751), .S(n4915), .Z(n4654) );
  OAI21_X1 U5203 ( .B1(n4746), .B2(n4754), .A(n4654), .ZN(U3544) );
  INV_X1 U5204 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4662) );
  AOI22_X1 U5205 ( .A1(n4656), .A2(n4738), .B1(n4724), .B2(n4655), .ZN(n4657)
         );
  OAI211_X1 U5206 ( .C1(n4659), .C2(n4726), .A(n4658), .B(n4657), .ZN(n4660)
         );
  AOI21_X1 U5207 ( .B1(n4661), .B2(n4900), .A(n4660), .ZN(n4755) );
  MUX2_X1 U5208 ( .A(n4662), .B(n4755), .S(n4915), .Z(n4663) );
  OAI21_X1 U5209 ( .B1(n4746), .B2(n4758), .A(n4663), .ZN(U3543) );
  AOI22_X1 U5210 ( .A1(n4665), .A2(n4738), .B1(n4724), .B2(n4664), .ZN(n4666)
         );
  OAI211_X1 U5211 ( .C1(n4668), .C2(n4726), .A(n4667), .B(n4666), .ZN(n4669)
         );
  AOI21_X1 U5212 ( .B1(n4670), .B2(n4900), .A(n4669), .ZN(n4759) );
  MUX2_X1 U5213 ( .A(n4671), .B(n4759), .S(n4915), .Z(n4672) );
  OAI21_X1 U5214 ( .B1(n4746), .B2(n4762), .A(n4672), .ZN(U3542) );
  AOI21_X1 U5215 ( .B1(n4674), .B2(n4900), .A(n4673), .ZN(n4764) );
  INV_X1 U5216 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4675) );
  MUX2_X1 U5217 ( .A(n4764), .B(n4675), .S(n4912), .Z(n4676) );
  OAI21_X1 U5218 ( .B1(n4746), .B2(n4766), .A(n4676), .ZN(U3541) );
  OAI21_X1 U5219 ( .B1(n4679), .B2(n4678), .A(n4677), .ZN(n4767) );
  MUX2_X1 U5220 ( .A(REG1_REG_22__SCAN_IN), .B(n4767), .S(n4915), .Z(n4680) );
  INV_X1 U5221 ( .A(n4680), .ZN(n4681) );
  OAI21_X1 U5222 ( .B1(n4746), .B2(n4770), .A(n4681), .ZN(U3540) );
  INV_X1 U5223 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4689) );
  AOI22_X1 U5224 ( .A1(n4683), .A2(n4738), .B1(n4682), .B2(n4724), .ZN(n4684)
         );
  OAI211_X1 U5225 ( .C1(n4686), .C2(n4726), .A(n4685), .B(n4684), .ZN(n4687)
         );
  AOI21_X1 U5226 ( .B1(n4688), .B2(n4900), .A(n4687), .ZN(n4771) );
  MUX2_X1 U5227 ( .A(n4689), .B(n4771), .S(n4915), .Z(n4690) );
  OAI21_X1 U5228 ( .B1(n4746), .B2(n4774), .A(n4690), .ZN(U3539) );
  INV_X1 U5229 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4694) );
  INV_X1 U5230 ( .A(n4691), .ZN(n4693) );
  AOI21_X1 U5231 ( .B1(n4896), .B2(n4693), .A(n4692), .ZN(n4775) );
  MUX2_X1 U5232 ( .A(n4694), .B(n4775), .S(n4915), .Z(n4695) );
  OAI21_X1 U5233 ( .B1(n4746), .B2(n4778), .A(n4695), .ZN(U3538) );
  AOI21_X1 U5234 ( .B1(n4900), .B2(n4697), .A(n4696), .ZN(n4779) );
  MUX2_X1 U5235 ( .A(n4368), .B(n4779), .S(n4915), .Z(n4698) );
  OAI21_X1 U5236 ( .B1(n4746), .B2(n4782), .A(n4698), .ZN(U3537) );
  NAND2_X1 U5237 ( .A1(n4699), .A2(n4900), .ZN(n4701) );
  NAND2_X1 U5238 ( .A1(n4701), .A2(n4700), .ZN(n4702) );
  MUX2_X1 U5239 ( .A(n4783), .B(REG1_REG_18__SCAN_IN), .S(n4912), .Z(U3536) );
  AOI22_X1 U5240 ( .A1(n4705), .A2(n4737), .B1(n4704), .B2(n4724), .ZN(n4706)
         );
  OAI21_X1 U5241 ( .B1(n4718), .B2(n4707), .A(n4706), .ZN(n4709) );
  AOI211_X1 U5242 ( .C1(n4710), .C2(n4900), .A(n4709), .B(n4708), .ZN(n4784)
         );
  MUX2_X1 U5243 ( .A(n2507), .B(n4784), .S(n4915), .Z(n4711) );
  OAI21_X1 U5244 ( .B1(n4746), .B2(n4787), .A(n4711), .ZN(U3535) );
  AOI21_X1 U5245 ( .B1(n4713), .B2(n4900), .A(n4712), .ZN(n4788) );
  MUX2_X1 U5246 ( .A(n2238), .B(n4788), .S(n4915), .Z(n4714) );
  OAI21_X1 U5247 ( .B1(n4746), .B2(n4791), .A(n4714), .ZN(U3534) );
  AOI22_X1 U5248 ( .A1(n4716), .A2(n4738), .B1(n4724), .B2(n4715), .ZN(n4717)
         );
  OAI21_X1 U5249 ( .B1(n4718), .B2(n4726), .A(n4717), .ZN(n4720) );
  AOI211_X1 U5250 ( .C1(n4900), .C2(n4721), .A(n4720), .B(n4719), .ZN(n4792)
         );
  MUX2_X1 U5251 ( .A(n2503), .B(n4792), .S(n4915), .Z(n4722) );
  OAI21_X1 U5252 ( .B1(n4746), .B2(n4795), .A(n4722), .ZN(U3533) );
  AOI22_X1 U5253 ( .A1(n4724), .A2(n4723), .B1(n4738), .B2(n4736), .ZN(n4725)
         );
  OAI21_X1 U5254 ( .B1(n4727), .B2(n4726), .A(n4725), .ZN(n4729) );
  AOI211_X1 U5255 ( .C1(n4896), .C2(n4730), .A(n4729), .B(n4728), .ZN(n4796)
         );
  MUX2_X1 U5256 ( .A(n4731), .B(n4796), .S(n4915), .Z(n4732) );
  OAI21_X1 U5257 ( .B1(n4746), .B2(n4799), .A(n4732), .ZN(U3532) );
  AOI21_X1 U5258 ( .B1(n4900), .B2(n4734), .A(n4733), .ZN(n4800) );
  MUX2_X1 U5259 ( .A(n2499), .B(n4800), .S(n4915), .Z(n4735) );
  OAI21_X1 U5260 ( .B1(n4746), .B2(n4803), .A(n4735), .ZN(U3531) );
  AOI22_X1 U5261 ( .A1(n4739), .A2(n4738), .B1(n4737), .B2(n4736), .ZN(n4740)
         );
  OAI21_X1 U5262 ( .B1(n2893), .B2(n4741), .A(n4740), .ZN(n4743) );
  AOI211_X1 U5263 ( .C1(n4900), .C2(n4744), .A(n4743), .B(n4742), .ZN(n4804)
         );
  MUX2_X1 U5264 ( .A(n2235), .B(n4804), .S(n4915), .Z(n4745) );
  OAI21_X1 U5265 ( .B1(n4746), .B2(n4808), .A(n4745), .ZN(U3530) );
  NAND2_X1 U5266 ( .A1(n4747), .A2(n4889), .ZN(n4749) );
  NAND2_X1 U5267 ( .A1(n4905), .A2(REG0_REG_30__SCAN_IN), .ZN(n4748) );
  OAI211_X1 U5268 ( .C1(n4750), .C2(n4905), .A(n4749), .B(n4748), .ZN(U3516)
         );
  INV_X1 U5269 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4752) );
  MUX2_X1 U5270 ( .A(n4752), .B(n4751), .S(n4907), .Z(n4753) );
  OAI21_X1 U5271 ( .B1(n4754), .B2(n4807), .A(n4753), .ZN(U3512) );
  INV_X1 U5272 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4756) );
  MUX2_X1 U5273 ( .A(n4756), .B(n4755), .S(n4907), .Z(n4757) );
  OAI21_X1 U5274 ( .B1(n4758), .B2(n4807), .A(n4757), .ZN(U3511) );
  INV_X1 U5275 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4760) );
  MUX2_X1 U5276 ( .A(n4760), .B(n4759), .S(n4907), .Z(n4761) );
  OAI21_X1 U5277 ( .B1(n4762), .B2(n4807), .A(n4761), .ZN(U3510) );
  INV_X1 U5278 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4763) );
  MUX2_X1 U5279 ( .A(n4764), .B(n4763), .S(n4905), .Z(n4765) );
  OAI21_X1 U5280 ( .B1(n4766), .B2(n4807), .A(n4765), .ZN(U3509) );
  MUX2_X1 U5281 ( .A(REG0_REG_22__SCAN_IN), .B(n4767), .S(n4907), .Z(n4768) );
  INV_X1 U5282 ( .A(n4768), .ZN(n4769) );
  OAI21_X1 U5283 ( .B1(n4770), .B2(n4807), .A(n4769), .ZN(U3508) );
  INV_X1 U5284 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4772) );
  MUX2_X1 U5285 ( .A(n4772), .B(n4771), .S(n4907), .Z(n4773) );
  OAI21_X1 U5286 ( .B1(n4774), .B2(n4807), .A(n4773), .ZN(U3507) );
  MUX2_X1 U5287 ( .A(n4776), .B(n4775), .S(n4907), .Z(n4777) );
  OAI21_X1 U5288 ( .B1(n4778), .B2(n4807), .A(n4777), .ZN(U3506) );
  INV_X1 U5289 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4780) );
  MUX2_X1 U5290 ( .A(n4780), .B(n4779), .S(n4907), .Z(n4781) );
  OAI21_X1 U5291 ( .B1(n4782), .B2(n4807), .A(n4781), .ZN(U3505) );
  MUX2_X1 U5292 ( .A(n4783), .B(REG0_REG_18__SCAN_IN), .S(n4905), .Z(U3503) );
  INV_X1 U5293 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4785) );
  MUX2_X1 U5294 ( .A(n4785), .B(n4784), .S(n4907), .Z(n4786) );
  OAI21_X1 U5295 ( .B1(n4787), .B2(n4807), .A(n4786), .ZN(U3501) );
  INV_X1 U5296 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4789) );
  MUX2_X1 U5297 ( .A(n4789), .B(n4788), .S(n4907), .Z(n4790) );
  OAI21_X1 U5298 ( .B1(n4791), .B2(n4807), .A(n4790), .ZN(U3499) );
  INV_X1 U5299 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4793) );
  MUX2_X1 U5300 ( .A(n4793), .B(n4792), .S(n4907), .Z(n4794) );
  OAI21_X1 U5301 ( .B1(n4795), .B2(n4807), .A(n4794), .ZN(U3497) );
  MUX2_X1 U5302 ( .A(n4797), .B(n4796), .S(n4907), .Z(n4798) );
  OAI21_X1 U5303 ( .B1(n4799), .B2(n4807), .A(n4798), .ZN(U3495) );
  INV_X1 U5304 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4801) );
  MUX2_X1 U5305 ( .A(n4801), .B(n4800), .S(n4907), .Z(n4802) );
  OAI21_X1 U5306 ( .B1(n4803), .B2(n4807), .A(n4802), .ZN(U3493) );
  INV_X1 U5307 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4805) );
  MUX2_X1 U5308 ( .A(n4805), .B(n4804), .S(n4907), .Z(n4806) );
  OAI21_X1 U5309 ( .B1(n4808), .B2(n4807), .A(n4806), .ZN(U3491) );
  MUX2_X1 U5310 ( .A(n4809), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5311 ( .A(DATAI_27_), .B(n4810), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5312 ( .A(n2862), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5313 ( .A(n4811), .B(DATAI_20_), .S(U3149), .Z(U3332) );
  MUX2_X1 U5314 ( .A(DATAI_19_), .B(n3181), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5315 ( .A(DATAI_14_), .B(n4812), .S(STATE_REG_SCAN_IN), .Z(U3338)
         );
  MUX2_X1 U5316 ( .A(n4813), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5317 ( .A(DATAI_12_), .B(n4814), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5318 ( .A(DATAI_11_), .B(n4815), .S(STATE_REG_SCAN_IN), .Z(U3341)
         );
  MUX2_X1 U5319 ( .A(n4816), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5320 ( .A(n4817), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5321 ( .A(DATAI_7_), .B(n4818), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5322 ( .A(n4819), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5323 ( .A(DATAI_4_), .B(n4820), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5324 ( .A(DATAI_2_), .B(n2010), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U5325 ( .A(n4821), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U5326 ( .A1(STATE_REG_SCAN_IN), .A2(n4822), .B1(n2780), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U5327 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4908) );
  AOI21_X1 U5328 ( .B1(n4908), .B2(n4824), .A(n4823), .ZN(n4825) );
  XNOR2_X1 U5329 ( .A(n4825), .B(n2379), .ZN(n4827) );
  AOI22_X1 U5330 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4846), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4826) );
  OAI21_X1 U5331 ( .B1(n4828), .B2(n4827), .A(n4826), .ZN(U3240) );
  AOI211_X1 U5332 ( .C1(n4831), .C2(n4830), .A(n4829), .B(n4840), .ZN(n4832)
         );
  AOI211_X1 U5333 ( .C1(ADDR_REG_15__SCAN_IN), .C2(n4846), .A(n4833), .B(n4832), .ZN(n4838) );
  OAI211_X1 U5334 ( .C1(n4836), .C2(n4835), .A(n4847), .B(n4834), .ZN(n4837)
         );
  OAI211_X1 U5335 ( .C1(n4852), .C2(n4879), .A(n4838), .B(n4837), .ZN(U3255)
         );
  INV_X1 U5336 ( .A(n4839), .ZN(n4845) );
  AOI221_X1 U5337 ( .B1(n4843), .B2(n4842), .C1(n4841), .C2(n4842), .A(n4840), 
        .ZN(n4844) );
  AOI211_X1 U5338 ( .C1(n4846), .C2(ADDR_REG_16__SCAN_IN), .A(n4845), .B(n4844), .ZN(n4851) );
  OAI221_X1 U5339 ( .B1(n4849), .B2(REG1_REG_16__SCAN_IN), .C1(n4849), .C2(
        n4848), .A(n4847), .ZN(n4850) );
  OAI211_X1 U5340 ( .C1(n4852), .C2(n4877), .A(n4851), .B(n4850), .ZN(U3256)
         );
  AOI22_X1 U5341 ( .A1(n4646), .A2(REG2_REG_3__SCAN_IN), .B1(n4859), .B2(n4853), .ZN(n4857) );
  AOI22_X1 U5342 ( .A1(n4862), .A2(n4855), .B1(n4861), .B2(n4854), .ZN(n4856)
         );
  OAI211_X1 U5343 ( .C1(n4646), .C2(n4858), .A(n4857), .B(n4856), .ZN(U3287)
         );
  AOI22_X1 U5344 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4646), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4859), .ZN(n4864) );
  AOI22_X1 U5345 ( .A1(n4862), .A2(n4888), .B1(n4861), .B2(n4860), .ZN(n4863)
         );
  OAI211_X1 U5346 ( .C1(n4646), .C2(n4865), .A(n4864), .B(n4863), .ZN(U3288)
         );
  AND2_X1 U5347 ( .A1(D_REG_31__SCAN_IN), .A2(n4870), .ZN(U3291) );
  INV_X1 U5348 ( .A(n4870), .ZN(n4872) );
  NOR2_X1 U5349 ( .A1(n4872), .A2(n4866), .ZN(U3292) );
  AND2_X1 U5350 ( .A1(D_REG_29__SCAN_IN), .A2(n4870), .ZN(U3293) );
  AND2_X1 U5351 ( .A1(D_REG_28__SCAN_IN), .A2(n4870), .ZN(U3294) );
  AND2_X1 U5352 ( .A1(D_REG_27__SCAN_IN), .A2(n4870), .ZN(U3295) );
  AND2_X1 U5353 ( .A1(D_REG_26__SCAN_IN), .A2(n4870), .ZN(U3296) );
  NOR2_X1 U5354 ( .A1(n4872), .A2(n4867), .ZN(U3297) );
  AND2_X1 U5355 ( .A1(D_REG_24__SCAN_IN), .A2(n4870), .ZN(U3298) );
  AND2_X1 U5356 ( .A1(D_REG_23__SCAN_IN), .A2(n4870), .ZN(U3299) );
  AND2_X1 U5357 ( .A1(D_REG_22__SCAN_IN), .A2(n4870), .ZN(U3300) );
  AND2_X1 U5358 ( .A1(D_REG_21__SCAN_IN), .A2(n4870), .ZN(U3301) );
  AND2_X1 U5359 ( .A1(D_REG_20__SCAN_IN), .A2(n4870), .ZN(U3302) );
  AND2_X1 U5360 ( .A1(D_REG_19__SCAN_IN), .A2(n4870), .ZN(U3303) );
  AND2_X1 U5361 ( .A1(D_REG_18__SCAN_IN), .A2(n4870), .ZN(U3304) );
  AND2_X1 U5362 ( .A1(D_REG_17__SCAN_IN), .A2(n4870), .ZN(U3305) );
  AND2_X1 U5363 ( .A1(D_REG_16__SCAN_IN), .A2(n4870), .ZN(U3306) );
  AND2_X1 U5364 ( .A1(D_REG_15__SCAN_IN), .A2(n4870), .ZN(U3307) );
  AND2_X1 U5365 ( .A1(D_REG_14__SCAN_IN), .A2(n4870), .ZN(U3308) );
  AND2_X1 U5366 ( .A1(D_REG_13__SCAN_IN), .A2(n4870), .ZN(U3309) );
  NOR2_X1 U5367 ( .A1(n4872), .A2(n4868), .ZN(U3310) );
  AND2_X1 U5368 ( .A1(D_REG_11__SCAN_IN), .A2(n4870), .ZN(U3311) );
  NOR2_X1 U5369 ( .A1(n4872), .A2(n4869), .ZN(U3312) );
  AND2_X1 U5370 ( .A1(D_REG_9__SCAN_IN), .A2(n4870), .ZN(U3313) );
  AND2_X1 U5371 ( .A1(D_REG_8__SCAN_IN), .A2(n4870), .ZN(U3314) );
  AND2_X1 U5372 ( .A1(D_REG_7__SCAN_IN), .A2(n4870), .ZN(U3315) );
  AND2_X1 U5373 ( .A1(D_REG_6__SCAN_IN), .A2(n4870), .ZN(U3316) );
  AND2_X1 U5374 ( .A1(D_REG_5__SCAN_IN), .A2(n4870), .ZN(U3317) );
  AND2_X1 U5375 ( .A1(D_REG_4__SCAN_IN), .A2(n4870), .ZN(U3318) );
  AND2_X1 U5376 ( .A1(D_REG_3__SCAN_IN), .A2(n4870), .ZN(U3319) );
  NOR2_X1 U5377 ( .A1(n4872), .A2(n4871), .ZN(U3320) );
  AOI21_X1 U5378 ( .B1(U3149), .B2(n2729), .A(n4873), .ZN(U3329) );
  AOI22_X1 U5379 ( .A1(STATE_REG_SCAN_IN), .A2(n4875), .B1(n4874), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5380 ( .A(DATAI_16_), .ZN(n4876) );
  AOI22_X1 U5381 ( .A1(STATE_REG_SCAN_IN), .A2(n4877), .B1(n4876), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5382 ( .A1(STATE_REG_SCAN_IN), .A2(n4879), .B1(n4878), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5383 ( .A1(STATE_REG_SCAN_IN), .A2(n2333), .B1(n2540), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5384 ( .A(n4880), .ZN(n4883) );
  INV_X1 U5385 ( .A(n4881), .ZN(n4882) );
  AOI211_X1 U5386 ( .C1(n4896), .C2(n4884), .A(n4883), .B(n4882), .ZN(n4909)
         );
  AOI22_X1 U5387 ( .A1(n4907), .A2(n4909), .B1(n4885), .B2(n4905), .ZN(U3467)
         );
  INV_X1 U5388 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4886) );
  AOI22_X1 U5389 ( .A1(n4907), .A2(n4887), .B1(n4886), .B2(n4905), .ZN(U3469)
         );
  AOI22_X1 U5390 ( .A1(n4890), .A2(n4907), .B1(n4889), .B2(n4888), .ZN(n4891)
         );
  OAI21_X1 U5391 ( .B1(n4907), .B2(n4892), .A(n4891), .ZN(U3471) );
  INV_X1 U5392 ( .A(n4893), .ZN(n4895) );
  AOI211_X1 U5393 ( .C1(n4897), .C2(n4896), .A(n4895), .B(n4894), .ZN(n4911)
         );
  AOI22_X1 U5394 ( .A1(n4907), .A2(n4911), .B1(n4898), .B2(n4905), .ZN(U3475)
         );
  AND3_X1 U5395 ( .A1(n4901), .A2(n4900), .A3(n4899), .ZN(n4902) );
  NOR3_X1 U5396 ( .A1(n4904), .A2(n4903), .A3(n4902), .ZN(n4914) );
  INV_X1 U5397 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4906) );
  AOI22_X1 U5398 ( .A1(n4907), .A2(n4914), .B1(n4906), .B2(n4905), .ZN(U3481)
         );
  AOI22_X1 U5399 ( .A1(n4915), .A2(n4909), .B1(n4908), .B2(n4912), .ZN(U3518)
         );
  AOI22_X1 U5400 ( .A1(n4915), .A2(n4911), .B1(n4910), .B2(n4912), .ZN(U3522)
         );
  AOI22_X1 U5401 ( .A1(n4915), .A2(n4914), .B1(n4913), .B2(n4912), .ZN(U3525)
         );
  CLKBUF_X3 U2251 ( .A(n4252), .Z(n2013) );
  CLKBUF_X1 U2295 ( .A(n2485), .Z(n2010) );
endmodule

