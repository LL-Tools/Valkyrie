

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5028, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11101;

  NAND2_X1 U5093 ( .A1(n6372), .A2(n6371), .ZN(n10455) );
  NAND2_X1 U5094 ( .A1(n5141), .A2(n5140), .ZN(n10894) );
  AOI21_X1 U5095 ( .B1(n5167), .B2(n7848), .A(n7025), .ZN(n7738) );
  NAND2_X1 U5096 ( .A1(n6473), .A2(n8779), .ZN(n6906) );
  NAND2_X1 U5097 ( .A1(n8256), .A2(n8800), .ZN(n8920) );
  NAND2_X1 U5098 ( .A1(n5937), .A2(n5936), .ZN(n5959) );
  CLKBUF_X2 U5099 ( .A(n6573), .Z(n5030) );
  AND2_X1 U5100 ( .A1(n6508), .A2(n6524), .ZN(n10683) );
  AND2_X2 U5101 ( .A1(n6373), .A2(n5687), .ZN(n6063) );
  NAND2_X2 U5102 ( .A1(n7425), .A2(n7424), .ZN(n10545) );
  INV_X1 U5103 ( .A(n11101), .ZN(n5028) );
  INV_X2 U5104 ( .A(n5028), .ZN(P1_U3084) );
  INV_X1 U5105 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n11101) );
  NAND2_X1 U5106 ( .A1(n7026), .A2(n7222), .ZN(n7787) );
  INV_X1 U5107 ( .A(n5030), .ZN(n6768) );
  AND2_X1 U5108 ( .A1(n10103), .A2(n6240), .ZN(n6263) );
  INV_X1 U5109 ( .A(n6342), .ZN(n5686) );
  INV_X1 U5111 ( .A(n8780), .ZN(n6521) );
  NAND2_X1 U5112 ( .A1(n9062), .A2(n6820), .ZN(n9109) );
  NOR2_X1 U5114 ( .A1(n9919), .A2(n9300), .ZN(n9285) );
  INV_X1 U5115 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n10002) );
  CLKBUF_X2 U5116 ( .A(n5758), .Z(n6303) );
  NAND4_X2 U5117 ( .A1(n5723), .A2(n5722), .A3(n5721), .A4(n5720), .ZN(n5727)
         );
  OR2_X2 U5118 ( .A1(n5959), .A2(n5313), .ZN(n5312) );
  NAND2_X2 U5119 ( .A1(n6138), .A2(n6137), .ZN(n6168) );
  OAI21_X4 U5120 ( .B1(n7787), .B2(n7028), .A(n7027), .ZN(n7901) );
  AND2_X4 U5121 ( .A1(n8697), .A2(n6483), .ZN(n6533) );
  INV_X1 U5122 ( .A(n5727), .ZN(n7745) );
  AOI22_X2 U5123 ( .A1(n5282), .A2(n5799), .B1(n5283), .B2(n5280), .ZN(n5821)
         );
  XNOR2_X1 U5124 ( .A(n8094), .B(n10168), .ZN(n8084) );
  NAND2_X2 U5125 ( .A1(n5942), .A2(n5941), .ZN(n8094) );
  INV_X2 U5127 ( .A(n8188), .ZN(n8190) );
  AND2_X1 U5128 ( .A1(n6373), .A2(n5687), .ZN(n5031) );
  NOR2_X1 U5129 ( .A1(n9361), .A2(n9360), .ZN(n9359) );
  INV_X1 U5130 ( .A(n7930), .ZN(n10825) );
  INV_X1 U5131 ( .A(n10174), .ZN(n7772) );
  CLKBUF_X2 U5132 ( .A(n5688), .Z(n6384) );
  INV_X1 U5134 ( .A(n7015), .ZN(n5175) );
  XNOR2_X1 U5136 ( .A(n5677), .B(n9808), .ZN(n7264) );
  AND2_X1 U5137 ( .A1(n5182), .A2(n5181), .ZN(n5676) );
  AOI21_X1 U5139 ( .B1(n5376), .B2(n11009), .A(n5117), .ZN(n10453) );
  NAND2_X1 U5140 ( .A1(n5227), .A2(n9259), .ZN(n9316) );
  NAND2_X1 U5141 ( .A1(n6191), .A2(n6190), .ZN(n10037) );
  NAND2_X1 U5142 ( .A1(n9359), .A2(n9256), .ZN(n5228) );
  AND2_X1 U5143 ( .A1(n5378), .A2(n5190), .ZN(n10337) );
  NAND2_X1 U5144 ( .A1(n9836), .A2(n9835), .ZN(n9834) );
  AND2_X1 U5145 ( .A1(n5207), .A2(n5206), .ZN(n9836) );
  NAND2_X1 U5146 ( .A1(n5209), .A2(n5208), .ZN(n8677) );
  NAND2_X1 U5147 ( .A1(n6822), .A2(n6821), .ZN(n9945) );
  NAND2_X1 U5148 ( .A1(n8477), .A2(n6674), .ZN(n8720) );
  NAND2_X1 U5149 ( .A1(n6272), .A2(n6271), .ZN(n10476) );
  NAND2_X1 U5150 ( .A1(n6810), .A2(n6809), .ZN(n9950) );
  OAI21_X1 U5151 ( .B1(n5607), .B2(n5604), .A(n9250), .ZN(n5603) );
  OAI21_X1 U5152 ( .B1(n8454), .B2(n5219), .A(n5217), .ZN(n5226) );
  OR2_X1 U5153 ( .A1(n8641), .A2(n11051), .ZN(n8642) );
  AOI21_X1 U5154 ( .B1(n5417), .B2(n5039), .A(n5116), .ZN(n5416) );
  NAND2_X1 U5155 ( .A1(n6738), .A2(n6737), .ZN(n9977) );
  NAND2_X1 U5156 ( .A1(n5409), .A2(n5408), .ZN(n7979) );
  NAND2_X1 U5157 ( .A1(n8027), .A2(n6546), .ZN(n8028) );
  NAND2_X1 U5158 ( .A1(n5470), .A2(n5468), .ZN(n9888) );
  OAI21_X1 U5159 ( .B1(n7664), .B2(n5504), .A(n5505), .ZN(n5806) );
  NAND2_X1 U5160 ( .A1(n6069), .A2(n6068), .ZN(n10135) );
  OR2_X1 U5161 ( .A1(n7942), .A2(n8076), .ZN(n8165) );
  NAND2_X2 U5162 ( .A1(n8203), .A2(n9849), .ZN(n10957) );
  XNOR2_X1 U5163 ( .A(n6044), .B(n6040), .ZN(n7659) );
  NAND2_X1 U5164 ( .A1(n5312), .A2(n5316), .ZN(n6019) );
  NAND2_X1 U5165 ( .A1(n5894), .A2(n5893), .ZN(n8076) );
  INV_X2 U5166 ( .A(n10869), .ZN(n11027) );
  AND2_X1 U5167 ( .A1(n7221), .A2(n7220), .ZN(n5167) );
  NAND2_X2 U5168 ( .A1(n7696), .A2(n10865), .ZN(n10869) );
  INV_X1 U5169 ( .A(n8331), .ZN(n8241) );
  NAND2_X1 U5170 ( .A1(n6528), .A2(n6527), .ZN(n8331) );
  OAI211_X1 U5171 ( .C1(n7470), .C2(n7419), .A(n5826), .B(n5825), .ZN(n7930)
         );
  AND3_X1 U5172 ( .A1(n5779), .A2(n5778), .A3(n5777), .ZN(n10758) );
  NAND2_X1 U5173 ( .A1(n5561), .A2(n5174), .ZN(n7024) );
  NAND2_X1 U5174 ( .A1(n5175), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5174) );
  OAI211_X1 U5175 ( .C1(n7470), .C2(n7405), .A(n5744), .B(n5743), .ZN(n10738)
         );
  NAND4_X2 U5176 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), .ZN(n5704)
         );
  NAND2_X1 U5177 ( .A1(n5484), .A2(n6395), .ZN(n7497) );
  AND2_X1 U5178 ( .A1(n8696), .A2(n8709), .ZN(n5790) );
  INV_X2 U5179 ( .A(n5763), .ZN(n7005) );
  AND2_X1 U5180 ( .A1(n8696), .A2(n5650), .ZN(n5758) );
  NAND2_X2 U5181 ( .A1(n6416), .A2(n7264), .ZN(n7470) );
  INV_X1 U5182 ( .A(n8594), .ZN(n5032) );
  NAND2_X1 U5183 ( .A1(n5642), .A2(n5629), .ZN(n10535) );
  INV_X2 U5184 ( .A(n8294), .ZN(n5033) );
  NAND2_X1 U5185 ( .A1(n6921), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6456) );
  NAND2_X2 U5186 ( .A1(n5768), .A2(P1_U3084), .ZN(n9004) );
  NAND2_X2 U5187 ( .A1(n5671), .A2(n5670), .ZN(n5768) );
  NOR2_X1 U5188 ( .A1(n5587), .A2(n5056), .ZN(n5586) );
  AND2_X1 U5189 ( .A1(n5620), .A2(n6440), .ZN(n5229) );
  AND2_X1 U5190 ( .A1(n9591), .A2(n9799), .ZN(n5588) );
  AND2_X1 U5191 ( .A1(n5166), .A2(n5165), .ZN(n5636) );
  AND3_X1 U5192 ( .A1(n5663), .A2(n9797), .A3(n9796), .ZN(n5641) );
  AND2_X1 U5193 ( .A1(n6457), .A2(n5230), .ZN(n5619) );
  AND2_X1 U5194 ( .A1(n5234), .A2(n5235), .ZN(n5620) );
  INV_X1 U5195 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5663) );
  NOR2_X1 U5196 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5166) );
  NOR2_X1 U5197 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5323) );
  INV_X1 U5198 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10687) );
  NOR2_X1 U5199 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5165) );
  NOR2_X1 U5200 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5324) );
  INV_X1 U5201 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9591) );
  INV_X1 U5202 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9798) );
  INV_X1 U5203 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9799) );
  INV_X4 U5204 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5205 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9796) );
  INV_X1 U5206 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6471) );
  INV_X1 U5207 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6469) );
  INV_X1 U5208 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9558) );
  INV_X1 U5209 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5771) );
  INV_X1 U5210 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9785) );
  NAND2_X1 U5211 ( .A1(n6416), .A2(n7264), .ZN(n5034) );
  NAND2_X1 U5212 ( .A1(n6416), .A2(n7264), .ZN(n5035) );
  XNOR2_X2 U5213 ( .A(n6456), .B(n6455), .ZN(n7287) );
  NOR2_X4 U5214 ( .A1(n8165), .A2(n8475), .ZN(n8164) );
  OR2_X1 U5215 ( .A1(n9970), .A2(n9876), .ZN(n9837) );
  OR2_X1 U5216 ( .A1(n9960), .A2(n9842), .ZN(n8792) );
  NAND2_X1 U5217 ( .A1(n5614), .A2(n5213), .ZN(n5212) );
  AND2_X1 U5218 ( .A1(n8930), .A2(n8536), .ZN(n5615) );
  AND3_X1 U5219 ( .A1(n5362), .A2(n5361), .A3(n5360), .ZN(n6441) );
  INV_X1 U5220 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5362) );
  OR2_X1 U5221 ( .A1(n10461), .A2(n10305), .ZN(n7196) );
  INV_X1 U5222 ( .A(n5520), .ZN(n5184) );
  NAND2_X1 U5223 ( .A1(n5160), .A2(n5159), .ZN(n9838) );
  AOI21_X1 U5224 ( .B1(n5455), .B2(n5458), .A(n9860), .ZN(n5159) );
  NAND2_X1 U5225 ( .A1(n7306), .A2(n6995), .ZN(n6540) );
  OR2_X1 U5226 ( .A1(n8971), .A2(n8992), .ZN(n10268) );
  AOI21_X1 U5227 ( .B1(n7912), .B2(n5583), .A(n7911), .ZN(n5580) );
  INV_X1 U5228 ( .A(n7908), .ZN(n5583) );
  AND2_X1 U5229 ( .A1(n5531), .A2(n6045), .ZN(n5530) );
  INV_X1 U5230 ( .A(n6064), .ZN(n6045) );
  OR2_X1 U5231 ( .A1(n5533), .A2(n5532), .ZN(n5531) );
  XNOR2_X1 U5232 ( .A(n6906), .B(n8193), .ZN(n6497) );
  NAND2_X1 U5233 ( .A1(n5449), .A2(n6838), .ZN(n5448) );
  OR2_X1 U5234 ( .A1(n6826), .A2(n5451), .ZN(n5450) );
  INV_X1 U5235 ( .A(n6836), .ZN(n5449) );
  OR2_X1 U5236 ( .A1(n6898), .A2(n6897), .ZN(n6965) );
  OR2_X1 U5237 ( .A1(n9939), .A2(n9092), .ZN(n8888) );
  NAND2_X1 U5238 ( .A1(n6666), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6681) );
  NAND2_X1 U5239 ( .A1(n9893), .A2(n10817), .ZN(n8812) );
  AND2_X1 U5240 ( .A1(n5043), .A2(n5085), .ZN(n5514) );
  NOR2_X1 U5241 ( .A1(n5386), .A2(n8983), .ZN(n5385) );
  INV_X1 U5242 ( .A(n8980), .ZN(n5386) );
  NOR2_X1 U5243 ( .A1(n10358), .A2(n5383), .ZN(n5382) );
  INV_X1 U5244 ( .A(n8982), .ZN(n5383) );
  OR2_X1 U5245 ( .A1(n10481), .A2(n10371), .ZN(n8984) );
  NOR2_X1 U5246 ( .A1(n8581), .A2(n8583), .ZN(n5630) );
  NAND2_X1 U5247 ( .A1(n5053), .A2(n8584), .ZN(n5558) );
  NAND2_X1 U5248 ( .A1(n8171), .A2(n5063), .ZN(n5572) );
  NAND2_X1 U5249 ( .A1(n5572), .A2(n5570), .ZN(n8387) );
  NOR2_X1 U5250 ( .A1(n8176), .A2(n5571), .ZN(n5570) );
  INV_X1 U5251 ( .A(n5573), .ZN(n5571) );
  NAND2_X1 U5252 ( .A1(n8291), .A2(n10344), .ZN(n7110) );
  INV_X1 U5253 ( .A(n5588), .ZN(n5587) );
  NAND2_X1 U5254 ( .A1(n5130), .A2(n6051), .ZN(n6090) );
  INV_X1 U5255 ( .A(n6052), .ZN(n6051) );
  INV_X1 U5256 ( .A(n6053), .ZN(n5130) );
  NAND2_X1 U5257 ( .A1(n5958), .A2(n5985), .ZN(n5313) );
  XNOR2_X1 U5258 ( .A(n6041), .B(n6020), .ZN(n6040) );
  NAND2_X1 U5259 ( .A1(n5322), .A2(n5958), .ZN(n5321) );
  OR2_X1 U5260 ( .A1(n5866), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U5261 ( .A1(n5366), .A2(n5369), .ZN(n5886) );
  AOI21_X1 U5262 ( .B1(n5860), .B2(n5370), .A(n5078), .ZN(n5369) );
  NAND2_X1 U5263 ( .A1(n5259), .A2(n5258), .ZN(n8948) );
  NAND2_X1 U5264 ( .A1(n8913), .A2(n8914), .ZN(n5258) );
  INV_X1 U5265 ( .A(n6549), .ZN(n6969) );
  OR2_X1 U5266 ( .A1(n9936), .A2(n9258), .ZN(n9259) );
  NAND2_X1 U5267 ( .A1(n5228), .A2(n5589), .ZN(n5227) );
  INV_X1 U5268 ( .A(n5590), .ZN(n5589) );
  OR2_X1 U5269 ( .A1(n9391), .A2(n5090), .ZN(n8760) );
  NAND2_X1 U5270 ( .A1(n9859), .A2(n9876), .ZN(n5206) );
  NAND2_X1 U5271 ( .A1(n9854), .A2(n9860), .ZN(n5207) );
  NAND2_X1 U5272 ( .A1(n5461), .A2(n5460), .ZN(n5459) );
  INV_X1 U5273 ( .A(n5464), .ZN(n5460) );
  INV_X1 U5274 ( .A(n5462), .ZN(n5461) );
  AOI21_X1 U5275 ( .B1(n5210), .B2(n8636), .A(n5038), .ZN(n5208) );
  NAND2_X1 U5276 ( .A1(n5613), .A2(n5210), .ZN(n5209) );
  NOR2_X1 U5277 ( .A1(n10909), .A2(n8448), .ZN(n5222) );
  NAND2_X1 U5278 ( .A1(n8454), .A2(n5224), .ZN(n5223) );
  NAND2_X1 U5279 ( .A1(n10765), .A2(n8249), .ZN(n10801) );
  XNOR2_X1 U5280 ( .A(n6476), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6483) );
  AND2_X1 U5281 ( .A1(n6477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6481) );
  MUX2_X1 U5282 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6452), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5137) );
  XNOR2_X1 U5283 ( .A(n6468), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U5284 ( .A1(n5644), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5677) );
  INV_X1 U5285 ( .A(n7470), .ZN(n6142) );
  AOI21_X1 U5286 ( .B1(n5567), .B2(n5304), .A(n5075), .ZN(n5303) );
  AND2_X1 U5287 ( .A1(n7195), .A2(n8989), .ZN(n10306) );
  AND2_X1 U5288 ( .A1(n6358), .A2(n6357), .ZN(n10305) );
  INV_X1 U5289 ( .A(n10052), .ZN(n10323) );
  NAND2_X1 U5290 ( .A1(n5297), .A2(n5296), .ZN(n8966) );
  AND2_X1 U5291 ( .A1(n5298), .A2(n5094), .ZN(n5296) );
  OR2_X1 U5292 ( .A1(n10507), .A2(n10430), .ZN(n8975) );
  INV_X1 U5293 ( .A(n8973), .ZN(n8630) );
  NAND2_X1 U5294 ( .A1(n7802), .A2(n5584), .ZN(n7909) );
  NAND2_X2 U5295 ( .A1(n5034), .A2(n6995), .ZN(n7015) );
  NAND2_X1 U5296 ( .A1(n7011), .A2(SI_29_), .ZN(n7014) );
  NAND2_X1 U5297 ( .A1(n6488), .A2(n9846), .ZN(n8955) );
  XNOR2_X1 U5298 ( .A(n5205), .B(n5128), .ZN(n5204) );
  NAND2_X1 U5299 ( .A1(n9231), .A2(n5129), .ZN(n5205) );
  NAND2_X1 U5300 ( .A1(n10268), .A2(n8972), .ZN(n10459) );
  OAI21_X1 U5301 ( .B1(n5255), .B2(n5254), .A(n5252), .ZN(n8827) );
  NOR2_X1 U5302 ( .A1(n5253), .A2(n5225), .ZN(n5252) );
  NAND2_X1 U5303 ( .A1(n8819), .A2(n8925), .ZN(n5254) );
  AOI21_X1 U5304 ( .B1(n8810), .B2(n8812), .A(n5256), .ZN(n5255) );
  INV_X1 U5305 ( .A(n8853), .ZN(n5250) );
  AND2_X1 U5306 ( .A1(n5249), .A2(n5095), .ZN(n5248) );
  OR2_X1 U5307 ( .A1(n5251), .A2(n8840), .ZN(n5249) );
  NAND2_X1 U5308 ( .A1(n5274), .A2(n9250), .ZN(n5273) );
  INV_X1 U5309 ( .A(n8868), .ZN(n5274) );
  AND2_X1 U5310 ( .A1(n5277), .A2(n5269), .ZN(n5268) );
  NAND2_X1 U5311 ( .A1(n5271), .A2(n5270), .ZN(n5269) );
  AND2_X1 U5312 ( .A1(n9839), .A2(n8870), .ZN(n5277) );
  INV_X1 U5313 ( .A(n5275), .ZN(n5270) );
  NOR2_X1 U5314 ( .A1(n5244), .A2(n8938), .ZN(n5239) );
  NAND2_X1 U5315 ( .A1(n8885), .A2(n9346), .ZN(n5245) );
  AND2_X1 U5316 ( .A1(n8895), .A2(n8894), .ZN(n8898) );
  NAND2_X1 U5317 ( .A1(n5546), .A2(n5068), .ZN(n5545) );
  INV_X1 U5318 ( .A(n8909), .ZN(n5263) );
  OR2_X1 U5319 ( .A1(n9244), .A2(n9271), .ZN(n8911) );
  INV_X1 U5320 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6450) );
  NOR2_X1 U5321 ( .A1(n5541), .A2(n5537), .ZN(n5536) );
  INV_X1 U5322 ( .A(n6194), .ZN(n5537) );
  OAI21_X1 U5323 ( .B1(n5541), .B2(n5542), .A(n6267), .ZN(n5540) );
  INV_X1 U5324 ( .A(n6042), .ZN(n5532) );
  INV_X1 U5325 ( .A(n5317), .ZN(n5316) );
  OAI21_X1 U5326 ( .B1(n5319), .B2(n5318), .A(n5633), .ZN(n5317) );
  NAND2_X1 U5327 ( .A1(n5912), .A2(n9644), .ZN(n5936) );
  NAND2_X1 U5328 ( .A1(n5889), .A2(n9448), .ZN(n5909) );
  OAI21_X1 U5329 ( .B1(n5157), .B2(n5154), .A(n5158), .ZN(n5153) );
  NAND2_X1 U5330 ( .A1(n9241), .A2(n8947), .ZN(n5158) );
  NAND2_X1 U5331 ( .A1(n8911), .A2(n5155), .ZN(n5154) );
  INV_X1 U5332 ( .A(n8907), .ZN(n5155) );
  NAND2_X1 U5333 ( .A1(n8908), .A2(n8911), .ZN(n5156) );
  OR2_X1 U5334 ( .A1(n9919), .A2(n9309), .ZN(n8904) );
  AND2_X1 U5335 ( .A1(n5599), .A2(n9307), .ZN(n5598) );
  NAND2_X1 U5336 ( .A1(n5600), .A2(n9261), .ZN(n5599) );
  INV_X1 U5337 ( .A(n9319), .ZN(n5600) );
  INV_X1 U5338 ( .A(n8896), .ZN(n5147) );
  OR2_X1 U5339 ( .A1(n9924), .A2(n9262), .ZN(n8901) );
  INV_X1 U5340 ( .A(n9349), .ZN(n5593) );
  OR2_X1 U5341 ( .A1(n6811), .A2(n9113), .ZN(n6828) );
  OR2_X1 U5342 ( .A1(n6799), .A2(n9681), .ZN(n6811) );
  NOR2_X1 U5343 ( .A1(n9960), .A2(n9967), .ZN(n5359) );
  NAND2_X1 U5344 ( .A1(n9869), .A2(n5608), .ZN(n5607) );
  INV_X1 U5345 ( .A(n5626), .ZN(n5608) );
  OR2_X1 U5346 ( .A1(n8735), .A2(n8670), .ZN(n8860) );
  OR2_X1 U5347 ( .A1(n8535), .A2(n5352), .ZN(n5351) );
  OR2_X1 U5348 ( .A1(n6652), .A2(n7866), .ZN(n6667) );
  AND2_X1 U5349 ( .A1(n8255), .A2(n5225), .ZN(n5224) );
  OR2_X1 U5350 ( .A1(n10938), .A2(n8423), .ZN(n8828) );
  INV_X1 U5351 ( .A(n8811), .ZN(n5472) );
  NAND2_X1 U5352 ( .A1(n9838), .A2(n8757), .ZN(n5161) );
  OR2_X1 U5353 ( .A1(n9893), .A2(n10804), .ZN(n5216) );
  NAND2_X1 U5354 ( .A1(n8193), .A2(n7959), .ZN(n8204) );
  NOR2_X1 U5355 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6440) );
  NOR2_X1 U5356 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5230) );
  NOR2_X1 U5357 ( .A1(n6108), .A2(n5517), .ZN(n5516) );
  NOR2_X1 U5358 ( .A1(n10125), .A2(n5512), .ZN(n5510) );
  INV_X1 U5359 ( .A(n10125), .ZN(n5508) );
  AND2_X1 U5360 ( .A1(n5491), .A2(n6039), .ZN(n5490) );
  NAND2_X1 U5361 ( .A1(n10337), .A2(n5304), .ZN(n5390) );
  OR2_X1 U5362 ( .A1(n6300), .A2(n6299), .ZN(n6332) );
  OR2_X1 U5363 ( .A1(n10493), .A2(n10402), .ZN(n8980) );
  OR2_X1 U5364 ( .A1(n10496), .A2(n10431), .ZN(n8978) );
  OR2_X1 U5365 ( .A1(n10514), .A2(n8626), .ZN(n8617) );
  NOR2_X1 U5366 ( .A1(n8385), .A2(n8094), .ZN(n5340) );
  NAND2_X1 U5367 ( .A1(n10965), .A2(n8309), .ZN(n5573) );
  NAND2_X1 U5368 ( .A1(n8158), .A2(n8078), .ZN(n8171) );
  INV_X1 U5369 ( .A(n7904), .ZN(n5180) );
  AND2_X1 U5370 ( .A1(n10848), .A2(n10844), .ZN(n7903) );
  NOR2_X1 U5371 ( .A1(n7806), .A2(n5585), .ZN(n5584) );
  INV_X1 U5372 ( .A(n7801), .ZN(n5585) );
  NAND2_X1 U5373 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  OAI21_X1 U5374 ( .B1(n6987), .B2(n6986), .A(n6985), .ZN(n6990) );
  OAI21_X1 U5375 ( .B1(n6293), .B2(n6292), .A(n6291), .ZN(n6318) );
  OAI21_X1 U5376 ( .B1(n6168), .B2(n6167), .A(n6166), .ZN(n6193) );
  AND2_X1 U5377 ( .A1(n6194), .A2(n6171), .ZN(n6192) );
  NOR2_X1 U5378 ( .A1(n5553), .A2(n5552), .ZN(n5551) );
  NOR2_X1 U5379 ( .A1(n6043), .A2(n5534), .ZN(n5533) );
  NOR2_X1 U5380 ( .A1(n5534), .A2(n5318), .ZN(n5314) );
  NOR2_X1 U5381 ( .A1(n5986), .A2(n5320), .ZN(n5319) );
  INV_X1 U5382 ( .A(n5961), .ZN(n5320) );
  INV_X1 U5383 ( .A(SI_11_), .ZN(n5938) );
  INV_X1 U5384 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9570) );
  OAI21_X1 U5385 ( .B1(n5886), .B2(n5292), .A(n5290), .ZN(n5915) );
  INV_X1 U5386 ( .A(n5293), .ZN(n5292) );
  AOI21_X1 U5387 ( .B1(n5884), .B2(n5293), .A(n5291), .ZN(n5290) );
  AND2_X1 U5388 ( .A1(n5294), .A2(n5888), .ZN(n5293) );
  OR3_X1 U5389 ( .A1(n5863), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        P1_IR_REG_7__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U5390 ( .A1(n5741), .A2(n5799), .ZN(n5281) );
  OAI21_X1 U5391 ( .B1(n5768), .B2(n5287), .A(n5286), .ZN(n5766) );
  NAND2_X1 U5392 ( .A1(n5768), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5286) );
  INV_X1 U5393 ( .A(n7999), .ZN(n5397) );
  AOI21_X1 U5394 ( .B1(n7948), .B2(n6599), .A(n5127), .ZN(n5398) );
  INV_X1 U5395 ( .A(n10707), .ZN(n7959) );
  OR2_X1 U5396 ( .A1(n8000), .A2(n7999), .ZN(n8045) );
  NAND2_X1 U5397 ( .A1(n6511), .A2(n6510), .ZN(n6512) );
  INV_X1 U5398 ( .A(n5424), .ZN(n5423) );
  NAND2_X1 U5399 ( .A1(n5424), .A2(n5422), .ZN(n5421) );
  NOR2_X1 U5400 ( .A1(n9088), .A2(n5425), .ZN(n5424) );
  INV_X1 U5401 ( .A(n6735), .ZN(n5425) );
  INV_X1 U5402 ( .A(n6548), .ZN(n5412) );
  INV_X1 U5403 ( .A(n6864), .ZN(n5443) );
  AND2_X1 U5404 ( .A1(n6947), .A2(n8947), .ZN(n7285) );
  NAND2_X1 U5405 ( .A1(n7830), .A2(n8947), .ZN(n8779) );
  OAI21_X1 U5406 ( .B1(n6467), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6914) );
  OR2_X1 U5407 ( .A1(n7344), .A2(n7343), .ZN(n5195) );
  OR2_X1 U5408 ( .A1(n7332), .A2(n7331), .ZN(n5201) );
  AND2_X1 U5409 ( .A1(n6899), .A2(n6965), .ZN(n9286) );
  INV_X1 U5410 ( .A(n9265), .ZN(n9290) );
  OR2_X1 U5411 ( .A1(n9306), .A2(n9307), .ZN(n9311) );
  NAND2_X1 U5412 ( .A1(n8918), .A2(n8917), .ZN(n9319) );
  NAND2_X1 U5413 ( .A1(n6841), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6852) );
  INV_X1 U5414 ( .A(n9257), .ZN(n9331) );
  AOI21_X1 U5415 ( .B1(n9334), .B2(n6550), .A(n6847), .ZN(n9350) );
  NAND2_X1 U5416 ( .A1(n5594), .A2(n5592), .ZN(n9339) );
  OR2_X1 U5417 ( .A1(n9950), .A2(n9065), .ZN(n8881) );
  AND2_X1 U5418 ( .A1(n8882), .A2(n9346), .ZN(n9360) );
  NAND2_X1 U5419 ( .A1(n8760), .A2(n5478), .ZN(n9380) );
  AND2_X1 U5420 ( .A1(n9254), .A2(n8759), .ZN(n5478) );
  AND2_X1 U5421 ( .A1(n6835), .A2(n6834), .ZN(n9378) );
  NOR2_X1 U5422 ( .A1(n9390), .A2(n9252), .ZN(n5612) );
  NAND2_X1 U5423 ( .A1(n9834), .A2(n5106), .ZN(n9399) );
  NAND2_X1 U5424 ( .A1(n9399), .A2(n9406), .ZN(n9398) );
  AND3_X1 U5425 ( .A1(n6791), .A2(n6790), .A3(n6789), .ZN(n9842) );
  AOI21_X1 U5426 ( .B1(n5457), .B2(n5462), .A(n5071), .ZN(n5455) );
  OAI21_X1 U5427 ( .B1(n8755), .B2(n5463), .A(n8864), .ZN(n5462) );
  NAND2_X1 U5428 ( .A1(n8679), .A2(n8859), .ZN(n5463) );
  NOR2_X1 U5429 ( .A1(n8755), .A2(n5465), .ZN(n5464) );
  INV_X1 U5430 ( .A(n8859), .ZN(n5465) );
  INV_X1 U5431 ( .A(n5607), .ZN(n5605) );
  INV_X1 U5432 ( .A(n9249), .ZN(n5606) );
  AND2_X1 U5433 ( .A1(n9250), .A2(n8867), .ZN(n9869) );
  AND2_X1 U5434 ( .A1(n8864), .A2(n8863), .ZN(n8935) );
  NOR2_X1 U5435 ( .A1(n8677), .A2(n8935), .ZN(n9249) );
  AND2_X1 U5436 ( .A1(n8860), .A2(n8859), .ZN(n8934) );
  NAND2_X1 U5437 ( .A1(n6680), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6695) );
  AOI21_X1 U5438 ( .B1(n5615), .B2(n8844), .A(n5086), .ZN(n5614) );
  OR2_X1 U5439 ( .A1(n5214), .A2(n5212), .ZN(n5211) );
  INV_X1 U5440 ( .A(n5613), .ZN(n5214) );
  NAND2_X1 U5441 ( .A1(n5132), .A2(n5133), .ZN(n5131) );
  NAND2_X1 U5442 ( .A1(n5467), .A2(n8544), .ZN(n5132) );
  NAND2_X1 U5443 ( .A1(n5354), .A2(n5353), .ZN(n5352) );
  NOR2_X1 U5444 ( .A1(n10933), .A2(n5351), .ZN(n8569) );
  NOR2_X1 U5445 ( .A1(n8925), .A2(n5618), .ZN(n5617) );
  INV_X1 U5446 ( .A(n8254), .ZN(n5618) );
  NAND2_X1 U5447 ( .A1(n9888), .A2(n8818), .ZN(n5142) );
  XNOR2_X1 U5448 ( .A(n9891), .B(n10873), .ZN(n8925) );
  NAND2_X1 U5449 ( .A1(n8248), .A2(n8247), .ZN(n8811) );
  AND2_X1 U5450 ( .A1(n8815), .A2(n8812), .ZN(n10808) );
  OAI211_X1 U5451 ( .C1(n6540), .C2(n7417), .A(n6543), .B(n5074), .ZN(n10769)
         );
  OR2_X1 U5452 ( .A1(n10773), .A2(n8258), .ZN(n10775) );
  NAND2_X1 U5453 ( .A1(n9161), .A2(n10707), .ZN(n8191) );
  AND2_X1 U5454 ( .A1(n7285), .A2(n6975), .ZN(n9890) );
  INV_X1 U5455 ( .A(n11070), .ZN(n10892) );
  NOR2_X1 U5456 ( .A1(n7821), .A2(n7820), .ZN(n7835) );
  NAND2_X1 U5457 ( .A1(n10945), .A2(n7826), .ZN(n11074) );
  INV_X1 U5458 ( .A(n5407), .ZN(n5406) );
  OAI21_X1 U5459 ( .B1(n6466), .B2(n10002), .A(n6469), .ZN(n5407) );
  NOR3_X1 U5460 ( .A1(n6662), .A2(P2_IR_REG_12__SCAN_IN), .A3(n6460), .ZN(
        n6721) );
  INV_X1 U5461 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U5462 ( .A1(n5842), .A2(n5841), .ZN(n7910) );
  AOI21_X1 U5463 ( .B1(n5044), .B2(n5502), .A(n5082), .ZN(n5500) );
  NAND2_X1 U5464 ( .A1(n10038), .A2(n10036), .ZN(n5496) );
  NAND2_X1 U5465 ( .A1(n5498), .A2(n6211), .ZN(n10040) );
  INV_X1 U5466 ( .A(n10037), .ZN(n5498) );
  INV_X1 U5467 ( .A(n6087), .ZN(n5519) );
  NAND2_X1 U5468 ( .A1(n10084), .A2(n10085), .ZN(n10083) );
  OR2_X1 U5469 ( .A1(n6430), .A2(n7577), .ZN(n6426) );
  OAI22_X1 U5470 ( .A1(n7112), .A2(n7111), .B1(n7142), .B2(n7110), .ZN(n7116)
         );
  AND2_X1 U5471 ( .A1(n6393), .A2(n5032), .ZN(n5484) );
  NOR2_X1 U5472 ( .A1(n10288), .A2(n10455), .ZN(n10256) );
  NAND2_X1 U5473 ( .A1(n8970), .A2(n8969), .ZN(n8971) );
  AND2_X1 U5474 ( .A1(n10296), .A2(n5303), .ZN(n5301) );
  NAND2_X1 U5475 ( .A1(n10311), .A2(n10293), .ZN(n10288) );
  OR2_X1 U5476 ( .A1(n10318), .A2(n5568), .ZN(n5302) );
  NAND2_X1 U5477 ( .A1(n5390), .A2(n5388), .ZN(n10303) );
  NOR2_X1 U5478 ( .A1(n5391), .A2(n5389), .ZN(n5388) );
  INV_X1 U5479 ( .A(n10306), .ZN(n5389) );
  NOR2_X1 U5480 ( .A1(n5387), .A2(n5391), .ZN(n10304) );
  INV_X1 U5481 ( .A(n5390), .ZN(n5387) );
  NOR2_X1 U5482 ( .A1(n10337), .A2(n8987), .ZN(n10322) );
  OAI21_X1 U5483 ( .B1(n8981), .B2(n5381), .A(n5379), .ZN(n5378) );
  AOI21_X1 U5484 ( .B1(n5382), .B2(n5380), .A(n8985), .ZN(n5379) );
  INV_X1 U5485 ( .A(n5382), .ZN(n5381) );
  AOI21_X1 U5486 ( .B1(n8964), .B2(n5299), .A(n5073), .ZN(n5298) );
  INV_X1 U5487 ( .A(n8963), .ZN(n5299) );
  OR2_X1 U5488 ( .A1(n10367), .A2(n5300), .ZN(n5297) );
  INV_X1 U5489 ( .A(n8964), .ZN(n5300) );
  NAND2_X1 U5490 ( .A1(n8981), .A2(n5385), .ZN(n5384) );
  AND2_X1 U5491 ( .A1(n5384), .A2(n5382), .ZN(n10356) );
  INV_X1 U5492 ( .A(n10485), .ZN(n10375) );
  NAND2_X1 U5493 ( .A1(n5563), .A2(n5565), .ZN(n10365) );
  AOI21_X1 U5494 ( .B1(n10385), .B2(n5566), .A(n5070), .ZN(n5565) );
  INV_X1 U5495 ( .A(n6176), .ZN(n6174) );
  NAND2_X1 U5496 ( .A1(n10404), .A2(n10403), .ZN(n10405) );
  AND2_X1 U5497 ( .A1(n8975), .A2(n7175), .ZN(n8973) );
  OAI21_X1 U5498 ( .B1(n10999), .B2(n5081), .A(n5556), .ZN(n8600) );
  NAND2_X1 U5499 ( .A1(n5558), .A2(n8598), .ZN(n5556) );
  NAND2_X1 U5500 ( .A1(n8600), .A2(n8607), .ZN(n8629) );
  AND2_X1 U5501 ( .A1(n6127), .A2(n6126), .ZN(n10430) );
  NAND2_X1 U5502 ( .A1(n8602), .A2(n8601), .ZN(n5176) );
  NAND2_X1 U5503 ( .A1(n5560), .A2(n5630), .ZN(n5559) );
  INV_X1 U5504 ( .A(n10999), .ZN(n5560) );
  INV_X1 U5505 ( .A(n5558), .ZN(n5557) );
  NAND2_X1 U5506 ( .A1(n7765), .A2(n7764), .ZN(n7802) );
  NAND2_X1 U5507 ( .A1(n7633), .A2(n7271), .ZN(n10849) );
  AND2_X1 U5508 ( .A1(n7216), .A2(n7724), .ZN(n7742) );
  NAND2_X1 U5509 ( .A1(n5331), .A2(n7404), .ZN(n5330) );
  INV_X1 U5510 ( .A(n7431), .ZN(n5331) );
  NAND2_X1 U5511 ( .A1(n5036), .A2(n7271), .ZN(n10851) );
  AND2_X1 U5512 ( .A1(n5869), .A2(n5868), .ZN(n10882) );
  AND2_X1 U5513 ( .A1(n5183), .A2(n5586), .ZN(n5185) );
  INV_X1 U5514 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9808) );
  NAND2_X1 U5515 ( .A1(n10535), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5643) );
  AND2_X1 U5516 ( .A1(n5648), .A2(n10535), .ZN(n5649) );
  OAI21_X1 U5517 ( .B1(n5676), .B2(n5647), .A(n5646), .ZN(n5648) );
  NAND2_X1 U5518 ( .A1(n9813), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U5519 ( .A1(n5625), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5647) );
  XNOR2_X1 U5520 ( .A(n6990), .B(n6988), .ZN(n7011) );
  XNOR2_X1 U5521 ( .A(n6987), .B(n6986), .ZN(n9002) );
  XNOR2_X1 U5522 ( .A(n6365), .B(n6366), .ZN(n8690) );
  NAND2_X1 U5523 ( .A1(n5656), .A2(n9798), .ZN(n5660) );
  OAI21_X1 U5524 ( .B1(n6220), .B2(n6219), .A(n6218), .ZN(n6243) );
  XNOR2_X1 U5525 ( .A(n5680), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U5526 ( .A1(n6090), .A2(n6089), .ZN(n6110) );
  NAND2_X1 U5527 ( .A1(n5283), .A2(n5741), .ZN(n5765) );
  NAND2_X1 U5528 ( .A1(n6694), .A2(n6693), .ZN(n11051) );
  NAND2_X1 U5529 ( .A1(n6798), .A2(n6797), .ZN(n9955) );
  INV_X1 U5530 ( .A(n8687), .ZN(n9982) );
  NAND2_X1 U5531 ( .A1(n6849), .A2(n6848), .ZN(n9939) );
  AND4_X1 U5532 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n8448)
         );
  INV_X1 U5533 ( .A(n5435), .ZN(n5434) );
  AOI21_X1 U5534 ( .B1(n5435), .B2(n5433), .A(n5432), .ZN(n5431) );
  NAND2_X1 U5535 ( .A1(n5525), .A2(n5524), .ZN(n5523) );
  INV_X1 U5536 ( .A(n9092), .ZN(n9357) );
  INV_X1 U5537 ( .A(n9065), .ZN(n9393) );
  AND4_X1 U5538 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n9876)
         );
  INV_X1 U5539 ( .A(n8449), .ZN(n9157) );
  NOR2_X1 U5540 ( .A1(n10676), .A2(n10675), .ZN(n10674) );
  AND2_X1 U5541 ( .A1(n5195), .A2(n5194), .ZN(n7355) );
  NAND2_X1 U5542 ( .A1(n7293), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5194) );
  AND2_X1 U5543 ( .A1(n5197), .A2(n5196), .ZN(n7392) );
  NAND2_X1 U5544 ( .A1(n7394), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U5545 ( .A1(n10684), .A2(n10902), .ZN(n5203) );
  NAND2_X1 U5546 ( .A1(n7303), .A2(n7302), .ZN(n10677) );
  AND2_X1 U5547 ( .A1(n8767), .A2(n8766), .ZN(n9279) );
  OR2_X1 U5548 ( .A1(n8764), .A2(n6540), .ZN(n8767) );
  NAND2_X1 U5549 ( .A1(n5058), .A2(n5479), .ZN(n9050) );
  NAND2_X1 U5550 ( .A1(n7306), .A2(n5480), .ZN(n5479) );
  OAI21_X1 U5551 ( .B1(n7431), .B2(n7404), .A(n5481), .ZN(n5480) );
  NAND2_X1 U5552 ( .A1(n5405), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6470) );
  AND2_X1 U5553 ( .A1(n6282), .A2(n6281), .ZN(n10359) );
  INV_X1 U5554 ( .A(n11084), .ZN(n10069) );
  AND2_X1 U5555 ( .A1(n6258), .A2(n6257), .ZN(n10371) );
  XNOR2_X1 U5556 ( .A(n5682), .B(P1_IR_REG_22__SCAN_IN), .ZN(n7716) );
  OR2_X1 U5557 ( .A1(n10127), .A2(n6334), .ZN(n6340) );
  OR2_X1 U5558 ( .A1(n8764), .A2(n5763), .ZN(n7017) );
  AOI21_X1 U5559 ( .B1(n8995), .B2(n11009), .A(n5188), .ZN(n10458) );
  OAI21_X1 U5560 ( .B1(n10459), .B2(n11013), .A(n5189), .ZN(n5188) );
  INV_X1 U5561 ( .A(n8994), .ZN(n5189) );
  NAND2_X1 U5562 ( .A1(n5569), .A2(n8967), .ZN(n10307) );
  NAND2_X1 U5563 ( .A1(n10318), .A2(n10321), .ZN(n5569) );
  NAND2_X1 U5564 ( .A1(n10509), .A2(n8960), .ZN(n10423) );
  INV_X1 U5565 ( .A(n10392), .ZN(n10344) );
  NAND2_X1 U5566 ( .A1(n5372), .A2(n5309), .ZN(n5375) );
  INV_X1 U5567 ( .A(n5310), .ZN(n5309) );
  NAND2_X1 U5568 ( .A1(n5373), .A2(n11089), .ZN(n5372) );
  OAI21_X1 U5569 ( .B1(n5326), .B2(n11085), .A(n5325), .ZN(n5310) );
  INV_X1 U5570 ( .A(n8823), .ZN(n5253) );
  AOI21_X1 U5571 ( .B1(n8868), .B2(n8867), .A(n5276), .ZN(n5275) );
  INV_X1 U5572 ( .A(n8865), .ZN(n5276) );
  AOI21_X1 U5573 ( .B1(n5248), .B2(n5251), .A(n5088), .ZN(n5247) );
  AND2_X1 U5574 ( .A1(n5064), .A2(n5267), .ZN(n5266) );
  NAND2_X1 U5575 ( .A1(n5268), .A2(n5272), .ZN(n5267) );
  NOR2_X1 U5576 ( .A1(n5244), .A2(n5243), .ZN(n5242) );
  INV_X1 U5577 ( .A(n8878), .ZN(n5243) );
  INV_X1 U5578 ( .A(n5238), .ZN(n5237) );
  OAI21_X1 U5579 ( .B1(n5239), .B2(n5245), .A(n8886), .ZN(n5238) );
  INV_X1 U5580 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9764) );
  INV_X1 U5581 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U5582 ( .A1(n7748), .A2(n5111), .ZN(n7121) );
  AOI21_X1 U5583 ( .B1(n8899), .B2(n5061), .A(n9307), .ZN(n5547) );
  NAND2_X1 U5584 ( .A1(n5550), .A2(n5549), .ZN(n5548) );
  NOR2_X1 U5585 ( .A1(n5148), .A2(n8912), .ZN(n5549) );
  OAI21_X1 U5586 ( .B1(n8898), .B2(n5257), .A(n8896), .ZN(n5550) );
  INV_X1 U5587 ( .A(n8897), .ZN(n5257) );
  INV_X1 U5588 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9742) );
  INV_X1 U5589 ( .A(SI_9_), .ZN(n9448) );
  INV_X1 U5590 ( .A(n9018), .ZN(n5451) );
  INV_X1 U5591 ( .A(n8912), .ZN(n8906) );
  OR2_X1 U5592 ( .A1(n8818), .A2(n5144), .ZN(n5143) );
  NAND2_X1 U5593 ( .A1(n6139), .A2(n9631), .ZN(n6166) );
  INV_X1 U5594 ( .A(n6089), .ZN(n5552) );
  INV_X1 U5595 ( .A(n5910), .ZN(n5294) );
  INV_X1 U5596 ( .A(n5909), .ZN(n5291) );
  INV_X1 U5597 ( .A(n5838), .ZN(n5370) );
  INV_X1 U5598 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5668) );
  INV_X1 U5599 ( .A(n6906), .ZN(n6907) );
  NAND2_X1 U5600 ( .A1(n5264), .A2(n5261), .ZN(n5260) );
  NOR2_X1 U5601 ( .A1(n5263), .A2(n5262), .ZN(n5261) );
  NAND2_X1 U5602 ( .A1(n8911), .A2(n8910), .ZN(n5262) );
  MUX2_X1 U5603 ( .A(n8787), .B(n8944), .S(n8906), .Z(n8915) );
  OAI21_X1 U5604 ( .B1(n5592), .B2(n5591), .A(n9257), .ZN(n5590) );
  OR2_X1 U5605 ( .A1(n9945), .A2(n9378), .ZN(n8882) );
  INV_X1 U5606 ( .A(n6787), .ZN(n6786) );
  AOI21_X1 U5607 ( .B1(n5212), .B2(n8635), .A(n8934), .ZN(n5210) );
  INV_X1 U5608 ( .A(n8846), .ZN(n5136) );
  INV_X1 U5609 ( .A(n5224), .ZN(n5218) );
  NOR2_X1 U5610 ( .A1(n8926), .A2(n5222), .ZN(n5221) );
  AND2_X1 U5611 ( .A1(n5143), .A2(n8925), .ZN(n5139) );
  NOR2_X1 U5612 ( .A1(n8201), .A2(n9846), .ZN(n8786) );
  NAND2_X1 U5613 ( .A1(n8193), .A2(n9159), .ZN(n8209) );
  INV_X1 U5614 ( .A(n9279), .ZN(n9918) );
  NAND2_X1 U5615 ( .A1(n9855), .A2(n9843), .ZN(n9845) );
  NOR2_X1 U5616 ( .A1(n8683), .A2(n9982), .ZN(n9877) );
  NAND2_X1 U5617 ( .A1(n8417), .A2(n5134), .ZN(n10935) );
  NOR2_X1 U5618 ( .A1(n10931), .A2(n5135), .ZN(n5134) );
  INV_X1 U5619 ( .A(n8828), .ZN(n5135) );
  NAND2_X1 U5620 ( .A1(n8190), .A2(n8189), .ZN(n8323) );
  AOI221_X1 U5621 ( .B1(P2_B_REG_SCAN_IN), .B2(n6928), .C1(n6927), .C2(n8462), 
        .A(n6944), .ZN(n6931) );
  INV_X1 U5622 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6478) );
  INV_X1 U5623 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5621) );
  AND2_X1 U5624 ( .A1(n5164), .A2(n6455), .ZN(n5163) );
  AND2_X1 U5625 ( .A1(n6449), .A2(n6441), .ZN(n5475) );
  INV_X1 U5626 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5164) );
  INV_X1 U5627 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5234) );
  INV_X1 U5628 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5235) );
  NOR2_X1 U5629 ( .A1(n5041), .A2(n5488), .ZN(n5487) );
  NAND2_X1 U5630 ( .A1(n5665), .A2(n7497), .ZN(n5688) );
  INV_X1 U5631 ( .A(n5503), .ZN(n5505) );
  INV_X1 U5632 ( .A(n5957), .ZN(n5502) );
  OR2_X1 U5633 ( .A1(n8223), .A2(n5502), .ZN(n5501) );
  NAND2_X1 U5634 ( .A1(n10283), .A2(n10157), .ZN(n7212) );
  NAND2_X1 U5635 ( .A1(n10255), .A2(n8993), .ZN(n7250) );
  OR2_X1 U5636 ( .A1(n10455), .A2(n10297), .ZN(n7211) );
  INV_X1 U5637 ( .A(n5385), .ZN(n5380) );
  NOR2_X1 U5638 ( .A1(n10375), .A2(n5335), .ZN(n5334) );
  INV_X1 U5639 ( .A(n5336), .ZN(n5335) );
  NOR2_X1 U5640 ( .A1(n10493), .A2(n10496), .ZN(n5336) );
  NOR2_X1 U5641 ( .A1(n10388), .A2(n10399), .ZN(n5564) );
  INV_X1 U5642 ( .A(n8962), .ZN(n5566) );
  OR2_X1 U5643 ( .A1(n8524), .A2(n11007), .ZN(n8581) );
  OR2_X1 U5644 ( .A1(n10135), .A2(n10067), .ZN(n8576) );
  NAND2_X1 U5645 ( .A1(n8387), .A2(n8386), .ZN(n10999) );
  OR2_X1 U5646 ( .A1(n8087), .A2(n5172), .ZN(n5170) );
  INV_X1 U5647 ( .A(n8174), .ZN(n5172) );
  AOI21_X1 U5648 ( .B1(n7802), .B2(n5581), .A(n5579), .ZN(n7933) );
  NOR2_X1 U5649 ( .A1(n10848), .A2(n5582), .ZN(n5581) );
  INV_X1 U5650 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5843) );
  NOR2_X1 U5651 ( .A1(n5844), .A2(n5843), .ZN(n5870) );
  NAND2_X1 U5652 ( .A1(n10433), .A2(n10414), .ZN(n10416) );
  NAND2_X1 U5653 ( .A1(n7014), .A2(n6991), .ZN(n7002) );
  NAND2_X1 U5654 ( .A1(n5535), .A2(n5539), .ZN(n6270) );
  INV_X1 U5655 ( .A(n5540), .ZN(n5539) );
  NAND2_X1 U5656 ( .A1(n5544), .A2(n6218), .ZN(n5543) );
  INV_X1 U5657 ( .A(n6242), .ZN(n5544) );
  NAND2_X1 U5658 ( .A1(n6193), .A2(n6192), .ZN(n6195) );
  NAND2_X1 U5659 ( .A1(n6048), .A2(n9439), .ZN(n6089) );
  AOI21_X1 U5660 ( .B1(n5530), .B2(n5532), .A(n5076), .ZN(n5527) );
  NAND2_X1 U5661 ( .A1(n5288), .A2(n5669), .ZN(n5670) );
  INV_X1 U5662 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U5663 ( .A1(n5667), .A2(n5668), .ZN(n5288) );
  INV_X1 U5664 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U5665 ( .A1(n5289), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U5666 ( .A1(n10687), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U5667 ( .A1(n5444), .A2(n5057), .ZN(n9072) );
  NAND2_X1 U5668 ( .A1(n5446), .A2(n5445), .ZN(n5444) );
  INV_X1 U5669 ( .A(n9109), .ZN(n5446) );
  NAND2_X1 U5670 ( .A1(n5438), .A2(n5437), .ZN(n9026) );
  INV_X1 U5671 ( .A(n6780), .ZN(n5437) );
  INV_X1 U5672 ( .A(n9027), .ZN(n5438) );
  INV_X1 U5673 ( .A(n9028), .ZN(n5433) );
  INV_X1 U5674 ( .A(n6796), .ZN(n5432) );
  AND2_X1 U5675 ( .A1(n9103), .A2(n5436), .ZN(n5435) );
  NAND2_X1 U5676 ( .A1(n6780), .A2(n9028), .ZN(n5436) );
  INV_X1 U5677 ( .A(n8191), .ZN(n5429) );
  AND2_X1 U5678 ( .A1(n8743), .A2(n5418), .ZN(n5417) );
  OR2_X1 U5679 ( .A1(n8715), .A2(n5039), .ZN(n5418) );
  INV_X1 U5680 ( .A(n5153), .ZN(n5152) );
  AND4_X1 U5681 ( .A1(n8787), .A2(n8944), .A3(n9267), .A4(n5628), .ZN(n8945)
         );
  XNOR2_X1 U5682 ( .A(n8951), .B(n5526), .ZN(n5525) );
  INV_X1 U5683 ( .A(n8950), .ZN(n5526) );
  NOR2_X1 U5684 ( .A1(n10706), .A2(n7830), .ZN(n5524) );
  AND3_X1 U5685 ( .A1(n8771), .A2(n8770), .A3(n8769), .ZN(n9241) );
  AND4_X1 U5686 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n8418)
         );
  AND4_X1 U5687 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n10938)
         );
  AND4_X1 U5688 ( .A1(n6520), .A2(n6519), .A3(n6518), .A4(n6517), .ZN(n8240)
         );
  OR2_X1 U5689 ( .A1(n7318), .A2(n7317), .ZN(n5199) );
  OR2_X1 U5690 ( .A1(n7368), .A2(n7367), .ZN(n5197) );
  NOR2_X1 U5691 ( .A1(n7982), .A2(n5120), .ZN(n8007) );
  NAND2_X1 U5692 ( .A1(n8007), .A2(n8006), .ZN(n8005) );
  INV_X1 U5693 ( .A(n7285), .ZN(n7824) );
  NAND2_X1 U5694 ( .A1(n8754), .A2(n8753), .ZN(n9244) );
  AND2_X1 U5695 ( .A1(n8908), .A2(n8907), .ZN(n9267) );
  AOI21_X1 U5696 ( .B1(n5598), .B2(n5601), .A(n5109), .ZN(n5596) );
  INV_X1 U5697 ( .A(n9261), .ZN(n5601) );
  NOR2_X1 U5698 ( .A1(n5147), .A2(n9331), .ZN(n5146) );
  AND2_X1 U5699 ( .A1(n6905), .A2(n6904), .ZN(n9309) );
  NOR2_X1 U5700 ( .A1(n5055), .A2(n5344), .ZN(n5343) );
  NAND2_X1 U5701 ( .A1(n9305), .A2(n9238), .ZN(n5344) );
  NOR2_X1 U5702 ( .A1(n5342), .A2(n9362), .ZN(n9323) );
  OR2_X1 U5703 ( .A1(n5055), .A2(n9930), .ZN(n5342) );
  OR2_X1 U5704 ( .A1(n9936), .A2(n9350), .ZN(n9318) );
  NAND2_X1 U5705 ( .A1(n6868), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U5706 ( .A1(n9347), .A2(n8888), .ZN(n9330) );
  NAND2_X1 U5707 ( .A1(n9330), .A2(n9331), .ZN(n9317) );
  NAND2_X1 U5708 ( .A1(n8888), .A2(n8788), .ZN(n9349) );
  NAND2_X1 U5709 ( .A1(n9380), .A2(n5476), .ZN(n9356) );
  NOR2_X1 U5710 ( .A1(n8942), .A2(n5477), .ZN(n5476) );
  INV_X1 U5711 ( .A(n8881), .ZN(n5477) );
  NOR2_X1 U5712 ( .A1(n9955), .A2(n5358), .ZN(n5357) );
  INV_X1 U5713 ( .A(n5359), .ZN(n5358) );
  AND2_X1 U5714 ( .A1(n9855), .A2(n5355), .ZN(n9372) );
  NOR2_X1 U5715 ( .A1(n9950), .A2(n5356), .ZN(n5355) );
  INV_X1 U5716 ( .A(n5357), .ZN(n5356) );
  NAND2_X1 U5717 ( .A1(n5611), .A2(n5609), .ZN(n9371) );
  NAND2_X1 U5718 ( .A1(n5610), .A2(n8938), .ZN(n5609) );
  NAND2_X1 U5719 ( .A1(n9399), .A2(n5065), .ZN(n5611) );
  INV_X1 U5720 ( .A(n5612), .ZN(n5610) );
  NAND2_X1 U5721 ( .A1(n9855), .A2(n5359), .ZN(n9400) );
  AND2_X1 U5722 ( .A1(n9877), .A2(n9884), .ZN(n9878) );
  AND2_X1 U5723 ( .A1(n9878), .A2(n9859), .ZN(n9855) );
  NAND2_X1 U5724 ( .A1(n6710), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6725) );
  OR2_X1 U5725 ( .A1(n6725), .A2(n9483), .ZN(n6741) );
  OR2_X1 U5726 ( .A1(n8642), .A2(n8735), .ZN(n8683) );
  OR2_X1 U5727 ( .A1(n6695), .A2(n9472), .ZN(n6711) );
  OR2_X1 U5728 ( .A1(n8426), .A2(n8844), .ZN(n5616) );
  NOR2_X1 U5729 ( .A1(n5351), .A2(n8714), .ZN(n5350) );
  NAND2_X1 U5730 ( .A1(n5466), .A2(n8543), .ZN(n8564) );
  OR2_X1 U5731 ( .A1(n6636), .A2(n9672), .ZN(n6652) );
  AOI21_X1 U5732 ( .B1(n10894), .B2(n10895), .A(n5473), .ZN(n8261) );
  INV_X1 U5733 ( .A(n8824), .ZN(n5473) );
  NAND2_X1 U5734 ( .A1(n8785), .A2(n8201), .ZN(n7831) );
  NOR2_X1 U5735 ( .A1(n9894), .A2(n10873), .ZN(n10891) );
  AND4_X1 U5736 ( .A1(n6571), .A2(n6570), .A3(n6569), .A4(n6568), .ZN(n8449)
         );
  NAND2_X1 U5737 ( .A1(n5348), .A2(n8251), .ZN(n9894) );
  INV_X1 U5738 ( .A(n10802), .ZN(n5348) );
  AOI21_X1 U5739 ( .B1(n5471), .B2(n8258), .A(n5469), .ZN(n5468) );
  NOR2_X1 U5740 ( .A1(n8259), .A2(n5472), .ZN(n5471) );
  NOR2_X1 U5741 ( .A1(n10770), .A2(n8264), .ZN(n10803) );
  NAND2_X1 U5742 ( .A1(n10803), .A2(n10817), .ZN(n10802) );
  AND2_X1 U5743 ( .A1(n6526), .A2(n5062), .ZN(n6527) );
  NAND2_X1 U5744 ( .A1(n5453), .A2(n8256), .ZN(n8325) );
  NOR2_X1 U5745 ( .A1(n8212), .A2(n8920), .ZN(n8211) );
  NAND2_X1 U5746 ( .A1(n7404), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U5747 ( .A1(n9276), .A2(n5363), .ZN(n9916) );
  OR2_X1 U5748 ( .A1(n9285), .A2(n9279), .ZN(n5363) );
  NAND2_X1 U5749 ( .A1(n6884), .A2(n6883), .ZN(n9924) );
  NAND2_X1 U5750 ( .A1(n6785), .A2(n6784), .ZN(n9960) );
  AND2_X1 U5751 ( .A1(n5161), .A2(n8871), .ZN(n9407) );
  NAND2_X1 U5752 ( .A1(n6753), .A2(n6752), .ZN(n9970) );
  NAND2_X1 U5753 ( .A1(n5616), .A2(n5615), .ZN(n11040) );
  OR2_X1 U5754 ( .A1(n7831), .A2(n7830), .ZN(n11070) );
  INV_X1 U5755 ( .A(n10975), .ZN(n11069) );
  NOR2_X1 U5756 ( .A1(n8652), .A2(n6931), .ZN(n10546) );
  INV_X1 U5757 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6455) );
  AND2_X1 U5758 ( .A1(n6922), .A2(n6921), .ZN(n6932) );
  NAND2_X1 U5759 ( .A1(n6915), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U5760 ( .A1(n6914), .A2(n6913), .ZN(n6915) );
  INV_X1 U5761 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6945) );
  INV_X1 U5762 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6917) );
  NOR2_X1 U5763 ( .A1(n5439), .A2(n5279), .ZN(n5278) );
  INV_X1 U5764 ( .A(n6441), .ZN(n5279) );
  NAND2_X1 U5765 ( .A1(n6461), .A2(n5047), .ZN(n5439) );
  NOR2_X1 U5766 ( .A1(n6541), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U5767 ( .A1(n5486), .A2(n5485), .ZN(n8468) );
  AOI21_X1 U5768 ( .B1(n8018), .B2(n5908), .A(n5105), .ZN(n5485) );
  AOI21_X1 U5769 ( .B1(n5087), .B2(n10112), .A(n5516), .ZN(n5515) );
  NAND2_X1 U5770 ( .A1(n5509), .A2(n5506), .ZN(n8699) );
  AOI21_X1 U5771 ( .B1(n5508), .B2(n5107), .A(n5507), .ZN(n5506) );
  NOR2_X1 U5772 ( .A1(n6346), .A2(n6347), .ZN(n5507) );
  INV_X1 U5773 ( .A(n6063), .ZN(n6390) );
  INV_X4 U5774 ( .A(n5688), .ZN(n6388) );
  OR2_X1 U5775 ( .A1(n5896), .A2(n5895), .ZN(n5922) );
  OR2_X1 U5776 ( .A1(n6000), .A2(n5999), .ZN(n6027) );
  OR2_X1 U5777 ( .A1(n6226), .A2(n10106), .ZN(n6251) );
  OR2_X1 U5778 ( .A1(n5922), .A2(n7568), .ZN(n5944) );
  NOR2_X1 U5779 ( .A1(n5944), .A2(n5943), .ZN(n5972) );
  NAND2_X1 U5780 ( .A1(n5662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5680) );
  OR2_X1 U5781 ( .A1(n7114), .A2(n7113), .ZN(n7256) );
  NOR2_X1 U5782 ( .A1(n10255), .A2(n10280), .ZN(n10279) );
  AND2_X1 U5783 ( .A1(n6377), .A2(n6418), .ZN(n8997) );
  NOR2_X1 U5784 ( .A1(n10295), .A2(n10296), .ZN(n10294) );
  AND2_X1 U5785 ( .A1(n8996), .A2(n10314), .ZN(n10311) );
  AND2_X1 U5786 ( .A1(n6332), .A2(n6301), .ZN(n10327) );
  AND2_X1 U5787 ( .A1(n10433), .A2(n5332), .ZN(n10352) );
  NOR2_X1 U5788 ( .A1(n10481), .A2(n5333), .ZN(n5332) );
  INV_X1 U5789 ( .A(n5334), .ZN(n5333) );
  NAND2_X1 U5790 ( .A1(n10433), .A2(n5336), .ZN(n5623) );
  NAND2_X1 U5791 ( .A1(n8981), .A2(n8980), .ZN(n10368) );
  AND2_X1 U5792 ( .A1(n6154), .A2(n6153), .ZN(n10401) );
  NAND2_X1 U5793 ( .A1(n6145), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6176) );
  AND2_X1 U5794 ( .A1(n6183), .A2(n6182), .ZN(n10431) );
  NAND2_X1 U5795 ( .A1(n8974), .A2(n8973), .ZN(n5392) );
  AND2_X1 U5796 ( .A1(n10432), .A2(n10435), .ZN(n10433) );
  NAND2_X1 U5797 ( .A1(n5576), .A2(n5574), .ZN(n10422) );
  INV_X1 U5798 ( .A(n5575), .ZN(n5574) );
  OAI21_X1 U5799 ( .B1(n8630), .B2(n5577), .A(n10427), .ZN(n5575) );
  NOR2_X1 U5800 ( .A1(n6071), .A2(n8065), .ZN(n6100) );
  AND2_X1 U5801 ( .A1(n8576), .A2(n7149), .ZN(n8528) );
  NAND2_X1 U5802 ( .A1(n8164), .A2(n5046), .ZN(n8516) );
  AOI21_X1 U5803 ( .B1(n11008), .B2(n11007), .A(n7057), .ZN(n5622) );
  NAND2_X1 U5804 ( .A1(n5622), .A2(n8392), .ZN(n8512) );
  NAND2_X1 U5805 ( .A1(n8164), .A2(n5042), .ZN(n11001) );
  NAND2_X1 U5806 ( .A1(n8390), .A2(n8389), .ZN(n11008) );
  AND2_X1 U5807 ( .A1(n7162), .A2(n8391), .ZN(n11007) );
  NAND2_X1 U5808 ( .A1(n8164), .A2(n5340), .ZN(n11000) );
  OAI21_X1 U5809 ( .B1(n8152), .B2(n5170), .A(n5168), .ZN(n8390) );
  INV_X1 U5810 ( .A(n5169), .ZN(n5168) );
  OAI21_X1 U5811 ( .B1(n5170), .B2(n8088), .A(n8176), .ZN(n5169) );
  NAND2_X1 U5812 ( .A1(n5173), .A2(n5171), .ZN(n8175) );
  INV_X1 U5813 ( .A(n5170), .ZN(n5171) );
  NAND2_X1 U5814 ( .A1(n5572), .A2(n5573), .ZN(n8172) );
  AND2_X1 U5815 ( .A1(n8164), .A2(n10965), .ZN(n8181) );
  NAND2_X1 U5816 ( .A1(n8152), .A2(n8088), .ZN(n5173) );
  AND2_X1 U5817 ( .A1(n7154), .A2(n8085), .ZN(n8160) );
  AOI21_X1 U5818 ( .B1(n5180), .B2(n7905), .A(n5179), .ZN(n5178) );
  INV_X1 U5819 ( .A(n7906), .ZN(n5179) );
  NAND2_X1 U5820 ( .A1(n10846), .A2(n7904), .ZN(n7936) );
  AND2_X1 U5821 ( .A1(n10841), .A2(n10863), .ZN(n10843) );
  NOR2_X1 U5822 ( .A1(n7811), .A2(n7930), .ZN(n10841) );
  NAND2_X1 U5823 ( .A1(n7909), .A2(n7908), .ZN(n10840) );
  OR2_X1 U5824 ( .A1(n7782), .A2(n7800), .ZN(n7811) );
  AND2_X1 U5825 ( .A1(n7227), .A2(n7230), .ZN(n7768) );
  NOR2_X1 U5826 ( .A1(n7856), .A2(n10738), .ZN(n7783) );
  INV_X1 U5827 ( .A(n5167), .ZN(n7850) );
  CLKBUF_X1 U5828 ( .A(n7120), .Z(n7715) );
  NAND2_X1 U5829 ( .A1(n7007), .A2(n7006), .ZN(n10449) );
  INV_X1 U5830 ( .A(n10452), .ZN(n5326) );
  NAND2_X1 U5831 ( .A1(n10255), .A2(n10739), .ZN(n5325) );
  INV_X1 U5832 ( .A(n10454), .ZN(n5373) );
  AND2_X1 U5833 ( .A1(n6057), .A2(n6056), .ZN(n11084) );
  INV_X1 U5834 ( .A(n7024), .ZN(n10724) );
  INV_X1 U5835 ( .A(n10739), .ZN(n11083) );
  AND2_X1 U5836 ( .A1(n7004), .A2(n7003), .ZN(n8752) );
  OR2_X1 U5837 ( .A1(n7002), .A2(n7001), .ZN(n7004) );
  NAND2_X1 U5838 ( .A1(n10534), .A2(n5645), .ZN(n5181) );
  CLKBUF_X1 U5839 ( .A(n7264), .Z(n10259) );
  OR2_X1 U5840 ( .A1(n5658), .A2(n10534), .ZN(n5659) );
  AND3_X1 U5841 ( .A1(n5183), .A2(n5554), .A3(n5521), .ZN(n5658) );
  OAI21_X1 U5842 ( .B1(n5543), .B2(n6216), .A(n6241), .ZN(n5541) );
  INV_X1 U5843 ( .A(n5543), .ZN(n5542) );
  AND2_X1 U5844 ( .A1(n6269), .A2(n6246), .ZN(n6267) );
  NAND2_X1 U5845 ( .A1(n5529), .A2(n6042), .ZN(n6065) );
  NAND2_X1 U5846 ( .A1(n6019), .A2(n5533), .ZN(n5529) );
  INV_X1 U5847 ( .A(n5311), .ZN(n6044) );
  OAI21_X1 U5848 ( .B1(n5959), .B2(n5084), .A(n5048), .ZN(n5311) );
  NAND2_X1 U5849 ( .A1(n5315), .A2(n5985), .ZN(n6017) );
  NAND2_X1 U5850 ( .A1(n5321), .A2(n5319), .ZN(n5315) );
  NAND2_X1 U5851 ( .A1(n5321), .A2(n5961), .ZN(n5987) );
  XNOR2_X1 U5852 ( .A(n5959), .B(n5958), .ZN(n7555) );
  AND2_X1 U5853 ( .A1(n5919), .A2(n5939), .ZN(n7606) );
  OR2_X1 U5854 ( .A1(n5915), .A2(n5632), .ZN(n5916) );
  NAND2_X1 U5855 ( .A1(n5295), .A2(n5888), .ZN(n5911) );
  NAND2_X1 U5856 ( .A1(n5886), .A2(n5885), .ZN(n5295) );
  AND2_X1 U5857 ( .A1(n5867), .A2(n5917), .ZN(n7488) );
  NAND2_X1 U5858 ( .A1(n5371), .A2(n5838), .ZN(n5861) );
  AND2_X1 U5859 ( .A1(n5839), .A2(n5819), .ZN(n10595) );
  NOR2_X1 U5860 ( .A1(n5281), .A2(n5365), .ZN(n5280) );
  INV_X1 U5861 ( .A(n5767), .ZN(n5365) );
  NOR2_X1 U5862 ( .A1(n5773), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5817) );
  NOR2_X1 U5863 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5712) );
  NOR2_X1 U5864 ( .A1(n10561), .A2(n8348), .ZN(n8349) );
  OR2_X1 U5865 ( .A1(n7949), .A2(n7948), .ZN(n9038) );
  NAND2_X1 U5866 ( .A1(n5415), .A2(n5417), .ZN(n8751) );
  OR2_X1 U5867 ( .A1(n6687), .A2(n5039), .ZN(n5415) );
  AND4_X1 U5868 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n8744)
         );
  NAND2_X1 U5869 ( .A1(n9109), .A2(n6826), .ZN(n9016) );
  NAND2_X1 U5870 ( .A1(n5447), .A2(n6838), .ZN(n9017) );
  NAND2_X1 U5871 ( .A1(n9109), .A2(n6836), .ZN(n5447) );
  OR2_X1 U5872 ( .A1(n8232), .A2(n8231), .ZN(n8403) );
  AND4_X1 U5873 ( .A1(n6539), .A2(n6538), .A3(n6537), .A4(n6536), .ZN(n8326)
         );
  NAND2_X1 U5874 ( .A1(n6953), .A2(n6952), .ZN(n9919) );
  AND2_X1 U5875 ( .A1(n6818), .A2(n6817), .ZN(n9065) );
  AND4_X1 U5876 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n10940)
         );
  NAND2_X1 U5877 ( .A1(n6731), .A2(n8669), .ZN(n8675) );
  NAND2_X1 U5878 ( .A1(n8675), .A2(n6735), .ZN(n9087) );
  NAND2_X1 U5879 ( .A1(n5430), .A2(n5435), .ZN(n9102) );
  NAND2_X1 U5880 ( .A1(n9027), .A2(n9028), .ZN(n5430) );
  AND4_X1 U5881 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n8716)
         );
  NAND2_X1 U5882 ( .A1(n5402), .A2(n5400), .ZN(n8477) );
  AND2_X1 U5883 ( .A1(n5401), .A2(n8401), .ZN(n5400) );
  NAND2_X1 U5884 ( .A1(n8231), .A2(n6646), .ZN(n5401) );
  NAND2_X1 U5885 ( .A1(n6515), .A2(n6516), .ZN(n7999) );
  AND2_X1 U5886 ( .A1(n6762), .A2(n5421), .ZN(n5420) );
  NAND2_X1 U5887 ( .A1(n8675), .A2(n5424), .ZN(n9121) );
  AOI21_X1 U5888 ( .B1(n5411), .B2(n5413), .A(n5126), .ZN(n5408) );
  NAND2_X1 U5889 ( .A1(n8028), .A2(n5411), .ZN(n5409) );
  AOI21_X1 U5890 ( .B1(n5412), .B2(n7966), .A(n5079), .ZN(n5411) );
  AND2_X1 U5891 ( .A1(n6557), .A2(n6556), .ZN(n8250) );
  AND3_X1 U5892 ( .A1(n6555), .A2(n6554), .A3(n6553), .ZN(n6557) );
  OR2_X1 U5893 ( .A1(n9080), .A2(n10939), .ZN(n9127) );
  AND2_X1 U5894 ( .A1(n9049), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9129) );
  NAND2_X1 U5895 ( .A1(n5410), .A2(n7966), .ZN(n7976) );
  NAND2_X1 U5896 ( .A1(n8028), .A2(n6548), .ZN(n5410) );
  AOI21_X1 U5897 ( .B1(n5040), .B2(n5452), .A(n5442), .ZN(n5441) );
  INV_X1 U5898 ( .A(n6863), .ZN(n5442) );
  AND2_X1 U5899 ( .A1(n6974), .A2(n6949), .ZN(n9135) );
  NAND2_X1 U5900 ( .A1(n6956), .A2(n9849), .ZN(n9098) );
  INV_X1 U5901 ( .A(n9135), .ZN(n9086) );
  NAND2_X1 U5902 ( .A1(n7274), .A2(n10648), .ZN(n10547) );
  INV_X1 U5903 ( .A(n8250), .ZN(n9893) );
  NAND4_X1 U5904 ( .A1(n6504), .A2(n6503), .A3(n6502), .A4(n6501), .ZN(n9158)
         );
  NAND2_X1 U5905 ( .A1(n5060), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6503) );
  NAND4_X1 U5906 ( .A1(n6492), .A2(n6491), .A3(n6490), .A4(n6489), .ZN(n9161)
         );
  INV_X2 U5907 ( .A(P2_U3966), .ZN(n9160) );
  NOR2_X1 U5908 ( .A1(n10674), .A2(n5069), .ZN(n7344) );
  INV_X1 U5909 ( .A(n5195), .ZN(n7342) );
  NOR2_X1 U5910 ( .A1(n7353), .A2(n5108), .ZN(n7332) );
  INV_X1 U5911 ( .A(n5201), .ZN(n7330) );
  NOR2_X1 U5912 ( .A1(n7380), .A2(n7379), .ZN(n7378) );
  AND2_X1 U5913 ( .A1(n5201), .A2(n5200), .ZN(n7380) );
  NAND2_X1 U5914 ( .A1(n7297), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5200) );
  INV_X1 U5915 ( .A(n5199), .ZN(n7365) );
  AND2_X1 U5916 ( .A1(n5199), .A2(n5198), .ZN(n7368) );
  NAND2_X1 U5917 ( .A1(n7370), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5198) );
  INV_X1 U5918 ( .A(n5197), .ZN(n7389) );
  NOR2_X1 U5919 ( .A1(n7867), .A2(n5121), .ZN(n7870) );
  NOR2_X1 U5920 ( .A1(n7870), .A2(n7869), .ZN(n7982) );
  AND2_X1 U5921 ( .A1(n7303), .A2(n6975), .ZN(n10684) );
  INV_X1 U5922 ( .A(n10677), .ZN(n10651) );
  NAND2_X1 U5923 ( .A1(n8777), .A2(n8776), .ZN(n9907) );
  NAND2_X1 U5924 ( .A1(n8774), .A2(n6511), .ZN(n8777) );
  INV_X1 U5925 ( .A(n9244), .ZN(n9914) );
  OR2_X1 U5926 ( .A1(n9244), .A2(n9276), .ZN(n9911) );
  AND2_X1 U5927 ( .A1(n9295), .A2(n9294), .ZN(n9922) );
  INV_X1 U5928 ( .A(n9924), .ZN(n9305) );
  NAND2_X1 U5929 ( .A1(n5597), .A2(n9261), .ZN(n9299) );
  AND2_X1 U5930 ( .A1(n6869), .A2(n6843), .ZN(n9334) );
  NAND2_X1 U5931 ( .A1(n9339), .A2(n9256), .ZN(n9329) );
  INV_X1 U5932 ( .A(n9945), .ZN(n9367) );
  NAND2_X1 U5933 ( .A1(n8760), .A2(n8759), .ZN(n9376) );
  NAND2_X1 U5934 ( .A1(n9398), .A2(n9253), .ZN(n9385) );
  NAND2_X1 U5935 ( .A1(n5162), .A2(n5455), .ZN(n9861) );
  OR2_X1 U5936 ( .A1(n5454), .A2(n5458), .ZN(n5162) );
  INV_X1 U5937 ( .A(n9970), .ZN(n9859) );
  AOI21_X1 U5938 ( .B1(n8680), .B2(n5464), .A(n5462), .ZN(n5456) );
  NOR2_X1 U5939 ( .A1(n9249), .A2(n5626), .ZN(n9870) );
  AND2_X1 U5940 ( .A1(n6724), .A2(n6723), .ZN(n8687) );
  OAI21_X1 U5941 ( .B1(n8680), .B2(n8679), .A(n8859), .ZN(n8756) );
  AND2_X1 U5942 ( .A1(n5211), .A2(n8635), .ZN(n8676) );
  INV_X1 U5943 ( .A(n5211), .ZN(n8637) );
  NOR2_X1 U5944 ( .A1(n10933), .A2(n5352), .ZN(n8428) );
  INV_X1 U5945 ( .A(n5222), .ZN(n5220) );
  NAND2_X1 U5946 ( .A1(n9898), .A2(n8254), .ZN(n8456) );
  NAND2_X1 U5947 ( .A1(n10775), .A2(n8811), .ZN(n10809) );
  INV_X1 U5948 ( .A(n10769), .ZN(n8247) );
  INV_X1 U5949 ( .A(n9849), .ZN(n10962) );
  OR2_X1 U5950 ( .A1(n8203), .A2(n8780), .ZN(n10952) );
  INV_X1 U5951 ( .A(n10956), .ZN(n9901) );
  INV_X1 U5952 ( .A(n10952), .ZN(n9897) );
  NAND2_X1 U5953 ( .A1(n10957), .A2(n10904), .ZN(n9887) );
  AND2_X2 U5954 ( .A1(n7835), .A2(n8198), .ZN(n11078) );
  NAND2_X1 U5955 ( .A1(n5232), .A2(n5231), .ZN(n9987) );
  NOR2_X1 U5956 ( .A1(n9917), .A2(n5233), .ZN(n5232) );
  NAND2_X1 U5957 ( .A1(n9915), .A2(n11074), .ZN(n5231) );
  OAI21_X1 U5958 ( .B1(n9916), .B2(n11070), .A(n5080), .ZN(n5233) );
  AND2_X2 U5959 ( .A1(n7835), .A2(n7822), .ZN(n11082) );
  INV_X1 U5960 ( .A(n6483), .ZN(n10008) );
  INV_X1 U5961 ( .A(n6932), .ZN(n8652) );
  XNOR2_X1 U5962 ( .A(n6918), .B(n6917), .ZN(n8462) );
  NAND2_X1 U5963 ( .A1(n6916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U5964 ( .A1(n6946), .A2(n6945), .ZN(n6916) );
  INV_X1 U5965 ( .A(n8947), .ZN(n8201) );
  AOI21_X1 U5966 ( .B1(n5406), .B2(n10002), .A(n10002), .ZN(n5403) );
  INV_X1 U5967 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7538) );
  INV_X1 U5968 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7451) );
  NAND2_X1 U5969 ( .A1(n6458), .A2(n5191), .ZN(n7430) );
  AOI22_X1 U5970 ( .A1(n5083), .A2(P2_IR_REG_0__SCAN_IN), .B1(n5193), .B2(
        n5192), .ZN(n5191) );
  INV_X1 U5971 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5193) );
  INV_X1 U5972 ( .A(n7910), .ZN(n10863) );
  INV_X1 U5973 ( .A(n7734), .ZN(n10850) );
  OR2_X1 U5974 ( .A1(n6426), .A2(n6425), .ZN(n10118) );
  NAND2_X1 U5975 ( .A1(n6352), .A2(n6351), .ZN(n10461) );
  NAND2_X1 U5976 ( .A1(n8553), .A2(n5059), .ZN(n8654) );
  NAND2_X1 U5977 ( .A1(n8553), .A2(n8554), .ZN(n5494) );
  NAND2_X1 U5978 ( .A1(n6144), .A2(n6143), .ZN(n10503) );
  NAND2_X1 U5979 ( .A1(n6298), .A2(n6297), .ZN(n10471) );
  NAND2_X1 U5980 ( .A1(n6088), .A2(n6087), .ZN(n10075) );
  NAND2_X1 U5981 ( .A1(n6097), .A2(n6096), .ZN(n10514) );
  NAND2_X1 U5982 ( .A1(n5489), .A2(n10028), .ZN(n10092) );
  AND2_X1 U5983 ( .A1(n6205), .A2(n6204), .ZN(n10402) );
  NAND2_X1 U5984 ( .A1(n10040), .A2(n10036), .ZN(n10102) );
  CLKBUF_X1 U5985 ( .A(n8220), .Z(n8221) );
  NAND2_X1 U5986 ( .A1(n8221), .A2(n8223), .ZN(n8222) );
  NAND2_X1 U5987 ( .A1(n5735), .A2(n5732), .ZN(n7653) );
  INV_X1 U5988 ( .A(n10118), .ZN(n10147) );
  NAND2_X1 U5989 ( .A1(n6088), .A2(n5043), .ZN(n5518) );
  NAND2_X1 U5990 ( .A1(n6118), .A2(n6117), .ZN(n10507) );
  NAND2_X1 U5991 ( .A1(n6415), .A2(n10865), .ZN(n10131) );
  AOI21_X1 U5992 ( .B1(n10083), .B2(n5511), .A(n5107), .ZN(n10124) );
  OR2_X1 U5993 ( .A1(n6426), .A2(n6412), .ZN(n10133) );
  OR2_X1 U5994 ( .A1(n6426), .A2(n6417), .ZN(n10149) );
  INV_X1 U5995 ( .A(n10133), .ZN(n10143) );
  OR2_X1 U5996 ( .A1(n6431), .A2(n7597), .ZN(n10152) );
  INV_X1 U5997 ( .A(n10359), .ZN(n10159) );
  INV_X1 U5998 ( .A(n10402), .ZN(n10162) );
  OR2_X1 U5999 ( .A1(n7497), .A2(n7270), .ZN(n10176) );
  AOI21_X1 U6000 ( .B1(n8774), .B2(n7005), .A(n7000), .ZN(n10445) );
  XNOR2_X1 U6001 ( .A(n5284), .B(n10272), .ZN(n10454) );
  NAND2_X1 U6002 ( .A1(n10268), .A2(n5285), .ZN(n5284) );
  NAND2_X1 U6003 ( .A1(n10455), .A2(n10274), .ZN(n5285) );
  NAND2_X1 U6004 ( .A1(n5302), .A2(n5303), .ZN(n10287) );
  AOI211_X1 U6005 ( .C1(n11009), .C2(n10310), .A(n10309), .B(n10308), .ZN(
        n10468) );
  NOR2_X1 U6006 ( .A1(n10322), .A2(n10321), .ZN(n10320) );
  INV_X1 U6007 ( .A(n5378), .ZN(n10339) );
  NAND2_X1 U6008 ( .A1(n5297), .A2(n5298), .ZN(n10333) );
  NAND2_X1 U6009 ( .A1(n5384), .A2(n8982), .ZN(n10357) );
  NAND2_X1 U6010 ( .A1(n10367), .A2(n8963), .ZN(n10351) );
  AND2_X1 U6011 ( .A1(n6225), .A2(n6224), .ZN(n10485) );
  NAND2_X1 U6012 ( .A1(n10386), .A2(n10385), .ZN(n10384) );
  NAND2_X1 U6013 ( .A1(n10405), .A2(n8962), .ZN(n10386) );
  INV_X1 U6014 ( .A(n8631), .ZN(n5578) );
  NAND2_X1 U6015 ( .A1(n5176), .A2(n8603), .ZN(n8606) );
  NAND2_X1 U6016 ( .A1(n5557), .A2(n5559), .ZN(n8599) );
  AND2_X1 U6017 ( .A1(n5559), .A2(n5053), .ZN(n8585) );
  NAND2_X1 U6018 ( .A1(n10869), .A2(n7701), .ZN(n11029) );
  NAND2_X1 U6019 ( .A1(n7802), .A2(n7801), .ZN(n7804) );
  NAND2_X1 U6020 ( .A1(n5329), .A2(n7470), .ZN(n5328) );
  OR2_X1 U6021 ( .A1(n7470), .A2(n10625), .ZN(n5327) );
  NAND2_X1 U6022 ( .A1(n5330), .A2(n5049), .ZN(n5329) );
  OR2_X1 U6023 ( .A1(n7575), .A2(n7577), .ZN(n10865) );
  INV_X1 U6024 ( .A(n11029), .ZN(n10413) );
  AND2_X1 U6025 ( .A1(n10439), .A2(n10515), .ZN(n11022) );
  INV_X1 U6026 ( .A(n10453), .ZN(n5308) );
  NAND2_X1 U6027 ( .A1(n10458), .A2(n5186), .ZN(n10522) );
  AND2_X1 U6028 ( .A1(n5187), .A2(n10457), .ZN(n5186) );
  OR2_X1 U6029 ( .A1(n10459), .A2(n10741), .ZN(n5187) );
  AND2_X1 U6030 ( .A1(n7495), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7426) );
  NAND2_X1 U6031 ( .A1(n5660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5661) );
  INV_X1 U6032 ( .A(n5644), .ZN(n5642) );
  NAND2_X1 U6033 ( .A1(n7014), .A2(n7013), .ZN(n8764) );
  OR2_X1 U6034 ( .A1(n5656), .A2(n9798), .ZN(n5657) );
  INV_X1 U6035 ( .A(n6393), .ZN(n8416) );
  INV_X1 U6036 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9737) );
  INV_X1 U6037 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9736) );
  OR2_X1 U6038 ( .A1(n5967), .A2(n5555), .ZN(n5683) );
  INV_X1 U6039 ( .A(n5631), .ZN(n5555) );
  AND2_X1 U6040 ( .A1(n6024), .A2(n6066), .ZN(n10217) );
  INV_X1 U6041 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7540) );
  INV_X1 U6042 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U6043 ( .A1(n5364), .A2(n5767), .ZN(n5797) );
  NAND2_X1 U6044 ( .A1(n5765), .A2(n5764), .ZN(n5364) );
  NOR2_X1 U6045 ( .A1(n8370), .A2(n8369), .ZN(n10578) );
  NOR2_X1 U6046 ( .A1(n10576), .A2(n10575), .ZN(n8369) );
  AOI21_X1 U6047 ( .B1(n5204), .B2(n10649), .A(n5202), .ZN(n9236) );
  OAI21_X1 U6048 ( .B1(n7263), .B2(n8040), .A(n7262), .ZN(n7269) );
  NAND2_X1 U6049 ( .A1(n5375), .A2(n11093), .ZN(n5374) );
  NAND2_X1 U6050 ( .A1(n5307), .A2(n5305), .ZN(P1_U3520) );
  OR2_X1 U6051 ( .A1(n11097), .A2(n5306), .ZN(n5305) );
  OAI21_X1 U6052 ( .B1(n5375), .B2(n5308), .A(n11097), .ZN(n5307) );
  INV_X1 U6053 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5306) );
  INV_X1 U6054 ( .A(n6533), .ZN(n6590) );
  AND2_X2 U6055 ( .A1(n6482), .A2(n6483), .ZN(n6550) );
  OAI21_X1 U6056 ( .B1(n10321), .B2(n8986), .A(n8988), .ZN(n5391) );
  AND2_X1 U6057 ( .A1(n5215), .A2(n8670), .ZN(n5038) );
  NOR2_X2 U6058 ( .A1(n6482), .A2(n6483), .ZN(n5060) );
  AND2_X1 U6059 ( .A1(n8745), .A2(n6689), .ZN(n5039) );
  OR2_X1 U6060 ( .A1(n11051), .A2(n9150), .ZN(n8635) );
  AND2_X1 U6061 ( .A1(n8845), .A2(n8541), .ZN(n8844) );
  AND2_X1 U6062 ( .A1(n5057), .A2(n5443), .ZN(n5040) );
  XNOR2_X1 U6063 ( .A(n5960), .B(n5938), .ZN(n5958) );
  INV_X1 U6064 ( .A(n10321), .ZN(n5304) );
  AND2_X1 U6065 ( .A1(n10094), .A2(n10093), .ZN(n5041) );
  AND2_X1 U6066 ( .A1(n5340), .A2(n5339), .ZN(n5042) );
  INV_X1 U6067 ( .A(n5458), .ZN(n5457) );
  NAND2_X1 U6068 ( .A1(n9873), .A2(n5459), .ZN(n5458) );
  NOR2_X1 U6069 ( .A1(n6109), .A2(n5519), .ZN(n5043) );
  AND2_X1 U6070 ( .A1(n5501), .A2(n5982), .ZN(n5044) );
  INV_X1 U6071 ( .A(n8815), .ZN(n5469) );
  AND2_X1 U6072 ( .A1(n8816), .A2(n8818), .ZN(n9900) );
  NOR2_X1 U6073 ( .A1(n6474), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5045) );
  INV_X1 U6074 ( .A(n8094), .ZN(n10965) );
  NOR2_X1 U6075 ( .A1(n9362), .A2(n5055), .ZN(n5345) );
  AND2_X1 U6076 ( .A1(n5042), .A2(n5338), .ZN(n5046) );
  AND4_X1 U6077 ( .A1(n6487), .A2(n6486), .A3(n6485), .A4(n6484), .ZN(n8194)
         );
  INV_X1 U6078 ( .A(n8194), .ZN(n9159) );
  AND2_X1 U6079 ( .A1(n6462), .A2(n6442), .ZN(n5047) );
  OR2_X1 U6080 ( .A1(n5316), .A2(n5534), .ZN(n5048) );
  NAND2_X1 U6081 ( .A1(n6995), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5049) );
  NAND3_X1 U6082 ( .A1(n5554), .A2(n5631), .A3(n5097), .ZN(n5050) );
  OR2_X1 U6083 ( .A1(n10476), .A2(n10359), .ZN(n8986) );
  NOR2_X1 U6084 ( .A1(n5146), .A2(n5148), .ZN(n5051) );
  NAND2_X1 U6085 ( .A1(n6840), .A2(n6839), .ZN(n9936) );
  INV_X1 U6086 ( .A(n9254), .ZN(n5244) );
  NAND2_X1 U6087 ( .A1(n5223), .A2(n5220), .ZN(n8422) );
  INV_X1 U6088 ( .A(n9238), .ZN(n9930) );
  NAND2_X1 U6089 ( .A1(n6477), .A2(n5137), .ZN(n6975) );
  INV_X1 U6090 ( .A(n10932), .ZN(n5353) );
  INV_X1 U6091 ( .A(n7966), .ZN(n5413) );
  NAND2_X1 U6092 ( .A1(n5173), .A2(n8086), .ZN(n5052) );
  INV_X4 U6093 ( .A(n6540), .ZN(n6511) );
  CLKBUF_X3 U6094 ( .A(n5790), .Z(n6302) );
  OR2_X1 U6095 ( .A1(n8583), .A2(n8582), .ZN(n5053) );
  NAND2_X1 U6096 ( .A1(n6488), .A2(n5427), .ZN(n8780) );
  XOR2_X1 U6097 ( .A(n8664), .B(n11004), .Z(n5054) );
  OR2_X1 U6098 ( .A1(n9936), .A2(n9939), .ZN(n5055) );
  NAND2_X1 U6099 ( .A1(n5035), .A2(n7404), .ZN(n5763) );
  NAND2_X1 U6100 ( .A1(n9807), .A2(n9798), .ZN(n5056) );
  AND2_X1 U6101 ( .A1(n5450), .A2(n5448), .ZN(n5057) );
  INV_X1 U6102 ( .A(n8816), .ZN(n5144) );
  NOR2_X1 U6103 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6457) );
  INV_X1 U6104 ( .A(n6995), .ZN(n7404) );
  OR2_X1 U6105 ( .A1(n7306), .A2(n7430), .ZN(n5058) );
  AND2_X1 U6106 ( .A1(n7017), .A2(n7016), .ZN(n10283) );
  AND2_X1 U6107 ( .A1(n6039), .A2(n8554), .ZN(n5059) );
  NAND2_X1 U6108 ( .A1(n10083), .A2(n6288), .ZN(n10048) );
  AOI21_X1 U6109 ( .B1(n6481), .B2(P2_IR_REG_29__SCAN_IN), .A(n6480), .ZN(
        n6482) );
  AND2_X1 U6110 ( .A1(n8918), .A2(n8912), .ZN(n5061) );
  XNOR2_X1 U6111 ( .A(n6998), .B(n6997), .ZN(n8774) );
  NAND2_X1 U6112 ( .A1(n5392), .A2(n8975), .ZN(n10424) );
  NAND2_X1 U6113 ( .A1(n6770), .A2(n6769), .ZN(n9967) );
  OR2_X1 U6114 ( .A1(n7306), .A2(n7408), .ZN(n5062) );
  NAND2_X1 U6115 ( .A1(n9930), .A2(n9308), .ZN(n8917) );
  INV_X1 U6116 ( .A(n6018), .ZN(n5534) );
  OR2_X1 U6117 ( .A1(n10965), .A2(n8309), .ZN(n5063) );
  AND2_X1 U6118 ( .A1(n8940), .A2(n8873), .ZN(n5064) );
  INV_X1 U6119 ( .A(n5619), .ZN(n6541) );
  NAND2_X1 U6120 ( .A1(n5619), .A2(n5620), .ZN(n6572) );
  AND2_X1 U6121 ( .A1(n8938), .A2(n9406), .ZN(n5065) );
  NAND2_X1 U6122 ( .A1(n7306), .A2(n7404), .ZN(n6573) );
  NAND2_X1 U6123 ( .A1(n6173), .A2(n6172), .ZN(n10496) );
  NAND2_X1 U6124 ( .A1(n5971), .A2(n5970), .ZN(n8385) );
  INV_X1 U6125 ( .A(n5452), .ZN(n5445) );
  NOR2_X1 U6126 ( .A1(n6838), .A2(n9018), .ZN(n5452) );
  AND2_X1 U6127 ( .A1(n9380), .A2(n8881), .ZN(n5066) );
  INV_X1 U6128 ( .A(n8996), .ZN(n10319) );
  NOR2_X1 U6129 ( .A1(n10334), .A2(n10471), .ZN(n8996) );
  AND2_X1 U6130 ( .A1(n9052), .A2(n5428), .ZN(n5067) );
  INV_X1 U6131 ( .A(n5345), .ZN(n5347) );
  INV_X1 U6132 ( .A(n10388), .ZN(n10385) );
  AND2_X1 U6133 ( .A1(n8980), .A2(n7074), .ZN(n10388) );
  AND2_X1 U6134 ( .A1(n6867), .A2(n6866), .ZN(n9238) );
  AND2_X1 U6135 ( .A1(n9290), .A2(n8902), .ZN(n5068) );
  AND2_X1 U6136 ( .A1(n10683), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5069) );
  INV_X1 U6137 ( .A(n5985), .ZN(n5318) );
  NAND2_X1 U6138 ( .A1(n5964), .A2(n5963), .ZN(n5985) );
  AND2_X1 U6139 ( .A1(n10493), .A2(n10162), .ZN(n5070) );
  AND2_X1 U6140 ( .A1(n9884), .A2(n9862), .ZN(n5071) );
  OR2_X1 U6141 ( .A1(n8701), .A2(n6413), .ZN(n5072) );
  AND2_X1 U6142 ( .A1(n8828), .A2(n8829), .ZN(n8926) );
  AND2_X1 U6143 ( .A1(n10481), .A2(n10160), .ZN(n5073) );
  AND2_X1 U6144 ( .A1(n7159), .A2(n8389), .ZN(n8176) );
  OR2_X1 U6145 ( .A1(n9977), .A2(n9862), .ZN(n9250) );
  OR2_X1 U6146 ( .A1(n7306), .A2(n7418), .ZN(n5074) );
  AND2_X1 U6147 ( .A1(n10465), .A2(n10052), .ZN(n5075) );
  INV_X1 U6148 ( .A(n5272), .ZN(n5271) );
  NAND2_X1 U6149 ( .A1(n9853), .A2(n5273), .ZN(n5272) );
  NOR2_X1 U6150 ( .A1(n9405), .A2(n9842), .ZN(n9252) );
  INV_X1 U6151 ( .A(n5884), .ZN(n5885) );
  XNOR2_X1 U6152 ( .A(n5887), .B(SI_8_), .ZN(n5884) );
  OR2_X1 U6153 ( .A1(n9955), .A2(n9408), .ZN(n8938) );
  AND2_X1 U6154 ( .A1(n6046), .A2(SI_15_), .ZN(n5076) );
  OR2_X1 U6155 ( .A1(n6662), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5077) );
  AND2_X1 U6156 ( .A1(n5862), .A2(SI_7_), .ZN(n5078) );
  AND2_X1 U6157 ( .A1(n6563), .A2(n7974), .ZN(n5079) );
  NAND2_X1 U6158 ( .A1(n9918), .A2(n10975), .ZN(n5080) );
  NAND2_X1 U6159 ( .A1(n5630), .A2(n8598), .ZN(n5081) );
  AND2_X1 U6160 ( .A1(n5984), .A2(n8302), .ZN(n5082) );
  NAND2_X1 U6161 ( .A1(n7677), .A2(n5756), .ZN(n5504) );
  AND2_X1 U6162 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5083) );
  NAND2_X1 U6163 ( .A1(n5958), .A2(n5314), .ZN(n5084) );
  OR2_X1 U6164 ( .A1(n10112), .A2(n10113), .ZN(n5085) );
  NOR2_X1 U6165 ( .A1(n11036), .A2(n8744), .ZN(n5086) );
  NAND2_X1 U6166 ( .A1(n6108), .A2(n5517), .ZN(n5087) );
  OR2_X1 U6167 ( .A1(n5250), .A2(n5213), .ZN(n5088) );
  INV_X1 U6168 ( .A(n8908), .ZN(n5157) );
  INV_X1 U6169 ( .A(n6460), .ZN(n6461) );
  NAND3_X1 U6170 ( .A1(n5637), .A2(n5636), .A3(n5641), .ZN(n5522) );
  INV_X1 U6171 ( .A(n5522), .ZN(n5183) );
  AND3_X1 U6172 ( .A1(n5229), .A2(n5163), .A3(n5619), .ZN(n5089) );
  NOR2_X1 U6173 ( .A1(n9955), .A2(n9377), .ZN(n5090) );
  AND2_X1 U6174 ( .A1(n5496), .A2(n10104), .ZN(n5091) );
  NAND2_X1 U6175 ( .A1(n7196), .A2(n7143), .ZN(n10296) );
  INV_X1 U6176 ( .A(n10314), .ZN(n10465) );
  AND2_X1 U6177 ( .A1(n6329), .A2(n6328), .ZN(n10314) );
  AND2_X1 U6178 ( .A1(n8604), .A2(n8603), .ZN(n5092) );
  AND2_X1 U6179 ( .A1(n8940), .A2(n8871), .ZN(n5093) );
  NAND2_X1 U6180 ( .A1(n8901), .A2(n8900), .ZN(n9307) );
  NAND2_X1 U6181 ( .A1(n10476), .A2(n10159), .ZN(n5094) );
  AND2_X1 U6182 ( .A1(n8849), .A2(n8850), .ZN(n5095) );
  AND2_X1 U6183 ( .A1(n5242), .A2(n8886), .ZN(n5096) );
  AND2_X1 U6184 ( .A1(n5637), .A2(n5636), .ZN(n5097) );
  AND2_X1 U6185 ( .A1(n9267), .A2(n8905), .ZN(n5098) );
  AND2_X1 U6186 ( .A1(n7211), .A2(n10270), .ZN(n8992) );
  AND2_X1 U6187 ( .A1(n7131), .A2(n8975), .ZN(n5099) );
  AND2_X1 U6188 ( .A1(n8881), .A2(n8883), .ZN(n9254) );
  AND2_X1 U6189 ( .A1(n8787), .A2(n9914), .ZN(n5100) );
  AND2_X1 U6190 ( .A1(n5152), .A2(n8787), .ZN(n5101) );
  INV_X1 U6191 ( .A(n5568), .ZN(n5567) );
  NAND2_X1 U6192 ( .A1(n5627), .A2(n8967), .ZN(n5568) );
  NAND2_X1 U6193 ( .A1(n8896), .A2(n8888), .ZN(n5102) );
  NOR2_X1 U6194 ( .A1(n9155), .A2(n8423), .ZN(n5103) );
  AND2_X1 U6195 ( .A1(n6450), .A2(n5621), .ZN(n5104) );
  INV_X1 U6196 ( .A(n9936), .ZN(n5346) );
  INV_X1 U6197 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U6198 ( .A1(n10935), .A2(n8836), .ZN(n8539) );
  INV_X1 U6199 ( .A(n10036), .ZN(n5497) );
  NAND2_X1 U6200 ( .A1(n9026), .A2(n9028), .ZN(n9025) );
  XOR2_X1 U6201 ( .A(n5930), .B(n5686), .Z(n5105) );
  OR2_X1 U6202 ( .A1(n9843), .A2(n9251), .ZN(n5106) );
  AND2_X1 U6203 ( .A1(n6315), .A2(n6314), .ZN(n5107) );
  INV_X1 U6204 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5287) );
  AND2_X1 U6205 ( .A1(n7295), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6206 ( .A1(n5518), .A2(n6108), .ZN(n10111) );
  INV_X1 U6207 ( .A(n5456), .ZN(n9872) );
  NAND2_X1 U6208 ( .A1(n8222), .A2(n5957), .ZN(n8301) );
  INV_X1 U6209 ( .A(n10113), .ZN(n5517) );
  AND2_X1 U6210 ( .A1(n9305), .A2(n9262), .ZN(n5109) );
  INV_X1 U6211 ( .A(n10338), .ZN(n5190) );
  INV_X1 U6212 ( .A(n10028), .ZN(n5488) );
  NAND2_X1 U6213 ( .A1(n5606), .A2(n5605), .ZN(n9868) );
  INV_X1 U6214 ( .A(n5226), .ZN(n10929) );
  OR2_X1 U6215 ( .A1(n9362), .A2(n9939), .ZN(n5110) );
  AND3_X1 U6216 ( .A1(n5167), .A2(n7583), .A3(n7715), .ZN(n5111) );
  NAND2_X1 U6217 ( .A1(n6615), .A2(n6441), .ZN(n6662) );
  NAND2_X1 U6218 ( .A1(n5229), .A2(n5619), .ZN(n6607) );
  AND2_X1 U6219 ( .A1(n6383), .A2(n6382), .ZN(n10297) );
  AND2_X1 U6220 ( .A1(n6469), .A2(n6471), .ZN(n5112) );
  NAND2_X1 U6221 ( .A1(n10433), .A2(n5334), .ZN(n5337) );
  INV_X1 U6222 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5360) );
  INV_X1 U6223 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6224 ( .A1(n9855), .A2(n5357), .ZN(n5113) );
  AND2_X1 U6225 ( .A1(n9398), .A2(n5612), .ZN(n5114) );
  INV_X1 U6226 ( .A(n9256), .ZN(n5591) );
  OR2_X1 U6227 ( .A1(n9939), .A2(n9357), .ZN(n9256) );
  NAND2_X1 U6228 ( .A1(n8158), .A2(n8157), .ZN(n5115) );
  INV_X1 U6229 ( .A(n5512), .ZN(n5511) );
  NAND2_X1 U6230 ( .A1(n5634), .A2(n6288), .ZN(n5512) );
  AND2_X1 U6231 ( .A1(n6702), .A2(n6701), .ZN(n5116) );
  NAND2_X1 U6232 ( .A1(n10278), .A2(n10277), .ZN(n5117) );
  OR2_X1 U6233 ( .A1(n8539), .A2(n8846), .ZN(n5466) );
  AND2_X1 U6234 ( .A1(n5616), .A2(n8536), .ZN(n5118) );
  NAND2_X1 U6235 ( .A1(n5278), .A2(n6615), .ZN(n5119) );
  NAND2_X1 U6236 ( .A1(n5998), .A2(n5997), .ZN(n8552) );
  INV_X1 U6237 ( .A(n8552), .ZN(n5339) );
  INV_X1 U6238 ( .A(n8669), .ZN(n5422) );
  NAND2_X1 U6239 ( .A1(n6026), .A2(n6025), .ZN(n8664) );
  INV_X1 U6240 ( .A(n8664), .ZN(n5338) );
  INV_X1 U6241 ( .A(n8554), .ZN(n5493) );
  NAND2_X1 U6242 ( .A1(n5399), .A2(n5398), .ZN(n8135) );
  NAND2_X1 U6243 ( .A1(n6709), .A2(n6708), .ZN(n8735) );
  INV_X1 U6244 ( .A(n8735), .ZN(n5215) );
  AND2_X1 U6245 ( .A1(n5396), .A2(n5394), .ZN(n8027) );
  XNOR2_X1 U6246 ( .A(n5661), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6395) );
  AND2_X1 U6247 ( .A1(n7991), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5120) );
  AND2_X1 U6248 ( .A1(n7663), .A2(n5756), .ZN(n7678) );
  AND2_X1 U6249 ( .A1(n7873), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6250 ( .A1(n5142), .A2(n8816), .ZN(n8447) );
  NAND2_X1 U6251 ( .A1(n5883), .A2(n8127), .ZN(n8017) );
  NAND2_X1 U6252 ( .A1(n8475), .A2(n8226), .ZN(n8085) );
  INV_X1 U6253 ( .A(n8085), .ZN(n5393) );
  OR2_X1 U6254 ( .A1(n10933), .A2(n10932), .ZN(n5122) );
  XNOR2_X1 U6255 ( .A(n6914), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6947) );
  INV_X1 U6256 ( .A(n6475), .ZN(n6921) );
  NAND2_X1 U6257 ( .A1(n10845), .A2(n7903), .ZN(n10846) );
  AND2_X1 U6258 ( .A1(n5475), .A2(n6615), .ZN(n6923) );
  NAND2_X1 U6259 ( .A1(n7664), .A2(n7665), .ZN(n7663) );
  AND2_X1 U6260 ( .A1(n7233), .A2(n7227), .ZN(n5123) );
  AND2_X1 U6261 ( .A1(n8417), .A2(n8828), .ZN(n5124) );
  NOR2_X1 U6262 ( .A1(n8422), .A2(n8926), .ZN(n5125) );
  NAND2_X1 U6263 ( .A1(n5393), .A2(n8084), .ZN(n8086) );
  INV_X1 U6264 ( .A(n10974), .ZN(n5354) );
  AND2_X2 U6265 ( .A1(n7588), .A2(n7702), .ZN(n11093) );
  OR2_X1 U6266 ( .A1(n7290), .A2(n9239), .ZN(n10673) );
  AND2_X1 U6267 ( .A1(n7705), .A2(n8040), .ZN(n10515) );
  INV_X1 U6268 ( .A(n10515), .ZN(n11085) );
  XOR2_X1 U6269 ( .A(n6579), .B(n6577), .Z(n5126) );
  NAND2_X1 U6270 ( .A1(n6626), .A2(n6614), .ZN(n5127) );
  INV_X1 U6271 ( .A(n8258), .ZN(n10768) );
  NAND2_X1 U6272 ( .A1(n8811), .A2(n8809), .ZN(n8258) );
  XOR2_X1 U6273 ( .A(n9846), .B(n9233), .Z(n5128) );
  OR2_X1 U6274 ( .A1(n9232), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6275 ( .A1(n5692), .A2(n7628), .ZN(n7592) );
  NOR2_X1 U6276 ( .A1(n8699), .A2(n8698), .ZN(n8701) );
  OAI22_X1 U6277 ( .A1(n8553), .A2(n5490), .B1(n5059), .B2(n5491), .ZN(n10058)
         );
  NAND2_X1 U6278 ( .A1(n5545), .A2(n5098), .ZN(n5264) );
  NAND2_X1 U6279 ( .A1(n5260), .A2(n8915), .ZN(n5259) );
  INV_X1 U6280 ( .A(n8948), .ZN(n8951) );
  NAND2_X1 U6281 ( .A1(n5528), .A2(n5527), .ZN(n6053) );
  NAND2_X1 U6282 ( .A1(n5915), .A2(n5632), .ZN(n5937) );
  NAND2_X1 U6283 ( .A1(n8952), .A2(n5523), .ZN(n8953) );
  NOR2_X1 U6284 ( .A1(n5859), .A2(n5368), .ZN(n5367) );
  NAND2_X1 U6285 ( .A1(n5548), .A2(n5547), .ZN(n5546) );
  AOI21_X1 U6286 ( .B1(n6220), .B2(n5542), .A(n5541), .ZN(n5538) );
  INV_X1 U6287 ( .A(n5538), .ZN(n6268) );
  NAND2_X1 U6288 ( .A1(n8261), .A2(n8926), .ZN(n8417) );
  OAI21_X1 U6289 ( .B1(n5467), .B2(n10935), .A(n5131), .ZN(n8639) );
  NAND3_X1 U6290 ( .A1(n8544), .A2(n5136), .A3(n8836), .ZN(n5133) );
  NAND2_X4 U6291 ( .A1(n6975), .A2(n7287), .ZN(n7306) );
  AND2_X1 U6292 ( .A1(n5138), .A2(n8260), .ZN(n5140) );
  NAND3_X1 U6293 ( .A1(n5143), .A2(n8925), .A3(n5144), .ZN(n5138) );
  NAND2_X1 U6294 ( .A1(n9888), .A2(n5139), .ZN(n5141) );
  INV_X1 U6295 ( .A(n9347), .ZN(n5145) );
  OAI21_X1 U6296 ( .B1(n5145), .B2(n5102), .A(n5051), .ZN(n9306) );
  INV_X1 U6297 ( .A(n8917), .ZN(n5148) );
  NAND2_X1 U6298 ( .A1(n5149), .A2(n5101), .ZN(n5150) );
  OR2_X1 U6299 ( .A1(n9269), .A2(n5156), .ZN(n5149) );
  NAND2_X1 U6300 ( .A1(n8773), .A2(n5100), .ZN(n5151) );
  NAND3_X1 U6301 ( .A1(n5151), .A2(n8782), .A3(n5150), .ZN(n8778) );
  AOI21_X1 U6302 ( .B1(n9269), .B2(n8907), .A(n5157), .ZN(n8772) );
  NAND2_X1 U6303 ( .A1(n5161), .A2(n5093), .ZN(n8758) );
  NAND2_X1 U6304 ( .A1(n5454), .A2(n5455), .ZN(n5160) );
  AND3_X1 U6305 ( .A1(n6449), .A2(n6615), .A3(n5474), .ZN(n6475) );
  AND3_X2 U6306 ( .A1(n5229), .A2(n5164), .A3(n5619), .ZN(n6615) );
  NAND3_X1 U6307 ( .A1(n6449), .A2(n5474), .A3(n5089), .ZN(n6451) );
  NAND2_X1 U6308 ( .A1(n5176), .A2(n5092), .ZN(n8618) );
  NAND3_X1 U6309 ( .A1(n10845), .A2(n7905), .A3(n7903), .ZN(n5177) );
  NAND2_X1 U6310 ( .A1(n5177), .A2(n5178), .ZN(n8080) );
  NAND4_X1 U6311 ( .A1(n5184), .A2(n5183), .A3(n5645), .A4(n5586), .ZN(n5182)
         );
  NAND2_X1 U6312 ( .A1(n5184), .A2(n5185), .ZN(n5644) );
  NOR2_X1 U6313 ( .A1(n5520), .A2(n5522), .ZN(n6409) );
  MUX2_X1 U6314 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n7275), .S(n7430), .Z(n10661)
         );
  NAND3_X1 U6315 ( .A1(n5203), .A2(n9235), .A3(n9234), .ZN(n5202) );
  NAND2_X1 U6316 ( .A1(n5613), .A2(n5614), .ZN(n8538) );
  INV_X1 U6317 ( .A(n8932), .ZN(n5213) );
  OAI21_X1 U6318 ( .B1(n10801), .B2(n10808), .A(n5216), .ZN(n9899) );
  NAND2_X1 U6319 ( .A1(n10764), .A2(n8258), .ZN(n10765) );
  INV_X1 U6320 ( .A(n9899), .ZN(n8253) );
  AOI21_X1 U6321 ( .B1(n5218), .B2(n5221), .A(n5103), .ZN(n5217) );
  INV_X1 U6322 ( .A(n5221), .ZN(n5219) );
  NAND2_X1 U6323 ( .A1(n8454), .A2(n8255), .ZN(n10890) );
  INV_X1 U6324 ( .A(n10895), .ZN(n5225) );
  MUX2_X1 U6325 ( .A(P2_IR_REG_0__SCAN_IN), .B(n10014), .S(n7306), .Z(n10707)
         );
  NAND2_X1 U6326 ( .A1(n5236), .A2(n5237), .ZN(n5240) );
  OR2_X1 U6327 ( .A1(n8880), .A2(n5245), .ZN(n5236) );
  NAND2_X1 U6328 ( .A1(n8879), .A2(n5096), .ZN(n5241) );
  NAND3_X1 U6329 ( .A1(n5241), .A2(n9345), .A3(n5240), .ZN(n8887) );
  AND2_X1 U6330 ( .A1(n5241), .A2(n5240), .ZN(n8889) );
  NAND2_X1 U6331 ( .A1(n5246), .A2(n5247), .ZN(n8858) );
  NAND2_X1 U6332 ( .A1(n8833), .A2(n5248), .ZN(n5246) );
  NAND2_X1 U6333 ( .A1(n8843), .A2(n8844), .ZN(n5251) );
  NAND3_X1 U6334 ( .A1(n8814), .A2(n8815), .A3(n9900), .ZN(n5256) );
  NAND2_X1 U6335 ( .A1(n5265), .A2(n5266), .ZN(n8874) );
  NAND2_X1 U6336 ( .A1(n8866), .A2(n5268), .ZN(n5265) );
  NAND3_X1 U6337 ( .A1(n5278), .A2(n6463), .A3(n6615), .ZN(n6465) );
  MUX2_X1 U6338 ( .A(n8803), .B(n8802), .S(n8912), .Z(n8807) );
  AND2_X2 U6339 ( .A1(n8786), .A2(n8785), .ZN(n8912) );
  NAND2_X1 U6340 ( .A1(n5739), .A2(n5738), .ZN(n5283) );
  OAI21_X1 U6341 ( .B1(n5764), .B2(n5365), .A(n5796), .ZN(n5282) );
  NAND2_X1 U6342 ( .A1(n5302), .A2(n5301), .ZN(n8970) );
  INV_X1 U6343 ( .A(n5959), .ZN(n5322) );
  AND3_X2 U6344 ( .A1(n5324), .A2(n5323), .A3(n5771), .ZN(n5637) );
  NAND2_X2 U6345 ( .A1(n5328), .A2(n5327), .ZN(n7216) );
  INV_X1 U6346 ( .A(n5337), .ZN(n10376) );
  INV_X1 U6347 ( .A(n9362), .ZN(n5341) );
  NAND2_X1 U6348 ( .A1(n5343), .A2(n5341), .ZN(n9300) );
  INV_X1 U6349 ( .A(n10933), .ZN(n5349) );
  NAND2_X1 U6350 ( .A1(n5349), .A2(n5350), .ZN(n8641) );
  NAND2_X1 U6351 ( .A1(n5836), .A2(n5835), .ZN(n5371) );
  NAND2_X1 U6352 ( .A1(n5836), .A2(n5367), .ZN(n5366) );
  INV_X1 U6353 ( .A(n5835), .ZN(n5368) );
  XNOR2_X1 U6354 ( .A(n10273), .B(n7139), .ZN(n5376) );
  OAI211_X1 U6355 ( .C1(n10453), .C2(n11091), .A(n5377), .B(n5374), .ZN(
        P1_U3552) );
  OR2_X1 U6356 ( .A1(n11093), .A2(n6421), .ZN(n5377) );
  NAND2_X1 U6357 ( .A1(n5392), .A2(n5099), .ZN(n10425) );
  NOR2_X1 U6358 ( .A1(n10294), .A2(n8990), .ZN(n8991) );
  NAND2_X1 U6359 ( .A1(n8513), .A2(n8528), .ZN(n8602) );
  NAND2_X1 U6360 ( .A1(n8618), .A2(n8617), .ZN(n8974) );
  NAND2_X1 U6361 ( .A1(n7555), .A2(n7005), .ZN(n5942) );
  NAND2_X1 U6362 ( .A1(n5824), .A2(n5823), .ZN(n5836) );
  NAND2_X1 U6363 ( .A1(n7745), .A2(n7024), .ZN(n7220) );
  AND4_X2 U6364 ( .A1(n5640), .A2(n5639), .A3(n5638), .A4(n9785), .ZN(n5631)
         );
  NAND2_X1 U6365 ( .A1(n6495), .A2(n5698), .ZN(n5716) );
  NAND2_X1 U6366 ( .A1(n9051), .A2(n6500), .ZN(n8000) );
  NAND2_X1 U6367 ( .A1(n8043), .A2(n5395), .ZN(n5394) );
  INV_X1 U6368 ( .A(n6516), .ZN(n5395) );
  NAND4_X1 U6369 ( .A1(n5397), .A2(n6500), .A3(n8043), .A4(n9051), .ZN(n5396)
         );
  NAND2_X1 U6370 ( .A1(n7949), .A2(n6599), .ZN(n5399) );
  NAND2_X1 U6371 ( .A1(n8232), .A2(n6646), .ZN(n5402) );
  NAND2_X1 U6372 ( .A1(n6751), .A2(n6466), .ZN(n5405) );
  NAND2_X1 U6373 ( .A1(n5404), .A2(n5403), .ZN(n6472) );
  NAND2_X1 U6374 ( .A1(n6751), .A2(n5406), .ZN(n5404) );
  NAND2_X1 U6375 ( .A1(n5414), .A2(n5416), .ZN(n6717) );
  NAND2_X1 U6376 ( .A1(n6687), .A2(n5417), .ZN(n5414) );
  NAND2_X1 U6377 ( .A1(n6687), .A2(n8715), .ZN(n8748) );
  OR2_X1 U6378 ( .A1(n6731), .A2(n5423), .ZN(n5419) );
  NAND2_X1 U6379 ( .A1(n5419), .A2(n5420), .ZN(n9120) );
  NAND2_X1 U6380 ( .A1(n8201), .A2(n9846), .ZN(n5426) );
  NOR2_X1 U6381 ( .A1(n6947), .A2(n5426), .ZN(n5427) );
  NAND2_X1 U6382 ( .A1(n8780), .A2(n5429), .ZN(n5428) );
  OAI21_X1 U6383 ( .B1(n9027), .B2(n5434), .A(n5431), .ZN(n6808) );
  NAND2_X1 U6384 ( .A1(n9109), .A2(n5040), .ZN(n5440) );
  NAND2_X1 U6385 ( .A1(n5440), .A2(n5441), .ZN(n9137) );
  INV_X1 U6386 ( .A(n8211), .ZN(n5453) );
  INV_X1 U6387 ( .A(n8680), .ZN(n5454) );
  INV_X1 U6388 ( .A(n8543), .ZN(n5467) );
  NAND2_X1 U6389 ( .A1(n10773), .A2(n5471), .ZN(n5470) );
  AND2_X1 U6390 ( .A1(n6441), .A2(n5104), .ZN(n5474) );
  INV_X1 U6391 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5483) );
  INV_X1 U6392 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5482) );
  AND3_X2 U6393 ( .A1(n9558), .A2(n5483), .A3(n5482), .ZN(n5772) );
  OAI21_X1 U6394 ( .B1(n8017), .B2(n8018), .A(n5908), .ZN(n5933) );
  NAND2_X1 U6395 ( .A1(n8017), .A2(n5908), .ZN(n5486) );
  NAND2_X1 U6396 ( .A1(n5489), .A2(n5487), .ZN(n6191) );
  NAND2_X1 U6397 ( .A1(n6161), .A2(n6160), .ZN(n5489) );
  AOI21_X1 U6398 ( .B1(n5493), .B2(n6038), .A(n5492), .ZN(n5491) );
  INV_X1 U6399 ( .A(n8656), .ZN(n5492) );
  NAND2_X1 U6400 ( .A1(n5494), .A2(n6038), .ZN(n8653) );
  NAND2_X1 U6401 ( .A1(n10037), .A2(n10036), .ZN(n5495) );
  NAND2_X1 U6402 ( .A1(n5495), .A2(n5091), .ZN(n10103) );
  NAND2_X1 U6403 ( .A1(n8220), .A2(n5044), .ZN(n5499) );
  NAND2_X1 U6404 ( .A1(n5499), .A2(n5500), .ZN(n8555) );
  OAI21_X1 U6405 ( .B1(n5504), .B2(n7665), .A(n7676), .ZN(n5503) );
  NAND2_X1 U6406 ( .A1(n10083), .A2(n5510), .ZN(n5509) );
  NAND2_X1 U6407 ( .A1(n6088), .A2(n5514), .ZN(n5513) );
  NAND2_X1 U6408 ( .A1(n5513), .A2(n5515), .ZN(n10027) );
  NAND2_X1 U6409 ( .A1(n5554), .A2(n5631), .ZN(n5520) );
  AND2_X1 U6410 ( .A1(n5631), .A2(n9591), .ZN(n5521) );
  NAND2_X1 U6411 ( .A1(n6019), .A2(n5530), .ZN(n5528) );
  NAND2_X1 U6412 ( .A1(n6195), .A2(n6194), .ZN(n6220) );
  NAND2_X1 U6413 ( .A1(n6195), .A2(n5536), .ZN(n5535) );
  NAND2_X1 U6414 ( .A1(n6090), .A2(n5551), .ZN(n6114) );
  INV_X1 U6415 ( .A(n6111), .ZN(n5553) );
  NAND3_X1 U6416 ( .A1(n5671), .A2(n5670), .A3(n5672), .ZN(n5698) );
  AND2_X2 U6417 ( .A1(n5772), .A2(n9587), .ZN(n5554) );
  NAND3_X1 U6418 ( .A1(n5637), .A2(n5772), .A3(n5636), .ZN(n5967) );
  INV_X1 U6419 ( .A(n5562), .ZN(n5561) );
  OAI22_X1 U6420 ( .A1(n5763), .A2(n7422), .B1(n7470), .B2(n7478), .ZN(n5562)
         );
  NAND2_X1 U6421 ( .A1(n10404), .A2(n5564), .ZN(n5563) );
  NAND2_X1 U6422 ( .A1(n8631), .A2(n8960), .ZN(n5576) );
  INV_X1 U6423 ( .A(n8960), .ZN(n5577) );
  NAND2_X1 U6424 ( .A1(n5578), .A2(n8630), .ZN(n10509) );
  INV_X1 U6425 ( .A(n5580), .ZN(n5579) );
  INV_X1 U6426 ( .A(n5584), .ZN(n5582) );
  NAND2_X1 U6427 ( .A1(n6409), .A2(n5588), .ZN(n5655) );
  INV_X1 U6428 ( .A(n6482), .ZN(n8697) );
  INV_X1 U6429 ( .A(n9359), .ZN(n5594) );
  NOR2_X1 U6430 ( .A1(n9359), .A2(n9255), .ZN(n9340) );
  NOR2_X1 U6431 ( .A1(n5593), .A2(n9255), .ZN(n5592) );
  NAND2_X1 U6432 ( .A1(n9316), .A2(n5598), .ZN(n5595) );
  NAND2_X1 U6433 ( .A1(n5595), .A2(n5596), .ZN(n9284) );
  NAND2_X1 U6434 ( .A1(n9316), .A2(n9319), .ZN(n5597) );
  INV_X1 U6435 ( .A(n5602), .ZN(n9854) );
  AOI21_X1 U6436 ( .B1(n8677), .B2(n5605), .A(n5603), .ZN(n5602) );
  INV_X1 U6437 ( .A(n8935), .ZN(n5604) );
  NAND2_X1 U6438 ( .A1(n8426), .A2(n5615), .ZN(n5613) );
  INV_X1 U6439 ( .A(n8426), .ZN(n8537) );
  NAND2_X1 U6440 ( .A1(n9898), .A2(n5617), .ZN(n8454) );
  NAND2_X1 U6441 ( .A1(n6923), .A2(n6450), .ZN(n6919) );
  NAND3_X1 U6442 ( .A1(n5679), .A2(n5624), .A3(n5678), .ZN(n7629) );
  OR2_X1 U6443 ( .A1(n7021), .A2(n6341), .ZN(n5678) );
  NOR2_X2 U6444 ( .A1(n7119), .A2(n7021), .ZN(n7714) );
  NAND2_X1 U6445 ( .A1(n9053), .A2(n5067), .ZN(n9051) );
  AND2_X1 U6446 ( .A1(n8955), .A2(n7285), .ZN(n7817) );
  INV_X1 U6447 ( .A(n9846), .ZN(n10902) );
  NAND2_X1 U6448 ( .A1(n6326), .A2(n6325), .ZN(n6349) );
  INV_X1 U6449 ( .A(n6326), .ZN(n6323) );
  OAI21_X1 U6450 ( .B1(n6318), .B2(n6317), .A(n6316), .ZN(n6326) );
  XNOR2_X1 U6451 ( .A(n6318), .B(n6317), .ZN(n8593) );
  INV_X1 U6452 ( .A(n5806), .ZN(n5809) );
  INV_X1 U6453 ( .A(n5879), .ZN(n5882) );
  NAND2_X1 U6454 ( .A1(n7763), .A2(n7762), .ZN(n7767) );
  OR2_X1 U6455 ( .A1(n10999), .A2(n11007), .ZN(n10997) );
  NAND2_X1 U6456 ( .A1(n10001), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U6457 ( .A1(n10001), .A2(n6479), .ZN(n6480) );
  NAND2_X1 U6458 ( .A1(n6475), .A2(n5045), .ZN(n10001) );
  NAND2_X1 U6459 ( .A1(n5655), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5656) );
  INV_X1 U6460 ( .A(n7101), .ZN(n6422) );
  NAND2_X1 U6461 ( .A1(n7101), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5695) );
  INV_X1 U6462 ( .A(n9161), .ZN(n7827) );
  AND2_X2 U6463 ( .A1(n10008), .A2(n6482), .ZN(n6549) );
  NAND2_X1 U6464 ( .A1(n6424), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5653) );
  INV_X1 U6465 ( .A(n5650), .ZN(n8709) );
  NAND2_X1 U6466 ( .A1(n8194), .A2(n9050), .ZN(n8798) );
  NAND2_X1 U6467 ( .A1(n5715), .A2(n5714), .ZN(n5718) );
  OAI21_X1 U6468 ( .B1(n5768), .B2(n7421), .A(n5699), .ZN(n5714) );
  BUF_X4 U6469 ( .A(n5768), .Z(n6995) );
  OR2_X1 U6470 ( .A1(n7497), .A2(n5666), .ZN(n5624) );
  NAND2_X1 U6471 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5625) );
  AND2_X1 U6472 ( .A1(n9982), .A2(n9248), .ZN(n5626) );
  OR2_X1 U6473 ( .A1(n10465), .A2(n10052), .ZN(n5627) );
  AND4_X1 U6474 ( .A1(n9290), .A2(n8763), .A3(n9331), .A4(n8943), .ZN(n5628)
         );
  AND3_X1 U6475 ( .A1(n9812), .A2(n9808), .A3(n9813), .ZN(n5629) );
  AND2_X1 U6476 ( .A1(n5936), .A2(n5914), .ZN(n5632) );
  AND2_X1 U6477 ( .A1(n6018), .A2(n5992), .ZN(n5633) );
  INV_X1 U6478 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10534) );
  OR2_X1 U6479 ( .A1(n7713), .A2(n7712), .ZN(n11013) );
  NAND2_X1 U6480 ( .A1(n7212), .A2(n7250), .ZN(n10272) );
  INV_X1 U6481 ( .A(n10283), .ZN(n10255) );
  INV_X1 U6482 ( .A(n9307), .ZN(n8763) );
  NAND2_X1 U6483 ( .A1(n10929), .A2(n10931), .ZN(n10930) );
  NAND2_X1 U6484 ( .A1(n10050), .A2(n10049), .ZN(n5634) );
  NOR2_X1 U6485 ( .A1(n8611), .A2(n10514), .ZN(n8610) );
  AND2_X1 U6486 ( .A1(n8780), .A2(n8779), .ZN(n5635) );
  AND2_X1 U6487 ( .A1(n8779), .A2(n8950), .ZN(n10811) );
  INV_X1 U6488 ( .A(n10811), .ZN(n10942) );
  INV_X1 U6489 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9797) );
  NOR2_X1 U6490 ( .A1(n8784), .A2(n8783), .ZN(n8944) );
  INV_X1 U6491 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9807) );
  INV_X1 U6492 ( .A(n6667), .ZN(n6666) );
  INV_X1 U6493 ( .A(n6711), .ZN(n6710) );
  INV_X1 U6494 ( .A(n5880), .ZN(n5881) );
  INV_X1 U6495 ( .A(n6251), .ZN(n6249) );
  INV_X1 U6496 ( .A(n6332), .ZN(n6330) );
  INV_X1 U6497 ( .A(n8086), .ZN(n8087) );
  INV_X1 U6498 ( .A(n6828), .ZN(n6827) );
  INV_X1 U6499 ( .A(n9050), .ZN(n8193) );
  INV_X1 U6500 ( .A(n6850), .ZN(n6841) );
  INV_X1 U6501 ( .A(n6741), .ZN(n6739) );
  NAND2_X1 U6502 ( .A1(n9356), .A2(n8762), .ZN(n9347) );
  INV_X1 U6503 ( .A(n6773), .ZN(n6771) );
  OR2_X1 U6504 ( .A1(n6755), .A2(n6754), .ZN(n6773) );
  INV_X1 U6505 ( .A(n9900), .ZN(n8252) );
  INV_X1 U6506 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U6507 ( .A1(n7216), .A2(n6373), .ZN(n5701) );
  NAND2_X1 U6508 ( .A1(n5882), .A2(n5881), .ZN(n8127) );
  NAND2_X1 U6509 ( .A1(n6249), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6275) );
  INV_X1 U6510 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U6511 ( .A1(n6330), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6376) );
  INV_X1 U6512 ( .A(n8607), .ZN(n8604) );
  OR2_X1 U6513 ( .A1(n6990), .A2(n6989), .ZN(n6991) );
  INV_X1 U6514 ( .A(n6133), .ZN(n6134) );
  INV_X1 U6515 ( .A(SI_10_), .ZN(n9644) );
  INV_X1 U6516 ( .A(n6869), .ZN(n6868) );
  NAND2_X1 U6517 ( .A1(n6827), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6850) );
  INV_X1 U6518 ( .A(n9158), .ZN(n8189) );
  NAND2_X1 U6519 ( .A1(n6786), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6799) );
  OR2_X1 U6520 ( .A1(n6852), .A2(n6842), .ZN(n6869) );
  NAND2_X1 U6521 ( .A1(n6739), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6755) );
  NAND2_X1 U6522 ( .A1(n6771), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6787) );
  INV_X1 U6523 ( .A(n7306), .ZN(n6767) );
  AND2_X1 U6524 ( .A1(n8824), .A2(n8825), .ZN(n10895) );
  NAND2_X1 U6525 ( .A1(n8196), .A2(n8195), .ZN(n8238) );
  OR2_X1 U6526 ( .A1(n7629), .A2(n5686), .ZN(n5692) );
  INV_X1 U6527 ( .A(n10038), .ZN(n6211) );
  INV_X1 U6528 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U6529 ( .A1(n6174), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6198) );
  INV_X1 U6530 ( .A(n5729), .ZN(n5730) );
  NOR2_X1 U6531 ( .A1(n6027), .A2(n8658), .ZN(n6070) );
  OR2_X1 U6532 ( .A1(n6376), .A2(n6375), .ZN(n6418) );
  INV_X1 U6533 ( .A(n6424), .ZN(n6334) );
  OR2_X1 U6534 ( .A1(n6198), .A2(n10042), .ZN(n6226) );
  INV_X1 U6535 ( .A(n7768), .ZN(n7764) );
  NAND2_X1 U6536 ( .A1(n7003), .A2(n6994), .ZN(n6998) );
  NAND2_X1 U6537 ( .A1(n6349), .A2(n6348), .ZN(n6365) );
  INV_X1 U6538 ( .A(SI_17_), .ZN(n9636) );
  NAND2_X1 U6539 ( .A1(n5990), .A2(n5989), .ZN(n6018) );
  INV_X1 U6540 ( .A(n9260), .ZN(n9308) );
  INV_X1 U6541 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9672) );
  INV_X1 U6542 ( .A(n9863), .ZN(n9251) );
  INV_X1 U6543 ( .A(n9129), .ZN(n9141) );
  AND2_X1 U6544 ( .A1(n8198), .A2(n6943), .ZN(n6974) );
  INV_X1 U6545 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U6546 ( .A1(n7827), .A2(n10707), .ZN(n8273) );
  INV_X1 U6547 ( .A(n9890), .ZN(n10939) );
  AND2_X1 U6548 ( .A1(n8955), .A2(n10706), .ZN(n10975) );
  AOI21_X1 U6549 ( .B1(n10546), .B2(n10548), .A(n10549), .ZN(n7820) );
  XNOR2_X1 U6550 ( .A(n5703), .B(n5686), .ZN(n7593) );
  AND3_X1 U6551 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U6552 ( .A1(n5809), .A2(n5808), .ZN(n7729) );
  AND2_X1 U6553 ( .A1(n7716), .A2(n7718), .ZN(n7271) );
  OAI21_X1 U6554 ( .B1(n7260), .B2(n7717), .A(n7259), .ZN(n7261) );
  INV_X1 U6555 ( .A(n10865), .ZN(n11025) );
  OR2_X1 U6556 ( .A1(n10741), .A2(n7718), .ZN(n7575) );
  AND2_X1 U6557 ( .A1(n7705), .A2(n7580), .ZN(n10739) );
  AND2_X1 U6558 ( .A1(n8529), .A2(n8528), .ZN(n11060) );
  INV_X1 U6559 ( .A(n10169), .ZN(n8226) );
  OR2_X1 U6560 ( .A1(n7578), .A2(n7596), .ZN(n7694) );
  XNOR2_X1 U6561 ( .A(n6112), .B(n9636), .ZN(n6111) );
  INV_X1 U6562 ( .A(SI_6_), .ZN(n9655) );
  NAND2_X1 U6563 ( .A1(n5768), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5699) );
  OR3_X1 U6564 ( .A1(n8462), .A2(n8597), .A3(n8652), .ZN(n7274) );
  NAND2_X1 U6565 ( .A1(n9135), .A2(n8780), .ZN(n9122) );
  OR2_X1 U6566 ( .A1(n9080), .A2(n10937), .ZN(n9104) );
  OR2_X1 U6567 ( .A1(n7824), .A2(n6975), .ZN(n10937) );
  AND2_X1 U6568 ( .A1(n6858), .A2(n6857), .ZN(n9092) );
  AND4_X1 U6569 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n8670)
         );
  NAND2_X1 U6570 ( .A1(n7308), .A2(n7307), .ZN(n9217) );
  INV_X1 U6571 ( .A(n10673), .ZN(n10649) );
  INV_X1 U6572 ( .A(n10937), .ZN(n9892) );
  OR2_X1 U6573 ( .A1(n10547), .A2(n7818), .ZN(n9849) );
  AND2_X1 U6574 ( .A1(n10644), .A2(n6930), .ZN(n8198) );
  INV_X1 U6575 ( .A(n11074), .ZN(n11034) );
  AND3_X1 U6576 ( .A1(n6488), .A2(n10902), .A3(n8785), .ZN(n10948) );
  INV_X1 U6577 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6706) );
  INV_X1 U6578 ( .A(n7261), .ZN(n7262) );
  AND2_X1 U6579 ( .A1(n6309), .A2(n6308), .ZN(n10340) );
  OR2_X1 U6580 ( .A1(n7494), .A2(n7493), .ZN(n7562) );
  OR2_X1 U6581 ( .A1(n10186), .A2(n10187), .ZN(n10188) );
  INV_X1 U6582 ( .A(n10695), .ZN(n10635) );
  INV_X1 U6583 ( .A(n10849), .ZN(n11006) );
  AND2_X1 U6584 ( .A1(n7233), .A2(n7231), .ZN(n7806) );
  AOI21_X1 U6585 ( .B1(n6407), .B2(n9817), .A(n7440), .ZN(n7702) );
  AND2_X1 U6586 ( .A1(n11013), .A2(n10741), .ZN(n11059) );
  OR2_X1 U6587 ( .A1(n7110), .A2(n7717), .ZN(n10741) );
  NOR2_X1 U6588 ( .A1(n7579), .A2(n7694), .ZN(n7588) );
  AND2_X1 U6589 ( .A1(n6095), .A2(n6115), .ZN(n10227) );
  INV_X1 U6590 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n8340) );
  NOR2_X1 U6591 ( .A1(n10574), .A2(n10573), .ZN(n8366) );
  INV_X1 U6592 ( .A(n9217), .ZN(n10672) );
  NOR2_X1 U6593 ( .A1(n6979), .A2(n6978), .ZN(n6980) );
  INV_X1 U6594 ( .A(n9098), .ZN(n9146) );
  NAND2_X1 U6595 ( .A1(n6876), .A2(n6875), .ZN(n9260) );
  OR2_X1 U6596 ( .A1(n6779), .A2(n6778), .ZN(n9863) );
  INV_X1 U6597 ( .A(n10684), .ZN(n10653) );
  NAND2_X1 U6598 ( .A1(n10957), .A2(n10899), .ZN(n10956) );
  INV_X2 U6599 ( .A(n10957), .ZN(n10906) );
  INV_X1 U6600 ( .A(n11078), .ZN(n11076) );
  INV_X1 U6601 ( .A(n11082), .ZN(n11079) );
  OR2_X1 U6602 ( .A1(n10547), .A2(n10546), .ZN(n10645) );
  AND2_X1 U6603 ( .A1(n7283), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10648) );
  INV_X1 U6604 ( .A(n6947), .ZN(n8785) );
  INV_X1 U6605 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7661) );
  INV_X1 U6606 ( .A(n10476), .ZN(n10347) );
  INV_X1 U6607 ( .A(n10131), .ZN(n10156) );
  INV_X1 U6608 ( .A(n10340), .ZN(n10158) );
  INV_X1 U6609 ( .A(n10401), .ZN(n10164) );
  OR2_X1 U6610 ( .A1(P1_U3083), .A2(n7498), .ZN(n10631) );
  OR2_X1 U6611 ( .A1(n10593), .A2(n10590), .ZN(n10695) );
  INV_X1 U6612 ( .A(n11093), .ZN(n11091) );
  INV_X1 U6613 ( .A(n11097), .ZN(n11094) );
  AND2_X2 U6614 ( .A1(n7588), .A2(n7695), .ZN(n11097) );
  INV_X1 U6615 ( .A(n5649), .ZN(n8696) );
  INV_X1 U6616 ( .A(n7716), .ZN(n8291) );
  INV_X1 U6617 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7627) );
  NOR2_X1 U6618 ( .A1(n8367), .A2(n8366), .ZN(n10576) );
  AND2_X1 U6619 ( .A1(n7282), .A2(n10648), .ZN(P2_U3966) );
  INV_X1 U6620 ( .A(n10176), .ZN(P1_U4006) );
  NOR2_X1 U6621 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5640) );
  NOR2_X1 U6622 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5639) );
  NOR2_X1 U6623 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5638) );
  INV_X1 U6624 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9812) );
  INV_X1 U6625 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9813) );
  INV_X1 U6626 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9605) );
  XNOR2_X2 U6627 ( .A(n5643), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U6628 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5645) );
  AND2_X4 U6629 ( .A1(n8709), .A2(n5649), .ZN(n7101) );
  NAND2_X1 U6630 ( .A1(n7101), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5654) );
  AND2_X4 U6631 ( .A1(n5649), .A2(n5650), .ZN(n6424) );
  NAND2_X1 U6632 ( .A1(n5790), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U6633 ( .A1(n5758), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5651) );
  NAND4_X2 U6634 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), .ZN(n7119)
         );
  NAND2_X2 U6635 ( .A1(n5660), .A2(n5657), .ZN(n8594) );
  XNOR2_X1 U6636 ( .A(n5659), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U6637 ( .A1(n5050), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U6638 ( .A1(n5664), .A2(n5663), .ZN(n5662) );
  XNOR2_X1 U6639 ( .A(n5664), .B(n5663), .ZN(n8040) );
  NAND2_X1 U6640 ( .A1(n7718), .A2(n8040), .ZN(n7710) );
  INV_X1 U6641 ( .A(n7710), .ZN(n5665) );
  NAND2_X1 U6642 ( .A1(n7119), .A2(n6388), .ZN(n5679) );
  INV_X1 U6643 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5666) );
  INV_X1 U6644 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10633) );
  AND2_X1 U6645 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5672) );
  INV_X1 U6646 ( .A(SI_0_), .ZN(n5674) );
  INV_X1 U6647 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5673) );
  OAI21_X1 U6648 ( .B1(n6995), .B2(n5674), .A(n5673), .ZN(n5675) );
  NAND2_X1 U6649 ( .A1(n5698), .A2(n5675), .ZN(n10540) );
  XNOR2_X2 U6650 ( .A(n5676), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6416) );
  MUX2_X1 U6651 ( .A(n10633), .B(n10540), .S(n7470), .Z(n7021) );
  AND2_X4 U6652 ( .A1(n7710), .A2(n7497), .ZN(n6373) );
  NAND2_X1 U6653 ( .A1(n5680), .A2(n9796), .ZN(n5681) );
  NAND2_X1 U6654 ( .A1(n5681), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U6655 ( .A1(n5683), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5684) );
  INV_X1 U6656 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9587) );
  XNOR2_X2 U6657 ( .A(n5684), .B(n9587), .ZN(n10392) );
  NAND2_X1 U6658 ( .A1(n7716), .A2(n10392), .ZN(n5685) );
  NAND2_X2 U6659 ( .A1(n7710), .A2(n5685), .ZN(n6342) );
  NAND2_X1 U6660 ( .A1(n8040), .A2(n10392), .ZN(n7580) );
  OR2_X1 U6661 ( .A1(n7716), .A2(n7580), .ZN(n5687) );
  NAND2_X1 U6662 ( .A1(n7119), .A2(n5031), .ZN(n5691) );
  OR2_X1 U6663 ( .A1(n7021), .A2(n6384), .ZN(n5690) );
  OR2_X1 U6664 ( .A1(n7497), .A2(n10633), .ZN(n5689) );
  AND3_X1 U6665 ( .A1(n5691), .A2(n5690), .A3(n5689), .ZN(n7630) );
  NAND2_X1 U6666 ( .A1(n7630), .A2(n7629), .ZN(n7628) );
  NAND2_X1 U6667 ( .A1(n6424), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U6668 ( .A1(n5790), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U6669 ( .A1(n5758), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U6670 ( .A1(n5704), .A2(n6388), .ZN(n5702) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7421) );
  AND2_X1 U6672 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U6673 ( .A1(n5768), .A2(n5697), .ZN(n6495) );
  INV_X1 U6674 ( .A(SI_1_), .ZN(n9462) );
  XNOR2_X1 U6675 ( .A(n5716), .B(n9462), .ZN(n5715) );
  XNOR2_X1 U6676 ( .A(n5715), .B(n5714), .ZN(n7431) );
  INV_X1 U6677 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9759) );
  NAND2_X1 U6678 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5700) );
  XNOR2_X1 U6679 ( .A(n9759), .B(n5700), .ZN(n10625) );
  NAND2_X1 U6680 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  NAND2_X1 U6681 ( .A1(n7592), .A2(n7593), .ZN(n5707) );
  NAND2_X1 U6682 ( .A1(n5704), .A2(n6063), .ZN(n5706) );
  NAND2_X1 U6683 ( .A1(n7216), .A2(n6388), .ZN(n5705) );
  NAND2_X1 U6684 ( .A1(n5706), .A2(n5705), .ZN(n7591) );
  NAND2_X1 U6685 ( .A1(n5707), .A2(n7591), .ZN(n5711) );
  INV_X1 U6686 ( .A(n7592), .ZN(n5709) );
  INV_X1 U6687 ( .A(n7593), .ZN(n5708) );
  NAND2_X1 U6688 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  NAND2_X1 U6689 ( .A1(n5711), .A2(n5710), .ZN(n7652) );
  INV_X1 U6690 ( .A(n7652), .ZN(n5734) );
  OR2_X1 U6691 ( .A1(n5712), .A2(n10534), .ZN(n5713) );
  XNOR2_X1 U6692 ( .A(n5713), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10691) );
  INV_X1 U6693 ( .A(n10691), .ZN(n7478) );
  NAND2_X1 U6694 ( .A1(n5716), .A2(SI_1_), .ZN(n5717) );
  NAND2_X1 U6695 ( .A1(n5718), .A2(n5717), .ZN(n5739) );
  MUX2_X1 U6696 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n5768), .Z(n5740) );
  INV_X1 U6697 ( .A(SI_2_), .ZN(n5719) );
  XNOR2_X1 U6698 ( .A(n5740), .B(n5719), .ZN(n5738) );
  XNOR2_X1 U6699 ( .A(n5739), .B(n5738), .ZN(n7422) );
  NAND2_X1 U6700 ( .A1(n7024), .A2(n6373), .ZN(n5725) );
  NAND2_X1 U6701 ( .A1(n6424), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U6702 ( .A1(n7101), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U6703 ( .A1(n5790), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U6704 ( .A1(n5758), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U6705 ( .A1(n5727), .A2(n6388), .ZN(n5724) );
  NAND2_X1 U6706 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  XNOR2_X1 U6707 ( .A(n5726), .B(n5686), .ZN(n5728) );
  AOI22_X1 U6708 ( .A1(n5727), .A2(n6063), .B1(n6388), .B2(n7024), .ZN(n5729)
         );
  NAND2_X1 U6709 ( .A1(n5728), .A2(n5729), .ZN(n5735) );
  INV_X1 U6710 ( .A(n5728), .ZN(n5731) );
  NAND2_X1 U6711 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  INV_X1 U6712 ( .A(n7653), .ZN(n5733) );
  NAND2_X1 U6713 ( .A1(n5734), .A2(n5733), .ZN(n7650) );
  NAND2_X1 U6714 ( .A1(n7650), .A2(n5735), .ZN(n7664) );
  OR3_X1 U6715 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_IR_REG_1__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U6716 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5736), .ZN(n5737) );
  XNOR2_X1 U6717 ( .A(n5737), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10610) );
  INV_X1 U6718 ( .A(n10610), .ZN(n7405) );
  NAND2_X1 U6719 ( .A1(n5740), .A2(SI_2_), .ZN(n5741) );
  INV_X1 U6720 ( .A(SI_3_), .ZN(n5742) );
  XNOR2_X1 U6721 ( .A(n5766), .B(n5742), .ZN(n5764) );
  XNOR2_X1 U6722 ( .A(n5765), .B(n5764), .ZN(n7409) );
  OR2_X1 U6723 ( .A1(n5763), .A2(n7409), .ZN(n5744) );
  OR2_X1 U6724 ( .A1(n7015), .A2(n5287), .ZN(n5743) );
  NAND2_X1 U6725 ( .A1(n10738), .A2(n6373), .ZN(n5751) );
  NAND2_X1 U6726 ( .A1(n7101), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5749) );
  INV_X1 U6727 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U6728 ( .A1(n6424), .A2(n5745), .ZN(n5748) );
  NAND2_X1 U6729 ( .A1(n5790), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U6730 ( .A1(n5758), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5746) );
  NAND4_X1 U6731 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n10175)
         );
  NAND2_X1 U6732 ( .A1(n10175), .A2(n6388), .ZN(n5750) );
  NAND2_X1 U6733 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  XNOR2_X1 U6734 ( .A(n5752), .B(n6342), .ZN(n5753) );
  AOI22_X1 U6735 ( .A1(n10175), .A2(n6063), .B1(n6388), .B2(n10738), .ZN(n5754) );
  XNOR2_X1 U6736 ( .A(n5753), .B(n5754), .ZN(n7665) );
  INV_X1 U6737 ( .A(n5753), .ZN(n5755) );
  NAND2_X1 U6738 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  NAND2_X1 U6739 ( .A1(n7101), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5762) );
  INV_X1 U6740 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5757) );
  XNOR2_X1 U6741 ( .A(n5757), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U6742 ( .A1(n6424), .A2(n7784), .ZN(n5761) );
  NAND2_X1 U6743 ( .A1(n6302), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U6744 ( .A1(n6303), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5759) );
  NAND4_X1 U6745 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n10174)
         );
  NAND2_X1 U6746 ( .A1(n10174), .A2(n6388), .ZN(n5781) );
  NAND2_X1 U6747 ( .A1(n5766), .A2(SI_3_), .ZN(n5767) );
  MUX2_X1 U6748 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n5768), .Z(n5798) );
  INV_X1 U6749 ( .A(SI_4_), .ZN(n5769) );
  XNOR2_X1 U6750 ( .A(n5798), .B(n5769), .ZN(n5796) );
  XNOR2_X1 U6751 ( .A(n5797), .B(n5796), .ZN(n7417) );
  OR2_X1 U6752 ( .A1(n5763), .A2(n7417), .ZN(n5779) );
  INV_X1 U6753 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5770) );
  OR2_X1 U6754 ( .A1(n7015), .A2(n5770), .ZN(n5778) );
  NAND2_X1 U6755 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  INV_X1 U6756 ( .A(n5817), .ZN(n5776) );
  NAND2_X1 U6757 ( .A1(n5773), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5774) );
  MUX2_X1 U6758 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5774), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5775) );
  NAND2_X1 U6759 ( .A1(n5776), .A2(n5775), .ZN(n7480) );
  OR2_X1 U6760 ( .A1(n7470), .A2(n7480), .ZN(n5777) );
  OR2_X1 U6761 ( .A1(n10758), .A2(n6341), .ZN(n5780) );
  NAND2_X1 U6762 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  XNOR2_X1 U6763 ( .A(n5782), .B(n5686), .ZN(n5785) );
  INV_X1 U6764 ( .A(n10758), .ZN(n7785) );
  NAND2_X1 U6765 ( .A1(n7785), .A2(n6388), .ZN(n5784) );
  NAND2_X1 U6766 ( .A1(n10174), .A2(n6063), .ZN(n5783) );
  AND2_X1 U6767 ( .A1(n5784), .A2(n5783), .ZN(n5786) );
  NAND2_X1 U6768 ( .A1(n5785), .A2(n5786), .ZN(n7677) );
  INV_X1 U6769 ( .A(n5785), .ZN(n5788) );
  INV_X1 U6770 ( .A(n5786), .ZN(n5787) );
  NAND2_X1 U6771 ( .A1(n5788), .A2(n5787), .ZN(n7676) );
  NAND2_X1 U6772 ( .A1(n7101), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5794) );
  AOI21_X1 U6773 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5789) );
  NOR2_X1 U6774 ( .A1(n5789), .A2(n5811), .ZN(n7770) );
  NAND2_X1 U6775 ( .A1(n6424), .A2(n7770), .ZN(n5793) );
  NAND2_X1 U6776 ( .A1(n6302), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U6777 ( .A1(n6303), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5791) );
  NAND4_X1 U6778 ( .A1(n5794), .A2(n5793), .A3(n5792), .A4(n5791), .ZN(n10173)
         );
  NAND2_X1 U6779 ( .A1(n10173), .A2(n6388), .ZN(n5804) );
  OR2_X1 U6780 ( .A1(n5817), .A2(n10534), .ZN(n5795) );
  XNOR2_X1 U6781 ( .A(n5795), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7532) );
  INV_X1 U6782 ( .A(n7532), .ZN(n7406) );
  NAND2_X1 U6783 ( .A1(n5798), .A2(SI_4_), .ZN(n5799) );
  MUX2_X1 U6784 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6995), .Z(n5822) );
  INV_X1 U6785 ( .A(SI_5_), .ZN(n5800) );
  XNOR2_X1 U6786 ( .A(n5822), .B(n5800), .ZN(n5820) );
  XNOR2_X1 U6787 ( .A(n5821), .B(n5820), .ZN(n7412) );
  OR2_X1 U6788 ( .A1(n5763), .A2(n7412), .ZN(n5802) );
  INV_X1 U6789 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7407) );
  OR2_X1 U6790 ( .A1(n7015), .A2(n7407), .ZN(n5801) );
  OAI211_X1 U6791 ( .C1(n5035), .C2(n7406), .A(n5802), .B(n5801), .ZN(n7800)
         );
  NAND2_X1 U6792 ( .A1(n7800), .A2(n6373), .ZN(n5803) );
  NAND2_X1 U6793 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  XNOR2_X1 U6794 ( .A(n5805), .B(n6342), .ZN(n5807) );
  NAND2_X1 U6795 ( .A1(n5806), .A2(n5807), .ZN(n7728) );
  AOI22_X1 U6796 ( .A1(n10173), .A2(n6063), .B1(n6388), .B2(n7800), .ZN(n7730)
         );
  NAND2_X1 U6797 ( .A1(n7728), .A2(n7730), .ZN(n5810) );
  INV_X1 U6798 ( .A(n5807), .ZN(n5808) );
  NAND2_X1 U6799 ( .A1(n5810), .A2(n7729), .ZN(n7925) );
  NAND2_X1 U6800 ( .A1(n7101), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U6801 ( .A1(n5811), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5844) );
  OAI21_X1 U6802 ( .B1(n5811), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5844), .ZN(
        n7810) );
  INV_X1 U6803 ( .A(n7810), .ZN(n7920) );
  NAND2_X1 U6804 ( .A1(n6424), .A2(n7920), .ZN(n5814) );
  NAND2_X1 U6805 ( .A1(n6302), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U6806 ( .A1(n6303), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5812) );
  NAND4_X1 U6807 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n7734)
         );
  NAND2_X1 U6808 ( .A1(n7734), .A2(n6388), .ZN(n5828) );
  INV_X1 U6809 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U6810 ( .A1(n5817), .A2(n5816), .ZN(n5863) );
  NAND2_X1 U6811 ( .A1(n5863), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5818) );
  INV_X1 U6812 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U6813 ( .A1(n5818), .A2(n9772), .ZN(n5839) );
  OR2_X1 U6814 ( .A1(n5818), .A2(n9772), .ZN(n5819) );
  INV_X1 U6815 ( .A(n10595), .ZN(n7419) );
  NAND2_X1 U6816 ( .A1(n5821), .A2(n5820), .ZN(n5824) );
  NAND2_X1 U6817 ( .A1(n5822), .A2(SI_5_), .ZN(n5823) );
  MUX2_X1 U6818 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6995), .Z(n5837) );
  XNOR2_X1 U6819 ( .A(n5837), .B(n9655), .ZN(n5835) );
  XNOR2_X1 U6820 ( .A(n5836), .B(n5835), .ZN(n7432) );
  OR2_X1 U6821 ( .A1(n7432), .A2(n5763), .ZN(n5826) );
  INV_X1 U6822 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7420) );
  OR2_X1 U6823 ( .A1(n7015), .A2(n7420), .ZN(n5825) );
  NAND2_X1 U6824 ( .A1(n7930), .A2(n6373), .ZN(n5827) );
  NAND2_X1 U6825 ( .A1(n5828), .A2(n5827), .ZN(n5829) );
  XNOR2_X1 U6826 ( .A(n5829), .B(n6342), .ZN(n5830) );
  AOI22_X1 U6827 ( .A1(n7734), .A2(n6063), .B1(n6388), .B2(n7930), .ZN(n5831)
         );
  XNOR2_X1 U6828 ( .A(n5830), .B(n5831), .ZN(n7926) );
  NAND2_X1 U6829 ( .A1(n7925), .A2(n7926), .ZN(n5834) );
  INV_X1 U6830 ( .A(n5830), .ZN(n5832) );
  NAND2_X1 U6831 ( .A1(n5832), .A2(n5831), .ZN(n5833) );
  NAND2_X1 U6832 ( .A1(n5834), .A2(n5833), .ZN(n7838) );
  NAND2_X1 U6833 ( .A1(n5837), .A2(SI_6_), .ZN(n5838) );
  MUX2_X1 U6834 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n5768), .Z(n5862) );
  XNOR2_X1 U6835 ( .A(n5862), .B(SI_7_), .ZN(n5859) );
  XNOR2_X1 U6836 ( .A(n5861), .B(n5859), .ZN(n7434) );
  NAND2_X1 U6837 ( .A1(n7434), .A2(n7005), .ZN(n5842) );
  NAND2_X1 U6838 ( .A1(n5839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U6839 ( .A(n5840), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7510) );
  AOI22_X1 U6840 ( .A1(n5037), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6142), .B2(
        n7510), .ZN(n5841) );
  NAND2_X1 U6841 ( .A1(n7910), .A2(n6373), .ZN(n5851) );
  NAND2_X1 U6842 ( .A1(n7101), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5849) );
  AND2_X1 U6843 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  NOR2_X1 U6844 ( .A1(n5870), .A2(n5845), .ZN(n10864) );
  NAND2_X1 U6845 ( .A1(n6424), .A2(n10864), .ZN(n5848) );
  NAND2_X1 U6846 ( .A1(n6302), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U6847 ( .A1(n6303), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5846) );
  NAND4_X1 U6848 ( .A1(n5849), .A2(n5848), .A3(n5847), .A4(n5846), .ZN(n10172)
         );
  NAND2_X1 U6849 ( .A1(n10172), .A2(n6388), .ZN(n5850) );
  NAND2_X1 U6850 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  XNOR2_X1 U6851 ( .A(n5852), .B(n5686), .ZN(n5857) );
  NAND2_X1 U6852 ( .A1(n7910), .A2(n6388), .ZN(n5854) );
  NAND2_X1 U6853 ( .A1(n10172), .A2(n6063), .ZN(n5853) );
  NAND2_X1 U6854 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  XNOR2_X1 U6855 ( .A(n5857), .B(n5855), .ZN(n7840) );
  NAND2_X1 U6856 ( .A1(n7838), .A2(n7840), .ZN(n7839) );
  INV_X1 U6857 ( .A(n5855), .ZN(n5856) );
  NAND2_X1 U6858 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  NAND2_X1 U6859 ( .A1(n7839), .A2(n5858), .ZN(n5879) );
  INV_X1 U6860 ( .A(n5859), .ZN(n5860) );
  MUX2_X1 U6861 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6995), .Z(n5887) );
  XNOR2_X1 U6862 ( .A(n5886), .B(n5884), .ZN(n7444) );
  NAND2_X1 U6863 ( .A1(n7444), .A2(n7005), .ZN(n5869) );
  NAND2_X1 U6864 ( .A1(n5866), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5865) );
  MUX2_X1 U6865 ( .A(n5865), .B(P1_IR_REG_31__SCAN_IN), .S(n5864), .Z(n5867)
         );
  AOI22_X1 U6866 ( .A1(n5037), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6142), .B2(
        n7488), .ZN(n5868) );
  OR2_X1 U6867 ( .A1(n10882), .A2(n6384), .ZN(n5877) );
  NAND2_X1 U6868 ( .A1(n7101), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U6869 ( .A1(n5870), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5896) );
  OR2_X1 U6870 ( .A1(n5870), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5871) );
  AND2_X1 U6871 ( .A1(n5896), .A2(n5871), .ZN(n8121) );
  NAND2_X1 U6872 ( .A1(n6424), .A2(n8121), .ZN(n5874) );
  NAND2_X1 U6873 ( .A1(n6302), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U6874 ( .A1(n6303), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5872) );
  NAND4_X1 U6875 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n10171)
         );
  NAND2_X1 U6876 ( .A1(n10171), .A2(n6063), .ZN(n5876) );
  AND2_X1 U6877 ( .A1(n5877), .A2(n5876), .ZN(n5880) );
  NAND2_X1 U6878 ( .A1(n5879), .A2(n5880), .ZN(n8126) );
  INV_X1 U6879 ( .A(n10171), .ZN(n10852) );
  OAI22_X1 U6880 ( .A1(n10882), .A2(n6341), .B1(n10852), .B2(n6384), .ZN(n5878) );
  XNOR2_X1 U6881 ( .A(n5878), .B(n6342), .ZN(n8129) );
  NAND2_X1 U6882 ( .A1(n8126), .A2(n8129), .ZN(n5883) );
  NAND2_X1 U6883 ( .A1(n5887), .A2(SI_8_), .ZN(n5888) );
  MUX2_X1 U6884 ( .A(n9750), .B(n7451), .S(n6995), .Z(n5889) );
  INV_X1 U6885 ( .A(n5889), .ZN(n5890) );
  NAND2_X1 U6886 ( .A1(n5890), .A2(SI_9_), .ZN(n5891) );
  NAND2_X1 U6887 ( .A1(n5909), .A2(n5891), .ZN(n5910) );
  XNOR2_X1 U6888 ( .A(n5911), .B(n5910), .ZN(n7450) );
  NAND2_X1 U6889 ( .A1(n7450), .A2(n7005), .ZN(n5894) );
  NAND2_X1 U6890 ( .A1(n5917), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5892) );
  XNOR2_X1 U6891 ( .A(n5892), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7500) );
  AOI22_X1 U6892 ( .A1(n5037), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6142), .B2(
        n7500), .ZN(n5893) );
  NAND2_X1 U6893 ( .A1(n8076), .A2(n6373), .ZN(n5903) );
  NAND2_X1 U6894 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  AND2_X1 U6895 ( .A1(n5922), .A2(n5897), .ZN(n8022) );
  NAND2_X1 U6896 ( .A1(n6424), .A2(n8022), .ZN(n5901) );
  NAND2_X1 U6897 ( .A1(n7101), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U6898 ( .A1(n6302), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U6899 ( .A1(n6303), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5898) );
  NAND4_X1 U6900 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n10170)
         );
  NAND2_X1 U6901 ( .A1(n10170), .A2(n6388), .ZN(n5902) );
  NAND2_X1 U6902 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  XNOR2_X1 U6903 ( .A(n5904), .B(n5686), .ZN(n5907) );
  AND2_X1 U6904 ( .A1(n10170), .A2(n6063), .ZN(n5905) );
  AOI21_X1 U6905 ( .B1(n8076), .B2(n6388), .A(n5905), .ZN(n5906) );
  XNOR2_X1 U6906 ( .A(n5907), .B(n5906), .ZN(n8018) );
  NAND2_X1 U6907 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  MUX2_X1 U6908 ( .A(n7540), .B(n7538), .S(n6995), .Z(n5912) );
  INV_X1 U6909 ( .A(n5912), .ZN(n5913) );
  NAND2_X1 U6910 ( .A1(n5913), .A2(SI_10_), .ZN(n5914) );
  NAND2_X1 U6911 ( .A1(n5937), .A2(n5916), .ZN(n7536) );
  NAND2_X1 U6912 ( .A1(n7536), .A2(n7005), .ZN(n5921) );
  OAI21_X1 U6913 ( .B1(n5917), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5918) );
  OR2_X1 U6914 ( .A1(n5918), .A2(n9570), .ZN(n5919) );
  NAND2_X1 U6915 ( .A1(n5918), .A2(n9570), .ZN(n5939) );
  AOI22_X1 U6916 ( .A1(n5037), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6142), .B2(
        n7606), .ZN(n5920) );
  NAND2_X2 U6917 ( .A1(n5921), .A2(n5920), .ZN(n8475) );
  NAND2_X1 U6918 ( .A1(n8475), .A2(n6373), .ZN(n5929) );
  NAND2_X1 U6919 ( .A1(n7101), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U6920 ( .A1(n5922), .A2(n7568), .ZN(n5923) );
  AND2_X1 U6921 ( .A1(n5944), .A2(n5923), .ZN(n8463) );
  NAND2_X1 U6922 ( .A1(n6424), .A2(n8463), .ZN(n5926) );
  NAND2_X1 U6923 ( .A1(n6302), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U6924 ( .A1(n6303), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5924) );
  NAND4_X1 U6925 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .ZN(n10169)
         );
  NAND2_X1 U6926 ( .A1(n10169), .A2(n6388), .ZN(n5928) );
  NAND2_X1 U6927 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  NAND2_X1 U6928 ( .A1(n8475), .A2(n6388), .ZN(n5932) );
  NAND2_X1 U6929 ( .A1(n10169), .A2(n6063), .ZN(n5931) );
  NAND2_X1 U6930 ( .A1(n5932), .A2(n5931), .ZN(n8471) );
  NAND2_X1 U6931 ( .A1(n8468), .A2(n8471), .ZN(n5935) );
  INV_X1 U6932 ( .A(n5933), .ZN(n5934) );
  NAND2_X1 U6933 ( .A1(n5934), .A2(n5105), .ZN(n8469) );
  NAND2_X1 U6934 ( .A1(n5935), .A2(n8469), .ZN(n8220) );
  MUX2_X1 U6935 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n6995), .Z(n5960) );
  NAND2_X1 U6936 ( .A1(n5939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5940) );
  XNOR2_X1 U6937 ( .A(n5940), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7881) );
  AOI22_X1 U6938 ( .A1(n5037), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6142), .B2(
        n7881), .ZN(n5941) );
  NAND2_X1 U6939 ( .A1(n8094), .A2(n6373), .ZN(n5951) );
  NAND2_X1 U6940 ( .A1(n7101), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5949) );
  INV_X1 U6941 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5943) );
  AND2_X1 U6942 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  NOR2_X1 U6943 ( .A1(n5972), .A2(n5945), .ZN(n8228) );
  NAND2_X1 U6944 ( .A1(n6424), .A2(n8228), .ZN(n5948) );
  NAND2_X1 U6945 ( .A1(n6302), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U6946 ( .A1(n6303), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5946) );
  NAND4_X1 U6947 ( .A1(n5949), .A2(n5948), .A3(n5947), .A4(n5946), .ZN(n10168)
         );
  NAND2_X1 U6948 ( .A1(n10168), .A2(n6388), .ZN(n5950) );
  NAND2_X1 U6949 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  XNOR2_X1 U6950 ( .A(n5952), .B(n6342), .ZN(n5956) );
  AND2_X1 U6951 ( .A1(n10168), .A2(n6063), .ZN(n5953) );
  AOI21_X1 U6952 ( .B1(n8094), .B2(n6388), .A(n5953), .ZN(n5954) );
  XNOR2_X1 U6953 ( .A(n5956), .B(n5954), .ZN(n8223) );
  INV_X1 U6954 ( .A(n5954), .ZN(n5955) );
  NAND2_X1 U6955 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  NAND2_X1 U6956 ( .A1(n5960), .A2(SI_11_), .ZN(n5961) );
  INV_X1 U6957 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5962) );
  MUX2_X1 U6958 ( .A(n7627), .B(n5962), .S(n6995), .Z(n5964) );
  INV_X1 U6959 ( .A(SI_12_), .ZN(n5963) );
  INV_X1 U6960 ( .A(n5964), .ZN(n5965) );
  NAND2_X1 U6961 ( .A1(n5965), .A2(SI_12_), .ZN(n5966) );
  NAND2_X1 U6962 ( .A1(n5985), .A2(n5966), .ZN(n5986) );
  XNOR2_X1 U6963 ( .A(n5987), .B(n5986), .ZN(n7624) );
  NAND2_X1 U6964 ( .A1(n7624), .A2(n7005), .ZN(n5971) );
  NAND2_X1 U6965 ( .A1(n5967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  MUX2_X1 U6966 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5968), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5969) );
  OR2_X1 U6967 ( .A1(n5967), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5995) );
  AND2_X1 U6968 ( .A1(n5969), .A2(n5995), .ZN(n10185) );
  AOI22_X1 U6969 ( .A1(n5037), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6142), .B2(
        n10185), .ZN(n5970) );
  NAND2_X1 U6970 ( .A1(n8385), .A2(n6373), .ZN(n5979) );
  OR2_X1 U6971 ( .A1(n5972), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U6972 ( .A1(n5972), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6000) );
  AND2_X1 U6973 ( .A1(n5973), .A2(n6000), .ZN(n8305) );
  NAND2_X1 U6974 ( .A1(n6424), .A2(n8305), .ZN(n5977) );
  NAND2_X1 U6975 ( .A1(n7101), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U6976 ( .A1(n6302), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U6977 ( .A1(n6303), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5974) );
  NAND4_X1 U6978 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n11005)
         );
  NAND2_X1 U6979 ( .A1(n11005), .A2(n6388), .ZN(n5978) );
  NAND2_X1 U6980 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  XNOR2_X1 U6981 ( .A(n5980), .B(n5686), .ZN(n8303) );
  AND2_X1 U6982 ( .A1(n11005), .A2(n6063), .ZN(n5981) );
  AOI21_X1 U6983 ( .B1(n8385), .B2(n6388), .A(n5981), .ZN(n5983) );
  NAND2_X1 U6984 ( .A1(n8303), .A2(n5983), .ZN(n5982) );
  INV_X1 U6985 ( .A(n8303), .ZN(n5984) );
  INV_X1 U6986 ( .A(n5983), .ZN(n8302) );
  INV_X1 U6987 ( .A(n8555), .ZN(n6012) );
  INV_X1 U6988 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5988) );
  MUX2_X1 U6989 ( .A(n5988), .B(n7661), .S(n6995), .Z(n5990) );
  INV_X1 U6990 ( .A(SI_13_), .ZN(n5989) );
  INV_X1 U6991 ( .A(n5990), .ZN(n5991) );
  NAND2_X1 U6992 ( .A1(n5991), .A2(SI_13_), .ZN(n5992) );
  XNOR2_X1 U6993 ( .A(n6017), .B(n5633), .ZN(n7657) );
  NAND2_X1 U6994 ( .A1(n7657), .A2(n7005), .ZN(n5998) );
  NAND2_X1 U6995 ( .A1(n5995), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5993) );
  MUX2_X1 U6996 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5993), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n5994) );
  INV_X1 U6997 ( .A(n5994), .ZN(n5996) );
  NOR2_X1 U6998 ( .A1(n5995), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6023) );
  NOR2_X1 U6999 ( .A1(n5996), .A2(n6023), .ZN(n10201) );
  AOI22_X1 U7000 ( .A1(n5037), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6142), .B2(
        n10201), .ZN(n5997) );
  NAND2_X1 U7001 ( .A1(n8552), .A2(n6373), .ZN(n6007) );
  NAND2_X1 U7002 ( .A1(n7101), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6005) );
  INV_X1 U7003 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7004 ( .A1(n6000), .A2(n5999), .ZN(n6001) );
  AND2_X1 U7005 ( .A1(n6027), .A2(n6001), .ZN(n11026) );
  NAND2_X1 U7006 ( .A1(n6424), .A2(n11026), .ZN(n6004) );
  NAND2_X1 U7007 ( .A1(n6302), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7008 ( .A1(n6303), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6002) );
  NAND4_X1 U7009 ( .A1(n6005), .A2(n6004), .A3(n6003), .A4(n6002), .ZN(n10167)
         );
  NAND2_X1 U7010 ( .A1(n10167), .A2(n6388), .ZN(n6006) );
  NAND2_X1 U7011 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  XNOR2_X1 U7012 ( .A(n6008), .B(n6342), .ZN(n6013) );
  NAND2_X1 U7013 ( .A1(n8552), .A2(n6388), .ZN(n6010) );
  NAND2_X1 U7014 ( .A1(n10167), .A2(n6063), .ZN(n6009) );
  NAND2_X1 U7015 ( .A1(n6010), .A2(n6009), .ZN(n6014) );
  AND2_X1 U7016 ( .A1(n6013), .A2(n6014), .ZN(n8556) );
  INV_X1 U7017 ( .A(n8556), .ZN(n6011) );
  NAND2_X1 U7018 ( .A1(n6012), .A2(n6011), .ZN(n8553) );
  INV_X1 U7019 ( .A(n6013), .ZN(n6016) );
  INV_X1 U7020 ( .A(n6014), .ZN(n6015) );
  NAND2_X1 U7021 ( .A1(n6016), .A2(n6015), .ZN(n8554) );
  MUX2_X1 U7022 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n6995), .Z(n6041) );
  INV_X1 U7023 ( .A(SI_14_), .ZN(n6020) );
  NAND2_X1 U7024 ( .A1(n7659), .A2(n7005), .ZN(n6026) );
  NOR2_X1 U7025 ( .A1(n6023), .A2(n10534), .ZN(n6021) );
  MUX2_X1 U7026 ( .A(n10534), .B(n6021), .S(P1_IR_REG_14__SCAN_IN), .Z(n6022)
         );
  INV_X1 U7027 ( .A(n6022), .ZN(n6024) );
  INV_X1 U7028 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U7029 ( .A1(n6023), .A2(n9578), .ZN(n6066) );
  AOI22_X1 U7030 ( .A1(n5037), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6142), .B2(
        n10217), .ZN(n6025) );
  NAND2_X1 U7031 ( .A1(n8664), .A2(n6373), .ZN(n6034) );
  NAND2_X1 U7032 ( .A1(n7101), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6032) );
  INV_X1 U7033 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8658) );
  AND2_X1 U7034 ( .A1(n6027), .A2(n8658), .ZN(n6028) );
  NOR2_X1 U7035 ( .A1(n6070), .A2(n6028), .ZN(n8657) );
  NAND2_X1 U7036 ( .A1(n6424), .A2(n8657), .ZN(n6031) );
  NAND2_X1 U7037 ( .A1(n6302), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7038 ( .A1(n6303), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6029) );
  NAND4_X1 U7039 ( .A1(n6032), .A2(n6031), .A3(n6030), .A4(n6029), .ZN(n11004)
         );
  NAND2_X1 U7040 ( .A1(n11004), .A2(n6388), .ZN(n6033) );
  NAND2_X1 U7041 ( .A1(n6034), .A2(n6033), .ZN(n6035) );
  XNOR2_X1 U7042 ( .A(n6035), .B(n5686), .ZN(n6038) );
  NAND2_X1 U7043 ( .A1(n8664), .A2(n6388), .ZN(n6037) );
  NAND2_X1 U7044 ( .A1(n11004), .A2(n6063), .ZN(n6036) );
  NAND2_X1 U7045 ( .A1(n6037), .A2(n6036), .ZN(n8656) );
  INV_X1 U7046 ( .A(n6038), .ZN(n6039) );
  INV_X1 U7047 ( .A(n6040), .ZN(n6043) );
  NAND2_X1 U7048 ( .A1(n6041), .A2(SI_14_), .ZN(n6042) );
  MUX2_X1 U7049 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6995), .Z(n6046) );
  XNOR2_X1 U7050 ( .A(n6046), .B(SI_15_), .ZN(n6064) );
  INV_X1 U7051 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6047) );
  MUX2_X1 U7052 ( .A(n9742), .B(n6047), .S(n6995), .Z(n6048) );
  INV_X1 U7053 ( .A(SI_16_), .ZN(n9439) );
  INV_X1 U7054 ( .A(n6048), .ZN(n6049) );
  NAND2_X1 U7055 ( .A1(n6049), .A2(SI_16_), .ZN(n6050) );
  NAND2_X1 U7056 ( .A1(n6089), .A2(n6050), .ZN(n6052) );
  NAND2_X1 U7057 ( .A1(n6053), .A2(n6052), .ZN(n6054) );
  NAND2_X1 U7058 ( .A1(n6090), .A2(n6054), .ZN(n7690) );
  NAND2_X1 U7059 ( .A1(n7690), .A2(n7005), .ZN(n6057) );
  OR2_X1 U7060 ( .A1(n6066), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7061 ( .A1(n6055), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6092) );
  XNOR2_X1 U7062 ( .A(n6092), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8499) );
  AOI22_X1 U7063 ( .A1(n5037), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6142), .B2(
        n8499), .ZN(n6056) );
  NAND2_X1 U7064 ( .A1(n7101), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7065 ( .A1(n6070), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6071) );
  INV_X1 U7066 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8065) );
  AOI21_X1 U7067 ( .B1(n6071), .B2(n8065), .A(n6100), .ZN(n10064) );
  NAND2_X1 U7068 ( .A1(n6424), .A2(n10064), .ZN(n6060) );
  NAND2_X1 U7069 ( .A1(n6302), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7070 ( .A1(n6303), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6058) );
  NAND4_X1 U7071 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6058), .ZN(n10146)
         );
  INV_X1 U7072 ( .A(n10146), .ZN(n10076) );
  OAI22_X1 U7073 ( .A1(n11084), .A2(n6341), .B1(n10076), .B2(n6384), .ZN(n6062) );
  XNOR2_X1 U7074 ( .A(n6062), .B(n6342), .ZN(n6083) );
  OAI22_X1 U7075 ( .A1(n11084), .A2(n6384), .B1(n10076), .B2(n6390), .ZN(
        n10061) );
  XNOR2_X1 U7076 ( .A(n6065), .B(n6064), .ZN(n7686) );
  NAND2_X1 U7077 ( .A1(n7686), .A2(n7005), .ZN(n6069) );
  NAND2_X1 U7078 ( .A1(n6066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U7079 ( .A(n6067), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8061) );
  AOI22_X1 U7080 ( .A1(n5037), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6142), .B2(
        n8061), .ZN(n6068) );
  NAND2_X1 U7081 ( .A1(n10135), .A2(n6388), .ZN(n6078) );
  NAND2_X1 U7082 ( .A1(n7101), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6076) );
  OR2_X1 U7083 ( .A1(n6070), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6072) );
  AND2_X1 U7084 ( .A1(n6072), .A2(n6071), .ZN(n10153) );
  NAND2_X1 U7085 ( .A1(n6424), .A2(n10153), .ZN(n6075) );
  NAND2_X1 U7086 ( .A1(n6302), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7087 ( .A1(n6303), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6073) );
  NAND4_X1 U7088 ( .A1(n6076), .A2(n6075), .A3(n6074), .A4(n6073), .ZN(n8659)
         );
  NAND2_X1 U7089 ( .A1(n8659), .A2(n6063), .ZN(n6077) );
  NAND2_X1 U7090 ( .A1(n6078), .A2(n6077), .ZN(n10137) );
  NAND2_X1 U7091 ( .A1(n10135), .A2(n6373), .ZN(n6080) );
  NAND2_X1 U7092 ( .A1(n8659), .A2(n6388), .ZN(n6079) );
  NAND2_X1 U7093 ( .A1(n6080), .A2(n6079), .ZN(n6081) );
  XNOR2_X1 U7094 ( .A(n6081), .B(n6342), .ZN(n6084) );
  AOI22_X1 U7095 ( .A1(n6083), .A2(n10061), .B1(n10137), .B2(n6084), .ZN(n6082) );
  NAND2_X1 U7096 ( .A1(n10058), .A2(n6082), .ZN(n6088) );
  INV_X1 U7097 ( .A(n6083), .ZN(n10062) );
  OAI21_X1 U7098 ( .B1(n6084), .B2(n10137), .A(n10061), .ZN(n6086) );
  NOR2_X1 U7099 ( .A1(n10061), .A2(n10137), .ZN(n6085) );
  INV_X1 U7100 ( .A(n6084), .ZN(n10059) );
  AOI22_X1 U7101 ( .A1(n10062), .A2(n6086), .B1(n6085), .B2(n10059), .ZN(n6087) );
  MUX2_X1 U7102 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n6995), .Z(n6112) );
  XNOR2_X1 U7103 ( .A(n6110), .B(n6111), .ZN(n7796) );
  NAND2_X1 U7104 ( .A1(n7796), .A2(n7005), .ZN(n6097) );
  INV_X1 U7105 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6091) );
  AOI21_X1 U7106 ( .B1(n6092), .B2(n6091), .A(n10534), .ZN(n6093) );
  NAND2_X1 U7107 ( .A1(n6093), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6095) );
  INV_X1 U7108 ( .A(n6093), .ZN(n6094) );
  INV_X1 U7109 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U7110 ( .A1(n6094), .A2(n9583), .ZN(n6115) );
  AOI22_X1 U7111 ( .A1(n5037), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6142), .B2(
        n10227), .ZN(n6096) );
  NAND2_X1 U7112 ( .A1(n10514), .A2(n6373), .ZN(n6105) );
  INV_X1 U7113 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8502) );
  NAND2_X1 U7114 ( .A1(n6302), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7115 ( .A1(n6303), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6098) );
  OAI211_X1 U7116 ( .C1(n6422), .C2(n8502), .A(n6099), .B(n6098), .ZN(n6103)
         );
  NAND2_X1 U7117 ( .A1(n6100), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6124) );
  OR2_X1 U7118 ( .A1(n6100), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7119 ( .A1(n6124), .A2(n6101), .ZN(n10079) );
  NOR2_X1 U7120 ( .A1(n10079), .A2(n6334), .ZN(n6102) );
  NOR2_X1 U7121 ( .A1(n6103), .A2(n6102), .ZN(n8626) );
  OR2_X1 U7122 ( .A1(n8626), .A2(n6384), .ZN(n6104) );
  NAND2_X1 U7123 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  XNOR2_X1 U7124 ( .A(n6106), .B(n5686), .ZN(n10073) );
  NOR2_X1 U7125 ( .A1(n8626), .A2(n6390), .ZN(n6107) );
  AOI21_X1 U7126 ( .B1(n10514), .B2(n6388), .A(n6107), .ZN(n10072) );
  AND2_X1 U7127 ( .A1(n10073), .A2(n10072), .ZN(n6109) );
  OR2_X1 U7128 ( .A1(n10073), .A2(n10072), .ZN(n6108) );
  NAND2_X1 U7129 ( .A1(n6112), .A2(SI_17_), .ZN(n6113) );
  NAND2_X1 U7130 ( .A1(n6114), .A2(n6113), .ZN(n6135) );
  MUX2_X1 U7131 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n6995), .Z(n6136) );
  XNOR2_X1 U7132 ( .A(n6136), .B(SI_18_), .ZN(n6133) );
  XNOR2_X1 U7133 ( .A(n6135), .B(n6133), .ZN(n7864) );
  NAND2_X1 U7134 ( .A1(n7864), .A2(n7005), .ZN(n6118) );
  NAND2_X1 U7135 ( .A1(n6115), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6116) );
  XNOR2_X1 U7136 ( .A(n6116), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U7137 ( .A1(n5037), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6142), .B2(
        n10244), .ZN(n6117) );
  NAND2_X1 U7138 ( .A1(n10507), .A2(n6388), .ZN(n6129) );
  INV_X1 U7139 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8497) );
  NAND2_X1 U7140 ( .A1(n6303), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7141 ( .A1(n6302), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6119) );
  OAI211_X1 U7142 ( .C1(n6422), .C2(n8497), .A(n6120), .B(n6119), .ZN(n6121)
         );
  INV_X1 U7143 ( .A(n6121), .ZN(n6127) );
  INV_X1 U7144 ( .A(n6124), .ZN(n6122) );
  NAND2_X1 U7145 ( .A1(n6122), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6147) );
  INV_X1 U7146 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7147 ( .A1(n6124), .A2(n6123), .ZN(n6125) );
  AND2_X1 U7148 ( .A1(n6147), .A2(n6125), .ZN(n10120) );
  NAND2_X1 U7149 ( .A1(n10120), .A2(n6424), .ZN(n6126) );
  INV_X1 U7150 ( .A(n10430), .ZN(n10165) );
  NAND2_X1 U7151 ( .A1(n10165), .A2(n6063), .ZN(n6128) );
  NAND2_X1 U7152 ( .A1(n6129), .A2(n6128), .ZN(n10113) );
  NAND2_X1 U7153 ( .A1(n10507), .A2(n6373), .ZN(n6131) );
  NAND2_X1 U7154 ( .A1(n10165), .A2(n6388), .ZN(n6130) );
  NAND2_X1 U7155 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  XNOR2_X1 U7156 ( .A(n6132), .B(n6342), .ZN(n10112) );
  INV_X1 U7157 ( .A(n10027), .ZN(n6161) );
  NAND2_X1 U7158 ( .A1(n6135), .A2(n6134), .ZN(n6138) );
  NAND2_X1 U7159 ( .A1(n6136), .A2(SI_18_), .ZN(n6137) );
  INV_X1 U7160 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7957) );
  MUX2_X1 U7161 ( .A(n9736), .B(n7957), .S(n6995), .Z(n6139) );
  INV_X1 U7162 ( .A(SI_19_), .ZN(n9631) );
  INV_X1 U7163 ( .A(n6139), .ZN(n6140) );
  NAND2_X1 U7164 ( .A1(n6140), .A2(SI_19_), .ZN(n6141) );
  NAND2_X1 U7165 ( .A1(n6166), .A2(n6141), .ZN(n6167) );
  XNOR2_X1 U7166 ( .A(n6168), .B(n6167), .ZN(n7956) );
  NAND2_X1 U7167 ( .A1(n7956), .A2(n7005), .ZN(n6144) );
  AOI22_X1 U7168 ( .A1(n5037), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10344), 
        .B2(n6142), .ZN(n6143) );
  NAND2_X1 U7169 ( .A1(n10503), .A2(n6373), .ZN(n6156) );
  INV_X1 U7170 ( .A(n6147), .ZN(n6145) );
  INV_X1 U7171 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7172 ( .A1(n6147), .A2(n6146), .ZN(n6148) );
  NAND2_X1 U7173 ( .A1(n6176), .A2(n6148), .ZN(n10436) );
  OR2_X1 U7174 ( .A1(n10436), .A2(n6334), .ZN(n6154) );
  INV_X1 U7175 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7176 ( .A1(n6303), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7177 ( .A1(n6302), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6149) );
  OAI211_X1 U7178 ( .C1(n6422), .C2(n6151), .A(n6150), .B(n6149), .ZN(n6152)
         );
  INV_X1 U7179 ( .A(n6152), .ZN(n6153) );
  NAND2_X1 U7180 ( .A1(n10164), .A2(n6388), .ZN(n6155) );
  NAND2_X1 U7181 ( .A1(n6156), .A2(n6155), .ZN(n6157) );
  XNOR2_X1 U7182 ( .A(n6157), .B(n6342), .ZN(n6162) );
  NAND2_X1 U7183 ( .A1(n10503), .A2(n6388), .ZN(n6159) );
  NAND2_X1 U7184 ( .A1(n10164), .A2(n6063), .ZN(n6158) );
  NAND2_X1 U7185 ( .A1(n6159), .A2(n6158), .ZN(n6163) );
  AND2_X1 U7186 ( .A1(n6162), .A2(n6163), .ZN(n10029) );
  INV_X1 U7187 ( .A(n10029), .ZN(n6160) );
  INV_X1 U7188 ( .A(n6162), .ZN(n6165) );
  INV_X1 U7189 ( .A(n6163), .ZN(n6164) );
  NAND2_X1 U7190 ( .A1(n6165), .A2(n6164), .ZN(n10028) );
  INV_X1 U7191 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8149) );
  MUX2_X1 U7192 ( .A(n9737), .B(n8149), .S(n6995), .Z(n6169) );
  INV_X1 U7193 ( .A(SI_20_), .ZN(n9431) );
  NAND2_X1 U7194 ( .A1(n6169), .A2(n9431), .ZN(n6194) );
  INV_X1 U7195 ( .A(n6169), .ZN(n6170) );
  NAND2_X1 U7196 ( .A1(n6170), .A2(SI_20_), .ZN(n6171) );
  XNOR2_X1 U7197 ( .A(n6193), .B(n6192), .ZN(n8039) );
  NAND2_X1 U7198 ( .A1(n8039), .A2(n7005), .ZN(n6173) );
  OR2_X1 U7199 ( .A1(n7015), .A2(n9737), .ZN(n6172) );
  NAND2_X1 U7200 ( .A1(n10496), .A2(n6373), .ZN(n6185) );
  INV_X1 U7201 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7202 ( .A1(n6176), .A2(n6175), .ZN(n6177) );
  NAND2_X1 U7203 ( .A1(n6198), .A2(n6177), .ZN(n10410) );
  OR2_X1 U7204 ( .A1(n10410), .A2(n6334), .ZN(n6183) );
  INV_X1 U7205 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7206 ( .A1(n6303), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7207 ( .A1(n6302), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6178) );
  OAI211_X1 U7208 ( .C1(n6422), .C2(n6180), .A(n6179), .B(n6178), .ZN(n6181)
         );
  INV_X1 U7209 ( .A(n6181), .ZN(n6182) );
  INV_X1 U7210 ( .A(n10431), .ZN(n10163) );
  NAND2_X1 U7211 ( .A1(n10163), .A2(n6388), .ZN(n6184) );
  NAND2_X1 U7212 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  XNOR2_X1 U7213 ( .A(n6186), .B(n5686), .ZN(n10094) );
  NOR2_X1 U7214 ( .A1(n10431), .A2(n6390), .ZN(n6187) );
  AOI21_X1 U7215 ( .B1(n10496), .B2(n6388), .A(n6187), .ZN(n10093) );
  INV_X1 U7216 ( .A(n10094), .ZN(n6189) );
  INV_X1 U7217 ( .A(n10093), .ZN(n6188) );
  NAND2_X1 U7218 ( .A1(n6189), .A2(n6188), .ZN(n6190) );
  MUX2_X1 U7219 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6995), .Z(n6217) );
  INV_X1 U7220 ( .A(SI_21_), .ZN(n9630) );
  XNOR2_X1 U7221 ( .A(n6217), .B(n9630), .ZN(n6216) );
  XNOR2_X1 U7222 ( .A(n6220), .B(n6216), .ZN(n8100) );
  NAND2_X1 U7223 ( .A1(n8100), .A2(n7005), .ZN(n6197) );
  INV_X1 U7224 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8101) );
  OR2_X1 U7225 ( .A1(n7015), .A2(n8101), .ZN(n6196) );
  NAND2_X2 U7226 ( .A1(n6197), .A2(n6196), .ZN(n10493) );
  NAND2_X1 U7227 ( .A1(n10493), .A2(n6373), .ZN(n6207) );
  INV_X1 U7228 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U7229 ( .A1(n6198), .A2(n10042), .ZN(n6199) );
  NAND2_X1 U7230 ( .A1(n6226), .A2(n6199), .ZN(n10394) );
  OR2_X1 U7231 ( .A1(n10394), .A2(n6334), .ZN(n6205) );
  INV_X1 U7232 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7233 ( .A1(n6302), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7234 ( .A1(n6303), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6200) );
  OAI211_X1 U7235 ( .C1(n6422), .C2(n6202), .A(n6201), .B(n6200), .ZN(n6203)
         );
  INV_X1 U7236 ( .A(n6203), .ZN(n6204) );
  NAND2_X1 U7237 ( .A1(n10162), .A2(n6388), .ZN(n6206) );
  NAND2_X1 U7238 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  XNOR2_X1 U7239 ( .A(n6208), .B(n6342), .ZN(n6212) );
  NAND2_X1 U7240 ( .A1(n10493), .A2(n6388), .ZN(n6210) );
  NAND2_X1 U7241 ( .A1(n10162), .A2(n6063), .ZN(n6209) );
  NAND2_X1 U7242 ( .A1(n6210), .A2(n6209), .ZN(n6213) );
  AND2_X1 U7243 ( .A1(n6212), .A2(n6213), .ZN(n10038) );
  INV_X1 U7244 ( .A(n6212), .ZN(n6215) );
  INV_X1 U7245 ( .A(n6213), .ZN(n6214) );
  NAND2_X1 U7246 ( .A1(n6215), .A2(n6214), .ZN(n10036) );
  INV_X1 U7247 ( .A(n6216), .ZN(n6219) );
  NAND2_X1 U7248 ( .A1(n6217), .A2(SI_21_), .ZN(n6218) );
  INV_X1 U7249 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9530) );
  INV_X1 U7250 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8292) );
  MUX2_X1 U7251 ( .A(n9530), .B(n8292), .S(n6995), .Z(n6221) );
  INV_X1 U7252 ( .A(SI_22_), .ZN(n9623) );
  NAND2_X1 U7253 ( .A1(n6221), .A2(n9623), .ZN(n6241) );
  INV_X1 U7254 ( .A(n6221), .ZN(n6222) );
  NAND2_X1 U7255 ( .A1(n6222), .A2(SI_22_), .ZN(n6223) );
  NAND2_X1 U7256 ( .A1(n6241), .A2(n6223), .ZN(n6242) );
  XNOR2_X1 U7257 ( .A(n6243), .B(n6242), .ZN(n8290) );
  NAND2_X1 U7258 ( .A1(n8290), .A2(n7005), .ZN(n6225) );
  OR2_X1 U7259 ( .A1(n7015), .A2(n9530), .ZN(n6224) );
  INV_X1 U7260 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n10106) );
  NAND2_X1 U7261 ( .A1(n6226), .A2(n10106), .ZN(n6227) );
  AND2_X1 U7262 ( .A1(n6251), .A2(n6227), .ZN(n10379) );
  NAND2_X1 U7263 ( .A1(n10379), .A2(n6424), .ZN(n6233) );
  INV_X1 U7264 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7265 ( .A1(n6302), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7266 ( .A1(n6303), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6228) );
  OAI211_X1 U7267 ( .C1(n6422), .C2(n6230), .A(n6229), .B(n6228), .ZN(n6231)
         );
  INV_X1 U7268 ( .A(n6231), .ZN(n6232) );
  NAND2_X1 U7269 ( .A1(n6233), .A2(n6232), .ZN(n10161) );
  INV_X1 U7270 ( .A(n10161), .ZN(n10390) );
  OAI22_X1 U7271 ( .A1(n10485), .A2(n6341), .B1(n10390), .B2(n6384), .ZN(n6234) );
  XNOR2_X1 U7272 ( .A(n6234), .B(n5686), .ZN(n6239) );
  OR2_X1 U7273 ( .A1(n10485), .A2(n6384), .ZN(n6236) );
  NAND2_X1 U7274 ( .A1(n10161), .A2(n6063), .ZN(n6235) );
  NAND2_X1 U7275 ( .A1(n6236), .A2(n6235), .ZN(n6237) );
  XNOR2_X1 U7276 ( .A(n6239), .B(n6237), .ZN(n10104) );
  INV_X1 U7277 ( .A(n6237), .ZN(n6238) );
  NAND2_X1 U7278 ( .A1(n6239), .A2(n6238), .ZN(n6240) );
  INV_X1 U7279 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9731) );
  INV_X1 U7280 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8300) );
  MUX2_X1 U7281 ( .A(n9731), .B(n8300), .S(n6995), .Z(n6244) );
  INV_X1 U7282 ( .A(SI_23_), .ZN(n9424) );
  NAND2_X1 U7283 ( .A1(n6244), .A2(n9424), .ZN(n6269) );
  INV_X1 U7284 ( .A(n6244), .ZN(n6245) );
  NAND2_X1 U7285 ( .A1(n6245), .A2(SI_23_), .ZN(n6246) );
  XNOR2_X1 U7286 ( .A(n6268), .B(n6267), .ZN(n8298) );
  NAND2_X1 U7287 ( .A1(n8298), .A2(n7005), .ZN(n6248) );
  OR2_X1 U7288 ( .A1(n7015), .A2(n9731), .ZN(n6247) );
  NAND2_X2 U7289 ( .A1(n6248), .A2(n6247), .ZN(n10481) );
  NAND2_X1 U7290 ( .A1(n10481), .A2(n6373), .ZN(n6260) );
  INV_X1 U7291 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7292 ( .A1(n6251), .A2(n6250), .ZN(n6252) );
  NAND2_X1 U7293 ( .A1(n6275), .A2(n6252), .ZN(n10022) );
  OR2_X1 U7294 ( .A1(n10022), .A2(n6334), .ZN(n6258) );
  INV_X1 U7295 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7296 ( .A1(n6303), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7297 ( .A1(n6302), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6253) );
  OAI211_X1 U7298 ( .C1(n6422), .C2(n6255), .A(n6254), .B(n6253), .ZN(n6256)
         );
  INV_X1 U7299 ( .A(n6256), .ZN(n6257) );
  INV_X1 U7300 ( .A(n10371), .ZN(n10160) );
  NAND2_X1 U7301 ( .A1(n10160), .A2(n6388), .ZN(n6259) );
  NAND2_X1 U7302 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  XNOR2_X1 U7303 ( .A(n6261), .B(n6342), .ZN(n6264) );
  NAND2_X1 U7304 ( .A1(n6263), .A2(n6264), .ZN(n10019) );
  NOR2_X1 U7305 ( .A1(n10371), .A2(n6390), .ZN(n6262) );
  AOI21_X1 U7306 ( .B1(n10481), .B2(n6388), .A(n6262), .ZN(n10017) );
  NAND2_X1 U7307 ( .A1(n10019), .A2(n10017), .ZN(n10016) );
  INV_X1 U7308 ( .A(n6263), .ZN(n6266) );
  INV_X1 U7309 ( .A(n6264), .ZN(n6265) );
  NAND2_X1 U7310 ( .A1(n6266), .A2(n6265), .ZN(n10018) );
  NAND2_X1 U7311 ( .A1(n10016), .A2(n10018), .ZN(n10084) );
  NAND2_X1 U7312 ( .A1(n6270), .A2(n6269), .ZN(n6293) );
  MUX2_X1 U7313 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6995), .Z(n6290) );
  INV_X1 U7314 ( .A(SI_24_), .ZN(n9622) );
  XNOR2_X1 U7315 ( .A(n6290), .B(n9622), .ZN(n6289) );
  XNOR2_X1 U7316 ( .A(n6293), .B(n6289), .ZN(n8414) );
  NAND2_X1 U7317 ( .A1(n8414), .A2(n7005), .ZN(n6272) );
  INV_X1 U7318 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8415) );
  OR2_X1 U7319 ( .A1(n7015), .A2(n8415), .ZN(n6271) );
  INV_X1 U7320 ( .A(n6275), .ZN(n6273) );
  NAND2_X1 U7321 ( .A1(n6273), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6300) );
  INV_X1 U7322 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7323 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  NAND2_X1 U7324 ( .A1(n6300), .A2(n6276), .ZN(n10087) );
  OR2_X1 U7325 ( .A1(n10087), .A2(n6334), .ZN(n6282) );
  INV_X1 U7326 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7327 ( .A1(n6303), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7328 ( .A1(n6302), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6277) );
  OAI211_X1 U7329 ( .C1(n6422), .C2(n6279), .A(n6278), .B(n6277), .ZN(n6280)
         );
  INV_X1 U7330 ( .A(n6280), .ZN(n6281) );
  OAI22_X1 U7331 ( .A1(n10347), .A2(n6384), .B1(n10359), .B2(n6390), .ZN(n6286) );
  NAND2_X1 U7332 ( .A1(n10476), .A2(n6373), .ZN(n6284) );
  NAND2_X1 U7333 ( .A1(n10159), .A2(n6388), .ZN(n6283) );
  NAND2_X1 U7334 ( .A1(n6284), .A2(n6283), .ZN(n6285) );
  XNOR2_X1 U7335 ( .A(n6285), .B(n6342), .ZN(n6287) );
  XOR2_X1 U7336 ( .A(n6286), .B(n6287), .Z(n10085) );
  OR2_X1 U7337 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  INV_X1 U7338 ( .A(n6289), .ZN(n6292) );
  NAND2_X1 U7339 ( .A1(n6290), .A2(SI_24_), .ZN(n6291) );
  INV_X1 U7340 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9526) );
  INV_X1 U7341 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8595) );
  MUX2_X1 U7342 ( .A(n9526), .B(n8595), .S(n6995), .Z(n6294) );
  INV_X1 U7343 ( .A(SI_25_), .ZN(n9621) );
  NAND2_X1 U7344 ( .A1(n6294), .A2(n9621), .ZN(n6316) );
  INV_X1 U7345 ( .A(n6294), .ZN(n6295) );
  NAND2_X1 U7346 ( .A1(n6295), .A2(SI_25_), .ZN(n6296) );
  NAND2_X1 U7347 ( .A1(n6316), .A2(n6296), .ZN(n6317) );
  NAND2_X1 U7348 ( .A1(n8593), .A2(n7005), .ZN(n6298) );
  OR2_X1 U7349 ( .A1(n7015), .A2(n9526), .ZN(n6297) );
  NAND2_X1 U7350 ( .A1(n10471), .A2(n6373), .ZN(n6311) );
  INV_X1 U7351 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7352 ( .A1(n6300), .A2(n6299), .ZN(n6301) );
  NAND2_X1 U7353 ( .A1(n10327), .A2(n6424), .ZN(n6309) );
  INV_X1 U7354 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7355 ( .A1(n6302), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7356 ( .A1(n6303), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6304) );
  OAI211_X1 U7357 ( .C1(n6422), .C2(n6306), .A(n6305), .B(n6304), .ZN(n6307)
         );
  INV_X1 U7358 ( .A(n6307), .ZN(n6308) );
  NAND2_X1 U7359 ( .A1(n10158), .A2(n6388), .ZN(n6310) );
  NAND2_X1 U7360 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  XNOR2_X1 U7361 ( .A(n6312), .B(n5686), .ZN(n10050) );
  NOR2_X1 U7362 ( .A1(n10340), .A2(n6390), .ZN(n6313) );
  AOI21_X1 U7363 ( .B1(n10471), .B2(n6388), .A(n6313), .ZN(n10049) );
  INV_X1 U7364 ( .A(n10050), .ZN(n6315) );
  INV_X1 U7365 ( .A(n10049), .ZN(n6314) );
  INV_X1 U7366 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9525) );
  INV_X1 U7367 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6865) );
  MUX2_X1 U7368 ( .A(n9525), .B(n6865), .S(n6995), .Z(n6320) );
  INV_X1 U7369 ( .A(SI_26_), .ZN(n6319) );
  NAND2_X1 U7370 ( .A1(n6320), .A2(n6319), .ZN(n6348) );
  INV_X1 U7371 ( .A(n6320), .ZN(n6321) );
  NAND2_X1 U7372 ( .A1(n6321), .A2(SI_26_), .ZN(n6322) );
  NAND2_X1 U7373 ( .A1(n6348), .A2(n6322), .ZN(n6324) );
  NAND2_X1 U7374 ( .A1(n6323), .A2(n6324), .ZN(n6327) );
  INV_X1 U7375 ( .A(n6324), .ZN(n6325) );
  NAND2_X1 U7376 ( .A1(n6327), .A2(n6349), .ZN(n8649) );
  NAND2_X1 U7377 ( .A1(n8649), .A2(n7005), .ZN(n6329) );
  OR2_X1 U7378 ( .A1(n7015), .A2(n9525), .ZN(n6328) );
  INV_X1 U7379 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7380 ( .A1(n6332), .A2(n6331), .ZN(n6333) );
  NAND2_X1 U7381 ( .A1(n6376), .A2(n6333), .ZN(n10127) );
  INV_X1 U7382 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7383 ( .A1(n6302), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7384 ( .A1(n6303), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6335) );
  OAI211_X1 U7385 ( .C1(n6422), .C2(n6337), .A(n6336), .B(n6335), .ZN(n6338)
         );
  INV_X1 U7386 ( .A(n6338), .ZN(n6339) );
  NAND2_X1 U7387 ( .A1(n6340), .A2(n6339), .ZN(n10052) );
  OAI22_X1 U7388 ( .A1(n10314), .A2(n6341), .B1(n10323), .B2(n6384), .ZN(n6343) );
  XNOR2_X1 U7389 ( .A(n6343), .B(n6342), .ZN(n6345) );
  OAI22_X1 U7390 ( .A1(n10314), .A2(n6384), .B1(n10323), .B2(n6390), .ZN(n6344) );
  XNOR2_X1 U7391 ( .A(n6345), .B(n6344), .ZN(n10125) );
  INV_X1 U7392 ( .A(n6344), .ZN(n6347) );
  INV_X1 U7393 ( .A(n6345), .ZN(n6346) );
  MUX2_X1 U7394 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n6995), .Z(n6368) );
  INV_X1 U7395 ( .A(SI_27_), .ZN(n9418) );
  XNOR2_X1 U7396 ( .A(n6368), .B(n9418), .ZN(n6366) );
  NAND2_X1 U7397 ( .A1(n8690), .A2(n7005), .ZN(n6352) );
  INV_X1 U7398 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n6350) );
  OR2_X1 U7399 ( .A1(n7015), .A2(n6350), .ZN(n6351) );
  NAND2_X1 U7400 ( .A1(n10461), .A2(n6373), .ZN(n6360) );
  XNOR2_X1 U7401 ( .A(n6376), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U7402 ( .A1(n10291), .A2(n6424), .ZN(n6358) );
  INV_X1 U7403 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U7404 ( .A1(n6303), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7405 ( .A1(n6302), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6353) );
  OAI211_X1 U7406 ( .C1(n6422), .C2(n6355), .A(n6354), .B(n6353), .ZN(n6356)
         );
  INV_X1 U7407 ( .A(n6356), .ZN(n6357) );
  OR2_X1 U7408 ( .A1(n10305), .A2(n6384), .ZN(n6359) );
  NAND2_X1 U7409 ( .A1(n6360), .A2(n6359), .ZN(n6361) );
  XNOR2_X1 U7410 ( .A(n6361), .B(n5686), .ZN(n6364) );
  NOR2_X1 U7411 ( .A1(n10305), .A2(n6390), .ZN(n6362) );
  AOI21_X1 U7412 ( .B1(n10461), .B2(n6388), .A(n6362), .ZN(n6363) );
  NAND2_X1 U7413 ( .A1(n6364), .A2(n6363), .ZN(n6434) );
  OAI21_X1 U7414 ( .B1(n6364), .B2(n6363), .A(n6434), .ZN(n8698) );
  INV_X1 U7415 ( .A(n6365), .ZN(n6367) );
  NAND2_X1 U7416 ( .A1(n6367), .A2(n6366), .ZN(n6370) );
  NAND2_X1 U7417 ( .A1(n6368), .A2(SI_27_), .ZN(n6369) );
  NAND2_X1 U7418 ( .A1(n6370), .A2(n6369), .ZN(n6987) );
  MUX2_X1 U7419 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n6995), .Z(n6983) );
  XNOR2_X1 U7420 ( .A(n6983), .B(SI_28_), .ZN(n6986) );
  NAND2_X1 U7421 ( .A1(n9002), .A2(n7005), .ZN(n6372) );
  INV_X1 U7422 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9003) );
  OR2_X1 U7423 ( .A1(n7015), .A2(n9003), .ZN(n6371) );
  NAND2_X1 U7424 ( .A1(n10455), .A2(n6373), .ZN(n6386) );
  INV_X1 U7425 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8702) );
  INV_X1 U7426 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6374) );
  OAI21_X1 U7427 ( .B1(n6376), .B2(n8702), .A(n6374), .ZN(n6377) );
  NAND2_X1 U7428 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6375) );
  NAND2_X1 U7429 ( .A1(n8997), .A2(n6424), .ZN(n6383) );
  INV_X1 U7430 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U7431 ( .A1(n6303), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U7432 ( .A1(n6302), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6378) );
  OAI211_X1 U7433 ( .C1(n6422), .C2(n6380), .A(n6379), .B(n6378), .ZN(n6381)
         );
  INV_X1 U7434 ( .A(n6381), .ZN(n6382) );
  OR2_X1 U7435 ( .A1(n10297), .A2(n6384), .ZN(n6385) );
  NAND2_X1 U7436 ( .A1(n6386), .A2(n6385), .ZN(n6387) );
  XNOR2_X1 U7437 ( .A(n6387), .B(n5686), .ZN(n6392) );
  NAND2_X1 U7438 ( .A1(n10455), .A2(n6388), .ZN(n6389) );
  OAI21_X1 U7439 ( .B1(n10297), .B2(n6390), .A(n6389), .ZN(n6391) );
  XNOR2_X1 U7440 ( .A(n6392), .B(n6391), .ZN(n6414) );
  INV_X1 U7441 ( .A(n6414), .ZN(n6435) );
  NAND2_X1 U7442 ( .A1(n8594), .A2(P1_B_REG_SCAN_IN), .ZN(n6394) );
  MUX2_X1 U7443 ( .A(n6394), .B(P1_B_REG_SCAN_IN), .S(n6393), .Z(n6396) );
  NAND2_X1 U7444 ( .A1(n6396), .A2(n6395), .ZN(n7424) );
  OAI22_X1 U7445 ( .A1(n7424), .A2(P1_D_REG_1__SCAN_IN), .B1(n6395), .B2(n5032), .ZN(n7693) );
  NOR4_X1 U7446 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6405) );
  NOR4_X1 U7447 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6404) );
  OR4_X1 U7448 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6402) );
  NOR4_X1 U7449 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6400) );
  NOR4_X1 U7450 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6399) );
  NOR4_X1 U7451 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6398) );
  NOR4_X1 U7452 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6397) );
  NAND4_X1 U7453 ( .A1(n6400), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(n6401)
         );
  NOR4_X1 U7454 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        n6402), .A4(n6401), .ZN(n6403) );
  AND3_X1 U7455 ( .A1(n6405), .A2(n6404), .A3(n6403), .ZN(n6406) );
  NOR2_X1 U7456 ( .A1(n7424), .A2(n6406), .ZN(n7578) );
  NOR2_X1 U7457 ( .A1(n7693), .A2(n7578), .ZN(n6408) );
  INV_X1 U7458 ( .A(n7424), .ZN(n6407) );
  INV_X1 U7459 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9817) );
  INV_X1 U7460 ( .A(n6395), .ZN(n8650) );
  AND2_X1 U7461 ( .A1(n8650), .A2(n8416), .ZN(n7440) );
  NAND2_X1 U7462 ( .A1(n6408), .A2(n7702), .ZN(n6430) );
  INV_X1 U7463 ( .A(n6409), .ZN(n6410) );
  NAND2_X1 U7464 ( .A1(n6410), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6411) );
  XNOR2_X1 U7465 ( .A(n6411), .B(n9591), .ZN(n7495) );
  NAND2_X1 U7466 ( .A1(n7497), .A2(n7426), .ZN(n7577) );
  INV_X1 U7467 ( .A(n7718), .ZN(n8102) );
  NAND2_X1 U7468 ( .A1(n8291), .A2(n8102), .ZN(n7585) );
  INV_X1 U7469 ( .A(n7585), .ZN(n7705) );
  OR2_X1 U7470 ( .A1(n10739), .A2(n7271), .ZN(n6412) );
  NAND3_X1 U7471 ( .A1(n6435), .A2(n10143), .A3(n6434), .ZN(n6413) );
  NAND3_X1 U7472 ( .A1(n8701), .A2(n10143), .A3(n6414), .ZN(n6439) );
  OR2_X1 U7473 ( .A1(n7585), .A2(n8040), .ZN(n7700) );
  OR2_X1 U7474 ( .A1(n6426), .A2(n7700), .ZN(n6415) );
  INV_X1 U7475 ( .A(n8040), .ZN(n7717) );
  INV_X1 U7476 ( .A(n5036), .ZN(n7633) );
  OR2_X1 U7477 ( .A1(n10849), .A2(n7580), .ZN(n6417) );
  INV_X1 U7478 ( .A(n6418), .ZN(n10281) );
  INV_X1 U7479 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U7480 ( .A1(n6302), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U7481 ( .A1(n6303), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6419) );
  OAI211_X1 U7482 ( .C1(n6422), .C2(n6421), .A(n6420), .B(n6419), .ZN(n6423)
         );
  AOI21_X1 U7483 ( .B1(n10281), .B2(n6424), .A(n6423), .ZN(n8993) );
  INV_X1 U7484 ( .A(n8993), .ZN(n10157) );
  OR2_X1 U7485 ( .A1(n10851), .A2(n7580), .ZN(n6425) );
  NAND2_X1 U7486 ( .A1(n10157), .A2(n10147), .ZN(n6433) );
  NAND2_X1 U7487 ( .A1(n6430), .A2(n11083), .ZN(n7595) );
  AND2_X1 U7488 ( .A1(n7271), .A2(n7580), .ZN(n7576) );
  INV_X1 U7489 ( .A(n7576), .ZN(n6427) );
  AND3_X1 U7490 ( .A1(n6427), .A2(n7497), .A3(n7495), .ZN(n6428) );
  AOI21_X1 U7491 ( .B1(n7595), .B2(n6428), .A(P1_U3084), .ZN(n6431) );
  NOR2_X1 U7492 ( .A1(n7577), .A2(n7700), .ZN(n6429) );
  AND2_X1 U7493 ( .A1(n6430), .A2(n6429), .ZN(n7597) );
  AOI22_X1 U7494 ( .A1(n8997), .A2(n10152), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6432) );
  OAI211_X1 U7495 ( .C1(n10305), .C2(n10149), .A(n6433), .B(n6432), .ZN(n6437)
         );
  NOR3_X1 U7496 ( .A1(n6435), .A2(n10133), .A3(n6434), .ZN(n6436) );
  AOI211_X1 U7497 ( .C1(n10455), .C2(n10131), .A(n6437), .B(n6436), .ZN(n6438)
         );
  NAND3_X1 U7498 ( .A1(n5072), .A2(n6439), .A3(n6438), .ZN(P1_U3218) );
  INV_X1 U7499 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6442) );
  NAND4_X1 U7500 ( .A1(n5112), .A2(n6917), .A3(n6945), .A4(n6442), .ZN(n6448)
         );
  NOR2_X1 U7501 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6446) );
  NOR2_X1 U7502 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6445) );
  NOR2_X1 U7503 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6444) );
  NOR2_X1 U7504 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6443) );
  NAND4_X1 U7505 ( .A1(n6446), .A2(n6445), .A3(n6444), .A4(n6443), .ZN(n6447)
         );
  NOR2_X1 U7506 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  NAND2_X1 U7507 ( .A1(n6451), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6452) );
  INV_X1 U7508 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U7509 ( .A1(n6455), .A2(n6453), .ZN(n6474) );
  INV_X1 U7510 ( .A(n6474), .ZN(n6454) );
  NAND2_X1 U7511 ( .A1(n6475), .A2(n6454), .ZN(n6477) );
  INV_X1 U7512 ( .A(n6457), .ZN(n6458) );
  INV_X1 U7513 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6459) );
  INV_X1 U7514 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6690) );
  INV_X1 U7515 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6703) );
  NAND3_X1 U7516 ( .A1(n6690), .A2(n6703), .A3(n6706), .ZN(n6460) );
  INV_X1 U7517 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6463) );
  INV_X1 U7518 ( .A(n6465), .ZN(n6464) );
  NAND3_X1 U7519 ( .A1(n6464), .A2(n6466), .A3(n5112), .ZN(n6467) );
  NAND2_X1 U7520 ( .A1(n6465), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6751) );
  INV_X1 U7521 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6466) );
  XNOR2_X2 U7522 ( .A(n6470), .B(n6469), .ZN(n9846) );
  NAND2_X1 U7523 ( .A1(n6947), .A2(n9846), .ZN(n7823) );
  NAND2_X1 U7524 ( .A1(n6467), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U7525 ( .A1(n7823), .A2(n8201), .ZN(n6473) );
  XNOR2_X1 U7526 ( .A(n6472), .B(n6471), .ZN(n6488) );
  INV_X1 U7527 ( .A(n6488), .ZN(n7830) );
  NAND2_X1 U7528 ( .A1(n6478), .A2(n10002), .ZN(n6479) );
  NAND2_X1 U7529 ( .A1(n5060), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7530 ( .A1(n6549), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7531 ( .A1(n6533), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U7532 ( .A1(n6550), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U7533 ( .A1(n9159), .A2(n8780), .ZN(n6498) );
  XNOR2_X1 U7534 ( .A(n6497), .B(n6498), .ZN(n9053) );
  NAND2_X1 U7535 ( .A1(n6550), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U7536 ( .A1(n6549), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U7537 ( .A1(n5060), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U7538 ( .A1(n6533), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U7539 ( .A1(n6995), .A2(SI_0_), .ZN(n6494) );
  INV_X1 U7540 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U7541 ( .A1(n6494), .A2(n6493), .ZN(n6496) );
  AND2_X1 U7542 ( .A1(n6496), .A2(n6495), .ZN(n10014) );
  NAND2_X1 U7543 ( .A1(n7959), .A2(n6906), .ZN(n9052) );
  INV_X1 U7544 ( .A(n6497), .ZN(n6499) );
  NAND2_X1 U7545 ( .A1(n6499), .A2(n6498), .ZN(n6500) );
  NAND2_X1 U7546 ( .A1(n6549), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U7547 ( .A1(n6550), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U7548 ( .A1(n6533), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6501) );
  NOR2_X1 U7549 ( .A1(n8189), .A2(n6521), .ZN(n6514) );
  OR2_X1 U7550 ( .A1(n6457), .A2(n10002), .ZN(n6507) );
  INV_X1 U7551 ( .A(n6507), .ZN(n6505) );
  NAND2_X1 U7552 ( .A1(n6505), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n6508) );
  INV_X1 U7553 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U7554 ( .A1(n6507), .A2(n6506), .ZN(n6524) );
  INV_X1 U7555 ( .A(n10683), .ZN(n7414) );
  AND2_X1 U7556 ( .A1(n7404), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U7557 ( .A1(n7306), .A2(n6509), .ZN(n6513) );
  INV_X1 U7558 ( .A(n7422), .ZN(n6510) );
  OAI211_X1 U7559 ( .C1(n7306), .C2(n7414), .A(n6513), .B(n6512), .ZN(n8188)
         );
  XNOR2_X1 U7560 ( .A(n8190), .B(n6906), .ZN(n8046) );
  NAND2_X1 U7561 ( .A1(n6514), .A2(n8046), .ZN(n6516) );
  OR2_X1 U7562 ( .A1(n6514), .A2(n8046), .ZN(n6515) );
  INV_X1 U7563 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U7564 ( .A1(n6550), .A2(n6535), .ZN(n6520) );
  NAND2_X1 U7565 ( .A1(n6549), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U7566 ( .A1(n5060), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U7567 ( .A1(n6533), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6517) );
  NOR2_X1 U7568 ( .A1(n8240), .A2(n6521), .ZN(n6529) );
  NAND2_X1 U7569 ( .A1(n6768), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6528) );
  INV_X1 U7570 ( .A(n7409), .ZN(n6522) );
  AND2_X1 U7571 ( .A1(n6995), .A2(n6522), .ZN(n6523) );
  NAND2_X1 U7572 ( .A1(n7306), .A2(n6523), .ZN(n6526) );
  NAND2_X1 U7573 ( .A1(n6524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6525) );
  XNOR2_X1 U7574 ( .A(n6525), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7293) );
  INV_X1 U7575 ( .A(n7293), .ZN(n7408) );
  XNOR2_X1 U7576 ( .A(n8241), .B(n6906), .ZN(n6530) );
  NAND2_X1 U7577 ( .A1(n6529), .A2(n6530), .ZN(n6544) );
  INV_X1 U7578 ( .A(n6529), .ZN(n6531) );
  INV_X1 U7579 ( .A(n6530), .ZN(n8033) );
  NAND2_X1 U7580 ( .A1(n6531), .A2(n8033), .ZN(n6532) );
  AND2_X1 U7581 ( .A1(n6544), .A2(n6532), .ZN(n8043) );
  NAND2_X1 U7582 ( .A1(n6533), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U7583 ( .A1(n5060), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U7584 ( .A1(n6549), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6537) );
  INV_X1 U7585 ( .A(n6550), .ZN(n6534) );
  XNOR2_X1 U7586 ( .A(n6535), .B(P2_REG3_REG_4__SCAN_IN), .ZN(n10786) );
  NAND2_X1 U7587 ( .A1(n6550), .A2(n10786), .ZN(n6536) );
  OR2_X1 U7588 ( .A1(n8326), .A2(n6521), .ZN(n6547) );
  INV_X1 U7589 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7416) );
  OR2_X1 U7590 ( .A1(n5030), .A2(n7416), .ZN(n6543) );
  NAND2_X1 U7591 ( .A1(n6541), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6542) );
  XNOR2_X1 U7592 ( .A(n6542), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7295) );
  INV_X1 U7593 ( .A(n7295), .ZN(n7418) );
  XNOR2_X1 U7594 ( .A(n6906), .B(n10769), .ZN(n7967) );
  XNOR2_X1 U7595 ( .A(n6547), .B(n7967), .ZN(n8026) );
  INV_X1 U7596 ( .A(n6544), .ZN(n6545) );
  NOR2_X1 U7597 ( .A1(n8026), .A2(n6545), .ZN(n6546) );
  NAND2_X1 U7598 ( .A1(n6547), .A2(n7967), .ZN(n6548) );
  NAND2_X1 U7599 ( .A1(n6549), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7600 ( .A1(n5060), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6554) );
  NAND3_X1 U7601 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .A3(P2_REG3_REG_3__SCAN_IN), .ZN(n6566) );
  INV_X1 U7602 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U7603 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6551) );
  NAND2_X1 U7604 ( .A1(n9694), .A2(n6551), .ZN(n6552) );
  AND2_X1 U7605 ( .A1(n6566), .A2(n6552), .ZN(n10805) );
  NAND2_X1 U7606 ( .A1(n6550), .A2(n10805), .ZN(n6553) );
  NAND2_X1 U7607 ( .A1(n6533), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6556) );
  OR2_X1 U7608 ( .A1(n8250), .A2(n6521), .ZN(n6563) );
  OR2_X1 U7609 ( .A1(n6558), .A2(n10002), .ZN(n6559) );
  XNOR2_X1 U7610 ( .A(n6559), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7297) );
  INV_X1 U7611 ( .A(n7297), .ZN(n7413) );
  OR2_X1 U7612 ( .A1(n6540), .A2(n7412), .ZN(n6561) );
  INV_X1 U7613 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7411) );
  OR2_X1 U7614 ( .A1(n5030), .A2(n7411), .ZN(n6560) );
  OAI211_X1 U7615 ( .C1(n7306), .C2(n7413), .A(n6561), .B(n6560), .ZN(n10804)
         );
  INV_X1 U7616 ( .A(n10804), .ZN(n10817) );
  XNOR2_X1 U7617 ( .A(n10817), .B(n6906), .ZN(n6562) );
  XNOR2_X1 U7618 ( .A(n6563), .B(n6562), .ZN(n7966) );
  INV_X1 U7619 ( .A(n6562), .ZN(n7974) );
  INV_X1 U7620 ( .A(n6566), .ZN(n6564) );
  NAND2_X1 U7621 ( .A1(n6564), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6588) );
  INV_X1 U7622 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U7623 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  AND2_X1 U7624 ( .A1(n6588), .A2(n6567), .ZN(n9896) );
  NAND2_X1 U7625 ( .A1(n6550), .A2(n9896), .ZN(n6571) );
  NAND2_X1 U7626 ( .A1(n6549), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U7627 ( .A1(n6533), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U7628 ( .A1(n5060), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6568) );
  OR2_X1 U7629 ( .A1(n8449), .A2(n6521), .ZN(n6579) );
  NAND2_X1 U7630 ( .A1(n6572), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6582) );
  INV_X1 U7631 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6581) );
  XNOR2_X1 U7632 ( .A(n6582), .B(n6581), .ZN(n7433) );
  INV_X1 U7633 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6574) );
  OR2_X1 U7634 ( .A1(n5030), .A2(n6574), .ZN(n6576) );
  OR2_X1 U7635 ( .A1(n6540), .A2(n7432), .ZN(n6575) );
  OAI211_X1 U7636 ( .C1(n7306), .C2(n7433), .A(n6576), .B(n6575), .ZN(n10832)
         );
  INV_X1 U7637 ( .A(n10832), .ZN(n8251) );
  XNOR2_X1 U7638 ( .A(n8251), .B(n6906), .ZN(n6577) );
  INV_X1 U7639 ( .A(n6577), .ZN(n6578) );
  NAND2_X1 U7640 ( .A1(n6579), .A2(n6578), .ZN(n6580) );
  NAND2_X1 U7641 ( .A1(n7979), .A2(n6580), .ZN(n7949) );
  NAND2_X1 U7642 ( .A1(n6582), .A2(n6581), .ZN(n6583) );
  NAND2_X1 U7643 ( .A1(n6583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6584) );
  XNOR2_X1 U7644 ( .A(n6584), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7320) );
  INV_X1 U7645 ( .A(n7320), .ZN(n7436) );
  NAND2_X1 U7646 ( .A1(n7434), .A2(n6511), .ZN(n6586) );
  INV_X1 U7647 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7435) );
  OR2_X1 U7648 ( .A1(n5030), .A2(n7435), .ZN(n6585) );
  OAI211_X1 U7649 ( .C1(n7306), .C2(n7436), .A(n6586), .B(n6585), .ZN(n10873)
         );
  XNOR2_X1 U7650 ( .A(n6907), .B(n10873), .ZN(n6595) );
  INV_X1 U7651 ( .A(n6588), .ZN(n6587) );
  NAND2_X1 U7652 ( .A1(n6587), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6601) );
  INV_X1 U7653 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U7654 ( .A1(n6588), .A2(n7951), .ZN(n6589) );
  AND2_X1 U7655 ( .A1(n6601), .A2(n6589), .ZN(n8452) );
  NAND2_X1 U7656 ( .A1(n6550), .A2(n8452), .ZN(n6594) );
  NAND2_X1 U7657 ( .A1(n6549), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U7658 ( .A1(n6885), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U7659 ( .A1(n6533), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6591) );
  NAND4_X1 U7660 ( .A1(n6594), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(n9891)
         );
  AND2_X1 U7661 ( .A1(n9891), .A2(n8780), .ZN(n6596) );
  NAND2_X1 U7662 ( .A1(n6595), .A2(n6596), .ZN(n6599) );
  INV_X1 U7663 ( .A(n6595), .ZN(n9039) );
  INV_X1 U7664 ( .A(n6596), .ZN(n6597) );
  NAND2_X1 U7665 ( .A1(n9039), .A2(n6597), .ZN(n6598) );
  NAND2_X1 U7666 ( .A1(n6599), .A2(n6598), .ZN(n7948) );
  INV_X1 U7667 ( .A(n6601), .ZN(n6600) );
  NAND2_X1 U7668 ( .A1(n6600), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6620) );
  INV_X1 U7669 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U7670 ( .A1(n6601), .A2(n9481), .ZN(n6602) );
  AND2_X1 U7671 ( .A1(n6620), .A2(n6602), .ZN(n10900) );
  NAND2_X1 U7672 ( .A1(n6550), .A2(n10900), .ZN(n6606) );
  NAND2_X1 U7673 ( .A1(n6549), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U7674 ( .A1(n6885), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U7675 ( .A1(n6533), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6603) );
  NOR2_X1 U7676 ( .A1(n8448), .A2(n6521), .ZN(n6612) );
  NAND2_X1 U7677 ( .A1(n7444), .A2(n6511), .ZN(n6610) );
  NAND2_X1 U7678 ( .A1(n6607), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6608) );
  XNOR2_X1 U7679 ( .A(n6608), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7370) );
  AOI22_X1 U7680 ( .A1(n6768), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6767), .B2(
        n7370), .ZN(n6609) );
  NAND2_X1 U7681 ( .A1(n6610), .A2(n6609), .ZN(n10898) );
  XNOR2_X1 U7682 ( .A(n10898), .B(n6907), .ZN(n6611) );
  NAND2_X1 U7683 ( .A1(n6612), .A2(n6611), .ZN(n6626) );
  INV_X1 U7684 ( .A(n6611), .ZN(n8136) );
  INV_X1 U7685 ( .A(n6612), .ZN(n6613) );
  NAND2_X1 U7686 ( .A1(n8136), .A2(n6613), .ZN(n6614) );
  NAND2_X1 U7687 ( .A1(n7450), .A2(n6511), .ZN(n6617) );
  OR2_X1 U7688 ( .A1(n6615), .A2(n10002), .ZN(n6632) );
  XNOR2_X1 U7689 ( .A(n6632), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7394) );
  AOI22_X1 U7690 ( .A1(n6768), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6767), .B2(
        n7394), .ZN(n6616) );
  NAND2_X1 U7691 ( .A1(n6617), .A2(n6616), .ZN(n8423) );
  XNOR2_X1 U7692 ( .A(n8423), .B(n6906), .ZN(n6630) );
  INV_X1 U7693 ( .A(n6620), .ZN(n6618) );
  NAND2_X1 U7694 ( .A1(n6618), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6636) );
  INV_X1 U7695 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U7696 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  AND2_X1 U7697 ( .A1(n6636), .A2(n6621), .ZN(n8267) );
  NAND2_X1 U7698 ( .A1(n6550), .A2(n8267), .ZN(n6625) );
  NAND2_X1 U7699 ( .A1(n6549), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6624) );
  NAND2_X1 U7700 ( .A1(n6885), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U7701 ( .A1(n6533), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6622) );
  NOR2_X1 U7702 ( .A1(n10938), .A2(n6521), .ZN(n6628) );
  XNOR2_X1 U7703 ( .A(n6630), .B(n6628), .ZN(n8147) );
  AND2_X1 U7704 ( .A1(n8147), .A2(n6626), .ZN(n6627) );
  NAND2_X1 U7705 ( .A1(n8135), .A2(n6627), .ZN(n8139) );
  INV_X1 U7706 ( .A(n6628), .ZN(n6629) );
  NAND2_X1 U7707 ( .A1(n6630), .A2(n6629), .ZN(n6631) );
  NAND2_X1 U7708 ( .A1(n8139), .A2(n6631), .ZN(n8232) );
  NAND2_X1 U7709 ( .A1(n7536), .A2(n6511), .ZN(n6635) );
  NAND2_X1 U7710 ( .A1(n6632), .A2(n5360), .ZN(n6633) );
  NAND2_X1 U7711 ( .A1(n6633), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6647) );
  XNOR2_X1 U7712 ( .A(n6647), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7873) );
  AOI22_X1 U7713 ( .A1(n6768), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6767), .B2(
        n7873), .ZN(n6634) );
  NAND2_X1 U7714 ( .A1(n6635), .A2(n6634), .ZN(n10932) );
  XNOR2_X1 U7715 ( .A(n10932), .B(n6907), .ZN(n6642) );
  NAND2_X1 U7716 ( .A1(n6549), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U7717 ( .A1(n6636), .A2(n9672), .ZN(n6637) );
  AND2_X1 U7718 ( .A1(n6652), .A2(n6637), .ZN(n10961) );
  NAND2_X1 U7719 ( .A1(n6550), .A2(n10961), .ZN(n6640) );
  NAND2_X1 U7720 ( .A1(n6533), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U7721 ( .A1(n6885), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6638) );
  NOR2_X1 U7722 ( .A1(n8418), .A2(n6521), .ZN(n6643) );
  NAND2_X1 U7723 ( .A1(n6642), .A2(n6643), .ZN(n6646) );
  INV_X1 U7724 ( .A(n6642), .ZN(n8404) );
  INV_X1 U7725 ( .A(n6643), .ZN(n6644) );
  NAND2_X1 U7726 ( .A1(n8404), .A2(n6644), .ZN(n6645) );
  NAND2_X1 U7727 ( .A1(n6646), .A2(n6645), .ZN(n8231) );
  NAND2_X1 U7728 ( .A1(n7555), .A2(n6511), .ZN(n6651) );
  NAND2_X1 U7729 ( .A1(n6647), .A2(n5361), .ZN(n6648) );
  NAND2_X1 U7730 ( .A1(n6648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6649) );
  XNOR2_X1 U7731 ( .A(n6649), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7991) );
  AOI22_X1 U7732 ( .A1(n6768), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6767), .B2(
        n7991), .ZN(n6650) );
  NAND2_X1 U7733 ( .A1(n6651), .A2(n6650), .ZN(n10974) );
  XNOR2_X1 U7734 ( .A(n10974), .B(n6907), .ZN(n6658) );
  NAND2_X1 U7735 ( .A1(n6652), .A2(n7866), .ZN(n6653) );
  AND2_X1 U7736 ( .A1(n6667), .A2(n6653), .ZN(n8440) );
  NAND2_X1 U7737 ( .A1(n6550), .A2(n8440), .ZN(n6657) );
  NAND2_X1 U7738 ( .A1(n6549), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U7739 ( .A1(n6885), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U7740 ( .A1(n6533), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6654) );
  NOR2_X1 U7741 ( .A1(n10940), .A2(n6521), .ZN(n6659) );
  NAND2_X1 U7742 ( .A1(n6658), .A2(n6659), .ZN(n6673) );
  INV_X1 U7743 ( .A(n6658), .ZN(n8478) );
  INV_X1 U7744 ( .A(n6659), .ZN(n6660) );
  NAND2_X1 U7745 ( .A1(n8478), .A2(n6660), .ZN(n6661) );
  AND2_X1 U7746 ( .A1(n6673), .A2(n6661), .ZN(n8401) );
  NAND2_X1 U7747 ( .A1(n7624), .A2(n6511), .ZN(n6665) );
  NAND2_X1 U7748 ( .A1(n6662), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6663) );
  XNOR2_X1 U7749 ( .A(n6663), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8015) );
  AOI22_X1 U7750 ( .A1(n6768), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6767), .B2(
        n8015), .ZN(n6664) );
  NAND2_X1 U7751 ( .A1(n6665), .A2(n6664), .ZN(n8535) );
  XNOR2_X1 U7752 ( .A(n8535), .B(n6906), .ZN(n8717) );
  NAND2_X1 U7753 ( .A1(n6549), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6672) );
  INV_X1 U7754 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9482) );
  NAND2_X1 U7755 ( .A1(n6667), .A2(n9482), .ZN(n6668) );
  AND2_X1 U7756 ( .A1(n6681), .A2(n6668), .ZN(n8481) );
  NAND2_X1 U7757 ( .A1(n6550), .A2(n8481), .ZN(n6671) );
  NAND2_X1 U7758 ( .A1(n6533), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6670) );
  NAND2_X1 U7759 ( .A1(n6885), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6669) );
  NOR2_X1 U7760 ( .A1(n8716), .A2(n6521), .ZN(n6675) );
  XNOR2_X1 U7761 ( .A(n8717), .B(n6675), .ZN(n8490) );
  AND2_X1 U7762 ( .A1(n8490), .A2(n6673), .ZN(n6674) );
  INV_X1 U7763 ( .A(n6675), .ZN(n6676) );
  NAND2_X1 U7764 ( .A1(n8717), .A2(n6676), .ZN(n6677) );
  NAND2_X1 U7765 ( .A1(n8720), .A2(n6677), .ZN(n6687) );
  NAND2_X1 U7766 ( .A1(n7657), .A2(n6511), .ZN(n6679) );
  NAND2_X1 U7767 ( .A1(n5077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6691) );
  XNOR2_X1 U7768 ( .A(n6691), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8110) );
  AOI22_X1 U7769 ( .A1(n6768), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6767), .B2(
        n8110), .ZN(n6678) );
  NAND2_X1 U7770 ( .A1(n6679), .A2(n6678), .ZN(n8714) );
  XNOR2_X1 U7771 ( .A(n8714), .B(n6906), .ZN(n8745) );
  NAND2_X1 U7772 ( .A1(n6549), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6686) );
  INV_X1 U7773 ( .A(n6681), .ZN(n6680) );
  INV_X1 U7774 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U7775 ( .A1(n6681), .A2(n9704), .ZN(n6682) );
  AND2_X1 U7776 ( .A1(n6695), .A2(n6682), .ZN(n8710) );
  NAND2_X1 U7777 ( .A1(n6550), .A2(n8710), .ZN(n6685) );
  NAND2_X1 U7778 ( .A1(n6533), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U7779 ( .A1(n6885), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6683) );
  NOR2_X1 U7780 ( .A1(n8744), .A2(n6521), .ZN(n6688) );
  XNOR2_X1 U7781 ( .A(n8745), .B(n6688), .ZN(n8715) );
  INV_X1 U7782 ( .A(n6688), .ZN(n6689) );
  NAND2_X1 U7783 ( .A1(n7659), .A2(n6511), .ZN(n6694) );
  NAND2_X1 U7784 ( .A1(n6691), .A2(n6690), .ZN(n6692) );
  NAND2_X1 U7785 ( .A1(n6692), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6704) );
  XNOR2_X1 U7786 ( .A(n6704), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9170) );
  AOI22_X1 U7787 ( .A1(n6768), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6767), .B2(
        n9170), .ZN(n6693) );
  XNOR2_X1 U7788 ( .A(n11051), .B(n6907), .ZN(n8729) );
  INV_X1 U7789 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U7790 ( .A1(n6695), .A2(n9472), .ZN(n6696) );
  AND2_X1 U7791 ( .A1(n6711), .A2(n6696), .ZN(n8738) );
  NAND2_X1 U7792 ( .A1(n6550), .A2(n8738), .ZN(n6700) );
  NAND2_X1 U7793 ( .A1(n6549), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U7794 ( .A1(n6885), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U7795 ( .A1(n6533), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6697) );
  NAND4_X1 U7796 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n9150)
         );
  NAND2_X1 U7797 ( .A1(n9150), .A2(n8780), .ZN(n6701) );
  XNOR2_X1 U7798 ( .A(n8729), .B(n6701), .ZN(n8743) );
  INV_X1 U7799 ( .A(n8729), .ZN(n6702) );
  NAND2_X1 U7800 ( .A1(n7686), .A2(n6511), .ZN(n6709) );
  NAND2_X1 U7801 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  NAND2_X1 U7802 ( .A1(n6705), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6707) );
  XNOR2_X1 U7803 ( .A(n6707), .B(n6706), .ZN(n9187) );
  INV_X1 U7804 ( .A(n9187), .ZN(n9168) );
  AOI22_X1 U7805 ( .A1(n6768), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6767), .B2(
        n9168), .ZN(n6708) );
  XNOR2_X1 U7806 ( .A(n8735), .B(n6906), .ZN(n8671) );
  INV_X1 U7807 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U7808 ( .A1(n6711), .A2(n9514), .ZN(n6712) );
  AND2_X1 U7809 ( .A1(n6725), .A2(n6712), .ZN(n8727) );
  NAND2_X1 U7810 ( .A1(n6550), .A2(n8727), .ZN(n6716) );
  NAND2_X1 U7811 ( .A1(n6549), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6715) );
  NAND2_X1 U7812 ( .A1(n6533), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U7813 ( .A1(n6885), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6713) );
  NOR2_X1 U7814 ( .A1(n8670), .A2(n6521), .ZN(n6718) );
  XNOR2_X1 U7815 ( .A(n8671), .B(n6718), .ZN(n8731) );
  NAND2_X1 U7816 ( .A1(n6717), .A2(n8731), .ZN(n8737) );
  INV_X1 U7817 ( .A(n6718), .ZN(n6719) );
  NAND2_X1 U7818 ( .A1(n8671), .A2(n6719), .ZN(n6720) );
  NAND2_X1 U7819 ( .A1(n8737), .A2(n6720), .ZN(n6731) );
  NAND2_X1 U7820 ( .A1(n7690), .A2(n6511), .ZN(n6724) );
  OR2_X1 U7821 ( .A1(n6721), .A2(n10002), .ZN(n6722) );
  XNOR2_X1 U7822 ( .A(n6722), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9202) );
  AOI22_X1 U7823 ( .A1(n6768), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6767), .B2(
        n9202), .ZN(n6723) );
  XNOR2_X1 U7824 ( .A(n8687), .B(n6906), .ZN(n6732) );
  NAND2_X1 U7825 ( .A1(n6549), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6730) );
  INV_X1 U7826 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U7827 ( .A1(n6725), .A2(n9483), .ZN(n6726) );
  AND2_X1 U7828 ( .A1(n6741), .A2(n6726), .ZN(n8684) );
  NAND2_X1 U7829 ( .A1(n6550), .A2(n8684), .ZN(n6729) );
  NAND2_X1 U7830 ( .A1(n6533), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U7831 ( .A1(n6885), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6727) );
  NAND4_X1 U7832 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n9248)
         );
  NAND2_X1 U7833 ( .A1(n9248), .A2(n8780), .ZN(n6733) );
  XNOR2_X1 U7834 ( .A(n6732), .B(n6733), .ZN(n8669) );
  INV_X1 U7835 ( .A(n6732), .ZN(n6734) );
  NAND2_X1 U7836 ( .A1(n6734), .A2(n6733), .ZN(n6735) );
  NAND2_X1 U7837 ( .A1(n7796), .A2(n6511), .ZN(n6738) );
  NAND2_X1 U7838 ( .A1(n5119), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6736) );
  XNOR2_X1 U7839 ( .A(n6736), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9221) );
  AOI22_X1 U7840 ( .A1(n6768), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6767), .B2(
        n9221), .ZN(n6737) );
  XNOR2_X1 U7841 ( .A(n9977), .B(n6907), .ZN(n6747) );
  NAND2_X1 U7842 ( .A1(n6549), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6746) );
  INV_X1 U7843 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U7844 ( .A1(n6741), .A2(n6740), .ZN(n6742) );
  AND2_X1 U7845 ( .A1(n6755), .A2(n6742), .ZN(n9881) );
  NAND2_X1 U7846 ( .A1(n6550), .A2(n9881), .ZN(n6745) );
  NAND2_X1 U7847 ( .A1(n6533), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U7848 ( .A1(n6885), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6743) );
  NAND4_X1 U7849 ( .A1(n6746), .A2(n6745), .A3(n6744), .A4(n6743), .ZN(n9862)
         );
  AND2_X1 U7850 ( .A1(n9862), .A2(n8780), .ZN(n6748) );
  NAND2_X1 U7851 ( .A1(n6747), .A2(n6748), .ZN(n6761) );
  INV_X1 U7852 ( .A(n6747), .ZN(n9123) );
  INV_X1 U7853 ( .A(n6748), .ZN(n6749) );
  NAND2_X1 U7854 ( .A1(n9123), .A2(n6749), .ZN(n6750) );
  NAND2_X1 U7855 ( .A1(n6761), .A2(n6750), .ZN(n9088) );
  NAND2_X1 U7856 ( .A1(n7864), .A2(n6511), .ZN(n6753) );
  XNOR2_X1 U7857 ( .A(n6751), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9232) );
  AOI22_X1 U7858 ( .A1(n6768), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6767), .B2(
        n9232), .ZN(n6752) );
  XNOR2_X1 U7859 ( .A(n9970), .B(n6906), .ZN(n6765) );
  INV_X1 U7860 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U7861 ( .A1(n6755), .A2(n6754), .ZN(n6756) );
  AND2_X1 U7862 ( .A1(n6773), .A2(n6756), .ZN(n9857) );
  NAND2_X1 U7863 ( .A1(n6550), .A2(n9857), .ZN(n6760) );
  NAND2_X1 U7864 ( .A1(n6549), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U7865 ( .A1(n6885), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U7866 ( .A1(n6533), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6757) );
  NOR2_X1 U7867 ( .A1(n9876), .A2(n6521), .ZN(n6763) );
  XNOR2_X1 U7868 ( .A(n6765), .B(n6763), .ZN(n9124) );
  AND2_X1 U7869 ( .A1(n9124), .A2(n6761), .ZN(n6762) );
  INV_X1 U7870 ( .A(n6763), .ZN(n6764) );
  NAND2_X1 U7871 ( .A1(n6765), .A2(n6764), .ZN(n6766) );
  NAND2_X1 U7872 ( .A1(n9120), .A2(n6766), .ZN(n9027) );
  NAND2_X1 U7873 ( .A1(n7956), .A2(n6511), .ZN(n6770) );
  AOI22_X1 U7874 ( .A1(n6768), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10902), 
        .B2(n6767), .ZN(n6769) );
  XNOR2_X1 U7875 ( .A(n9967), .B(n6906), .ZN(n6781) );
  INV_X1 U7876 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U7877 ( .A1(n6773), .A2(n6772), .ZN(n6774) );
  NAND2_X1 U7878 ( .A1(n6787), .A2(n6774), .ZN(n9848) );
  INV_X1 U7879 ( .A(n6885), .ZN(n6776) );
  INV_X1 U7880 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n6775) );
  OAI22_X1 U7881 ( .A1(n9848), .A2(n6534), .B1(n6776), .B2(n6775), .ZN(n6779)
         );
  INV_X1 U7882 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9233) );
  INV_X1 U7883 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6777) );
  OAI22_X1 U7884 ( .A1(n6969), .A2(n9233), .B1(n6590), .B2(n6777), .ZN(n6778)
         );
  NAND2_X1 U7885 ( .A1(n9863), .A2(n8780), .ZN(n6782) );
  AND2_X1 U7886 ( .A1(n6781), .A2(n6782), .ZN(n6780) );
  INV_X1 U7887 ( .A(n6781), .ZN(n9031) );
  INV_X1 U7888 ( .A(n6782), .ZN(n6783) );
  NAND2_X1 U7889 ( .A1(n9031), .A2(n6783), .ZN(n9028) );
  NAND2_X1 U7890 ( .A1(n8039), .A2(n6511), .ZN(n6785) );
  OR2_X1 U7891 ( .A1(n5030), .A2(n8149), .ZN(n6784) );
  XNOR2_X1 U7892 ( .A(n9960), .B(n6907), .ZN(n6792) );
  INV_X1 U7893 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U7894 ( .A1(n6787), .A2(n9703), .ZN(n6788) );
  NAND2_X1 U7895 ( .A1(n6799), .A2(n6788), .ZN(n9402) );
  OR2_X1 U7896 ( .A1(n9402), .A2(n6534), .ZN(n6791) );
  AOI22_X1 U7897 ( .A1(n6549), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6533), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U7898 ( .A1(n6885), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6789) );
  NOR2_X1 U7899 ( .A1(n9842), .A2(n6521), .ZN(n6793) );
  NAND2_X1 U7900 ( .A1(n6792), .A2(n6793), .ZN(n6796) );
  INV_X1 U7901 ( .A(n6792), .ZN(n9061) );
  INV_X1 U7902 ( .A(n6793), .ZN(n6794) );
  NAND2_X1 U7903 ( .A1(n9061), .A2(n6794), .ZN(n6795) );
  AND2_X1 U7904 ( .A1(n6796), .A2(n6795), .ZN(n9103) );
  NAND2_X1 U7905 ( .A1(n8100), .A2(n6511), .ZN(n6798) );
  INV_X1 U7906 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8119) );
  OR2_X1 U7907 ( .A1(n5030), .A2(n8119), .ZN(n6797) );
  XNOR2_X1 U7908 ( .A(n9955), .B(n6907), .ZN(n6804) );
  INV_X1 U7909 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6803) );
  INV_X1 U7910 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9681) );
  NAND2_X1 U7911 ( .A1(n6799), .A2(n9681), .ZN(n6800) );
  NAND2_X1 U7912 ( .A1(n6811), .A2(n6800), .ZN(n9386) );
  OR2_X1 U7913 ( .A1(n9386), .A2(n6534), .ZN(n6802) );
  AOI22_X1 U7914 ( .A1(n6533), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n5060), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6801) );
  OAI211_X1 U7915 ( .C1(n6969), .C2(n6803), .A(n6802), .B(n6801), .ZN(n9408)
         );
  AND2_X1 U7916 ( .A1(n9408), .A2(n8780), .ZN(n6805) );
  NAND2_X1 U7917 ( .A1(n6804), .A2(n6805), .ZN(n6819) );
  INV_X1 U7918 ( .A(n6804), .ZN(n9110) );
  INV_X1 U7919 ( .A(n6805), .ZN(n6806) );
  NAND2_X1 U7920 ( .A1(n9110), .A2(n6806), .ZN(n6807) );
  AND2_X1 U7921 ( .A1(n6819), .A2(n6807), .ZN(n9059) );
  NAND2_X1 U7922 ( .A1(n6808), .A2(n9059), .ZN(n9062) );
  NAND2_X1 U7923 ( .A1(n8290), .A2(n6511), .ZN(n6810) );
  OR2_X1 U7924 ( .A1(n5030), .A2(n8292), .ZN(n6809) );
  XNOR2_X1 U7925 ( .A(n9950), .B(n6907), .ZN(n6823) );
  INV_X1 U7926 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U7927 ( .A1(n6811), .A2(n9113), .ZN(n6812) );
  AND2_X1 U7928 ( .A1(n6828), .A2(n6812), .ZN(n9373) );
  NAND2_X1 U7929 ( .A1(n9373), .A2(n6550), .ZN(n6818) );
  INV_X1 U7930 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6815) );
  NAND2_X1 U7931 ( .A1(n6885), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U7932 ( .A1(n6533), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6813) );
  OAI211_X1 U7933 ( .C1(n6815), .C2(n6969), .A(n6814), .B(n6813), .ZN(n6816)
         );
  INV_X1 U7934 ( .A(n6816), .ZN(n6817) );
  NAND2_X1 U7935 ( .A1(n9393), .A2(n8780), .ZN(n6824) );
  XNOR2_X1 U7936 ( .A(n6823), .B(n6824), .ZN(n9111) );
  AND2_X1 U7937 ( .A1(n9111), .A2(n6819), .ZN(n6820) );
  NAND2_X1 U7938 ( .A1(n8298), .A2(n6511), .ZN(n6822) );
  OR2_X1 U7939 ( .A1(n5030), .A2(n8300), .ZN(n6821) );
  XNOR2_X1 U7940 ( .A(n9945), .B(n6907), .ZN(n6837) );
  INV_X1 U7941 ( .A(n6823), .ZN(n6825) );
  NAND2_X1 U7942 ( .A1(n6825), .A2(n6824), .ZN(n6836) );
  AND2_X1 U7943 ( .A1(n6837), .A2(n6836), .ZN(n6826) );
  INV_X1 U7944 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U7945 ( .A1(n6828), .A2(n9473), .ZN(n6829) );
  NAND2_X1 U7946 ( .A1(n6850), .A2(n6829), .ZN(n9364) );
  OR2_X1 U7947 ( .A1(n9364), .A2(n6534), .ZN(n6835) );
  INV_X1 U7948 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U7949 ( .A1(n6885), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U7950 ( .A1(n6533), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6830) );
  OAI211_X1 U7951 ( .C1(n6832), .C2(n6969), .A(n6831), .B(n6830), .ZN(n6833)
         );
  INV_X1 U7952 ( .A(n6833), .ZN(n6834) );
  INV_X1 U7953 ( .A(n9378), .ZN(n9148) );
  NAND2_X1 U7954 ( .A1(n9148), .A2(n8780), .ZN(n9018) );
  INV_X1 U7955 ( .A(n6837), .ZN(n6838) );
  NAND2_X1 U7956 ( .A1(n8593), .A2(n6511), .ZN(n6840) );
  OR2_X1 U7957 ( .A1(n5030), .A2(n8595), .ZN(n6839) );
  XNOR2_X1 U7958 ( .A(n9936), .B(n6907), .ZN(n9075) );
  INV_X1 U7959 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6842) );
  NAND2_X1 U7960 ( .A1(n6852), .A2(n6842), .ZN(n6843) );
  INV_X1 U7961 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U7962 ( .A1(n6533), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U7963 ( .A1(n5060), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6844) );
  OAI211_X1 U7964 ( .C1(n6846), .C2(n6969), .A(n6845), .B(n6844), .ZN(n6847)
         );
  OR2_X1 U7965 ( .A1(n9350), .A2(n6521), .ZN(n9074) );
  INV_X1 U7966 ( .A(n9074), .ZN(n6860) );
  NAND2_X1 U7967 ( .A1(n8414), .A2(n6511), .ZN(n6849) );
  INV_X1 U7968 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8460) );
  OR2_X1 U7969 ( .A1(n5030), .A2(n8460), .ZN(n6848) );
  XNOR2_X1 U7970 ( .A(n9939), .B(n6907), .ZN(n9070) );
  INV_X1 U7971 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9692) );
  NAND2_X1 U7972 ( .A1(n6850), .A2(n9692), .ZN(n6851) );
  NAND2_X1 U7973 ( .A1(n6852), .A2(n6851), .ZN(n9342) );
  OR2_X1 U7974 ( .A1(n9342), .A2(n6534), .ZN(n6858) );
  INV_X1 U7975 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U7976 ( .A1(n6885), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6854) );
  NAND2_X1 U7977 ( .A1(n6533), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6853) );
  OAI211_X1 U7978 ( .C1(n6855), .C2(n6969), .A(n6854), .B(n6853), .ZN(n6856)
         );
  INV_X1 U7979 ( .A(n6856), .ZN(n6857) );
  NOR2_X1 U7980 ( .A1(n9092), .A2(n6521), .ZN(n9071) );
  OAI22_X1 U7981 ( .A1(n9075), .A2(n6860), .B1(n9070), .B2(n9071), .ZN(n6864)
         );
  NAND2_X1 U7982 ( .A1(n9070), .A2(n9071), .ZN(n6859) );
  NAND2_X1 U7983 ( .A1(n6859), .A2(n9074), .ZN(n6862) );
  INV_X1 U7984 ( .A(n6859), .ZN(n6861) );
  AOI22_X1 U7985 ( .A1(n9075), .A2(n6862), .B1(n6861), .B2(n6860), .ZN(n6863)
         );
  NAND2_X1 U7986 ( .A1(n8649), .A2(n6511), .ZN(n6867) );
  OR2_X1 U7987 ( .A1(n5030), .A2(n6865), .ZN(n6866) );
  XNOR2_X1 U7988 ( .A(n9238), .B(n6906), .ZN(n6877) );
  INV_X1 U7989 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9713) );
  NAND2_X1 U7990 ( .A1(n6869), .A2(n9713), .ZN(n6870) );
  NAND2_X1 U7991 ( .A1(n6898), .A2(n6870), .ZN(n9325) );
  OR2_X1 U7992 ( .A1(n9325), .A2(n6534), .ZN(n6876) );
  INV_X1 U7993 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U7994 ( .A1(n6533), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U7995 ( .A1(n6885), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6871) );
  OAI211_X1 U7996 ( .C1(n6873), .C2(n6969), .A(n6872), .B(n6871), .ZN(n6874)
         );
  INV_X1 U7997 ( .A(n6874), .ZN(n6875) );
  AND2_X1 U7998 ( .A1(n9260), .A2(n8780), .ZN(n6878) );
  NAND2_X1 U7999 ( .A1(n6877), .A2(n6878), .ZN(n6881) );
  INV_X1 U8000 ( .A(n6877), .ZN(n9007) );
  INV_X1 U8001 ( .A(n6878), .ZN(n6879) );
  NAND2_X1 U8002 ( .A1(n9007), .A2(n6879), .ZN(n6880) );
  AND2_X1 U8003 ( .A1(n6881), .A2(n6880), .ZN(n9138) );
  NAND2_X1 U8004 ( .A1(n9137), .A2(n9138), .ZN(n9136) );
  NAND2_X1 U8005 ( .A1(n9136), .A2(n6881), .ZN(n6895) );
  NAND2_X1 U8006 ( .A1(n8690), .A2(n6511), .ZN(n6884) );
  INV_X1 U8007 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6882) );
  OR2_X1 U8008 ( .A1(n5030), .A2(n6882), .ZN(n6883) );
  XNOR2_X1 U8009 ( .A(n9924), .B(n6907), .ZN(n6890) );
  XNOR2_X1 U8010 ( .A(n6898), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9303) );
  INV_X1 U8011 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6888) );
  NAND2_X1 U8012 ( .A1(n6533), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U8013 ( .A1(n6885), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6886) );
  OAI211_X1 U8014 ( .C1(n6888), .C2(n6969), .A(n6887), .B(n6886), .ZN(n6889)
         );
  AOI21_X1 U8015 ( .B1(n9303), .B2(n6550), .A(n6889), .ZN(n9262) );
  NOR2_X1 U8016 ( .A1(n9262), .A2(n6521), .ZN(n6891) );
  NAND2_X1 U8017 ( .A1(n6890), .A2(n6891), .ZN(n6896) );
  INV_X1 U8018 ( .A(n6890), .ZN(n6893) );
  INV_X1 U8019 ( .A(n6891), .ZN(n6892) );
  NAND2_X1 U8020 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  AND2_X1 U8021 ( .A1(n6896), .A2(n6894), .ZN(n9005) );
  NAND2_X1 U8022 ( .A1(n6895), .A2(n9005), .ZN(n9008) );
  NAND2_X1 U8023 ( .A1(n9008), .A2(n6896), .ZN(n6912) );
  INV_X1 U8024 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9011) );
  INV_X1 U8025 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9680) );
  OAI21_X1 U8026 ( .B1(n6898), .B2(n9011), .A(n9680), .ZN(n6899) );
  NAND2_X1 U8027 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6897) );
  NAND2_X1 U8028 ( .A1(n9286), .A2(n6550), .ZN(n6905) );
  INV_X1 U8029 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6902) );
  NAND2_X1 U8030 ( .A1(n6533), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6901) );
  NAND2_X1 U8031 ( .A1(n5060), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6900) );
  OAI211_X1 U8032 ( .C1(n6969), .C2(n6902), .A(n6901), .B(n6900), .ZN(n6903)
         );
  INV_X1 U8033 ( .A(n6903), .ZN(n6904) );
  NAND2_X1 U8034 ( .A1(n8780), .A2(n6906), .ZN(n6909) );
  NAND2_X1 U8035 ( .A1(n9309), .A2(n6907), .ZN(n6908) );
  OAI21_X1 U8036 ( .B1(n9309), .B2(n6909), .A(n6908), .ZN(n6910) );
  INV_X1 U8037 ( .A(n6910), .ZN(n6911) );
  XNOR2_X1 U8038 ( .A(n6912), .B(n6911), .ZN(n6957) );
  INV_X1 U8039 ( .A(n6957), .ZN(n6950) );
  INV_X1 U8040 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U8041 ( .A1(n6919), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6920) );
  MUX2_X1 U8042 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6920), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6922) );
  NAND2_X1 U8043 ( .A1(n8462), .A2(n8652), .ZN(n10644) );
  INV_X1 U8044 ( .A(n8462), .ZN(n6928) );
  INV_X1 U8045 ( .A(P2_B_REG_SCAN_IN), .ZN(n6927) );
  NOR2_X1 U8046 ( .A1(n6923), .A2(n10002), .ZN(n6924) );
  MUX2_X1 U8047 ( .A(n10002), .B(n6924), .S(P2_IR_REG_25__SCAN_IN), .Z(n6925)
         );
  INV_X1 U8048 ( .A(n6925), .ZN(n6926) );
  AND2_X1 U8049 ( .A1(n6919), .A2(n6926), .ZN(n6944) );
  NOR2_X1 U8050 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n6931), .ZN(n6929) );
  NAND2_X1 U8051 ( .A1(n6932), .A2(n6929), .ZN(n6930) );
  INV_X1 U8052 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10548) );
  NOR2_X1 U8053 ( .A1(n6944), .A2(n6932), .ZN(n10549) );
  NOR4_X1 U8054 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6936) );
  NOR4_X1 U8055 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6935) );
  NOR4_X1 U8056 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6934) );
  NOR4_X1 U8057 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6933) );
  NAND4_X1 U8058 ( .A1(n6936), .A2(n6935), .A3(n6934), .A4(n6933), .ZN(n6942)
         );
  NOR2_X1 U8059 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6940) );
  NOR4_X1 U8060 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6939) );
  NOR4_X1 U8061 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6938) );
  NOR4_X1 U8062 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6937) );
  NAND4_X1 U8063 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6941)
         );
  OAI21_X1 U8064 ( .B1(n6942), .B2(n6941), .A(n10546), .ZN(n7819) );
  NAND2_X1 U8065 ( .A1(n7820), .A2(n7819), .ZN(n8197) );
  INV_X1 U8066 ( .A(n8197), .ZN(n6943) );
  INV_X1 U8067 ( .A(n6944), .ZN(n8597) );
  XNOR2_X1 U8068 ( .A(n6946), .B(n6945), .ZN(n7283) );
  INV_X1 U8069 ( .A(n7831), .ZN(n10706) );
  OR2_X1 U8070 ( .A1(n10975), .A2(n7285), .ZN(n6948) );
  NOR2_X1 U8071 ( .A1(n10547), .A2(n6948), .ZN(n6949) );
  NAND2_X1 U8072 ( .A1(n6950), .A2(n9135), .ZN(n6982) );
  NAND2_X1 U8073 ( .A1(n9002), .A2(n6511), .ZN(n6953) );
  INV_X1 U8074 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6951) );
  OR2_X1 U8075 ( .A1(n5030), .A2(n6951), .ZN(n6952) );
  NOR2_X1 U8076 ( .A1(n7831), .A2(n6488), .ZN(n10899) );
  INV_X1 U8077 ( .A(n10899), .ZN(n6954) );
  NOR2_X1 U8078 ( .A1(n10547), .A2(n6954), .ZN(n6955) );
  NAND2_X1 U8079 ( .A1(n6974), .A2(n6955), .ZN(n6956) );
  NAND2_X1 U8080 ( .A1(n10948), .A2(n8201), .ZN(n7818) );
  AOI21_X1 U8081 ( .B1(n6957), .B2(n9135), .A(n9098), .ZN(n6958) );
  INV_X1 U8082 ( .A(n6958), .ZN(n6959) );
  NAND2_X1 U8083 ( .A1(n6959), .A2(n9919), .ZN(n6981) );
  INV_X1 U8084 ( .A(n6974), .ZN(n6960) );
  NAND2_X1 U8085 ( .A1(n6960), .A2(n7818), .ZN(n6964) );
  INV_X1 U8086 ( .A(n7283), .ZN(n6961) );
  NOR2_X1 U8087 ( .A1(n7817), .A2(n6961), .ZN(n6962) );
  AND2_X1 U8088 ( .A1(n6962), .A2(n7274), .ZN(n6963) );
  NAND2_X1 U8089 ( .A1(n6964), .A2(n6963), .ZN(n9049) );
  INV_X1 U8090 ( .A(n6965), .ZN(n9277) );
  NAND2_X1 U8091 ( .A1(n9277), .A2(n6550), .ZN(n6972) );
  INV_X1 U8092 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6968) );
  NAND2_X1 U8093 ( .A1(n6533), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U8094 ( .A1(n5060), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6966) );
  OAI211_X1 U8095 ( .C1(n6969), .C2(n6968), .A(n6967), .B(n6966), .ZN(n6970)
         );
  INV_X1 U8096 ( .A(n6970), .ZN(n6971) );
  NAND2_X1 U8097 ( .A1(n6972), .A2(n6971), .ZN(n9292) );
  INV_X1 U8098 ( .A(n9292), .ZN(n8768) );
  NOR2_X1 U8099 ( .A1(n10547), .A2(n8955), .ZN(n6973) );
  NAND2_X1 U8100 ( .A1(n6974), .A2(n6973), .ZN(n9080) );
  OAI22_X1 U8101 ( .A1(n8768), .A2(n9127), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9680), .ZN(n6976) );
  AOI21_X1 U8102 ( .B1(n9286), .B2(n9129), .A(n6976), .ZN(n6977) );
  INV_X1 U8103 ( .A(n6977), .ZN(n6979) );
  NOR2_X1 U8104 ( .A1(n9262), .A2(n9104), .ZN(n6978) );
  OAI211_X1 U8105 ( .C1(n6982), .C2(n9919), .A(n6981), .B(n6980), .ZN(P2_U3222) );
  AND2_X1 U8106 ( .A1(n7271), .A2(n10344), .ZN(n7117) );
  INV_X1 U8107 ( .A(n7110), .ZN(n7107) );
  INV_X1 U8108 ( .A(n6983), .ZN(n6984) );
  INV_X1 U8109 ( .A(SI_28_), .ZN(n9419) );
  NAND2_X1 U8110 ( .A1(n6984), .A2(n9419), .ZN(n6985) );
  MUX2_X1 U8111 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n6995), .Z(n6988) );
  INV_X1 U8112 ( .A(n6988), .ZN(n6989) );
  MUX2_X1 U8113 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6995), .Z(n6992) );
  NAND2_X1 U8114 ( .A1(n6992), .A2(SI_30_), .ZN(n6994) );
  OAI21_X1 U8115 ( .B1(n6992), .B2(SI_30_), .A(n6994), .ZN(n6993) );
  INV_X1 U8116 ( .A(n6993), .ZN(n7001) );
  MUX2_X1 U8117 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6995), .Z(n6996) );
  XNOR2_X1 U8118 ( .A(n6996), .B(SI_31_), .ZN(n6997) );
  INV_X1 U8119 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6999) );
  NOR2_X1 U8120 ( .A1(n7015), .A2(n6999), .ZN(n7000) );
  NAND2_X1 U8121 ( .A1(n8752), .A2(n7005), .ZN(n7007) );
  INV_X1 U8122 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8708) );
  OR2_X1 U8123 ( .A1(n7015), .A2(n8708), .ZN(n7006) );
  NAND2_X1 U8124 ( .A1(n7101), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7010) );
  NAND2_X1 U8125 ( .A1(n6303), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7009) );
  NAND2_X1 U8126 ( .A1(n6302), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7008) );
  NAND3_X1 U8127 ( .A1(n7010), .A2(n7009), .A3(n7008), .ZN(n10276) );
  INV_X1 U8128 ( .A(n10276), .ZN(n7118) );
  OR2_X1 U8129 ( .A1(n10449), .A2(n7118), .ZN(n7253) );
  INV_X1 U8130 ( .A(n7011), .ZN(n7012) );
  INV_X1 U8131 ( .A(SI_29_), .ZN(n9413) );
  NAND2_X1 U8132 ( .A1(n7012), .A2(n9413), .ZN(n7013) );
  INV_X1 U8133 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8695) );
  OR2_X1 U8134 ( .A1(n7015), .A2(n8695), .ZN(n7016) );
  NAND2_X1 U8135 ( .A1(n10455), .A2(n10297), .ZN(n10270) );
  NAND2_X1 U8136 ( .A1(n10461), .A2(n10305), .ZN(n7143) );
  NAND2_X1 U8137 ( .A1(n8986), .A2(n8984), .ZN(n7213) );
  NAND2_X1 U8138 ( .A1(n10375), .A2(n10390), .ZN(n8982) );
  OR2_X1 U8139 ( .A1(n7213), .A2(n8982), .ZN(n7018) );
  AND2_X1 U8140 ( .A1(n10485), .A2(n10161), .ZN(n8983) );
  INV_X1 U8141 ( .A(n8983), .ZN(n7184) );
  MUX2_X1 U8142 ( .A(n7018), .B(n7184), .S(n7110), .Z(n7086) );
  NAND2_X1 U8143 ( .A1(n7213), .A2(n7107), .ZN(n7083) );
  NAND2_X1 U8144 ( .A1(n10481), .A2(n10371), .ZN(n7188) );
  NAND2_X1 U8145 ( .A1(n8984), .A2(n7188), .ZN(n10358) );
  INV_X1 U8146 ( .A(n10358), .ZN(n7080) );
  NAND2_X1 U8147 ( .A1(n7184), .A2(n8982), .ZN(n10369) );
  INV_X1 U8148 ( .A(n10369), .ZN(n7134) );
  NAND2_X1 U8149 ( .A1(n8980), .A2(n8978), .ZN(n7181) );
  NAND2_X1 U8150 ( .A1(n10493), .A2(n10402), .ZN(n7074) );
  NAND2_X1 U8151 ( .A1(n7181), .A2(n7074), .ZN(n7020) );
  NAND2_X1 U8152 ( .A1(n10496), .A2(n10431), .ZN(n7075) );
  NAND2_X1 U8153 ( .A1(n7074), .A2(n7075), .ZN(n7019) );
  NAND2_X1 U8154 ( .A1(n7019), .A2(n8980), .ZN(n7144) );
  MUX2_X1 U8155 ( .A(n7020), .B(n7144), .S(n7110), .Z(n7078) );
  XNOR2_X1 U8156 ( .A(n5704), .B(n7216), .ZN(n7120) );
  NAND2_X1 U8157 ( .A1(n7120), .A2(n7714), .ZN(n7023) );
  INV_X1 U8158 ( .A(n5704), .ZN(n7851) );
  NAND2_X1 U8159 ( .A1(n7851), .A2(n7216), .ZN(n7022) );
  NAND2_X1 U8160 ( .A1(n7023), .A2(n7022), .ZN(n7848) );
  NAND2_X1 U8161 ( .A1(n5727), .A2(n10724), .ZN(n7221) );
  INV_X1 U8162 ( .A(n7220), .ZN(n7025) );
  INV_X1 U8163 ( .A(n10175), .ZN(n7852) );
  NAND2_X1 U8164 ( .A1(n7852), .A2(n10738), .ZN(n7224) );
  NAND2_X1 U8165 ( .A1(n7738), .A2(n7224), .ZN(n7026) );
  INV_X1 U8166 ( .A(n10738), .ZN(n7759) );
  NAND2_X1 U8167 ( .A1(n10175), .A2(n7759), .ZN(n7222) );
  AND2_X1 U8168 ( .A1(n10174), .A2(n10758), .ZN(n7028) );
  NAND2_X1 U8169 ( .A1(n7772), .A2(n7785), .ZN(n7027) );
  XNOR2_X1 U8170 ( .A(n7901), .B(n7107), .ZN(n7032) );
  INV_X1 U8171 ( .A(n10173), .ZN(n7924) );
  NAND2_X1 U8172 ( .A1(n7924), .A2(n7800), .ZN(n7227) );
  INV_X1 U8173 ( .A(n7800), .ZN(n10794) );
  NAND2_X1 U8174 ( .A1(n10173), .A2(n10794), .ZN(n7230) );
  NAND2_X1 U8175 ( .A1(n10850), .A2(n7930), .ZN(n7233) );
  NAND2_X1 U8176 ( .A1(n7734), .A2(n10825), .ZN(n7231) );
  INV_X1 U8177 ( .A(n10172), .ZN(n8125) );
  NAND2_X1 U8178 ( .A1(n8125), .A2(n7910), .ZN(n7904) );
  NAND2_X1 U8179 ( .A1(n10863), .A2(n10172), .ZN(n7234) );
  AND2_X2 U8180 ( .A1(n7904), .A2(n7234), .ZN(n10848) );
  NAND3_X1 U8181 ( .A1(n7924), .A2(n7107), .A3(n7800), .ZN(n7030) );
  NAND3_X1 U8182 ( .A1(n10173), .A2(n10794), .A3(n7110), .ZN(n7029) );
  NAND4_X1 U8183 ( .A1(n7806), .A2(n10848), .A3(n7030), .A4(n7029), .ZN(n7031)
         );
  AOI21_X1 U8184 ( .B1(n7032), .B2(n7768), .A(n7031), .ZN(n7038) );
  NAND2_X1 U8185 ( .A1(n7233), .A2(n7904), .ZN(n7033) );
  NAND2_X1 U8186 ( .A1(n7033), .A2(n7234), .ZN(n7035) );
  NAND2_X1 U8187 ( .A1(n7234), .A2(n7231), .ZN(n7190) );
  NAND2_X1 U8188 ( .A1(n7190), .A2(n7904), .ZN(n7034) );
  MUX2_X1 U8189 ( .A(n7035), .B(n7034), .S(n7107), .Z(n7036) );
  INV_X1 U8190 ( .A(n7036), .ZN(n7037) );
  NAND2_X1 U8191 ( .A1(n10882), .A2(n10171), .ZN(n7905) );
  INV_X1 U8192 ( .A(n10882), .ZN(n8133) );
  NAND2_X1 U8193 ( .A1(n8133), .A2(n10852), .ZN(n7906) );
  NAND2_X1 U8194 ( .A1(n7905), .A2(n7906), .ZN(n7932) );
  INV_X1 U8195 ( .A(n7932), .ZN(n7935) );
  OAI21_X1 U8196 ( .B1(n7038), .B2(n7037), .A(n7935), .ZN(n7044) );
  XNOR2_X1 U8197 ( .A(n8076), .B(n10170), .ZN(n8079) );
  MUX2_X1 U8198 ( .A(n7906), .B(n7905), .S(n7107), .Z(n7039) );
  AND2_X1 U8199 ( .A1(n8079), .A2(n7039), .ZN(n7043) );
  OR2_X1 U8200 ( .A1(n8475), .A2(n8226), .ZN(n7154) );
  INV_X1 U8201 ( .A(n10170), .ZN(n8467) );
  OR2_X1 U8202 ( .A1(n8076), .A2(n8467), .ZN(n7151) );
  NAND2_X1 U8203 ( .A1(n7154), .A2(n7151), .ZN(n7041) );
  NAND2_X1 U8204 ( .A1(n8076), .A2(n8467), .ZN(n8081) );
  INV_X1 U8205 ( .A(n8081), .ZN(n7040) );
  MUX2_X1 U8206 ( .A(n7041), .B(n7040), .S(n7107), .Z(n7042) );
  AOI21_X1 U8207 ( .B1(n7044), .B2(n7043), .A(n7042), .ZN(n7045) );
  MUX2_X1 U8208 ( .A(n7110), .B(n7045), .S(n8085), .Z(n7047) );
  OAI21_X1 U8209 ( .B1(n7110), .B2(n7154), .A(n8084), .ZN(n7046) );
  OR2_X1 U8210 ( .A1(n7047), .A2(n7046), .ZN(n7050) );
  INV_X1 U8211 ( .A(n11005), .ZN(n8560) );
  OR2_X1 U8212 ( .A1(n8385), .A2(n8560), .ZN(n7159) );
  NAND2_X1 U8213 ( .A1(n8385), .A2(n8560), .ZN(n8389) );
  INV_X1 U8214 ( .A(n10168), .ZN(n8309) );
  NAND2_X1 U8215 ( .A1(n8094), .A2(n8309), .ZN(n8174) );
  OR2_X1 U8216 ( .A1(n8094), .A2(n8309), .ZN(n7158) );
  MUX2_X1 U8217 ( .A(n8174), .B(n7158), .S(n7110), .Z(n7048) );
  AND2_X1 U8218 ( .A1(n8176), .A2(n7048), .ZN(n7049) );
  NAND2_X1 U8219 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  INV_X1 U8220 ( .A(n10167), .ZN(n8662) );
  NAND2_X1 U8221 ( .A1(n8552), .A2(n8662), .ZN(n8391) );
  INV_X1 U8222 ( .A(n8391), .ZN(n7057) );
  AOI21_X1 U8223 ( .B1(n7051), .B2(n7159), .A(n7057), .ZN(n7053) );
  OR2_X1 U8224 ( .A1(n8552), .A2(n8662), .ZN(n7162) );
  INV_X1 U8225 ( .A(n7162), .ZN(n7055) );
  AOI21_X1 U8226 ( .B1(n7051), .B2(n8389), .A(n7055), .ZN(n7052) );
  MUX2_X1 U8227 ( .A(n7053), .B(n7052), .S(n7110), .Z(n7054) );
  INV_X1 U8228 ( .A(n5054), .ZN(n8392) );
  NAND2_X1 U8229 ( .A1(n7054), .A2(n8392), .ZN(n7063) );
  INV_X1 U8230 ( .A(n8659), .ZN(n10067) );
  NAND2_X1 U8231 ( .A1(n10135), .A2(n10067), .ZN(n7149) );
  INV_X1 U8232 ( .A(n11004), .ZN(n10150) );
  NAND2_X1 U8233 ( .A1(n8664), .A2(n10150), .ZN(n7148) );
  NAND2_X1 U8234 ( .A1(n7148), .A2(n7055), .ZN(n7056) );
  OR2_X1 U8235 ( .A1(n8664), .A2(n10150), .ZN(n8511) );
  NAND2_X1 U8236 ( .A1(n7056), .A2(n8511), .ZN(n7060) );
  NAND2_X1 U8237 ( .A1(n8511), .A2(n7057), .ZN(n7058) );
  NAND2_X1 U8238 ( .A1(n7058), .A2(n7148), .ZN(n7059) );
  MUX2_X1 U8239 ( .A(n7060), .B(n7059), .S(n7110), .Z(n7061) );
  INV_X1 U8240 ( .A(n7061), .ZN(n7062) );
  NAND3_X1 U8241 ( .A1(n7063), .A2(n8528), .A3(n7062), .ZN(n7065) );
  NAND2_X1 U8242 ( .A1(n11084), .A2(n10146), .ZN(n7147) );
  NAND2_X1 U8243 ( .A1(n10069), .A2(n10076), .ZN(n8603) );
  NAND2_X1 U8244 ( .A1(n7147), .A2(n8603), .ZN(n8584) );
  INV_X1 U8245 ( .A(n8584), .ZN(n7128) );
  MUX2_X1 U8246 ( .A(n7149), .B(n8576), .S(n7110), .Z(n7064) );
  NAND3_X1 U8247 ( .A1(n7065), .A2(n7128), .A3(n7064), .ZN(n7067) );
  MUX2_X1 U8248 ( .A(n7147), .B(n8603), .S(n7110), .Z(n7066) );
  NAND2_X1 U8249 ( .A1(n10514), .A2(n8626), .ZN(n7145) );
  NAND2_X1 U8250 ( .A1(n8617), .A2(n7145), .ZN(n8607) );
  AOI21_X1 U8251 ( .B1(n7067), .B2(n7066), .A(n8607), .ZN(n7071) );
  NAND2_X1 U8252 ( .A1(n10507), .A2(n10430), .ZN(n7175) );
  MUX2_X1 U8253 ( .A(n8617), .B(n7145), .S(n7110), .Z(n7068) );
  NAND2_X1 U8254 ( .A1(n8973), .A2(n7068), .ZN(n7070) );
  OR2_X1 U8255 ( .A1(n10503), .A2(n10401), .ZN(n7178) );
  NAND2_X1 U8256 ( .A1(n10503), .A2(n10401), .ZN(n10398) );
  NAND2_X1 U8257 ( .A1(n7178), .A2(n10398), .ZN(n10427) );
  INV_X1 U8258 ( .A(n10427), .ZN(n7131) );
  MUX2_X1 U8259 ( .A(n8975), .B(n7175), .S(n7107), .Z(n7069) );
  OAI211_X1 U8260 ( .C1(n7071), .C2(n7070), .A(n7131), .B(n7069), .ZN(n7073)
         );
  MUX2_X1 U8261 ( .A(n7178), .B(n10398), .S(n7110), .Z(n7072) );
  NAND2_X1 U8262 ( .A1(n7073), .A2(n7072), .ZN(n7076) );
  NAND2_X1 U8263 ( .A1(n8978), .A2(n7075), .ZN(n10403) );
  INV_X1 U8264 ( .A(n10403), .ZN(n10399) );
  NAND3_X1 U8265 ( .A1(n7076), .A2(n10388), .A3(n10399), .ZN(n7077) );
  NAND3_X1 U8266 ( .A1(n7134), .A2(n7078), .A3(n7077), .ZN(n7079) );
  NAND2_X1 U8267 ( .A1(n7080), .A2(n7079), .ZN(n7082) );
  NAND2_X1 U8268 ( .A1(n10476), .A2(n10359), .ZN(n7193) );
  INV_X1 U8269 ( .A(n7193), .ZN(n7081) );
  AOI21_X1 U8270 ( .B1(n7083), .B2(n7082), .A(n7081), .ZN(n7085) );
  AOI21_X1 U8271 ( .B1(n7193), .B2(n7188), .A(n7107), .ZN(n7084) );
  AOI21_X1 U8272 ( .B1(n7086), .B2(n7085), .A(n7084), .ZN(n7090) );
  OR2_X1 U8273 ( .A1(n10471), .A2(n10340), .ZN(n8988) );
  NAND2_X1 U8274 ( .A1(n10471), .A2(n10340), .ZN(n7194) );
  NAND2_X1 U8275 ( .A1(n8988), .A2(n7194), .ZN(n10321) );
  NOR2_X1 U8276 ( .A1(n8986), .A2(n7107), .ZN(n7087) );
  OR2_X1 U8277 ( .A1(n10321), .A2(n7087), .ZN(n7089) );
  NAND2_X1 U8278 ( .A1(n10314), .A2(n10052), .ZN(n7195) );
  NAND2_X1 U8279 ( .A1(n10465), .A2(n10323), .ZN(n8989) );
  MUX2_X1 U8280 ( .A(n8988), .B(n7194), .S(n7110), .Z(n7088) );
  OAI211_X1 U8281 ( .C1(n7090), .C2(n7089), .A(n10306), .B(n7088), .ZN(n7092)
         );
  MUX2_X1 U8282 ( .A(n8989), .B(n7195), .S(n7110), .Z(n7091) );
  NAND3_X1 U8283 ( .A1(n8968), .A2(n7092), .A3(n7091), .ZN(n7094) );
  MUX2_X1 U8284 ( .A(n7196), .B(n7143), .S(n7110), .Z(n7093) );
  AND3_X1 U8285 ( .A1(n8992), .A2(n7094), .A3(n7093), .ZN(n7097) );
  INV_X1 U8286 ( .A(n7097), .ZN(n7095) );
  NAND3_X1 U8287 ( .A1(n7250), .A2(n10270), .A3(n7095), .ZN(n7096) );
  NAND2_X1 U8288 ( .A1(n7096), .A2(n7212), .ZN(n7099) );
  NAND2_X1 U8289 ( .A1(n7212), .A2(n7211), .ZN(n7202) );
  OAI21_X1 U8290 ( .B1(n7202), .B2(n7097), .A(n7250), .ZN(n7098) );
  MUX2_X1 U8291 ( .A(n7099), .B(n7098), .S(n7110), .Z(n7100) );
  OAI21_X1 U8292 ( .B1(n10445), .B2(n7253), .A(n7100), .ZN(n7106) );
  NAND2_X1 U8293 ( .A1(n7101), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7104) );
  NAND2_X1 U8294 ( .A1(n6303), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7103) );
  NAND2_X1 U8295 ( .A1(n6302), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7102) );
  NAND3_X1 U8296 ( .A1(n7104), .A2(n7103), .A3(n7102), .ZN(n10261) );
  NAND2_X1 U8297 ( .A1(n10261), .A2(n10276), .ZN(n7105) );
  NAND2_X1 U8298 ( .A1(n10449), .A2(n7105), .ZN(n7200) );
  MUX2_X2 U8299 ( .A(n7107), .B(n7106), .S(n7200), .Z(n7112) );
  INV_X1 U8300 ( .A(n10445), .ZN(n7114) );
  INV_X1 U8301 ( .A(n10261), .ZN(n7113) );
  NAND2_X1 U8302 ( .A1(n7114), .A2(n7113), .ZN(n7255) );
  INV_X1 U8303 ( .A(n7255), .ZN(n7111) );
  INV_X1 U8304 ( .A(n7253), .ZN(n7108) );
  NAND2_X1 U8305 ( .A1(n7108), .A2(n10261), .ZN(n7109) );
  AND2_X1 U8306 ( .A1(n7109), .A2(n7255), .ZN(n7142) );
  OAI21_X1 U8307 ( .B1(n7716), .B2(n8102), .A(n7116), .ZN(n7115) );
  OAI211_X1 U8308 ( .C1(n7117), .C2(n7116), .A(n7115), .B(n7256), .ZN(n7210)
         );
  INV_X1 U8309 ( .A(n10272), .ZN(n7139) );
  NAND2_X1 U8310 ( .A1(n10449), .A2(n7118), .ZN(n7249) );
  NAND2_X1 U8311 ( .A1(n8986), .A2(n7193), .ZN(n10338) );
  AND2_X1 U8312 ( .A1(n7119), .A2(n7021), .ZN(n7215) );
  NOR2_X1 U8313 ( .A1(n7714), .A2(n7215), .ZN(n7583) );
  NAND2_X1 U8314 ( .A1(n7224), .A2(n7222), .ZN(n7757) );
  INV_X1 U8315 ( .A(n7757), .ZN(n7748) );
  NOR2_X1 U8316 ( .A1(n7121), .A2(n7764), .ZN(n7122) );
  XNOR2_X1 U8317 ( .A(n10174), .B(n10758), .ZN(n7788) );
  INV_X1 U8318 ( .A(n7788), .ZN(n7780) );
  NAND4_X1 U8319 ( .A1(n7122), .A2(n7806), .A3(n10848), .A4(n7780), .ZN(n7123)
         );
  NOR2_X1 U8320 ( .A1(n7123), .A2(n7932), .ZN(n7124) );
  AND4_X1 U8321 ( .A1(n8176), .A2(n8160), .A3(n7124), .A4(n8079), .ZN(n7125)
         );
  NAND3_X1 U8322 ( .A1(n11007), .A2(n7125), .A3(n8084), .ZN(n7126) );
  NOR2_X1 U8323 ( .A1(n5054), .A2(n7126), .ZN(n7127) );
  NAND3_X1 U8324 ( .A1(n7128), .A2(n8528), .A3(n7127), .ZN(n7129) );
  NOR2_X1 U8325 ( .A1(n8607), .A2(n7129), .ZN(n7130) );
  NAND3_X1 U8326 ( .A1(n7131), .A2(n8973), .A3(n7130), .ZN(n7132) );
  NOR2_X1 U8327 ( .A1(n7132), .A2(n10403), .ZN(n7133) );
  NAND3_X1 U8328 ( .A1(n7134), .A2(n10388), .A3(n7133), .ZN(n7135) );
  NOR2_X1 U8329 ( .A1(n10358), .A2(n7135), .ZN(n7136) );
  NAND4_X1 U8330 ( .A1(n10306), .A2(n5304), .A3(n5190), .A4(n7136), .ZN(n7137)
         );
  NOR2_X1 U8331 ( .A1(n10296), .A2(n7137), .ZN(n7138) );
  AND4_X1 U8332 ( .A1(n7139), .A2(n7249), .A3(n8992), .A4(n7138), .ZN(n7140)
         );
  NAND4_X1 U8333 ( .A1(n7256), .A2(n7140), .A3(n7255), .A4(n7253), .ZN(n7141)
         );
  NAND2_X1 U8334 ( .A1(n7141), .A2(n8102), .ZN(n7208) );
  INV_X1 U8335 ( .A(n7142), .ZN(n7205) );
  INV_X1 U8336 ( .A(n7196), .ZN(n8990) );
  OAI211_X1 U8337 ( .C1(n8990), .C2(n8989), .A(n10270), .B(n7143), .ZN(n7247)
         );
  NAND2_X1 U8338 ( .A1(n8982), .A2(n7144), .ZN(n7186) );
  AND2_X1 U8339 ( .A1(n7145), .A2(n8603), .ZN(n7146) );
  NAND2_X1 U8340 ( .A1(n7175), .A2(n7146), .ZN(n7171) );
  AND2_X1 U8341 ( .A1(n7147), .A2(n8576), .ZN(n8601) );
  NAND2_X1 U8342 ( .A1(n7149), .A2(n7148), .ZN(n7170) );
  INV_X1 U8343 ( .A(n7905), .ZN(n7150) );
  NAND2_X1 U8344 ( .A1(n8081), .A2(n7150), .ZN(n7152) );
  NAND2_X1 U8345 ( .A1(n7152), .A2(n7151), .ZN(n7153) );
  NAND2_X1 U8346 ( .A1(n7153), .A2(n8085), .ZN(n7155) );
  NAND2_X1 U8347 ( .A1(n7155), .A2(n7154), .ZN(n7156) );
  NAND2_X1 U8348 ( .A1(n8174), .A2(n7156), .ZN(n7157) );
  NAND3_X1 U8349 ( .A1(n7159), .A2(n7158), .A3(n7157), .ZN(n7160) );
  NAND2_X1 U8350 ( .A1(n7160), .A2(n8389), .ZN(n7161) );
  NAND2_X1 U8351 ( .A1(n7162), .A2(n7161), .ZN(n7163) );
  NAND2_X1 U8352 ( .A1(n7163), .A2(n8391), .ZN(n7164) );
  AND2_X1 U8353 ( .A1(n8511), .A2(n7164), .ZN(n7165) );
  OR2_X1 U8354 ( .A1(n7170), .A2(n7165), .ZN(n7166) );
  AND2_X1 U8355 ( .A1(n8601), .A2(n7166), .ZN(n7167) );
  OR2_X1 U8356 ( .A1(n7171), .A2(n7167), .ZN(n7236) );
  AND4_X1 U8357 ( .A1(n8085), .A2(n8081), .A3(n7906), .A4(n7904), .ZN(n7168)
         );
  NAND4_X1 U8358 ( .A1(n8391), .A2(n7168), .A3(n8389), .A4(n8174), .ZN(n7169)
         );
  OR3_X1 U8359 ( .A1(n7171), .A2(n7170), .A3(n7169), .ZN(n7172) );
  NAND2_X1 U8360 ( .A1(n7236), .A2(n7172), .ZN(n7173) );
  NAND2_X1 U8361 ( .A1(n7173), .A2(n10398), .ZN(n7185) );
  INV_X1 U8362 ( .A(n8617), .ZN(n7174) );
  NAND2_X1 U8363 ( .A1(n7175), .A2(n7174), .ZN(n7176) );
  NAND2_X1 U8364 ( .A1(n7176), .A2(n8975), .ZN(n7177) );
  NAND2_X1 U8365 ( .A1(n10398), .A2(n7177), .ZN(n7179) );
  NAND2_X1 U8366 ( .A1(n7179), .A2(n7178), .ZN(n7180) );
  NOR2_X1 U8367 ( .A1(n7181), .A2(n7180), .ZN(n7182) );
  OR2_X1 U8368 ( .A1(n7186), .A2(n7182), .ZN(n7183) );
  AND2_X1 U8369 ( .A1(n7184), .A2(n7183), .ZN(n7214) );
  OAI21_X1 U8370 ( .B1(n7186), .B2(n7185), .A(n7214), .ZN(n7187) );
  AND2_X1 U8371 ( .A1(n7188), .A2(n7187), .ZN(n7237) );
  INV_X1 U8372 ( .A(n7227), .ZN(n7189) );
  AOI21_X1 U8373 ( .B1(n7901), .B2(n7768), .A(n7189), .ZN(n7805) );
  AOI21_X1 U8374 ( .B1(n7805), .B2(n7233), .A(n7190), .ZN(n7191) );
  NAND3_X1 U8375 ( .A1(n7214), .A2(n7191), .A3(n7236), .ZN(n7192) );
  AOI21_X1 U8376 ( .B1(n7237), .B2(n7192), .A(n7213), .ZN(n7197) );
  NAND2_X1 U8377 ( .A1(n7194), .A2(n7193), .ZN(n7240) );
  AND2_X1 U8378 ( .A1(n7195), .A2(n8988), .ZN(n7243) );
  OAI211_X1 U8379 ( .C1(n7197), .C2(n7240), .A(n7196), .B(n7243), .ZN(n7198)
         );
  INV_X1 U8380 ( .A(n7198), .ZN(n7199) );
  NOR2_X1 U8381 ( .A1(n7247), .A2(n7199), .ZN(n7201) );
  OAI211_X1 U8382 ( .C1(n7202), .C2(n7201), .A(n7200), .B(n7250), .ZN(n7203)
         );
  INV_X1 U8383 ( .A(n7203), .ZN(n7204) );
  OAI211_X1 U8384 ( .C1(n7205), .C2(n7204), .A(n7718), .B(n7256), .ZN(n7206)
         );
  NAND2_X1 U8385 ( .A1(n7206), .A2(n7208), .ZN(n7207) );
  MUX2_X1 U8386 ( .A(n7208), .B(n7207), .S(n10392), .Z(n7209) );
  NAND2_X1 U8387 ( .A1(n7210), .A2(n7209), .ZN(n7263) );
  AND2_X1 U8388 ( .A1(n7212), .A2(n7211), .ZN(n7248) );
  INV_X1 U8389 ( .A(n7213), .ZN(n7242) );
  INV_X1 U8390 ( .A(n7214), .ZN(n7239) );
  INV_X1 U8391 ( .A(n7215), .ZN(n7218) );
  INV_X1 U8392 ( .A(n7216), .ZN(n10716) );
  NAND2_X1 U8393 ( .A1(n5704), .A2(n10716), .ZN(n7217) );
  NAND3_X1 U8394 ( .A1(n7218), .A2(n7718), .A3(n7217), .ZN(n7219) );
  NAND2_X1 U8395 ( .A1(n7220), .A2(n7219), .ZN(n7223) );
  OAI211_X1 U8396 ( .C1(n7848), .C2(n7223), .A(n7222), .B(n7221), .ZN(n7225)
         );
  NAND2_X1 U8397 ( .A1(n7225), .A2(n7224), .ZN(n7226) );
  AOI21_X1 U8398 ( .B1(n7226), .B2(n7785), .A(n7772), .ZN(n7229) );
  NOR2_X1 U8399 ( .A1(n7226), .A2(n7785), .ZN(n7228) );
  OAI21_X1 U8400 ( .B1(n7229), .B2(n7228), .A(n5123), .ZN(n7235) );
  NAND2_X1 U8401 ( .A1(n7231), .A2(n7230), .ZN(n7232) );
  NAND2_X1 U8402 ( .A1(n7233), .A2(n7232), .ZN(n10844) );
  NAND4_X1 U8403 ( .A1(n7236), .A2(n7235), .A3(n7234), .A4(n10844), .ZN(n7238)
         );
  OAI21_X1 U8404 ( .B1(n7239), .B2(n7238), .A(n7237), .ZN(n7241) );
  AOI21_X1 U8405 ( .B1(n7242), .B2(n7241), .A(n7240), .ZN(n7245) );
  INV_X1 U8406 ( .A(n7243), .ZN(n7244) );
  NOR2_X1 U8407 ( .A1(n7245), .A2(n7244), .ZN(n7246) );
  NAND3_X1 U8408 ( .A1(n7248), .A2(n8968), .A3(n7246), .ZN(n7252) );
  NAND2_X1 U8409 ( .A1(n7248), .A2(n7247), .ZN(n7251) );
  NAND4_X1 U8410 ( .A1(n7252), .A2(n7251), .A3(n7250), .A4(n7249), .ZN(n7254)
         );
  NAND3_X1 U8411 ( .A1(n7255), .A2(n7254), .A3(n7253), .ZN(n7257) );
  NAND2_X1 U8412 ( .A1(n7257), .A2(n7256), .ZN(n7258) );
  XNOR2_X1 U8413 ( .A(n7258), .B(n10392), .ZN(n7260) );
  OR2_X1 U8414 ( .A1(n7495), .A2(P1_U3084), .ZN(n8295) );
  INV_X1 U8415 ( .A(n8295), .ZN(n7259) );
  OR3_X1 U8416 ( .A1(n10849), .A2(n7580), .A3(n10259), .ZN(n7265) );
  NOR2_X1 U8417 ( .A1(n7265), .A2(n7577), .ZN(n7267) );
  OAI21_X1 U8418 ( .B1(n7716), .B2(n8295), .A(P1_B_REG_SCAN_IN), .ZN(n7266) );
  OR2_X1 U8419 ( .A1(n7267), .A2(n7266), .ZN(n7268) );
  NAND2_X1 U8420 ( .A1(n7269), .A2(n7268), .ZN(P1_U3240) );
  INV_X1 U8421 ( .A(n7426), .ZN(n7270) );
  INV_X1 U8422 ( .A(n7271), .ZN(n7581) );
  NAND2_X1 U8423 ( .A1(n7497), .A2(n7581), .ZN(n7272) );
  NAND2_X1 U8424 ( .A1(n7272), .A2(n7495), .ZN(n7492) );
  NAND2_X1 U8425 ( .A1(n7492), .A2(n7470), .ZN(n7273) );
  NAND2_X1 U8426 ( .A1(n7273), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8427 ( .A(n7274), .ZN(n7282) );
  INV_X1 U8428 ( .A(n7433), .ZN(n7300) );
  INV_X1 U8429 ( .A(n7430), .ZN(n10668) );
  INV_X1 U8430 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U8431 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10662) );
  NOR2_X1 U8432 ( .A1(n10661), .A2(n10662), .ZN(n10660) );
  AOI21_X1 U8433 ( .B1(n10668), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10660), .ZN(
        n10676) );
  NAND2_X1 U8434 ( .A1(n10683), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7276) );
  OAI21_X1 U8435 ( .B1(n10683), .B2(P2_REG1_REG_2__SCAN_IN), .A(n7276), .ZN(
        n10675) );
  NAND2_X1 U8436 ( .A1(n7293), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7277) );
  OAI21_X1 U8437 ( .B1(n7293), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7277), .ZN(
        n7343) );
  NAND2_X1 U8438 ( .A1(n7295), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7278) );
  OAI21_X1 U8439 ( .B1(n7295), .B2(P2_REG1_REG_4__SCAN_IN), .A(n7278), .ZN(
        n7354) );
  NOR2_X1 U8440 ( .A1(n7355), .A2(n7354), .ZN(n7353) );
  NAND2_X1 U8441 ( .A1(n7297), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7279) );
  OAI21_X1 U8442 ( .B1(n7297), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7279), .ZN(
        n7331) );
  INV_X1 U8443 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7280) );
  MUX2_X1 U8444 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7280), .S(n7433), .Z(n7379)
         );
  AOI21_X1 U8445 ( .B1(n7300), .B2(P2_REG1_REG_6__SCAN_IN), .A(n7378), .ZN(
        n7289) );
  NAND2_X1 U8446 ( .A1(n7320), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7281) );
  OAI21_X1 U8447 ( .B1(n7320), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7281), .ZN(
        n7288) );
  NOR2_X1 U8448 ( .A1(n7289), .A2(n7288), .ZN(n7315) );
  NOR2_X1 U8449 ( .A1(n6975), .A2(P2_U3152), .ZN(n10009) );
  NAND2_X1 U8450 ( .A1(n7282), .A2(n10009), .ZN(n7284) );
  OR2_X1 U8451 ( .A1(n7283), .A2(P2_U3152), .ZN(n8958) );
  OAI211_X1 U8452 ( .C1(n10547), .C2(n7285), .A(n7284), .B(n8958), .ZN(n7286)
         );
  NAND2_X1 U8453 ( .A1(n7286), .A2(n7306), .ZN(n7290) );
  INV_X1 U8454 ( .A(n7287), .ZN(n9239) );
  AOI211_X1 U8455 ( .C1(n7289), .C2(n7288), .A(n7315), .B(n10673), .ZN(n7314)
         );
  NAND2_X1 U8456 ( .A1(n7290), .A2(n9160), .ZN(n7303) );
  NOR2_X1 U8457 ( .A1(n10653), .A2(n7436), .ZN(n7313) );
  INV_X1 U8458 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8286) );
  MUX2_X1 U8459 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n8286), .S(n7430), .Z(n10664)
         );
  NAND2_X1 U8460 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10665) );
  NOR2_X1 U8461 ( .A1(n10664), .A2(n10665), .ZN(n10663) );
  AOI21_X1 U8462 ( .B1(n10668), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10663), .ZN(
        n10680) );
  NAND2_X1 U8463 ( .A1(n10683), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7291) );
  OAI21_X1 U8464 ( .B1(n10683), .B2(P2_REG2_REG_2__SCAN_IN), .A(n7291), .ZN(
        n10679) );
  NOR2_X1 U8465 ( .A1(n10680), .A2(n10679), .ZN(n10678) );
  NAND2_X1 U8466 ( .A1(n7293), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7292) );
  OAI21_X1 U8467 ( .B1(n7293), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7292), .ZN(
        n7346) );
  NOR2_X1 U8468 ( .A1(n7347), .A2(n7346), .ZN(n7345) );
  AOI21_X1 U8469 ( .B1(n7293), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7345), .ZN(
        n7358) );
  NAND2_X1 U8470 ( .A1(n7295), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7294) );
  OAI21_X1 U8471 ( .B1(n7295), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7294), .ZN(
        n7357) );
  NOR2_X1 U8472 ( .A1(n7358), .A2(n7357), .ZN(n7356) );
  AOI21_X1 U8473 ( .B1(n7295), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7356), .ZN(
        n7335) );
  NAND2_X1 U8474 ( .A1(n7297), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7296) );
  OAI21_X1 U8475 ( .B1(n7297), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7296), .ZN(
        n7334) );
  NOR2_X1 U8476 ( .A1(n7335), .A2(n7334), .ZN(n7333) );
  AOI21_X1 U8477 ( .B1(n7297), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7333), .ZN(
        n7383) );
  INV_X1 U8478 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7298) );
  MUX2_X1 U8479 ( .A(n7298), .B(P2_REG2_REG_6__SCAN_IN), .S(n7433), .Z(n7299)
         );
  INV_X1 U8480 ( .A(n7299), .ZN(n7382) );
  NOR2_X1 U8481 ( .A1(n7383), .A2(n7382), .ZN(n7381) );
  AOI21_X1 U8482 ( .B1(n7300), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7381), .ZN(
        n7305) );
  NAND2_X1 U8483 ( .A1(n7320), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7301) );
  OAI21_X1 U8484 ( .B1(n7320), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7301), .ZN(
        n7304) );
  NOR2_X1 U8485 ( .A1(n7305), .A2(n7304), .ZN(n7319) );
  NOR2_X1 U8486 ( .A1(n6975), .A2(n7287), .ZN(n7302) );
  AOI211_X1 U8487 ( .C1(n7305), .C2(n7304), .A(n7319), .B(n10677), .ZN(n7312)
         );
  OAI21_X1 U8488 ( .B1(n10547), .B2(n7824), .A(n7306), .ZN(n7308) );
  NAND2_X1 U8489 ( .A1(n10547), .A2(n8958), .ZN(n7307) );
  INV_X1 U8490 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7310) );
  NAND2_X1 U8491 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n7309) );
  OAI21_X1 U8492 ( .B1(n9217), .B2(n7310), .A(n7309), .ZN(n7311) );
  OR4_X1 U8493 ( .A1(n7314), .A2(n7313), .A3(n7312), .A4(n7311), .ZN(P2_U3252)
         );
  AOI21_X1 U8494 ( .B1(n7320), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7315), .ZN(
        n7318) );
  INV_X1 U8495 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7316) );
  MUX2_X1 U8496 ( .A(n7316), .B(P2_REG1_REG_8__SCAN_IN), .S(n7370), .Z(n7317)
         );
  AOI211_X1 U8497 ( .C1(n7318), .C2(n7317), .A(n7365), .B(n10673), .ZN(n7329)
         );
  INV_X1 U8498 ( .A(n7370), .ZN(n7448) );
  NOR2_X1 U8499 ( .A1(n10653), .A2(n7448), .ZN(n7328) );
  AOI21_X1 U8500 ( .B1(n7320), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7319), .ZN(
        n7323) );
  INV_X1 U8501 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7321) );
  MUX2_X1 U8502 ( .A(n7321), .B(P2_REG2_REG_8__SCAN_IN), .S(n7370), .Z(n7322)
         );
  NOR2_X1 U8503 ( .A1(n7323), .A2(n7322), .ZN(n7369) );
  AOI211_X1 U8504 ( .C1(n7323), .C2(n7322), .A(n7369), .B(n10677), .ZN(n7327)
         );
  INV_X1 U8505 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7325) );
  NAND2_X1 U8506 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7324) );
  OAI21_X1 U8507 ( .B1(n9217), .B2(n7325), .A(n7324), .ZN(n7326) );
  OR4_X1 U8508 ( .A1(n7329), .A2(n7328), .A3(n7327), .A4(n7326), .ZN(P2_U3253)
         );
  AOI211_X1 U8509 ( .C1(n7332), .C2(n7331), .A(n7330), .B(n10673), .ZN(n7341)
         );
  NOR2_X1 U8510 ( .A1(n10653), .A2(n7413), .ZN(n7340) );
  AOI211_X1 U8511 ( .C1(n7335), .C2(n7334), .A(n7333), .B(n10677), .ZN(n7339)
         );
  INV_X1 U8512 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7337) );
  NAND2_X1 U8513 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n7336) );
  OAI21_X1 U8514 ( .B1(n9217), .B2(n7337), .A(n7336), .ZN(n7338) );
  OR4_X1 U8515 ( .A1(n7341), .A2(n7340), .A3(n7339), .A4(n7338), .ZN(P2_U3250)
         );
  AOI211_X1 U8516 ( .C1(n7344), .C2(n7343), .A(n7342), .B(n10673), .ZN(n7352)
         );
  NOR2_X1 U8517 ( .A1(n10653), .A2(n7408), .ZN(n7351) );
  AOI211_X1 U8518 ( .C1(n7347), .C2(n7346), .A(n7345), .B(n10677), .ZN(n7350)
         );
  NAND2_X1 U8519 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n7348) );
  OAI21_X1 U8520 ( .B1(n9217), .B2(n8340), .A(n7348), .ZN(n7349) );
  OR4_X1 U8521 ( .A1(n7352), .A2(n7351), .A3(n7350), .A4(n7349), .ZN(P2_U3248)
         );
  AOI211_X1 U8522 ( .C1(n7355), .C2(n7354), .A(n7353), .B(n10673), .ZN(n7364)
         );
  NOR2_X1 U8523 ( .A1(n10653), .A2(n7418), .ZN(n7363) );
  AOI211_X1 U8524 ( .C1(n7358), .C2(n7357), .A(n7356), .B(n10677), .ZN(n7362)
         );
  INV_X1 U8525 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7360) );
  NAND2_X1 U8526 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7359) );
  OAI21_X1 U8527 ( .B1(n9217), .B2(n7360), .A(n7359), .ZN(n7361) );
  OR4_X1 U8528 ( .A1(n7364), .A2(n7363), .A3(n7362), .A4(n7361), .ZN(P2_U3249)
         );
  INV_X1 U8529 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7366) );
  MUX2_X1 U8530 ( .A(n7366), .B(P2_REG1_REG_9__SCAN_IN), .S(n7394), .Z(n7367)
         );
  AOI211_X1 U8531 ( .C1(n7368), .C2(n7367), .A(n7389), .B(n10673), .ZN(n7377)
         );
  INV_X1 U8532 ( .A(n7394), .ZN(n7452) );
  NOR2_X1 U8533 ( .A1(n10653), .A2(n7452), .ZN(n7376) );
  AOI21_X1 U8534 ( .B1(n7370), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7369), .ZN(
        n7373) );
  NAND2_X1 U8535 ( .A1(n7394), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7371) );
  OAI21_X1 U8536 ( .B1(n7394), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7371), .ZN(
        n7372) );
  NOR2_X1 U8537 ( .A1(n7373), .A2(n7372), .ZN(n7393) );
  AOI211_X1 U8538 ( .C1(n7373), .C2(n7372), .A(n7393), .B(n10677), .ZN(n7375)
         );
  INV_X1 U8539 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10568) );
  NAND2_X1 U8540 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8142) );
  OAI21_X1 U8541 ( .B1(n9217), .B2(n10568), .A(n8142), .ZN(n7374) );
  OR4_X1 U8542 ( .A1(n7377), .A2(n7376), .A3(n7375), .A4(n7374), .ZN(P2_U3254)
         );
  AOI211_X1 U8543 ( .C1(n7380), .C2(n7379), .A(n7378), .B(n10673), .ZN(n7388)
         );
  NOR2_X1 U8544 ( .A1(n10653), .A2(n7433), .ZN(n7387) );
  AOI211_X1 U8545 ( .C1(n7383), .C2(n7382), .A(n7381), .B(n10677), .ZN(n7386)
         );
  INV_X1 U8546 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7384) );
  NAND2_X1 U8547 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7971) );
  OAI21_X1 U8548 ( .B1(n9217), .B2(n7384), .A(n7971), .ZN(n7385) );
  OR4_X1 U8549 ( .A1(n7388), .A2(n7387), .A3(n7386), .A4(n7385), .ZN(P2_U3251)
         );
  INV_X1 U8550 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7390) );
  MUX2_X1 U8551 ( .A(n7390), .B(P2_REG1_REG_10__SCAN_IN), .S(n7873), .Z(n7391)
         );
  NOR2_X1 U8552 ( .A1(n7392), .A2(n7391), .ZN(n7867) );
  AOI211_X1 U8553 ( .C1(n7392), .C2(n7391), .A(n7867), .B(n10673), .ZN(n7403)
         );
  INV_X1 U8554 ( .A(n7873), .ZN(n7537) );
  NOR2_X1 U8555 ( .A1(n10653), .A2(n7537), .ZN(n7402) );
  AOI21_X1 U8556 ( .B1(n7394), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7393), .ZN(
        n7398) );
  INV_X1 U8557 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7395) );
  MUX2_X1 U8558 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7395), .S(n7873), .Z(n7396)
         );
  INV_X1 U8559 ( .A(n7396), .ZN(n7397) );
  NOR2_X1 U8560 ( .A1(n7398), .A2(n7397), .ZN(n7872) );
  AOI211_X1 U8561 ( .C1(n7398), .C2(n7397), .A(n7872), .B(n10677), .ZN(n7401)
         );
  INV_X1 U8562 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U8563 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7399) );
  OAI21_X1 U8564 ( .B1(n9217), .B2(n8338), .A(n7399), .ZN(n7400) );
  OR4_X1 U8565 ( .A1(n7403), .A2(n7402), .A3(n7401), .A4(n7400), .ZN(P2_U3255)
         );
  AND2_X1 U8566 ( .A1(n7404), .A2(P1_U3084), .ZN(n8294) );
  OAI222_X1 U8567 ( .A1(n9004), .A2(n5287), .B1(n5033), .B2(n7409), .C1(
        P1_U3084), .C2(n7405), .ZN(P1_U3350) );
  OAI222_X1 U8568 ( .A1(n7480), .A2(P1_U3084), .B1(n5033), .B2(n7417), .C1(
        n9004), .C2(n5770), .ZN(P1_U3349) );
  OAI222_X1 U8569 ( .A1(n9004), .A2(n7407), .B1(n5033), .B2(n7412), .C1(
        P1_U3084), .C2(n7406), .ZN(P1_U3348) );
  NOR2_X1 U8570 ( .A1(n5768), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10010) );
  INV_X2 U8571 ( .A(n10010), .ZN(n10005) );
  INV_X1 U8572 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7410) );
  NAND2_X1 U8573 ( .A1(n5768), .A2(P2_U3152), .ZN(n10012) );
  OAI222_X1 U8574 ( .A1(n10005), .A2(n7410), .B1(n10012), .B2(n7409), .C1(
        n7408), .C2(P2_U3152), .ZN(P2_U3355) );
  OAI222_X1 U8575 ( .A1(n7413), .A2(P2_U3152), .B1(n10012), .B2(n7412), .C1(
        n7411), .C2(n10005), .ZN(P2_U3353) );
  INV_X1 U8576 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7415) );
  OAI222_X1 U8577 ( .A1(n10005), .A2(n7415), .B1(n10012), .B2(n7422), .C1(
        n7414), .C2(P2_U3152), .ZN(P2_U3356) );
  OAI222_X1 U8578 ( .A1(n7418), .A2(P2_U3152), .B1(n10012), .B2(n7417), .C1(
        n7416), .C2(n10005), .ZN(P2_U3354) );
  OAI222_X1 U8579 ( .A1(n9004), .A2(n7420), .B1(n5033), .B2(n7432), .C1(
        P1_U3084), .C2(n7419), .ZN(P1_U3347) );
  OAI222_X1 U8580 ( .A1(n9004), .A2(n7421), .B1(n5033), .B2(n7431), .C1(
        P1_U3084), .C2(n10625), .ZN(P1_U3352) );
  INV_X1 U8581 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7423) );
  OAI222_X1 U8582 ( .A1(n9004), .A2(n7423), .B1(n5033), .B2(n7422), .C1(
        P1_U3084), .C2(n7478), .ZN(P1_U3351) );
  INV_X1 U8583 ( .A(n7577), .ZN(n7425) );
  INV_X1 U8584 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n7429) );
  NAND2_X1 U8585 ( .A1(n8594), .A2(n7426), .ZN(n7427) );
  NOR2_X1 U8586 ( .A1(n6395), .A2(n7427), .ZN(n7428) );
  AOI21_X1 U8587 ( .B1(n10545), .B2(n7429), .A(n7428), .ZN(P1_U3441) );
  INV_X1 U8588 ( .A(n10012), .ZN(n8297) );
  INV_X1 U8589 ( .A(n8297), .ZN(n8693) );
  OAI222_X1 U8590 ( .A1(n10005), .A2(n6459), .B1(n8693), .B2(n7431), .C1(n7430), .C2(P2_U3152), .ZN(P2_U3357) );
  OAI222_X1 U8591 ( .A1(n7433), .A2(P2_U3152), .B1(n8693), .B2(n7432), .C1(
        n10005), .C2(n6574), .ZN(P2_U3352) );
  INV_X1 U8592 ( .A(n7434), .ZN(n7437) );
  OAI222_X1 U8593 ( .A1(n7436), .A2(P2_U3152), .B1(n10012), .B2(n7437), .C1(
        n7435), .C2(n10005), .ZN(P2_U3351) );
  INV_X1 U8594 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7438) );
  INV_X1 U8595 ( .A(n7510), .ZN(n7485) );
  OAI222_X1 U8596 ( .A1(n9004), .A2(n7438), .B1(n5033), .B2(n7437), .C1(
        P1_U3084), .C2(n7485), .ZN(P1_U3346) );
  NAND2_X1 U8597 ( .A1(n10545), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7439) );
  OAI21_X1 U8598 ( .B1(n10545), .B2(n7440), .A(n7439), .ZN(P1_U3440) );
  NAND2_X1 U8599 ( .A1(n7734), .A2(P1_U4006), .ZN(n7441) );
  OAI21_X1 U8600 ( .B1(P1_U4006), .B2(n6574), .A(n7441), .ZN(P1_U3561) );
  NAND2_X1 U8601 ( .A1(n10146), .A2(P1_U4006), .ZN(n7442) );
  OAI21_X1 U8602 ( .B1(n6047), .B2(P1_U4006), .A(n7442), .ZN(P1_U3571) );
  INV_X1 U8603 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U8604 ( .A1(n8659), .A2(P1_U4006), .ZN(n7443) );
  OAI21_X1 U8605 ( .B1(n7688), .B2(P1_U4006), .A(n7443), .ZN(P1_U3570) );
  INV_X1 U8606 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7445) );
  INV_X1 U8607 ( .A(n7444), .ZN(n7447) );
  INV_X1 U8608 ( .A(n7488), .ZN(n7546) );
  OAI222_X1 U8609 ( .A1(n9004), .A2(n7445), .B1(n5033), .B2(n7447), .C1(
        P1_U3084), .C2(n7546), .ZN(P1_U3345) );
  INV_X1 U8610 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7446) );
  OAI222_X1 U8611 ( .A1(n7448), .A2(P2_U3152), .B1(n10012), .B2(n7447), .C1(
        n7446), .C2(n10005), .ZN(P2_U3350) );
  INV_X1 U8612 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U8613 ( .A1(n11004), .A2(P1_U4006), .ZN(n7449) );
  OAI21_X1 U8614 ( .B1(n7671), .B2(P1_U4006), .A(n7449), .ZN(P1_U3569) );
  INV_X1 U8615 ( .A(n7450), .ZN(n7453) );
  OAI222_X1 U8616 ( .A1(n7452), .A2(P2_U3152), .B1(n8693), .B2(n7453), .C1(
        n7451), .C2(n10005), .ZN(P2_U3349) );
  INV_X1 U8617 ( .A(n7500), .ZN(n7563) );
  OAI222_X1 U8618 ( .A1(n9004), .A2(n9750), .B1(n5033), .B2(n7453), .C1(
        P1_U3084), .C2(n7563), .ZN(P1_U3344) );
  NOR2_X1 U8619 ( .A1(n7510), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7466) );
  NAND2_X1 U8620 ( .A1(n10595), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7464) );
  INV_X1 U8621 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7454) );
  MUX2_X1 U8622 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n7454), .S(n10595), .Z(n10602) );
  INV_X1 U8623 ( .A(n7480), .ZN(n7643) );
  NAND2_X1 U8624 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n10610), .ZN(n7459) );
  INV_X1 U8625 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7455) );
  MUX2_X1 U8626 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7455), .S(n10610), .Z(n10617) );
  NAND2_X1 U8627 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(n10691), .ZN(n7458) );
  INV_X1 U8628 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7456) );
  MUX2_X1 U8629 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n7456), .S(n10691), .Z(n10690) );
  INV_X1 U8630 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10720) );
  OR2_X1 U8631 ( .A1(n10625), .A2(n10720), .ZN(n7457) );
  MUX2_X1 U8632 ( .A(n10720), .B(P1_REG1_REG_1__SCAN_IN), .S(n10625), .Z(
        n10636) );
  NAND3_X1 U8633 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n10636), .ZN(n10634) );
  NAND2_X1 U8634 ( .A1(n7457), .A2(n10634), .ZN(n10689) );
  NAND2_X1 U8635 ( .A1(n10690), .A2(n10689), .ZN(n10688) );
  NAND2_X1 U8636 ( .A1(n7458), .A2(n10688), .ZN(n10618) );
  NAND2_X1 U8637 ( .A1(n10617), .A2(n10618), .ZN(n10616) );
  NAND2_X1 U8638 ( .A1(n7459), .A2(n10616), .ZN(n7637) );
  INV_X1 U8639 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7460) );
  MUX2_X1 U8640 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7460), .S(n7480), .Z(n7636)
         );
  NOR2_X1 U8641 ( .A1(n7637), .A2(n7636), .ZN(n7635) );
  INV_X1 U8642 ( .A(n7635), .ZN(n7461) );
  OAI21_X1 U8643 ( .B1(n7643), .B2(P1_REG1_REG_4__SCAN_IN), .A(n7461), .ZN(
        n7529) );
  INV_X1 U8644 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10798) );
  MUX2_X1 U8645 ( .A(n10798), .B(P1_REG1_REG_5__SCAN_IN), .S(n7532), .Z(n7528)
         );
  NOR2_X1 U8646 ( .A1(n7529), .A2(n7528), .ZN(n7527) );
  INV_X1 U8647 ( .A(n7527), .ZN(n7463) );
  NAND2_X1 U8648 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n7532), .ZN(n7462) );
  NAND2_X1 U8649 ( .A1(n7463), .A2(n7462), .ZN(n10603) );
  NAND2_X1 U8650 ( .A1(n10602), .A2(n10603), .ZN(n10601) );
  NAND2_X1 U8651 ( .A1(n7464), .A2(n10601), .ZN(n7515) );
  INV_X1 U8652 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7465) );
  MUX2_X1 U8653 ( .A(n7465), .B(P1_REG1_REG_7__SCAN_IN), .S(n7510), .Z(n7514)
         );
  NOR2_X1 U8654 ( .A1(n7515), .A2(n7514), .ZN(n7513) );
  OR2_X1 U8655 ( .A1(n7466), .A2(n7513), .ZN(n7549) );
  INV_X1 U8656 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10887) );
  MUX2_X1 U8657 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10887), .S(n7488), .Z(n7550)
         );
  NAND2_X1 U8658 ( .A1(n7549), .A2(n7550), .ZN(n7548) );
  NAND2_X1 U8659 ( .A1(n7546), .A2(n10887), .ZN(n7468) );
  INV_X1 U8660 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7467) );
  MUX2_X1 U8661 ( .A(n7467), .B(P1_REG1_REG_9__SCAN_IN), .S(n7500), .Z(n7469)
         );
  AOI21_X1 U8662 ( .B1(n7548), .B2(n7468), .A(n7469), .ZN(n7559) );
  AND3_X1 U8663 ( .A1(n7548), .A2(n7469), .A3(n7468), .ZN(n7472) );
  AND2_X1 U8664 ( .A1(n5035), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7471) );
  NAND2_X1 U8665 ( .A1(n7492), .A2(n7471), .ZN(n10593) );
  INV_X1 U8666 ( .A(n10259), .ZN(n10590) );
  OAI21_X1 U8667 ( .B1(n7559), .B2(n7472), .A(n10635), .ZN(n7506) );
  NOR2_X1 U8668 ( .A1(n7510), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7487) );
  NAND2_X1 U8669 ( .A1(n10595), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7484) );
  INV_X1 U8670 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7473) );
  MUX2_X1 U8671 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7473), .S(n10595), .Z(n10605) );
  NAND2_X1 U8672 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n10610), .ZN(n7479) );
  INV_X1 U8673 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7474) );
  MUX2_X1 U8674 ( .A(n7474), .B(P1_REG2_REG_3__SCAN_IN), .S(n10610), .Z(n7475)
         );
  INV_X1 U8675 ( .A(n7475), .ZN(n10620) );
  INV_X1 U8676 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7477) );
  XNOR2_X1 U8677 ( .A(n7478), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n10702) );
  INV_X1 U8678 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7476) );
  MUX2_X1 U8679 ( .A(n7476), .B(P1_REG2_REG_1__SCAN_IN), .S(n10625), .Z(n10639) );
  NAND3_X1 U8680 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .A3(n10639), .ZN(n10638) );
  OAI21_X1 U8681 ( .B1(n10625), .B2(n7476), .A(n10638), .ZN(n10701) );
  NAND2_X1 U8682 ( .A1(n10702), .A2(n10701), .ZN(n10699) );
  OAI21_X1 U8683 ( .B1(n7478), .B2(n7477), .A(n10699), .ZN(n10621) );
  NAND2_X1 U8684 ( .A1(n10620), .A2(n10621), .ZN(n10619) );
  NAND2_X1 U8685 ( .A1(n7479), .A2(n10619), .ZN(n7640) );
  INV_X1 U8686 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7481) );
  MUX2_X1 U8687 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7481), .S(n7480), .Z(n7639)
         );
  NOR2_X1 U8688 ( .A1(n7640), .A2(n7639), .ZN(n7638) );
  NOR2_X1 U8689 ( .A1(n7643), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7522) );
  INV_X1 U8690 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7775) );
  MUX2_X1 U8691 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7775), .S(n7532), .Z(n7521)
         );
  OAI21_X1 U8692 ( .B1(n7638), .B2(n7522), .A(n7521), .ZN(n7525) );
  INV_X1 U8693 ( .A(n7525), .ZN(n7483) );
  NOR2_X1 U8694 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n7532), .ZN(n7482) );
  NOR2_X1 U8695 ( .A1(n7483), .A2(n7482), .ZN(n10606) );
  NAND2_X1 U8696 ( .A1(n10605), .A2(n10606), .ZN(n10604) );
  NAND2_X1 U8697 ( .A1(n7484), .A2(n10604), .ZN(n7509) );
  INV_X1 U8698 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7486) );
  AOI22_X1 U8699 ( .A1(n7510), .A2(n7486), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n7485), .ZN(n7508) );
  NOR2_X1 U8700 ( .A1(n7509), .A2(n7508), .ZN(n7507) );
  NOR2_X1 U8701 ( .A1(n7487), .A2(n7507), .ZN(n7544) );
  INV_X1 U8702 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7489) );
  MUX2_X1 U8703 ( .A(n7489), .B(P1_REG2_REG_8__SCAN_IN), .S(n7488), .Z(n7543)
         );
  OR2_X1 U8704 ( .A1(n7544), .A2(n7543), .ZN(n7541) );
  NAND2_X1 U8705 ( .A1(n7546), .A2(n7489), .ZN(n7490) );
  NAND2_X1 U8706 ( .A1(n7541), .A2(n7490), .ZN(n7494) );
  INV_X1 U8707 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7491) );
  MUX2_X1 U8708 ( .A(n7491), .B(P1_REG2_REG_9__SCAN_IN), .S(n7500), .Z(n7493)
         );
  NOR2_X1 U8709 ( .A1(n10259), .A2(P1_U3084), .ZN(n8691) );
  NAND2_X1 U8710 ( .A1(n7492), .A2(n8691), .ZN(n7609) );
  OR2_X1 U8711 ( .A1(n7609), .A2(n5036), .ZN(n10248) );
  AOI21_X1 U8712 ( .B1(n7494), .B2(n7493), .A(n10248), .ZN(n7504) );
  INV_X1 U8713 ( .A(n7495), .ZN(n7496) );
  NOR2_X1 U8714 ( .A1(n7497), .A2(n7496), .ZN(n7498) );
  INV_X1 U8715 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7502) );
  INV_X1 U8716 ( .A(n7609), .ZN(n7499) );
  AND2_X1 U8717 ( .A1(n7499), .A2(n5036), .ZN(n10692) );
  NAND2_X1 U8718 ( .A1(n10692), .A2(n7500), .ZN(n7501) );
  NAND2_X1 U8719 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8019) );
  OAI211_X1 U8720 ( .C1(n10631), .C2(n7502), .A(n7501), .B(n8019), .ZN(n7503)
         );
  AOI21_X1 U8721 ( .B1(n7504), .B2(n7562), .A(n7503), .ZN(n7505) );
  NAND2_X1 U8722 ( .A1(n7506), .A2(n7505), .ZN(P1_U3250) );
  AOI21_X1 U8723 ( .B1(n7509), .B2(n7508), .A(n7507), .ZN(n7520) );
  INV_X1 U8724 ( .A(n10631), .ZN(n10698) );
  NAND2_X1 U8725 ( .A1(n10692), .A2(n7510), .ZN(n7512) );
  AND2_X1 U8726 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7842) );
  INV_X1 U8727 ( .A(n7842), .ZN(n7511) );
  NAND2_X1 U8728 ( .A1(n7512), .A2(n7511), .ZN(n7518) );
  AOI21_X1 U8729 ( .B1(n7515), .B2(n7514), .A(n7513), .ZN(n7516) );
  NOR2_X1 U8730 ( .A1(n7516), .A2(n10695), .ZN(n7517) );
  AOI211_X1 U8731 ( .C1(n10698), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7518), .B(
        n7517), .ZN(n7519) );
  OAI21_X1 U8732 ( .B1(n7520), .B2(n10248), .A(n7519), .ZN(P1_U3248) );
  INV_X1 U8733 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7535) );
  INV_X1 U8734 ( .A(n10248), .ZN(n10700) );
  INV_X1 U8735 ( .A(n7521), .ZN(n7524) );
  INV_X1 U8736 ( .A(n7522), .ZN(n7523) );
  NAND2_X1 U8737 ( .A1(n7524), .A2(n7523), .ZN(n7526) );
  OAI21_X1 U8738 ( .B1(n7638), .B2(n7526), .A(n7525), .ZN(n7531) );
  AOI211_X1 U8739 ( .C1(n7529), .C2(n7528), .A(n7527), .B(n10695), .ZN(n7530)
         );
  AOI21_X1 U8740 ( .B1(n10700), .B2(n7531), .A(n7530), .ZN(n7534) );
  AND2_X1 U8741 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7733) );
  AOI21_X1 U8742 ( .B1(n10692), .B2(n7532), .A(n7733), .ZN(n7533) );
  OAI211_X1 U8743 ( .C1(n7535), .C2(n10631), .A(n7534), .B(n7533), .ZN(
        P1_U3246) );
  INV_X1 U8744 ( .A(n7536), .ZN(n7539) );
  OAI222_X1 U8745 ( .A1(n10005), .A2(n7538), .B1(n8693), .B2(n7539), .C1(n7537), .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8746 ( .A(n7606), .ZN(n7603) );
  OAI222_X1 U8747 ( .A1(n9004), .A2(n7540), .B1(n5033), .B2(n7539), .C1(
        P1_U3084), .C2(n7603), .ZN(P1_U3343) );
  INV_X1 U8748 ( .A(n7541), .ZN(n7542) );
  AOI21_X1 U8749 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n7554) );
  INV_X1 U8750 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7545) );
  NOR2_X1 U8751 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7545), .ZN(n8122) );
  INV_X1 U8752 ( .A(n10692), .ZN(n10251) );
  NOR2_X1 U8753 ( .A1(n10251), .A2(n7546), .ZN(n7547) );
  AOI211_X1 U8754 ( .C1(n10698), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n8122), .B(
        n7547), .ZN(n7553) );
  OAI21_X1 U8755 ( .B1(n7550), .B2(n7549), .A(n7548), .ZN(n7551) );
  NAND2_X1 U8756 ( .A1(n7551), .A2(n10635), .ZN(n7552) );
  OAI211_X1 U8757 ( .C1(n7554), .C2(n10248), .A(n7553), .B(n7552), .ZN(
        P1_U3249) );
  INV_X1 U8758 ( .A(n7555), .ZN(n7558) );
  INV_X1 U8759 ( .A(n7881), .ZN(n7617) );
  INV_X1 U8760 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7556) );
  OAI222_X1 U8761 ( .A1(n5033), .A2(n7558), .B1(n7617), .B2(P1_U3084), .C1(
        n7556), .C2(n9004), .ZN(P1_U3342) );
  INV_X1 U8762 ( .A(n7991), .ZN(n7880) );
  INV_X1 U8763 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7557) );
  OAI222_X1 U8764 ( .A1(P2_U3152), .A2(n7880), .B1(n8693), .B2(n7558), .C1(
        n7557), .C2(n10005), .ZN(P2_U3347) );
  AOI21_X1 U8765 ( .B1(n7467), .B2(n7563), .A(n7559), .ZN(n7561) );
  INV_X1 U8766 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8318) );
  AOI22_X1 U8767 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n7603), .B1(n7606), .B2(
        n8318), .ZN(n7560) );
  NOR2_X1 U8768 ( .A1(n7561), .A2(n7560), .ZN(n7602) );
  AOI21_X1 U8769 ( .B1(n7561), .B2(n7560), .A(n7602), .ZN(n7574) );
  INV_X1 U8770 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7571) );
  OAI21_X1 U8771 ( .B1(n7563), .B2(n7491), .A(n7562), .ZN(n7567) );
  INV_X1 U8772 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7564) );
  MUX2_X1 U8773 ( .A(n7564), .B(P1_REG2_REG_10__SCAN_IN), .S(n7606), .Z(n7565)
         );
  INV_X1 U8774 ( .A(n7565), .ZN(n7566) );
  NAND2_X1 U8775 ( .A1(n7566), .A2(n7567), .ZN(n7607) );
  OAI211_X1 U8776 ( .C1(n7567), .C2(n7566), .A(n10700), .B(n7607), .ZN(n7570)
         );
  NOR2_X1 U8777 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7568), .ZN(n8464) );
  AOI21_X1 U8778 ( .B1(n10692), .B2(n7606), .A(n8464), .ZN(n7569) );
  OAI211_X1 U8779 ( .C1(n10631), .C2(n7571), .A(n7570), .B(n7569), .ZN(n7572)
         );
  INV_X1 U8780 ( .A(n7572), .ZN(n7573) );
  OAI21_X1 U8781 ( .B1(n7574), .B2(n10695), .A(n7573), .ZN(P1_U3251) );
  NAND2_X1 U8782 ( .A1(n7693), .A2(n7575), .ZN(n7579) );
  OR2_X1 U8783 ( .A1(n7577), .A2(n7576), .ZN(n7596) );
  INV_X1 U8784 ( .A(n7702), .ZN(n7695) );
  INV_X1 U8785 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7587) );
  OR2_X1 U8786 ( .A1(n7581), .A2(n7580), .ZN(n7582) );
  NAND2_X1 U8787 ( .A1(n7582), .A2(n7585), .ZN(n7713) );
  OAI22_X1 U8788 ( .A1(n7583), .A2(n7713), .B1(n7851), .B2(n10851), .ZN(n7699)
         );
  INV_X1 U8789 ( .A(n7699), .ZN(n7584) );
  OAI21_X1 U8790 ( .B1(n7021), .B2(n7585), .A(n7584), .ZN(n7589) );
  NAND2_X1 U8791 ( .A1(n7589), .A2(n11097), .ZN(n7586) );
  OAI21_X1 U8792 ( .B1(n11097), .B2(n7587), .A(n7586), .ZN(P1_U3454) );
  NAND2_X1 U8793 ( .A1(n7589), .A2(n11093), .ZN(n7590) );
  OAI21_X1 U8794 ( .B1(n11093), .B2(n5666), .A(n7590), .ZN(P1_U3523) );
  XNOR2_X1 U8795 ( .A(n7592), .B(n7591), .ZN(n7594) );
  XNOR2_X1 U8796 ( .A(n7594), .B(n5708), .ZN(n7601) );
  INV_X1 U8797 ( .A(n10149), .ZN(n10115) );
  AOI22_X1 U8798 ( .A1(n10147), .A2(n5727), .B1(n10115), .B2(n7119), .ZN(n7600) );
  INV_X1 U8799 ( .A(n7595), .ZN(n7598) );
  OR3_X1 U8800 ( .A1(n7598), .A2(n7597), .A3(n7596), .ZN(n8724) );
  AOI22_X1 U8801 ( .A1(n7216), .A2(n10131), .B1(n8724), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7599) );
  OAI211_X1 U8802 ( .C1(n7601), .C2(n10133), .A(n7600), .B(n7599), .ZN(
        P1_U3220) );
  AOI21_X1 U8803 ( .B1(n8318), .B2(n7603), .A(n7602), .ZN(n7605) );
  INV_X1 U8804 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U8805 ( .A1(n7881), .A2(n10970), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n7617), .ZN(n7604) );
  NOR2_X1 U8806 ( .A1(n7605), .A2(n7604), .ZN(n10179) );
  AOI21_X1 U8807 ( .B1(n7605), .B2(n7604), .A(n10179), .ZN(n7623) );
  NAND2_X1 U8808 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7606), .ZN(n7608) );
  NAND2_X1 U8809 ( .A1(n7608), .A2(n7607), .ZN(n7614) );
  NAND2_X1 U8810 ( .A1(n7614), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7613) );
  OAI21_X1 U8811 ( .B1(n7613), .B2(n7609), .A(n10251), .ZN(n7612) );
  AND2_X1 U8812 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8224) );
  INV_X1 U8813 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7610) );
  NOR2_X1 U8814 ( .A1(n10631), .A2(n7610), .ZN(n7611) );
  AOI211_X1 U8815 ( .C1(n7612), .C2(n7881), .A(n8224), .B(n7611), .ZN(n7622)
         );
  NAND2_X1 U8816 ( .A1(n7613), .A2(n7617), .ZN(n7616) );
  INV_X1 U8817 ( .A(n7614), .ZN(n7619) );
  INV_X1 U8818 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7618) );
  NAND2_X1 U8819 ( .A1(n7619), .A2(n7618), .ZN(n7615) );
  NAND2_X1 U8820 ( .A1(n7616), .A2(n7615), .ZN(n10186) );
  NAND3_X1 U8821 ( .A1(n7619), .A2(n7618), .A3(n7617), .ZN(n7620) );
  NAND3_X1 U8822 ( .A1(n10186), .A2(n10700), .A3(n7620), .ZN(n7621) );
  OAI211_X1 U8823 ( .C1(n7623), .C2(n10695), .A(n7622), .B(n7621), .ZN(
        P1_U3252) );
  INV_X1 U8824 ( .A(n7624), .ZN(n7626) );
  AOI22_X1 U8825 ( .A1(n8015), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n10010), .ZN(n7625) );
  OAI21_X1 U8826 ( .B1(n7626), .B2(n10012), .A(n7625), .ZN(P2_U3346) );
  INV_X1 U8827 ( .A(n10185), .ZN(n7882) );
  OAI222_X1 U8828 ( .A1(n9004), .A2(n7627), .B1(n5033), .B2(n7626), .C1(
        P1_U3084), .C2(n7882), .ZN(P1_U3341) );
  INV_X1 U8829 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7708) );
  NOR2_X1 U8830 ( .A1(n10633), .A2(n7708), .ZN(n10640) );
  OAI21_X1 U8831 ( .B1(n7630), .B2(n7629), .A(n7628), .ZN(n8723) );
  INV_X1 U8832 ( .A(n8723), .ZN(n7631) );
  MUX2_X1 U8833 ( .A(n10640), .B(n7631), .S(n10259), .Z(n7634) );
  AOI21_X1 U8834 ( .B1(n10590), .B2(n7708), .A(n5036), .ZN(n10589) );
  OAI21_X1 U8835 ( .B1(n10589), .B2(P1_IR_REG_0__SCAN_IN), .A(P1_U4006), .ZN(
        n7632) );
  AOI21_X1 U8836 ( .B1(n7634), .B2(n7633), .A(n7632), .ZN(n10696) );
  AOI21_X1 U8837 ( .B1(n7637), .B2(n7636), .A(n7635), .ZN(n7642) );
  AOI21_X1 U8838 ( .B1(n7640), .B2(n7639), .A(n7638), .ZN(n7641) );
  OAI22_X1 U8839 ( .A1(n7642), .A2(n10695), .B1(n10248), .B2(n7641), .ZN(n7646) );
  INV_X1 U8840 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8339) );
  AND2_X1 U8841 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7681) );
  AOI21_X1 U8842 ( .B1(n10692), .B2(n7643), .A(n7681), .ZN(n7644) );
  OAI21_X1 U8843 ( .B1(n8339), .B2(n10631), .A(n7644), .ZN(n7645) );
  OR3_X1 U8844 ( .A1(n10696), .A2(n7646), .A3(n7645), .ZN(P1_U3245) );
  INV_X1 U8845 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7899) );
  INV_X1 U8846 ( .A(n9876), .ZN(n7647) );
  NAND2_X1 U8847 ( .A1(n7647), .A2(P2_U3966), .ZN(n7648) );
  OAI21_X1 U8848 ( .B1(n7899), .B2(P2_U3966), .A(n7648), .ZN(P2_U3570) );
  INV_X1 U8849 ( .A(n8326), .ZN(n8248) );
  NAND2_X1 U8850 ( .A1(n8248), .A2(P2_U3966), .ZN(n7649) );
  OAI21_X1 U8851 ( .B1(n5770), .B2(P2_U3966), .A(n7649), .ZN(P2_U3556) );
  INV_X1 U8852 ( .A(n7650), .ZN(n7651) );
  AOI21_X1 U8853 ( .B1(n7653), .B2(n7652), .A(n7651), .ZN(n7656) );
  AOI22_X1 U8854 ( .A1(n10115), .A2(n5704), .B1(n10147), .B2(n10175), .ZN(
        n7655) );
  AOI22_X1 U8855 ( .A1(n7024), .A2(n10131), .B1(n8724), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7654) );
  OAI211_X1 U8856 ( .C1(n7656), .C2(n10133), .A(n7655), .B(n7654), .ZN(
        P1_U3235) );
  INV_X1 U8857 ( .A(n7657), .ZN(n7662) );
  INV_X1 U8858 ( .A(n9004), .ZN(n10537) );
  AOI22_X1 U8859 ( .A1(n10201), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10537), .ZN(n7658) );
  OAI21_X1 U8860 ( .B1(n7662), .B2(n5033), .A(n7658), .ZN(P1_U3340) );
  NOR2_X1 U8861 ( .A1(n10672), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8862 ( .A(n7659), .ZN(n7670) );
  AOI22_X1 U8863 ( .A1(n10217), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10537), .ZN(n7660) );
  OAI21_X1 U8864 ( .B1(n7670), .B2(n5033), .A(n7660), .ZN(P1_U3339) );
  INV_X1 U8865 ( .A(n8110), .ZN(n7997) );
  OAI222_X1 U8866 ( .A1(P2_U3152), .A2(n7997), .B1(n8693), .B2(n7662), .C1(
        n7661), .C2(n10005), .ZN(P2_U3345) );
  INV_X1 U8867 ( .A(n10152), .ZN(n10098) );
  OAI21_X1 U8868 ( .B1(n7665), .B2(n7664), .A(n7663), .ZN(n7666) );
  NAND2_X1 U8869 ( .A1(n7666), .A2(n10143), .ZN(n7669) );
  NOR2_X1 U8870 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5745), .ZN(n10611) );
  OAI22_X1 U8871 ( .A1(n10156), .A2(n7759), .B1(n7745), .B2(n10149), .ZN(n7667) );
  AOI211_X1 U8872 ( .C1(n10147), .C2(n10174), .A(n10611), .B(n7667), .ZN(n7668) );
  OAI211_X1 U8873 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n10098), .A(n7669), .B(
        n7668), .ZN(P1_U3216) );
  INV_X1 U8874 ( .A(n9170), .ZN(n8118) );
  OAI222_X1 U8875 ( .A1(n8118), .A2(P2_U3152), .B1(n10005), .B2(n7671), .C1(
        n7670), .C2(n10012), .ZN(P2_U3344) );
  NAND2_X1 U8876 ( .A1(n6549), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U8877 ( .A1(n5060), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U8878 ( .A1(n6533), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7672) );
  AND3_X1 U8879 ( .A1(n7674), .A2(n7673), .A3(n7672), .ZN(n9271) );
  NAND2_X1 U8880 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n9160), .ZN(n7675) );
  OAI21_X1 U8881 ( .B1(n9271), .B2(n9160), .A(n7675), .ZN(P2_U3582) );
  NAND2_X1 U8882 ( .A1(n7677), .A2(n7676), .ZN(n7679) );
  XOR2_X1 U8883 ( .A(n7679), .B(n7678), .Z(n7684) );
  OAI22_X1 U8884 ( .A1(n10156), .A2(n10758), .B1(n7852), .B2(n10149), .ZN(
        n7680) );
  AOI211_X1 U8885 ( .C1(n10147), .C2(n10173), .A(n7681), .B(n7680), .ZN(n7683)
         );
  NAND2_X1 U8886 ( .A1(n10152), .A2(n7784), .ZN(n7682) );
  OAI211_X1 U8887 ( .C1(n7684), .C2(n10133), .A(n7683), .B(n7682), .ZN(
        P1_U3228) );
  NAND2_X1 U8888 ( .A1(n10052), .A2(P1_U4006), .ZN(n7685) );
  OAI21_X1 U8889 ( .B1(n6865), .B2(P1_U4006), .A(n7685), .ZN(P1_U3581) );
  INV_X1 U8890 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7687) );
  INV_X1 U8891 ( .A(n7686), .ZN(n7689) );
  INV_X1 U8892 ( .A(n8061), .ZN(n8053) );
  OAI222_X1 U8893 ( .A1(n9004), .A2(n7687), .B1(n5033), .B2(n7689), .C1(
        P1_U3084), .C2(n8053), .ZN(P1_U3338) );
  OAI222_X1 U8894 ( .A1(n9187), .A2(P2_U3152), .B1(n8693), .B2(n7689), .C1(
        n10005), .C2(n7688), .ZN(P2_U3343) );
  INV_X1 U8895 ( .A(n7690), .ZN(n7692) );
  AOI22_X1 U8896 ( .A1(n8499), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10537), .ZN(n7691) );
  OAI21_X1 U8897 ( .B1(n7692), .B2(n5033), .A(n7691), .ZN(P1_U3337) );
  INV_X1 U8898 ( .A(n9202), .ZN(n9185) );
  OAI222_X1 U8899 ( .A1(n9185), .A2(P2_U3152), .B1(n8693), .B2(n7692), .C1(
        n10005), .C2(n6047), .ZN(P2_U3342) );
  NOR2_X1 U8900 ( .A1(n7694), .A2(n7693), .ZN(n7704) );
  NAND2_X1 U8901 ( .A1(n7704), .A2(n7695), .ZN(n7696) );
  INV_X1 U8902 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7697) );
  NOR2_X1 U8903 ( .A1(n10865), .A2(n7697), .ZN(n7698) );
  OAI21_X1 U8904 ( .B1(n7699), .B2(n7698), .A(n10869), .ZN(n7707) );
  INV_X1 U8905 ( .A(n7700), .ZN(n7701) );
  NOR2_X1 U8906 ( .A1(n7702), .A2(n10344), .ZN(n7703) );
  AND2_X1 U8907 ( .A1(n7704), .A2(n7703), .ZN(n10439) );
  INV_X1 U8908 ( .A(n7021), .ZN(n7724) );
  OAI21_X1 U8909 ( .B1(n10413), .B2(n11022), .A(n7724), .ZN(n7706) );
  OAI211_X1 U8910 ( .C1(n7708), .C2(n10869), .A(n7707), .B(n7706), .ZN(
        P1_U3291) );
  NAND2_X1 U8911 ( .A1(n7119), .A2(n7724), .ZN(n7709) );
  XNOR2_X1 U8912 ( .A(n7715), .B(n7709), .ZN(n10714) );
  NOR2_X1 U8913 ( .A1(n7710), .A2(n10392), .ZN(n7749) );
  NAND2_X1 U8914 ( .A1(n10869), .A2(n7749), .ZN(n10419) );
  NAND2_X1 U8915 ( .A1(n8291), .A2(n7710), .ZN(n7711) );
  NAND2_X1 U8916 ( .A1(n7711), .A2(n10392), .ZN(n7712) );
  INV_X1 U8917 ( .A(n10851), .ZN(n11003) );
  AOI22_X1 U8918 ( .A1(n11006), .A2(n7119), .B1(n5727), .B2(n11003), .ZN(n7723) );
  XNOR2_X1 U8919 ( .A(n7715), .B(n7714), .ZN(n7721) );
  NAND2_X1 U8920 ( .A1(n7716), .A2(n10344), .ZN(n7720) );
  NAND2_X1 U8921 ( .A1(n7718), .A2(n7717), .ZN(n7719) );
  NAND2_X1 U8922 ( .A1(n7720), .A2(n7719), .ZN(n11009) );
  NAND2_X1 U8923 ( .A1(n7721), .A2(n11009), .ZN(n7722) );
  OAI211_X1 U8924 ( .C1(n10714), .C2(n11013), .A(n7723), .B(n7722), .ZN(n10717) );
  NAND2_X1 U8925 ( .A1(n10716), .A2(n7021), .ZN(n7752) );
  INV_X1 U8926 ( .A(n7752), .ZN(n7857) );
  OR3_X1 U8927 ( .A1(n7857), .A2(n7742), .A3(n11085), .ZN(n10715) );
  INV_X1 U8928 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10627) );
  OAI22_X1 U8929 ( .A1(n10715), .A2(n10344), .B1(n10627), .B2(n10865), .ZN(
        n7725) );
  OAI21_X1 U8930 ( .B1(n10717), .B2(n7725), .A(n10869), .ZN(n7727) );
  AOI22_X1 U8931 ( .A1(n10413), .A2(n7216), .B1(n11027), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7726) );
  OAI211_X1 U8932 ( .C1(n10714), .C2(n10419), .A(n7727), .B(n7726), .ZN(
        P1_U3290) );
  NAND2_X1 U8933 ( .A1(n7729), .A2(n7728), .ZN(n7731) );
  XNOR2_X1 U8934 ( .A(n7731), .B(n7730), .ZN(n7737) );
  OAI22_X1 U8935 ( .A1(n10156), .A2(n10794), .B1(n7772), .B2(n10149), .ZN(
        n7732) );
  AOI211_X1 U8936 ( .C1(n10147), .C2(n7734), .A(n7733), .B(n7732), .ZN(n7736)
         );
  NAND2_X1 U8937 ( .A1(n10152), .A2(n7770), .ZN(n7735) );
  OAI211_X1 U8938 ( .C1(n7737), .C2(n10133), .A(n7736), .B(n7735), .ZN(
        P1_U3225) );
  XNOR2_X1 U8939 ( .A(n7738), .B(n7757), .ZN(n7739) );
  NAND2_X1 U8940 ( .A1(n7739), .A2(n11009), .ZN(n7741) );
  AOI22_X1 U8941 ( .A1(n11006), .A2(n5727), .B1(n10174), .B2(n11003), .ZN(
        n7740) );
  NAND2_X1 U8942 ( .A1(n7741), .A2(n7740), .ZN(n10744) );
  MUX2_X1 U8943 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10744), .S(n10869), .Z(n7756) );
  NAND2_X1 U8944 ( .A1(n7742), .A2(n7119), .ZN(n7743) );
  NAND2_X1 U8945 ( .A1(n7743), .A2(n7851), .ZN(n7744) );
  OAI211_X1 U8946 ( .C1(n7119), .C2(n7216), .A(n7744), .B(n7752), .ZN(n7849)
         );
  NAND2_X1 U8947 ( .A1(n7849), .A2(n7850), .ZN(n7747) );
  NAND2_X1 U8948 ( .A1(n7745), .A2(n10724), .ZN(n7746) );
  NAND2_X1 U8949 ( .A1(n7747), .A2(n7746), .ZN(n7758) );
  XNOR2_X1 U8950 ( .A(n7758), .B(n7748), .ZN(n10742) );
  INV_X1 U8951 ( .A(n7749), .ZN(n7750) );
  NAND2_X1 U8952 ( .A1(n11013), .A2(n7750), .ZN(n7751) );
  NAND2_X1 U8953 ( .A1(n10869), .A2(n7751), .ZN(n10442) );
  OR2_X1 U8954 ( .A1(n7752), .A2(n7024), .ZN(n7856) );
  AOI211_X1 U8955 ( .C1(n10738), .C2(n7856), .A(n11085), .B(n7783), .ZN(n10737) );
  NAND2_X1 U8956 ( .A1(n10737), .A2(n10439), .ZN(n7754) );
  AOI22_X1 U8957 ( .A1(n10413), .A2(n10738), .B1(n5745), .B2(n11025), .ZN(
        n7753) );
  OAI211_X1 U8958 ( .C1(n10742), .C2(n10442), .A(n7754), .B(n7753), .ZN(n7755)
         );
  OR2_X1 U8959 ( .A1(n7756), .A2(n7755), .ZN(P1_U3288) );
  INV_X1 U8960 ( .A(n11013), .ZN(n10746) );
  NAND2_X1 U8961 ( .A1(n7758), .A2(n7757), .ZN(n7761) );
  NAND2_X1 U8962 ( .A1(n7852), .A2(n7759), .ZN(n7760) );
  NAND2_X1 U8963 ( .A1(n7761), .A2(n7760), .ZN(n7781) );
  NAND2_X1 U8964 ( .A1(n7781), .A2(n7788), .ZN(n7763) );
  NAND2_X1 U8965 ( .A1(n7772), .A2(n10758), .ZN(n7762) );
  INV_X1 U8966 ( .A(n7767), .ZN(n7765) );
  INV_X1 U8967 ( .A(n7802), .ZN(n7766) );
  AOI21_X1 U8968 ( .B1(n7768), .B2(n7767), .A(n7766), .ZN(n10797) );
  NAND2_X1 U8969 ( .A1(n7783), .A2(n10758), .ZN(n7782) );
  AOI21_X1 U8970 ( .B1(n7782), .B2(n7800), .A(n11085), .ZN(n7769) );
  NAND2_X1 U8971 ( .A1(n7769), .A2(n7811), .ZN(n10793) );
  INV_X1 U8972 ( .A(n7770), .ZN(n7771) );
  OAI22_X1 U8973 ( .A1(n10793), .A2(n10344), .B1(n10865), .B2(n7771), .ZN(
        n7774) );
  XNOR2_X1 U8974 ( .A(n7901), .B(n7764), .ZN(n7773) );
  INV_X1 U8975 ( .A(n11009), .ZN(n10429) );
  OAI222_X1 U8976 ( .A1(n10851), .A2(n10850), .B1(n7773), .B2(n10429), .C1(
        n10849), .C2(n7772), .ZN(n10795) );
  AOI211_X1 U8977 ( .C1(n10746), .C2(n10797), .A(n7774), .B(n10795), .ZN(n7778) );
  INV_X1 U8978 ( .A(n10419), .ZN(n11023) );
  OAI22_X1 U8979 ( .A1(n11029), .A2(n10794), .B1(n7775), .B2(n10869), .ZN(
        n7776) );
  AOI21_X1 U8980 ( .B1(n10797), .B2(n11023), .A(n7776), .ZN(n7777) );
  OAI21_X1 U8981 ( .B1(n7778), .B2(n11027), .A(n7777), .ZN(P1_U3286) );
  INV_X1 U8982 ( .A(n10305), .ZN(n10126) );
  NAND2_X1 U8983 ( .A1(n10126), .A2(P1_U4006), .ZN(n7779) );
  OAI21_X1 U8984 ( .B1(n6882), .B2(P1_U4006), .A(n7779), .ZN(P1_U3582) );
  XNOR2_X1 U8985 ( .A(n7781), .B(n7780), .ZN(n7792) );
  INV_X1 U8986 ( .A(n7792), .ZN(n10761) );
  OAI211_X1 U8987 ( .C1(n7783), .C2(n10758), .A(n7782), .B(n10515), .ZN(n10757) );
  INV_X1 U8988 ( .A(n10439), .ZN(n7860) );
  AOI22_X1 U8989 ( .A1(n10413), .A2(n7785), .B1(n7784), .B2(n11025), .ZN(n7786) );
  OAI21_X1 U8990 ( .B1(n10757), .B2(n7860), .A(n7786), .ZN(n7794) );
  XNOR2_X1 U8991 ( .A(n7787), .B(n7788), .ZN(n7789) );
  NAND2_X1 U8992 ( .A1(n7789), .A2(n11009), .ZN(n7791) );
  AOI22_X1 U8993 ( .A1(n11006), .A2(n10175), .B1(n10173), .B2(n11003), .ZN(
        n7790) );
  OAI211_X1 U8994 ( .C1(n11013), .C2(n7792), .A(n7791), .B(n7790), .ZN(n10759)
         );
  MUX2_X1 U8995 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10759), .S(n10869), .Z(n7793) );
  AOI211_X1 U8996 ( .C1(n10761), .C2(n11023), .A(n7794), .B(n7793), .ZN(n7795)
         );
  INV_X1 U8997 ( .A(n7795), .ZN(P1_U3287) );
  INV_X1 U8998 ( .A(n7796), .ZN(n7799) );
  AOI22_X1 U8999 ( .A1(n9221), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n10010), .ZN(n7797) );
  OAI21_X1 U9000 ( .B1(n7799), .B2(n8693), .A(n7797), .ZN(P2_U3341) );
  AOI22_X1 U9001 ( .A1(n10227), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10537), .ZN(n7798) );
  OAI21_X1 U9002 ( .B1(n7799), .B2(n5033), .A(n7798), .ZN(P1_U3336) );
  NAND2_X1 U9003 ( .A1(n10173), .A2(n7800), .ZN(n7801) );
  INV_X1 U9004 ( .A(n7909), .ZN(n7803) );
  AOI21_X1 U9005 ( .B1(n7806), .B2(n7804), .A(n7803), .ZN(n10824) );
  AOI22_X1 U9006 ( .A1(n11006), .A2(n10173), .B1(n10172), .B2(n11003), .ZN(
        n7809) );
  XOR2_X1 U9007 ( .A(n7806), .B(n7805), .Z(n7807) );
  NAND2_X1 U9008 ( .A1(n7807), .A2(n11009), .ZN(n7808) );
  OAI211_X1 U9009 ( .C1(n10824), .C2(n11013), .A(n7809), .B(n7808), .ZN(n10827) );
  NAND2_X1 U9010 ( .A1(n10827), .A2(n10869), .ZN(n7816) );
  OAI22_X1 U9011 ( .A1(n10869), .A2(n7473), .B1(n7810), .B2(n10865), .ZN(n7814) );
  AND2_X1 U9012 ( .A1(n7811), .A2(n7930), .ZN(n7812) );
  OR2_X1 U9013 ( .A1(n7812), .A2(n10841), .ZN(n10826) );
  INV_X1 U9014 ( .A(n11022), .ZN(n10378) );
  NOR2_X1 U9015 ( .A1(n10826), .A2(n10378), .ZN(n7813) );
  AOI211_X1 U9016 ( .C1(n10413), .C2(n7930), .A(n7814), .B(n7813), .ZN(n7815)
         );
  OAI211_X1 U9017 ( .C1(n10824), .C2(n10419), .A(n7816), .B(n7815), .ZN(
        P1_U3285) );
  NOR2_X1 U9018 ( .A1(n10547), .A2(n7817), .ZN(n8200) );
  NAND3_X1 U9019 ( .A1(n7819), .A2(n8200), .A3(n7818), .ZN(n7821) );
  INV_X1 U9020 ( .A(n8198), .ZN(n7822) );
  INV_X1 U9021 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U9022 ( .A1(n8798), .A2(n8209), .ZN(n8919) );
  XOR2_X1 U9023 ( .A(n8191), .B(n8919), .Z(n8289) );
  OAI21_X1 U9024 ( .B1(n8955), .B2(n8201), .A(n7823), .ZN(n7825) );
  NAND2_X1 U9025 ( .A1(n7825), .A2(n7824), .ZN(n10945) );
  INV_X1 U9026 ( .A(n10948), .ZN(n7826) );
  XNOR2_X1 U9027 ( .A(n8273), .B(n8919), .ZN(n7828) );
  NAND2_X1 U9028 ( .A1(n6947), .A2(n10902), .ZN(n8950) );
  OAI22_X1 U9029 ( .A1(n7827), .A2(n10937), .B1(n8189), .B2(n10939), .ZN(n9048) );
  AOI21_X1 U9030 ( .B1(n7828), .B2(n10942), .A(n9048), .ZN(n8285) );
  NAND2_X1 U9031 ( .A1(n9050), .A2(n10707), .ZN(n7829) );
  AND2_X1 U9032 ( .A1(n8204), .A2(n7829), .ZN(n8282) );
  AOI22_X1 U9033 ( .A1(n8282), .A2(n10892), .B1(n10975), .B2(n9050), .ZN(n7832) );
  OAI211_X1 U9034 ( .C1(n8289), .C2(n11034), .A(n8285), .B(n7832), .ZN(n7836)
         );
  NAND2_X1 U9035 ( .A1(n11082), .A2(n7836), .ZN(n7833) );
  OAI21_X1 U9036 ( .B1(n11082), .B2(n7834), .A(n7833), .ZN(P2_U3454) );
  NAND2_X1 U9037 ( .A1(n11078), .A2(n7836), .ZN(n7837) );
  OAI21_X1 U9038 ( .B1(n11078), .B2(n7275), .A(n7837), .ZN(P2_U3521) );
  OAI21_X1 U9039 ( .B1(n7840), .B2(n7838), .A(n7839), .ZN(n7841) );
  NAND2_X1 U9040 ( .A1(n7841), .A2(n10143), .ZN(n7847) );
  NAND2_X1 U9041 ( .A1(n10152), .A2(n10864), .ZN(n7844) );
  AOI21_X1 U9042 ( .B1(n10147), .B2(n10171), .A(n7842), .ZN(n7843) );
  OAI211_X1 U9043 ( .C1(n10850), .C2(n10149), .A(n7844), .B(n7843), .ZN(n7845)
         );
  INV_X1 U9044 ( .A(n7845), .ZN(n7846) );
  OAI211_X1 U9045 ( .C1(n10863), .C2(n10156), .A(n7847), .B(n7846), .ZN(
        P1_U3211) );
  XNOR2_X1 U9046 ( .A(n7850), .B(n7848), .ZN(n7855) );
  XNOR2_X1 U9047 ( .A(n7850), .B(n7849), .ZN(n10727) );
  OAI22_X1 U9048 ( .A1(n7852), .A2(n10851), .B1(n7851), .B2(n10849), .ZN(n7853) );
  AOI21_X1 U9049 ( .B1(n10727), .B2(n10746), .A(n7853), .ZN(n7854) );
  OAI21_X1 U9050 ( .B1(n10429), .B2(n7855), .A(n7854), .ZN(n10725) );
  INV_X1 U9051 ( .A(n10725), .ZN(n7863) );
  OAI211_X1 U9052 ( .C1(n7857), .C2(n10724), .A(n10515), .B(n7856), .ZN(n10723) );
  AOI22_X1 U9053 ( .A1(n11027), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n11025), .ZN(n7859) );
  NAND2_X1 U9054 ( .A1(n10413), .A2(n7024), .ZN(n7858) );
  OAI211_X1 U9055 ( .C1(n10723), .C2(n7860), .A(n7859), .B(n7858), .ZN(n7861)
         );
  AOI21_X1 U9056 ( .B1(n10727), .B2(n11023), .A(n7861), .ZN(n7862) );
  OAI21_X1 U9057 ( .B1(n7863), .B2(n11027), .A(n7862), .ZN(P1_U3289) );
  INV_X1 U9058 ( .A(n7864), .ZN(n7900) );
  AOI22_X1 U9059 ( .A1(n9232), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n10010), .ZN(n7865) );
  OAI21_X1 U9060 ( .B1(n7900), .B2(n10012), .A(n7865), .ZN(P2_U3340) );
  NOR2_X1 U9061 ( .A1(n7866), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8411) );
  INV_X1 U9062 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7868) );
  MUX2_X1 U9063 ( .A(n7868), .B(P2_REG1_REG_11__SCAN_IN), .S(n7991), .Z(n7869)
         );
  AOI211_X1 U9064 ( .C1(n7870), .C2(n7869), .A(n7982), .B(n10673), .ZN(n7871)
         );
  AOI211_X1 U9065 ( .C1(n10672), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n8411), .B(
        n7871), .ZN(n7879) );
  AOI21_X1 U9066 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7873), .A(n7872), .ZN(
        n7876) );
  NOR2_X1 U9067 ( .A1(n7991), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7874) );
  AOI21_X1 U9068 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n7991), .A(n7874), .ZN(
        n7875) );
  NAND2_X1 U9069 ( .A1(n7876), .A2(n7875), .ZN(n7990) );
  OAI21_X1 U9070 ( .B1(n7876), .B2(n7875), .A(n7990), .ZN(n7877) );
  NAND2_X1 U9071 ( .A1(n7877), .A2(n10651), .ZN(n7878) );
  OAI211_X1 U9072 ( .C1(n10653), .C2(n7880), .A(n7879), .B(n7878), .ZN(
        P2_U3256) );
  NOR2_X1 U9073 ( .A1(n7881), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10178) );
  INV_X1 U9074 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10987) );
  MUX2_X1 U9075 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10987), .S(n10185), .Z(
        n10177) );
  OAI21_X1 U9076 ( .B1(n10179), .B2(n10178), .A(n10177), .ZN(n10196) );
  NAND2_X1 U9077 ( .A1(n7882), .A2(n10987), .ZN(n10194) );
  INV_X1 U9078 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11017) );
  NOR2_X1 U9079 ( .A1(n10201), .A2(n11017), .ZN(n7883) );
  AOI21_X1 U9080 ( .B1(n11017), .B2(n10201), .A(n7883), .ZN(n10195) );
  AOI21_X1 U9081 ( .B1(n10196), .B2(n10194), .A(n10195), .ZN(n10211) );
  NOR2_X1 U9082 ( .A1(n10201), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10210) );
  INV_X1 U9083 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U9084 ( .A1(n10217), .A2(n7885), .ZN(n7884) );
  OAI21_X1 U9085 ( .B1(n10217), .B2(n7885), .A(n7884), .ZN(n10209) );
  OAI21_X1 U9086 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(n10208) );
  OAI21_X1 U9087 ( .B1(n10217), .B2(P1_REG1_REG_14__SCAN_IN), .A(n10208), .ZN(
        n8052) );
  XOR2_X1 U9088 ( .A(n8061), .B(n8052), .Z(n8055) );
  XNOR2_X1 U9089 ( .A(n8055), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n7897) );
  INV_X1 U9090 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7887) );
  AND2_X1 U9091 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10145) );
  AOI21_X1 U9092 ( .B1(n10692), .B2(n8061), .A(n10145), .ZN(n7886) );
  OAI21_X1 U9093 ( .B1(n7887), .B2(n10631), .A(n7886), .ZN(n7896) );
  XNOR2_X1 U9094 ( .A(n10185), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U9095 ( .A1(n10185), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7888) );
  NAND2_X1 U9096 ( .A1(n10188), .A2(n7888), .ZN(n10204) );
  INV_X1 U9097 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7889) );
  XNOR2_X1 U9098 ( .A(n10201), .B(n7889), .ZN(n10203) );
  NAND2_X1 U9099 ( .A1(n10204), .A2(n10203), .ZN(n10202) );
  NAND2_X1 U9100 ( .A1(n10201), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U9101 ( .A1(n10202), .A2(n7890), .ZN(n10220) );
  OR2_X1 U9102 ( .A1(n10217), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U9103 ( .A1(n10217), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7892) );
  AND2_X1 U9104 ( .A1(n7891), .A2(n7892), .ZN(n10219) );
  NAND2_X1 U9105 ( .A1(n10220), .A2(n10219), .ZN(n10218) );
  NAND2_X1 U9106 ( .A1(n10218), .A2(n7892), .ZN(n8060) );
  XNOR2_X1 U9107 ( .A(n8060), .B(n8061), .ZN(n7894) );
  INV_X1 U9108 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7893) );
  NOR2_X1 U9109 ( .A1(n7894), .A2(n7893), .ZN(n8059) );
  AOI211_X1 U9110 ( .C1(n7894), .C2(n7893), .A(n10248), .B(n8059), .ZN(n7895)
         );
  AOI211_X1 U9111 ( .C1(n7897), .C2(n10635), .A(n7896), .B(n7895), .ZN(n7898)
         );
  INV_X1 U9112 ( .A(n7898), .ZN(P1_U3256) );
  INV_X1 U9113 ( .A(n10244), .ZN(n10239) );
  OAI222_X1 U9114 ( .A1(n10239), .A2(P1_U3084), .B1(n5033), .B2(n7900), .C1(
        n9004), .C2(n7899), .ZN(P1_U3335) );
  INV_X1 U9115 ( .A(n7901), .ZN(n7902) );
  NAND2_X1 U9116 ( .A1(n7902), .A2(n5123), .ZN(n10845) );
  XOR2_X1 U9117 ( .A(n8079), .B(n8080), .Z(n7907) );
  OAI222_X1 U9118 ( .A1(n10851), .A2(n8226), .B1(n10849), .B2(n10852), .C1(
        n10429), .C2(n7907), .ZN(n10916) );
  INV_X1 U9119 ( .A(n10916), .ZN(n7919) );
  NAND2_X1 U9120 ( .A1(n10850), .A2(n10825), .ZN(n7908) );
  INV_X1 U9121 ( .A(n10848), .ZN(n7912) );
  NOR2_X1 U9122 ( .A1(n7910), .A2(n10172), .ZN(n7911) );
  NAND2_X1 U9123 ( .A1(n7933), .A2(n7932), .ZN(n8154) );
  NAND2_X1 U9124 ( .A1(n8133), .A2(n10171), .ZN(n8073) );
  NAND2_X1 U9125 ( .A1(n8154), .A2(n8073), .ZN(n7913) );
  XNOR2_X1 U9126 ( .A(n7913), .B(n8079), .ZN(n10918) );
  INV_X1 U9127 ( .A(n10442), .ZN(n8632) );
  NAND2_X1 U9128 ( .A1(n10843), .A2(n10882), .ZN(n7942) );
  INV_X1 U9129 ( .A(n7942), .ZN(n7914) );
  INV_X1 U9130 ( .A(n8076), .ZN(n10914) );
  OAI21_X1 U9131 ( .B1(n7914), .B2(n10914), .A(n8165), .ZN(n10915) );
  AOI22_X1 U9132 ( .A1(n11027), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8022), .B2(
        n11025), .ZN(n7916) );
  NAND2_X1 U9133 ( .A1(n10413), .A2(n8076), .ZN(n7915) );
  OAI211_X1 U9134 ( .C1(n10915), .C2(n10378), .A(n7916), .B(n7915), .ZN(n7917)
         );
  AOI21_X1 U9135 ( .B1(n10918), .B2(n8632), .A(n7917), .ZN(n7918) );
  OAI21_X1 U9136 ( .B1(n7919), .B2(n11027), .A(n7918), .ZN(P1_U3282) );
  NAND2_X1 U9137 ( .A1(n10152), .A2(n7920), .ZN(n7923) );
  INV_X1 U9138 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7921) );
  NOR2_X1 U9139 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7921), .ZN(n10596) );
  AOI21_X1 U9140 ( .B1(n10147), .B2(n10172), .A(n10596), .ZN(n7922) );
  OAI211_X1 U9141 ( .C1(n7924), .C2(n10149), .A(n7923), .B(n7922), .ZN(n7929)
         );
  XOR2_X1 U9142 ( .A(n7925), .B(n7926), .Z(n7927) );
  NOR2_X1 U9143 ( .A1(n7927), .A2(n10133), .ZN(n7928) );
  AOI211_X1 U9144 ( .C1(n7930), .C2(n10131), .A(n7929), .B(n7928), .ZN(n7931)
         );
  INV_X1 U9145 ( .A(n7931), .ZN(P1_U3237) );
  OR2_X1 U9146 ( .A1(n7933), .A2(n7932), .ZN(n7934) );
  NAND2_X1 U9147 ( .A1(n8154), .A2(n7934), .ZN(n7940) );
  AOI22_X1 U9148 ( .A1(n11006), .A2(n10172), .B1(n10170), .B2(n11003), .ZN(
        n7939) );
  XNOR2_X1 U9149 ( .A(n7936), .B(n7935), .ZN(n7937) );
  NAND2_X1 U9150 ( .A1(n7937), .A2(n11009), .ZN(n7938) );
  OAI211_X1 U9151 ( .C1(n7940), .C2(n11013), .A(n7939), .B(n7938), .ZN(n10884)
         );
  INV_X1 U9152 ( .A(n10884), .ZN(n7947) );
  INV_X1 U9153 ( .A(n7940), .ZN(n10886) );
  OR2_X1 U9154 ( .A1(n10843), .A2(n10882), .ZN(n7941) );
  NAND2_X1 U9155 ( .A1(n7942), .A2(n7941), .ZN(n10883) );
  AOI22_X1 U9156 ( .A1(n11027), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8121), .B2(
        n11025), .ZN(n7944) );
  NAND2_X1 U9157 ( .A1(n10413), .A2(n8133), .ZN(n7943) );
  OAI211_X1 U9158 ( .C1(n10883), .C2(n10378), .A(n7944), .B(n7943), .ZN(n7945)
         );
  AOI21_X1 U9159 ( .B1(n10886), .B2(n11023), .A(n7945), .ZN(n7946) );
  OAI21_X1 U9160 ( .B1(n7947), .B2(n11027), .A(n7946), .ZN(P1_U3283) );
  AOI21_X1 U9161 ( .B1(n7949), .B2(n7948), .A(n9086), .ZN(n7950) );
  NAND2_X1 U9162 ( .A1(n7950), .A2(n9038), .ZN(n7955) );
  OAI22_X1 U9163 ( .A1(n9127), .A2(n8448), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7951), .ZN(n7953) );
  INV_X1 U9164 ( .A(n10873), .ZN(n8820) );
  OAI22_X1 U9165 ( .A1(n9146), .A2(n8820), .B1(n9104), .B2(n8449), .ZN(n7952)
         );
  AOI211_X1 U9166 ( .C1(n8452), .C2(n9129), .A(n7953), .B(n7952), .ZN(n7954)
         );
  NAND2_X1 U9167 ( .A1(n7955), .A2(n7954), .ZN(P2_U3215) );
  INV_X1 U9168 ( .A(n7956), .ZN(n7958) );
  OAI222_X1 U9169 ( .A1(n9004), .A2(n9736), .B1(n5033), .B2(n7958), .C1(
        P1_U3084), .C2(n10392), .ZN(P1_U3334) );
  OAI222_X1 U9170 ( .A1(n9846), .A2(P2_U3152), .B1(n8693), .B2(n7958), .C1(
        n7957), .C2(n10005), .ZN(P2_U3339) );
  INV_X1 U9171 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8277) );
  NOR2_X1 U9172 ( .A1(n9049), .A2(P2_U3152), .ZN(n7963) );
  INV_X1 U9173 ( .A(n9122), .ZN(n9093) );
  NAND2_X1 U9174 ( .A1(n9161), .A2(n7959), .ZN(n8793) );
  INV_X1 U9175 ( .A(n8793), .ZN(n8274) );
  INV_X1 U9176 ( .A(n9127), .ZN(n8739) );
  AOI22_X1 U9177 ( .A1(n9093), .A2(n8274), .B1(n8739), .B2(n9159), .ZN(n7962)
         );
  OAI21_X1 U9178 ( .B1(n7959), .B2(n8780), .A(n8273), .ZN(n7960) );
  AOI22_X1 U9179 ( .A1(n10707), .A2(n9098), .B1(n9135), .B2(n7960), .ZN(n7961)
         );
  OAI211_X1 U9180 ( .C1(n8277), .C2(n7963), .A(n7962), .B(n7961), .ZN(P2_U3234) );
  AOI22_X1 U9181 ( .A1(n9892), .A2(n8248), .B1(n9157), .B2(n9890), .ZN(n10810)
         );
  OAI22_X1 U9182 ( .A1(n10810), .A2(n9080), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9694), .ZN(n7965) );
  NOR2_X1 U9183 ( .A1(n9146), .A2(n10817), .ZN(n7964) );
  AOI211_X1 U9184 ( .C1(n9129), .C2(n10805), .A(n7965), .B(n7964), .ZN(n7970)
         );
  OAI22_X1 U9185 ( .A1(n8326), .A2(n9122), .B1(n9086), .B2(n7967), .ZN(n7968)
         );
  NAND3_X1 U9186 ( .A1(n8028), .A2(n5413), .A3(n7968), .ZN(n7969) );
  OAI211_X1 U9187 ( .C1(n7976), .C2(n9086), .A(n7970), .B(n7969), .ZN(P2_U3229) );
  OAI21_X1 U9188 ( .B1(n9146), .B2(n8251), .A(n7971), .ZN(n7973) );
  INV_X1 U9189 ( .A(n9891), .ZN(n9042) );
  OAI22_X1 U9190 ( .A1(n9042), .A2(n9127), .B1(n9104), .B2(n8250), .ZN(n7972)
         );
  AOI211_X1 U9191 ( .C1(n9896), .C2(n9129), .A(n7973), .B(n7972), .ZN(n7978)
         );
  OAI22_X1 U9192 ( .A1(n8250), .A2(n9122), .B1(n9086), .B2(n7974), .ZN(n7975)
         );
  NAND3_X1 U9193 ( .A1(n7976), .A2(n5126), .A3(n7975), .ZN(n7977) );
  OAI211_X1 U9194 ( .C1(n7979), .C2(n9086), .A(n7978), .B(n7977), .ZN(P2_U3241) );
  INV_X1 U9195 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7980) );
  MUX2_X1 U9196 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n7980), .S(n8110), .Z(n7984)
         );
  INV_X1 U9197 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7981) );
  MUX2_X1 U9198 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7981), .S(n8015), .Z(n8006)
         );
  OAI21_X1 U9199 ( .B1(n8015), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8005), .ZN(
        n7983) );
  NAND2_X1 U9200 ( .A1(n7984), .A2(n7983), .ZN(n8104) );
  OAI21_X1 U9201 ( .B1(n7984), .B2(n7983), .A(n8104), .ZN(n7986) );
  INV_X1 U9202 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U9203 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8711) );
  OAI21_X1 U9204 ( .B1(n9217), .B2(n8368), .A(n8711), .ZN(n7985) );
  AOI21_X1 U9205 ( .B1(n10649), .B2(n7986), .A(n7985), .ZN(n7996) );
  INV_X1 U9206 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7987) );
  MUX2_X1 U9207 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n7987), .S(n8110), .Z(n7993)
         );
  INV_X1 U9208 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7988) );
  MUX2_X1 U9209 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7988), .S(n8015), .Z(n7989)
         );
  INV_X1 U9210 ( .A(n7989), .ZN(n8011) );
  OAI21_X1 U9211 ( .B1(n7991), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7990), .ZN(
        n8012) );
  NOR2_X1 U9212 ( .A1(n8011), .A2(n8012), .ZN(n8010) );
  AOI21_X1 U9213 ( .B1(n8015), .B2(P2_REG2_REG_12__SCAN_IN), .A(n8010), .ZN(
        n7992) );
  NAND2_X1 U9214 ( .A1(n7992), .A2(n7993), .ZN(n8111) );
  OAI21_X1 U9215 ( .B1(n7993), .B2(n7992), .A(n8111), .ZN(n7994) );
  NAND2_X1 U9216 ( .A1(n10651), .A2(n7994), .ZN(n7995) );
  OAI211_X1 U9217 ( .C1(n10653), .C2(n7997), .A(n7996), .B(n7995), .ZN(
        P2_U3258) );
  INV_X1 U9218 ( .A(n8045), .ZN(n7998) );
  AOI211_X1 U9219 ( .C1(n8000), .C2(n7999), .A(n9086), .B(n7998), .ZN(n8004)
         );
  INV_X1 U9220 ( .A(n8240), .ZN(n8242) );
  AOI22_X1 U9221 ( .A1(n8739), .A2(n8242), .B1(n8188), .B2(n9098), .ZN(n8002)
         );
  AND2_X1 U9222 ( .A1(P2_U3152), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n10671) );
  AOI21_X1 U9223 ( .B1(n9049), .B2(P2_REG3_REG_2__SCAN_IN), .A(n10671), .ZN(
        n8001) );
  OAI211_X1 U9224 ( .C1(n8194), .C2(n9104), .A(n8002), .B(n8001), .ZN(n8003)
         );
  OR2_X1 U9225 ( .A1(n8004), .A2(n8003), .ZN(P2_U3239) );
  INV_X1 U9226 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8365) );
  OAI21_X1 U9227 ( .B1(n8007), .B2(n8006), .A(n8005), .ZN(n8008) );
  NAND2_X1 U9228 ( .A1(n10649), .A2(n8008), .ZN(n8009) );
  NAND2_X1 U9229 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n8484) );
  OAI211_X1 U9230 ( .C1(n8365), .C2(n9217), .A(n8009), .B(n8484), .ZN(n8014)
         );
  AOI211_X1 U9231 ( .C1(n8012), .C2(n8011), .A(n8010), .B(n10677), .ZN(n8013)
         );
  AOI211_X1 U9232 ( .C1(n10684), .C2(n8015), .A(n8014), .B(n8013), .ZN(n8016)
         );
  INV_X1 U9233 ( .A(n8016), .ZN(P2_U3257) );
  XOR2_X1 U9234 ( .A(n8017), .B(n8018), .Z(n8025) );
  NAND2_X1 U9235 ( .A1(n10115), .A2(n10171), .ZN(n8020) );
  OAI211_X1 U9236 ( .C1(n8226), .C2(n10118), .A(n8020), .B(n8019), .ZN(n8021)
         );
  AOI21_X1 U9237 ( .B1(n8022), .B2(n10152), .A(n8021), .ZN(n8024) );
  NAND2_X1 U9238 ( .A1(n8076), .A2(n10131), .ZN(n8023) );
  OAI211_X1 U9239 ( .C1(n8025), .C2(n10133), .A(n8024), .B(n8023), .ZN(
        P1_U3229) );
  INV_X1 U9240 ( .A(n8026), .ZN(n8034) );
  OAI21_X1 U9241 ( .B1(n8034), .B2(n8027), .A(n8028), .ZN(n8037) );
  INV_X1 U9242 ( .A(n9080), .ZN(n9143) );
  OR2_X1 U9243 ( .A1(n8250), .A2(n10939), .ZN(n8030) );
  OR2_X1 U9244 ( .A1(n8240), .A2(n10937), .ZN(n8029) );
  NAND2_X1 U9245 ( .A1(n8030), .A2(n8029), .ZN(n10774) );
  AOI22_X1 U9246 ( .A1(n9143), .A2(n10774), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n8032) );
  NAND2_X1 U9247 ( .A1(n9129), .A2(n10786), .ZN(n8031) );
  OAI211_X1 U9248 ( .C1(n8247), .C2(n9146), .A(n8032), .B(n8031), .ZN(n8036)
         );
  NOR4_X1 U9249 ( .A1(n9122), .A2(n8034), .A3(n8240), .A4(n8033), .ZN(n8035)
         );
  AOI211_X1 U9250 ( .C1(n8037), .C2(n9135), .A(n8036), .B(n8035), .ZN(n8038)
         );
  INV_X1 U9251 ( .A(n8038), .ZN(P2_U3232) );
  INV_X1 U9252 ( .A(n8039), .ZN(n8150) );
  OAI222_X1 U9253 ( .A1(n5033), .A2(n8150), .B1(n8040), .B2(P1_U3084), .C1(
        n9737), .C2(n9004), .ZN(P1_U3333) );
  INV_X1 U9254 ( .A(n9104), .ZN(n9125) );
  MUX2_X1 U9255 ( .A(n9129), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n8042) );
  OAI22_X1 U9256 ( .A1(n9146), .A2(n8241), .B1(n9127), .B2(n8326), .ZN(n8041)
         );
  AOI211_X1 U9257 ( .C1(n9125), .C2(n9158), .A(n8042), .B(n8041), .ZN(n8051)
         );
  INV_X1 U9258 ( .A(n8043), .ZN(n8044) );
  AOI21_X1 U9259 ( .B1(n8045), .B2(n8044), .A(n9086), .ZN(n8049) );
  INV_X1 U9260 ( .A(n8046), .ZN(n8047) );
  NOR3_X1 U9261 ( .A1(n9122), .A2(n8189), .A3(n8047), .ZN(n8048) );
  OAI21_X1 U9262 ( .B1(n8049), .B2(n8048), .A(n8027), .ZN(n8050) );
  NAND2_X1 U9263 ( .A1(n8051), .A2(n8050), .ZN(P2_U3220) );
  INV_X1 U9264 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8054) );
  OAI22_X1 U9265 ( .A1(n8055), .A2(n8054), .B1(n8053), .B2(n8052), .ZN(n8058)
         );
  NOR2_X1 U9266 ( .A1(n8499), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8056) );
  AOI21_X1 U9267 ( .B1(n8499), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8056), .ZN(
        n8057) );
  NAND2_X1 U9268 ( .A1(n8057), .A2(n8058), .ZN(n8500) );
  OAI211_X1 U9269 ( .C1(n8058), .C2(n8057), .A(n10635), .B(n8500), .ZN(n8071)
         );
  AOI21_X1 U9270 ( .B1(n8061), .B2(n8060), .A(n8059), .ZN(n8064) );
  NAND2_X1 U9271 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8499), .ZN(n8062) );
  OAI21_X1 U9272 ( .B1(n8499), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8062), .ZN(
        n8063) );
  NOR2_X1 U9273 ( .A1(n8064), .A2(n8063), .ZN(n8493) );
  AOI211_X1 U9274 ( .C1(n8064), .C2(n8063), .A(n8493), .B(n10248), .ZN(n8069)
         );
  INV_X1 U9275 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n8376) );
  NOR2_X1 U9276 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8065), .ZN(n8066) );
  AOI21_X1 U9277 ( .B1(n10692), .B2(n8499), .A(n8066), .ZN(n8067) );
  OAI21_X1 U9278 ( .B1(n8376), .B2(n10631), .A(n8067), .ZN(n8068) );
  NOR2_X1 U9279 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  NAND2_X1 U9280 ( .A1(n8071), .A2(n8070), .ZN(P1_U3257) );
  NAND2_X1 U9281 ( .A1(n8076), .A2(n10170), .ZN(n8072) );
  AND2_X1 U9282 ( .A1(n8073), .A2(n8072), .ZN(n8153) );
  INV_X1 U9283 ( .A(n8160), .ZN(n8074) );
  AND2_X1 U9284 ( .A1(n8153), .A2(n8074), .ZN(n8075) );
  NAND2_X1 U9285 ( .A1(n8154), .A2(n8075), .ZN(n8158) );
  OR2_X1 U9286 ( .A1(n8475), .A2(n10169), .ZN(n8077) );
  OR2_X1 U9287 ( .A1(n8076), .A2(n10170), .ZN(n8155) );
  OR2_X1 U9288 ( .A1(n8160), .A2(n8155), .ZN(n8157) );
  AND2_X1 U9289 ( .A1(n8077), .A2(n8157), .ZN(n8078) );
  XNOR2_X1 U9290 ( .A(n8171), .B(n8084), .ZN(n8092) );
  AOI22_X1 U9291 ( .A1(n11006), .A2(n10169), .B1(n11005), .B2(n11003), .ZN(
        n8091) );
  NAND2_X1 U9292 ( .A1(n8080), .A2(n8079), .ZN(n8082) );
  NAND2_X1 U9293 ( .A1(n8082), .A2(n8081), .ZN(n8152) );
  NAND2_X1 U9294 ( .A1(n8152), .A2(n8160), .ZN(n8151) );
  INV_X1 U9295 ( .A(n8151), .ZN(n8083) );
  NOR3_X1 U9296 ( .A1(n8083), .A2(n5393), .A3(n8084), .ZN(n8089) );
  AND2_X1 U9297 ( .A1(n8160), .A2(n8084), .ZN(n8088) );
  OAI21_X1 U9298 ( .B1(n8089), .B2(n5052), .A(n11009), .ZN(n8090) );
  OAI211_X1 U9299 ( .C1(n8092), .C2(n11013), .A(n8091), .B(n8090), .ZN(n10967)
         );
  INV_X1 U9300 ( .A(n10967), .ZN(n8099) );
  INV_X1 U9301 ( .A(n8092), .ZN(n10969) );
  NOR2_X1 U9302 ( .A1(n8164), .A2(n10965), .ZN(n8093) );
  OR2_X1 U9303 ( .A1(n8181), .A2(n8093), .ZN(n10966) );
  AOI22_X1 U9304 ( .A1(n11027), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8228), .B2(
        n11025), .ZN(n8096) );
  NAND2_X1 U9305 ( .A1(n8094), .A2(n10413), .ZN(n8095) );
  OAI211_X1 U9306 ( .C1(n10966), .C2(n10378), .A(n8096), .B(n8095), .ZN(n8097)
         );
  AOI21_X1 U9307 ( .B1(n10969), .B2(n11023), .A(n8097), .ZN(n8098) );
  OAI21_X1 U9308 ( .B1(n8099), .B2(n11027), .A(n8098), .ZN(P1_U3280) );
  INV_X1 U9309 ( .A(n8100), .ZN(n8120) );
  OAI222_X1 U9310 ( .A1(n5033), .A2(n8120), .B1(n8102), .B2(P1_U3084), .C1(
        n8101), .C2(n9004), .ZN(P1_U3332) );
  INV_X1 U9311 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8103) );
  MUX2_X1 U9312 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8103), .S(n9170), .Z(n8106)
         );
  OAI21_X1 U9313 ( .B1(n8110), .B2(P2_REG1_REG_13__SCAN_IN), .A(n8104), .ZN(
        n8105) );
  NAND2_X1 U9314 ( .A1(n8106), .A2(n8105), .ZN(n9164) );
  OAI21_X1 U9315 ( .B1(n8106), .B2(n8105), .A(n9164), .ZN(n8108) );
  INV_X1 U9316 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U9317 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8740) );
  OAI21_X1 U9318 ( .B1(n9217), .B2(n8371), .A(n8740), .ZN(n8107) );
  AOI21_X1 U9319 ( .B1(n10649), .B2(n8108), .A(n8107), .ZN(n8117) );
  INV_X1 U9320 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8109) );
  MUX2_X1 U9321 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n8109), .S(n9170), .Z(n8114)
         );
  OR2_X1 U9322 ( .A1(n8110), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U9323 ( .A1(n8112), .A2(n8111), .ZN(n8113) );
  NAND2_X1 U9324 ( .A1(n8114), .A2(n8113), .ZN(n9169) );
  OAI21_X1 U9325 ( .B1(n8114), .B2(n8113), .A(n9169), .ZN(n8115) );
  NAND2_X1 U9326 ( .A1(n10651), .A2(n8115), .ZN(n8116) );
  OAI211_X1 U9327 ( .C1(n10653), .C2(n8118), .A(n8117), .B(n8116), .ZN(
        P2_U3259) );
  OAI222_X1 U9328 ( .A1(P2_U3152), .A2(n8201), .B1(n8693), .B2(n8120), .C1(
        n8119), .C2(n10005), .ZN(P2_U3337) );
  NAND2_X1 U9329 ( .A1(n10152), .A2(n8121), .ZN(n8124) );
  AOI21_X1 U9330 ( .B1(n10147), .B2(n10170), .A(n8122), .ZN(n8123) );
  OAI211_X1 U9331 ( .C1(n8125), .C2(n10149), .A(n8124), .B(n8123), .ZN(n8132)
         );
  NAND2_X1 U9332 ( .A1(n8127), .A2(n8126), .ZN(n8128) );
  XOR2_X1 U9333 ( .A(n8129), .B(n8128), .Z(n8130) );
  NOR2_X1 U9334 ( .A1(n8130), .A2(n10133), .ZN(n8131) );
  AOI211_X1 U9335 ( .C1(n8133), .C2(n10131), .A(n8132), .B(n8131), .ZN(n8134)
         );
  INV_X1 U9336 ( .A(n8134), .ZN(P1_U3219) );
  INV_X1 U9337 ( .A(n8135), .ZN(n8138) );
  NOR3_X1 U9338 ( .A1(n9122), .A2(n8448), .A3(n8136), .ZN(n8137) );
  AOI21_X1 U9339 ( .B1(n8138), .B2(n9135), .A(n8137), .ZN(n8148) );
  INV_X1 U9340 ( .A(n8139), .ZN(n8145) );
  INV_X1 U9341 ( .A(n8418), .ZN(n9154) );
  AOI22_X1 U9342 ( .A1(n8739), .A2(n9154), .B1(n9129), .B2(n8267), .ZN(n8143)
         );
  NAND2_X1 U9343 ( .A1(n9098), .A2(n8423), .ZN(n8141) );
  INV_X1 U9344 ( .A(n8448), .ZN(n9156) );
  NAND2_X1 U9345 ( .A1(n9125), .A2(n9156), .ZN(n8140) );
  NAND4_X1 U9346 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n8144)
         );
  AOI21_X1 U9347 ( .B1(n8145), .B2(n9135), .A(n8144), .ZN(n8146) );
  OAI21_X1 U9348 ( .B1(n8148), .B2(n8147), .A(n8146), .ZN(P2_U3233) );
  OAI222_X1 U9349 ( .A1(P2_U3152), .A2(n6488), .B1(n8693), .B2(n8150), .C1(
        n8149), .C2(n10005), .ZN(P2_U3338) );
  OAI21_X1 U9350 ( .B1(n8160), .B2(n8152), .A(n8151), .ZN(n8163) );
  OAI22_X1 U9351 ( .A1(n8309), .A2(n10851), .B1(n8467), .B2(n10849), .ZN(n8162) );
  NAND2_X1 U9352 ( .A1(n8154), .A2(n8153), .ZN(n8156) );
  AND2_X1 U9353 ( .A1(n8156), .A2(n8155), .ZN(n8159) );
  AOI21_X1 U9354 ( .B1(n8160), .B2(n8159), .A(n5115), .ZN(n8316) );
  NOR2_X1 U9355 ( .A1(n8316), .A2(n11013), .ZN(n8161) );
  AOI211_X1 U9356 ( .C1(n11009), .C2(n8163), .A(n8162), .B(n8161), .ZN(n8315)
         );
  AOI21_X1 U9357 ( .B1(n8475), .B2(n8165), .A(n8164), .ZN(n8313) );
  INV_X1 U9358 ( .A(n8475), .ZN(n8167) );
  AOI22_X1 U9359 ( .A1(n11027), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8463), .B2(
        n11025), .ZN(n8166) );
  OAI21_X1 U9360 ( .B1(n8167), .B2(n11029), .A(n8166), .ZN(n8169) );
  NOR2_X1 U9361 ( .A1(n8316), .A2(n10419), .ZN(n8168) );
  AOI211_X1 U9362 ( .C1(n8313), .C2(n11022), .A(n8169), .B(n8168), .ZN(n8170)
         );
  OAI21_X1 U9363 ( .B1(n8315), .B2(n11027), .A(n8170), .ZN(P1_U3281) );
  NAND2_X1 U9364 ( .A1(n8172), .A2(n8176), .ZN(n8173) );
  NAND2_X1 U9365 ( .A1(n8387), .A2(n8173), .ZN(n8180) );
  OAI21_X1 U9366 ( .B1(n8176), .B2(n8175), .A(n8390), .ZN(n8178) );
  OAI22_X1 U9367 ( .A1(n8662), .A2(n10851), .B1(n8309), .B2(n10849), .ZN(n8177) );
  AOI21_X1 U9368 ( .B1(n8178), .B2(n11009), .A(n8177), .ZN(n8179) );
  OAI21_X1 U9369 ( .B1(n8180), .B2(n11013), .A(n8179), .ZN(n10984) );
  INV_X1 U9370 ( .A(n10984), .ZN(n8187) );
  INV_X1 U9371 ( .A(n8180), .ZN(n10986) );
  INV_X1 U9372 ( .A(n8385), .ZN(n10982) );
  OR2_X1 U9373 ( .A1(n8181), .A2(n10982), .ZN(n8182) );
  NAND2_X1 U9374 ( .A1(n11000), .A2(n8182), .ZN(n10983) );
  AOI22_X1 U9375 ( .A1(n11027), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8305), .B2(
        n11025), .ZN(n8184) );
  NAND2_X1 U9376 ( .A1(n8385), .A2(n10413), .ZN(n8183) );
  OAI211_X1 U9377 ( .C1(n10983), .C2(n10378), .A(n8184), .B(n8183), .ZN(n8185)
         );
  AOI21_X1 U9378 ( .B1(n10986), .B2(n11023), .A(n8185), .ZN(n8186) );
  OAI21_X1 U9379 ( .B1(n8187), .B2(n11027), .A(n8186), .ZN(P1_U3279) );
  NAND2_X1 U9380 ( .A1(n8189), .A2(n8188), .ZN(n8256) );
  NAND2_X1 U9381 ( .A1(n9158), .A2(n8190), .ZN(n8800) );
  NAND2_X1 U9382 ( .A1(n9159), .A2(n9050), .ZN(n8192) );
  NAND2_X1 U9383 ( .A1(n8192), .A2(n8191), .ZN(n8196) );
  NAND2_X1 U9384 ( .A1(n8194), .A2(n8193), .ZN(n8195) );
  XNOR2_X1 U9385 ( .A(n8920), .B(n8238), .ZN(n10733) );
  INV_X1 U9386 ( .A(n10733), .ZN(n8219) );
  NOR2_X1 U9387 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  NAND2_X1 U9388 ( .A1(n8200), .A2(n8199), .ZN(n8203) );
  NAND2_X1 U9389 ( .A1(n8786), .A2(n6488), .ZN(n8276) );
  INV_X1 U9390 ( .A(n8276), .ZN(n8202) );
  NAND2_X1 U9391 ( .A1(n10957), .A2(n8202), .ZN(n10953) );
  OR2_X1 U9392 ( .A1(n8204), .A2(n8188), .ZN(n10770) );
  NAND2_X1 U9393 ( .A1(n8204), .A2(n8188), .ZN(n8205) );
  NAND2_X1 U9394 ( .A1(n10770), .A2(n8205), .ZN(n10730) );
  INV_X1 U9395 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8206) );
  OAI22_X1 U9396 ( .A1(n10952), .A2(n10730), .B1(n8206), .B2(n9849), .ZN(n8208) );
  NOR2_X1 U9397 ( .A1(n10956), .A2(n8190), .ZN(n8207) );
  AOI211_X1 U9398 ( .C1(n10906), .C2(P2_REG2_REG_2__SCAN_IN), .A(n8208), .B(
        n8207), .ZN(n8218) );
  NAND2_X1 U9399 ( .A1(n8273), .A2(n8798), .ZN(n8210) );
  NAND2_X1 U9400 ( .A1(n8210), .A2(n8209), .ZN(n8212) );
  AOI21_X1 U9401 ( .B1(n8920), .B2(n8212), .A(n8211), .ZN(n8216) );
  AOI22_X1 U9402 ( .A1(n8242), .A2(n9890), .B1(n9892), .B2(n9159), .ZN(n8215)
         );
  INV_X1 U9403 ( .A(n10945), .ZN(n8213) );
  NAND2_X1 U9404 ( .A1(n10733), .A2(n8213), .ZN(n8214) );
  OAI211_X1 U9405 ( .C1(n8216), .C2(n10811), .A(n8215), .B(n8214), .ZN(n10731)
         );
  NAND2_X1 U9406 ( .A1(n10731), .A2(n10957), .ZN(n8217) );
  OAI211_X1 U9407 ( .C1(n8219), .C2(n10953), .A(n8218), .B(n8217), .ZN(
        P2_U3294) );
  OAI211_X1 U9408 ( .C1(n8221), .C2(n8223), .A(n8222), .B(n10143), .ZN(n8230)
         );
  AOI21_X1 U9409 ( .B1(n10147), .B2(n11005), .A(n8224), .ZN(n8225) );
  OAI21_X1 U9410 ( .B1(n8226), .B2(n10149), .A(n8225), .ZN(n8227) );
  AOI21_X1 U9411 ( .B1(n8228), .B2(n10152), .A(n8227), .ZN(n8229) );
  OAI211_X1 U9412 ( .C1(n10965), .C2(n10156), .A(n8230), .B(n8229), .ZN(
        P1_U3234) );
  AOI21_X1 U9413 ( .B1(n8232), .B2(n8231), .A(n9086), .ZN(n8233) );
  NAND2_X1 U9414 ( .A1(n8233), .A2(n8403), .ZN(n8237) );
  NOR2_X1 U9415 ( .A1(n9104), .A2(n10938), .ZN(n8235) );
  OAI22_X1 U9416 ( .A1(n9127), .A2(n10940), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9672), .ZN(n8234) );
  AOI211_X1 U9417 ( .C1(n9129), .C2(n10961), .A(n8235), .B(n8234), .ZN(n8236)
         );
  OAI211_X1 U9418 ( .C1(n5353), .C2(n9146), .A(n8237), .B(n8236), .ZN(P2_U3219) );
  NAND2_X1 U9419 ( .A1(n8423), .A2(n10938), .ZN(n8829) );
  NAND2_X1 U9420 ( .A1(n8920), .A2(n8238), .ZN(n8322) );
  NAND2_X1 U9421 ( .A1(n8240), .A2(n8241), .ZN(n8244) );
  AND2_X1 U9422 ( .A1(n8323), .A2(n8244), .ZN(n8239) );
  NAND2_X1 U9423 ( .A1(n8322), .A2(n8239), .ZN(n8246) );
  NAND2_X1 U9424 ( .A1(n8240), .A2(n8331), .ZN(n8804) );
  NAND2_X1 U9425 ( .A1(n8242), .A2(n8241), .ZN(n8805) );
  NAND2_X1 U9426 ( .A1(n8804), .A2(n8805), .ZN(n8921) );
  INV_X1 U9427 ( .A(n8921), .ZN(n8243) );
  NAND2_X1 U9428 ( .A1(n8244), .A2(n8243), .ZN(n8245) );
  NAND2_X1 U9429 ( .A1(n8246), .A2(n8245), .ZN(n10764) );
  NAND2_X1 U9430 ( .A1(n8326), .A2(n10769), .ZN(n8809) );
  NAND2_X1 U9431 ( .A1(n8248), .A2(n10769), .ZN(n8249) );
  NAND2_X1 U9432 ( .A1(n8250), .A2(n10804), .ZN(n8815) );
  NAND2_X1 U9433 ( .A1(n8449), .A2(n10832), .ZN(n8816) );
  NAND2_X1 U9434 ( .A1(n9157), .A2(n8251), .ZN(n8818) );
  NAND2_X1 U9435 ( .A1(n8253), .A2(n8252), .ZN(n9898) );
  NAND2_X1 U9436 ( .A1(n9157), .A2(n10832), .ZN(n8254) );
  NAND2_X1 U9437 ( .A1(n9042), .A2(n8820), .ZN(n8255) );
  NAND2_X1 U9438 ( .A1(n8448), .A2(n10898), .ZN(n8824) );
  INV_X1 U9439 ( .A(n10898), .ZN(n10909) );
  NAND2_X1 U9440 ( .A1(n10909), .A2(n9156), .ZN(n8825) );
  AOI21_X1 U9441 ( .B1(n8926), .B2(n8422), .A(n5125), .ZN(n10921) );
  AOI22_X1 U9442 ( .A1(n9892), .A2(n9156), .B1(n9154), .B2(n9890), .ZN(n8263)
         );
  NAND2_X1 U9443 ( .A1(n8325), .A2(n8243), .ZN(n8257) );
  NAND2_X1 U9444 ( .A1(n8257), .A2(n8804), .ZN(n10773) );
  INV_X1 U9445 ( .A(n8812), .ZN(n8259) );
  NAND2_X1 U9446 ( .A1(n9042), .A2(n10873), .ZN(n8260) );
  OAI211_X1 U9447 ( .C1(n8261), .C2(n8926), .A(n10942), .B(n8417), .ZN(n8262)
         );
  OAI211_X1 U9448 ( .C1(n10921), .C2(n10945), .A(n8263), .B(n8262), .ZN(n10924) );
  NAND2_X1 U9449 ( .A1(n10924), .A2(n10957), .ZN(n8272) );
  NAND2_X1 U9450 ( .A1(n8247), .A2(n8241), .ZN(n8264) );
  AND2_X1 U9451 ( .A1(n10891), .A2(n10909), .ZN(n8265) );
  INV_X1 U9452 ( .A(n8423), .ZN(n10922) );
  NAND2_X1 U9453 ( .A1(n8265), .A2(n10922), .ZN(n10933) );
  OR2_X1 U9454 ( .A1(n8265), .A2(n10922), .ZN(n8266) );
  NAND2_X1 U9455 ( .A1(n10933), .A2(n8266), .ZN(n10923) );
  INV_X1 U9456 ( .A(n10923), .ZN(n8270) );
  AOI22_X1 U9457 ( .A1(n10906), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n8267), .B2(
        n10962), .ZN(n8268) );
  OAI21_X1 U9458 ( .B1(n10922), .B2(n10956), .A(n8268), .ZN(n8269) );
  AOI21_X1 U9459 ( .B1(n8270), .B2(n9897), .A(n8269), .ZN(n8271) );
  OAI211_X1 U9460 ( .C1(n10921), .C2(n10953), .A(n8272), .B(n8271), .ZN(
        P2_U3287) );
  INV_X1 U9461 ( .A(n8273), .ZN(n8275) );
  NOR2_X1 U9462 ( .A1(n8275), .A2(n8274), .ZN(n8922) );
  NAND2_X1 U9463 ( .A1(n10945), .A2(n8276), .ZN(n10904) );
  INV_X1 U9464 ( .A(n8922), .ZN(n10708) );
  AOI22_X1 U9465 ( .A1(n10708), .A2(n10942), .B1(n9890), .B2(n9159), .ZN(
        n10710) );
  OAI21_X1 U9466 ( .B1(n8277), .B2(n9849), .A(n10710), .ZN(n8279) );
  INV_X1 U9467 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10650) );
  NOR2_X1 U9468 ( .A1(n10957), .A2(n10650), .ZN(n8278) );
  AOI21_X1 U9469 ( .B1(n8279), .B2(n10957), .A(n8278), .ZN(n8281) );
  OAI21_X1 U9470 ( .B1(n9901), .B2(n9897), .A(n10707), .ZN(n8280) );
  OAI211_X1 U9471 ( .C1(n8922), .C2(n9887), .A(n8281), .B(n8280), .ZN(P2_U3296) );
  INV_X1 U9472 ( .A(n8282), .ZN(n8283) );
  INV_X1 U9473 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9047) );
  OAI22_X1 U9474 ( .A1(n10952), .A2(n8283), .B1(n9047), .B2(n9849), .ZN(n8284)
         );
  AOI21_X1 U9475 ( .B1(n9901), .B2(n9050), .A(n8284), .ZN(n8288) );
  MUX2_X1 U9476 ( .A(n8286), .B(n8285), .S(n10957), .Z(n8287) );
  OAI211_X1 U9477 ( .C1(n8289), .C2(n9887), .A(n8288), .B(n8287), .ZN(P2_U3295) );
  INV_X1 U9478 ( .A(n8290), .ZN(n8293) );
  OAI222_X1 U9479 ( .A1(n9004), .A2(n9530), .B1(n5033), .B2(n8293), .C1(
        P1_U3084), .C2(n8291), .ZN(P1_U3331) );
  OAI222_X1 U9480 ( .A1(n8785), .A2(P2_U3152), .B1(n8693), .B2(n8293), .C1(
        n8292), .C2(n10005), .ZN(P2_U3336) );
  NAND2_X1 U9481 ( .A1(n8298), .A2(n8294), .ZN(n8296) );
  OAI211_X1 U9482 ( .C1(n9731), .C2(n9004), .A(n8296), .B(n8295), .ZN(P1_U3330) );
  NAND2_X1 U9483 ( .A1(n8298), .A2(n8297), .ZN(n8299) );
  OAI211_X1 U9484 ( .C1(n8300), .C2(n10005), .A(n8299), .B(n8958), .ZN(
        P2_U3335) );
  XNOR2_X1 U9485 ( .A(n8303), .B(n8302), .ZN(n8304) );
  XNOR2_X1 U9486 ( .A(n8301), .B(n8304), .ZN(n8312) );
  NAND2_X1 U9487 ( .A1(n10152), .A2(n8305), .ZN(n8308) );
  INV_X1 U9488 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8306) );
  NOR2_X1 U9489 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8306), .ZN(n10184) );
  AOI21_X1 U9490 ( .B1(n10147), .B2(n10167), .A(n10184), .ZN(n8307) );
  OAI211_X1 U9491 ( .C1(n8309), .C2(n10149), .A(n8308), .B(n8307), .ZN(n8310)
         );
  AOI21_X1 U9492 ( .B1(n8385), .B2(n10131), .A(n8310), .ZN(n8311) );
  OAI21_X1 U9493 ( .B1(n8312), .B2(n10133), .A(n8311), .ZN(P1_U3222) );
  AOI22_X1 U9494 ( .A1(n8313), .A2(n10515), .B1(n10739), .B2(n8475), .ZN(n8314) );
  OAI211_X1 U9495 ( .C1(n8316), .C2(n10741), .A(n8315), .B(n8314), .ZN(n8319)
         );
  NAND2_X1 U9496 ( .A1(n8319), .A2(n11093), .ZN(n8317) );
  OAI21_X1 U9497 ( .B1(n11093), .B2(n8318), .A(n8317), .ZN(P1_U3533) );
  INV_X1 U9498 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U9499 ( .A1(n8319), .A2(n11097), .ZN(n8320) );
  OAI21_X1 U9500 ( .B1(n11097), .B2(n8321), .A(n8320), .ZN(P1_U3484) );
  NAND2_X1 U9501 ( .A1(n8322), .A2(n8323), .ZN(n8324) );
  XNOR2_X1 U9502 ( .A(n8324), .B(n8243), .ZN(n10749) );
  XNOR2_X1 U9503 ( .A(n8325), .B(n8243), .ZN(n8328) );
  OAI22_X1 U9504 ( .A1(n8326), .A2(n10939), .B1(n8189), .B2(n10937), .ZN(n8327) );
  AOI21_X1 U9505 ( .B1(n8328), .B2(n10942), .A(n8327), .ZN(n8329) );
  OAI21_X1 U9506 ( .B1(n10749), .B2(n10945), .A(n8329), .ZN(n10751) );
  INV_X1 U9507 ( .A(n10751), .ZN(n8337) );
  NOR2_X1 U9508 ( .A1(n10749), .A2(n10953), .ZN(n8335) );
  NOR2_X1 U9509 ( .A1(n10956), .A2(n8241), .ZN(n8334) );
  INV_X1 U9510 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8330) );
  OAI22_X1 U9511 ( .A1(n10957), .A2(n8330), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9849), .ZN(n8333) );
  XNOR2_X1 U9512 ( .A(n10770), .B(n8331), .ZN(n10750) );
  NOR2_X1 U9513 ( .A1(n10952), .A2(n10750), .ZN(n8332) );
  NOR4_X1 U9514 ( .A1(n8335), .A2(n8334), .A3(n8333), .A4(n8332), .ZN(n8336)
         );
  OAI21_X1 U9515 ( .B1(n10906), .B2(n8337), .A(n8336), .ZN(P2_U3293) );
  NOR2_X1 U9516 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8380) );
  NOR2_X1 U9517 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8378) );
  NOR2_X1 U9518 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8375) );
  NOR2_X1 U9519 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8373) );
  NOR2_X1 U9520 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8370) );
  NOR2_X1 U9521 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8367) );
  NAND2_X1 U9522 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8364) );
  XOR2_X1 U9523 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10572) );
  NAND2_X1 U9524 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8362) );
  XNOR2_X1 U9525 ( .A(n8338), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n10570) );
  NOR2_X1 U9526 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8346) );
  XOR2_X1 U9527 ( .A(n8339), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10560) );
  NAND2_X1 U9528 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8344) );
  XNOR2_X1 U9529 ( .A(n8340), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n10558) );
  NAND2_X1 U9530 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n8342) );
  XOR2_X1 U9531 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10556) );
  AOI21_X1 U9532 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10550) );
  INV_X1 U9533 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10554) );
  NAND3_X1 U9534 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10552) );
  OAI21_X1 U9535 ( .B1(n10550), .B2(n10554), .A(n10552), .ZN(n10555) );
  NAND2_X1 U9536 ( .A1(n10556), .A2(n10555), .ZN(n8341) );
  NAND2_X1 U9537 ( .A1(n8342), .A2(n8341), .ZN(n10557) );
  NAND2_X1 U9538 ( .A1(n10558), .A2(n10557), .ZN(n8343) );
  NAND2_X1 U9539 ( .A1(n8344), .A2(n8343), .ZN(n10559) );
  NOR2_X1 U9540 ( .A1(n10560), .A2(n10559), .ZN(n8345) );
  NOR2_X1 U9541 ( .A1(n8346), .A2(n8345), .ZN(n8347) );
  NOR2_X1 U9542 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8347), .ZN(n10561) );
  AND2_X1 U9543 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8347), .ZN(n10562) );
  NOR2_X1 U9544 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10562), .ZN(n8348) );
  NAND2_X1 U9545 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n8349), .ZN(n8351) );
  XOR2_X1 U9546 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n8349), .Z(n10564) );
  NAND2_X1 U9547 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10564), .ZN(n8350) );
  NAND2_X1 U9548 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  NAND2_X1 U9549 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n8352), .ZN(n8354) );
  XOR2_X1 U9550 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n8352), .Z(n10565) );
  NAND2_X1 U9551 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10565), .ZN(n8353) );
  NAND2_X1 U9552 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  NAND2_X1 U9553 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n8355), .ZN(n8357) );
  XOR2_X1 U9554 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n8355), .Z(n10566) );
  NAND2_X1 U9555 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10566), .ZN(n8356) );
  NAND2_X1 U9556 ( .A1(n8357), .A2(n8356), .ZN(n8358) );
  NAND2_X1 U9557 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n8358), .ZN(n8360) );
  XOR2_X1 U9558 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n8358), .Z(n10567) );
  NAND2_X1 U9559 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10567), .ZN(n8359) );
  NAND2_X1 U9560 ( .A1(n8360), .A2(n8359), .ZN(n10569) );
  NAND2_X1 U9561 ( .A1(n10570), .A2(n10569), .ZN(n8361) );
  NAND2_X1 U9562 ( .A1(n8362), .A2(n8361), .ZN(n10571) );
  NAND2_X1 U9563 ( .A1(n10572), .A2(n10571), .ZN(n8363) );
  NAND2_X1 U9564 ( .A1(n8364), .A2(n8363), .ZN(n10574) );
  XOR2_X1 U9565 ( .A(n8365), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n10573) );
  XOR2_X1 U9566 ( .A(n8368), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n10575) );
  XOR2_X1 U9567 ( .A(n8371), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n10577) );
  NOR2_X1 U9568 ( .A1(n10578), .A2(n10577), .ZN(n8372) );
  NOR2_X1 U9569 ( .A1(n8373), .A2(n8372), .ZN(n10580) );
  INV_X1 U9570 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9163) );
  XOR2_X1 U9571 ( .A(n9163), .B(P1_ADDR_REG_15__SCAN_IN), .Z(n10579) );
  NOR2_X1 U9572 ( .A1(n10580), .A2(n10579), .ZN(n8374) );
  NOR2_X1 U9573 ( .A1(n8375), .A2(n8374), .ZN(n10582) );
  XOR2_X1 U9574 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n8376), .Z(n10581) );
  NOR2_X1 U9575 ( .A1(n10582), .A2(n10581), .ZN(n8377) );
  NOR2_X1 U9576 ( .A1(n8378), .A2(n8377), .ZN(n10584) );
  INV_X1 U9577 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9208) );
  XOR2_X1 U9578 ( .A(n9208), .B(P1_ADDR_REG_17__SCAN_IN), .Z(n10583) );
  NOR2_X1 U9579 ( .A1(n10584), .A2(n10583), .ZN(n8379) );
  NOR2_X1 U9580 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  AND2_X1 U9581 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8381), .ZN(n10585) );
  NOR2_X1 U9582 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10585), .ZN(n8382) );
  NOR2_X1 U9583 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n8381), .ZN(n10586) );
  NOR2_X1 U9584 ( .A1(n8382), .A2(n10586), .ZN(n8384) );
  XNOR2_X1 U9585 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8383) );
  XNOR2_X1 U9586 ( .A(n8384), .B(n8383), .ZN(ADD_1071_U4) );
  NAND2_X1 U9587 ( .A1(n8385), .A2(n11005), .ZN(n8386) );
  OR2_X1 U9588 ( .A1(n8552), .A2(n10167), .ZN(n8522) );
  NAND2_X1 U9589 ( .A1(n10997), .A2(n8522), .ZN(n8388) );
  XNOR2_X1 U9590 ( .A(n8388), .B(n5054), .ZN(n11047) );
  INV_X1 U9591 ( .A(n11047), .ZN(n8400) );
  OAI211_X1 U9592 ( .C1(n5622), .C2(n8392), .A(n8512), .B(n11009), .ZN(n8394)
         );
  AOI22_X1 U9593 ( .A1(n11006), .A2(n10167), .B1(n8659), .B2(n11003), .ZN(
        n8393) );
  NAND2_X1 U9594 ( .A1(n8394), .A2(n8393), .ZN(n11045) );
  INV_X1 U9595 ( .A(n11001), .ZN(n8395) );
  OAI21_X1 U9596 ( .B1(n8395), .B2(n5338), .A(n8516), .ZN(n11044) );
  AOI22_X1 U9597 ( .A1(n11027), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8657), .B2(
        n11025), .ZN(n8397) );
  NAND2_X1 U9598 ( .A1(n8664), .A2(n10413), .ZN(n8396) );
  OAI211_X1 U9599 ( .C1(n11044), .C2(n10378), .A(n8397), .B(n8396), .ZN(n8398)
         );
  AOI21_X1 U9600 ( .B1(n11045), .B2(n10869), .A(n8398), .ZN(n8399) );
  OAI21_X1 U9601 ( .B1(n8400), .B2(n10442), .A(n8399), .ZN(P1_U3277) );
  INV_X1 U9602 ( .A(n8401), .ZN(n8402) );
  AOI21_X1 U9603 ( .B1(n8403), .B2(n8402), .A(n9086), .ZN(n8406) );
  NOR3_X1 U9604 ( .A1(n8404), .A2(n9122), .A3(n8418), .ZN(n8405) );
  OAI21_X1 U9605 ( .B1(n8406), .B2(n8405), .A(n8477), .ZN(n8413) );
  OR2_X1 U9606 ( .A1(n8716), .A2(n10939), .ZN(n8408) );
  OR2_X1 U9607 ( .A1(n8418), .A2(n10937), .ZN(n8407) );
  NAND2_X1 U9608 ( .A1(n8408), .A2(n8407), .ZN(n8437) );
  INV_X1 U9609 ( .A(n8440), .ZN(n8409) );
  NOR2_X1 U9610 ( .A1(n9141), .A2(n8409), .ZN(n8410) );
  AOI211_X1 U9611 ( .C1(n9143), .C2(n8437), .A(n8411), .B(n8410), .ZN(n8412)
         );
  OAI211_X1 U9612 ( .C1(n5354), .C2(n9146), .A(n8413), .B(n8412), .ZN(P2_U3238) );
  INV_X1 U9613 ( .A(n8414), .ZN(n8461) );
  OAI222_X1 U9614 ( .A1(n5033), .A2(n8461), .B1(P1_U3084), .B2(n8416), .C1(
        n8415), .C2(n9004), .ZN(P1_U3329) );
  OR2_X1 U9615 ( .A1(n10932), .A2(n8418), .ZN(n8834) );
  NAND2_X1 U9616 ( .A1(n10932), .A2(n8418), .ZN(n8836) );
  NAND2_X1 U9617 ( .A1(n8834), .A2(n8836), .ZN(n10931) );
  NAND2_X1 U9618 ( .A1(n10974), .A2(n10940), .ZN(n8837) );
  INV_X1 U9619 ( .A(n8837), .ZN(n8419) );
  OR2_X1 U9620 ( .A1(n10974), .A2(n10940), .ZN(n8835) );
  OAI21_X1 U9621 ( .B1(n8539), .B2(n8419), .A(n8835), .ZN(n8420) );
  OR2_X1 U9622 ( .A1(n8535), .A2(n8716), .ZN(n8845) );
  NAND2_X1 U9623 ( .A1(n8535), .A2(n8716), .ZN(n8541) );
  XNOR2_X1 U9624 ( .A(n8420), .B(n8844), .ZN(n8421) );
  OAI222_X1 U9625 ( .A1(n10939), .A2(n8744), .B1(n10937), .B2(n10940), .C1(
        n10811), .C2(n8421), .ZN(n10992) );
  INV_X1 U9626 ( .A(n10992), .ZN(n8435) );
  INV_X1 U9627 ( .A(n10938), .ZN(n9155) );
  NAND2_X1 U9628 ( .A1(n10932), .A2(n9154), .ZN(n8424) );
  NAND2_X1 U9629 ( .A1(n10930), .A2(n8424), .ZN(n8443) );
  NAND2_X1 U9630 ( .A1(n8835), .A2(n8837), .ZN(n8928) );
  NAND2_X1 U9631 ( .A1(n8443), .A2(n8928), .ZN(n8442) );
  INV_X1 U9632 ( .A(n10940), .ZN(n9153) );
  NAND2_X1 U9633 ( .A1(n10974), .A2(n9153), .ZN(n8425) );
  NAND2_X1 U9634 ( .A1(n8442), .A2(n8425), .ZN(n8426) );
  INV_X1 U9635 ( .A(n8844), .ZN(n8929) );
  OR2_X1 U9636 ( .A1(n8426), .A2(n8844), .ZN(n8427) );
  OAI21_X1 U9637 ( .B1(n8537), .B2(n8929), .A(n8427), .ZN(n10994) );
  INV_X1 U9638 ( .A(n9887), .ZN(n10790) );
  INV_X1 U9639 ( .A(n8535), .ZN(n10990) );
  NOR2_X1 U9640 ( .A1(n8428), .A2(n10990), .ZN(n8429) );
  OR2_X1 U9641 ( .A1(n8569), .A2(n8429), .ZN(n10991) );
  INV_X1 U9642 ( .A(n8481), .ZN(n8430) );
  OAI22_X1 U9643 ( .A1(n10957), .A2(n7988), .B1(n8430), .B2(n9849), .ZN(n8431)
         );
  AOI21_X1 U9644 ( .B1(n9901), .B2(n8535), .A(n8431), .ZN(n8432) );
  OAI21_X1 U9645 ( .B1(n10991), .B2(n10952), .A(n8432), .ZN(n8433) );
  AOI21_X1 U9646 ( .B1(n10994), .B2(n10790), .A(n8433), .ZN(n8434) );
  OAI21_X1 U9647 ( .B1(n8435), .B2(n10906), .A(n8434), .ZN(P2_U3284) );
  INV_X1 U9648 ( .A(n8928), .ZN(n8436) );
  XNOR2_X1 U9649 ( .A(n8539), .B(n8436), .ZN(n8438) );
  AOI21_X1 U9650 ( .B1(n8438), .B2(n10942), .A(n8437), .ZN(n10977) );
  AND2_X1 U9651 ( .A1(n10957), .A2(n9846), .ZN(n9880) );
  XNOR2_X1 U9652 ( .A(n5122), .B(n10974), .ZN(n8439) );
  NOR2_X1 U9653 ( .A1(n8439), .A2(n11070), .ZN(n10973) );
  AOI22_X1 U9654 ( .A1(n10906), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8440), .B2(
        n10962), .ZN(n8441) );
  OAI21_X1 U9655 ( .B1(n5354), .B2(n10956), .A(n8441), .ZN(n8445) );
  OAI21_X1 U9656 ( .B1(n8443), .B2(n8928), .A(n8442), .ZN(n10978) );
  NOR2_X1 U9657 ( .A1(n10978), .A2(n9887), .ZN(n8444) );
  AOI211_X1 U9658 ( .C1(n9880), .C2(n10973), .A(n8445), .B(n8444), .ZN(n8446)
         );
  OAI21_X1 U9659 ( .B1(n10906), .B2(n10977), .A(n8446), .ZN(P2_U3285) );
  XNOR2_X1 U9660 ( .A(n8447), .B(n8925), .ZN(n8451) );
  OAI22_X1 U9661 ( .A1(n8449), .A2(n10937), .B1(n8448), .B2(n10939), .ZN(n8450) );
  AOI21_X1 U9662 ( .B1(n8451), .B2(n10942), .A(n8450), .ZN(n10876) );
  AOI21_X1 U9663 ( .B1(n10873), .B2(n9894), .A(n10891), .ZN(n10874) );
  AOI22_X1 U9664 ( .A1(n10906), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n8452), .B2(
        n10962), .ZN(n8453) );
  OAI21_X1 U9665 ( .B1(n8820), .B2(n10956), .A(n8453), .ZN(n8458) );
  INV_X1 U9666 ( .A(n8454), .ZN(n8455) );
  AOI21_X1 U9667 ( .B1(n8925), .B2(n8456), .A(n8455), .ZN(n10877) );
  NOR2_X1 U9668 ( .A1(n10877), .A2(n9887), .ZN(n8457) );
  AOI211_X1 U9669 ( .C1(n9897), .C2(n10874), .A(n8458), .B(n8457), .ZN(n8459)
         );
  OAI21_X1 U9670 ( .B1(n10906), .B2(n10876), .A(n8459), .ZN(P2_U3289) );
  OAI222_X1 U9671 ( .A1(n8462), .A2(P2_U3152), .B1(n8693), .B2(n8461), .C1(
        n8460), .C2(n10005), .ZN(P2_U3334) );
  NAND2_X1 U9672 ( .A1(n10152), .A2(n8463), .ZN(n8466) );
  AOI21_X1 U9673 ( .B1(n10147), .B2(n10168), .A(n8464), .ZN(n8465) );
  OAI211_X1 U9674 ( .C1(n8467), .C2(n10149), .A(n8466), .B(n8465), .ZN(n8474)
         );
  NAND2_X1 U9675 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  XOR2_X1 U9676 ( .A(n8471), .B(n8470), .Z(n8472) );
  NOR2_X1 U9677 ( .A1(n8472), .A2(n10133), .ZN(n8473) );
  AOI211_X1 U9678 ( .C1(n8475), .C2(n10131), .A(n8474), .B(n8473), .ZN(n8476)
         );
  INV_X1 U9679 ( .A(n8476), .ZN(P1_U3215) );
  INV_X1 U9680 ( .A(n8477), .ZN(n8480) );
  NOR3_X1 U9681 ( .A1(n8478), .A2(n10940), .A3(n9122), .ZN(n8479) );
  AOI21_X1 U9682 ( .B1(n8480), .B2(n9135), .A(n8479), .ZN(n8489) );
  INV_X1 U9683 ( .A(n8720), .ZN(n8487) );
  INV_X1 U9684 ( .A(n8744), .ZN(n9151) );
  AOI22_X1 U9685 ( .A1(n8739), .A2(n9151), .B1(n9129), .B2(n8481), .ZN(n8485)
         );
  NAND2_X1 U9686 ( .A1(n8535), .A2(n9098), .ZN(n8483) );
  NAND2_X1 U9687 ( .A1(n9125), .A2(n9153), .ZN(n8482) );
  NAND4_X1 U9688 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n8486)
         );
  AOI21_X1 U9689 ( .B1(n8487), .B2(n9135), .A(n8486), .ZN(n8488) );
  OAI21_X1 U9690 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(P2_U3226) );
  INV_X1 U9691 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8492) );
  NOR2_X1 U9692 ( .A1(n10244), .A2(n8492), .ZN(n8491) );
  AOI21_X1 U9693 ( .B1(n10244), .B2(n8492), .A(n8491), .ZN(n8496) );
  AOI21_X1 U9694 ( .B1(n8499), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8493), .ZN(
        n10230) );
  NAND2_X1 U9695 ( .A1(n10227), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8494) );
  OAI21_X1 U9696 ( .B1(n10227), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8494), .ZN(
        n10229) );
  NOR2_X1 U9697 ( .A1(n10230), .A2(n10229), .ZN(n10228) );
  AOI21_X1 U9698 ( .B1(n10227), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10228), .ZN(
        n8495) );
  NOR2_X1 U9699 ( .A1(n8495), .A2(n8496), .ZN(n10243) );
  AOI211_X1 U9700 ( .C1(n8496), .C2(n8495), .A(n10243), .B(n10248), .ZN(n8510)
         );
  NOR2_X1 U9701 ( .A1(n10244), .A2(n8497), .ZN(n8498) );
  AOI21_X1 U9702 ( .B1(n8497), .B2(n10244), .A(n8498), .ZN(n8505) );
  INV_X1 U9703 ( .A(n10227), .ZN(n8503) );
  XNOR2_X1 U9704 ( .A(n8503), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10234) );
  INV_X1 U9705 ( .A(n8499), .ZN(n8501) );
  INV_X1 U9706 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11092) );
  OAI21_X1 U9707 ( .B1(n8501), .B2(n11092), .A(n8500), .ZN(n10233) );
  NAND2_X1 U9708 ( .A1(n10234), .A2(n10233), .ZN(n10232) );
  OAI21_X1 U9709 ( .B1(n8503), .B2(n8502), .A(n10232), .ZN(n8504) );
  NOR2_X1 U9710 ( .A1(n8504), .A2(n8505), .ZN(n10238) );
  AOI21_X1 U9711 ( .B1(n8505), .B2(n8504), .A(n10238), .ZN(n8506) );
  NOR2_X1 U9712 ( .A1(n8506), .A2(n10695), .ZN(n8509) );
  INV_X1 U9713 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U9714 ( .A1(n10692), .A2(n10244), .ZN(n8507) );
  NAND2_X1 U9715 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10116) );
  OAI211_X1 U9716 ( .C1(n10631), .C2(n10588), .A(n8507), .B(n10116), .ZN(n8508) );
  OR3_X1 U9717 ( .A1(n8510), .A2(n8509), .A3(n8508), .ZN(P1_U3259) );
  NAND2_X1 U9718 ( .A1(n8512), .A2(n8511), .ZN(n8513) );
  OAI211_X1 U9719 ( .C1(n8528), .C2(n8513), .A(n8602), .B(n11009), .ZN(n8515)
         );
  AOI22_X1 U9720 ( .A1(n11006), .A2(n11004), .B1(n10146), .B2(n11003), .ZN(
        n8514) );
  NAND2_X1 U9721 ( .A1(n8515), .A2(n8514), .ZN(n11063) );
  AND2_X1 U9722 ( .A1(n8516), .A2(n10135), .ZN(n8517) );
  NOR2_X2 U9723 ( .A1(n8516), .A2(n10135), .ZN(n8587) );
  OR2_X1 U9724 ( .A1(n8517), .A2(n8587), .ZN(n11062) );
  AOI22_X1 U9725 ( .A1(n11027), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10153), 
        .B2(n11025), .ZN(n8519) );
  NAND2_X1 U9726 ( .A1(n10135), .A2(n10413), .ZN(n8518) );
  OAI211_X1 U9727 ( .C1(n11062), .C2(n10378), .A(n8519), .B(n8518), .ZN(n8532)
         );
  OR2_X1 U9728 ( .A1(n8664), .A2(n11004), .ZN(n8521) );
  INV_X1 U9729 ( .A(n8521), .ZN(n8520) );
  NOR2_X1 U9730 ( .A1(n8520), .A2(n5054), .ZN(n8524) );
  OR2_X1 U9731 ( .A1(n10999), .A2(n8581), .ZN(n8527) );
  INV_X1 U9732 ( .A(n8528), .ZN(n8525) );
  AND2_X1 U9733 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  OR2_X1 U9734 ( .A1(n8524), .A2(n8523), .ZN(n8526) );
  AND2_X1 U9735 ( .A1(n8525), .A2(n8526), .ZN(n8582) );
  NAND2_X1 U9736 ( .A1(n8527), .A2(n8582), .ZN(n11065) );
  INV_X1 U9737 ( .A(n11065), .ZN(n8530) );
  NAND2_X1 U9738 ( .A1(n8527), .A2(n8526), .ZN(n8529) );
  NOR3_X1 U9739 ( .A1(n8530), .A2(n11060), .A3(n10442), .ZN(n8531) );
  AOI211_X1 U9740 ( .C1(n10869), .C2(n11063), .A(n8532), .B(n8531), .ZN(n8533)
         );
  INV_X1 U9741 ( .A(n8533), .ZN(P1_U3276) );
  NAND2_X1 U9742 ( .A1(n11051), .A2(n9150), .ZN(n8534) );
  NAND2_X1 U9743 ( .A1(n8635), .A2(n8534), .ZN(n8932) );
  INV_X1 U9744 ( .A(n8714), .ZN(n11036) );
  INV_X1 U9745 ( .A(n8716), .ZN(n9152) );
  OR2_X1 U9746 ( .A1(n8535), .A2(n9152), .ZN(n8536) );
  OR2_X1 U9747 ( .A1(n8714), .A2(n8744), .ZN(n8852) );
  NAND2_X1 U9748 ( .A1(n8714), .A2(n8744), .ZN(n8851) );
  NAND2_X1 U9749 ( .A1(n8852), .A2(n8851), .ZN(n8930) );
  AOI21_X1 U9750 ( .B1(n8932), .B2(n8538), .A(n8637), .ZN(n11050) );
  NAND2_X1 U9751 ( .A1(n8541), .A2(n8837), .ZN(n8846) );
  INV_X1 U9752 ( .A(n8835), .ZN(n8540) );
  NAND2_X1 U9753 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U9754 ( .A1(n8542), .A2(n8845), .ZN(n8565) );
  NOR2_X1 U9755 ( .A1(n8930), .A2(n8565), .ZN(n8543) );
  AND2_X1 U9756 ( .A1(n8564), .A2(n8851), .ZN(n8545) );
  AND2_X1 U9757 ( .A1(n8932), .A2(n8851), .ZN(n8544) );
  OAI211_X1 U9758 ( .C1(n8545), .C2(n8932), .A(n10942), .B(n8639), .ZN(n8547)
         );
  OR2_X1 U9759 ( .A1(n8670), .A2(n10939), .ZN(n8546) );
  OAI211_X1 U9760 ( .C1(n8744), .C2(n10937), .A(n8547), .B(n8546), .ZN(n11055)
         );
  XNOR2_X1 U9761 ( .A(n8641), .B(n11051), .ZN(n11053) );
  AOI22_X1 U9762 ( .A1(n10906), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8738), .B2(
        n10962), .ZN(n8549) );
  NAND2_X1 U9763 ( .A1(n11051), .A2(n9901), .ZN(n8548) );
  OAI211_X1 U9764 ( .C1(n11053), .C2(n10952), .A(n8549), .B(n8548), .ZN(n8550)
         );
  AOI21_X1 U9765 ( .B1(n11055), .B2(n10957), .A(n8550), .ZN(n8551) );
  OAI21_X1 U9766 ( .B1(n11050), .B2(n9887), .A(n8551), .ZN(P2_U3282) );
  OAI21_X1 U9767 ( .B1(n5493), .B2(n8556), .A(n8555), .ZN(n8557) );
  OAI21_X1 U9768 ( .B1(n8553), .B2(n5493), .A(n8557), .ZN(n8558) );
  NAND2_X1 U9769 ( .A1(n8558), .A2(n10143), .ZN(n8563) );
  AND2_X1 U9770 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10200) );
  AOI21_X1 U9771 ( .B1(n10147), .B2(n11004), .A(n10200), .ZN(n8559) );
  OAI21_X1 U9772 ( .B1(n8560), .B2(n10149), .A(n8559), .ZN(n8561) );
  AOI21_X1 U9773 ( .B1(n11026), .B2(n10152), .A(n8561), .ZN(n8562) );
  OAI211_X1 U9774 ( .C1(n5339), .C2(n10156), .A(n8563), .B(n8562), .ZN(
        P1_U3232) );
  INV_X1 U9775 ( .A(n9150), .ZN(n8854) );
  INV_X1 U9776 ( .A(n8564), .ZN(n8567) );
  INV_X1 U9777 ( .A(n8565), .ZN(n8847) );
  INV_X1 U9778 ( .A(n8930), .ZN(n8850) );
  AOI21_X1 U9779 ( .B1(n5466), .B2(n8847), .A(n8850), .ZN(n8566) );
  NOR2_X1 U9780 ( .A1(n8567), .A2(n8566), .ZN(n8568) );
  OAI222_X1 U9781 ( .A1(n10939), .A2(n8854), .B1(n10937), .B2(n8716), .C1(
        n10811), .C2(n8568), .ZN(n11038) );
  OAI21_X1 U9782 ( .B1(n8569), .B2(n11036), .A(n8641), .ZN(n11037) );
  AOI22_X1 U9783 ( .A1(n10906), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8710), .B2(
        n10962), .ZN(n8571) );
  NAND2_X1 U9784 ( .A1(n8714), .A2(n9901), .ZN(n8570) );
  OAI211_X1 U9785 ( .C1(n11037), .C2(n10952), .A(n8571), .B(n8570), .ZN(n8574)
         );
  NOR2_X1 U9786 ( .A1(n5118), .A2(n8930), .ZN(n11035) );
  INV_X1 U9787 ( .A(n11040), .ZN(n8572) );
  NOR3_X1 U9788 ( .A1(n11035), .A2(n8572), .A3(n9887), .ZN(n8573) );
  AOI211_X1 U9789 ( .C1(n10957), .C2(n11038), .A(n8574), .B(n8573), .ZN(n8575)
         );
  INV_X1 U9790 ( .A(n8575), .ZN(P2_U3283) );
  NAND2_X1 U9791 ( .A1(n8602), .A2(n8576), .ZN(n8577) );
  XNOR2_X1 U9792 ( .A(n8577), .B(n8584), .ZN(n8578) );
  NAND2_X1 U9793 ( .A1(n8578), .A2(n11009), .ZN(n8580) );
  INV_X1 U9794 ( .A(n8626), .ZN(n10166) );
  AOI22_X1 U9795 ( .A1(n10166), .A2(n11003), .B1(n11006), .B2(n8659), .ZN(
        n8579) );
  NAND2_X1 U9796 ( .A1(n8580), .A2(n8579), .ZN(n11087) );
  INV_X1 U9797 ( .A(n11087), .ZN(n8592) );
  AND2_X1 U9798 ( .A1(n10135), .A2(n8659), .ZN(n8583) );
  OAI21_X1 U9799 ( .B1(n8585), .B2(n8584), .A(n8599), .ZN(n8586) );
  INV_X1 U9800 ( .A(n8586), .ZN(n11090) );
  NAND2_X1 U9801 ( .A1(n8587), .A2(n11084), .ZN(n8611) );
  OAI21_X1 U9802 ( .B1(n8587), .B2(n11084), .A(n8611), .ZN(n11086) );
  AOI22_X1 U9803 ( .A1(n11027), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10064), 
        .B2(n11025), .ZN(n8589) );
  NAND2_X1 U9804 ( .A1(n10069), .A2(n10413), .ZN(n8588) );
  OAI211_X1 U9805 ( .C1(n11086), .C2(n10378), .A(n8589), .B(n8588), .ZN(n8590)
         );
  AOI21_X1 U9806 ( .B1(n11090), .B2(n8632), .A(n8590), .ZN(n8591) );
  OAI21_X1 U9807 ( .B1(n11027), .B2(n8592), .A(n8591), .ZN(P1_U3275) );
  INV_X1 U9808 ( .A(n8593), .ZN(n8596) );
  OAI222_X1 U9809 ( .A1(n9004), .A2(n9526), .B1(n5033), .B2(n8596), .C1(n8594), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9810 ( .A1(P2_U3152), .A2(n8597), .B1(n10012), .B2(n8596), .C1(
        n8595), .C2(n10005), .ZN(P2_U3333) );
  NAND2_X1 U9811 ( .A1(n10069), .A2(n10146), .ZN(n8598) );
  OAI21_X1 U9812 ( .B1(n8600), .B2(n8607), .A(n8629), .ZN(n10513) );
  OAI22_X1 U9813 ( .A1(n10430), .A2(n10851), .B1(n10076), .B2(n10849), .ZN(
        n8609) );
  INV_X1 U9814 ( .A(n8618), .ZN(n8605) );
  AOI211_X1 U9815 ( .C1(n8607), .C2(n8606), .A(n10429), .B(n8605), .ZN(n8608)
         );
  AOI211_X1 U9816 ( .C1(n10746), .C2(n10513), .A(n8609), .B(n8608), .ZN(n10518) );
  INV_X1 U9817 ( .A(n8610), .ZN(n8620) );
  AOI21_X1 U9818 ( .B1(n10514), .B2(n8611), .A(n8610), .ZN(n10516) );
  INV_X1 U9819 ( .A(n10514), .ZN(n8627) );
  NOR2_X1 U9820 ( .A1(n8627), .A2(n11029), .ZN(n8614) );
  INV_X1 U9821 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8612) );
  OAI22_X1 U9822 ( .A1(n10869), .A2(n8612), .B1(n10079), .B2(n10865), .ZN(
        n8613) );
  AOI211_X1 U9823 ( .C1(n10516), .C2(n11022), .A(n8614), .B(n8613), .ZN(n8616)
         );
  NAND2_X1 U9824 ( .A1(n10513), .A2(n11023), .ZN(n8615) );
  OAI211_X1 U9825 ( .C1(n10518), .C2(n11027), .A(n8616), .B(n8615), .ZN(
        P1_U3274) );
  XOR2_X1 U9826 ( .A(n8974), .B(n8973), .Z(n8619) );
  AOI222_X1 U9827 ( .A1(n11009), .A2(n8619), .B1(n10164), .B2(n11003), .C1(
        n10166), .C2(n11006), .ZN(n10512) );
  NOR2_X2 U9828 ( .A1(n8620), .A2(n10507), .ZN(n10432) );
  NAND2_X1 U9829 ( .A1(n8620), .A2(n10507), .ZN(n8621) );
  NAND2_X1 U9830 ( .A1(n8621), .A2(n10515), .ZN(n8622) );
  NOR2_X1 U9831 ( .A1(n10432), .A2(n8622), .ZN(n10506) );
  NAND2_X1 U9832 ( .A1(n10507), .A2(n10413), .ZN(n8624) );
  AOI22_X1 U9833 ( .A1(n11027), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10120), 
        .B2(n11025), .ZN(n8623) );
  NAND2_X1 U9834 ( .A1(n8624), .A2(n8623), .ZN(n8625) );
  AOI21_X1 U9835 ( .B1(n10506), .B2(n10439), .A(n8625), .ZN(n8634) );
  NAND2_X1 U9836 ( .A1(n8627), .A2(n8626), .ZN(n8628) );
  NAND2_X1 U9837 ( .A1(n8629), .A2(n8628), .ZN(n8631) );
  NAND2_X1 U9838 ( .A1(n8631), .A2(n8973), .ZN(n10508) );
  NAND3_X1 U9839 ( .A1(n10509), .A2(n10508), .A3(n8632), .ZN(n8633) );
  OAI211_X1 U9840 ( .C1(n10512), .C2(n11027), .A(n8634), .B(n8633), .ZN(
        P1_U3273) );
  INV_X1 U9841 ( .A(n8635), .ZN(n8636) );
  NAND2_X1 U9842 ( .A1(n8735), .A2(n8670), .ZN(n8859) );
  XNOR2_X1 U9843 ( .A(n8676), .B(n8934), .ZN(n11075) );
  INV_X1 U9844 ( .A(n11075), .ZN(n8648) );
  INV_X1 U9845 ( .A(n9248), .ZN(n9874) );
  OR2_X1 U9846 ( .A1(n11051), .A2(n8854), .ZN(n8638) );
  NAND2_X1 U9847 ( .A1(n8639), .A2(n8638), .ZN(n8680) );
  XNOR2_X1 U9848 ( .A(n8680), .B(n8934), .ZN(n8640) );
  OAI222_X1 U9849 ( .A1(n10939), .A2(n9874), .B1(n10937), .B2(n8854), .C1(
        n10811), .C2(n8640), .ZN(n11073) );
  INV_X1 U9850 ( .A(n8642), .ZN(n8643) );
  OAI21_X1 U9851 ( .B1(n8643), .B2(n5215), .A(n8683), .ZN(n11071) );
  AOI22_X1 U9852 ( .A1(n10906), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8727), .B2(
        n10962), .ZN(n8645) );
  NAND2_X1 U9853 ( .A1(n8735), .A2(n9901), .ZN(n8644) );
  OAI211_X1 U9854 ( .C1(n11071), .C2(n10952), .A(n8645), .B(n8644), .ZN(n8646)
         );
  AOI21_X1 U9855 ( .B1(n11073), .B2(n10957), .A(n8646), .ZN(n8647) );
  OAI21_X1 U9856 ( .B1(n8648), .B2(n9887), .A(n8647), .ZN(P2_U3281) );
  INV_X1 U9857 ( .A(n8649), .ZN(n8651) );
  OAI222_X1 U9858 ( .A1(n9004), .A2(n9525), .B1(n5033), .B2(n8651), .C1(n8650), 
        .C2(P1_U3084), .ZN(P1_U3327) );
  OAI222_X1 U9859 ( .A1(P2_U3152), .A2(n8652), .B1(n10012), .B2(n8651), .C1(
        n10005), .C2(n6865), .ZN(P2_U3332) );
  NAND2_X1 U9860 ( .A1(n8654), .A2(n8653), .ZN(n8655) );
  XOR2_X1 U9861 ( .A(n8656), .B(n8655), .Z(n8666) );
  NAND2_X1 U9862 ( .A1(n10152), .A2(n8657), .ZN(n8661) );
  NOR2_X1 U9863 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8658), .ZN(n10216) );
  AOI21_X1 U9864 ( .B1(n10147), .B2(n8659), .A(n10216), .ZN(n8660) );
  OAI211_X1 U9865 ( .C1(n8662), .C2(n10149), .A(n8661), .B(n8660), .ZN(n8663)
         );
  AOI21_X1 U9866 ( .B1(n8664), .B2(n10131), .A(n8663), .ZN(n8665) );
  OAI21_X1 U9867 ( .B1(n8666), .B2(n10133), .A(n8665), .ZN(P1_U3213) );
  INV_X1 U9868 ( .A(n8670), .ZN(n9149) );
  AOI22_X1 U9869 ( .A1(n9149), .A2(n9892), .B1(n9890), .B2(n9862), .ZN(n8681)
         );
  NAND2_X1 U9870 ( .A1(n9129), .A2(n8684), .ZN(n8667) );
  NAND2_X1 U9871 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9184) );
  OAI211_X1 U9872 ( .C1(n8681), .C2(n9080), .A(n8667), .B(n9184), .ZN(n8668)
         );
  AOI21_X1 U9873 ( .B1(n9982), .B2(n9098), .A(n8668), .ZN(n8674) );
  OAI22_X1 U9874 ( .A1(n8671), .A2(n9086), .B1(n8670), .B2(n9122), .ZN(n8672)
         );
  NAND3_X1 U9875 ( .A1(n8737), .A2(n5422), .A3(n8672), .ZN(n8673) );
  OAI211_X1 U9876 ( .C1(n8675), .C2(n9086), .A(n8674), .B(n8673), .ZN(P2_U3228) );
  NAND2_X1 U9877 ( .A1(n8687), .A2(n9248), .ZN(n8864) );
  NAND2_X1 U9878 ( .A1(n9982), .A2(n9874), .ZN(n8863) );
  AOI21_X1 U9879 ( .B1(n8935), .B2(n8677), .A(n9249), .ZN(n8678) );
  INV_X1 U9880 ( .A(n8678), .ZN(n9984) );
  INV_X1 U9881 ( .A(n8860), .ZN(n8679) );
  XOR2_X1 U9882 ( .A(n8756), .B(n8935), .Z(n8682) );
  OAI21_X1 U9883 ( .B1(n8682), .B2(n10811), .A(n8681), .ZN(n9980) );
  AOI211_X1 U9884 ( .C1(n9982), .C2(n8683), .A(n11070), .B(n9877), .ZN(n9981)
         );
  NAND2_X1 U9885 ( .A1(n9981), .A2(n9880), .ZN(n8686) );
  AOI22_X1 U9886 ( .A1(n10906), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8684), .B2(
        n10962), .ZN(n8685) );
  OAI211_X1 U9887 ( .C1(n8687), .C2(n10956), .A(n8686), .B(n8685), .ZN(n8688)
         );
  AOI21_X1 U9888 ( .B1(n9980), .B2(n10957), .A(n8688), .ZN(n8689) );
  OAI21_X1 U9889 ( .B1(n9984), .B2(n9887), .A(n8689), .ZN(P2_U3280) );
  INV_X1 U9890 ( .A(n8690), .ZN(n8694) );
  AOI21_X1 U9891 ( .B1(n10537), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n8691), .ZN(
        n8692) );
  OAI21_X1 U9892 ( .B1(n8694), .B2(n5033), .A(n8692), .ZN(P1_U3326) );
  OAI222_X1 U9893 ( .A1(n7287), .A2(P2_U3152), .B1(n10005), .B2(n6882), .C1(
        n8694), .C2(n8693), .ZN(P2_U3331) );
  OAI222_X1 U9894 ( .A1(n5033), .A2(n8764), .B1(n8696), .B2(P1_U3084), .C1(
        n8695), .C2(n9004), .ZN(P1_U3324) );
  INV_X1 U9895 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8765) );
  OAI222_X1 U9896 ( .A1(P2_U3152), .A2(n8697), .B1(n10012), .B2(n8764), .C1(
        n8765), .C2(n10005), .ZN(P2_U3329) );
  AND2_X1 U9897 ( .A1(n8699), .A2(n8698), .ZN(n8700) );
  NOR2_X1 U9898 ( .A1(n8701), .A2(n8700), .ZN(n8707) );
  OAI22_X1 U9899 ( .A1(n10323), .A2(n10149), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8702), .ZN(n8703) );
  AOI21_X1 U9900 ( .B1(n10291), .B2(n10152), .A(n8703), .ZN(n8704) );
  OAI21_X1 U9901 ( .B1(n10297), .B2(n10118), .A(n8704), .ZN(n8705) );
  AOI21_X1 U9902 ( .B1(n10461), .B2(n10131), .A(n8705), .ZN(n8706) );
  OAI21_X1 U9903 ( .B1(n8707), .B2(n10133), .A(n8706), .ZN(P1_U3212) );
  INV_X1 U9904 ( .A(n8752), .ZN(n10007) );
  OAI222_X1 U9905 ( .A1(n5033), .A2(n10007), .B1(n8709), .B2(P1_U3084), .C1(
        n8708), .C2(n9004), .ZN(P1_U3323) );
  AOI22_X1 U9906 ( .A1(n8739), .A2(n9150), .B1(n9129), .B2(n8710), .ZN(n8712)
         );
  OAI211_X1 U9907 ( .C1(n8716), .C2(n9104), .A(n8712), .B(n8711), .ZN(n8713)
         );
  AOI21_X1 U9908 ( .B1(n8714), .B2(n9098), .A(n8713), .ZN(n8722) );
  INV_X1 U9909 ( .A(n8715), .ZN(n8719) );
  OAI22_X1 U9910 ( .A1(n8717), .A2(n9086), .B1(n8716), .B2(n9122), .ZN(n8718)
         );
  NAND3_X1 U9911 ( .A1(n8720), .A2(n8719), .A3(n8718), .ZN(n8721) );
  OAI211_X1 U9912 ( .C1(n8748), .C2(n9086), .A(n8722), .B(n8721), .ZN(P2_U3236) );
  NAND2_X1 U9913 ( .A1(n8723), .A2(n10143), .ZN(n8726) );
  AOI22_X1 U9914 ( .A1(n10147), .A2(n5704), .B1(n8724), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n8725) );
  OAI211_X1 U9915 ( .C1(n10156), .C2(n7021), .A(n8726), .B(n8725), .ZN(
        P1_U3230) );
  AOI22_X1 U9916 ( .A1(n8739), .A2(n9248), .B1(n9129), .B2(n8727), .ZN(n8728)
         );
  NAND2_X1 U9917 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n9162) );
  OAI211_X1 U9918 ( .C1(n8854), .C2(n9104), .A(n8728), .B(n9162), .ZN(n8734)
         );
  INV_X1 U9919 ( .A(n8751), .ZN(n8732) );
  AOI22_X1 U9920 ( .A1(n8729), .A2(n9135), .B1(n9093), .B2(n9150), .ZN(n8730)
         );
  NOR3_X1 U9921 ( .A1(n8732), .A2(n8731), .A3(n8730), .ZN(n8733) );
  AOI211_X1 U9922 ( .C1(n8735), .C2(n9098), .A(n8734), .B(n8733), .ZN(n8736)
         );
  OAI21_X1 U9923 ( .B1(n8737), .B2(n9086), .A(n8736), .ZN(P2_U3243) );
  AOI22_X1 U9924 ( .A1(n8739), .A2(n9149), .B1(n9129), .B2(n8738), .ZN(n8741)
         );
  OAI211_X1 U9925 ( .C1(n8744), .C2(n9104), .A(n8741), .B(n8740), .ZN(n8742)
         );
  AOI21_X1 U9926 ( .B1(n11051), .B2(n9098), .A(n8742), .ZN(n8750) );
  INV_X1 U9927 ( .A(n8743), .ZN(n8747) );
  OAI22_X1 U9928 ( .A1(n8745), .A2(n9086), .B1(n8744), .B2(n9122), .ZN(n8746)
         );
  NAND3_X1 U9929 ( .A1(n8748), .A2(n8747), .A3(n8746), .ZN(n8749) );
  OAI211_X1 U9930 ( .C1(n8751), .C2(n9086), .A(n8750), .B(n8749), .ZN(P2_U3217) );
  NAND2_X1 U9931 ( .A1(n8752), .A2(n6511), .ZN(n8754) );
  INV_X1 U9932 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10006) );
  OR2_X1 U9933 ( .A1(n5030), .A2(n10006), .ZN(n8753) );
  INV_X1 U9934 ( .A(n8863), .ZN(n8755) );
  NAND2_X1 U9935 ( .A1(n9977), .A2(n9862), .ZN(n8867) );
  INV_X1 U9936 ( .A(n9869), .ZN(n9873) );
  INV_X1 U9937 ( .A(n9977), .ZN(n9884) );
  NAND2_X1 U9938 ( .A1(n9970), .A2(n9876), .ZN(n8869) );
  NAND2_X1 U9939 ( .A1(n9837), .A2(n8869), .ZN(n9860) );
  INV_X1 U9940 ( .A(n9860), .ZN(n9853) );
  OR2_X1 U9941 ( .A1(n9967), .A2(n9251), .ZN(n8872) );
  AND2_X1 U9942 ( .A1(n9837), .A2(n8872), .ZN(n8757) );
  NAND2_X1 U9943 ( .A1(n9967), .A2(n9251), .ZN(n8871) );
  NAND2_X1 U9944 ( .A1(n9960), .A2(n9842), .ZN(n8791) );
  NAND2_X1 U9945 ( .A1(n8792), .A2(n8791), .ZN(n9406) );
  INV_X1 U9946 ( .A(n9406), .ZN(n8940) );
  NAND2_X1 U9947 ( .A1(n8758), .A2(n8792), .ZN(n9391) );
  INV_X1 U9948 ( .A(n9408), .ZN(n9377) );
  NAND2_X1 U9949 ( .A1(n9955), .A2(n9377), .ZN(n8759) );
  NAND2_X1 U9950 ( .A1(n9950), .A2(n9065), .ZN(n8883) );
  NAND2_X1 U9951 ( .A1(n9945), .A2(n9378), .ZN(n9346) );
  INV_X1 U9952 ( .A(n9360), .ZN(n8942) );
  NAND2_X1 U9953 ( .A1(n9939), .A2(n9092), .ZN(n8788) );
  INV_X1 U9954 ( .A(n9346), .ZN(n8761) );
  NOR2_X1 U9955 ( .A1(n9349), .A2(n8761), .ZN(n8762) );
  NAND2_X1 U9956 ( .A1(n9936), .A2(n9350), .ZN(n8897) );
  NAND2_X1 U9957 ( .A1(n9318), .A2(n8897), .ZN(n9257) );
  NAND2_X1 U9958 ( .A1(n9238), .A2(n9260), .ZN(n8918) );
  AND2_X1 U9959 ( .A1(n8918), .A2(n9318), .ZN(n8896) );
  NAND2_X1 U9960 ( .A1(n9924), .A2(n9262), .ZN(n8900) );
  NAND2_X1 U9961 ( .A1(n9311), .A2(n8901), .ZN(n9291) );
  NAND2_X1 U9962 ( .A1(n9919), .A2(n9309), .ZN(n8903) );
  NAND2_X1 U9963 ( .A1(n8904), .A2(n8903), .ZN(n9265) );
  NAND2_X1 U9964 ( .A1(n9291), .A2(n9290), .ZN(n9289) );
  NAND2_X1 U9965 ( .A1(n9289), .A2(n8904), .ZN(n9269) );
  OR2_X1 U9966 ( .A1(n5030), .A2(n8765), .ZN(n8766) );
  NAND2_X1 U9967 ( .A1(n9918), .A2(n8768), .ZN(n8907) );
  NAND2_X1 U9968 ( .A1(n9279), .A2(n9292), .ZN(n8908) );
  INV_X1 U9969 ( .A(n8772), .ZN(n8773) );
  NAND2_X1 U9970 ( .A1(n6549), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U9971 ( .A1(n6533), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U9972 ( .A1(n5060), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8769) );
  INV_X1 U9973 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8775) );
  OR2_X1 U9974 ( .A1(n5030), .A2(n8775), .ZN(n8776) );
  NAND2_X1 U9975 ( .A1(n9244), .A2(n9271), .ZN(n8910) );
  OAI21_X1 U9976 ( .B1(n9907), .B2(n9241), .A(n8910), .ZN(n8916) );
  NAND2_X1 U9977 ( .A1(n9907), .A2(n9241), .ZN(n8782) );
  XNOR2_X1 U9978 ( .A(n8778), .B(n9846), .ZN(n8781) );
  NOR2_X1 U9979 ( .A1(n8781), .A2(n5635), .ZN(n8954) );
  INV_X1 U9980 ( .A(n8916), .ZN(n8787) );
  INV_X1 U9981 ( .A(n8782), .ZN(n8784) );
  INV_X1 U9982 ( .A(n8911), .ZN(n8783) );
  AND2_X1 U9983 ( .A1(n8788), .A2(n9346), .ZN(n8790) );
  AND2_X1 U9984 ( .A1(n8888), .A2(n8882), .ZN(n8789) );
  MUX2_X1 U9985 ( .A(n8790), .B(n8789), .S(n8912), .Z(n8886) );
  MUX2_X1 U9986 ( .A(n8792), .B(n8791), .S(n8906), .Z(n8875) );
  INV_X1 U9987 ( .A(n8325), .ZN(n8796) );
  INV_X1 U9988 ( .A(n8920), .ZN(n8794) );
  AND2_X1 U9989 ( .A1(n8209), .A2(n8793), .ZN(n8797) );
  NAND3_X1 U9990 ( .A1(n8794), .A2(n8947), .A3(n8797), .ZN(n8795) );
  NAND2_X1 U9991 ( .A1(n8796), .A2(n8795), .ZN(n8803) );
  INV_X1 U9992 ( .A(n8797), .ZN(n8799) );
  NAND2_X1 U9993 ( .A1(n8799), .A2(n8798), .ZN(n8801) );
  OAI21_X1 U9994 ( .B1(n8920), .B2(n8801), .A(n8800), .ZN(n8802) );
  MUX2_X1 U9995 ( .A(n8805), .B(n8804), .S(n8912), .Z(n8806) );
  OAI211_X1 U9996 ( .C1(n8807), .C2(n8921), .A(n10768), .B(n8806), .ZN(n8808)
         );
  OAI21_X1 U9997 ( .B1(n8912), .B2(n8809), .A(n8808), .ZN(n8810) );
  NAND2_X1 U9998 ( .A1(n8812), .A2(n8811), .ZN(n8813) );
  NAND2_X1 U9999 ( .A1(n8813), .A2(n8912), .ZN(n8814) );
  AOI21_X1 U10000 ( .B1(n9900), .B2(n5469), .A(n5144), .ZN(n8817) );
  MUX2_X1 U10001 ( .A(n8818), .B(n8817), .S(n8912), .Z(n8819) );
  NAND2_X1 U10002 ( .A1(n10873), .A2(n8906), .ZN(n8822) );
  NAND2_X1 U10003 ( .A1(n8820), .A2(n8912), .ZN(n8821) );
  MUX2_X1 U10004 ( .A(n8822), .B(n8821), .S(n9891), .Z(n8823) );
  MUX2_X1 U10005 ( .A(n8825), .B(n8824), .S(n8912), .Z(n8826) );
  NAND3_X1 U10006 ( .A1(n8827), .A2(n8828), .A3(n8826), .ZN(n8833) );
  NAND2_X1 U10007 ( .A1(n8834), .A2(n8828), .ZN(n8830) );
  INV_X1 U10008 ( .A(n8829), .ZN(n8839) );
  MUX2_X1 U10009 ( .A(n8830), .B(n8839), .S(n8906), .Z(n8832) );
  INV_X1 U10010 ( .A(n8836), .ZN(n8831) );
  NOR2_X1 U10011 ( .A1(n8832), .A2(n8831), .ZN(n8840) );
  AND2_X1 U10012 ( .A1(n8835), .A2(n8834), .ZN(n8842) );
  NAND2_X1 U10013 ( .A1(n8837), .A2(n8836), .ZN(n8838) );
  AOI21_X1 U10014 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8841) );
  MUX2_X1 U10015 ( .A(n8842), .B(n8841), .S(n8912), .Z(n8843) );
  NAND2_X1 U10016 ( .A1(n8846), .A2(n8845), .ZN(n8848) );
  MUX2_X1 U10017 ( .A(n8848), .B(n8847), .S(n8912), .Z(n8849) );
  MUX2_X1 U10018 ( .A(n8852), .B(n8851), .S(n8912), .Z(n8853) );
  NAND2_X1 U10019 ( .A1(n9150), .A2(n8912), .ZN(n8856) );
  NAND2_X1 U10020 ( .A1(n8854), .A2(n8906), .ZN(n8855) );
  MUX2_X1 U10021 ( .A(n8856), .B(n8855), .S(n11051), .Z(n8857) );
  NAND3_X1 U10022 ( .A1(n8858), .A2(n8934), .A3(n8857), .ZN(n8862) );
  MUX2_X1 U10023 ( .A(n8860), .B(n8859), .S(n8912), .Z(n8861) );
  NAND3_X1 U10024 ( .A1(n8862), .A2(n8935), .A3(n8861), .ZN(n8866) );
  MUX2_X1 U10025 ( .A(n8864), .B(n8863), .S(n8906), .Z(n8865) );
  MUX2_X1 U10026 ( .A(n9977), .B(n9862), .S(n8912), .Z(n8868) );
  NAND2_X1 U10027 ( .A1(n8872), .A2(n8871), .ZN(n9835) );
  INV_X1 U10028 ( .A(n9835), .ZN(n9839) );
  MUX2_X1 U10029 ( .A(n9837), .B(n8869), .S(n8906), .Z(n8870) );
  MUX2_X1 U10030 ( .A(n8872), .B(n8871), .S(n8912), .Z(n8873) );
  AND2_X1 U10031 ( .A1(n8875), .A2(n8874), .ZN(n8880) );
  INV_X1 U10032 ( .A(n8880), .ZN(n8877) );
  NAND2_X1 U10033 ( .A1(n9955), .A2(n9408), .ZN(n8937) );
  INV_X1 U10034 ( .A(n8937), .ZN(n8876) );
  NAND2_X1 U10035 ( .A1(n8877), .A2(n8876), .ZN(n8879) );
  MUX2_X1 U10036 ( .A(n9408), .B(n9955), .S(n8912), .Z(n8878) );
  AND2_X1 U10037 ( .A1(n8882), .A2(n8881), .ZN(n8884) );
  MUX2_X1 U10038 ( .A(n8884), .B(n8883), .S(n8912), .Z(n8885) );
  INV_X1 U10039 ( .A(n9939), .ZN(n9345) );
  NAND2_X1 U10040 ( .A1(n8887), .A2(n9318), .ZN(n8892) );
  NAND2_X1 U10041 ( .A1(n8892), .A2(n8912), .ZN(n8891) );
  NAND2_X1 U10042 ( .A1(n8889), .A2(n8888), .ZN(n8890) );
  NAND2_X1 U10043 ( .A1(n8891), .A2(n8890), .ZN(n8895) );
  INV_X1 U10044 ( .A(n8892), .ZN(n8893) );
  NAND3_X1 U10045 ( .A1(n8893), .A2(n8912), .A3(n9092), .ZN(n8894) );
  NAND3_X1 U10046 ( .A1(n8898), .A2(n8917), .A3(n8897), .ZN(n8899) );
  MUX2_X1 U10047 ( .A(n8901), .B(n8900), .S(n8906), .Z(n8902) );
  MUX2_X1 U10048 ( .A(n8904), .B(n8903), .S(n8912), .Z(n8905) );
  MUX2_X1 U10049 ( .A(n8908), .B(n8907), .S(n8906), .Z(n8909) );
  INV_X1 U10050 ( .A(n9241), .ZN(n9147) );
  NAND2_X1 U10051 ( .A1(n9907), .A2(n9147), .ZN(n8914) );
  MUX2_X1 U10052 ( .A(n9147), .B(n9907), .S(n8912), .Z(n8913) );
  NOR4_X1 U10053 ( .A1(n8921), .A2(n8920), .A3(n8919), .A4(n6488), .ZN(n8923)
         );
  NAND4_X1 U10054 ( .A1(n8923), .A2(n10768), .A3(n10808), .A4(n8922), .ZN(
        n8924) );
  NOR3_X1 U10055 ( .A1(n8924), .A2(n8252), .A3(n5225), .ZN(n8927) );
  INV_X1 U10056 ( .A(n10931), .ZN(n10936) );
  NAND4_X1 U10057 ( .A1(n8927), .A2(n8926), .A3(n10936), .A4(n8925), .ZN(n8931) );
  NOR4_X1 U10058 ( .A1(n8931), .A2(n8930), .A3(n8929), .A4(n8928), .ZN(n8933)
         );
  NAND4_X1 U10059 ( .A1(n8935), .A2(n8934), .A3(n8933), .A4(n8932), .ZN(n8936)
         );
  NOR4_X1 U10060 ( .A1(n9835), .A2(n9860), .A3(n9869), .A4(n8936), .ZN(n8939)
         );
  NAND2_X1 U10061 ( .A1(n8938), .A2(n8937), .ZN(n9390) );
  NAND4_X1 U10062 ( .A1(n9254), .A2(n8940), .A3(n8939), .A4(n9390), .ZN(n8941)
         );
  NOR4_X1 U10063 ( .A1(n9319), .A2(n8942), .A3(n9349), .A4(n8941), .ZN(n8943)
         );
  XNOR2_X1 U10064 ( .A(n8945), .B(n10902), .ZN(n8946) );
  AOI211_X1 U10065 ( .C1(n6488), .C2(n8948), .A(n8947), .B(n8946), .ZN(n8949)
         );
  INV_X1 U10066 ( .A(n8949), .ZN(n8952) );
  NOR2_X1 U10067 ( .A1(n8954), .A2(n8953), .ZN(n8959) );
  NOR4_X1 U10068 ( .A1(n10547), .A2(n8955), .A3(n7287), .A4(n10937), .ZN(n8957) );
  OAI21_X1 U10069 ( .B1(n8958), .B2(n6947), .A(P2_B_REG_SCAN_IN), .ZN(n8956)
         );
  OAI22_X1 U10070 ( .A1(n8959), .A2(n8958), .B1(n8957), .B2(n8956), .ZN(
        P2_U3244) );
  NAND2_X1 U10071 ( .A1(n10507), .A2(n10165), .ZN(n8960) );
  NAND2_X1 U10072 ( .A1(n10503), .A2(n10164), .ZN(n8961) );
  NAND2_X1 U10073 ( .A1(n10422), .A2(n8961), .ZN(n10404) );
  NAND2_X1 U10074 ( .A1(n10496), .A2(n10163), .ZN(n8962) );
  NAND2_X1 U10075 ( .A1(n10365), .A2(n10369), .ZN(n10367) );
  NAND2_X1 U10076 ( .A1(n10375), .A2(n10161), .ZN(n8963) );
  OR2_X1 U10077 ( .A1(n10481), .A2(n10160), .ZN(n8964) );
  OR2_X1 U10078 ( .A1(n10476), .A2(n10159), .ZN(n8965) );
  NAND2_X1 U10079 ( .A1(n8966), .A2(n8965), .ZN(n10318) );
  OR2_X1 U10080 ( .A1(n10471), .A2(n10158), .ZN(n8967) );
  INV_X1 U10081 ( .A(n10296), .ZN(n8968) );
  OR2_X1 U10082 ( .A1(n10461), .A2(n10126), .ZN(n8969) );
  NAND2_X1 U10083 ( .A1(n8971), .A2(n8992), .ZN(n8972) );
  INV_X1 U10084 ( .A(n10398), .ZN(n8976) );
  NOR2_X1 U10085 ( .A1(n10403), .A2(n8976), .ZN(n8977) );
  NAND2_X1 U10086 ( .A1(n10425), .A2(n8977), .ZN(n8979) );
  NAND2_X1 U10087 ( .A1(n8979), .A2(n8978), .ZN(n10387) );
  NAND2_X1 U10088 ( .A1(n10387), .A2(n10388), .ZN(n8981) );
  INV_X1 U10089 ( .A(n8984), .ZN(n8985) );
  INV_X1 U10090 ( .A(n8986), .ZN(n8987) );
  NAND2_X1 U10091 ( .A1(n10303), .A2(n8989), .ZN(n10295) );
  NAND2_X1 U10092 ( .A1(n8991), .A2(n8992), .ZN(n10271) );
  OAI21_X1 U10093 ( .B1(n8992), .B2(n8991), .A(n10271), .ZN(n8995) );
  OAI22_X1 U10094 ( .A1(n10305), .A2(n10849), .B1(n8993), .B2(n10851), .ZN(
        n8994) );
  INV_X1 U10095 ( .A(n10461), .ZN(n10293) );
  INV_X1 U10096 ( .A(n10481), .ZN(n10355) );
  INV_X1 U10097 ( .A(n10503), .ZN(n10435) );
  INV_X1 U10098 ( .A(n10496), .ZN(n10414) );
  NAND2_X1 U10099 ( .A1(n10347), .A2(n10352), .ZN(n10334) );
  AOI21_X1 U10100 ( .B1(n10455), .B2(n10288), .A(n10256), .ZN(n10456) );
  INV_X1 U10101 ( .A(n10455), .ZN(n10269) );
  AOI22_X1 U10102 ( .A1(n8997), .A2(n11025), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n11027), .ZN(n8998) );
  OAI21_X1 U10103 ( .B1(n10269), .B2(n11029), .A(n8998), .ZN(n9000) );
  NOR2_X1 U10104 ( .A1(n10459), .A2(n10419), .ZN(n8999) );
  AOI211_X1 U10105 ( .C1(n11022), .C2(n10456), .A(n9000), .B(n8999), .ZN(n9001) );
  OAI21_X1 U10106 ( .B1(n10458), .B2(n11027), .A(n9001), .ZN(P1_U3263) );
  INV_X1 U10107 ( .A(n9002), .ZN(n10013) );
  OAI222_X1 U10108 ( .A1(n9004), .A2(n9003), .B1(n5033), .B2(n10013), .C1(
        P1_U3084), .C2(n5036), .ZN(P1_U3325) );
  INV_X1 U10109 ( .A(n9005), .ZN(n9006) );
  AOI21_X1 U10110 ( .B1(n9136), .B2(n9006), .A(n9086), .ZN(n9010) );
  NOR3_X1 U10111 ( .A1(n9007), .A2(n9308), .A3(n9122), .ZN(n9009) );
  OAI21_X1 U10112 ( .B1(n9010), .B2(n9009), .A(n9008), .ZN(n9015) );
  OAI22_X1 U10113 ( .A1(n9308), .A2(n9104), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9011), .ZN(n9013) );
  NOR2_X1 U10114 ( .A1(n9309), .A2(n9127), .ZN(n9012) );
  AOI211_X1 U10115 ( .C1(n9129), .C2(n9303), .A(n9013), .B(n9012), .ZN(n9014)
         );
  OAI211_X1 U10116 ( .C1(n9305), .C2(n9146), .A(n9015), .B(n9014), .ZN(
        P2_U3216) );
  NAND2_X1 U10117 ( .A1(n9017), .A2(n9016), .ZN(n9024) );
  NAND2_X1 U10118 ( .A1(n9018), .A2(n9135), .ZN(n9023) );
  NAND3_X1 U10119 ( .A1(n9024), .A2(n9093), .A3(n9148), .ZN(n9022) );
  OAI22_X1 U10120 ( .A1(n9104), .A2(n9065), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9473), .ZN(n9020) );
  OAI22_X1 U10121 ( .A1(n9364), .A2(n9141), .B1(n9092), .B2(n9127), .ZN(n9019)
         );
  AOI211_X1 U10122 ( .C1(n9945), .C2(n9098), .A(n9020), .B(n9019), .ZN(n9021)
         );
  OAI211_X1 U10123 ( .C1(n9024), .C2(n9023), .A(n9022), .B(n9021), .ZN(
        P2_U3218) );
  INV_X1 U10124 ( .A(n9025), .ZN(n9034) );
  INV_X1 U10125 ( .A(n9026), .ZN(n9029) );
  AOI21_X1 U10126 ( .B1(n9029), .B2(n9028), .A(n9027), .ZN(n9030) );
  AOI21_X1 U10127 ( .B1(n9034), .B2(n9031), .A(n9030), .ZN(n9037) );
  NAND2_X1 U10128 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9235) );
  OAI21_X1 U10129 ( .B1(n9104), .B2(n9876), .A(n9235), .ZN(n9033) );
  OAI22_X1 U10130 ( .A1(n9141), .A2(n9848), .B1(n9842), .B2(n9127), .ZN(n9032)
         );
  AOI211_X1 U10131 ( .C1(n9967), .C2(n9098), .A(n9033), .B(n9032), .ZN(n9036)
         );
  NAND3_X1 U10132 ( .A1(n9034), .A2(n9093), .A3(n9863), .ZN(n9035) );
  OAI211_X1 U10133 ( .C1(n9037), .C2(n9086), .A(n9036), .B(n9035), .ZN(
        P2_U3221) );
  AOI21_X1 U10134 ( .B1(n9038), .B2(n5127), .A(n9086), .ZN(n9041) );
  NOR3_X1 U10135 ( .A1(n9122), .A2(n9042), .A3(n9039), .ZN(n9040) );
  OAI21_X1 U10136 ( .B1(n9041), .B2(n9040), .A(n8135), .ZN(n9046) );
  OAI22_X1 U10137 ( .A1(n9042), .A2(n10937), .B1(n10938), .B2(n10939), .ZN(
        n10896) );
  AOI22_X1 U10138 ( .A1(n9143), .A2(n10896), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n9045) );
  NAND2_X1 U10139 ( .A1(n9098), .A2(n10898), .ZN(n9044) );
  NAND2_X1 U10140 ( .A1(n9129), .A2(n10900), .ZN(n9043) );
  NAND4_X1 U10141 ( .A1(n9046), .A2(n9045), .A3(n9044), .A4(n9043), .ZN(
        P2_U3223) );
  OR3_X1 U10142 ( .A1(n9122), .A2(n9053), .A3(n8191), .ZN(n9058) );
  NOR2_X1 U10143 ( .A1(n9047), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10659) );
  AOI21_X1 U10144 ( .B1(n9143), .B2(n9048), .A(n10659), .ZN(n9057) );
  AOI22_X1 U10145 ( .A1(n9098), .A2(n9050), .B1(n9049), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n9056) );
  OAI21_X1 U10146 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(n9054) );
  NAND2_X1 U10147 ( .A1(n9054), .A2(n9135), .ZN(n9055) );
  NAND4_X1 U10148 ( .A1(n9058), .A2(n9057), .A3(n9056), .A4(n9055), .ZN(
        P2_U3224) );
  INV_X1 U10149 ( .A(n9059), .ZN(n9060) );
  AOI21_X1 U10150 ( .B1(n9102), .B2(n9060), .A(n9086), .ZN(n9064) );
  NOR3_X1 U10151 ( .A1(n9061), .A2(n9842), .A3(n9122), .ZN(n9063) );
  OAI21_X1 U10152 ( .B1(n9064), .B2(n9063), .A(n9062), .ZN(n9069) );
  OAI22_X1 U10153 ( .A1(n9127), .A2(n9065), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9681), .ZN(n9067) );
  OAI22_X1 U10154 ( .A1(n9141), .A2(n9386), .B1(n9842), .B2(n9104), .ZN(n9066)
         );
  AOI211_X1 U10155 ( .C1(n9955), .C2(n9098), .A(n9067), .B(n9066), .ZN(n9068)
         );
  NAND2_X1 U10156 ( .A1(n9069), .A2(n9068), .ZN(P2_U3225) );
  INV_X1 U10157 ( .A(n9070), .ZN(n9073) );
  XNOR2_X1 U10158 ( .A(n9072), .B(n9070), .ZN(n9094) );
  NAND2_X1 U10159 ( .A1(n9094), .A2(n9071), .ZN(n9095) );
  OAI21_X1 U10160 ( .B1(n9073), .B2(n9072), .A(n9095), .ZN(n9077) );
  XNOR2_X1 U10161 ( .A(n9075), .B(n9074), .ZN(n9076) );
  XNOR2_X1 U10162 ( .A(n9077), .B(n9076), .ZN(n9083) );
  NOR2_X1 U10163 ( .A1(n9092), .A2(n10937), .ZN(n9078) );
  AOI21_X1 U10164 ( .B1(n9260), .B2(n9890), .A(n9078), .ZN(n9332) );
  AOI22_X1 U10165 ( .A1(n9334), .A2(n9129), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n9079) );
  OAI21_X1 U10166 ( .B1(n9332), .B2(n9080), .A(n9079), .ZN(n9081) );
  AOI21_X1 U10167 ( .B1(n9936), .B2(n9098), .A(n9081), .ZN(n9082) );
  OAI21_X1 U10168 ( .B1(n9083), .B2(n9086), .A(n9082), .ZN(P2_U3227) );
  AOI22_X1 U10169 ( .A1(n9125), .A2(n9248), .B1(n9129), .B2(n9881), .ZN(n9084)
         );
  NAND2_X1 U10170 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9206) );
  OAI211_X1 U10171 ( .C1(n9876), .C2(n9127), .A(n9084), .B(n9206), .ZN(n9090)
         );
  INV_X1 U10172 ( .A(n9121), .ZN(n9085) );
  AOI211_X1 U10173 ( .C1(n9088), .C2(n9087), .A(n9086), .B(n9085), .ZN(n9089)
         );
  AOI211_X1 U10174 ( .C1(n9977), .C2(n9098), .A(n9090), .B(n9089), .ZN(n9091)
         );
  INV_X1 U10175 ( .A(n9091), .ZN(P2_U3230) );
  AOI22_X1 U10176 ( .A1(n9094), .A2(n9135), .B1(n9093), .B2(n9357), .ZN(n9101)
         );
  INV_X1 U10177 ( .A(n9095), .ZN(n9100) );
  OAI22_X1 U10178 ( .A1(n9350), .A2(n9127), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9692), .ZN(n9097) );
  OAI22_X1 U10179 ( .A1(n9141), .A2(n9342), .B1(n9378), .B2(n9104), .ZN(n9096)
         );
  AOI211_X1 U10180 ( .C1(n9939), .C2(n9098), .A(n9097), .B(n9096), .ZN(n9099)
         );
  OAI21_X1 U10181 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(P2_U3231) );
  INV_X1 U10182 ( .A(n9960), .ZN(n9405) );
  OAI211_X1 U10183 ( .C1(n9103), .C2(n9025), .A(n9102), .B(n9135), .ZN(n9108)
         );
  NOR2_X1 U10184 ( .A1(n9127), .A2(n9377), .ZN(n9106) );
  OAI22_X1 U10185 ( .A1(n9141), .A2(n9402), .B1(n9251), .B2(n9104), .ZN(n9105)
         );
  AOI211_X1 U10186 ( .C1(P2_REG3_REG_20__SCAN_IN), .C2(P2_U3152), .A(n9106), 
        .B(n9105), .ZN(n9107) );
  OAI211_X1 U10187 ( .C1(n9405), .C2(n9146), .A(n9108), .B(n9107), .ZN(
        P2_U3235) );
  OAI21_X1 U10188 ( .B1(n9111), .B2(n9062), .A(n9109), .ZN(n9118) );
  INV_X1 U10189 ( .A(n9950), .ZN(n9375) );
  NOR3_X1 U10190 ( .A1(n9111), .A2(n9110), .A3(n9122), .ZN(n9112) );
  OAI21_X1 U10191 ( .B1(n9112), .B2(n9125), .A(n9408), .ZN(n9116) );
  OAI22_X1 U10192 ( .A1(n9378), .A2(n9127), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9113), .ZN(n9114) );
  AOI21_X1 U10193 ( .B1(n9373), .B2(n9129), .A(n9114), .ZN(n9115) );
  OAI211_X1 U10194 ( .C1(n9375), .C2(n9146), .A(n9116), .B(n9115), .ZN(n9117)
         );
  AOI21_X1 U10195 ( .B1(n9118), .B2(n9135), .A(n9117), .ZN(n9119) );
  INV_X1 U10196 ( .A(n9119), .ZN(P2_U3237) );
  OAI21_X1 U10197 ( .B1(n9124), .B2(n9121), .A(n9120), .ZN(n9133) );
  NOR3_X1 U10198 ( .A1(n9124), .A2(n9123), .A3(n9122), .ZN(n9126) );
  OAI21_X1 U10199 ( .B1(n9126), .B2(n9125), .A(n9862), .ZN(n9131) );
  NAND2_X1 U10200 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9215) );
  OAI21_X1 U10201 ( .B1(n9127), .B2(n9251), .A(n9215), .ZN(n9128) );
  AOI21_X1 U10202 ( .B1(n9857), .B2(n9129), .A(n9128), .ZN(n9130) );
  OAI211_X1 U10203 ( .C1(n9859), .C2(n9146), .A(n9131), .B(n9130), .ZN(n9132)
         );
  AOI21_X1 U10204 ( .B1(n9133), .B2(n9135), .A(n9132), .ZN(n9134) );
  INV_X1 U10205 ( .A(n9134), .ZN(P2_U3240) );
  OAI211_X1 U10206 ( .C1(n9138), .C2(n9137), .A(n9136), .B(n9135), .ZN(n9145)
         );
  OR2_X1 U10207 ( .A1(n9262), .A2(n10939), .ZN(n9140) );
  OR2_X1 U10208 ( .A1(n9350), .A2(n10937), .ZN(n9139) );
  NAND2_X1 U10209 ( .A1(n9140), .A2(n9139), .ZN(n9321) );
  OAI22_X1 U10210 ( .A1(n9325), .A2(n9141), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9713), .ZN(n9142) );
  AOI21_X1 U10211 ( .B1(n9321), .B2(n9143), .A(n9142), .ZN(n9144) );
  OAI211_X1 U10212 ( .C1(n9238), .C2(n9146), .A(n9145), .B(n9144), .ZN(
        P2_U3242) );
  MUX2_X1 U10213 ( .A(n9147), .B(P2_DATAO_REG_31__SCAN_IN), .S(n9160), .Z(
        P2_U3583) );
  MUX2_X1 U10214 ( .A(n9292), .B(P2_DATAO_REG_29__SCAN_IN), .S(n9160), .Z(
        P2_U3581) );
  INV_X1 U10215 ( .A(n9309), .ZN(n9263) );
  MUX2_X1 U10216 ( .A(n9263), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9160), .Z(
        P2_U3580) );
  INV_X1 U10217 ( .A(n9262), .ZN(n9293) );
  MUX2_X1 U10218 ( .A(n9293), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9160), .Z(
        P2_U3579) );
  MUX2_X1 U10219 ( .A(n9260), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9160), .Z(
        P2_U3578) );
  INV_X1 U10220 ( .A(n9350), .ZN(n9258) );
  MUX2_X1 U10221 ( .A(n9258), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9160), .Z(
        P2_U3577) );
  MUX2_X1 U10222 ( .A(n9357), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9160), .Z(
        P2_U3576) );
  MUX2_X1 U10223 ( .A(n9148), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9160), .Z(
        P2_U3575) );
  MUX2_X1 U10224 ( .A(n9393), .B(P2_DATAO_REG_22__SCAN_IN), .S(n9160), .Z(
        P2_U3574) );
  MUX2_X1 U10225 ( .A(n9408), .B(P2_DATAO_REG_21__SCAN_IN), .S(n9160), .Z(
        P2_U3573) );
  INV_X1 U10226 ( .A(n9842), .ZN(n9394) );
  MUX2_X1 U10227 ( .A(n9394), .B(P2_DATAO_REG_20__SCAN_IN), .S(n9160), .Z(
        P2_U3572) );
  MUX2_X1 U10228 ( .A(n9863), .B(P2_DATAO_REG_19__SCAN_IN), .S(n9160), .Z(
        P2_U3571) );
  MUX2_X1 U10229 ( .A(n9862), .B(P2_DATAO_REG_17__SCAN_IN), .S(n9160), .Z(
        P2_U3569) );
  MUX2_X1 U10230 ( .A(n9248), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9160), .Z(
        P2_U3568) );
  MUX2_X1 U10231 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9149), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10232 ( .A(n9150), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9160), .Z(
        P2_U3566) );
  MUX2_X1 U10233 ( .A(n9151), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9160), .Z(
        P2_U3565) );
  MUX2_X1 U10234 ( .A(n9152), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9160), .Z(
        P2_U3564) );
  MUX2_X1 U10235 ( .A(n9153), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9160), .Z(
        P2_U3563) );
  MUX2_X1 U10236 ( .A(n9154), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9160), .Z(
        P2_U3562) );
  MUX2_X1 U10237 ( .A(n9155), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9160), .Z(
        P2_U3561) );
  MUX2_X1 U10238 ( .A(n9156), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9160), .Z(
        P2_U3560) );
  MUX2_X1 U10239 ( .A(n9891), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9160), .Z(
        P2_U3559) );
  MUX2_X1 U10240 ( .A(n9157), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9160), .Z(
        P2_U3558) );
  MUX2_X1 U10241 ( .A(n9893), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9160), .Z(
        P2_U3557) );
  MUX2_X1 U10242 ( .A(n8242), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9160), .Z(
        P2_U3555) );
  MUX2_X1 U10243 ( .A(n9158), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9160), .Z(
        P2_U3554) );
  MUX2_X1 U10244 ( .A(n9159), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9160), .Z(
        P2_U3553) );
  MUX2_X1 U10245 ( .A(n9161), .B(P2_DATAO_REG_0__SCAN_IN), .S(n9160), .Z(
        P2_U3552) );
  OAI21_X1 U10246 ( .B1(n9217), .B2(n9163), .A(n9162), .ZN(n9167) );
  OAI21_X1 U10247 ( .B1(n9170), .B2(P2_REG1_REG_14__SCAN_IN), .A(n9164), .ZN(
        n9177) );
  XNOR2_X1 U10248 ( .A(n9187), .B(n9177), .ZN(n9165) );
  INV_X1 U10249 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11077) );
  NOR2_X1 U10250 ( .A1(n11077), .A2(n9165), .ZN(n9178) );
  AOI211_X1 U10251 ( .C1(n9165), .C2(n11077), .A(n9178), .B(n10673), .ZN(n9166) );
  AOI211_X1 U10252 ( .C1(n10684), .C2(n9168), .A(n9167), .B(n9166), .ZN(n9176)
         );
  OAI21_X1 U10253 ( .B1(n9170), .B2(P2_REG2_REG_14__SCAN_IN), .A(n9169), .ZN(
        n9186) );
  INV_X1 U10254 ( .A(n9186), .ZN(n9171) );
  XNOR2_X1 U10255 ( .A(n9187), .B(n9171), .ZN(n9173) );
  INV_X1 U10256 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U10257 ( .A1(n9173), .A2(n9172), .ZN(n9188) );
  OAI21_X1 U10258 ( .B1(n9173), .B2(n9172), .A(n9188), .ZN(n9174) );
  NAND2_X1 U10259 ( .A1(n10651), .A2(n9174), .ZN(n9175) );
  NAND2_X1 U10260 ( .A1(n9176), .A2(n9175), .ZN(P2_U3260) );
  NOR2_X1 U10261 ( .A1(n9187), .A2(n9177), .ZN(n9179) );
  NOR2_X1 U10262 ( .A1(n9179), .A2(n9178), .ZN(n9182) );
  INV_X1 U10263 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9180) );
  AOI22_X1 U10264 ( .A1(n9202), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9180), .B2(
        n9185), .ZN(n9181) );
  NAND2_X1 U10265 ( .A1(n9182), .A2(n9181), .ZN(n9198) );
  OAI21_X1 U10266 ( .B1(n9182), .B2(n9181), .A(n9198), .ZN(n9196) );
  NAND2_X1 U10267 ( .A1(n10672), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n9183) );
  OAI211_X1 U10268 ( .C1(n10653), .C2(n9185), .A(n9184), .B(n9183), .ZN(n9195)
         );
  NAND2_X1 U10269 ( .A1(n9187), .A2(n9186), .ZN(n9189) );
  NAND2_X1 U10270 ( .A1(n9189), .A2(n9188), .ZN(n9193) );
  INV_X1 U10271 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9190) );
  MUX2_X1 U10272 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n9190), .S(n9202), .Z(n9191) );
  INV_X1 U10273 ( .A(n9191), .ZN(n9192) );
  NOR2_X1 U10274 ( .A1(n9193), .A2(n9192), .ZN(n9201) );
  AOI211_X1 U10275 ( .C1(n9193), .C2(n9192), .A(n9201), .B(n10677), .ZN(n9194)
         );
  AOI211_X1 U10276 ( .C1(n9196), .C2(n10649), .A(n9195), .B(n9194), .ZN(n9197)
         );
  INV_X1 U10277 ( .A(n9197), .ZN(P2_U3261) );
  OAI21_X1 U10278 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n9202), .A(n9198), .ZN(
        n9200) );
  XNOR2_X1 U10279 ( .A(n9221), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9199) );
  NOR2_X1 U10280 ( .A1(n9199), .A2(n9200), .ZN(n9212) );
  AOI211_X1 U10281 ( .C1(n9200), .C2(n9199), .A(n9212), .B(n10673), .ZN(n9211)
         );
  AOI21_X1 U10282 ( .B1(n9202), .B2(P2_REG2_REG_16__SCAN_IN), .A(n9201), .ZN(
        n9205) );
  NAND2_X1 U10283 ( .A1(n9221), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n9203) );
  OAI21_X1 U10284 ( .B1(n9221), .B2(P2_REG2_REG_17__SCAN_IN), .A(n9203), .ZN(
        n9204) );
  NOR2_X1 U10285 ( .A1(n9205), .A2(n9204), .ZN(n9220) );
  AOI211_X1 U10286 ( .C1(n9205), .C2(n9204), .A(n9220), .B(n10677), .ZN(n9210)
         );
  NAND2_X1 U10287 ( .A1(n10684), .A2(n9221), .ZN(n9207) );
  OAI211_X1 U10288 ( .C1(n9208), .C2(n9217), .A(n9207), .B(n9206), .ZN(n9209)
         );
  OR3_X1 U10289 ( .A1(n9211), .A2(n9210), .A3(n9209), .ZN(P2_U3262) );
  INV_X1 U10290 ( .A(n9232), .ZN(n9227) );
  XOR2_X1 U10291 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9232), .Z(n9214) );
  AOI21_X1 U10292 ( .B1(n9221), .B2(P2_REG1_REG_17__SCAN_IN), .A(n9212), .ZN(
        n9213) );
  NAND2_X1 U10293 ( .A1(n9214), .A2(n9213), .ZN(n9231) );
  OAI21_X1 U10294 ( .B1(n9214), .B2(n9213), .A(n9231), .ZN(n9219) );
  INV_X1 U10295 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9216) );
  OAI21_X1 U10296 ( .B1(n9217), .B2(n9216), .A(n9215), .ZN(n9218) );
  AOI21_X1 U10297 ( .B1(n10649), .B2(n9219), .A(n9218), .ZN(n9226) );
  XOR2_X1 U10298 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n9232), .Z(n9223) );
  AOI21_X1 U10299 ( .B1(n9221), .B2(P2_REG2_REG_17__SCAN_IN), .A(n9220), .ZN(
        n9222) );
  NAND2_X1 U10300 ( .A1(n9223), .A2(n9222), .ZN(n9228) );
  OAI21_X1 U10301 ( .B1(n9223), .B2(n9222), .A(n9228), .ZN(n9224) );
  NAND2_X1 U10302 ( .A1(n10651), .A2(n9224), .ZN(n9225) );
  OAI211_X1 U10303 ( .C1(n10653), .C2(n9227), .A(n9226), .B(n9225), .ZN(
        P2_U3263) );
  OAI21_X1 U10304 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n9232), .A(n9228), .ZN(
        n9230) );
  MUX2_X1 U10305 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n6777), .S(n9846), .Z(n9229) );
  XNOR2_X1 U10306 ( .A(n9230), .B(n9229), .ZN(n9237) );
  NAND2_X1 U10307 ( .A1(n10672), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9234) );
  OAI21_X1 U10308 ( .B1(n9237), .B2(n10677), .A(n9236), .ZN(P2_U3264) );
  INV_X1 U10309 ( .A(n9967), .ZN(n9843) );
  NAND2_X1 U10310 ( .A1(n9367), .A2(n9372), .ZN(n9362) );
  NAND2_X1 U10311 ( .A1(n9279), .A2(n9285), .ZN(n9276) );
  XNOR2_X1 U10312 ( .A(n9907), .B(n9911), .ZN(n9909) );
  NAND2_X1 U10313 ( .A1(n9239), .A2(P2_B_REG_SCAN_IN), .ZN(n9240) );
  NAND2_X1 U10314 ( .A1(n9890), .A2(n9240), .ZN(n9272) );
  NOR2_X1 U10315 ( .A1(n9241), .A2(n9272), .ZN(n9906) );
  INV_X1 U10316 ( .A(n9906), .ZN(n9912) );
  NOR2_X1 U10317 ( .A1(n10906), .A2(n9912), .ZN(n9245) );
  AOI21_X1 U10318 ( .B1(n10906), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9245), .ZN(
        n9243) );
  NAND2_X1 U10319 ( .A1(n9907), .A2(n9901), .ZN(n9242) );
  OAI211_X1 U10320 ( .C1(n9909), .C2(n10952), .A(n9243), .B(n9242), .ZN(
        P2_U3265) );
  NAND2_X1 U10321 ( .A1(n9244), .A2(n9276), .ZN(n9910) );
  NAND3_X1 U10322 ( .A1(n9911), .A2(n9910), .A3(n9897), .ZN(n9247) );
  AOI21_X1 U10323 ( .B1(n10906), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9245), .ZN(
        n9246) );
  OAI211_X1 U10324 ( .C1(n9914), .C2(n10956), .A(n9247), .B(n9246), .ZN(
        P2_U3266) );
  INV_X1 U10325 ( .A(n9252), .ZN(n9253) );
  OAI22_X1 U10326 ( .A1(n9371), .A2(n9254), .B1(n9393), .B2(n9950), .ZN(n9361)
         );
  NOR2_X1 U10327 ( .A1(n9367), .A2(n9378), .ZN(n9255) );
  NAND2_X1 U10328 ( .A1(n9238), .A2(n9308), .ZN(n9261) );
  NOR2_X1 U10329 ( .A1(n9919), .A2(n9263), .ZN(n9264) );
  AOI21_X1 U10330 ( .B1(n9284), .B2(n9265), .A(n9264), .ZN(n9266) );
  XNOR2_X1 U10331 ( .A(n9266), .B(n9267), .ZN(n9915) );
  INV_X1 U10332 ( .A(n9915), .ZN(n9283) );
  INV_X1 U10333 ( .A(n9267), .ZN(n9268) );
  XNOR2_X1 U10334 ( .A(n9269), .B(n9268), .ZN(n9270) );
  NAND2_X1 U10335 ( .A1(n9270), .A2(n10942), .ZN(n9275) );
  OAI22_X1 U10336 ( .A1(n9309), .A2(n10937), .B1(n9272), .B2(n9271), .ZN(n9273) );
  INV_X1 U10337 ( .A(n9273), .ZN(n9274) );
  NAND2_X1 U10338 ( .A1(n9275), .A2(n9274), .ZN(n9917) );
  NOR2_X1 U10339 ( .A1(n9916), .A2(n10952), .ZN(n9281) );
  AOI22_X1 U10340 ( .A1(n9277), .A2(n10962), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n10906), .ZN(n9278) );
  OAI21_X1 U10341 ( .B1(n9279), .B2(n10956), .A(n9278), .ZN(n9280) );
  AOI211_X1 U10342 ( .C1(n9917), .C2(n10957), .A(n9281), .B(n9280), .ZN(n9282)
         );
  OAI21_X1 U10343 ( .B1(n9283), .B2(n9887), .A(n9282), .ZN(P2_U3267) );
  XNOR2_X1 U10344 ( .A(n9284), .B(n9290), .ZN(n9923) );
  AOI21_X1 U10345 ( .B1(n9919), .B2(n9300), .A(n9285), .ZN(n9920) );
  INV_X1 U10346 ( .A(n9919), .ZN(n9288) );
  AOI22_X1 U10347 ( .A1(n9286), .A2(n10962), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n10906), .ZN(n9287) );
  OAI21_X1 U10348 ( .B1(n9288), .B2(n10956), .A(n9287), .ZN(n9297) );
  OAI211_X1 U10349 ( .C1(n9291), .C2(n9290), .A(n9289), .B(n10942), .ZN(n9295)
         );
  AOI22_X1 U10350 ( .A1(n9293), .A2(n9892), .B1(n9890), .B2(n9292), .ZN(n9294)
         );
  NOR2_X1 U10351 ( .A1(n9922), .A2(n10906), .ZN(n9296) );
  AOI211_X1 U10352 ( .C1(n9897), .C2(n9920), .A(n9297), .B(n9296), .ZN(n9298)
         );
  OAI21_X1 U10353 ( .B1(n9923), .B2(n9887), .A(n9298), .ZN(P2_U3268) );
  XOR2_X1 U10354 ( .A(n9307), .B(n9299), .Z(n9928) );
  INV_X1 U10355 ( .A(n9323), .ZN(n9302) );
  INV_X1 U10356 ( .A(n9300), .ZN(n9301) );
  AOI21_X1 U10357 ( .B1(n9924), .B2(n9302), .A(n9301), .ZN(n9925) );
  AOI22_X1 U10358 ( .A1(n9303), .A2(n10962), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10906), .ZN(n9304) );
  OAI21_X1 U10359 ( .B1(n9305), .B2(n10956), .A(n9304), .ZN(n9314) );
  AOI21_X1 U10360 ( .B1(n9306), .B2(n9307), .A(n10811), .ZN(n9312) );
  OAI22_X1 U10361 ( .A1(n9309), .A2(n10939), .B1(n9308), .B2(n10937), .ZN(
        n9310) );
  AOI21_X1 U10362 ( .B1(n9312), .B2(n9311), .A(n9310), .ZN(n9927) );
  NOR2_X1 U10363 ( .A1(n9927), .A2(n10906), .ZN(n9313) );
  AOI211_X1 U10364 ( .C1(n9897), .C2(n9925), .A(n9314), .B(n9313), .ZN(n9315)
         );
  OAI21_X1 U10365 ( .B1(n9928), .B2(n9887), .A(n9315), .ZN(P2_U3269) );
  XOR2_X1 U10366 ( .A(n9319), .B(n9316), .Z(n9933) );
  AOI22_X1 U10367 ( .A1(n9930), .A2(n9901), .B1(n10906), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U10368 ( .A1(n9317), .A2(n9318), .ZN(n9320) );
  XNOR2_X1 U10369 ( .A(n9320), .B(n9319), .ZN(n9322) );
  AOI21_X1 U10370 ( .B1(n9322), .B2(n10942), .A(n9321), .ZN(n9932) );
  AOI211_X1 U10371 ( .C1(n9930), .C2(n5347), .A(n11070), .B(n9323), .ZN(n9929)
         );
  NAND2_X1 U10372 ( .A1(n9929), .A2(n9846), .ZN(n9324) );
  OAI211_X1 U10373 ( .C1(n9849), .C2(n9325), .A(n9932), .B(n9324), .ZN(n9326)
         );
  NAND2_X1 U10374 ( .A1(n9326), .A2(n10957), .ZN(n9327) );
  OAI211_X1 U10375 ( .C1(n9933), .C2(n9887), .A(n9328), .B(n9327), .ZN(
        P2_U3270) );
  XNOR2_X1 U10376 ( .A(n9329), .B(n9331), .ZN(n9938) );
  OAI211_X1 U10377 ( .C1(n9331), .C2(n9330), .A(n9317), .B(n10942), .ZN(n9333)
         );
  NAND2_X1 U10378 ( .A1(n9333), .A2(n9332), .ZN(n9934) );
  AOI211_X1 U10379 ( .C1(n9936), .C2(n5110), .A(n11070), .B(n5345), .ZN(n9935)
         );
  NAND2_X1 U10380 ( .A1(n9935), .A2(n9880), .ZN(n9336) );
  AOI22_X1 U10381 ( .A1(n10906), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n9334), 
        .B2(n10962), .ZN(n9335) );
  OAI211_X1 U10382 ( .C1(n5346), .C2(n10956), .A(n9336), .B(n9335), .ZN(n9337)
         );
  AOI21_X1 U10383 ( .B1(n9934), .B2(n10957), .A(n9337), .ZN(n9338) );
  OAI21_X1 U10384 ( .B1(n9938), .B2(n9887), .A(n9338), .ZN(P2_U3271) );
  OAI21_X1 U10385 ( .B1(n9340), .B2(n9349), .A(n9339), .ZN(n9341) );
  INV_X1 U10386 ( .A(n9341), .ZN(n9943) );
  XNOR2_X1 U10387 ( .A(n9345), .B(n9362), .ZN(n9940) );
  INV_X1 U10388 ( .A(n9342), .ZN(n9343) );
  AOI22_X1 U10389 ( .A1(n10906), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9343), 
        .B2(n10962), .ZN(n9344) );
  OAI21_X1 U10390 ( .B1(n9345), .B2(n10956), .A(n9344), .ZN(n9354) );
  NAND2_X1 U10391 ( .A1(n9356), .A2(n9346), .ZN(n9348) );
  AOI211_X1 U10392 ( .C1(n9349), .C2(n9348), .A(n10811), .B(n5145), .ZN(n9352)
         );
  OAI22_X1 U10393 ( .A1(n9350), .A2(n10939), .B1(n9378), .B2(n10937), .ZN(
        n9351) );
  NOR2_X1 U10394 ( .A1(n9352), .A2(n9351), .ZN(n9942) );
  NOR2_X1 U10395 ( .A1(n9942), .A2(n10906), .ZN(n9353) );
  AOI211_X1 U10396 ( .C1(n9940), .C2(n9897), .A(n9354), .B(n9353), .ZN(n9355)
         );
  OAI21_X1 U10397 ( .B1(n9943), .B2(n9887), .A(n9355), .ZN(P2_U3272) );
  OAI21_X1 U10398 ( .B1(n5066), .B2(n9360), .A(n9356), .ZN(n9358) );
  AOI222_X1 U10399 ( .A1(n10942), .A2(n9358), .B1(n9357), .B2(n9890), .C1(
        n9393), .C2(n9892), .ZN(n9948) );
  NAND2_X1 U10400 ( .A1(n9361), .A2(n9360), .ZN(n9944) );
  NAND3_X1 U10401 ( .A1(n5594), .A2(n10790), .A3(n9944), .ZN(n9370) );
  INV_X1 U10402 ( .A(n9372), .ZN(n9363) );
  AOI21_X1 U10403 ( .B1(n9945), .B2(n9363), .A(n5341), .ZN(n9946) );
  INV_X1 U10404 ( .A(n9364), .ZN(n9365) );
  AOI22_X1 U10405 ( .A1(n10906), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9365), 
        .B2(n10962), .ZN(n9366) );
  OAI21_X1 U10406 ( .B1(n9367), .B2(n10956), .A(n9366), .ZN(n9368) );
  AOI21_X1 U10407 ( .B1(n9946), .B2(n9897), .A(n9368), .ZN(n9369) );
  OAI211_X1 U10408 ( .C1(n10906), .C2(n9948), .A(n9370), .B(n9369), .ZN(
        P2_U3273) );
  XNOR2_X1 U10409 ( .A(n9371), .B(n5244), .ZN(n9954) );
  AOI21_X1 U10410 ( .B1(n9950), .B2(n5113), .A(n9372), .ZN(n9951) );
  AOI22_X1 U10411 ( .A1(n10906), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9373), 
        .B2(n10962), .ZN(n9374) );
  OAI21_X1 U10412 ( .B1(n9375), .B2(n10956), .A(n9374), .ZN(n9383) );
  AOI21_X1 U10413 ( .B1(n9376), .B2(n5244), .A(n10811), .ZN(n9381) );
  OAI22_X1 U10414 ( .A1(n9378), .A2(n10939), .B1(n9377), .B2(n10937), .ZN(
        n9379) );
  AOI21_X1 U10415 ( .B1(n9381), .B2(n9380), .A(n9379), .ZN(n9953) );
  NOR2_X1 U10416 ( .A1(n9953), .A2(n10906), .ZN(n9382) );
  AOI211_X1 U10417 ( .C1(n9951), .C2(n9897), .A(n9383), .B(n9382), .ZN(n9384)
         );
  OAI21_X1 U10418 ( .B1(n9954), .B2(n9887), .A(n9384), .ZN(P2_U3274) );
  AOI21_X1 U10419 ( .B1(n9390), .B2(n9385), .A(n5114), .ZN(n9959) );
  XOR2_X1 U10420 ( .A(n9955), .B(n9400), .Z(n9956) );
  INV_X1 U10421 ( .A(n9955), .ZN(n9389) );
  INV_X1 U10422 ( .A(n9386), .ZN(n9387) );
  AOI22_X1 U10423 ( .A1(n10906), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9387), 
        .B2(n10962), .ZN(n9388) );
  OAI21_X1 U10424 ( .B1(n9389), .B2(n10956), .A(n9388), .ZN(n9396) );
  XOR2_X1 U10425 ( .A(n9391), .B(n9390), .Z(n9392) );
  AOI222_X1 U10426 ( .A1(n9394), .A2(n9892), .B1(n9393), .B2(n9890), .C1(
        n10942), .C2(n9392), .ZN(n9958) );
  NOR2_X1 U10427 ( .A1(n9958), .A2(n10906), .ZN(n9395) );
  AOI211_X1 U10428 ( .C1(n9956), .C2(n9897), .A(n9396), .B(n9395), .ZN(n9397)
         );
  OAI21_X1 U10429 ( .B1(n9959), .B2(n9887), .A(n9397), .ZN(P2_U3275) );
  OAI21_X1 U10430 ( .B1(n9399), .B2(n9406), .A(n9398), .ZN(n9964) );
  INV_X1 U10431 ( .A(n9400), .ZN(n9401) );
  AOI21_X1 U10432 ( .B1(n9960), .B2(n9845), .A(n9401), .ZN(n9961) );
  INV_X1 U10433 ( .A(n9402), .ZN(n9403) );
  AOI22_X1 U10434 ( .A1(n10906), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9403), 
        .B2(n10962), .ZN(n9404) );
  OAI21_X1 U10435 ( .B1(n9405), .B2(n10956), .A(n9404), .ZN(n9411) );
  XNOR2_X1 U10436 ( .A(n9407), .B(n9406), .ZN(n9409) );
  AOI222_X1 U10437 ( .A1(n10942), .A2(n9409), .B1(n9408), .B2(n9890), .C1(
        n9863), .C2(n9892), .ZN(n9963) );
  NOR2_X1 U10438 ( .A1(n9963), .A2(n10906), .ZN(n9410) );
  AOI211_X1 U10439 ( .C1(n9961), .C2(n9897), .A(n9411), .B(n9410), .ZN(n9412)
         );
  OAI21_X1 U10440 ( .B1(n9964), .B2(n9887), .A(n9412), .ZN(n9833) );
  XOR2_X1 U10441 ( .A(SI_31_), .B(keyinput_1), .Z(n9417) );
  XOR2_X1 U10442 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n9416) );
  XNOR2_X1 U10443 ( .A(SI_30_), .B(keyinput_2), .ZN(n9415) );
  XNOR2_X1 U10444 ( .A(n9413), .B(keyinput_3), .ZN(n9414) );
  AOI211_X1 U10445 ( .C1(n9417), .C2(n9416), .A(n9415), .B(n9414), .ZN(n9423)
         );
  XNOR2_X1 U10446 ( .A(n9418), .B(keyinput_5), .ZN(n9422) );
  XNOR2_X1 U10447 ( .A(n9419), .B(keyinput_4), .ZN(n9421) );
  XNOR2_X1 U10448 ( .A(SI_26_), .B(keyinput_6), .ZN(n9420) );
  NOR4_X1 U10449 ( .A1(n9423), .A2(n9422), .A3(n9421), .A4(n9420), .ZN(n9430)
         );
  XNOR2_X1 U10450 ( .A(SI_25_), .B(keyinput_7), .ZN(n9429) );
  XNOR2_X1 U10451 ( .A(n9622), .B(keyinput_8), .ZN(n9427) );
  XNOR2_X1 U10452 ( .A(n9424), .B(keyinput_9), .ZN(n9426) );
  XNOR2_X1 U10453 ( .A(SI_22_), .B(keyinput_10), .ZN(n9425) );
  NOR3_X1 U10454 ( .A1(n9427), .A2(n9426), .A3(n9425), .ZN(n9428) );
  OAI21_X1 U10455 ( .B1(n9430), .B2(n9429), .A(n9428), .ZN(n9438) );
  XOR2_X1 U10456 ( .A(SI_18_), .B(keyinput_14), .Z(n9435) );
  XNOR2_X1 U10457 ( .A(n9431), .B(keyinput_12), .ZN(n9434) );
  XNOR2_X1 U10458 ( .A(SI_21_), .B(keyinput_11), .ZN(n9433) );
  XNOR2_X1 U10459 ( .A(SI_19_), .B(keyinput_13), .ZN(n9432) );
  NOR4_X1 U10460 ( .A1(n9435), .A2(n9434), .A3(n9433), .A4(n9432), .ZN(n9437)
         );
  XNOR2_X1 U10461 ( .A(n9636), .B(keyinput_15), .ZN(n9436) );
  AOI21_X1 U10462 ( .B1(n9438), .B2(n9437), .A(n9436), .ZN(n9443) );
  XNOR2_X1 U10463 ( .A(n9439), .B(keyinput_16), .ZN(n9442) );
  XNOR2_X1 U10464 ( .A(SI_14_), .B(keyinput_18), .ZN(n9441) );
  XNOR2_X1 U10465 ( .A(SI_15_), .B(keyinput_17), .ZN(n9440) );
  OAI211_X1 U10466 ( .C1(n9443), .C2(n9442), .A(n9441), .B(n9440), .ZN(n9451)
         );
  XNOR2_X1 U10467 ( .A(SI_10_), .B(keyinput_22), .ZN(n9447) );
  XNOR2_X1 U10468 ( .A(SI_11_), .B(keyinput_21), .ZN(n9446) );
  XNOR2_X1 U10469 ( .A(SI_13_), .B(keyinput_19), .ZN(n9445) );
  XNOR2_X1 U10470 ( .A(SI_12_), .B(keyinput_20), .ZN(n9444) );
  NOR4_X1 U10471 ( .A1(n9447), .A2(n9446), .A3(n9445), .A4(n9444), .ZN(n9450)
         );
  XNOR2_X1 U10472 ( .A(n9448), .B(keyinput_23), .ZN(n9449) );
  AOI21_X1 U10473 ( .B1(n9451), .B2(n9450), .A(n9449), .ZN(n9454) );
  XNOR2_X1 U10474 ( .A(SI_8_), .B(keyinput_24), .ZN(n9453) );
  XOR2_X1 U10475 ( .A(SI_7_), .B(keyinput_25), .Z(n9452) );
  OAI21_X1 U10476 ( .B1(n9454), .B2(n9453), .A(n9452), .ZN(n9458) );
  XNOR2_X1 U10477 ( .A(n9655), .B(keyinput_26), .ZN(n9457) );
  XNOR2_X1 U10478 ( .A(SI_5_), .B(keyinput_27), .ZN(n9456) );
  XNOR2_X1 U10479 ( .A(SI_4_), .B(keyinput_28), .ZN(n9455) );
  NAND4_X1 U10480 ( .A1(n9458), .A2(n9457), .A3(n9456), .A4(n9455), .ZN(n9461)
         );
  XNOR2_X1 U10481 ( .A(SI_3_), .B(keyinput_29), .ZN(n9460) );
  XNOR2_X1 U10482 ( .A(SI_2_), .B(keyinput_30), .ZN(n9459) );
  NAND3_X1 U10483 ( .A1(n9461), .A2(n9460), .A3(n9459), .ZN(n9468) );
  XNOR2_X1 U10484 ( .A(n9462), .B(keyinput_31), .ZN(n9467) );
  XNOR2_X1 U10485 ( .A(P2_U3152), .B(keyinput_34), .ZN(n9465) );
  XNOR2_X1 U10486 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n9464) );
  XNOR2_X1 U10487 ( .A(SI_0_), .B(keyinput_32), .ZN(n9463) );
  NAND3_X1 U10488 ( .A1(n9465), .A2(n9464), .A3(n9463), .ZN(n9466) );
  AOI21_X1 U10489 ( .B1(n9468), .B2(n9467), .A(n9466), .ZN(n9471) );
  XNOR2_X1 U10490 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n9470) );
  XOR2_X1 U10491 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .Z(n9469) );
  OAI21_X1 U10492 ( .B1(n9471), .B2(n9470), .A(n9469), .ZN(n9477) );
  XNOR2_X1 U10493 ( .A(n9472), .B(keyinput_37), .ZN(n9476) );
  XNOR2_X1 U10494 ( .A(n9473), .B(keyinput_38), .ZN(n9475) );
  XNOR2_X1 U10495 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n9474)
         );
  NAND4_X1 U10496 ( .A1(n9477), .A2(n9476), .A3(n9475), .A4(n9474), .ZN(n9480)
         );
  XNOR2_X1 U10497 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n9479) );
  XNOR2_X1 U10498 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_41), .ZN(n9478)
         );
  NAND3_X1 U10499 ( .A1(n9480), .A2(n9479), .A3(n9478), .ZN(n9493) );
  XNOR2_X1 U10500 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n9492)
         );
  XOR2_X1 U10501 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n9490) );
  XNOR2_X1 U10502 ( .A(n9481), .B(keyinput_43), .ZN(n9489) );
  XNOR2_X1 U10503 ( .A(n9482), .B(keyinput_46), .ZN(n9487) );
  XNOR2_X1 U10504 ( .A(n9483), .B(keyinput_48), .ZN(n9486) );
  XNOR2_X1 U10505 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n9485)
         );
  XNOR2_X1 U10506 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n9484)
         );
  NOR4_X1 U10507 ( .A1(n9487), .A2(n9486), .A3(n9485), .A4(n9484), .ZN(n9488)
         );
  NAND3_X1 U10508 ( .A1(n9490), .A2(n9489), .A3(n9488), .ZN(n9491) );
  AOI21_X1 U10509 ( .B1(n9493), .B2(n9492), .A(n9491), .ZN(n9497) );
  XNOR2_X1 U10510 ( .A(n9692), .B(keyinput_51), .ZN(n9496) );
  XNOR2_X1 U10511 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n9495)
         );
  XNOR2_X1 U10512 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n9494) );
  NOR4_X1 U10513 ( .A1(n9497), .A2(n9496), .A3(n9495), .A4(n9494), .ZN(n9501)
         );
  XOR2_X1 U10514 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .Z(n9500) );
  XOR2_X1 U10515 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n9499) );
  XNOR2_X1 U10516 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n9498) );
  OAI211_X1 U10517 ( .C1(n9501), .C2(n9500), .A(n9499), .B(n9498), .ZN(n9504)
         );
  XNOR2_X1 U10518 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n9503)
         );
  XNOR2_X1 U10519 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .ZN(n9502)
         );
  AOI21_X1 U10520 ( .B1(n9504), .B2(n9503), .A(n9502), .ZN(n9507) );
  XNOR2_X1 U10521 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n9506)
         );
  XNOR2_X1 U10522 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n9505)
         );
  OAI21_X1 U10523 ( .B1(n9507), .B2(n9506), .A(n9505), .ZN(n9510) );
  XNOR2_X1 U10524 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .ZN(n9509)
         );
  XNOR2_X1 U10525 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n9508) );
  NAND3_X1 U10526 ( .A1(n9510), .A2(n9509), .A3(n9508), .ZN(n9513) );
  XNOR2_X1 U10527 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n9512) );
  XNOR2_X1 U10528 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n9511)
         );
  NAND3_X1 U10529 ( .A1(n9513), .A2(n9512), .A3(n9511), .ZN(n9524) );
  XNOR2_X1 U10530 ( .A(n9514), .B(keyinput_63), .ZN(n9523) );
  XOR2_X1 U10531 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n9518) );
  XNOR2_X1 U10532 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n9517)
         );
  XOR2_X1 U10533 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .Z(n9516) );
  XOR2_X1 U10534 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n9515) );
  NOR4_X1 U10535 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n9515), .ZN(n9521)
         );
  XOR2_X1 U10536 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .Z(n9520) );
  XOR2_X1 U10537 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n9519) );
  NAND3_X1 U10538 ( .A1(n9521), .A2(n9520), .A3(n9519), .ZN(n9522) );
  AOI21_X1 U10539 ( .B1(n9524), .B2(n9523), .A(n9522), .ZN(n9529) );
  XNOR2_X1 U10540 ( .A(n9525), .B(keyinput_70), .ZN(n9528) );
  XNOR2_X1 U10541 ( .A(n9526), .B(keyinput_71), .ZN(n9527) );
  OAI21_X1 U10542 ( .B1(n9529), .B2(n9528), .A(n9527), .ZN(n9534) );
  XOR2_X1 U10543 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n9533) );
  XNOR2_X1 U10544 ( .A(n9530), .B(keyinput_74), .ZN(n9532) );
  XNOR2_X1 U10545 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n9531)
         );
  NAND4_X1 U10546 ( .A1(n9534), .A2(n9533), .A3(n9532), .A4(n9531), .ZN(n9545)
         );
  XNOR2_X1 U10547 ( .A(n9737), .B(keyinput_76), .ZN(n9538) );
  XNOR2_X1 U10548 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n9537)
         );
  XNOR2_X1 U10549 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n9536)
         );
  XNOR2_X1 U10550 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .ZN(n9535)
         );
  NOR4_X1 U10551 ( .A1(n9538), .A2(n9537), .A3(n9536), .A4(n9535), .ZN(n9544)
         );
  XOR2_X1 U10552 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .Z(n9542) );
  XOR2_X1 U10553 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n9541) );
  XNOR2_X1 U10554 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n9540)
         );
  XNOR2_X1 U10555 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n9539)
         );
  NAND4_X1 U10556 ( .A1(n9542), .A2(n9541), .A3(n9540), .A4(n9539), .ZN(n9543)
         );
  AOI21_X1 U10557 ( .B1(n9545), .B2(n9544), .A(n9543), .ZN(n9553) );
  XNOR2_X1 U10558 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n9552)
         );
  XNOR2_X1 U10559 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n9551)
         );
  XNOR2_X1 U10560 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .ZN(n9549)
         );
  XNOR2_X1 U10561 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n9548)
         );
  XNOR2_X1 U10562 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n9547)
         );
  XNOR2_X1 U10563 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n9546)
         );
  NAND4_X1 U10564 ( .A1(n9549), .A2(n9548), .A3(n9547), .A4(n9546), .ZN(n9550)
         );
  NOR4_X1 U10565 ( .A1(n9553), .A2(n9552), .A3(n9551), .A4(n9550), .ZN(n9565)
         );
  XOR2_X1 U10566 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .Z(n9557) );
  XOR2_X1 U10567 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .Z(n9556) );
  XNOR2_X1 U10568 ( .A(n10633), .B(keyinput_91), .ZN(n9555) );
  XNOR2_X1 U10569 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_92), .ZN(n9554) );
  NAND4_X1 U10570 ( .A1(n9557), .A2(n9556), .A3(n9555), .A4(n9554), .ZN(n9564)
         );
  XNOR2_X1 U10571 ( .A(n9558), .B(keyinput_94), .ZN(n9562) );
  XNOR2_X1 U10572 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .ZN(n9561) );
  XNOR2_X1 U10573 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_93), .ZN(n9560) );
  XNOR2_X1 U10574 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_95), .ZN(n9559) );
  NOR4_X1 U10575 ( .A1(n9562), .A2(n9561), .A3(n9560), .A4(n9559), .ZN(n9563)
         );
  OAI21_X1 U10576 ( .B1(n9565), .B2(n9564), .A(n9563), .ZN(n9569) );
  XNOR2_X1 U10577 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_97), .ZN(n9568) );
  XNOR2_X1 U10578 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_98), .ZN(n9567) );
  XNOR2_X1 U10579 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_99), .ZN(n9566) );
  AOI211_X1 U10580 ( .C1(n9569), .C2(n9568), .A(n9567), .B(n9566), .ZN(n9577)
         );
  XNOR2_X1 U10581 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_100), .ZN(n9576) );
  XOR2_X1 U10582 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_103), .Z(n9574) );
  XNOR2_X1 U10583 ( .A(n9570), .B(keyinput_101), .ZN(n9573) );
  XNOR2_X1 U10584 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_102), .ZN(n9572) );
  XNOR2_X1 U10585 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_104), .ZN(n9571) );
  NOR4_X1 U10586 ( .A1(n9574), .A2(n9573), .A3(n9572), .A4(n9571), .ZN(n9575)
         );
  OAI21_X1 U10587 ( .B1(n9577), .B2(n9576), .A(n9575), .ZN(n9582) );
  XNOR2_X1 U10588 ( .A(n9578), .B(keyinput_105), .ZN(n9581) );
  XNOR2_X1 U10589 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_106), .ZN(n9580) );
  XNOR2_X1 U10590 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_107), .ZN(n9579) );
  NAND4_X1 U10591 ( .A1(n9582), .A2(n9581), .A3(n9580), .A4(n9579), .ZN(n9586)
         );
  XNOR2_X1 U10592 ( .A(n9583), .B(keyinput_108), .ZN(n9585) );
  XNOR2_X1 U10593 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_109), .ZN(n9584) );
  AOI21_X1 U10594 ( .B1(n9586), .B2(n9585), .A(n9584), .ZN(n9590) );
  XNOR2_X1 U10595 ( .A(n9587), .B(keyinput_110), .ZN(n9589) );
  XNOR2_X1 U10596 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_111), .ZN(n9588) );
  OAI21_X1 U10597 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9598) );
  XNOR2_X1 U10598 ( .A(n9796), .B(keyinput_112), .ZN(n9597) );
  XNOR2_X1 U10599 ( .A(n9797), .B(keyinput_113), .ZN(n9595) );
  XNOR2_X1 U10600 ( .A(n9799), .B(keyinput_115), .ZN(n9594) );
  XNOR2_X1 U10601 ( .A(n9591), .B(keyinput_114), .ZN(n9593) );
  XNOR2_X1 U10602 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_116), .ZN(n9592) );
  NAND4_X1 U10603 ( .A1(n9595), .A2(n9594), .A3(n9593), .A4(n9592), .ZN(n9596)
         );
  AOI21_X1 U10604 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n9601) );
  XNOR2_X1 U10605 ( .A(n9807), .B(keyinput_117), .ZN(n9600) );
  XNOR2_X1 U10606 ( .A(n9808), .B(keyinput_118), .ZN(n9599) );
  NOR3_X1 U10607 ( .A1(n9601), .A2(n9600), .A3(n9599), .ZN(n9604) );
  XNOR2_X1 U10608 ( .A(n9812), .B(keyinput_119), .ZN(n9603) );
  XNOR2_X1 U10609 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_120), .ZN(n9602) );
  OAI21_X1 U10610 ( .B1(n9604), .B2(n9603), .A(n9602), .ZN(n9609) );
  XNOR2_X1 U10611 ( .A(n9605), .B(keyinput_121), .ZN(n9608) );
  XNOR2_X1 U10612 ( .A(n9817), .B(keyinput_123), .ZN(n9607) );
  XOR2_X1 U10613 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .Z(n9606) );
  NAND4_X1 U10614 ( .A1(n9609), .A2(n9608), .A3(n9607), .A4(n9606), .ZN(n9612)
         );
  XNOR2_X1 U10615 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_124), .ZN(n9611) );
  INV_X1 U10616 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10542) );
  XNOR2_X1 U10617 ( .A(n10542), .B(keyinput_125), .ZN(n9610) );
  AOI21_X1 U10618 ( .B1(n9612), .B2(n9611), .A(n9610), .ZN(n9831) );
  INV_X1 U10619 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10543) );
  XNOR2_X1 U10620 ( .A(n10543), .B(keyinput_126), .ZN(n9830) );
  XNOR2_X1 U10621 ( .A(SI_31_), .B(keyinput_129), .ZN(n9616) );
  XNOR2_X1 U10622 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .ZN(n9615) );
  XOR2_X1 U10623 ( .A(SI_30_), .B(keyinput_130), .Z(n9614) );
  XNOR2_X1 U10624 ( .A(SI_29_), .B(keyinput_131), .ZN(n9613) );
  OAI211_X1 U10625 ( .C1(n9616), .C2(n9615), .A(n9614), .B(n9613), .ZN(n9620)
         );
  XNOR2_X1 U10626 ( .A(SI_26_), .B(keyinput_134), .ZN(n9619) );
  XNOR2_X1 U10627 ( .A(SI_28_), .B(keyinput_132), .ZN(n9618) );
  XNOR2_X1 U10628 ( .A(SI_27_), .B(keyinput_133), .ZN(n9617) );
  NAND4_X1 U10629 ( .A1(n9620), .A2(n9619), .A3(n9618), .A4(n9617), .ZN(n9629)
         );
  XNOR2_X1 U10630 ( .A(n9621), .B(keyinput_135), .ZN(n9628) );
  XNOR2_X1 U10631 ( .A(n9622), .B(keyinput_136), .ZN(n9626) );
  XNOR2_X1 U10632 ( .A(n9623), .B(keyinput_138), .ZN(n9625) );
  XNOR2_X1 U10633 ( .A(SI_23_), .B(keyinput_137), .ZN(n9624) );
  NAND3_X1 U10634 ( .A1(n9626), .A2(n9625), .A3(n9624), .ZN(n9627) );
  AOI21_X1 U10635 ( .B1(n9629), .B2(n9628), .A(n9627), .ZN(n9639) );
  XNOR2_X1 U10636 ( .A(n9630), .B(keyinput_139), .ZN(n9635) );
  XNOR2_X1 U10637 ( .A(n9631), .B(keyinput_141), .ZN(n9634) );
  XNOR2_X1 U10638 ( .A(SI_18_), .B(keyinput_142), .ZN(n9633) );
  XNOR2_X1 U10639 ( .A(SI_20_), .B(keyinput_140), .ZN(n9632) );
  NAND4_X1 U10640 ( .A1(n9635), .A2(n9634), .A3(n9633), .A4(n9632), .ZN(n9638)
         );
  XNOR2_X1 U10641 ( .A(n9636), .B(keyinput_143), .ZN(n9637) );
  OAI21_X1 U10642 ( .B1(n9639), .B2(n9638), .A(n9637), .ZN(n9643) );
  XNOR2_X1 U10643 ( .A(SI_16_), .B(keyinput_144), .ZN(n9642) );
  XOR2_X1 U10644 ( .A(SI_15_), .B(keyinput_145), .Z(n9641) );
  XNOR2_X1 U10645 ( .A(SI_14_), .B(keyinput_146), .ZN(n9640) );
  AOI211_X1 U10646 ( .C1(n9643), .C2(n9642), .A(n9641), .B(n9640), .ZN(n9651)
         );
  XNOR2_X1 U10647 ( .A(n9644), .B(keyinput_150), .ZN(n9648) );
  XNOR2_X1 U10648 ( .A(SI_12_), .B(keyinput_148), .ZN(n9647) );
  XNOR2_X1 U10649 ( .A(SI_13_), .B(keyinput_147), .ZN(n9646) );
  XNOR2_X1 U10650 ( .A(SI_11_), .B(keyinput_149), .ZN(n9645) );
  NAND4_X1 U10651 ( .A1(n9648), .A2(n9647), .A3(n9646), .A4(n9645), .ZN(n9650)
         );
  XNOR2_X1 U10652 ( .A(SI_9_), .B(keyinput_151), .ZN(n9649) );
  OAI21_X1 U10653 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9654) );
  XNOR2_X1 U10654 ( .A(SI_8_), .B(keyinput_152), .ZN(n9653) );
  XOR2_X1 U10655 ( .A(SI_7_), .B(keyinput_153), .Z(n9652) );
  AOI21_X1 U10656 ( .B1(n9654), .B2(n9653), .A(n9652), .ZN(n9659) );
  XNOR2_X1 U10657 ( .A(n9655), .B(keyinput_154), .ZN(n9658) );
  XNOR2_X1 U10658 ( .A(SI_5_), .B(keyinput_155), .ZN(n9657) );
  XNOR2_X1 U10659 ( .A(SI_4_), .B(keyinput_156), .ZN(n9656) );
  NOR4_X1 U10660 ( .A1(n9659), .A2(n9658), .A3(n9657), .A4(n9656), .ZN(n9662)
         );
  XNOR2_X1 U10661 ( .A(SI_3_), .B(keyinput_157), .ZN(n9661) );
  XNOR2_X1 U10662 ( .A(SI_2_), .B(keyinput_158), .ZN(n9660) );
  NOR3_X1 U10663 ( .A1(n9662), .A2(n9661), .A3(n9660), .ZN(n9668) );
  XNOR2_X1 U10664 ( .A(SI_1_), .B(keyinput_159), .ZN(n9667) );
  XNOR2_X1 U10665 ( .A(n10687), .B(keyinput_161), .ZN(n9665) );
  XNOR2_X1 U10666 ( .A(P2_U3152), .B(keyinput_162), .ZN(n9664) );
  XNOR2_X1 U10667 ( .A(SI_0_), .B(keyinput_160), .ZN(n9663) );
  NOR3_X1 U10668 ( .A1(n9665), .A2(n9664), .A3(n9663), .ZN(n9666) );
  OAI21_X1 U10669 ( .B1(n9668), .B2(n9667), .A(n9666), .ZN(n9671) );
  XNOR2_X1 U10670 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n9670)
         );
  XOR2_X1 U10671 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .Z(n9669) );
  AOI21_X1 U10672 ( .B1(n9671), .B2(n9670), .A(n9669), .ZN(n9676) );
  XNOR2_X1 U10673 ( .A(n9672), .B(keyinput_167), .ZN(n9675) );
  XNOR2_X1 U10674 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n9674)
         );
  XNOR2_X1 U10675 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n9673)
         );
  NOR4_X1 U10676 ( .A1(n9676), .A2(n9675), .A3(n9674), .A4(n9673), .ZN(n9679)
         );
  XNOR2_X1 U10677 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n9678)
         );
  XNOR2_X1 U10678 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n9677)
         );
  NOR3_X1 U10679 ( .A1(n9679), .A2(n9678), .A3(n9677), .ZN(n9691) );
  XNOR2_X1 U10680 ( .A(n9680), .B(keyinput_170), .ZN(n9690) );
  XNOR2_X1 U10681 ( .A(n9681), .B(keyinput_173), .ZN(n9685) );
  XNOR2_X1 U10682 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n9684)
         );
  XNOR2_X1 U10683 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n9683)
         );
  XNOR2_X1 U10684 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_174), .ZN(n9682)
         );
  NAND4_X1 U10685 ( .A1(n9685), .A2(n9684), .A3(n9683), .A4(n9682), .ZN(n9688)
         );
  XNOR2_X1 U10686 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n9687)
         );
  XNOR2_X1 U10687 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n9686)
         );
  NOR3_X1 U10688 ( .A1(n9688), .A2(n9687), .A3(n9686), .ZN(n9689) );
  OAI21_X1 U10689 ( .B1(n9691), .B2(n9690), .A(n9689), .ZN(n9698) );
  XNOR2_X1 U10690 ( .A(n9692), .B(keyinput_179), .ZN(n9697) );
  OAI22_X1 U10691 ( .A1(n9694), .A2(keyinput_177), .B1(keyinput_178), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n9693) );
  AOI21_X1 U10692 ( .B1(n9694), .B2(keyinput_177), .A(n9693), .ZN(n9696) );
  NAND2_X1 U10693 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_178), .ZN(n9695) );
  NAND4_X1 U10694 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(n9702)
         );
  XOR2_X1 U10695 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .Z(n9701) );
  XNOR2_X1 U10696 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_181), .ZN(n9700)
         );
  XNOR2_X1 U10697 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n9699)
         );
  AOI211_X1 U10698 ( .C1(n9702), .C2(n9701), .A(n9700), .B(n9699), .ZN(n9707)
         );
  XNOR2_X1 U10699 ( .A(n9703), .B(keyinput_183), .ZN(n9706) );
  XNOR2_X1 U10700 ( .A(n9704), .B(keyinput_184), .ZN(n9705) );
  OAI21_X1 U10701 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9710) );
  XNOR2_X1 U10702 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_185), .ZN(n9709)
         );
  XNOR2_X1 U10703 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n9708)
         );
  AOI21_X1 U10704 ( .B1(n9710), .B2(n9709), .A(n9708), .ZN(n9717) );
  XOR2_X1 U10705 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .Z(n9712) );
  XNOR2_X1 U10706 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n9711)
         );
  NAND2_X1 U10707 ( .A1(n9712), .A2(n9711), .ZN(n9716) );
  XNOR2_X1 U10708 ( .A(n9713), .B(keyinput_190), .ZN(n9715) );
  XNOR2_X1 U10709 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n9714)
         );
  OAI211_X1 U10710 ( .C1(n9717), .C2(n9716), .A(n9715), .B(n9714), .ZN(n9727)
         );
  XNOR2_X1 U10711 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_191), .ZN(n9726)
         );
  XOR2_X1 U10712 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .Z(n9721) );
  XOR2_X1 U10713 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .Z(n9720)
         );
  XOR2_X1 U10714 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .Z(n9719)
         );
  XOR2_X1 U10715 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .Z(n9718)
         );
  NOR4_X1 U10716 ( .A1(n9721), .A2(n9720), .A3(n9719), .A4(n9718), .ZN(n9724)
         );
  XOR2_X1 U10717 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .Z(n9723)
         );
  XOR2_X1 U10718 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .Z(n9722)
         );
  NAND3_X1 U10719 ( .A1(n9724), .A2(n9723), .A3(n9722), .ZN(n9725) );
  AOI21_X1 U10720 ( .B1(n9727), .B2(n9726), .A(n9725), .ZN(n9730) );
  XNOR2_X1 U10721 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .ZN(n9729)
         );
  XNOR2_X1 U10722 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_199), .ZN(n9728)
         );
  OAI21_X1 U10723 ( .B1(n9730), .B2(n9729), .A(n9728), .ZN(n9735) );
  XNOR2_X1 U10724 ( .A(n9731), .B(keyinput_201), .ZN(n9734) );
  XNOR2_X1 U10725 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n9733)
         );
  XNOR2_X1 U10726 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n9732)
         );
  NAND4_X1 U10727 ( .A1(n9735), .A2(n9734), .A3(n9733), .A4(n9732), .ZN(n9749)
         );
  XOR2_X1 U10728 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n9741)
         );
  XNOR2_X1 U10729 ( .A(n9736), .B(keyinput_205), .ZN(n9740) );
  XNOR2_X1 U10730 ( .A(n9737), .B(keyinput_204), .ZN(n9739) );
  XNOR2_X1 U10731 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .ZN(n9738)
         );
  NOR4_X1 U10732 ( .A1(n9741), .A2(n9740), .A3(n9739), .A4(n9738), .ZN(n9748)
         );
  XOR2_X1 U10733 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_210), .Z(n9746)
         );
  XNOR2_X1 U10734 ( .A(n9742), .B(keyinput_208), .ZN(n9745) );
  XNOR2_X1 U10735 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n9744)
         );
  XNOR2_X1 U10736 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n9743)
         );
  NAND4_X1 U10737 ( .A1(n9746), .A2(n9745), .A3(n9744), .A4(n9743), .ZN(n9747)
         );
  AOI21_X1 U10738 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(n9758) );
  XNOR2_X1 U10739 ( .A(n9750), .B(keyinput_215), .ZN(n9757) );
  XNOR2_X1 U10740 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .ZN(n9756)
         );
  XNOR2_X1 U10741 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .ZN(n9754)
         );
  XNOR2_X1 U10742 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n9753)
         );
  XNOR2_X1 U10743 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n9752)
         );
  XNOR2_X1 U10744 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .ZN(n9751)
         );
  NAND4_X1 U10745 ( .A1(n9754), .A2(n9753), .A3(n9752), .A4(n9751), .ZN(n9755)
         );
  NOR4_X1 U10746 ( .A1(n9758), .A2(n9757), .A3(n9756), .A4(n9755), .ZN(n9771)
         );
  XNOR2_X1 U10747 ( .A(n9759), .B(keyinput_220), .ZN(n9763) );
  XNOR2_X1 U10748 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_218), .ZN(n9762)
         );
  XNOR2_X1 U10749 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_219), .ZN(n9761) );
  XNOR2_X1 U10750 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .ZN(n9760)
         );
  NAND4_X1 U10751 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n9770)
         );
  XNOR2_X1 U10752 ( .A(n9764), .B(keyinput_223), .ZN(n9768) );
  XNOR2_X1 U10753 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_222), .ZN(n9767) );
  XNOR2_X1 U10754 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_224), .ZN(n9766) );
  XNOR2_X1 U10755 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_221), .ZN(n9765) );
  NOR4_X1 U10756 ( .A1(n9768), .A2(n9767), .A3(n9766), .A4(n9765), .ZN(n9769)
         );
  OAI21_X1 U10757 ( .B1(n9771), .B2(n9770), .A(n9769), .ZN(n9776) );
  XNOR2_X1 U10758 ( .A(n9772), .B(keyinput_225), .ZN(n9775) );
  XNOR2_X1 U10759 ( .A(n5864), .B(keyinput_227), .ZN(n9774) );
  XNOR2_X1 U10760 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_226), .ZN(n9773) );
  AOI211_X1 U10761 ( .C1(n9776), .C2(n9775), .A(n9774), .B(n9773), .ZN(n9784)
         );
  XNOR2_X1 U10762 ( .A(n9777), .B(keyinput_228), .ZN(n9783) );
  XOR2_X1 U10763 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_232), .Z(n9781) );
  XOR2_X1 U10764 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_231), .Z(n9780) );
  XNOR2_X1 U10765 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_229), .ZN(n9779) );
  XNOR2_X1 U10766 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_230), .ZN(n9778) );
  NOR4_X1 U10767 ( .A1(n9781), .A2(n9780), .A3(n9779), .A4(n9778), .ZN(n9782)
         );
  OAI21_X1 U10768 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9789) );
  XNOR2_X1 U10769 ( .A(n9785), .B(keyinput_234), .ZN(n9788) );
  XNOR2_X1 U10770 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_235), .ZN(n9787) );
  XNOR2_X1 U10771 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_233), .ZN(n9786) );
  NAND4_X1 U10772 ( .A1(n9789), .A2(n9788), .A3(n9787), .A4(n9786), .ZN(n9792)
         );
  XNOR2_X1 U10773 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_236), .ZN(n9791) );
  XNOR2_X1 U10774 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_237), .ZN(n9790) );
  AOI21_X1 U10775 ( .B1(n9792), .B2(n9791), .A(n9790), .ZN(n9795) );
  XNOR2_X1 U10776 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_238), .ZN(n9794) );
  XNOR2_X1 U10777 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_239), .ZN(n9793) );
  OAI21_X1 U10778 ( .B1(n9795), .B2(n9794), .A(n9793), .ZN(n9806) );
  XNOR2_X1 U10779 ( .A(n9796), .B(keyinput_240), .ZN(n9805) );
  XNOR2_X1 U10780 ( .A(n9797), .B(keyinput_241), .ZN(n9803) );
  XNOR2_X1 U10781 ( .A(n9798), .B(keyinput_244), .ZN(n9802) );
  XNOR2_X1 U10782 ( .A(n9799), .B(keyinput_243), .ZN(n9801) );
  XNOR2_X1 U10783 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_242), .ZN(n9800) );
  NAND4_X1 U10784 ( .A1(n9803), .A2(n9802), .A3(n9801), .A4(n9800), .ZN(n9804)
         );
  AOI21_X1 U10785 ( .B1(n9806), .B2(n9805), .A(n9804), .ZN(n9811) );
  XNOR2_X1 U10786 ( .A(n9807), .B(keyinput_245), .ZN(n9810) );
  XNOR2_X1 U10787 ( .A(n9808), .B(keyinput_246), .ZN(n9809) );
  NOR3_X1 U10788 ( .A1(n9811), .A2(n9810), .A3(n9809), .ZN(n9816) );
  XNOR2_X1 U10789 ( .A(n9812), .B(keyinput_247), .ZN(n9815) );
  XNOR2_X1 U10790 ( .A(n9813), .B(keyinput_248), .ZN(n9814) );
  OAI21_X1 U10791 ( .B1(n9816), .B2(n9815), .A(n9814), .ZN(n9821) );
  XOR2_X1 U10792 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_250), .Z(n9820) );
  XNOR2_X1 U10793 ( .A(n9817), .B(keyinput_251), .ZN(n9819) );
  XNOR2_X1 U10794 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_249), .ZN(n9818) );
  NAND4_X1 U10795 ( .A1(n9821), .A2(n9820), .A3(n9819), .A4(n9818), .ZN(n9824)
         );
  XOR2_X1 U10796 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_252), .Z(n9823) );
  XNOR2_X1 U10797 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_253), .ZN(n9822) );
  AOI21_X1 U10798 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9827) );
  XNOR2_X1 U10799 ( .A(n10543), .B(keyinput_254), .ZN(n9826) );
  XOR2_X1 U10800 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_255), .Z(n9825) );
  OAI21_X1 U10801 ( .B1(n9827), .B2(n9826), .A(n9825), .ZN(n9829) );
  XOR2_X1 U10802 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_127), .Z(n9828) );
  OAI211_X1 U10803 ( .C1(n9831), .C2(n9830), .A(n9829), .B(n9828), .ZN(n9832)
         );
  XNOR2_X1 U10804 ( .A(n9833), .B(n9832), .ZN(P2_U3276) );
  OAI21_X1 U10805 ( .B1(n9836), .B2(n9835), .A(n9834), .ZN(n9969) );
  AOI22_X1 U10806 ( .A1(n9967), .A2(n9901), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n10906), .ZN(n9852) );
  NAND2_X1 U10807 ( .A1(n9838), .A2(n9837), .ZN(n9840) );
  XNOR2_X1 U10808 ( .A(n9840), .B(n9839), .ZN(n9841) );
  OAI222_X1 U10809 ( .A1(n10939), .A2(n9842), .B1(n10937), .B2(n9876), .C1(
        n10811), .C2(n9841), .ZN(n9965) );
  OR2_X1 U10810 ( .A1(n9855), .A2(n9843), .ZN(n9844) );
  AND3_X1 U10811 ( .A1(n9845), .A2(n9844), .A3(n10892), .ZN(n9966) );
  NAND2_X1 U10812 ( .A1(n9966), .A2(n9846), .ZN(n9847) );
  OAI21_X1 U10813 ( .B1(n9849), .B2(n9848), .A(n9847), .ZN(n9850) );
  OAI21_X1 U10814 ( .B1(n9965), .B2(n9850), .A(n10957), .ZN(n9851) );
  OAI211_X1 U10815 ( .C1(n9969), .C2(n9887), .A(n9852), .B(n9851), .ZN(
        P2_U3277) );
  XNOR2_X1 U10816 ( .A(n9854), .B(n9853), .ZN(n9974) );
  INV_X1 U10817 ( .A(n9878), .ZN(n9856) );
  AOI21_X1 U10818 ( .B1(n9970), .B2(n9856), .A(n9855), .ZN(n9971) );
  AOI22_X1 U10819 ( .A1(n10906), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9857), 
        .B2(n10962), .ZN(n9858) );
  OAI21_X1 U10820 ( .B1(n9859), .B2(n10956), .A(n9858), .ZN(n9866) );
  XNOR2_X1 U10821 ( .A(n9861), .B(n9860), .ZN(n9864) );
  AOI222_X1 U10822 ( .A1(n10942), .A2(n9864), .B1(n9863), .B2(n9890), .C1(
        n9862), .C2(n9892), .ZN(n9973) );
  NOR2_X1 U10823 ( .A1(n9973), .A2(n10906), .ZN(n9865) );
  AOI211_X1 U10824 ( .C1(n9971), .C2(n9897), .A(n9866), .B(n9865), .ZN(n9867)
         );
  OAI21_X1 U10825 ( .B1(n9974), .B2(n9887), .A(n9867), .ZN(P2_U3278) );
  OAI21_X1 U10826 ( .B1(n9870), .B2(n9869), .A(n9868), .ZN(n9871) );
  INV_X1 U10827 ( .A(n9871), .ZN(n9979) );
  XNOR2_X1 U10828 ( .A(n9872), .B(n9873), .ZN(n9875) );
  OAI222_X1 U10829 ( .A1(n10939), .A2(n9876), .B1(n9875), .B2(n10811), .C1(
        n10937), .C2(n9874), .ZN(n9975) );
  INV_X1 U10830 ( .A(n9877), .ZN(n9879) );
  AOI211_X1 U10831 ( .C1(n9977), .C2(n9879), .A(n11070), .B(n9878), .ZN(n9976)
         );
  NAND2_X1 U10832 ( .A1(n9976), .A2(n9880), .ZN(n9883) );
  AOI22_X1 U10833 ( .A1(n10906), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9881), 
        .B2(n10962), .ZN(n9882) );
  OAI211_X1 U10834 ( .C1(n9884), .C2(n10956), .A(n9883), .B(n9882), .ZN(n9885)
         );
  AOI21_X1 U10835 ( .B1(n9975), .B2(n10957), .A(n9885), .ZN(n9886) );
  OAI21_X1 U10836 ( .B1(n9979), .B2(n9887), .A(n9886), .ZN(P2_U3279) );
  XNOR2_X1 U10837 ( .A(n9888), .B(n9900), .ZN(n9889) );
  AOI222_X1 U10838 ( .A1(n9893), .A2(n9892), .B1(n9891), .B2(n9890), .C1(
        n10942), .C2(n9889), .ZN(n10837) );
  MUX2_X1 U10839 ( .A(n7298), .B(n10837), .S(n10957), .Z(n9905) );
  INV_X1 U10840 ( .A(n9894), .ZN(n9895) );
  AOI21_X1 U10841 ( .B1(n10832), .B2(n10802), .A(n9895), .ZN(n10833) );
  AOI22_X1 U10842 ( .A1(n10833), .A2(n9897), .B1(n9896), .B2(n10962), .ZN(
        n9904) );
  NAND2_X1 U10843 ( .A1(n9899), .A2(n9900), .ZN(n10834) );
  NAND3_X1 U10844 ( .A1(n9898), .A2(n10834), .A3(n10790), .ZN(n9903) );
  NAND2_X1 U10845 ( .A1(n9901), .A2(n10832), .ZN(n9902) );
  NAND4_X1 U10846 ( .A1(n9905), .A2(n9904), .A3(n9903), .A4(n9902), .ZN(
        P2_U3290) );
  AOI21_X1 U10847 ( .B1(n9907), .B2(n10975), .A(n9906), .ZN(n9908) );
  OAI21_X1 U10848 ( .B1(n9909), .B2(n11070), .A(n9908), .ZN(n9985) );
  MUX2_X1 U10849 ( .A(n9985), .B(P2_REG1_REG_31__SCAN_IN), .S(n11076), .Z(
        P2_U3551) );
  NAND3_X1 U10850 ( .A1(n9911), .A2(n10892), .A3(n9910), .ZN(n9913) );
  OAI211_X1 U10851 ( .C1(n9914), .C2(n11069), .A(n9913), .B(n9912), .ZN(n9986)
         );
  MUX2_X1 U10852 ( .A(n9986), .B(P2_REG1_REG_30__SCAN_IN), .S(n11076), .Z(
        P2_U3550) );
  MUX2_X1 U10853 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9987), .S(n11078), .Z(
        P2_U3549) );
  AOI22_X1 U10854 ( .A1(n9920), .A2(n10892), .B1(n10975), .B2(n9919), .ZN(
        n9921) );
  OAI211_X1 U10855 ( .C1(n9923), .C2(n11034), .A(n9922), .B(n9921), .ZN(n9988)
         );
  MUX2_X1 U10856 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9988), .S(n11078), .Z(
        P2_U3548) );
  AOI22_X1 U10857 ( .A1(n9925), .A2(n10892), .B1(n10975), .B2(n9924), .ZN(
        n9926) );
  OAI211_X1 U10858 ( .C1(n9928), .C2(n11034), .A(n9927), .B(n9926), .ZN(n9989)
         );
  MUX2_X1 U10859 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9989), .S(n11078), .Z(
        P2_U3547) );
  AOI21_X1 U10860 ( .B1(n10975), .B2(n9930), .A(n9929), .ZN(n9931) );
  OAI211_X1 U10861 ( .C1(n9933), .C2(n11034), .A(n9932), .B(n9931), .ZN(n9990)
         );
  MUX2_X1 U10862 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9990), .S(n11078), .Z(
        P2_U3546) );
  AOI211_X1 U10863 ( .C1(n10975), .C2(n9936), .A(n9935), .B(n9934), .ZN(n9937)
         );
  OAI21_X1 U10864 ( .B1(n9938), .B2(n11034), .A(n9937), .ZN(n9991) );
  MUX2_X1 U10865 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9991), .S(n11078), .Z(
        P2_U3545) );
  AOI22_X1 U10866 ( .A1(n9940), .A2(n10892), .B1(n10975), .B2(n9939), .ZN(
        n9941) );
  OAI211_X1 U10867 ( .C1(n9943), .C2(n11034), .A(n9942), .B(n9941), .ZN(n9992)
         );
  MUX2_X1 U10868 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9992), .S(n11078), .Z(
        P2_U3544) );
  NAND2_X1 U10869 ( .A1(n9944), .A2(n11074), .ZN(n9949) );
  AOI22_X1 U10870 ( .A1(n9946), .A2(n10892), .B1(n10975), .B2(n9945), .ZN(
        n9947) );
  OAI211_X1 U10871 ( .C1(n9359), .C2(n9949), .A(n9948), .B(n9947), .ZN(n9993)
         );
  MUX2_X1 U10872 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9993), .S(n11078), .Z(
        P2_U3543) );
  AOI22_X1 U10873 ( .A1(n9951), .A2(n10892), .B1(n10975), .B2(n9950), .ZN(
        n9952) );
  OAI211_X1 U10874 ( .C1(n9954), .C2(n11034), .A(n9953), .B(n9952), .ZN(n9994)
         );
  MUX2_X1 U10875 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9994), .S(n11078), .Z(
        P2_U3542) );
  AOI22_X1 U10876 ( .A1(n9956), .A2(n10892), .B1(n10975), .B2(n9955), .ZN(
        n9957) );
  OAI211_X1 U10877 ( .C1(n9959), .C2(n11034), .A(n9958), .B(n9957), .ZN(n9995)
         );
  MUX2_X1 U10878 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9995), .S(n11078), .Z(
        P2_U3541) );
  AOI22_X1 U10879 ( .A1(n9961), .A2(n10892), .B1(n10975), .B2(n9960), .ZN(
        n9962) );
  OAI211_X1 U10880 ( .C1(n9964), .C2(n11034), .A(n9963), .B(n9962), .ZN(n9996)
         );
  MUX2_X1 U10881 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9996), .S(n11078), .Z(
        P2_U3540) );
  AOI211_X1 U10882 ( .C1(n10975), .C2(n9967), .A(n9966), .B(n9965), .ZN(n9968)
         );
  OAI21_X1 U10883 ( .B1(n9969), .B2(n11034), .A(n9968), .ZN(n9997) );
  MUX2_X1 U10884 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9997), .S(n11078), .Z(
        P2_U3539) );
  AOI22_X1 U10885 ( .A1(n9971), .A2(n10892), .B1(n10975), .B2(n9970), .ZN(
        n9972) );
  OAI211_X1 U10886 ( .C1(n9974), .C2(n11034), .A(n9973), .B(n9972), .ZN(n9998)
         );
  MUX2_X1 U10887 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9998), .S(n11078), .Z(
        P2_U3538) );
  AOI211_X1 U10888 ( .C1(n10975), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9978)
         );
  OAI21_X1 U10889 ( .B1(n9979), .B2(n11034), .A(n9978), .ZN(n9999) );
  MUX2_X1 U10890 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9999), .S(n11078), .Z(
        P2_U3537) );
  AOI211_X1 U10891 ( .C1(n10975), .C2(n9982), .A(n9981), .B(n9980), .ZN(n9983)
         );
  OAI21_X1 U10892 ( .B1(n9984), .B2(n11034), .A(n9983), .ZN(n10000) );
  MUX2_X1 U10893 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n10000), .S(n11078), .Z(
        P2_U3536) );
  MUX2_X1 U10894 ( .A(n9985), .B(P2_REG0_REG_31__SCAN_IN), .S(n11079), .Z(
        P2_U3519) );
  MUX2_X1 U10895 ( .A(n9986), .B(P2_REG0_REG_30__SCAN_IN), .S(n11079), .Z(
        P2_U3518) );
  MUX2_X1 U10896 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9987), .S(n11082), .Z(
        P2_U3517) );
  MUX2_X1 U10897 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9988), .S(n11082), .Z(
        P2_U3516) );
  MUX2_X1 U10898 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9989), .S(n11082), .Z(
        P2_U3515) );
  MUX2_X1 U10899 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9990), .S(n11082), .Z(
        P2_U3514) );
  MUX2_X1 U10900 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9991), .S(n11082), .Z(
        P2_U3513) );
  MUX2_X1 U10901 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9992), .S(n11082), .Z(
        P2_U3512) );
  MUX2_X1 U10902 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9993), .S(n11082), .Z(
        P2_U3511) );
  MUX2_X1 U10903 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9994), .S(n11082), .Z(
        P2_U3510) );
  MUX2_X1 U10904 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9995), .S(n11082), .Z(
        P2_U3509) );
  MUX2_X1 U10905 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9996), .S(n11082), .Z(
        P2_U3508) );
  MUX2_X1 U10906 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9997), .S(n11082), .Z(
        P2_U3507) );
  MUX2_X1 U10907 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9998), .S(n11082), .Z(
        P2_U3505) );
  MUX2_X1 U10908 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9999), .S(n11082), .Z(
        P2_U3502) );
  MUX2_X1 U10909 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n10000), .S(n11082), .Z(
        P2_U3499) );
  INV_X1 U10910 ( .A(n8774), .ZN(n10539) );
  NOR4_X1 U10911 ( .A1(n10001), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), 
        .A4(n10002), .ZN(n10003) );
  AOI21_X1 U10912 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n10010), .A(n10003), 
        .ZN(n10004) );
  OAI21_X1 U10913 ( .B1(n10539), .B2(n10012), .A(n10004), .ZN(P2_U3327) );
  OAI222_X1 U10914 ( .A1(P2_U3152), .A2(n10008), .B1(n10012), .B2(n10007), 
        .C1(n10006), .C2(n10005), .ZN(P2_U3328) );
  AOI21_X1 U10915 ( .B1(n10010), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n10009), 
        .ZN(n10011) );
  OAI21_X1 U10916 ( .B1(n10013), .B2(n10012), .A(n10011), .ZN(P2_U3330) );
  MUX2_X1 U10917 ( .A(n10014), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10918 ( .A(n10018), .ZN(n10015) );
  NOR2_X1 U10919 ( .A1(n10016), .A2(n10015), .ZN(n10021) );
  AOI21_X1 U10920 ( .B1(n10019), .B2(n10018), .A(n10017), .ZN(n10020) );
  OAI21_X1 U10921 ( .B1(n10021), .B2(n10020), .A(n10143), .ZN(n10026) );
  INV_X1 U10922 ( .A(n10022), .ZN(n10353) );
  AOI22_X1 U10923 ( .A1(n10353), .A2(n10152), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10023) );
  OAI21_X1 U10924 ( .B1(n10390), .B2(n10149), .A(n10023), .ZN(n10024) );
  AOI21_X1 U10925 ( .B1(n10159), .B2(n10147), .A(n10024), .ZN(n10025) );
  OAI211_X1 U10926 ( .C1(n10355), .C2(n10156), .A(n10026), .B(n10025), .ZN(
        P1_U3214) );
  NOR2_X1 U10927 ( .A1(n5488), .A2(n10029), .ZN(n10030) );
  XNOR2_X1 U10928 ( .A(n10027), .B(n10030), .ZN(n10035) );
  NAND2_X1 U10929 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10250)
         );
  OAI21_X1 U10930 ( .B1(n10149), .B2(n10430), .A(n10250), .ZN(n10031) );
  AOI21_X1 U10931 ( .B1(n10163), .B2(n10147), .A(n10031), .ZN(n10032) );
  OAI21_X1 U10932 ( .B1(n10098), .B2(n10436), .A(n10032), .ZN(n10033) );
  AOI21_X1 U10933 ( .B1(n10503), .B2(n10131), .A(n10033), .ZN(n10034) );
  OAI21_X1 U10934 ( .B1(n10035), .B2(n10133), .A(n10034), .ZN(P1_U3217) );
  INV_X1 U10935 ( .A(n10493), .ZN(n10047) );
  OAI21_X1 U10936 ( .B1(n5497), .B2(n10038), .A(n10037), .ZN(n10039) );
  OAI21_X1 U10937 ( .B1(n10040), .B2(n5497), .A(n10039), .ZN(n10041) );
  NAND2_X1 U10938 ( .A1(n10041), .A2(n10143), .ZN(n10046) );
  OAI22_X1 U10939 ( .A1(n10431), .A2(n10149), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10042), .ZN(n10044) );
  NOR2_X1 U10940 ( .A1(n10098), .A2(n10394), .ZN(n10043) );
  AOI211_X1 U10941 ( .C1(n10147), .C2(n10161), .A(n10044), .B(n10043), .ZN(
        n10045) );
  OAI211_X1 U10942 ( .C1(n10047), .C2(n10156), .A(n10046), .B(n10045), .ZN(
        P1_U3221) );
  XNOR2_X1 U10943 ( .A(n10050), .B(n10049), .ZN(n10051) );
  XNOR2_X1 U10944 ( .A(n10048), .B(n10051), .ZN(n10057) );
  NAND2_X1 U10945 ( .A1(n10052), .A2(n10147), .ZN(n10054) );
  AOI22_X1 U10946 ( .A1(n10327), .A2(n10152), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10053) );
  OAI211_X1 U10947 ( .C1(n10359), .C2(n10149), .A(n10054), .B(n10053), .ZN(
        n10055) );
  AOI21_X1 U10948 ( .B1(n10471), .B2(n10131), .A(n10055), .ZN(n10056) );
  OAI21_X1 U10949 ( .B1(n10057), .B2(n10133), .A(n10056), .ZN(P1_U3223) );
  NAND2_X1 U10950 ( .A1(n10058), .A2(n10059), .ZN(n10136) );
  NAND2_X1 U10951 ( .A1(n10136), .A2(n10137), .ZN(n10138) );
  NOR2_X1 U10952 ( .A1(n10058), .A2(n10059), .ZN(n10139) );
  INV_X1 U10953 ( .A(n10139), .ZN(n10060) );
  NAND2_X1 U10954 ( .A1(n10138), .A2(n10060), .ZN(n10142) );
  XNOR2_X1 U10955 ( .A(n10062), .B(n10061), .ZN(n10063) );
  XNOR2_X1 U10956 ( .A(n10142), .B(n10063), .ZN(n10071) );
  AOI22_X1 U10957 ( .A1(n10147), .A2(n10166), .B1(P1_REG3_REG_16__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10066) );
  NAND2_X1 U10958 ( .A1(n10152), .A2(n10064), .ZN(n10065) );
  OAI211_X1 U10959 ( .C1(n10067), .C2(n10149), .A(n10066), .B(n10065), .ZN(
        n10068) );
  AOI21_X1 U10960 ( .B1(n10069), .B2(n10131), .A(n10068), .ZN(n10070) );
  OAI21_X1 U10961 ( .B1(n10071), .B2(n10133), .A(n10070), .ZN(P1_U3224) );
  XNOR2_X1 U10962 ( .A(n10073), .B(n10072), .ZN(n10074) );
  XNOR2_X1 U10963 ( .A(n10075), .B(n10074), .ZN(n10082) );
  AND2_X1 U10964 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U10965 ( .A1(n10149), .A2(n10076), .ZN(n10077) );
  AOI211_X1 U10966 ( .C1(n10147), .C2(n10165), .A(n10226), .B(n10077), .ZN(
        n10078) );
  OAI21_X1 U10967 ( .B1(n10098), .B2(n10079), .A(n10078), .ZN(n10080) );
  AOI21_X1 U10968 ( .B1(n10514), .B2(n10131), .A(n10080), .ZN(n10081) );
  OAI21_X1 U10969 ( .B1(n10082), .B2(n10133), .A(n10081), .ZN(P1_U3226) );
  OAI21_X1 U10970 ( .B1(n10085), .B2(n10084), .A(n10083), .ZN(n10086) );
  NAND2_X1 U10971 ( .A1(n10086), .A2(n10143), .ZN(n10091) );
  INV_X1 U10972 ( .A(n10087), .ZN(n10345) );
  AOI22_X1 U10973 ( .A1(n10345), .A2(n10152), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10088) );
  OAI21_X1 U10974 ( .B1(n10371), .B2(n10149), .A(n10088), .ZN(n10089) );
  AOI21_X1 U10975 ( .B1(n10158), .B2(n10147), .A(n10089), .ZN(n10090) );
  OAI211_X1 U10976 ( .C1(n10347), .C2(n10156), .A(n10091), .B(n10090), .ZN(
        P1_U3227) );
  XNOR2_X1 U10977 ( .A(n10094), .B(n10093), .ZN(n10095) );
  XNOR2_X1 U10978 ( .A(n10092), .B(n10095), .ZN(n10101) );
  NAND2_X1 U10979 ( .A1(n10162), .A2(n10147), .ZN(n10097) );
  AOI22_X1 U10980 ( .A1(n10164), .A2(n10115), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10096) );
  OAI211_X1 U10981 ( .C1(n10098), .C2(n10410), .A(n10097), .B(n10096), .ZN(
        n10099) );
  AOI21_X1 U10982 ( .B1(n10496), .B2(n10131), .A(n10099), .ZN(n10100) );
  OAI21_X1 U10983 ( .B1(n10101), .B2(n10133), .A(n10100), .ZN(P1_U3231) );
  OAI21_X1 U10984 ( .B1(n10104), .B2(n10102), .A(n10103), .ZN(n10105) );
  NAND2_X1 U10985 ( .A1(n10105), .A2(n10143), .ZN(n10110) );
  OAI22_X1 U10986 ( .A1(n10402), .A2(n10149), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10106), .ZN(n10108) );
  NOR2_X1 U10987 ( .A1(n10371), .A2(n10118), .ZN(n10107) );
  AOI211_X1 U10988 ( .C1(n10379), .C2(n10152), .A(n10108), .B(n10107), .ZN(
        n10109) );
  OAI211_X1 U10989 ( .C1(n10485), .C2(n10156), .A(n10110), .B(n10109), .ZN(
        P1_U3233) );
  XOR2_X1 U10990 ( .A(n10113), .B(n10112), .Z(n10114) );
  XNOR2_X1 U10991 ( .A(n10111), .B(n10114), .ZN(n10123) );
  NAND2_X1 U10992 ( .A1(n10115), .A2(n10166), .ZN(n10117) );
  OAI211_X1 U10993 ( .C1(n10401), .C2(n10118), .A(n10117), .B(n10116), .ZN(
        n10119) );
  AOI21_X1 U10994 ( .B1(n10120), .B2(n10152), .A(n10119), .ZN(n10122) );
  NAND2_X1 U10995 ( .A1(n10507), .A2(n10131), .ZN(n10121) );
  OAI211_X1 U10996 ( .C1(n10123), .C2(n10133), .A(n10122), .B(n10121), .ZN(
        P1_U3236) );
  XNOR2_X1 U10997 ( .A(n10124), .B(n10125), .ZN(n10134) );
  NAND2_X1 U10998 ( .A1(n10126), .A2(n10147), .ZN(n10129) );
  INV_X1 U10999 ( .A(n10127), .ZN(n10312) );
  AOI22_X1 U11000 ( .A1(n10312), .A2(n10152), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3084), .ZN(n10128) );
  OAI211_X1 U11001 ( .C1(n10340), .C2(n10149), .A(n10129), .B(n10128), .ZN(
        n10130) );
  AOI21_X1 U11002 ( .B1(n10465), .B2(n10131), .A(n10130), .ZN(n10132) );
  OAI21_X1 U11003 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(P1_U3238) );
  INV_X1 U11004 ( .A(n10135), .ZN(n11061) );
  INV_X1 U11005 ( .A(n10136), .ZN(n10141) );
  OAI21_X1 U11006 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(n10140) );
  OAI21_X1 U11007 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(n10144) );
  NAND2_X1 U11008 ( .A1(n10144), .A2(n10143), .ZN(n10155) );
  AOI21_X1 U11009 ( .B1(n10147), .B2(n10146), .A(n10145), .ZN(n10148) );
  OAI21_X1 U11010 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(n10151) );
  AOI21_X1 U11011 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(n10154) );
  OAI211_X1 U11012 ( .C1(n11061), .C2(n10156), .A(n10155), .B(n10154), .ZN(
        P1_U3239) );
  MUX2_X1 U11013 ( .A(n10261), .B(P1_DATAO_REG_31__SCAN_IN), .S(n10176), .Z(
        P1_U3586) );
  MUX2_X1 U11014 ( .A(n10276), .B(P1_DATAO_REG_30__SCAN_IN), .S(n10176), .Z(
        P1_U3585) );
  MUX2_X1 U11015 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n10157), .S(P1_U4006), .Z(
        P1_U3584) );
  INV_X1 U11016 ( .A(n10297), .ZN(n10274) );
  MUX2_X1 U11017 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10274), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U11018 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10158), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U11019 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10159), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U11020 ( .A(n10160), .B(P1_DATAO_REG_23__SCAN_IN), .S(n10176), .Z(
        P1_U3578) );
  MUX2_X1 U11021 ( .A(n10161), .B(P1_DATAO_REG_22__SCAN_IN), .S(n10176), .Z(
        P1_U3577) );
  MUX2_X1 U11022 ( .A(n10162), .B(P1_DATAO_REG_21__SCAN_IN), .S(n10176), .Z(
        P1_U3576) );
  MUX2_X1 U11023 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10163), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U11024 ( .A(n10164), .B(P1_DATAO_REG_19__SCAN_IN), .S(n10176), .Z(
        P1_U3574) );
  MUX2_X1 U11025 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10165), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U11026 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10166), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U11027 ( .A(n10167), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10176), .Z(
        P1_U3568) );
  MUX2_X1 U11028 ( .A(n11005), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10176), .Z(
        P1_U3567) );
  MUX2_X1 U11029 ( .A(n10168), .B(P1_DATAO_REG_11__SCAN_IN), .S(n10176), .Z(
        P1_U3566) );
  MUX2_X1 U11030 ( .A(n10169), .B(P1_DATAO_REG_10__SCAN_IN), .S(n10176), .Z(
        P1_U3565) );
  MUX2_X1 U11031 ( .A(n10170), .B(P1_DATAO_REG_9__SCAN_IN), .S(n10176), .Z(
        P1_U3564) );
  MUX2_X1 U11032 ( .A(n10171), .B(P1_DATAO_REG_8__SCAN_IN), .S(n10176), .Z(
        P1_U3563) );
  MUX2_X1 U11033 ( .A(n10172), .B(P1_DATAO_REG_7__SCAN_IN), .S(n10176), .Z(
        P1_U3562) );
  MUX2_X1 U11034 ( .A(n10173), .B(P1_DATAO_REG_5__SCAN_IN), .S(n10176), .Z(
        P1_U3560) );
  MUX2_X1 U11035 ( .A(n10174), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10176), .Z(
        P1_U3559) );
  MUX2_X1 U11036 ( .A(n10175), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10176), .Z(
        P1_U3558) );
  MUX2_X1 U11037 ( .A(n5727), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10176), .Z(
        P1_U3557) );
  MUX2_X1 U11038 ( .A(n5704), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10176), .Z(
        P1_U3556) );
  MUX2_X1 U11039 ( .A(n7119), .B(P1_DATAO_REG_0__SCAN_IN), .S(n10176), .Z(
        P1_U3555) );
  INV_X1 U11040 ( .A(n10196), .ZN(n10181) );
  NOR3_X1 U11041 ( .A1(n10179), .A2(n10178), .A3(n10177), .ZN(n10180) );
  OAI21_X1 U11042 ( .B1(n10181), .B2(n10180), .A(n10635), .ZN(n10193) );
  INV_X1 U11043 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10182) );
  NOR2_X1 U11044 ( .A1(n10631), .A2(n10182), .ZN(n10183) );
  AOI211_X1 U11045 ( .C1(n10185), .C2(n10692), .A(n10184), .B(n10183), .ZN(
        n10192) );
  INV_X1 U11046 ( .A(n10186), .ZN(n10190) );
  INV_X1 U11047 ( .A(n10187), .ZN(n10189) );
  OAI211_X1 U11048 ( .C1(n10190), .C2(n10189), .A(n10700), .B(n10188), .ZN(
        n10191) );
  NAND3_X1 U11049 ( .A1(n10193), .A2(n10192), .A3(n10191), .ZN(P1_U3253) );
  AND3_X1 U11050 ( .A1(n10196), .A2(n10195), .A3(n10194), .ZN(n10197) );
  OAI21_X1 U11051 ( .B1(n10211), .B2(n10197), .A(n10635), .ZN(n10207) );
  INV_X1 U11052 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U11053 ( .A1(n10631), .A2(n10198), .ZN(n10199) );
  AOI211_X1 U11054 ( .C1(n10201), .C2(n10692), .A(n10200), .B(n10199), .ZN(
        n10206) );
  OAI211_X1 U11055 ( .C1(n10204), .C2(n10203), .A(n10202), .B(n10700), .ZN(
        n10205) );
  NAND3_X1 U11056 ( .A1(n10207), .A2(n10206), .A3(n10205), .ZN(P1_U3254) );
  INV_X1 U11057 ( .A(n10208), .ZN(n10213) );
  NOR3_X1 U11058 ( .A1(n10211), .A2(n10210), .A3(n10209), .ZN(n10212) );
  OAI21_X1 U11059 ( .B1(n10213), .B2(n10212), .A(n10635), .ZN(n10223) );
  INV_X1 U11060 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U11061 ( .A1(n10631), .A2(n10214), .ZN(n10215) );
  AOI211_X1 U11062 ( .C1(n10217), .C2(n10692), .A(n10216), .B(n10215), .ZN(
        n10222) );
  OAI211_X1 U11063 ( .C1(n10220), .C2(n10219), .A(n10218), .B(n10700), .ZN(
        n10221) );
  NAND3_X1 U11064 ( .A1(n10223), .A2(n10222), .A3(n10221), .ZN(P1_U3255) );
  INV_X1 U11065 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U11066 ( .A1(n10631), .A2(n10224), .ZN(n10225) );
  AOI211_X1 U11067 ( .C1(n10227), .C2(n10692), .A(n10226), .B(n10225), .ZN(
        n10237) );
  AOI211_X1 U11068 ( .C1(n10230), .C2(n10229), .A(n10228), .B(n10248), .ZN(
        n10231) );
  INV_X1 U11069 ( .A(n10231), .ZN(n10236) );
  OAI211_X1 U11070 ( .C1(n10234), .C2(n10233), .A(n10635), .B(n10232), .ZN(
        n10235) );
  NAND3_X1 U11071 ( .A1(n10237), .A2(n10236), .A3(n10235), .ZN(P1_U3258) );
  AOI21_X1 U11072 ( .B1(n10239), .B2(n8497), .A(n10238), .ZN(n10241) );
  XNOR2_X1 U11073 ( .A(n10392), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10240) );
  XNOR2_X1 U11074 ( .A(n10241), .B(n10240), .ZN(n10249) );
  INV_X1 U11075 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10242) );
  MUX2_X1 U11076 ( .A(n10242), .B(P1_REG2_REG_19__SCAN_IN), .S(n10392), .Z(
        n10246) );
  AOI21_X1 U11077 ( .B1(n10244), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10243), 
        .ZN(n10245) );
  XOR2_X1 U11078 ( .A(n10246), .B(n10245), .Z(n10247) );
  OAI22_X1 U11079 ( .A1(n10695), .A2(n10249), .B1(n10248), .B2(n10247), .ZN(
        n10253) );
  OAI21_X1 U11080 ( .B1(n10251), .B2(n10392), .A(n10250), .ZN(n10252) );
  AOI211_X1 U11081 ( .C1(P1_ADDR_REG_19__SCAN_IN), .C2(n10698), .A(n10253), 
        .B(n10252), .ZN(n10254) );
  INV_X1 U11082 ( .A(n10254), .ZN(P1_U3260) );
  INV_X1 U11083 ( .A(n10449), .ZN(n10267) );
  INV_X1 U11084 ( .A(n10256), .ZN(n10280) );
  NAND2_X1 U11085 ( .A1(n10267), .A2(n10279), .ZN(n10257) );
  XNOR2_X1 U11086 ( .A(n10445), .B(n10257), .ZN(n10443) );
  NAND2_X1 U11087 ( .A1(n10443), .A2(n11022), .ZN(n10263) );
  INV_X1 U11088 ( .A(P1_B_REG_SCAN_IN), .ZN(n10258) );
  NOR2_X1 U11089 ( .A1(n10259), .A2(n10258), .ZN(n10260) );
  NOR2_X1 U11090 ( .A1(n10851), .A2(n10260), .ZN(n10275) );
  NAND2_X1 U11091 ( .A1(n10261), .A2(n10275), .ZN(n10447) );
  NOR2_X1 U11092 ( .A1(n11027), .A2(n10447), .ZN(n10264) );
  AOI21_X1 U11093 ( .B1(n11027), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10264), 
        .ZN(n10262) );
  OAI211_X1 U11094 ( .C1(n10445), .C2(n11029), .A(n10263), .B(n10262), .ZN(
        P1_U3261) );
  XNOR2_X1 U11095 ( .A(n10449), .B(n10279), .ZN(n10446) );
  NAND2_X1 U11096 ( .A1(n10446), .A2(n11022), .ZN(n10266) );
  AOI21_X1 U11097 ( .B1(n11027), .B2(P1_REG2_REG_30__SCAN_IN), .A(n10264), 
        .ZN(n10265) );
  OAI211_X1 U11098 ( .C1(n10267), .C2(n11029), .A(n10266), .B(n10265), .ZN(
        P1_U3262) );
  NAND2_X1 U11099 ( .A1(n10271), .A2(n10270), .ZN(n10273) );
  NAND2_X1 U11100 ( .A1(n10274), .A2(n11006), .ZN(n10278) );
  NAND2_X1 U11101 ( .A1(n10276), .A2(n10275), .ZN(n10277) );
  OR2_X1 U11102 ( .A1(n10453), .A2(n11027), .ZN(n10286) );
  AOI21_X1 U11103 ( .B1(n10255), .B2(n10280), .A(n10279), .ZN(n10452) );
  AOI22_X1 U11104 ( .A1(n10281), .A2(n11025), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n11027), .ZN(n10282) );
  OAI21_X1 U11105 ( .B1(n10283), .B2(n11029), .A(n10282), .ZN(n10284) );
  AOI21_X1 U11106 ( .B1(n10452), .B2(n11022), .A(n10284), .ZN(n10285) );
  OAI211_X1 U11107 ( .C1(n10442), .C2(n10454), .A(n10286), .B(n10285), .ZN(
        P1_U3355) );
  XNOR2_X1 U11108 ( .A(n10287), .B(n10296), .ZN(n10464) );
  INV_X1 U11109 ( .A(n10311), .ZN(n10290) );
  INV_X1 U11110 ( .A(n10288), .ZN(n10289) );
  AOI211_X1 U11111 ( .C1(n10461), .C2(n10290), .A(n11085), .B(n10289), .ZN(
        n10460) );
  AOI22_X1 U11112 ( .A1(n10291), .A2(n11025), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n11027), .ZN(n10292) );
  OAI21_X1 U11113 ( .B1(n10293), .B2(n11029), .A(n10292), .ZN(n10301) );
  AOI211_X1 U11114 ( .C1(n10296), .C2(n10295), .A(n10429), .B(n10294), .ZN(
        n10299) );
  OAI22_X1 U11115 ( .A1(n10297), .A2(n10851), .B1(n10323), .B2(n10849), .ZN(
        n10298) );
  NOR2_X1 U11116 ( .A1(n10299), .A2(n10298), .ZN(n10463) );
  NOR2_X1 U11117 ( .A1(n10463), .A2(n11027), .ZN(n10300) );
  AOI211_X1 U11118 ( .C1(n10439), .C2(n10460), .A(n10301), .B(n10300), .ZN(
        n10302) );
  OAI21_X1 U11119 ( .B1(n10464), .B2(n10442), .A(n10302), .ZN(P1_U3264) );
  OAI21_X1 U11120 ( .B1(n10306), .B2(n10304), .A(n10303), .ZN(n10310) );
  OAI22_X1 U11121 ( .A1(n10305), .A2(n10851), .B1(n10340), .B2(n10849), .ZN(
        n10309) );
  XNOR2_X1 U11122 ( .A(n10307), .B(n10306), .ZN(n10469) );
  NOR2_X1 U11123 ( .A1(n10469), .A2(n11013), .ZN(n10308) );
  AOI21_X1 U11124 ( .B1(n10465), .B2(n10319), .A(n10311), .ZN(n10466) );
  AOI22_X1 U11125 ( .A1(n10312), .A2(n11025), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n11027), .ZN(n10313) );
  OAI21_X1 U11126 ( .B1(n10314), .B2(n11029), .A(n10313), .ZN(n10316) );
  NOR2_X1 U11127 ( .A1(n10469), .A2(n10419), .ZN(n10315) );
  AOI211_X1 U11128 ( .C1(n10466), .C2(n11022), .A(n10316), .B(n10315), .ZN(
        n10317) );
  OAI21_X1 U11129 ( .B1(n10468), .B2(n11027), .A(n10317), .ZN(P1_U3265) );
  XNOR2_X1 U11130 ( .A(n10318), .B(n5304), .ZN(n10474) );
  AOI211_X1 U11131 ( .C1(n10471), .C2(n10334), .A(n11085), .B(n8996), .ZN(
        n10470) );
  INV_X1 U11132 ( .A(n10470), .ZN(n10326) );
  AOI211_X1 U11133 ( .C1(n10322), .C2(n10321), .A(n10429), .B(n10320), .ZN(
        n10325) );
  OAI22_X1 U11134 ( .A1(n10323), .A2(n10851), .B1(n10359), .B2(n10849), .ZN(
        n10324) );
  NOR2_X1 U11135 ( .A1(n10325), .A2(n10324), .ZN(n10473) );
  OAI21_X1 U11136 ( .B1(n10344), .B2(n10326), .A(n10473), .ZN(n10331) );
  INV_X1 U11137 ( .A(n10471), .ZN(n10329) );
  AOI22_X1 U11138 ( .A1(n10327), .A2(n11025), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n11027), .ZN(n10328) );
  OAI21_X1 U11139 ( .B1(n10329), .B2(n11029), .A(n10328), .ZN(n10330) );
  AOI21_X1 U11140 ( .B1(n10331), .B2(n10869), .A(n10330), .ZN(n10332) );
  OAI21_X1 U11141 ( .B1(n10474), .B2(n10442), .A(n10332), .ZN(P1_U3266) );
  XNOR2_X1 U11142 ( .A(n10333), .B(n10338), .ZN(n10479) );
  INV_X1 U11143 ( .A(n10352), .ZN(n10336) );
  INV_X1 U11144 ( .A(n10334), .ZN(n10335) );
  AOI211_X1 U11145 ( .C1(n10476), .C2(n10336), .A(n11085), .B(n10335), .ZN(
        n10475) );
  INV_X1 U11146 ( .A(n10475), .ZN(n10343) );
  AOI211_X1 U11147 ( .C1(n10339), .C2(n10338), .A(n10429), .B(n10337), .ZN(
        n10342) );
  OAI22_X1 U11148 ( .A1(n10340), .A2(n10851), .B1(n10371), .B2(n10849), .ZN(
        n10341) );
  NOR2_X1 U11149 ( .A1(n10342), .A2(n10341), .ZN(n10478) );
  OAI21_X1 U11150 ( .B1(n10344), .B2(n10343), .A(n10478), .ZN(n10349) );
  AOI22_X1 U11151 ( .A1(n10345), .A2(n11025), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n11027), .ZN(n10346) );
  OAI21_X1 U11152 ( .B1(n10347), .B2(n11029), .A(n10346), .ZN(n10348) );
  AOI21_X1 U11153 ( .B1(n10349), .B2(n10869), .A(n10348), .ZN(n10350) );
  OAI21_X1 U11154 ( .B1(n10442), .B2(n10479), .A(n10350), .ZN(P1_U3267) );
  XNOR2_X1 U11155 ( .A(n10351), .B(n10358), .ZN(n10484) );
  AOI211_X1 U11156 ( .C1(n10481), .C2(n5337), .A(n11085), .B(n10352), .ZN(
        n10480) );
  AOI22_X1 U11157 ( .A1(n10353), .A2(n11025), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n11027), .ZN(n10354) );
  OAI21_X1 U11158 ( .B1(n10355), .B2(n11029), .A(n10354), .ZN(n10363) );
  AOI211_X1 U11159 ( .C1(n10358), .C2(n10357), .A(n10429), .B(n10356), .ZN(
        n10361) );
  OAI22_X1 U11160 ( .A1(n10359), .A2(n10851), .B1(n10390), .B2(n10849), .ZN(
        n10360) );
  NOR2_X1 U11161 ( .A1(n10361), .A2(n10360), .ZN(n10483) );
  NOR2_X1 U11162 ( .A1(n10483), .A2(n11027), .ZN(n10362) );
  AOI211_X1 U11163 ( .C1(n10480), .C2(n10439), .A(n10363), .B(n10362), .ZN(
        n10364) );
  OAI21_X1 U11164 ( .B1(n10442), .B2(n10484), .A(n10364), .ZN(P1_U3268) );
  OR2_X1 U11165 ( .A1(n10365), .A2(n10369), .ZN(n10366) );
  NAND2_X1 U11166 ( .A1(n10367), .A2(n10366), .ZN(n10490) );
  XNOR2_X1 U11167 ( .A(n10368), .B(n10369), .ZN(n10370) );
  NAND2_X1 U11168 ( .A1(n10370), .A2(n11009), .ZN(n10374) );
  OAI22_X1 U11169 ( .A1(n10371), .A2(n10851), .B1(n10402), .B2(n10849), .ZN(
        n10372) );
  INV_X1 U11170 ( .A(n10372), .ZN(n10373) );
  NAND2_X1 U11171 ( .A1(n10374), .A2(n10373), .ZN(n10488) );
  AND2_X1 U11172 ( .A1(n10375), .A2(n5623), .ZN(n10377) );
  OR2_X1 U11173 ( .A1(n10377), .A2(n10376), .ZN(n10486) );
  NOR2_X1 U11174 ( .A1(n10486), .A2(n10378), .ZN(n10382) );
  AOI22_X1 U11175 ( .A1(n10379), .A2(n11025), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n11027), .ZN(n10380) );
  OAI21_X1 U11176 ( .B1(n10485), .B2(n11029), .A(n10380), .ZN(n10381) );
  AOI211_X1 U11177 ( .C1(n10488), .C2(n10869), .A(n10382), .B(n10381), .ZN(
        n10383) );
  OAI21_X1 U11178 ( .B1(n10490), .B2(n10442), .A(n10383), .ZN(P1_U3269) );
  OAI21_X1 U11179 ( .B1(n10386), .B2(n10385), .A(n10384), .ZN(n10495) );
  AOI22_X1 U11180 ( .A1(n10493), .A2(n10413), .B1(n11027), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n10397) );
  XNOR2_X1 U11181 ( .A(n10387), .B(n10388), .ZN(n10389) );
  OAI222_X1 U11182 ( .A1(n10851), .A2(n10390), .B1(n10849), .B2(n10431), .C1(
        n10429), .C2(n10389), .ZN(n10491) );
  AOI21_X1 U11183 ( .B1(n10416), .B2(n10493), .A(n11085), .ZN(n10391) );
  AND2_X1 U11184 ( .A1(n10391), .A2(n5623), .ZN(n10492) );
  NAND2_X1 U11185 ( .A1(n10492), .A2(n10392), .ZN(n10393) );
  OAI21_X1 U11186 ( .B1(n10865), .B2(n10394), .A(n10393), .ZN(n10395) );
  OAI21_X1 U11187 ( .B1(n10491), .B2(n10395), .A(n10869), .ZN(n10396) );
  OAI211_X1 U11188 ( .C1(n10495), .C2(n10442), .A(n10397), .B(n10396), .ZN(
        P1_U3270) );
  NAND2_X1 U11189 ( .A1(n10425), .A2(n10398), .ZN(n10400) );
  XNOR2_X1 U11190 ( .A(n10400), .B(n10399), .ZN(n10409) );
  OAI22_X1 U11191 ( .A1(n10402), .A2(n10851), .B1(n10401), .B2(n10849), .ZN(
        n10408) );
  OR2_X1 U11192 ( .A1(n10404), .A2(n10403), .ZN(n10406) );
  NAND2_X1 U11193 ( .A1(n10406), .A2(n10405), .ZN(n10500) );
  NOR2_X1 U11194 ( .A1(n10500), .A2(n11013), .ZN(n10407) );
  AOI211_X1 U11195 ( .C1(n10409), .C2(n11009), .A(n10408), .B(n10407), .ZN(
        n10499) );
  INV_X1 U11196 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10411) );
  OAI22_X1 U11197 ( .A1(n10869), .A2(n10411), .B1(n10410), .B2(n10865), .ZN(
        n10412) );
  AOI21_X1 U11198 ( .B1(n10496), .B2(n10413), .A(n10412), .ZN(n10418) );
  OR2_X1 U11199 ( .A1(n10433), .A2(n10414), .ZN(n10415) );
  AND2_X1 U11200 ( .A1(n10416), .A2(n10415), .ZN(n10497) );
  NAND2_X1 U11201 ( .A1(n10497), .A2(n11022), .ZN(n10417) );
  OAI211_X1 U11202 ( .C1(n10500), .C2(n10419), .A(n10418), .B(n10417), .ZN(
        n10420) );
  INV_X1 U11203 ( .A(n10420), .ZN(n10421) );
  OAI21_X1 U11204 ( .B1(n10499), .B2(n11027), .A(n10421), .ZN(P1_U3271) );
  OAI21_X1 U11205 ( .B1(n10423), .B2(n10427), .A(n10422), .ZN(n10505) );
  INV_X1 U11206 ( .A(n10425), .ZN(n10426) );
  AOI21_X1 U11207 ( .B1(n10427), .B2(n10424), .A(n10426), .ZN(n10428) );
  OAI222_X1 U11208 ( .A1(n10851), .A2(n10431), .B1(n10849), .B2(n10430), .C1(
        n10429), .C2(n10428), .ZN(n10501) );
  NAND2_X1 U11209 ( .A1(n10501), .A2(n10869), .ZN(n10441) );
  INV_X1 U11210 ( .A(n10432), .ZN(n10434) );
  AOI211_X1 U11211 ( .C1(n10503), .C2(n10434), .A(n11085), .B(n10433), .ZN(
        n10502) );
  NOR2_X1 U11212 ( .A1(n10435), .A2(n11029), .ZN(n10438) );
  OAI22_X1 U11213 ( .A1(n10869), .A2(n10242), .B1(n10436), .B2(n10865), .ZN(
        n10437) );
  AOI211_X1 U11214 ( .C1(n10502), .C2(n10439), .A(n10438), .B(n10437), .ZN(
        n10440) );
  OAI211_X1 U11215 ( .C1(n10505), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        P1_U3272) );
  NAND2_X1 U11216 ( .A1(n10443), .A2(n10515), .ZN(n10444) );
  OAI211_X1 U11217 ( .C1(n10445), .C2(n11083), .A(n10444), .B(n10447), .ZN(
        n10520) );
  MUX2_X1 U11218 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10520), .S(n11093), .Z(
        P1_U3554) );
  NAND2_X1 U11219 ( .A1(n10446), .A2(n10515), .ZN(n10451) );
  INV_X1 U11220 ( .A(n10447), .ZN(n10448) );
  AOI21_X1 U11221 ( .B1(n10449), .B2(n10739), .A(n10448), .ZN(n10450) );
  NAND2_X1 U11222 ( .A1(n10451), .A2(n10450), .ZN(n10521) );
  MUX2_X1 U11223 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10521), .S(n11093), .Z(
        P1_U3553) );
  AOI22_X1 U11224 ( .A1(n10456), .A2(n10515), .B1(n10739), .B2(n10455), .ZN(
        n10457) );
  MUX2_X1 U11225 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10522), .S(n11093), .Z(
        P1_U3551) );
  AOI21_X1 U11226 ( .B1(n10739), .B2(n10461), .A(n10460), .ZN(n10462) );
  OAI211_X1 U11227 ( .C1(n11059), .C2(n10464), .A(n10463), .B(n10462), .ZN(
        n10523) );
  MUX2_X1 U11228 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10523), .S(n11093), .Z(
        P1_U3550) );
  AOI22_X1 U11229 ( .A1(n10466), .A2(n10515), .B1(n10739), .B2(n10465), .ZN(
        n10467) );
  OAI211_X1 U11230 ( .C1(n10469), .C2(n10741), .A(n10468), .B(n10467), .ZN(
        n10524) );
  MUX2_X1 U11231 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10524), .S(n11093), .Z(
        P1_U3549) );
  AOI21_X1 U11232 ( .B1(n10739), .B2(n10471), .A(n10470), .ZN(n10472) );
  OAI211_X1 U11233 ( .C1(n11059), .C2(n10474), .A(n10473), .B(n10472), .ZN(
        n10525) );
  MUX2_X1 U11234 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10525), .S(n11093), .Z(
        P1_U3548) );
  AOI21_X1 U11235 ( .B1(n10739), .B2(n10476), .A(n10475), .ZN(n10477) );
  OAI211_X1 U11236 ( .C1(n11059), .C2(n10479), .A(n10478), .B(n10477), .ZN(
        n10526) );
  MUX2_X1 U11237 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10526), .S(n11093), .Z(
        P1_U3547) );
  AOI21_X1 U11238 ( .B1(n10739), .B2(n10481), .A(n10480), .ZN(n10482) );
  OAI211_X1 U11239 ( .C1(n10484), .C2(n11059), .A(n10483), .B(n10482), .ZN(
        n10527) );
  MUX2_X1 U11240 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10527), .S(n11093), .Z(
        P1_U3546) );
  OAI22_X1 U11241 ( .A1(n10486), .A2(n11085), .B1(n10485), .B2(n11083), .ZN(
        n10487) );
  NOR2_X1 U11242 ( .A1(n10488), .A2(n10487), .ZN(n10489) );
  OAI21_X1 U11243 ( .B1(n10490), .B2(n11059), .A(n10489), .ZN(n10528) );
  MUX2_X1 U11244 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10528), .S(n11093), .Z(
        P1_U3545) );
  AOI211_X1 U11245 ( .C1(n10739), .C2(n10493), .A(n10492), .B(n10491), .ZN(
        n10494) );
  OAI21_X1 U11246 ( .B1(n11059), .B2(n10495), .A(n10494), .ZN(n10529) );
  MUX2_X1 U11247 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10529), .S(n11093), .Z(
        P1_U3544) );
  AOI22_X1 U11248 ( .A1(n10497), .A2(n10515), .B1(n10739), .B2(n10496), .ZN(
        n10498) );
  OAI211_X1 U11249 ( .C1(n10741), .C2(n10500), .A(n10499), .B(n10498), .ZN(
        n10530) );
  MUX2_X1 U11250 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10530), .S(n11093), .Z(
        P1_U3543) );
  AOI211_X1 U11251 ( .C1(n10739), .C2(n10503), .A(n10502), .B(n10501), .ZN(
        n10504) );
  OAI21_X1 U11252 ( .B1(n11059), .B2(n10505), .A(n10504), .ZN(n10531) );
  MUX2_X1 U11253 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10531), .S(n11093), .Z(
        P1_U3542) );
  AOI21_X1 U11254 ( .B1(n10739), .B2(n10507), .A(n10506), .ZN(n10511) );
  INV_X1 U11255 ( .A(n11059), .ZN(n11089) );
  NAND3_X1 U11256 ( .A1(n10509), .A2(n11089), .A3(n10508), .ZN(n10510) );
  NAND3_X1 U11257 ( .A1(n10512), .A2(n10511), .A3(n10510), .ZN(n10532) );
  MUX2_X1 U11258 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10532), .S(n11093), .Z(
        P1_U3541) );
  INV_X1 U11259 ( .A(n10513), .ZN(n10519) );
  AOI22_X1 U11260 ( .A1(n10516), .A2(n10515), .B1(n10739), .B2(n10514), .ZN(
        n10517) );
  OAI211_X1 U11261 ( .C1(n10519), .C2(n10741), .A(n10518), .B(n10517), .ZN(
        n10533) );
  MUX2_X1 U11262 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10533), .S(n11093), .Z(
        P1_U3540) );
  MUX2_X1 U11263 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10520), .S(n11097), .Z(
        P1_U3522) );
  MUX2_X1 U11264 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10521), .S(n11097), .Z(
        P1_U3521) );
  MUX2_X1 U11265 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10522), .S(n11097), .Z(
        P1_U3519) );
  MUX2_X1 U11266 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10523), .S(n11097), .Z(
        P1_U3518) );
  MUX2_X1 U11267 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10524), .S(n11097), .Z(
        P1_U3517) );
  MUX2_X1 U11268 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10525), .S(n11097), .Z(
        P1_U3516) );
  MUX2_X1 U11269 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10526), .S(n11097), .Z(
        P1_U3515) );
  MUX2_X1 U11270 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10527), .S(n11097), .Z(
        P1_U3514) );
  MUX2_X1 U11271 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10528), .S(n11097), .Z(
        P1_U3513) );
  MUX2_X1 U11272 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10529), .S(n11097), .Z(
        P1_U3512) );
  MUX2_X1 U11273 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10530), .S(n11097), .Z(
        P1_U3511) );
  MUX2_X1 U11274 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10531), .S(n11097), .Z(
        P1_U3510) );
  MUX2_X1 U11275 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10532), .S(n11097), .Z(
        P1_U3508) );
  MUX2_X1 U11276 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10533), .S(n11097), .Z(
        P1_U3505) );
  NOR4_X1 U11277 ( .A1(n10535), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n10534), .ZN(n10536) );
  AOI21_X1 U11278 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10537), .A(n10536), 
        .ZN(n10538) );
  OAI21_X1 U11279 ( .B1(n10539), .B2(n5033), .A(n10538), .ZN(P1_U3322) );
  INV_X1 U11280 ( .A(n10540), .ZN(n10541) );
  MUX2_X1 U11281 ( .A(n10541), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11282 ( .A(n10545), .ZN(n10544) );
  NOR2_X1 U11283 ( .A1(n10544), .A2(n10542), .ZN(P1_U3321) );
  NOR2_X1 U11284 ( .A1(n10544), .A2(n10543), .ZN(P1_U3320) );
  AND2_X1 U11285 ( .A1(n10545), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  AND2_X1 U11286 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10545), .ZN(P1_U3318) );
  AND2_X1 U11287 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10545), .ZN(P1_U3317) );
  AND2_X1 U11288 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10545), .ZN(P1_U3316) );
  AND2_X1 U11289 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10545), .ZN(P1_U3315) );
  AND2_X1 U11290 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10545), .ZN(P1_U3314) );
  AND2_X1 U11291 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10545), .ZN(P1_U3313) );
  AND2_X1 U11292 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10545), .ZN(P1_U3312) );
  AND2_X1 U11293 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10545), .ZN(P1_U3311) );
  AND2_X1 U11294 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10545), .ZN(P1_U3310) );
  AND2_X1 U11295 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10545), .ZN(P1_U3309) );
  AND2_X1 U11296 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10545), .ZN(P1_U3308) );
  AND2_X1 U11297 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10545), .ZN(P1_U3307) );
  AND2_X1 U11298 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10545), .ZN(P1_U3306) );
  AND2_X1 U11299 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10545), .ZN(P1_U3305) );
  AND2_X1 U11300 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10545), .ZN(P1_U3304) );
  AND2_X1 U11301 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10545), .ZN(P1_U3303) );
  AND2_X1 U11302 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10545), .ZN(P1_U3302) );
  AND2_X1 U11303 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10545), .ZN(P1_U3301) );
  AND2_X1 U11304 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10545), .ZN(P1_U3300) );
  AND2_X1 U11305 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10545), .ZN(P1_U3299) );
  AND2_X1 U11306 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10545), .ZN(P1_U3298) );
  AND2_X1 U11307 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10545), .ZN(P1_U3297) );
  AND2_X1 U11308 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10545), .ZN(P1_U3296) );
  AND2_X1 U11309 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10545), .ZN(P1_U3295) );
  AND2_X1 U11310 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10545), .ZN(P1_U3294) );
  AND2_X1 U11311 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10545), .ZN(P1_U3293) );
  AND2_X1 U11312 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10545), .ZN(P1_U3292) );
  AOI22_X1 U11313 ( .A1(n10648), .A2(n10549), .B1(n10548), .B2(n10645), .ZN(
        P2_U3438) );
  AND2_X1 U11314 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10645), .ZN(P2_U3326) );
  AND2_X1 U11315 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10645), .ZN(P2_U3325) );
  AND2_X1 U11316 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10645), .ZN(P2_U3324) );
  AND2_X1 U11317 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10645), .ZN(P2_U3323) );
  AND2_X1 U11318 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10645), .ZN(P2_U3322) );
  AND2_X1 U11319 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10645), .ZN(P2_U3321) );
  AND2_X1 U11320 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10645), .ZN(P2_U3320) );
  AND2_X1 U11321 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10645), .ZN(P2_U3319) );
  AND2_X1 U11322 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10645), .ZN(P2_U3318) );
  AND2_X1 U11323 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10645), .ZN(P2_U3317) );
  AND2_X1 U11324 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10645), .ZN(P2_U3316) );
  AND2_X1 U11325 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10645), .ZN(P2_U3315) );
  AND2_X1 U11326 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10645), .ZN(P2_U3314) );
  AND2_X1 U11327 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10645), .ZN(P2_U3313) );
  AND2_X1 U11328 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10645), .ZN(P2_U3312) );
  AND2_X1 U11329 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10645), .ZN(P2_U3311) );
  AND2_X1 U11330 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10645), .ZN(P2_U3310) );
  AND2_X1 U11331 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10645), .ZN(P2_U3309) );
  AND2_X1 U11332 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10645), .ZN(P2_U3308) );
  AND2_X1 U11333 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10645), .ZN(P2_U3307) );
  AND2_X1 U11334 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10645), .ZN(P2_U3306) );
  AND2_X1 U11335 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10645), .ZN(P2_U3305) );
  AND2_X1 U11336 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10645), .ZN(P2_U3304) );
  AND2_X1 U11337 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10645), .ZN(P2_U3303) );
  AND2_X1 U11338 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10645), .ZN(P2_U3302) );
  AND2_X1 U11339 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10645), .ZN(P2_U3301) );
  AND2_X1 U11340 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10645), .ZN(P2_U3300) );
  AND2_X1 U11341 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10645), .ZN(P2_U3299) );
  AND2_X1 U11342 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10645), .ZN(P2_U3298) );
  AND2_X1 U11343 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10645), .ZN(P2_U3297) );
  XOR2_X1 U11344 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11345 ( .A(n10550), .ZN(n10551) );
  NAND2_X1 U11346 ( .A1(n10552), .A2(n10551), .ZN(n10553) );
  XOR2_X1 U11347 ( .A(n10554), .B(n10553), .Z(ADD_1071_U5) );
  XOR2_X1 U11348 ( .A(n10556), .B(n10555), .Z(ADD_1071_U54) );
  XOR2_X1 U11349 ( .A(n10558), .B(n10557), .Z(ADD_1071_U53) );
  XNOR2_X1 U11350 ( .A(n10560), .B(n10559), .ZN(ADD_1071_U52) );
  NOR2_X1 U11351 ( .A1(n10562), .A2(n10561), .ZN(n10563) );
  XOR2_X1 U11352 ( .A(n10563), .B(P2_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11353 ( .A(n10564), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U11354 ( .A(n10565), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11355 ( .A(n10566), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  XNOR2_X1 U11356 ( .A(n10568), .B(n10567), .ZN(ADD_1071_U47) );
  XOR2_X1 U11357 ( .A(n10570), .B(n10569), .Z(ADD_1071_U63) );
  XOR2_X1 U11358 ( .A(n10572), .B(n10571), .Z(ADD_1071_U62) );
  XNOR2_X1 U11359 ( .A(n10574), .B(n10573), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11360 ( .A(n10576), .B(n10575), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11361 ( .A(n10578), .B(n10577), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11362 ( .A(n10580), .B(n10579), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11363 ( .A(n10582), .B(n10581), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11364 ( .A(n10584), .B(n10583), .ZN(ADD_1071_U56) );
  NOR2_X1 U11365 ( .A1(n10586), .A2(n10585), .ZN(n10587) );
  XNOR2_X1 U11366 ( .A(n10588), .B(n10587), .ZN(ADD_1071_U55) );
  OAI21_X1 U11367 ( .B1(n10590), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10589), .ZN(
        n10591) );
  XNOR2_X1 U11368 ( .A(n10591), .B(n10633), .ZN(n10594) );
  AOI22_X1 U11369 ( .A1(n10698), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10592) );
  OAI21_X1 U11370 ( .B1(n10594), .B2(n10593), .A(n10592), .ZN(P1_U3241) );
  INV_X1 U11371 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U11372 ( .A1(n10692), .A2(n10595), .ZN(n10598) );
  INV_X1 U11373 ( .A(n10596), .ZN(n10597) );
  OAI211_X1 U11374 ( .C1(n10631), .C2(n10599), .A(n10598), .B(n10597), .ZN(
        n10600) );
  INV_X1 U11375 ( .A(n10600), .ZN(n10609) );
  OAI211_X1 U11376 ( .C1(n10603), .C2(n10602), .A(n10601), .B(n10635), .ZN(
        n10608) );
  OAI211_X1 U11377 ( .C1(n10606), .C2(n10605), .A(n10604), .B(n10700), .ZN(
        n10607) );
  NAND3_X1 U11378 ( .A1(n10609), .A2(n10608), .A3(n10607), .ZN(P1_U3247) );
  INV_X1 U11379 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U11380 ( .A1(n10692), .A2(n10610), .ZN(n10613) );
  INV_X1 U11381 ( .A(n10611), .ZN(n10612) );
  OAI211_X1 U11382 ( .C1(n10631), .C2(n10614), .A(n10613), .B(n10612), .ZN(
        n10615) );
  INV_X1 U11383 ( .A(n10615), .ZN(n10624) );
  OAI211_X1 U11384 ( .C1(n10618), .C2(n10617), .A(n10635), .B(n10616), .ZN(
        n10623) );
  OAI211_X1 U11385 ( .C1(n10621), .C2(n10620), .A(n10700), .B(n10619), .ZN(
        n10622) );
  NAND3_X1 U11386 ( .A1(n10624), .A2(n10623), .A3(n10622), .ZN(P1_U3244) );
  INV_X1 U11387 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10630) );
  INV_X1 U11388 ( .A(n10625), .ZN(n10626) );
  NAND2_X1 U11389 ( .A1(n10692), .A2(n10626), .ZN(n10629) );
  NAND2_X1 U11390 ( .A1(P1_U3084), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10628) );
  OAI211_X1 U11391 ( .C1(n10631), .C2(n10630), .A(n10629), .B(n10628), .ZN(
        n10632) );
  INV_X1 U11392 ( .A(n10632), .ZN(n10643) );
  NOR2_X1 U11393 ( .A1(n10633), .A2(n5666), .ZN(n10637) );
  OAI211_X1 U11394 ( .C1(n10637), .C2(n10636), .A(n10635), .B(n10634), .ZN(
        n10642) );
  OAI211_X1 U11395 ( .C1(n10640), .C2(n10639), .A(n10700), .B(n10638), .ZN(
        n10641) );
  NAND3_X1 U11396 ( .A1(n10643), .A2(n10642), .A3(n10641), .ZN(P1_U3242) );
  INV_X1 U11397 ( .A(n10644), .ZN(n10647) );
  INV_X1 U11398 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U11399 ( .A1(n10648), .A2(n10647), .B1(n10646), .B2(n10645), .ZN(
        P2_U3437) );
  AOI22_X1 U11400 ( .A1(n10651), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n10649), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U11401 ( .A1(n10672), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10656) );
  NAND2_X1 U11402 ( .A1(n10651), .A2(n10650), .ZN(n10652) );
  OAI211_X1 U11403 ( .C1(n10673), .C2(P2_REG1_REG_0__SCAN_IN), .A(n10653), .B(
        n10652), .ZN(n10654) );
  NAND2_X1 U11404 ( .A1(n10654), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10655) );
  OAI211_X1 U11405 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10657), .A(n10656), .B(
        n10655), .ZN(P2_U3245) );
  AOI21_X1 U11406 ( .B1(n10672), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n10659), .ZN(
        n10670) );
  AOI211_X1 U11407 ( .C1(n10662), .C2(n10661), .A(n10660), .B(n10673), .ZN(
        n10667) );
  AOI211_X1 U11408 ( .C1(n10665), .C2(n10664), .A(n10663), .B(n10677), .ZN(
        n10666) );
  AOI211_X1 U11409 ( .C1(n10684), .C2(n10668), .A(n10667), .B(n10666), .ZN(
        n10669) );
  NAND2_X1 U11410 ( .A1(n10670), .A2(n10669), .ZN(P2_U3246) );
  AOI21_X1 U11411 ( .B1(n10672), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n10671), .ZN(
        n10686) );
  AOI211_X1 U11412 ( .C1(n10676), .C2(n10675), .A(n10674), .B(n10673), .ZN(
        n10682) );
  AOI211_X1 U11413 ( .C1(n10680), .C2(n10679), .A(n10678), .B(n10677), .ZN(
        n10681) );
  AOI211_X1 U11414 ( .C1(n10684), .C2(n10683), .A(n10682), .B(n10681), .ZN(
        n10685) );
  NAND2_X1 U11415 ( .A1(n10686), .A2(n10685), .ZN(P2_U3247) );
  XOR2_X1 U11416 ( .A(n10687), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  INV_X1 U11417 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10705) );
  OAI21_X1 U11418 ( .B1(n10690), .B2(n10689), .A(n10688), .ZN(n10694) );
  NAND2_X1 U11419 ( .A1(n10692), .A2(n10691), .ZN(n10693) );
  OAI21_X1 U11420 ( .B1(n10695), .B2(n10694), .A(n10693), .ZN(n10697) );
  AOI211_X1 U11421 ( .C1(n10698), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n10697), .B(
        n10696), .ZN(n10704) );
  OAI211_X1 U11422 ( .C1(n10702), .C2(n10701), .A(n10700), .B(n10699), .ZN(
        n10703) );
  OAI211_X1 U11423 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n10705), .A(n10704), .B(
        n10703), .ZN(P1_U3243) );
  AOI22_X1 U11424 ( .A1(n10708), .A2(n11074), .B1(n10707), .B2(n10706), .ZN(
        n10709) );
  AND2_X1 U11425 ( .A1(n10710), .A2(n10709), .ZN(n10713) );
  INV_X1 U11426 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U11427 ( .A1(n11078), .A2(n10713), .B1(n10711), .B2(n11076), .ZN(
        P2_U3520) );
  INV_X1 U11428 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U11429 ( .A1(n11082), .A2(n10713), .B1(n10712), .B2(n11079), .ZN(
        P2_U3451) );
  INV_X1 U11430 ( .A(n10741), .ZN(n11016) );
  INV_X1 U11431 ( .A(n10714), .ZN(n10719) );
  OAI21_X1 U11432 ( .B1(n10716), .B2(n11083), .A(n10715), .ZN(n10718) );
  AOI211_X1 U11433 ( .C1(n11016), .C2(n10719), .A(n10718), .B(n10717), .ZN(
        n10722) );
  AOI22_X1 U11434 ( .A1(n11093), .A2(n10722), .B1(n10720), .B2(n11091), .ZN(
        P1_U3524) );
  INV_X1 U11435 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U11436 ( .A1(n11097), .A2(n10722), .B1(n10721), .B2(n11094), .ZN(
        P1_U3457) );
  OAI21_X1 U11437 ( .B1(n10724), .B2(n11083), .A(n10723), .ZN(n10726) );
  AOI211_X1 U11438 ( .C1(n11016), .C2(n10727), .A(n10726), .B(n10725), .ZN(
        n10729) );
  AOI22_X1 U11439 ( .A1(n11093), .A2(n10729), .B1(n7456), .B2(n11091), .ZN(
        P1_U3525) );
  INV_X1 U11440 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U11441 ( .A1(n11097), .A2(n10729), .B1(n10728), .B2(n11094), .ZN(
        P1_U3460) );
  OAI22_X1 U11442 ( .A1(n10730), .A2(n11070), .B1(n8190), .B2(n11069), .ZN(
        n10732) );
  AOI211_X1 U11443 ( .C1(n10948), .C2(n10733), .A(n10732), .B(n10731), .ZN(
        n10736) );
  INV_X1 U11444 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U11445 ( .A1(n11078), .A2(n10736), .B1(n10734), .B2(n11076), .ZN(
        P2_U3522) );
  INV_X1 U11446 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10735) );
  AOI22_X1 U11447 ( .A1(n11082), .A2(n10736), .B1(n10735), .B2(n11079), .ZN(
        P2_U3457) );
  INV_X1 U11448 ( .A(n10742), .ZN(n10745) );
  AOI21_X1 U11449 ( .B1(n10739), .B2(n10738), .A(n10737), .ZN(n10740) );
  OAI21_X1 U11450 ( .B1(n10742), .B2(n10741), .A(n10740), .ZN(n10743) );
  AOI211_X1 U11451 ( .C1(n10746), .C2(n10745), .A(n10744), .B(n10743), .ZN(
        n10748) );
  AOI22_X1 U11452 ( .A1(n11093), .A2(n10748), .B1(n7455), .B2(n11091), .ZN(
        P1_U3526) );
  INV_X1 U11453 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U11454 ( .A1(n11097), .A2(n10748), .B1(n10747), .B2(n11094), .ZN(
        P1_U3463) );
  INV_X1 U11455 ( .A(n10749), .ZN(n10753) );
  OAI22_X1 U11456 ( .A1(n10750), .A2(n11070), .B1(n8241), .B2(n11069), .ZN(
        n10752) );
  AOI211_X1 U11457 ( .C1(n10948), .C2(n10753), .A(n10752), .B(n10751), .ZN(
        n10756) );
  INV_X1 U11458 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U11459 ( .A1(n11078), .A2(n10756), .B1(n10754), .B2(n11076), .ZN(
        P2_U3523) );
  INV_X1 U11460 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U11461 ( .A1(n11082), .A2(n10756), .B1(n10755), .B2(n11079), .ZN(
        P2_U3460) );
  OAI21_X1 U11462 ( .B1(n10758), .B2(n11083), .A(n10757), .ZN(n10760) );
  AOI211_X1 U11463 ( .C1(n11016), .C2(n10761), .A(n10760), .B(n10759), .ZN(
        n10763) );
  AOI22_X1 U11464 ( .A1(n11093), .A2(n10763), .B1(n7460), .B2(n11091), .ZN(
        P1_U3527) );
  INV_X1 U11465 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U11466 ( .A1(n11097), .A2(n10763), .B1(n10762), .B2(n11094), .ZN(
        P1_U3466) );
  INV_X1 U11467 ( .A(n10764), .ZN(n10767) );
  INV_X1 U11468 ( .A(n10765), .ZN(n10766) );
  AOI21_X1 U11469 ( .B1(n10768), .B2(n10767), .A(n10766), .ZN(n10789) );
  OAI21_X1 U11470 ( .B1(n10770), .B2(n8331), .A(n10769), .ZN(n10771) );
  INV_X1 U11471 ( .A(n10771), .ZN(n10772) );
  OR2_X1 U11472 ( .A1(n10772), .A2(n10803), .ZN(n10783) );
  OAI22_X1 U11473 ( .A1(n10783), .A2(n11070), .B1(n8247), .B2(n11069), .ZN(
        n10778) );
  AOI21_X1 U11474 ( .B1(n10773), .B2(n8258), .A(n10811), .ZN(n10776) );
  AOI21_X1 U11475 ( .B1(n10776), .B2(n10775), .A(n10774), .ZN(n10792) );
  INV_X1 U11476 ( .A(n10792), .ZN(n10777) );
  AOI211_X1 U11477 ( .C1(n10789), .C2(n11074), .A(n10778), .B(n10777), .ZN(
        n10781) );
  INV_X1 U11478 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U11479 ( .A1(n11078), .A2(n10781), .B1(n10779), .B2(n11076), .ZN(
        P2_U3524) );
  INV_X1 U11480 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U11481 ( .A1(n11082), .A2(n10781), .B1(n10780), .B2(n11079), .ZN(
        P2_U3463) );
  INV_X1 U11482 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10782) );
  NOR2_X1 U11483 ( .A1(n10957), .A2(n10782), .ZN(n10785) );
  NOR2_X1 U11484 ( .A1(n10952), .A2(n10783), .ZN(n10784) );
  AOI211_X1 U11485 ( .C1(n10962), .C2(n10786), .A(n10785), .B(n10784), .ZN(
        n10787) );
  OAI21_X1 U11486 ( .B1(n8247), .B2(n10956), .A(n10787), .ZN(n10788) );
  AOI21_X1 U11487 ( .B1(n10790), .B2(n10789), .A(n10788), .ZN(n10791) );
  OAI21_X1 U11488 ( .B1(n10906), .B2(n10792), .A(n10791), .ZN(P2_U3292) );
  OAI21_X1 U11489 ( .B1(n10794), .B2(n11083), .A(n10793), .ZN(n10796) );
  AOI211_X1 U11490 ( .C1(n10797), .C2(n11089), .A(n10796), .B(n10795), .ZN(
        n10800) );
  AOI22_X1 U11491 ( .A1(n11093), .A2(n10800), .B1(n10798), .B2(n11091), .ZN(
        P1_U3528) );
  INV_X1 U11492 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U11493 ( .A1(n11097), .A2(n10800), .B1(n10799), .B2(n11094), .ZN(
        P1_U3469) );
  INV_X1 U11494 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10815) );
  XNOR2_X1 U11495 ( .A(n10801), .B(n10808), .ZN(n10820) );
  OAI211_X1 U11496 ( .C1(n10803), .C2(n10817), .A(n10802), .B(n10892), .ZN(
        n10816) );
  NAND2_X1 U11497 ( .A1(n10899), .A2(n10804), .ZN(n10807) );
  NAND2_X1 U11498 ( .A1(n10962), .A2(n10805), .ZN(n10806) );
  OAI211_X1 U11499 ( .C1(n10816), .C2(n10902), .A(n10807), .B(n10806), .ZN(
        n10813) );
  XNOR2_X1 U11500 ( .A(n10809), .B(n10808), .ZN(n10812) );
  OAI21_X1 U11501 ( .B1(n10812), .B2(n10811), .A(n10810), .ZN(n10818) );
  AOI211_X1 U11502 ( .C1(n10820), .C2(n10904), .A(n10813), .B(n10818), .ZN(
        n10814) );
  AOI22_X1 U11503 ( .A1(n10906), .A2(n10815), .B1(n10814), .B2(n10957), .ZN(
        P2_U3291) );
  OAI21_X1 U11504 ( .B1(n10817), .B2(n11069), .A(n10816), .ZN(n10819) );
  AOI211_X1 U11505 ( .C1(n10820), .C2(n11074), .A(n10819), .B(n10818), .ZN(
        n10823) );
  INV_X1 U11506 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U11507 ( .A1(n11078), .A2(n10823), .B1(n10821), .B2(n11076), .ZN(
        P2_U3525) );
  INV_X1 U11508 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U11509 ( .A1(n11082), .A2(n10823), .B1(n10822), .B2(n11079), .ZN(
        P2_U3466) );
  INV_X1 U11510 ( .A(n10824), .ZN(n10829) );
  OAI22_X1 U11511 ( .A1(n10826), .A2(n11085), .B1(n10825), .B2(n11083), .ZN(
        n10828) );
  AOI211_X1 U11512 ( .C1(n11016), .C2(n10829), .A(n10828), .B(n10827), .ZN(
        n10831) );
  AOI22_X1 U11513 ( .A1(n11093), .A2(n10831), .B1(n7454), .B2(n11091), .ZN(
        P1_U3529) );
  INV_X1 U11514 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U11515 ( .A1(n11097), .A2(n10831), .B1(n10830), .B2(n11094), .ZN(
        P1_U3472) );
  AOI22_X1 U11516 ( .A1(n10833), .A2(n10892), .B1(n10975), .B2(n10832), .ZN(
        n10836) );
  NAND3_X1 U11517 ( .A1(n9898), .A2(n10834), .A3(n11074), .ZN(n10835) );
  AND3_X1 U11518 ( .A1(n10837), .A2(n10836), .A3(n10835), .ZN(n10839) );
  AOI22_X1 U11519 ( .A1(n11078), .A2(n10839), .B1(n7280), .B2(n11076), .ZN(
        P2_U3526) );
  INV_X1 U11520 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U11521 ( .A1(n11082), .A2(n10839), .B1(n10838), .B2(n11079), .ZN(
        P2_U3469) );
  XNOR2_X1 U11522 ( .A(n10840), .B(n10848), .ZN(n10856) );
  INV_X1 U11523 ( .A(n10856), .ZN(n10862) );
  NOR2_X1 U11524 ( .A1(n10841), .A2(n10863), .ZN(n10842) );
  OR2_X1 U11525 ( .A1(n10843), .A2(n10842), .ZN(n10860) );
  OAI22_X1 U11526 ( .A1(n10860), .A2(n11085), .B1(n10863), .B2(n11083), .ZN(
        n10857) );
  AND2_X1 U11527 ( .A1(n10845), .A2(n10844), .ZN(n10847) );
  OAI21_X1 U11528 ( .B1(n10848), .B2(n10847), .A(n10846), .ZN(n10854) );
  OAI22_X1 U11529 ( .A1(n10852), .A2(n10851), .B1(n10850), .B2(n10849), .ZN(
        n10853) );
  AOI21_X1 U11530 ( .B1(n10854), .B2(n11009), .A(n10853), .ZN(n10855) );
  OAI21_X1 U11531 ( .B1(n10856), .B2(n11013), .A(n10855), .ZN(n10870) );
  AOI211_X1 U11532 ( .C1(n11016), .C2(n10862), .A(n10857), .B(n10870), .ZN(
        n10859) );
  AOI22_X1 U11533 ( .A1(n11093), .A2(n10859), .B1(n7465), .B2(n11091), .ZN(
        P1_U3530) );
  INV_X1 U11534 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U11535 ( .A1(n11097), .A2(n10859), .B1(n10858), .B2(n11094), .ZN(
        P1_U3475) );
  INV_X1 U11536 ( .A(n10860), .ZN(n10861) );
  AOI22_X1 U11537 ( .A1(n10862), .A2(n11023), .B1(n11022), .B2(n10861), .ZN(
        n10872) );
  NOR2_X1 U11538 ( .A1(n11029), .A2(n10863), .ZN(n10868) );
  INV_X1 U11539 ( .A(n10864), .ZN(n10866) );
  OAI22_X1 U11540 ( .A1(n10869), .A2(n7486), .B1(n10866), .B2(n10865), .ZN(
        n10867) );
  AOI211_X1 U11541 ( .C1(n10870), .C2(n10869), .A(n10868), .B(n10867), .ZN(
        n10871) );
  NAND2_X1 U11542 ( .A1(n10872), .A2(n10871), .ZN(P1_U3284) );
  AOI22_X1 U11543 ( .A1(n10874), .A2(n10892), .B1(n10975), .B2(n10873), .ZN(
        n10875) );
  OAI211_X1 U11544 ( .C1(n10877), .C2(n11034), .A(n10876), .B(n10875), .ZN(
        n10878) );
  INV_X1 U11545 ( .A(n10878), .ZN(n10881) );
  INV_X1 U11546 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U11547 ( .A1(n11078), .A2(n10881), .B1(n10879), .B2(n11076), .ZN(
        P2_U3527) );
  INV_X1 U11548 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U11549 ( .A1(n11082), .A2(n10881), .B1(n10880), .B2(n11079), .ZN(
        P2_U3472) );
  OAI22_X1 U11550 ( .A1(n10883), .A2(n11085), .B1(n10882), .B2(n11083), .ZN(
        n10885) );
  AOI211_X1 U11551 ( .C1(n11016), .C2(n10886), .A(n10885), .B(n10884), .ZN(
        n10889) );
  AOI22_X1 U11552 ( .A1(n11093), .A2(n10889), .B1(n10887), .B2(n11091), .ZN(
        P1_U3531) );
  INV_X1 U11553 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U11554 ( .A1(n11097), .A2(n10889), .B1(n10888), .B2(n11094), .ZN(
        P1_U3478) );
  XNOR2_X1 U11555 ( .A(n10890), .B(n5225), .ZN(n10911) );
  XNOR2_X1 U11556 ( .A(n10891), .B(n10898), .ZN(n10893) );
  NAND2_X1 U11557 ( .A1(n10893), .A2(n10892), .ZN(n10907) );
  XNOR2_X1 U11558 ( .A(n10894), .B(n10895), .ZN(n10897) );
  AOI21_X1 U11559 ( .B1(n10897), .B2(n10942), .A(n10896), .ZN(n10908) );
  AOI22_X1 U11560 ( .A1(n10962), .A2(n10900), .B1(n10899), .B2(n10898), .ZN(
        n10901) );
  OAI211_X1 U11561 ( .C1(n10902), .C2(n10907), .A(n10908), .B(n10901), .ZN(
        n10903) );
  AOI21_X1 U11562 ( .B1(n10904), .B2(n10911), .A(n10903), .ZN(n10905) );
  AOI22_X1 U11563 ( .A1(n10906), .A2(n7321), .B1(n10905), .B2(n10957), .ZN(
        P2_U3288) );
  OAI211_X1 U11564 ( .C1(n10909), .C2(n11069), .A(n10908), .B(n10907), .ZN(
        n10910) );
  AOI21_X1 U11565 ( .B1(n11074), .B2(n10911), .A(n10910), .ZN(n10913) );
  AOI22_X1 U11566 ( .A1(n11078), .A2(n10913), .B1(n7316), .B2(n11076), .ZN(
        P2_U3528) );
  INV_X1 U11567 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U11568 ( .A1(n11082), .A2(n10913), .B1(n10912), .B2(n11079), .ZN(
        P2_U3475) );
  OAI22_X1 U11569 ( .A1(n10915), .A2(n11085), .B1(n10914), .B2(n11083), .ZN(
        n10917) );
  AOI211_X1 U11570 ( .C1(n11089), .C2(n10918), .A(n10917), .B(n10916), .ZN(
        n10920) );
  AOI22_X1 U11571 ( .A1(n11093), .A2(n10920), .B1(n7467), .B2(n11091), .ZN(
        P1_U3532) );
  INV_X1 U11572 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U11573 ( .A1(n11097), .A2(n10920), .B1(n10919), .B2(n11094), .ZN(
        P1_U3481) );
  INV_X1 U11574 ( .A(n10921), .ZN(n10926) );
  OAI22_X1 U11575 ( .A1(n10923), .A2(n11070), .B1(n10922), .B2(n11069), .ZN(
        n10925) );
  AOI211_X1 U11576 ( .C1(n10948), .C2(n10926), .A(n10925), .B(n10924), .ZN(
        n10928) );
  AOI22_X1 U11577 ( .A1(n11078), .A2(n10928), .B1(n7366), .B2(n11076), .ZN(
        P2_U3529) );
  INV_X1 U11578 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U11579 ( .A1(n11082), .A2(n10928), .B1(n10927), .B2(n11079), .ZN(
        P2_U3478) );
  OAI21_X1 U11580 ( .B1(n10929), .B2(n10931), .A(n10930), .ZN(n10954) );
  INV_X1 U11581 ( .A(n10954), .ZN(n10947) );
  NAND2_X1 U11582 ( .A1(n10933), .A2(n10932), .ZN(n10934) );
  NAND2_X1 U11583 ( .A1(n5122), .A2(n10934), .ZN(n10951) );
  OAI22_X1 U11584 ( .A1(n10951), .A2(n11070), .B1(n5353), .B2(n11069), .ZN(
        n10946) );
  OAI21_X1 U11585 ( .B1(n5124), .B2(n10936), .A(n10935), .ZN(n10943) );
  OAI22_X1 U11586 ( .A1(n10940), .A2(n10939), .B1(n10938), .B2(n10937), .ZN(
        n10941) );
  AOI21_X1 U11587 ( .B1(n10943), .B2(n10942), .A(n10941), .ZN(n10944) );
  OAI21_X1 U11588 ( .B1(n10954), .B2(n10945), .A(n10944), .ZN(n10958) );
  AOI211_X1 U11589 ( .C1(n10948), .C2(n10947), .A(n10946), .B(n10958), .ZN(
        n10950) );
  AOI22_X1 U11590 ( .A1(n11078), .A2(n10950), .B1(n7390), .B2(n11076), .ZN(
        P2_U3530) );
  INV_X1 U11591 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U11592 ( .A1(n11082), .A2(n10950), .B1(n10949), .B2(n11079), .ZN(
        P2_U3481) );
  OAI22_X1 U11593 ( .A1(n10954), .A2(n10953), .B1(n10952), .B2(n10951), .ZN(
        n10955) );
  INV_X1 U11594 ( .A(n10955), .ZN(n10964) );
  NOR2_X1 U11595 ( .A1(n10956), .A2(n5353), .ZN(n10960) );
  MUX2_X1 U11596 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10958), .S(n10957), .Z(
        n10959) );
  AOI211_X1 U11597 ( .C1(n10962), .C2(n10961), .A(n10960), .B(n10959), .ZN(
        n10963) );
  NAND2_X1 U11598 ( .A1(n10964), .A2(n10963), .ZN(P2_U3286) );
  OAI22_X1 U11599 ( .A1(n10966), .A2(n11085), .B1(n10965), .B2(n11083), .ZN(
        n10968) );
  AOI211_X1 U11600 ( .C1(n11016), .C2(n10969), .A(n10968), .B(n10967), .ZN(
        n10972) );
  AOI22_X1 U11601 ( .A1(n11093), .A2(n10972), .B1(n10970), .B2(n11091), .ZN(
        P1_U3534) );
  INV_X1 U11602 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U11603 ( .A1(n11097), .A2(n10972), .B1(n10971), .B2(n11094), .ZN(
        P1_U3487) );
  AOI21_X1 U11604 ( .B1(n10975), .B2(n10974), .A(n10973), .ZN(n10976) );
  OAI211_X1 U11605 ( .C1(n10978), .C2(n11034), .A(n10977), .B(n10976), .ZN(
        n10979) );
  INV_X1 U11606 ( .A(n10979), .ZN(n10981) );
  AOI22_X1 U11607 ( .A1(n11078), .A2(n10981), .B1(n7868), .B2(n11076), .ZN(
        P2_U3531) );
  INV_X1 U11608 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U11609 ( .A1(n11082), .A2(n10981), .B1(n10980), .B2(n11079), .ZN(
        P2_U3484) );
  OAI22_X1 U11610 ( .A1(n10983), .A2(n11085), .B1(n10982), .B2(n11083), .ZN(
        n10985) );
  AOI211_X1 U11611 ( .C1(n11016), .C2(n10986), .A(n10985), .B(n10984), .ZN(
        n10989) );
  AOI22_X1 U11612 ( .A1(n11093), .A2(n10989), .B1(n10987), .B2(n11091), .ZN(
        P1_U3535) );
  INV_X1 U11613 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U11614 ( .A1(n11097), .A2(n10989), .B1(n10988), .B2(n11094), .ZN(
        P1_U3490) );
  OAI22_X1 U11615 ( .A1(n10991), .A2(n11070), .B1(n10990), .B2(n11069), .ZN(
        n10993) );
  AOI211_X1 U11616 ( .C1(n11074), .C2(n10994), .A(n10993), .B(n10992), .ZN(
        n10996) );
  AOI22_X1 U11617 ( .A1(n11078), .A2(n10996), .B1(n7981), .B2(n11076), .ZN(
        P2_U3532) );
  INV_X1 U11618 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U11619 ( .A1(n11082), .A2(n10996), .B1(n10995), .B2(n11079), .ZN(
        P2_U3487) );
  INV_X1 U11620 ( .A(n10997), .ZN(n10998) );
  AOI21_X1 U11621 ( .B1(n11007), .B2(n10999), .A(n10998), .ZN(n11014) );
  INV_X1 U11622 ( .A(n11014), .ZN(n11024) );
  INV_X1 U11623 ( .A(n11000), .ZN(n11002) );
  OAI21_X1 U11624 ( .B1(n11002), .B2(n5339), .A(n11001), .ZN(n11020) );
  OAI22_X1 U11625 ( .A1(n11020), .A2(n11085), .B1(n5339), .B2(n11083), .ZN(
        n11015) );
  AOI22_X1 U11626 ( .A1(n11006), .A2(n11005), .B1(n11004), .B2(n11003), .ZN(
        n11012) );
  XNOR2_X1 U11627 ( .A(n11008), .B(n11007), .ZN(n11010) );
  NAND2_X1 U11628 ( .A1(n11010), .A2(n11009), .ZN(n11011) );
  OAI211_X1 U11629 ( .C1(n11014), .C2(n11013), .A(n11012), .B(n11011), .ZN(
        n11031) );
  AOI211_X1 U11630 ( .C1(n11016), .C2(n11024), .A(n11015), .B(n11031), .ZN(
        n11019) );
  AOI22_X1 U11631 ( .A1(n11093), .A2(n11019), .B1(n11017), .B2(n11091), .ZN(
        P1_U3536) );
  INV_X1 U11632 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U11633 ( .A1(n11097), .A2(n11019), .B1(n11018), .B2(n11094), .ZN(
        P1_U3493) );
  INV_X1 U11634 ( .A(n11020), .ZN(n11021) );
  AOI22_X1 U11635 ( .A1(n11024), .A2(n11023), .B1(n11022), .B2(n11021), .ZN(
        n11033) );
  AOI22_X1 U11636 ( .A1(n11027), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n11026), 
        .B2(n11025), .ZN(n11028) );
  OAI21_X1 U11637 ( .B1(n5339), .B2(n11029), .A(n11028), .ZN(n11030) );
  AOI21_X1 U11638 ( .B1(n11031), .B2(n10869), .A(n11030), .ZN(n11032) );
  NAND2_X1 U11639 ( .A1(n11033), .A2(n11032), .ZN(P1_U3278) );
  NOR2_X1 U11640 ( .A1(n11035), .A2(n11034), .ZN(n11041) );
  OAI22_X1 U11641 ( .A1(n11037), .A2(n11070), .B1(n11036), .B2(n11069), .ZN(
        n11039) );
  AOI211_X1 U11642 ( .C1(n11041), .C2(n11040), .A(n11039), .B(n11038), .ZN(
        n11043) );
  AOI22_X1 U11643 ( .A1(n11078), .A2(n11043), .B1(n7980), .B2(n11076), .ZN(
        P2_U3533) );
  INV_X1 U11644 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U11645 ( .A1(n11082), .A2(n11043), .B1(n11042), .B2(n11079), .ZN(
        P2_U3490) );
  OAI22_X1 U11646 ( .A1(n11044), .A2(n11085), .B1(n5338), .B2(n11083), .ZN(
        n11046) );
  AOI211_X1 U11647 ( .C1(n11089), .C2(n11047), .A(n11046), .B(n11045), .ZN(
        n11049) );
  AOI22_X1 U11648 ( .A1(n11093), .A2(n11049), .B1(n7885), .B2(n11091), .ZN(
        P1_U3537) );
  INV_X1 U11649 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U11650 ( .A1(n11097), .A2(n11049), .B1(n11048), .B2(n11094), .ZN(
        P1_U3496) );
  INV_X1 U11651 ( .A(n11050), .ZN(n11056) );
  INV_X1 U11652 ( .A(n11051), .ZN(n11052) );
  OAI22_X1 U11653 ( .A1(n11053), .A2(n11070), .B1(n11052), .B2(n11069), .ZN(
        n11054) );
  AOI211_X1 U11654 ( .C1(n11056), .C2(n11074), .A(n11055), .B(n11054), .ZN(
        n11058) );
  AOI22_X1 U11655 ( .A1(n11078), .A2(n11058), .B1(n8103), .B2(n11076), .ZN(
        P2_U3534) );
  INV_X1 U11656 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U11657 ( .A1(n11082), .A2(n11058), .B1(n11057), .B2(n11079), .ZN(
        P2_U3493) );
  NOR2_X1 U11658 ( .A1(n11060), .A2(n11059), .ZN(n11066) );
  OAI22_X1 U11659 ( .A1(n11062), .A2(n11085), .B1(n11061), .B2(n11083), .ZN(
        n11064) );
  AOI211_X1 U11660 ( .C1(n11066), .C2(n11065), .A(n11064), .B(n11063), .ZN(
        n11068) );
  AOI22_X1 U11661 ( .A1(n11093), .A2(n11068), .B1(n8054), .B2(n11091), .ZN(
        P1_U3538) );
  INV_X1 U11662 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11067) );
  AOI22_X1 U11663 ( .A1(n11097), .A2(n11068), .B1(n11067), .B2(n11094), .ZN(
        P1_U3499) );
  OAI22_X1 U11664 ( .A1(n11071), .A2(n11070), .B1(n5215), .B2(n11069), .ZN(
        n11072) );
  AOI211_X1 U11665 ( .C1(n11075), .C2(n11074), .A(n11073), .B(n11072), .ZN(
        n11081) );
  AOI22_X1 U11666 ( .A1(n11078), .A2(n11081), .B1(n11077), .B2(n11076), .ZN(
        P2_U3535) );
  INV_X1 U11667 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U11668 ( .A1(n11082), .A2(n11081), .B1(n11080), .B2(n11079), .ZN(
        P2_U3496) );
  OAI22_X1 U11669 ( .A1(n11086), .A2(n11085), .B1(n11084), .B2(n11083), .ZN(
        n11088) );
  AOI211_X1 U11670 ( .C1(n11090), .C2(n11089), .A(n11088), .B(n11087), .ZN(
        n11096) );
  AOI22_X1 U11671 ( .A1(n11093), .A2(n11096), .B1(n11092), .B2(n11091), .ZN(
        P1_U3539) );
  INV_X1 U11672 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n11095) );
  AOI22_X1 U11673 ( .A1(n11097), .A2(n11096), .B1(n11095), .B2(n11094), .ZN(
        P1_U3502) );
  XNOR2_X1 U11674 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U5110 ( .A(n6373), .ZN(n6341) );
  CLKBUF_X1 U5113 ( .A(n5175), .Z(n5037) );
  CLKBUF_X1 U5126 ( .A(n5060), .Z(n6885) );
  AOI21_X1 U5133 ( .B1(n10683), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10678), .ZN(
        n7347) );
  CLKBUF_X1 U5135 ( .A(n6416), .Z(n5036) );
endmodule

