

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6428, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617;

  AOI211_X1 U7175 ( .C1(n15311), .C2(n15036), .A(n15035), .B(n15034), .ZN(
        n15038) );
  INV_X4 U7176 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X4 U7178 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OR2_X1 U7179 ( .A1(n8292), .A2(n8291), .ZN(n8306) );
  INV_X2 U7181 ( .A(n12728), .ZN(n6436) );
  NAND2_X1 U7182 ( .A1(n7906), .A2(n7905), .ZN(n11596) );
  OR2_X1 U7183 ( .A1(n15532), .A2(n11163), .ZN(n12408) );
  CLKBUF_X2 U7185 ( .A(n9015), .Z(n12367) );
  INV_X1 U7186 ( .A(n8471), .ZN(n8702) );
  INV_X2 U7187 ( .A(n12365), .ZN(n9813) );
  INV_X1 U7188 ( .A(n12394), .ZN(n12392) );
  INV_X1 U7189 ( .A(n7856), .ZN(n8166) );
  CLKBUF_X2 U7190 ( .A(n12376), .Z(n6435) );
  NAND2_X1 U7191 ( .A1(n8933), .A2(n8929), .ZN(n9425) );
  AND2_X4 U7192 ( .A1(n7778), .A2(n15160), .ZN(n7835) );
  XNOR2_X1 U7193 ( .A(n8432), .B(n8431), .ZN(n10417) );
  NAND2_X1 U7194 ( .A1(n6777), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7794) );
  CLKBUF_X1 U7195 ( .A(n13563), .Z(n6428) );
  NOR2_X1 U7196 ( .A1(n11782), .A2(n15541), .ZN(n13563) );
  AND2_X1 U7197 ( .A1(n13925), .A2(n7584), .ZN(n7581) );
  INV_X2 U7198 ( .A(n14414), .ZN(n14346) );
  NAND2_X1 U7199 ( .A1(n10383), .A2(n10380), .ZN(n10527) );
  OAI22_X1 U7200 ( .A1(n7278), .A2(n9624), .B1(n11413), .B2(n7276), .ZN(n9553)
         );
  AND2_X1 U7201 ( .A1(n9470), .A2(n12390), .ZN(n12391) );
  INV_X1 U7202 ( .A(n9726), .ZN(n9777) );
  AND2_X1 U7203 ( .A1(n7259), .A2(n7258), .ZN(n12978) );
  NAND2_X1 U7204 ( .A1(n11345), .A2(n11582), .ZN(n11697) );
  INV_X2 U7205 ( .A(n14359), .ZN(n11660) );
  AND2_X1 U7206 ( .A1(n9060), .A2(n10944), .ZN(n9077) );
  INV_X1 U7207 ( .A(n9425), .ZN(n9325) );
  NAND2_X1 U7208 ( .A1(n11414), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11413) );
  INV_X1 U7209 ( .A(n12543), .ZN(n13389) );
  NAND2_X1 U7210 ( .A1(n13577), .A2(n13428), .ZN(n12506) );
  AND2_X2 U7211 ( .A1(n8827), .A2(n11070), .ZN(n11176) );
  INV_X1 U7212 ( .A(n12692), .ZN(n15491) );
  INV_X1 U7213 ( .A(n14578), .ZN(n12041) );
  INV_X1 U7214 ( .A(n14576), .ZN(n14521) );
  NOR2_X2 U7215 ( .A1(n7740), .A2(n15117), .ZN(n12072) );
  INV_X1 U7216 ( .A(n7868), .ZN(n8167) );
  AND4_X1 U7217 ( .A1(n9405), .A2(n9404), .A3(n9403), .A4(n9402), .ZN(n13048)
         );
  NAND2_X1 U7218 ( .A1(n13511), .A2(n6675), .ZN(n13499) );
  AND2_X1 U7219 ( .A1(n9412), .A2(n6505), .ZN(n12582) );
  INV_X1 U7220 ( .A(n8440), .ZN(n12820) );
  AND4_X1 U7221 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), .ZN(n11316)
         );
  INV_X1 U7222 ( .A(n15437), .ZN(n14085) );
  NAND2_X1 U7223 ( .A1(n8825), .A2(n8824), .ZN(n14222) );
  AND4_X1 U7224 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7876), .ZN(n11284)
         );
  CLKBUF_X1 U7225 ( .A(n11032), .Z(n6434) );
  NAND2_X1 U7226 ( .A1(n8205), .A2(n8204), .ZN(n14888) );
  AOI211_X1 U7227 ( .C1(n13581), .C2(n13435), .A(n13434), .B(n13433), .ZN(
        n13584) );
  NAND2_X1 U7228 ( .A1(n13007), .A2(n6992), .ZN(n13016) );
  INV_X2 U7229 ( .A(n14064), .ZN(n6438) );
  AOI211_X1 U7230 ( .C1(n15273), .C2(n14774), .A(n14773), .B(n14772), .ZN(
        n14775) );
  NAND2_X1 U7231 ( .A1(n7360), .A2(n7361), .ZN(n11076) );
  AOI21_X2 U7232 ( .B1(n7243), .B2(n9030), .A(n10939), .ZN(n7239) );
  NAND2_X2 U7233 ( .A1(n7505), .A2(n11408), .ZN(n10048) );
  NAND4_X4 U7234 ( .A1(n8452), .A2(n8455), .A3(n8454), .A4(n8453), .ZN(n13866)
         );
  XNOR2_X1 U7235 ( .A(n6973), .B(n10088), .ZN(n9859) );
  BUF_X2 U7237 ( .A(n15310), .Z(n6430) );
  OAI211_X1 U7238 ( .C1(n7856), .C2(n14619), .A(n7870), .B(n7869), .ZN(n15310)
         );
  NAND2_X1 U7239 ( .A1(n7360), .A2(n7361), .ZN(n6431) );
  OAI21_X1 U7240 ( .B1(n7294), .B2(n10403), .A(n7293), .ZN(n13251) );
  NOR2_X4 U7241 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8467) );
  BUF_X2 U7242 ( .A(n8447), .Z(n8497) );
  AND2_X2 U7243 ( .A1(n9893), .A2(n8316), .ZN(n10517) );
  NOR2_X2 U7244 ( .A1(n9136), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9154) );
  OAI21_X2 U7245 ( .B1(n13770), .B2(n13766), .A(n13767), .ZN(n13733) );
  AOI21_X2 U7246 ( .B1(n7843), .B2(n7842), .A(n7841), .ZN(n7865) );
  NAND2_X2 U7247 ( .A1(n8395), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7502) );
  AND2_X1 U7248 ( .A1(n10371), .A2(n15297), .ZN(n14962) );
  NOR2_X2 U7249 ( .A1(n6690), .A2(n6687), .ZN(n9407) );
  AOI21_X2 U7250 ( .B1(n13232), .B2(n13230), .A(n13231), .ZN(n13234) );
  BUF_X1 U7251 ( .A(n11032), .Z(n6433) );
  OAI211_X1 U7252 ( .C1(n8262), .C2(n10276), .A(n7849), .B(n7848), .ZN(n11032)
         );
  NAND2_X2 U7253 ( .A1(n8354), .A2(n8353), .ZN(n14784) );
  XNOR2_X2 U7254 ( .A(n14115), .B(n13839), .ZN(n13925) );
  NAND2_X1 U7255 ( .A1(n8939), .A2(n10039), .ZN(n12376) );
  XNOR2_X2 U7256 ( .A(n7758), .B(P1_IR_REG_19__SCAN_IN), .ZN(n15296) );
  AOI21_X2 U7257 ( .B1(n11055), .B2(n8522), .A(n7736), .ZN(n11237) );
  NAND2_X2 U7258 ( .A1(n15439), .A2(n15440), .ZN(n11055) );
  NAND2_X2 U7259 ( .A1(n8510), .A2(n8511), .ZN(n12933) );
  INV_X2 U7260 ( .A(n14351), .ZN(n14413) );
  AND2_X1 U7261 ( .A1(n14750), .A2(n15027), .ZN(n12656) );
  NAND2_X1 U7262 ( .A1(n6975), .A2(n7433), .ZN(n6442) );
  AND2_X1 U7263 ( .A1(n9841), .A2(n9840), .ZN(n14768) );
  OR2_X1 U7264 ( .A1(n9425), .A2(n13371), .ZN(n9391) );
  AND2_X1 U7265 ( .A1(n8153), .A2(n8152), .ZN(n15144) );
  AND2_X1 U7266 ( .A1(n9551), .A2(n9623), .ZN(n6920) );
  AND2_X1 U7267 ( .A1(n6733), .A2(n11116), .ZN(n11218) );
  OR2_X1 U7268 ( .A1(n13420), .A2(n9425), .ZN(n9344) );
  NAND2_X1 U7269 ( .A1(n12407), .A2(n12402), .ZN(n15528) );
  INV_X4 U7270 ( .A(n14413), .ZN(n14295) );
  NAND2_X1 U7271 ( .A1(n12408), .A2(n12409), .ZN(n12548) );
  INV_X4 U7272 ( .A(n12524), .ZN(n12529) );
  NAND2_X1 U7273 ( .A1(n6660), .A2(n6661), .ZN(n15533) );
  NOR2_X4 U7274 ( .A1(n14414), .A2(n14962), .ZN(n10794) );
  INV_X1 U7275 ( .A(n13866), .ZN(n8458) );
  NAND4_X1 U7276 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n13213)
         );
  OR2_X2 U7277 ( .A1(n7768), .A2(n10380), .ZN(n14359) );
  CLKBUF_X2 U7278 ( .A(n9024), .Z(n9259) );
  INV_X2 U7279 ( .A(n12366), .ZN(n9093) );
  INV_X2 U7280 ( .A(n8262), .ZN(n10061) );
  NAND4_X1 U7281 ( .A1(n8464), .A2(n8463), .A3(n8462), .A4(n8461), .ZN(n13865)
         );
  NAND2_X1 U7282 ( .A1(n15297), .A2(n10092), .ZN(n10379) );
  INV_X2 U7283 ( .A(n12906), .ZN(n6437) );
  OAI21_X1 U7284 ( .B1(n6439), .B2(n7902), .A(n7901), .ZN(n7935) );
  OAI21_X1 U7285 ( .B1(n6439), .B2(n7867), .A(n7866), .ZN(n7897) );
  INV_X4 U7286 ( .A(n10193), .ZN(n10039) );
  AND2_X2 U7287 ( .A1(n9055), .A2(n6523), .ZN(n9112) );
  NAND2_X1 U7288 ( .A1(n6670), .A2(n6672), .ZN(n13399) );
  NAND2_X1 U7289 ( .A1(n9859), .A2(n14874), .ZN(n15037) );
  AOI21_X1 U7290 ( .B1(n12535), .B2(n12536), .A(n12534), .ZN(n12539) );
  OR2_X1 U7291 ( .A1(n13730), .A2(n6996), .ZN(n6995) );
  INV_X1 U7292 ( .A(n12978), .ZN(n13808) );
  AND2_X1 U7293 ( .A1(n15045), .A2(n6843), .ZN(n6842) );
  XNOR2_X1 U7294 ( .A(n9487), .B(n12568), .ZN(n9527) );
  NOR2_X1 U7295 ( .A1(n6552), .A2(n6709), .ZN(n6708) );
  AND2_X1 U7296 ( .A1(n14373), .A2(n14372), .ZN(n14417) );
  AND3_X1 U7297 ( .A1(n9824), .A2(n9823), .A3(n9822), .ZN(n13629) );
  OAI21_X1 U7298 ( .B1(n7318), .B2(n13179), .A(n13080), .ZN(n6911) );
  AND2_X1 U7299 ( .A1(n13427), .A2(n13426), .ZN(n13581) );
  NAND2_X1 U7300 ( .A1(n10143), .A2(n12542), .ZN(n10142) );
  OR2_X1 U7301 ( .A1(n9821), .A2(n6613), .ZN(n9822) );
  NAND2_X1 U7302 ( .A1(n6926), .A2(n7677), .ZN(n14109) );
  AND2_X1 U7303 ( .A1(n7321), .A2(n6592), .ZN(n7319) );
  OAI21_X1 U7304 ( .B1(n14450), .B2(n7616), .A(n6729), .ZN(n14538) );
  NAND2_X1 U7305 ( .A1(n8314), .A2(n8313), .ZN(n9878) );
  NAND2_X1 U7306 ( .A1(n10144), .A2(n9394), .ZN(n10146) );
  MUX2_X1 U7307 ( .A(n12654), .B(n12656), .S(n15319), .Z(n12655) );
  NAND2_X1 U7308 ( .A1(n6442), .A2(n8346), .ZN(n14838) );
  NAND2_X1 U7309 ( .A1(n9347), .A2(n13407), .ZN(n13415) );
  INV_X1 U7310 ( .A(n6971), .ZN(n6970) );
  NAND2_X1 U7311 ( .A1(n14424), .A2(n14425), .ZN(n6709) );
  NAND2_X1 U7312 ( .A1(n14813), .A2(n14812), .ZN(n14811) );
  NOR2_X1 U7313 ( .A1(n6960), .A2(n6956), .ZN(n6955) );
  AND3_X1 U7314 ( .A1(n7583), .A2(n7582), .A3(n7590), .ZN(n12958) );
  AOI21_X1 U7315 ( .B1(n7329), .B2(n7328), .A(n6532), .ZN(n7327) );
  NAND2_X1 U7316 ( .A1(n13984), .A2(n13986), .ZN(n13985) );
  NOR2_X1 U7317 ( .A1(n13251), .A2(n13561), .ZN(n13273) );
  OR2_X1 U7318 ( .A1(n14114), .A2(n6961), .ZN(n6960) );
  OAI21_X1 U7319 ( .B1(n14405), .B2(n7624), .A(n6726), .ZN(n14393) );
  AND2_X1 U7320 ( .A1(n9486), .A2(n12517), .ZN(n7175) );
  AOI21_X1 U7321 ( .B1(n7623), .B2(n6547), .A(n6727), .ZN(n6726) );
  NAND2_X1 U7322 ( .A1(n7294), .A2(n10403), .ZN(n7293) );
  AND2_X1 U7323 ( .A1(n13382), .A2(n13378), .ZN(n7176) );
  INV_X1 U7324 ( .A(n9838), .ZN(n6969) );
  NAND2_X1 U7325 ( .A1(n9399), .A2(n9398), .ZN(n13079) );
  XNOR2_X1 U7326 ( .A(n15036), .B(n10028), .ZN(n10088) );
  INV_X1 U7327 ( .A(n12512), .ZN(n13382) );
  NAND2_X1 U7328 ( .A1(n12252), .A2(n12251), .ZN(n13024) );
  NAND2_X1 U7329 ( .A1(n6751), .A2(n8697), .ZN(n14032) );
  NAND2_X1 U7330 ( .A1(n14528), .A2(n14529), .ZN(n14527) );
  OR2_X1 U7331 ( .A1(n13572), .A2(n13045), .ZN(n12517) );
  AND2_X1 U7332 ( .A1(n13403), .A2(n13416), .ZN(n12512) );
  AND2_X1 U7333 ( .A1(n8312), .A2(n8311), .ZN(n14543) );
  AND2_X1 U7334 ( .A1(n9865), .A2(n8362), .ZN(n14766) );
  AND2_X1 U7335 ( .A1(n7577), .A2(n13963), .ZN(n6460) );
  NOR2_X1 U7336 ( .A1(n14427), .A2(n7627), .ZN(n7626) );
  NAND2_X1 U7337 ( .A1(n6654), .A2(n9208), .ZN(n13514) );
  OAI21_X1 U7338 ( .B1(n13261), .B2(n7081), .A(n7079), .ZN(n9631) );
  AND2_X1 U7339 ( .A1(n7434), .A2(n8345), .ZN(n7433) );
  XNOR2_X1 U7340 ( .A(n6874), .B(n9383), .ZN(n13711) );
  NAND2_X1 U7341 ( .A1(n12812), .A2(n12811), .ZN(n12952) );
  AND2_X1 U7342 ( .A1(n7181), .A2(n12494), .ZN(n7180) );
  NAND2_X1 U7343 ( .A1(n9382), .A2(n9381), .ZN(n6874) );
  NAND2_X1 U7344 ( .A1(n7410), .A2(n7409), .ZN(n7408) );
  AOI21_X1 U7345 ( .B1(n14244), .B2(n10061), .A(n6616), .ZN(n12659) );
  OR2_X1 U7346 ( .A1(n9380), .A2(n9379), .ZN(n9382) );
  NAND2_X1 U7347 ( .A1(n8783), .A2(n8782), .ZN(n14115) );
  INV_X1 U7348 ( .A(n7411), .ZN(n7410) );
  OR2_X1 U7349 ( .A1(n7436), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U7350 ( .A1(n9338), .A2(n9337), .ZN(n13577) );
  NAND2_X1 U7351 ( .A1(n14316), .A2(n14315), .ZN(n14502) );
  NAND2_X1 U7352 ( .A1(n6440), .A2(n8330), .ZN(n11833) );
  INV_X1 U7353 ( .A(n13945), .ZN(n14119) );
  OR2_X1 U7354 ( .A1(n9425), .A2(n9505), .ZN(n9403) );
  AOI21_X1 U7355 ( .B1(n9351), .B2(n6482), .A(n6643), .ZN(n7532) );
  NAND2_X1 U7356 ( .A1(n8264), .A2(n8263), .ZN(n14833) );
  AND2_X1 U7357 ( .A1(n14873), .A2(n8341), .ZN(n14911) );
  OAI21_X1 U7358 ( .B1(n8794), .B2(n13712), .A(n8795), .ZN(n7140) );
  XNOR2_X1 U7359 ( .A(n8794), .B(SI_27_), .ZN(n15162) );
  AND2_X1 U7360 ( .A1(n8437), .A2(n8436), .ZN(n13945) );
  INV_X1 U7361 ( .A(n13385), .ZN(n13416) );
  INV_X1 U7362 ( .A(n11555), .ZN(n9688) );
  NAND2_X1 U7363 ( .A1(n8239), .A2(n8238), .ZN(n15061) );
  NAND2_X1 U7364 ( .A1(n6593), .A2(n11460), .ZN(n6441) );
  XNOR2_X1 U7365 ( .A(n9849), .B(n9843), .ZN(n8794) );
  AOI21_X1 U7366 ( .B1(n6940), .B2(n6534), .A(n6938), .ZN(n6937) );
  OAI21_X1 U7367 ( .B1(n11306), .B2(n11307), .A(n7282), .ZN(n7279) );
  OR2_X1 U7368 ( .A1(n9425), .A2(n13394), .ZN(n9374) );
  NAND2_X1 U7369 ( .A1(n8747), .A2(n8746), .ZN(n14138) );
  NAND4_X1 U7370 ( .A1(n9362), .A2(n9361), .A3(n9360), .A4(n9359), .ZN(n13385)
         );
  NAND2_X1 U7371 ( .A1(n6719), .A2(n6718), .ZN(n11476) );
  OR2_X1 U7372 ( .A1(n9425), .A2(n13400), .ZN(n9360) );
  CLKBUF_X1 U7373 ( .A(n11743), .Z(n6925) );
  OAI22_X2 U7374 ( .A1(n8302), .A2(n6769), .B1(n8300), .B2(n13718), .ZN(n9849)
         );
  NAND2_X1 U7375 ( .A1(n8724), .A2(n8723), .ZN(n14151) );
  NAND2_X1 U7376 ( .A1(n8738), .A2(n8737), .ZN(n14147) );
  NAND2_X1 U7377 ( .A1(n8704), .A2(n8703), .ZN(n14163) );
  NAND2_X1 U7378 ( .A1(n6443), .A2(n11279), .ZN(n11283) );
  NAND2_X1 U7379 ( .A1(n11560), .A2(n8568), .ZN(n11696) );
  XNOR2_X1 U7380 ( .A(n8237), .B(n8236), .ZN(n11733) );
  AND2_X1 U7381 ( .A1(n13022), .A2(n13559), .ZN(n7382) );
  AOI21_X1 U7382 ( .B1(n6988), .B2(n6990), .A(n6987), .ZN(n6986) );
  NAND2_X1 U7383 ( .A1(n8211), .A2(n8210), .ZN(n14910) );
  NAND2_X1 U7384 ( .A1(n8169), .A2(n8168), .ZN(n15088) );
  NAND2_X1 U7385 ( .A1(n11092), .A2(n11280), .ZN(n6443) );
  NAND2_X1 U7386 ( .A1(n7493), .A2(n8272), .ZN(n8287) );
  NAND2_X1 U7387 ( .A1(n8257), .A2(n8258), .ZN(n7493) );
  NAND2_X1 U7388 ( .A1(n8255), .A2(SI_24_), .ZN(n8272) );
  NAND2_X1 U7389 ( .A1(n6917), .A2(n9547), .ZN(n10836) );
  AND2_X1 U7390 ( .A1(n9978), .A2(n8334), .ZN(n7424) );
  NAND2_X1 U7391 ( .A1(n8256), .A2(n12296), .ZN(n8257) );
  OAI21_X1 U7392 ( .B1(n8253), .B2(n8252), .A(n7465), .ZN(n8256) );
  INV_X1 U7393 ( .A(n13064), .ZN(n13487) );
  NAND2_X1 U7394 ( .A1(n8223), .A2(n8222), .ZN(n8253) );
  NAND2_X1 U7395 ( .A1(n8633), .A2(n8632), .ZN(n14201) );
  AND2_X1 U7396 ( .A1(n8163), .A2(n8146), .ZN(n8147) );
  AND2_X1 U7397 ( .A1(n9282), .A2(n9281), .ZN(n13064) );
  NAND2_X1 U7398 ( .A1(n8659), .A2(n8658), .ZN(n14086) );
  NAND2_X1 U7399 ( .A1(n6767), .A2(n8202), .ZN(n8223) );
  INV_X1 U7400 ( .A(n11465), .ZN(n7698) );
  OAI21_X1 U7401 ( .B1(n7459), .B2(n6488), .A(n6765), .ZN(n6767) );
  NAND2_X1 U7402 ( .A1(n7461), .A2(n7462), .ZN(n8190) );
  NAND2_X1 U7403 ( .A1(n9786), .A2(n15434), .ZN(n15332) );
  NAND2_X2 U7404 ( .A1(n8581), .A2(n8580), .ZN(n12711) );
  NAND2_X1 U7405 ( .A1(n7974), .A2(n7975), .ZN(n12044) );
  OR2_X1 U7406 ( .A1(n8129), .A2(n7464), .ZN(n7461) );
  INV_X2 U7407 ( .A(n15305), .ZN(n15307) );
  OAI21_X2 U7408 ( .B1(n10392), .B2(n15291), .A(n14997), .ZN(n10393) );
  NAND2_X1 U7409 ( .A1(n8129), .A2(n6455), .ZN(n7459) );
  INV_X1 U7410 ( .A(n11213), .ZN(n11120) );
  INV_X2 U7411 ( .A(n9777), .ZN(n9771) );
  NAND2_X1 U7412 ( .A1(n12933), .A2(n6875), .ZN(n8836) );
  NAND2_X2 U7413 ( .A1(n14072), .A2(n12901), .ZN(n9726) );
  OR2_X1 U7414 ( .A1(n13211), .A2(n11372), .ZN(n12425) );
  OR2_X2 U7415 ( .A1(n14222), .A2(n11404), .ZN(n12728) );
  CLKBUF_X1 U7416 ( .A(n9657), .Z(n13017) );
  NAND2_X1 U7417 ( .A1(n12417), .A2(n12418), .ZN(n12547) );
  AND3_X1 U7418 ( .A1(n9028), .A2(n9027), .A3(n9026), .ZN(n11372) );
  AND2_X1 U7419 ( .A1(n9047), .A2(n9046), .ZN(n11673) );
  NAND3_X1 U7420 ( .A1(n7963), .A2(n7965), .A3(n7964), .ZN(n7968) );
  NAND2_X1 U7421 ( .A1(n6868), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8045) );
  NOR2_X1 U7422 ( .A1(n13214), .A2(n12579), .ZN(n13270) );
  NAND2_X1 U7423 ( .A1(n8503), .A2(n8504), .ZN(n12683) );
  CLKBUF_X1 U7424 ( .A(n15543), .Z(n15531) );
  AND3_X1 U7425 ( .A1(n8992), .A2(n8991), .A3(n8990), .ZN(n11328) );
  NOR2_X1 U7426 ( .A1(n8827), .A2(n11173), .ZN(n12663) );
  INV_X1 U7427 ( .A(n8029), .ZN(n6868) );
  NAND4_X2 U7428 ( .A1(n9020), .A2(n9019), .A3(n9018), .A4(n9017), .ZN(n13211)
         );
  NAND2_X2 U7429 ( .A1(n6487), .A2(n7855), .ZN(n14583) );
  NAND2_X2 U7430 ( .A1(n12582), .A2(n12394), .ZN(n12524) );
  NAND2_X1 U7431 ( .A1(n6761), .A2(n6758), .ZN(n6757) );
  NAND4_X2 U7432 ( .A1(n7805), .A2(n7806), .A3(n7803), .A4(n7804), .ZN(n14587)
         );
  NAND2_X2 U7433 ( .A1(n10379), .A2(n10383), .ZN(n14414) );
  AND3_X1 U7434 ( .A1(n8474), .A2(n8473), .A3(n8472), .ZN(n11397) );
  NAND2_X2 U7435 ( .A1(n6737), .A2(n6736), .ZN(n10383) );
  NAND2_X1 U7436 ( .A1(n10449), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10774) );
  INV_X1 U7437 ( .A(n10379), .ZN(n10380) );
  AOI21_X1 U7438 ( .B1(n8123), .B2(n6558), .A(n8122), .ZN(n8124) );
  INV_X2 U7439 ( .A(n7835), .ZN(n10032) );
  INV_X1 U7440 ( .A(n6435), .ZN(n9260) );
  AOI22_X1 U7441 ( .A1(n8702), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10412), .B2(
        n10499), .ZN(n8503) );
  AOI21_X1 U7442 ( .B1(n8143), .B2(n7463), .A(n6567), .ZN(n7462) );
  XNOR2_X1 U7443 ( .A(n9241), .B(n9240), .ZN(n11153) );
  NOR2_X1 U7444 ( .A1(n6759), .A2(n6755), .ZN(n6754) );
  XNOR2_X1 U7445 ( .A(n9433), .B(n9432), .ZN(n9446) );
  INV_X2 U7446 ( .A(n7833), .ZN(n9851) );
  CLKBUF_X1 U7447 ( .A(n8471), .Z(n12824) );
  AND2_X1 U7448 ( .A1(n10772), .A2(n9535), .ZN(n10449) );
  NAND2_X1 U7449 ( .A1(n15160), .A2(n7780), .ZN(n7836) );
  OR2_X1 U7450 ( .A1(n9534), .A2(n10462), .ZN(n9535) );
  INV_X1 U7451 ( .A(n8933), .ZN(n12617) );
  AND2_X1 U7452 ( .A1(n7778), .A2(n7779), .ZN(n7833) );
  OR2_X1 U7453 ( .A1(n8690), .A2(n11170), .ZN(n8453) );
  NAND2_X1 U7454 ( .A1(n8447), .A2(n10171), .ZN(n8757) );
  INV_X2 U7455 ( .A(n8485), .ZN(n12816) );
  XNOR2_X1 U7456 ( .A(n6662), .B(n11906), .ZN(n9422) );
  NAND2_X1 U7457 ( .A1(n8812), .A2(n8811), .ZN(n12906) );
  NAND2_X1 U7458 ( .A1(n7780), .A2(n7779), .ZN(n7871) );
  MUX2_X1 U7460 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8375), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n8376) );
  XNOR2_X1 U7461 ( .A(n8378), .B(P1_IR_REG_24__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U7462 ( .A1(n12355), .A2(n8420), .ZN(n8485) );
  AND2_X2 U7463 ( .A1(n12355), .A2(n8438), .ZN(n8440) );
  NAND2_X1 U7464 ( .A1(n6725), .A2(n6724), .ZN(n7765) );
  NOR2_X1 U7465 ( .A1(n8022), .A2(n7472), .ZN(n7471) );
  INV_X1 U7466 ( .A(n7987), .ZN(n7988) );
  OR2_X1 U7467 ( .A1(n7761), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U7468 ( .A1(n6703), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6662) );
  XNOR2_X1 U7469 ( .A(n8813), .B(P2_IR_REG_21__SCAN_IN), .ZN(n12899) );
  NAND2_X1 U7470 ( .A1(n7761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7758) );
  NAND2_X1 U7471 ( .A1(n13697), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8928) );
  MUX2_X1 U7472 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8810), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8812) );
  NAND2_X1 U7473 ( .A1(n10619), .A2(n9532), .ZN(n10564) );
  NAND2_X1 U7474 ( .A1(n7013), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U7475 ( .A1(n8815), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8813) );
  NAND2_X2 U7476 ( .A1(n10039), .A2(P1_U3086), .ZN(n15165) );
  NAND2_X1 U7477 ( .A1(n15152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7776) );
  XNOR2_X1 U7478 ( .A(n8435), .B(n8434), .ZN(n10420) );
  NAND2_X1 U7479 ( .A1(n9112), .A2(n6854), .ZN(n7350) );
  NOR2_X1 U7480 ( .A1(n8433), .A2(n6568), .ZN(n7062) );
  XNOR2_X1 U7481 ( .A(n8491), .B(n8490), .ZN(n15348) );
  NAND2_X1 U7482 ( .A1(n7923), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7947) );
  OR2_X1 U7483 ( .A1(n8819), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n8815) );
  NOR2_X1 U7484 ( .A1(n7774), .A2(n7759), .ZN(n7760) );
  AND2_X2 U7485 ( .A1(n7012), .A2(n6503), .ZN(n6717) );
  OR2_X1 U7486 ( .A1(n9004), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9041) );
  AND3_X1 U7487 ( .A1(n6609), .A2(n7284), .A3(n7283), .ZN(n9618) );
  NAND3_X1 U7488 ( .A1(n8418), .A2(n8809), .A3(n8498), .ZN(n8433) );
  AND2_X1 U7489 ( .A1(n8605), .A2(n6512), .ZN(n8617) );
  CLKBUF_X3 U7490 ( .A(n7790), .Z(n10193) );
  BUF_X4 U7491 ( .A(n7818), .Z(n6439) );
  OR2_X1 U7492 ( .A1(n9111), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9004) );
  AND2_X1 U7493 ( .A1(n7754), .A2(n7753), .ZN(n8080) );
  AND3_X1 U7494 ( .A1(n9530), .A2(n8921), .A3(n7188), .ZN(n8925) );
  AND4_X1 U7495 ( .A1(n6750), .A2(n6747), .A3(n8523), .A4(n6746), .ZN(n6745)
         );
  AND3_X1 U7496 ( .A1(n6653), .A2(n6652), .A3(n8920), .ZN(n9055) );
  AND4_X1 U7497 ( .A1(n7752), .A2(n7750), .A3(n7751), .A4(n11887), .ZN(n6775)
         );
  AND4_X2 U7498 ( .A1(n7825), .A2(n7755), .A3(n7756), .A4(n7011), .ZN(n7903)
         );
  MUX2_X1 U7499 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8940), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n8942) );
  NOR2_X1 U7500 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n7772) );
  NOR2_X1 U7501 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n6652) );
  NOR2_X1 U7502 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n6653) );
  INV_X1 U7503 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n11988) );
  NOR2_X1 U7504 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7755) );
  NOR2_X1 U7505 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n7756) );
  NOR2_X1 U7506 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7750) );
  NOR2_X1 U7507 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7751) );
  OR2_X1 U7508 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n8427) );
  INV_X1 U7509 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7796) );
  NOR2_X1 U7510 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6750) );
  INV_X1 U7511 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8417) );
  NOR2_X1 U7512 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n6692) );
  INV_X1 U7513 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9240) );
  INV_X1 U7514 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9237) );
  NOR2_X1 U7515 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n6747) );
  INV_X1 U7516 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9239) );
  INV_X1 U7517 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n11887) );
  NOR2_X1 U7518 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6746) );
  INV_X4 U7519 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7520 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n6688) );
  INV_X2 U7521 ( .A(n7871), .ZN(n7851) );
  XNOR2_X2 U7522 ( .A(n7776), .B(n7775), .ZN(n7780) );
  NAND2_X1 U7523 ( .A1(n7851), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7806) );
  NAND2_X1 U7524 ( .A1(n11833), .A2(n11836), .ZN(n8333) );
  NAND2_X1 U7525 ( .A1(n7416), .A2(n6441), .ZN(n6440) );
  NAND2_X1 U7526 ( .A1(n14859), .A2(n6442), .ZN(n14861) );
  NAND2_X2 U7527 ( .A1(n11093), .A2(n11099), .ZN(n11092) );
  INV_X1 U7528 ( .A(n8323), .ZN(n11093) );
  NAND3_X2 U7529 ( .A1(n6757), .A2(n6756), .A3(n6753), .ZN(n8120) );
  INV_X1 U7530 ( .A(n12366), .ZN(n6444) );
  OR2_X2 U7531 ( .A1(n13234), .A2(n7295), .ZN(n7294) );
  INV_X4 U7532 ( .A(n7871), .ZN(n9866) );
  NAND4_X4 U7533 ( .A1(n7784), .A2(n7783), .A3(n7782), .A4(n7781), .ZN(n10474)
         );
  NAND2_X1 U7534 ( .A1(n7833), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7782) );
  OAI21_X2 U7535 ( .B1(n13952), .B2(n8781), .A(n7685), .ZN(n6878) );
  NOR2_X1 U7536 ( .A1(n6994), .A2(n6993), .ZN(n6445) );
  NOR2_X1 U7537 ( .A1(n6994), .A2(n6993), .ZN(n15443) );
  INV_X2 U7538 ( .A(n6433), .ZN(n7686) );
  XNOR2_X1 U7539 ( .A(n14584), .B(n6433), .ZN(n10073) );
  OR2_X1 U7540 ( .A1(n14222), .A2(n11404), .ZN(n6446) );
  OR2_X2 U7541 ( .A1(n14222), .A2(n11404), .ZN(n6447) );
  AND2_X2 U7542 ( .A1(n8367), .A2(n8366), .ZN(n15033) );
  OAI22_X2 U7543 ( .A1(n14032), .A2(n8711), .B1(n13771), .B2(n14033), .ZN(
        n14023) );
  NOR2_X2 U7544 ( .A1(n9189), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9203) );
  OR2_X2 U7545 ( .A1(n9171), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9189) );
  INV_X2 U7546 ( .A(n14048), .ZN(n14173) );
  NAND2_X2 U7547 ( .A1(n8686), .A2(n8685), .ZN(n14048) );
  NOR2_X2 U7548 ( .A1(n9031), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9060) );
  OAI222_X1 U7549 ( .A1(P3_U3151), .A2(n10634), .B1(n13719), .B2(n10176), .C1(
        n13717), .C2(n10175), .ZN(P3_U3294) );
  INV_X2 U7550 ( .A(n13702), .ZN(n13717) );
  NAND2_X1 U7551 ( .A1(n12850), .A2(n7136), .ZN(n12853) );
  NAND2_X1 U7552 ( .A1(n12840), .A2(n12841), .ZN(n7136) );
  INV_X1 U7553 ( .A(n7371), .ZN(n7370) );
  OAI21_X1 U7554 ( .B1(n6461), .B2(n13038), .A(n6533), .ZN(n7371) );
  XNOR2_X1 U7555 ( .A(n13403), .B(n13385), .ZN(n12510) );
  AND2_X1 U7556 ( .A1(n13430), .A2(n9332), .ZN(n9347) );
  AND2_X1 U7557 ( .A1(n13630), .A2(n13077), .ZN(n12380) );
  AOI21_X1 U7558 ( .B1(n7650), .B2(n7653), .A(n6565), .ZN(n7649) );
  INV_X1 U7559 ( .A(n6808), .ZN(n6807) );
  OAI21_X1 U7560 ( .B1(n7547), .B2(n6809), .A(n9235), .ZN(n6808) );
  AND2_X1 U7561 ( .A1(n8858), .A2(n7599), .ZN(n7598) );
  NAND2_X1 U7562 ( .A1(n7601), .A2(n7600), .ZN(n7599) );
  NOR2_X1 U7563 ( .A1(n8301), .A2(SI_26_), .ZN(n6769) );
  OR2_X1 U7564 ( .A1(n13630), .A2(n13077), .ZN(n12527) );
  AND2_X1 U7565 ( .A1(n9225), .A2(n9224), .ZN(n13027) );
  NAND2_X1 U7566 ( .A1(n13499), .A2(n6530), .ZN(n7352) );
  INV_X1 U7567 ( .A(n12478), .ZN(n7353) );
  NOR2_X1 U7568 ( .A1(n7688), .A2(n14780), .ZN(n7687) );
  NAND2_X1 U7569 ( .A1(n14768), .A2(n10027), .ZN(n7688) );
  AOI21_X1 U7570 ( .B1(n7723), .B2(n7721), .A(n6556), .ZN(n14848) );
  NOR2_X1 U7571 ( .A1(n8234), .A2(n7722), .ZN(n7721) );
  INV_X1 U7572 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7011) );
  AOI21_X1 U7573 ( .B1(n9897), .B2(n9896), .A(n7735), .ZN(n9902) );
  NAND2_X1 U7574 ( .A1(n7052), .A2(n12705), .ZN(n7051) );
  NAND2_X1 U7575 ( .A1(n7455), .A2(n7055), .ZN(n7052) );
  AOI21_X1 U7576 ( .B1(n7128), .B2(n7126), .A(n7124), .ZN(n7123) );
  INV_X1 U7577 ( .A(n9930), .ZN(n7124) );
  NOR2_X1 U7578 ( .A1(n7117), .A2(n7116), .ZN(n7115) );
  AND2_X1 U7579 ( .A1(n9997), .A2(n9996), .ZN(n7117) );
  NOR2_X1 U7580 ( .A1(n12853), .A2(n12829), .ZN(n12833) );
  NAND2_X1 U7581 ( .A1(n7573), .A2(n7572), .ZN(n6931) );
  AND2_X1 U7582 ( .A1(n8836), .A2(n8835), .ZN(n7572) );
  AOI21_X1 U7583 ( .B1(n7509), .B2(n7508), .A(n6841), .ZN(n7506) );
  INV_X1 U7584 ( .A(n15048), .ZN(n9888) );
  NAND2_X1 U7585 ( .A1(n6511), .A2(n9991), .ZN(n7435) );
  INV_X1 U7586 ( .A(n8018), .ZN(n6783) );
  INV_X1 U7587 ( .A(n7487), .ZN(n7486) );
  OAI21_X1 U7588 ( .B1(n7491), .B2(n7488), .A(n10036), .ZN(n7487) );
  INV_X1 U7589 ( .A(n8074), .ZN(n8076) );
  NOR2_X1 U7590 ( .A1(n8073), .A2(n10469), .ZN(n8075) );
  AND2_X1 U7591 ( .A1(n7246), .A2(n7245), .ZN(n9619) );
  NAND2_X1 U7592 ( .A1(n10186), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7245) );
  INV_X1 U7593 ( .A(n9357), .ZN(n9356) );
  OR2_X1 U7594 ( .A1(n13639), .A2(n13429), .ZN(n12502) );
  AND2_X1 U7595 ( .A1(n13465), .A2(n12481), .ZN(n7351) );
  INV_X1 U7596 ( .A(n12465), .ZN(n12469) );
  NAND2_X1 U7597 ( .A1(n9422), .A2(n9424), .ZN(n8939) );
  AOI21_X1 U7598 ( .B1(n7344), .B2(n7341), .A(n12452), .ZN(n7338) );
  OR2_X1 U7599 ( .A1(n10271), .A2(n10268), .ZN(n9511) );
  NAND2_X1 U7600 ( .A1(n9336), .A2(n9335), .ZN(n9350) );
  INV_X1 U7601 ( .A(n9233), .ZN(n6809) );
  INV_X1 U7602 ( .A(n9071), .ZN(n7531) );
  NOR2_X1 U7603 ( .A1(n8772), .A2(n8771), .ZN(n7187) );
  INV_X1 U7604 ( .A(n11144), .ZN(n7151) );
  NAND2_X1 U7605 ( .A1(n8409), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8761) );
  INV_X1 U7606 ( .A(n8749), .ZN(n8409) );
  OR2_X1 U7607 ( .A1(n8761), .A2(n8760), .ZN(n8772) );
  INV_X1 U7608 ( .A(n12721), .ZN(n7602) );
  XNOR2_X1 U7609 ( .A(n12711), .B(n12262), .ZN(n12881) );
  NOR2_X1 U7610 ( .A1(n13925), .A2(n7679), .ZN(n7678) );
  INV_X1 U7611 ( .A(n7680), .ZN(n7679) );
  NAND2_X1 U7612 ( .A1(n14119), .A2(n13840), .ZN(n7683) );
  NOR2_X1 U7613 ( .A1(n8652), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8656) );
  INV_X1 U7614 ( .A(n7626), .ZN(n7625) );
  NAND2_X1 U7615 ( .A1(n14785), .A2(n8299), .ZN(n8356) );
  INV_X1 U7616 ( .A(n14989), .ZN(n7430) );
  AOI21_X1 U7617 ( .B1(n7715), .B2(n7719), .A(n6466), .ZN(n7714) );
  NAND2_X1 U7618 ( .A1(n12098), .A2(n7718), .ZN(n7717) );
  INV_X1 U7619 ( .A(n7986), .ZN(n7718) );
  NOR2_X1 U7620 ( .A1(n14770), .A2(n7710), .ZN(n7709) );
  INV_X1 U7621 ( .A(n9877), .ZN(n7710) );
  INV_X1 U7622 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7773) );
  OAI21_X2 U7623 ( .B1(n8287), .B2(n8286), .A(n8285), .ZN(n8302) );
  XNOR2_X1 U7624 ( .A(n8145), .B(SI_17_), .ZN(n8143) );
  NOR2_X1 U7625 ( .A1(n8072), .A2(SI_14_), .ZN(n8119) );
  NOR2_X1 U7626 ( .A1(n8076), .A2(n8075), .ZN(n8121) );
  XNOR2_X1 U7627 ( .A(n8019), .B(SI_11_), .ZN(n8022) );
  NAND3_X1 U7628 ( .A1(n10162), .A2(n10198), .A3(n7297), .ZN(n10223) );
  AOI21_X1 U7629 ( .B1(n11616), .B2(n11615), .A(n11614), .ZN(n11622) );
  INV_X1 U7630 ( .A(n13043), .ZN(n7365) );
  AOI21_X1 U7631 ( .B1(n7379), .B2(n7382), .A(n6569), .ZN(n7378) );
  INV_X1 U7632 ( .A(n7380), .ZN(n7379) );
  OAI21_X1 U7633 ( .B1(n13023), .B2(n7382), .A(n7381), .ZN(n7380) );
  INV_X1 U7634 ( .A(n13188), .ZN(n7381) );
  INV_X1 U7635 ( .A(n7376), .ZN(n7375) );
  OR2_X1 U7636 ( .A1(n13030), .A2(n13490), .ZN(n13031) );
  AND3_X1 U7637 ( .A1(n9207), .A2(n9206), .A3(n9205), .ZN(n13192) );
  NAND2_X1 U7638 ( .A1(n7088), .A2(n7087), .ZN(n10451) );
  OAI21_X1 U7639 ( .B1(n10566), .B2(n7089), .A(n10166), .ZN(n7088) );
  INV_X1 U7640 ( .A(n7092), .ZN(n7089) );
  NAND2_X1 U7641 ( .A1(n13219), .A2(n13218), .ZN(n13238) );
  OAI211_X1 U7642 ( .C1(n13300), .C2(n7232), .A(n13310), .B(n7231), .ZN(n13335) );
  OR2_X1 U7643 ( .A1(n13312), .A2(n13299), .ZN(n7232) );
  NAND2_X1 U7644 ( .A1(n9605), .A2(n7230), .ZN(n7231) );
  NOR2_X1 U7645 ( .A1(n13312), .A2(n10672), .ZN(n7230) );
  XNOR2_X1 U7646 ( .A(n7202), .B(n13354), .ZN(n13344) );
  AND2_X1 U7647 ( .A1(n9298), .A2(n9297), .ZN(n13474) );
  INV_X1 U7648 ( .A(n12547), .ZN(n6699) );
  NAND2_X1 U7649 ( .A1(n10146), .A2(n9406), .ZN(n9821) );
  NAND2_X1 U7650 ( .A1(n9650), .A2(n15596), .ZN(n6669) );
  AND2_X1 U7651 ( .A1(n9648), .A2(n9649), .ZN(n6672) );
  AOI21_X1 U7652 ( .B1(n9283), .B2(n6468), .A(n6571), .ZN(n7005) );
  OR2_X1 U7653 ( .A1(n12524), .A2(n10889), .ZN(n15508) );
  AND2_X1 U7654 ( .A1(n9481), .A2(n12473), .ZN(n6675) );
  NAND2_X1 U7655 ( .A1(n13531), .A2(n12468), .ZN(n13522) );
  AOI21_X1 U7656 ( .B1(n7652), .B2(n7651), .A(n6559), .ZN(n7650) );
  INV_X1 U7657 ( .A(n7744), .ZN(n7651) );
  AND2_X1 U7658 ( .A1(n6645), .A2(n9396), .ZN(n7560) );
  NAND2_X1 U7659 ( .A1(n6806), .A2(n6804), .ZN(n9305) );
  AOI21_X1 U7660 ( .B1(n6807), .B2(n6809), .A(n6805), .ZN(n6804) );
  NAND2_X1 U7661 ( .A1(n7549), .A2(n6807), .ZN(n6806) );
  INV_X1 U7662 ( .A(n9271), .ZN(n6805) );
  XNOR2_X1 U7663 ( .A(n9305), .B(n11383), .ZN(n9286) );
  AND2_X1 U7664 ( .A1(n9271), .A2(n9234), .ZN(n9235) );
  OAI21_X1 U7665 ( .B1(n7549), .B2(n6809), .A(n6807), .ZN(n9272) );
  NAND2_X1 U7666 ( .A1(n7549), .A2(n7547), .ZN(n9253) );
  OAI21_X1 U7667 ( .B1(n9196), .B2(n6813), .A(n6811), .ZN(n9212) );
  INV_X1 U7668 ( .A(n6812), .ZN(n6811) );
  OAI21_X1 U7669 ( .B1(n9195), .B2(n6813), .A(n9209), .ZN(n6812) );
  INV_X1 U7670 ( .A(n9197), .ZN(n6813) );
  NAND2_X1 U7671 ( .A1(n9146), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U7672 ( .A1(n7545), .A2(n7543), .ZN(n9143) );
  NOR2_X1 U7673 ( .A1(n9128), .A2(n7544), .ZN(n7543) );
  INV_X1 U7674 ( .A(n9124), .ZN(n7544) );
  AOI21_X1 U7675 ( .B1(n7527), .B2(n7530), .A(n6818), .ZN(n6817) );
  INV_X1 U7676 ( .A(n9103), .ZN(n6818) );
  INV_X1 U7677 ( .A(n7527), .ZN(n6819) );
  XNOR2_X1 U7678 ( .A(n9025), .B(P3_IR_REG_6__SCAN_IN), .ZN(n9620) );
  AND2_X1 U7679 ( .A1(n13809), .A2(n6519), .ZN(n7258) );
  INV_X1 U7680 ( .A(n9777), .ZN(n12992) );
  OR2_X1 U7681 ( .A1(n13726), .A2(n9759), .ZN(n9764) );
  XNOR2_X1 U7682 ( .A(n9726), .B(n12683), .ZN(n12927) );
  NAND2_X1 U7683 ( .A1(n6984), .A2(n6982), .ZN(n11312) );
  NOR2_X1 U7684 ( .A1(n15328), .A2(n6983), .ZN(n6982) );
  INV_X1 U7685 ( .A(n9668), .ZN(n6983) );
  INV_X1 U7686 ( .A(n7269), .ZN(n7267) );
  NAND2_X1 U7687 ( .A1(n13017), .A2(n11381), .ZN(n12905) );
  INV_X1 U7688 ( .A(n8690), .ZN(n8787) );
  INV_X1 U7689 ( .A(n12355), .ZN(n8450) );
  OAI21_X1 U7690 ( .B1(n8485), .B2(n8439), .A(n6739), .ZN(n6738) );
  NAND2_X1 U7691 ( .A1(n8420), .A2(n6740), .ZN(n6739) );
  NOR2_X1 U7692 ( .A1(n12355), .A2(n10636), .ZN(n6740) );
  NAND2_X1 U7693 ( .A1(n13838), .A2(n13801), .ZN(n12962) );
  INV_X1 U7694 ( .A(n8872), .ZN(n7590) );
  AOI21_X1 U7695 ( .B1(n6460), .B2(n7578), .A(n6548), .ZN(n7575) );
  XNOR2_X1 U7696 ( .A(n13970), .B(n13842), .ZN(n13963) );
  AOI21_X1 U7697 ( .B1(n6453), .B2(n8722), .A(n6557), .ZN(n7660) );
  AOI21_X1 U7698 ( .B1(n7646), .B2(n12885), .A(n6537), .ZN(n7644) );
  NAND2_X1 U7699 ( .A1(n9657), .A2(n8817), .ZN(n14072) );
  INV_X1 U7700 ( .A(n14186), .ZN(n15479) );
  NAND2_X1 U7701 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n7067) );
  AND2_X1 U7702 ( .A1(n14383), .A2(n6502), .ZN(n6731) );
  INV_X1 U7703 ( .A(n14768), .ZN(n15041) );
  NAND2_X1 U7704 ( .A1(n14450), .A2(n14451), .ZN(n14357) );
  AND2_X1 U7705 ( .A1(n14461), .A2(n14463), .ZN(n7620) );
  AND2_X1 U7706 ( .A1(n10382), .A2(n7629), .ZN(n10388) );
  NAND2_X1 U7707 ( .A1(n14587), .A2(n10794), .ZN(n7629) );
  NAND2_X1 U7708 ( .A1(n7021), .A2(n7023), .ZN(n7018) );
  NAND2_X1 U7709 ( .A1(n14462), .A2(n7021), .ZN(n7019) );
  INV_X1 U7710 ( .A(n10262), .ZN(n10390) );
  NOR2_X1 U7711 ( .A1(n10116), .A2(n7494), .ZN(n10141) );
  INV_X1 U7712 ( .A(n7495), .ZN(n7494) );
  AOI21_X1 U7713 ( .B1(n10114), .B2(n10115), .A(n11734), .ZN(n7495) );
  INV_X1 U7714 ( .A(n7836), .ZN(n10029) );
  NOR2_X1 U7715 ( .A1(n7008), .A2(n15157), .ZN(n9850) );
  OAI22_X1 U7716 ( .A1(n10090), .A2(n6972), .B1(n15041), .B2(n15033), .ZN(
        n6971) );
  NAND2_X1 U7717 ( .A1(n14763), .A2(n14768), .ZN(n14762) );
  AND2_X1 U7718 ( .A1(n14793), .A2(n14365), .ZN(n14763) );
  AND2_X1 U7719 ( .A1(n14806), .A2(n15048), .ZN(n14793) );
  AND2_X1 U7720 ( .A1(n14828), .A2(n14810), .ZN(n14806) );
  AND2_X1 U7721 ( .A1(n7693), .A2(n7692), .ZN(n7691) );
  INV_X1 U7722 ( .A(n15061), .ZN(n7692) );
  NOR2_X1 U7723 ( .A1(n8221), .A2(n7724), .ZN(n7720) );
  INV_X1 U7724 ( .A(n8179), .ZN(n7724) );
  NOR2_X1 U7725 ( .A1(n8371), .A2(n10092), .ZN(n10371) );
  NAND2_X1 U7726 ( .A1(n9878), .A2(n9877), .ZN(n14771) );
  INV_X1 U7727 ( .A(n15314), .ZN(n15078) );
  XNOR2_X1 U7728 ( .A(n8381), .B(P1_IR_REG_26__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U7729 ( .A1(n8257), .A2(n8272), .ZN(n8260) );
  NAND2_X1 U7730 ( .A1(n10960), .A2(n10302), .ZN(n10307) );
  NAND2_X1 U7731 ( .A1(n10299), .A2(n10959), .ZN(n10301) );
  NOR2_X1 U7732 ( .A1(n6450), .A2(n7308), .ZN(n7307) );
  NAND2_X1 U7733 ( .A1(n7320), .A2(n13169), .ZN(n7318) );
  XNOR2_X1 U7734 ( .A(n12385), .B(n11153), .ZN(n6679) );
  AND2_X1 U7735 ( .A1(n13392), .A2(n13393), .ZN(n13575) );
  INV_X1 U7736 ( .A(n13826), .ZN(n15325) );
  OAI21_X1 U7737 ( .B1(n10070), .B2(n10069), .A(n10026), .ZN(n7109) );
  OR2_X1 U7738 ( .A1(n6448), .A2(n15223), .ZN(n6825) );
  MUX2_X1 U7739 ( .A(n6447), .B(n12662), .S(n12661), .Z(n7437) );
  NOR2_X1 U7740 ( .A1(n7077), .A2(n12686), .ZN(n7074) );
  INV_X1 U7741 ( .A(n12684), .ZN(n7077) );
  INV_X1 U7742 ( .A(n12679), .ZN(n7441) );
  NOR2_X1 U7743 ( .A1(n12682), .A2(n12679), .ZN(n7442) );
  NOR2_X1 U7744 ( .A1(n7074), .A2(n7447), .ZN(n7073) );
  INV_X1 U7745 ( .A(n7446), .ZN(n7070) );
  NOR2_X1 U7746 ( .A1(n12691), .A2(n12688), .ZN(n7447) );
  NAND2_X1 U7747 ( .A1(n12691), .A2(n12688), .ZN(n7446) );
  INV_X1 U7748 ( .A(n7074), .ZN(n7072) );
  NAND2_X1 U7749 ( .A1(n9925), .A2(n7127), .ZN(n7126) );
  INV_X1 U7750 ( .A(n9921), .ZN(n7518) );
  NAND2_X1 U7751 ( .A1(n12701), .A2(n7056), .ZN(n7055) );
  INV_X1 U7752 ( .A(n7126), .ZN(n6882) );
  NOR2_X1 U7753 ( .A1(n7127), .A2(n9925), .ZN(n7128) );
  NOR2_X1 U7754 ( .A1(n12710), .A2(n12707), .ZN(n7454) );
  INV_X1 U7755 ( .A(n12707), .ZN(n7453) );
  NAND2_X1 U7756 ( .A1(n6880), .A2(n6541), .ZN(n7135) );
  NAND2_X1 U7757 ( .A1(n6840), .A2(n6839), .ZN(n6880) );
  INV_X1 U7758 ( .A(n7517), .ZN(n6839) );
  INV_X1 U7759 ( .A(n12780), .ZN(n7448) );
  NOR2_X1 U7760 ( .A1(n7450), .A2(n12780), .ZN(n7449) );
  NOR2_X1 U7761 ( .A1(n9997), .A2(n9996), .ZN(n7114) );
  NAND2_X1 U7762 ( .A1(n12792), .A2(n12794), .ZN(n7452) );
  NOR2_X1 U7763 ( .A1(n6496), .A2(n6472), .ZN(n7043) );
  NOR2_X1 U7764 ( .A1(n6471), .A2(n7121), .ZN(n7120) );
  NOR2_X1 U7765 ( .A1(n7519), .A2(n10005), .ZN(n7121) );
  INV_X1 U7766 ( .A(n10003), .ZN(n7519) );
  NAND2_X1 U7767 ( .A1(n12803), .A2(n7060), .ZN(n7059) );
  NAND2_X1 U7768 ( .A1(n7499), .A2(n7498), .ZN(n10107) );
  NAND2_X1 U7769 ( .A1(n10045), .A2(n9947), .ZN(n7498) );
  NAND2_X1 U7770 ( .A1(n14756), .A2(n10066), .ZN(n7499) );
  OR2_X1 U7771 ( .A1(n9887), .A2(n15297), .ZN(n7105) );
  AOI21_X1 U7772 ( .B1(n7421), .B2(n7419), .A(n6555), .ZN(n7418) );
  INV_X1 U7773 ( .A(n8325), .ZN(n7419) );
  INV_X1 U7774 ( .A(n7421), .ZN(n7420) );
  NOR2_X1 U7775 ( .A1(n7489), .A2(n9847), .ZN(n7483) );
  NAND2_X1 U7776 ( .A1(n6478), .A2(n7490), .ZN(n7489) );
  INV_X1 U7777 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6966) );
  INV_X1 U7778 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6963) );
  AOI21_X1 U7779 ( .B1(n6455), .B2(n7464), .A(n6553), .ZN(n7460) );
  INV_X1 U7780 ( .A(n8143), .ZN(n7464) );
  NAND2_X1 U7781 ( .A1(n7936), .A2(n7938), .ZN(n7962) );
  NAND2_X1 U7782 ( .A1(n10438), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10201) );
  INV_X1 U7783 ( .A(n7331), .ZN(n7328) );
  INV_X1 U7784 ( .A(n11076), .ZN(n13035) );
  OR2_X1 U7785 ( .A1(n13361), .A2(n13363), .ZN(n12533) );
  NAND2_X1 U7786 ( .A1(n7091), .A2(n7090), .ZN(n7093) );
  INV_X1 U7787 ( .A(n10567), .ZN(n7091) );
  NAND2_X1 U7788 ( .A1(n10580), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7092) );
  NAND2_X1 U7789 ( .A1(n10188), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7241) );
  OR2_X1 U7790 ( .A1(n11307), .A2(n9624), .ZN(n7276) );
  AOI21_X1 U7791 ( .B1(n11296), .B2(n11297), .A(n7103), .ZN(n9625) );
  NAND2_X1 U7792 ( .A1(n13244), .A2(n9627), .ZN(n9628) );
  OR2_X1 U7793 ( .A1(n13582), .A2(n13417), .ZN(n12498) );
  NOR2_X1 U7794 ( .A1(n7635), .A2(n7633), .ZN(n7632) );
  INV_X1 U7795 ( .A(n9318), .ZN(n7633) );
  AND2_X1 U7796 ( .A1(n12444), .A2(n12451), .ZN(n12557) );
  INV_X1 U7797 ( .A(n15544), .ZN(n6702) );
  NAND2_X1 U7798 ( .A1(n10884), .A2(n9470), .ZN(n15523) );
  AND2_X1 U7799 ( .A1(n9469), .A2(n11019), .ZN(n12393) );
  NAND2_X1 U7800 ( .A1(n15540), .A2(n15533), .ZN(n12390) );
  NAND2_X1 U7801 ( .A1(n13415), .A2(n6497), .ZN(n9647) );
  OR2_X1 U7802 ( .A1(n7351), .A2(n7182), .ZN(n7181) );
  INV_X1 U7803 ( .A(n12490), .ZN(n7182) );
  OR2_X1 U7804 ( .A1(n13645), .A2(n13474), .ZN(n12493) );
  NAND2_X1 U7805 ( .A1(n13534), .A2(n9194), .ZN(n7642) );
  NAND2_X1 U7806 ( .A1(n9177), .A2(n7638), .ZN(n6655) );
  NOR2_X1 U7807 ( .A1(n7643), .A2(n7639), .ZN(n7638) );
  INV_X1 U7808 ( .A(n9176), .ZN(n7639) );
  NOR2_X1 U7809 ( .A1(n7003), .A2(n6648), .ZN(n6647) );
  INV_X1 U7810 ( .A(n9102), .ZN(n6648) );
  INV_X1 U7811 ( .A(n7650), .ZN(n7003) );
  INV_X1 U7812 ( .A(n7341), .ZN(n7339) );
  AND2_X1 U7813 ( .A1(n12454), .A2(n12456), .ZN(n12559) );
  NAND2_X1 U7814 ( .A1(n11688), .A2(n11689), .ZN(n6649) );
  INV_X1 U7815 ( .A(n12440), .ZN(n7345) );
  NAND2_X1 U7816 ( .A1(n8927), .A2(n8926), .ZN(n6703) );
  INV_X1 U7817 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7188) );
  XNOR2_X1 U7818 ( .A(n9461), .B(n9460), .ZN(n10853) );
  NAND2_X1 U7819 ( .A1(n9409), .A2(n7391), .ZN(n7390) );
  INV_X1 U7820 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7391) );
  NOR2_X1 U7821 ( .A1(n7350), .A2(n9408), .ZN(n9416) );
  NOR2_X1 U7822 ( .A1(n9250), .A2(n7548), .ZN(n7547) );
  INV_X1 U7823 ( .A(n9229), .ZN(n7548) );
  NAND2_X1 U7824 ( .A1(n9143), .A2(n9142), .ZN(n9144) );
  INV_X1 U7825 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n6650) );
  INV_X1 U7826 ( .A(n9008), .ZN(n7526) );
  INV_X1 U7827 ( .A(n7525), .ZN(n7524) );
  OAI21_X1 U7828 ( .B1(n9006), .B2(n7526), .A(n9021), .ZN(n7525) );
  NOR2_X1 U7829 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n8921) );
  AND2_X1 U7830 ( .A1(n12833), .A2(n12831), .ZN(n12832) );
  INV_X1 U7831 ( .A(n10486), .ZN(n7171) );
  AND2_X1 U7832 ( .A1(n7171), .A2(n15365), .ZN(n7170) );
  INV_X1 U7833 ( .A(n11141), .ZN(n7157) );
  NAND2_X1 U7834 ( .A1(n11268), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7158) );
  OAI22_X1 U7835 ( .A1(n15404), .A2(n15405), .B1(n12324), .B2(n15407), .ZN(
        n13876) );
  NAND2_X1 U7836 ( .A1(n14057), .A2(n7601), .ZN(n7597) );
  NAND2_X1 U7837 ( .A1(n14173), .A2(n7402), .ZN(n7401) );
  INV_X1 U7838 ( .A(n14181), .ZN(n7402) );
  AND2_X1 U7839 ( .A1(n7591), .A2(n6941), .ZN(n6940) );
  INV_X1 U7840 ( .A(n7592), .ZN(n7591) );
  NAND2_X1 U7841 ( .A1(n6943), .A2(n8848), .ZN(n6941) );
  OAI21_X1 U7842 ( .B1(n7595), .B2(n6495), .A(n8854), .ZN(n7592) );
  AND2_X1 U7843 ( .A1(n14073), .A2(n8651), .ZN(n7646) );
  INV_X1 U7844 ( .A(n8616), .ZN(n7670) );
  INV_X1 U7845 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n11911) );
  OR2_X1 U7846 ( .A1(n8497), .A2(n15335), .ZN(n8475) );
  INV_X1 U7847 ( .A(n11795), .ZN(n8894) );
  INV_X1 U7848 ( .A(n8811), .ZN(n8896) );
  INV_X1 U7849 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U7850 ( .A1(n8699), .A2(n8698), .ZN(n8818) );
  INV_X1 U7851 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8640) );
  AOI21_X1 U7852 ( .B1(n14539), .B2(n7618), .A(n14363), .ZN(n7617) );
  NOR2_X1 U7853 ( .A1(n10105), .A2(n10104), .ZN(n10124) );
  AND3_X1 U7854 ( .A1(n6905), .A2(n10082), .A3(n6902), .ZN(n10084) );
  NOR2_X1 U7855 ( .A1(n10089), .A2(n10088), .ZN(n6774) );
  OAI21_X1 U7856 ( .B1(n10011), .B2(n7509), .A(n6575), .ZN(n10017) );
  NOR2_X1 U7857 ( .A1(n7435), .A2(n14929), .ZN(n6974) );
  AND2_X1 U7858 ( .A1(n14924), .A2(n9988), .ZN(n7436) );
  OR2_X1 U7859 ( .A1(n7714), .A2(n6783), .ZN(n6779) );
  NOR2_X1 U7860 ( .A1(n7716), .A2(n6783), .ZN(n6781) );
  NOR2_X1 U7861 ( .A1(n10081), .A2(n7707), .ZN(n7706) );
  NOR2_X1 U7862 ( .A1(n10080), .A2(n7708), .ZN(n7707) );
  INV_X1 U7863 ( .A(n8035), .ZN(n7708) );
  AOI21_X1 U7864 ( .B1(n6540), .B2(n10073), .A(n6469), .ZN(n7712) );
  INV_X1 U7865 ( .A(n9878), .ZN(n6793) );
  INV_X1 U7866 ( .A(n7709), .ZN(n6797) );
  AND2_X1 U7867 ( .A1(n9880), .A2(n6796), .ZN(n6795) );
  INV_X1 U7868 ( .A(n10088), .ZN(n6796) );
  INV_X1 U7869 ( .A(n9880), .ZN(n6790) );
  INV_X1 U7870 ( .A(n8206), .ZN(n8199) );
  INV_X1 U7871 ( .A(n6764), .ZN(n8198) );
  AOI21_X1 U7872 ( .B1(n7459), .B2(n7460), .A(n6488), .ZN(n6764) );
  INV_X1 U7873 ( .A(n8120), .ZN(n6886) );
  NOR2_X1 U7874 ( .A1(n8074), .A2(n8119), .ZN(n6885) );
  AOI21_X1 U7875 ( .B1(n8036), .B2(n6979), .A(n6573), .ZN(n6978) );
  INV_X1 U7876 ( .A(n8021), .ZN(n6979) );
  AND2_X1 U7877 ( .A1(n7475), .A2(n8036), .ZN(n6976) );
  NAND2_X1 U7878 ( .A1(n7141), .A2(SI_10_), .ZN(n8004) );
  NAND2_X1 U7879 ( .A1(n7467), .A2(n7989), .ZN(n7470) );
  INV_X1 U7880 ( .A(n7962), .ZN(n7960) );
  NAND2_X1 U7881 ( .A1(n7938), .A2(n7939), .ZN(n7958) );
  XNOR2_X1 U7882 ( .A(n7935), .B(SI_7_), .ZN(n7939) );
  XNOR2_X1 U7883 ( .A(n7900), .B(SI_6_), .ZN(n7907) );
  NAND2_X1 U7884 ( .A1(n7298), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10198) );
  INV_X1 U7885 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U7886 ( .A1(n7299), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n7297) );
  INV_X1 U7887 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n7299) );
  NAND2_X1 U7888 ( .A1(n10980), .A2(n10979), .ZN(n11616) );
  OR2_X1 U7889 ( .A1(n10978), .A2(n14657), .ZN(n10980) );
  AOI21_X1 U7890 ( .B1(n11854), .B2(n11853), .A(n11852), .ZN(n12333) );
  OAI22_X1 U7891 ( .A1(n15182), .A2(n15181), .B1(P1_ADDR_REG_12__SCAN_IN), 
        .B2(n15180), .ZN(n15194) );
  NAND2_X1 U7892 ( .A1(n9387), .A2(n9386), .ZN(n9400) );
  XNOR2_X1 U7893 ( .A(n11076), .B(n11037), .ZN(n11072) );
  NAND2_X1 U7894 ( .A1(n7323), .A2(n7322), .ZN(n7321) );
  OAI21_X1 U7895 ( .B1(n13073), .B2(n7329), .A(n7327), .ZN(n7322) );
  NAND2_X1 U7896 ( .A1(n7325), .A2(n7324), .ZN(n7323) );
  INV_X1 U7897 ( .A(n13073), .ZN(n7325) );
  XNOR2_X1 U7898 ( .A(n6431), .B(n12426), .ZN(n13081) );
  NAND2_X1 U7899 ( .A1(n12393), .A2(n12390), .ZN(n10884) );
  AND2_X1 U7900 ( .A1(n6525), .A2(n7386), .ZN(n7385) );
  OR2_X1 U7901 ( .A1(n11603), .A2(n7387), .ZN(n7386) );
  OR2_X1 U7902 ( .A1(n12172), .A2(n12448), .ZN(n12021) );
  INV_X1 U7903 ( .A(n12019), .ZN(n7387) );
  XNOR2_X1 U7904 ( .A(n11076), .B(n6700), .ZN(n11036) );
  OR2_X1 U7905 ( .A1(n10872), .A2(n10871), .ZN(n10890) );
  AND2_X1 U7906 ( .A1(n13624), .A2(n13363), .ZN(n7348) );
  INV_X1 U7907 ( .A(n11640), .ZN(n9513) );
  AND3_X1 U7908 ( .A1(n9175), .A2(n9174), .A3(n9173), .ZN(n12028) );
  AND4_X1 U7909 ( .A1(n9141), .A2(n9140), .A3(n9139), .A4(n9138), .ZN(n13161)
         );
  AND4_X1 U7910 ( .A1(n9122), .A2(n9121), .A3(n9120), .A4(n9119), .ZN(n13157)
         );
  NAND2_X1 U7911 ( .A1(n12617), .A2(n8932), .ZN(n9015) );
  NOR2_X1 U7912 ( .A1(n10663), .A2(n10621), .ZN(n10620) );
  NOR2_X1 U7913 ( .A1(n7228), .A2(n9581), .ZN(n7227) );
  INV_X1 U7914 ( .A(n10457), .ZN(n7228) );
  INV_X1 U7915 ( .A(n10769), .ZN(n7224) );
  NAND2_X1 U7916 ( .A1(n10741), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U7917 ( .A1(n7096), .A2(n10746), .ZN(n7099) );
  INV_X1 U7918 ( .A(n9619), .ZN(n7096) );
  NAND2_X1 U7919 ( .A1(n7095), .A2(n7094), .ZN(n7098) );
  NAND2_X1 U7920 ( .A1(n9619), .A2(n6489), .ZN(n7095) );
  OAI22_X1 U7921 ( .A1(n9619), .A2(n6549), .B1(n10825), .B2(n9584), .ZN(n7094)
         );
  NAND2_X1 U7922 ( .A1(n6474), .A2(n6641), .ZN(n7209) );
  INV_X1 U7923 ( .A(n11410), .ZN(n7212) );
  NOR2_X1 U7924 ( .A1(n7215), .A2(n7214), .ZN(n7213) );
  NAND2_X1 U7925 ( .A1(n7220), .A2(n11410), .ZN(n7214) );
  NAND2_X1 U7926 ( .A1(n7208), .A2(n7206), .ZN(n11298) );
  NOR2_X1 U7927 ( .A1(n7209), .A2(n7207), .ZN(n7206) );
  INV_X1 U7928 ( .A(n11300), .ZN(n7207) );
  NOR2_X1 U7929 ( .A1(n11418), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7102) );
  NAND2_X1 U7930 ( .A1(n7238), .A2(n7241), .ZN(n7235) );
  INV_X1 U7931 ( .A(n7239), .ZN(n7238) );
  INV_X1 U7932 ( .A(n7102), .ZN(n7101) );
  NAND2_X1 U7933 ( .A1(n13238), .A2(n6620), .ZN(n13255) );
  XNOR2_X1 U7934 ( .A(n9635), .B(n9634), .ZN(n13330) );
  NAND2_X1 U7935 ( .A1(n13347), .A2(n13346), .ZN(n7290) );
  NAND2_X1 U7936 ( .A1(n9323), .A2(n6908), .ZN(n9357) );
  INV_X1 U7937 ( .A(n6912), .ZN(n9265) );
  INV_X1 U7938 ( .A(n12557), .ZN(n11689) );
  AOI21_X1 U7939 ( .B1(n7636), .B2(n6563), .A(n6486), .ZN(n7000) );
  NAND2_X1 U7940 ( .A1(n9494), .A2(n9493), .ZN(n13435) );
  OAI22_X1 U7941 ( .A1(n12391), .A2(n15547), .B1(n6659), .B2(n15533), .ZN(
        n15529) );
  NOR2_X1 U7942 ( .A1(n9563), .A2(n15541), .ZN(n10869) );
  NAND2_X1 U7943 ( .A1(n6680), .A2(n7346), .ZN(n12381) );
  NAND2_X1 U7944 ( .A1(n6588), .A2(n12523), .ZN(n7346) );
  INV_X1 U7945 ( .A(n12570), .ZN(n9829) );
  NAND2_X1 U7946 ( .A1(n10148), .A2(n10147), .ZN(n7658) );
  OR2_X1 U7947 ( .A1(n10144), .A2(n9394), .ZN(n10145) );
  NAND2_X1 U7948 ( .A1(n13455), .A2(n9300), .ZN(n13445) );
  INV_X1 U7949 ( .A(n13454), .ZN(n9299) );
  AND2_X1 U7950 ( .A1(n13514), .A2(n9227), .ZN(n6921) );
  AND2_X1 U7951 ( .A1(n12493), .A2(n12494), .ZN(n13454) );
  NAND2_X1 U7952 ( .A1(n7352), .A2(n7351), .ZN(n13463) );
  NAND2_X1 U7953 ( .A1(n13514), .A2(n9227), .ZN(n7631) );
  INV_X1 U7954 ( .A(n13502), .ZN(n9481) );
  AND2_X1 U7955 ( .A1(n9226), .A2(n12473), .ZN(n13513) );
  NAND2_X1 U7956 ( .A1(n13522), .A2(n13523), .ZN(n9480) );
  NAND2_X1 U7957 ( .A1(n13510), .A2(n13513), .ZN(n13511) );
  AND2_X1 U7958 ( .A1(n12470), .A2(n12469), .ZN(n13523) );
  INV_X1 U7959 ( .A(n9194), .ZN(n7643) );
  NOR2_X1 U7960 ( .A1(n12524), .A2(n9430), .ZN(n15543) );
  NAND2_X1 U7961 ( .A1(n9177), .A2(n9176), .ZN(n13535) );
  INV_X1 U7962 ( .A(n12457), .ZN(n7392) );
  AND2_X1 U7963 ( .A1(n12458), .A2(n12457), .ZN(n13556) );
  INV_X1 U7964 ( .A(n11811), .ZN(n9123) );
  CLKBUF_X1 U7965 ( .A(n13553), .Z(n13554) );
  NAND2_X1 U7966 ( .A1(n9123), .A2(n7744), .ZN(n7654) );
  AND2_X1 U7967 ( .A1(n7654), .A2(n6504), .ZN(n12114) );
  INV_X1 U7968 ( .A(n15508), .ZN(n15546) );
  AOI21_X1 U7969 ( .B1(n7343), .B2(n9477), .A(n7342), .ZN(n7341) );
  INV_X1 U7970 ( .A(n12444), .ZN(n7342) );
  INV_X1 U7971 ( .A(n7741), .ZN(n6694) );
  AOI21_X1 U7972 ( .B1(n7741), .B2(n6470), .A(n6550), .ZN(n6693) );
  NAND2_X1 U7973 ( .A1(n10854), .A2(n10310), .ZN(n9563) );
  NOR2_X1 U7974 ( .A1(n9511), .A2(n9517), .ZN(n10868) );
  OR2_X1 U7975 ( .A1(n9518), .A2(n9517), .ZN(n10872) );
  NAND2_X1 U7976 ( .A1(n9490), .A2(n12392), .ZN(n15541) );
  AND2_X1 U7977 ( .A1(n8926), .A2(n11906), .ZN(n7666) );
  OAI21_X1 U7978 ( .B1(n12358), .B2(n12357), .A(n12356), .ZN(n12374) );
  NAND2_X1 U7979 ( .A1(n9349), .A2(n11797), .ZN(n7537) );
  NAND2_X1 U7980 ( .A1(n9413), .A2(n7389), .ZN(n9434) );
  NOR2_X1 U7981 ( .A1(n7390), .A2(P3_IR_REG_23__SCAN_IN), .ZN(n7389) );
  XNOR2_X1 U7982 ( .A(n9350), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n9349) );
  AOI21_X1 U7983 ( .B1(n7555), .B2(n7557), .A(n6644), .ZN(n7553) );
  AND2_X1 U7984 ( .A1(n9416), .A2(n9417), .ZN(n9413) );
  NAND2_X1 U7985 ( .A1(n6476), .A2(n6625), .ZN(n7558) );
  AND2_X1 U7986 ( .A1(n6476), .A2(n9271), .ZN(n7559) );
  NAND2_X1 U7987 ( .A1(n9212), .A2(n7550), .ZN(n7549) );
  NOR2_X1 U7988 ( .A1(n9230), .A2(n7551), .ZN(n7550) );
  INV_X1 U7989 ( .A(n9211), .ZN(n7551) );
  NAND3_X1 U7990 ( .A1(n7539), .A2(n7538), .A3(n9179), .ZN(n9196) );
  NAND2_X1 U7991 ( .A1(n9144), .A2(n10466), .ZN(n9161) );
  AND2_X1 U7992 ( .A1(n9145), .A2(n9161), .ZN(n9146) );
  NAND2_X1 U7993 ( .A1(n6844), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n9145) );
  INV_X1 U7994 ( .A(n9144), .ZN(n6844) );
  NAND2_X1 U7995 ( .A1(n6815), .A2(n6814), .ZN(n7545) );
  AOI21_X1 U7996 ( .B1(n6817), .B2(n6819), .A(n6587), .ZN(n6814) );
  INV_X1 U7997 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9105) );
  XNOR2_X1 U7998 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9103) );
  AOI21_X1 U7999 ( .B1(n7529), .B2(n7531), .A(n6583), .ZN(n7527) );
  INV_X1 U8000 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9087) );
  INV_X1 U8001 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9070) );
  XNOR2_X1 U8002 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9085) );
  XNOR2_X1 U8003 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n9068) );
  AND2_X1 U8004 ( .A1(n10275), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9039) );
  XNOR2_X1 U8005 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9021) );
  XNOR2_X1 U8006 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9006) );
  NAND2_X1 U8007 ( .A1(n8975), .A2(n6821), .ZN(n6820) );
  XNOR2_X1 U8008 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8973) );
  NAND2_X1 U8009 ( .A1(n9165), .A2(n8962), .ZN(n7283) );
  NAND2_X1 U8010 ( .A1(n8961), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7284) );
  INV_X1 U8011 ( .A(n7256), .ZN(n7255) );
  OAI21_X1 U8012 ( .B1(n9687), .B2(n7257), .A(n11384), .ZN(n7256) );
  INV_X1 U8013 ( .A(n9689), .ZN(n7257) );
  NAND2_X1 U8014 ( .A1(n7266), .A2(n7265), .ZN(n7264) );
  INV_X1 U8015 ( .A(n9734), .ZN(n7265) );
  NAND2_X1 U8016 ( .A1(n9674), .A2(n11312), .ZN(n11315) );
  OR2_X1 U8017 ( .A1(n8573), .A2(n11994), .ZN(n8582) );
  INV_X1 U8018 ( .A(n11070), .ZN(n11173) );
  AOI21_X1 U8019 ( .B1(n9734), .B2(n9735), .A(n6577), .ZN(n7269) );
  NAND2_X1 U8020 ( .A1(n12599), .A2(n9734), .ZN(n7268) );
  INV_X1 U8021 ( .A(n7187), .ZN(n8774) );
  INV_X1 U8022 ( .A(n13739), .ZN(n7260) );
  AND2_X1 U8023 ( .A1(n8426), .A2(n8425), .ZN(n12830) );
  OR2_X1 U8024 ( .A1(n13941), .A2(n8690), .ZN(n8426) );
  AND2_X1 U8025 ( .A1(n8696), .A2(n8695), .ZN(n12645) );
  AND2_X1 U8026 ( .A1(n8667), .A2(n8666), .ZN(n12719) );
  NAND2_X1 U8027 ( .A1(n7171), .A2(n7169), .ZN(n7168) );
  INV_X1 U8028 ( .A(n10487), .ZN(n7169) );
  NAND2_X1 U8029 ( .A1(n15364), .A2(n7170), .ZN(n7167) );
  OR2_X1 U8030 ( .A1(n10686), .A2(n10685), .ZN(n11136) );
  AND2_X1 U8031 ( .A1(n7155), .A2(n7159), .ZN(n7154) );
  OR2_X1 U8032 ( .A1(n11141), .A2(n7156), .ZN(n7155) );
  NAND2_X1 U8033 ( .A1(n10921), .A2(n7160), .ZN(n7156) );
  NAND2_X1 U8034 ( .A1(n10922), .A2(n6498), .ZN(n7152) );
  INV_X1 U8035 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6967) );
  AND2_X1 U8036 ( .A1(n8801), .A2(n8786), .ZN(n13934) );
  NAND2_X1 U8037 ( .A1(n14126), .A2(n13813), .ZN(n7685) );
  NOR2_X1 U8038 ( .A1(n8867), .A2(n7580), .ZN(n7579) );
  INV_X1 U8039 ( .A(n8864), .ZN(n7580) );
  OR2_X1 U8040 ( .A1(n12867), .A2(n12866), .ZN(n13981) );
  NAND2_X1 U8041 ( .A1(n13985), .A2(n7742), .ZN(n13974) );
  NAND2_X1 U8042 ( .A1(n8408), .A2(n7194), .ZN(n8749) );
  AND2_X1 U8043 ( .A1(n7195), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n7194) );
  OR2_X1 U8044 ( .A1(n8705), .A2(n11975), .ZN(n8714) );
  NAND2_X1 U8045 ( .A1(n7604), .A2(n6564), .ZN(n7603) );
  NAND2_X1 U8046 ( .A1(n6945), .A2(n6948), .ZN(n8850) );
  INV_X1 U8047 ( .A(n6944), .ZN(n6948) );
  NAND2_X1 U8048 ( .A1(n6947), .A2(n6946), .ZN(n6945) );
  NAND2_X1 U8049 ( .A1(n11698), .A2(n6527), .ZN(n7731) );
  AOI21_X1 U8050 ( .B1(n6485), .B2(n7674), .A(n7673), .ZN(n7672) );
  NOR2_X1 U8051 ( .A1(n14212), .A2(n13855), .ZN(n7673) );
  NOR2_X1 U8052 ( .A1(n8604), .A2(n7676), .ZN(n7675) );
  INV_X1 U8053 ( .A(n8591), .ZN(n7676) );
  NAND2_X1 U8054 ( .A1(n8406), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U8055 ( .A1(n7565), .A2(n6933), .ZN(n6932) );
  NAND2_X1 U8056 ( .A1(n15430), .A2(n15429), .ZN(n7573) );
  AND4_X1 U8057 ( .A1(n8508), .A2(n8507), .A3(n8506), .A4(n8505), .ZN(n11191)
         );
  NAND2_X1 U8058 ( .A1(n8440), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8505) );
  INV_X1 U8059 ( .A(n13801), .ZN(n13812) );
  NAND2_X1 U8060 ( .A1(n11173), .A2(n15466), .ZN(n11172) );
  INV_X1 U8061 ( .A(n6994), .ZN(n9784) );
  AND2_X1 U8062 ( .A1(n14099), .A2(n7396), .ZN(n14111) );
  NAND2_X1 U8063 ( .A1(n14100), .A2(n15472), .ZN(n7396) );
  AOI21_X1 U8064 ( .B1(n7678), .B2(n7681), .A(n6586), .ZN(n7677) );
  OR2_X1 U8065 ( .A1(n12965), .A2(n14102), .ZN(n14108) );
  OAI21_X1 U8066 ( .B1(n12151), .B2(n8893), .A(n12351), .ZN(n15449) );
  NAND2_X1 U8067 ( .A1(n14246), .A2(n8895), .ZN(n7066) );
  INV_X1 U8068 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8419) );
  AND2_X1 U8069 ( .A1(n8412), .A2(n8411), .ZN(n8429) );
  OR2_X1 U8070 ( .A1(n8888), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U8071 ( .A1(n8896), .A2(n8897), .ZN(n8888) );
  NAND2_X1 U8072 ( .A1(n11473), .A2(n11474), .ZN(n7612) );
  INV_X1 U8073 ( .A(n14503), .ZN(n6727) );
  INV_X1 U8074 ( .A(n6871), .ZN(n8171) );
  AND2_X1 U8075 ( .A1(n14369), .A2(n14368), .ZN(n14422) );
  INV_X1 U8076 ( .A(n14423), .ZN(n7028) );
  NOR2_X1 U8077 ( .A1(n14422), .A2(n14561), .ZN(n7027) );
  INV_X1 U8078 ( .A(n14372), .ZN(n6713) );
  NOR2_X1 U8079 ( .A1(n7617), .A2(n6713), .ZN(n6711) );
  NAND2_X1 U8080 ( .A1(n14357), .A2(n7615), .ZN(n7029) );
  NOR2_X1 U8081 ( .A1(n7619), .A2(n7616), .ZN(n7615) );
  INV_X1 U8082 ( .A(n14539), .ZN(n7619) );
  NAND2_X1 U8083 ( .A1(n11476), .A2(n7613), .ZN(n7609) );
  AND2_X1 U8084 ( .A1(n7022), .A2(n14474), .ZN(n7021) );
  NAND2_X1 U8085 ( .A1(n14278), .A2(n7016), .ZN(n7022) );
  NAND2_X1 U8086 ( .A1(n7024), .A2(n7016), .ZN(n7023) );
  INV_X1 U8087 ( .A(n7620), .ZN(n7024) );
  AND2_X1 U8088 ( .A1(n14451), .A2(n14344), .ZN(n14483) );
  NAND2_X1 U8089 ( .A1(n10388), .A2(n10471), .ZN(n10473) );
  AOI21_X1 U8090 ( .B1(n6731), .B2(n6715), .A(n6585), .ZN(n6714) );
  INV_X1 U8091 ( .A(n6731), .ZN(n6716) );
  AND2_X1 U8092 ( .A1(n14261), .A2(n14260), .ZN(n14463) );
  AND2_X1 U8093 ( .A1(n9858), .A2(n9857), .ZN(n10028) );
  NAND2_X1 U8094 ( .A1(n7835), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7415) );
  OR2_X1 U8095 ( .A1(n10335), .A2(n10336), .ZN(n10607) );
  NAND2_X1 U8096 ( .A1(n8374), .A2(n11988), .ZN(n7761) );
  NAND2_X1 U8097 ( .A1(n14811), .A2(n8282), .ZN(n14786) );
  INV_X1 U8098 ( .A(n8282), .ZN(n6778) );
  OR2_X1 U8099 ( .A1(n7008), .A2(n11797), .ZN(n8263) );
  NAND2_X1 U8100 ( .A1(n6871), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U8101 ( .A1(n8134), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8155) );
  OAI21_X1 U8102 ( .B1(n7429), .B2(n7430), .A(n8338), .ZN(n7426) );
  AND2_X1 U8103 ( .A1(n14964), .A2(n14955), .ZN(n14953) );
  NOR2_X1 U8104 ( .A1(n15000), .A2(n14981), .ZN(n14964) );
  NAND2_X1 U8105 ( .A1(n11743), .A2(n7715), .ZN(n6784) );
  NAND2_X1 U8106 ( .A1(n7945), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7978) );
  INV_X1 U8107 ( .A(n7947), .ZN(n7945) );
  XNOR2_X1 U8108 ( .A(n11723), .B(n12041), .ZN(n11719) );
  NAND2_X1 U8109 ( .A1(n11456), .A2(n14579), .ZN(n7931) );
  NAND2_X1 U8110 ( .A1(n11291), .A2(n11220), .ZN(n11456) );
  NOR2_X1 U8111 ( .A1(n11465), .A2(n11596), .ZN(n11716) );
  NAND2_X1 U8112 ( .A1(n7832), .A2(n7831), .ZN(n10706) );
  INV_X1 U8113 ( .A(n10073), .ZN(n10707) );
  AND2_X1 U8114 ( .A1(n10390), .A2(n7809), .ZN(n15008) );
  NAND2_X1 U8115 ( .A1(n9878), .A2(n7709), .ZN(n14769) );
  INV_X1 U8116 ( .A(n14955), .ZN(n15099) );
  NAND2_X1 U8117 ( .A1(n8062), .A2(n8061), .ZN(n15112) );
  NAND2_X1 U8118 ( .A1(n8011), .A2(n8010), .ZN(n15117) );
  AND2_X1 U8119 ( .A1(n8382), .A2(n8397), .ZN(n10251) );
  INV_X1 U8120 ( .A(n7479), .ZN(n7478) );
  XNOR2_X1 U8121 ( .A(n10042), .B(n10041), .ZN(n12809) );
  XNOR2_X1 U8122 ( .A(n7777), .B(P1_IR_REG_29__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U8123 ( .A1(n6855), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7777) );
  AND2_X1 U8124 ( .A1(n6459), .A2(n7903), .ZN(n6856) );
  INV_X1 U8125 ( .A(n7792), .ZN(n6776) );
  XNOR2_X1 U8126 ( .A(n8302), .B(n8288), .ZN(n12348) );
  INV_X1 U8127 ( .A(n8259), .ZN(n8258) );
  INV_X1 U8128 ( .A(n8256), .ZN(n8255) );
  INV_X1 U8129 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7762) );
  NOR2_X1 U8130 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n7763) );
  NAND2_X1 U8131 ( .A1(n8129), .A2(n8128), .ZN(n8144) );
  XNOR2_X1 U8132 ( .A(n8101), .B(n8100), .ZN(n10751) );
  AND2_X1 U8133 ( .A1(n8107), .A2(n8130), .ZN(n12087) );
  XNOR2_X1 U8134 ( .A(n6858), .B(n7939), .ZN(n10246) );
  NAND2_X1 U8135 ( .A1(n7937), .A2(n7936), .ZN(n6858) );
  XNOR2_X1 U8136 ( .A(n7907), .B(n7908), .ZN(n10243) );
  XNOR2_X1 U8137 ( .A(n7884), .B(n7883), .ZN(n10238) );
  AND2_X1 U8138 ( .A1(n7296), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10162) );
  NAND2_X1 U8139 ( .A1(n11621), .A2(n11620), .ZN(n6836) );
  NAND2_X1 U8140 ( .A1(n6456), .A2(n6561), .ZN(n7304) );
  INV_X1 U8141 ( .A(n15203), .ZN(n7305) );
  NAND2_X1 U8142 ( .A1(n11500), .A2(n11499), .ZN(n11604) );
  NAND2_X1 U8143 ( .A1(n7364), .A2(n7363), .ZN(n13100) );
  AOI21_X1 U8144 ( .B1(n6449), .B2(n13038), .A(n6584), .ZN(n7363) );
  AND3_X1 U8145 ( .A1(n9193), .A2(n9192), .A3(n9191), .ZN(n13113) );
  AND2_X1 U8146 ( .A1(n7373), .A2(n7374), .ZN(n13119) );
  AOI21_X1 U8147 ( .B1(n7376), .B2(n7380), .A(n6581), .ZN(n7374) );
  OR2_X1 U8148 ( .A1(n13024), .A2(n7375), .ZN(n7373) );
  AOI21_X1 U8149 ( .B1(n13060), .B2(n7358), .A(n6526), .ZN(n7357) );
  INV_X1 U8150 ( .A(n13031), .ZN(n7358) );
  AND2_X1 U8151 ( .A1(n9152), .A2(n9151), .ZN(n12029) );
  OR2_X1 U8152 ( .A1(n10404), .A2(n9149), .ZN(n9152) );
  INV_X1 U8153 ( .A(n13195), .ZN(n13184) );
  NAND2_X1 U8154 ( .A1(n6685), .A2(n15552), .ZN(n6684) );
  INV_X1 U8155 ( .A(n12539), .ZN(n6685) );
  NAND2_X1 U8156 ( .A1(n12577), .A2(n12583), .ZN(n6678) );
  INV_X1 U8157 ( .A(n13429), .ZN(n13457) );
  INV_X1 U8158 ( .A(n13490), .ZN(n13515) );
  INV_X1 U8159 ( .A(n13027), .ZN(n13525) );
  INV_X1 U8160 ( .A(n12028), .ZN(n13559) );
  INV_X1 U8161 ( .A(n13161), .ZN(n13558) );
  OR2_X2 U8162 ( .A1(n10854), .A2(n10270), .ZN(n13214) );
  CLKBUF_X1 U8163 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n6864) );
  NAND2_X1 U8164 ( .A1(n10456), .A2(n9580), .ZN(n7226) );
  NAND2_X1 U8165 ( .A1(n10570), .A2(n7227), .ZN(n7225) );
  AND2_X1 U8166 ( .A1(n7244), .A2(n7085), .ZN(n10780) );
  NAND2_X1 U8167 ( .A1(n7236), .A2(n7235), .ZN(n7104) );
  NAND2_X1 U8168 ( .A1(n7210), .A2(n7216), .ZN(n11412) );
  NAND2_X1 U8169 ( .A1(n10834), .A2(n7211), .ZN(n7210) );
  NAND2_X1 U8170 ( .A1(n13269), .A2(n7200), .ZN(n13271) );
  AND2_X1 U8171 ( .A1(n13267), .A2(n13268), .ZN(n7200) );
  AND2_X1 U8172 ( .A1(n7271), .A2(n9556), .ZN(n7273) );
  INV_X1 U8173 ( .A(n13337), .ZN(n7250) );
  AOI21_X1 U8174 ( .B1(n13338), .B2(n13339), .A(n7249), .ZN(n7248) );
  INV_X1 U8175 ( .A(n13332), .ZN(n7249) );
  NOR2_X1 U8176 ( .A1(n13329), .A2(n13517), .ZN(n13328) );
  XNOR2_X1 U8177 ( .A(n13330), .B(n13604), .ZN(n7251) );
  INV_X1 U8178 ( .A(n13341), .ZN(n13348) );
  INV_X1 U8179 ( .A(n13360), .ZN(n6866) );
  NOR2_X1 U8180 ( .A1(n13343), .A2(n7201), .ZN(n9610) );
  OR2_X1 U8181 ( .A1(n9641), .A2(n9567), .ZN(n13341) );
  NAND2_X1 U8182 ( .A1(n9368), .A2(n9367), .ZN(n13572) );
  NAND2_X1 U8183 ( .A1(n9354), .A2(n9353), .ZN(n13403) );
  NAND2_X1 U8184 ( .A1(n9274), .A2(n9273), .ZN(n13594) );
  NAND2_X1 U8185 ( .A1(n9809), .A2(n9808), .ZN(n13630) );
  OAI21_X1 U8186 ( .B1(n9527), .B2(n13620), .A(n9495), .ZN(n9496) );
  INV_X1 U8187 ( .A(n6669), .ZN(n6668) );
  NOR2_X1 U8188 ( .A1(n15600), .A2(n13628), .ZN(n6923) );
  OAI21_X1 U8189 ( .B1(n9421), .B2(n6800), .A(n6799), .ZN(n6798) );
  OR2_X1 U8190 ( .A1(n9420), .A2(n13472), .ZN(n6800) );
  AND2_X1 U8191 ( .A1(n13575), .A2(n13574), .ZN(n13633) );
  AND2_X1 U8192 ( .A1(n6672), .A2(n15600), .ZN(n6667) );
  NAND2_X1 U8193 ( .A1(n9309), .A2(n9308), .ZN(n13639) );
  NAND2_X1 U8194 ( .A1(n9243), .A2(n9242), .ZN(n13655) );
  NAND2_X1 U8195 ( .A1(n9262), .A2(n9261), .ZN(n13661) );
  NAND2_X1 U8196 ( .A1(n9202), .A2(n9201), .ZN(n13673) );
  NAND2_X1 U8197 ( .A1(n9168), .A2(n9167), .ZN(n13685) );
  NAND2_X1 U8198 ( .A1(n9135), .A2(n9134), .ZN(n12125) );
  OR2_X1 U8199 ( .A1(n10292), .A2(n9149), .ZN(n9135) );
  INV_X1 U8200 ( .A(n13654), .ZN(n13691) );
  OR2_X1 U8201 ( .A1(n15598), .A2(n15541), .ZN(n13654) );
  NAND2_X1 U8202 ( .A1(n9449), .A2(n9448), .ZN(n10268) );
  OR2_X1 U8203 ( .A1(n9447), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9449) );
  INV_X1 U8204 ( .A(n12977), .ZN(n9778) );
  AND2_X1 U8205 ( .A1(n13011), .A2(n9721), .ZN(n6992) );
  NAND2_X1 U8206 ( .A1(n6997), .A2(n13822), .ZN(n6996) );
  INV_X1 U8207 ( .A(n13755), .ZN(n6997) );
  XNOR2_X1 U8208 ( .A(n13728), .B(n13727), .ZN(n13730) );
  NAND2_X1 U8209 ( .A1(n13016), .A2(n9725), .ZN(n12599) );
  NAND2_X1 U8210 ( .A1(n12651), .A2(n9748), .ZN(n13770) );
  OR2_X1 U8211 ( .A1(n11382), .A2(n8757), .ZN(n8713) );
  XNOR2_X1 U8212 ( .A(n13726), .B(n13724), .ZN(n13792) );
  AND2_X1 U8213 ( .A1(n9789), .A2(n9788), .ZN(n13826) );
  NOR2_X1 U8214 ( .A1(n15327), .A2(n11066), .ZN(n13821) );
  NAND2_X1 U8215 ( .A1(n8644), .A2(n8643), .ZN(n13831) );
  INV_X1 U8216 ( .A(n12830), .ZN(n13840) );
  NAND2_X1 U8217 ( .A1(n8768), .A2(n8767), .ZN(n13842) );
  NAND2_X1 U8218 ( .A1(n8756), .A2(n8755), .ZN(n13843) );
  OR2_X1 U8219 ( .A1(n13721), .A2(n8690), .ZN(n8756) );
  OR2_X1 U8220 ( .A1(n8690), .A2(n11067), .ZN(n8442) );
  INV_X1 U8221 ( .A(n6738), .ZN(n8443) );
  NAND2_X1 U8222 ( .A1(n15364), .A2(n15365), .ZN(n15363) );
  NAND2_X1 U8223 ( .A1(n10683), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7160) );
  OR2_X1 U8224 ( .A1(n10922), .A2(n10921), .ZN(n7153) );
  OR2_X1 U8225 ( .A1(n10422), .A2(n12903), .ZN(n15392) );
  NAND2_X1 U8226 ( .A1(n6849), .A2(n6847), .ZN(n7174) );
  INV_X1 U8227 ( .A(n6848), .ZN(n6847) );
  NAND2_X1 U8228 ( .A1(n13915), .A2(n15423), .ZN(n6849) );
  OAI21_X1 U8229 ( .B1(n13914), .B2(n15392), .A(n15408), .ZN(n6848) );
  OAI21_X1 U8230 ( .B1(n15427), .B2(n6967), .A(n13918), .ZN(n7173) );
  NAND2_X1 U8231 ( .A1(n12962), .A2(n12961), .ZN(n12963) );
  NAND2_X1 U8232 ( .A1(n6949), .A2(n15479), .ZN(n6957) );
  INV_X1 U8233 ( .A(n13931), .ZN(n6949) );
  OR2_X1 U8234 ( .A1(n6438), .A2(n11171), .ZN(n15437) );
  INV_X1 U8235 ( .A(n14089), .ZN(n15445) );
  NAND2_X1 U8236 ( .A1(n12149), .A2(n11177), .ZN(n15446) );
  NAND2_X1 U8237 ( .A1(n9785), .A2(n15459), .ZN(n15434) );
  INV_X1 U8238 ( .A(n9792), .ZN(n9785) );
  NOR2_X1 U8239 ( .A1(n6953), .A2(n6626), .ZN(n6952) );
  NOR2_X1 U8240 ( .A1(n6955), .A2(n6954), .ZN(n6953) );
  INV_X1 U8241 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6959) );
  INV_X1 U8242 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11383) );
  AND2_X1 U8243 ( .A1(n8397), .A2(n11796), .ZN(n6737) );
  INV_X1 U8244 ( .A(n12154), .ZN(n6736) );
  AOI21_X1 U8245 ( .B1(n11476), .B2(n11475), .A(n7610), .ZN(n11657) );
  INV_X1 U8246 ( .A(n7612), .ZN(n7610) );
  AND4_X1 U8247 ( .A1(n8050), .A2(n8049), .A3(n8048), .A4(n8047), .ZN(n14386)
         );
  INV_X1 U8248 ( .A(n14981), .ZN(n15105) );
  NAND2_X1 U8249 ( .A1(n11023), .A2(n6734), .ZN(n6733) );
  INV_X1 U8250 ( .A(n14833), .ZN(n15057) );
  OR2_X1 U8251 ( .A1(n7868), .A2(n7867), .ZN(n7869) );
  OR2_X1 U8252 ( .A1(n7608), .A2(n12035), .ZN(n7605) );
  AOI21_X1 U8253 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(n6772) );
  AND2_X1 U8254 ( .A1(n10141), .A2(n10140), .ZN(n7107) );
  NAND2_X1 U8255 ( .A1(n8233), .A2(n8232), .ZN(n14879) );
  NAND2_X1 U8256 ( .A1(n8185), .A2(n8184), .ZN(n14901) );
  INV_X1 U8257 ( .A(n14386), .ZN(n15011) );
  AND2_X1 U8258 ( .A1(n7690), .A2(n7689), .ZN(n15034) );
  OR2_X1 U8259 ( .A1(n7008), .A2(n12945), .ZN(n9840) );
  XNOR2_X1 U8260 ( .A(n14758), .B(n14770), .ZN(n14761) );
  MUX2_X1 U8261 ( .A(n8358), .B(n8357), .S(n10090), .Z(n8370) );
  OR2_X1 U8262 ( .A1(n14793), .A2(n14792), .ZN(n15046) );
  NAND2_X1 U8263 ( .A1(n14851), .A2(n8250), .ZN(n14825) );
  OR2_X1 U8264 ( .A1(n7008), .A2(n11736), .ZN(n8238) );
  OR2_X1 U8265 ( .A1(n7008), .A2(n11380), .ZN(n8210) );
  NOR3_X1 U8266 ( .A1(n11723), .A2(n11465), .A3(n11596), .ZN(n11748) );
  NAND2_X1 U8267 ( .A1(n15305), .A2(n9864), .ZN(n15279) );
  AND2_X1 U8268 ( .A1(n15305), .A2(n8398), .ZN(n15273) );
  INV_X1 U8269 ( .A(n15320), .ZN(n6896) );
  INV_X1 U8270 ( .A(n11291), .ZN(n11429) );
  OR2_X1 U8271 ( .A1(n7868), .A2(n10250), .ZN(n7848) );
  OR2_X1 U8272 ( .A1(n7008), .A2(n15166), .ZN(n8303) );
  AND3_X2 U8273 ( .A1(n7802), .A2(n7801), .A3(n7800), .ZN(n15292) );
  NAND2_X1 U8274 ( .A1(n15319), .A2(n15311), .ZN(n15143) );
  INV_X1 U8275 ( .A(n15296), .ZN(n8398) );
  NAND2_X1 U8276 ( .A1(n10308), .A2(n10307), .ZN(n6832) );
  NAND2_X1 U8277 ( .A1(n6832), .A2(n10309), .ZN(n7310) );
  NAND2_X1 U8278 ( .A1(n11630), .A2(n11629), .ZN(n11849) );
  NAND2_X1 U8279 ( .A1(n6833), .A2(n11627), .ZN(n11848) );
  INV_X1 U8280 ( .A(n6836), .ZN(n6833) );
  NAND2_X1 U8281 ( .A1(n6836), .A2(n11628), .ZN(n11630) );
  XNOR2_X1 U8282 ( .A(n15178), .B(n15176), .ZN(n15175) );
  NOR2_X1 U8283 ( .A1(n15204), .A2(n15203), .ZN(n15208) );
  NOR2_X1 U8284 ( .A1(n6450), .A2(n15203), .ZN(n7306) );
  AND3_X1 U8285 ( .A1(n15241), .A2(n15244), .A3(n15428), .ZN(n15246) );
  INV_X1 U8286 ( .A(n9924), .ZN(n9898) );
  OAI21_X1 U8287 ( .B1(n7076), .B2(n7071), .A(n7069), .ZN(n12695) );
  AOI21_X1 U8288 ( .B1(n7073), .B2(n7078), .A(n7070), .ZN(n7069) );
  INV_X1 U8289 ( .A(n7073), .ZN(n7071) );
  AOI21_X1 U8290 ( .B1(n7447), .B2(n7446), .A(n7444), .ZN(n7443) );
  NAND2_X1 U8291 ( .A1(n7075), .A2(n7072), .ZN(n12689) );
  NOR2_X1 U8292 ( .A1(n7056), .A2(n12701), .ZN(n7455) );
  NOR2_X1 U8293 ( .A1(n7047), .A2(n7050), .ZN(n7046) );
  INV_X1 U8294 ( .A(n12704), .ZN(n7050) );
  NOR2_X1 U8295 ( .A1(n7051), .A2(n7055), .ZN(n7047) );
  OAI21_X1 U8296 ( .B1(n12702), .B2(n7455), .A(n7048), .ZN(n7053) );
  NOR2_X1 U8297 ( .A1(n7049), .A2(n12705), .ZN(n7048) );
  INV_X1 U8298 ( .A(n7055), .ZN(n7049) );
  NAND2_X1 U8299 ( .A1(n9932), .A2(n9931), .ZN(n9934) );
  OAI21_X1 U8300 ( .B1(n9926), .B2(n7128), .A(n6881), .ZN(n9931) );
  NOR2_X1 U8301 ( .A1(n6882), .A2(n9930), .ZN(n6881) );
  NAND2_X1 U8302 ( .A1(n7516), .A2(n9933), .ZN(n7515) );
  NOR2_X1 U8303 ( .A1(n7516), .A2(n9933), .ZN(n7517) );
  INV_X1 U8304 ( .A(n9934), .ZN(n6840) );
  NAND2_X1 U8305 ( .A1(n7184), .A2(n12529), .ZN(n6853) );
  NOR2_X1 U8306 ( .A1(n6454), .A2(n7040), .ZN(n7039) );
  INV_X1 U8307 ( .A(n12712), .ZN(n7040) );
  NOR2_X1 U8308 ( .A1(n6454), .A2(n12715), .ZN(n7037) );
  NAND2_X1 U8309 ( .A1(n9939), .A2(n7511), .ZN(n7510) );
  INV_X1 U8310 ( .A(n12781), .ZN(n7450) );
  INV_X1 U8311 ( .A(n9993), .ZN(n7116) );
  NAND2_X1 U8312 ( .A1(n12790), .A2(n7045), .ZN(n7044) );
  INV_X1 U8313 ( .A(n7114), .ZN(n7110) );
  NOR2_X1 U8314 ( .A1(n7114), .A2(n7112), .ZN(n7111) );
  INV_X1 U8315 ( .A(n10007), .ZN(n7122) );
  OAI21_X1 U8316 ( .B1(n13000), .B2(n6436), .A(n7137), .ZN(n12841) );
  NAND2_X1 U8317 ( .A1(n12828), .A2(n6436), .ZN(n7137) );
  OR2_X1 U8318 ( .A1(n8371), .A2(n15296), .ZN(n9884) );
  NOR2_X1 U8319 ( .A1(n7422), .A2(n11719), .ZN(n7421) );
  INV_X1 U8320 ( .A(n8326), .ZN(n7422) );
  NOR2_X1 U8321 ( .A1(n6928), .A2(n9394), .ZN(n6927) );
  INV_X1 U8322 ( .A(n12519), .ZN(n6928) );
  AND2_X1 U8323 ( .A1(n6604), .A2(n9378), .ZN(n6802) );
  AND2_X1 U8324 ( .A1(n13673), .A2(n13192), .ZN(n12465) );
  MUX2_X1 U8325 ( .A(n13837), .B(n14100), .S(n12728), .Z(n12838) );
  INV_X1 U8326 ( .A(n6564), .ZN(n7600) );
  INV_X1 U8327 ( .A(n8851), .ZN(n7593) );
  OR4_X1 U8328 ( .A1(n12075), .A2(n10078), .A3(n12098), .A4(n11719), .ZN(
        n10079) );
  NOR2_X1 U8329 ( .A1(n6904), .A2(n6903), .ZN(n6902) );
  NAND2_X1 U8330 ( .A1(n15020), .A2(n10081), .ZN(n6904) );
  NAND2_X1 U8331 ( .A1(n8337), .A2(n14948), .ZN(n6903) );
  NAND2_X1 U8332 ( .A1(n10010), .A2(n10013), .ZN(n7508) );
  AOI21_X1 U8333 ( .B1(n7120), .B2(n7520), .A(n6473), .ZN(n7118) );
  NOR2_X1 U8334 ( .A1(n10006), .A2(n10003), .ZN(n7520) );
  NOR2_X1 U8335 ( .A1(n10013), .A2(n10010), .ZN(n7509) );
  NAND2_X1 U8336 ( .A1(n8315), .A2(n9893), .ZN(n9892) );
  INV_X1 U8337 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n11953) );
  INV_X1 U8338 ( .A(n8128), .ZN(n7463) );
  INV_X1 U8339 ( .A(n6759), .ZN(n6758) );
  NAND2_X1 U8340 ( .A1(n6978), .A2(n8054), .ZN(n6761) );
  NAND2_X1 U8341 ( .A1(n6439), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7901) );
  AND2_X1 U8342 ( .A1(n7893), .A2(n7456), .ZN(n6857) );
  OAI22_X1 U8343 ( .A1(n10202), .A2(n6535), .B1(n7314), .B2(
        P3_ADDR_REG_3__SCAN_IN), .ZN(n10205) );
  NAND2_X1 U8344 ( .A1(n13180), .A2(n7331), .ZN(n7330) );
  OR2_X1 U8345 ( .A1(n13407), .A2(n12386), .ZN(n12544) );
  OAI21_X1 U8346 ( .B1(n13714), .B2(P3_REG2_REG_1__SCAN_IN), .A(n7199), .ZN(
        n7198) );
  NAND2_X1 U8347 ( .A1(n13714), .A2(n10627), .ZN(n7199) );
  NAND2_X1 U8348 ( .A1(n7198), .A2(n9568), .ZN(n9571) );
  NOR2_X1 U8349 ( .A1(n10942), .A2(n9550), .ZN(n9551) );
  INV_X1 U8350 ( .A(n6490), .ZN(n7215) );
  NAND2_X1 U8351 ( .A1(n13307), .A2(n9633), .ZN(n9635) );
  AND2_X1 U8352 ( .A1(n9830), .A2(n9401), .ZN(n9505) );
  OR2_X1 U8353 ( .A1(n13374), .A2(n13387), .ZN(n12520) );
  OR2_X1 U8354 ( .A1(n13577), .A2(n13428), .ZN(n12500) );
  NOR2_X1 U8355 ( .A1(n9263), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n6912) );
  NOR2_X1 U8356 ( .A1(n9095), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n6706) );
  INV_X1 U8357 ( .A(n15506), .ZN(n15504) );
  INV_X1 U8358 ( .A(n11673), .ZN(n12428) );
  NAND2_X1 U8359 ( .A1(n11252), .A2(n9011), .ZN(n11448) );
  INV_X1 U8360 ( .A(n15528), .ZN(n12400) );
  OR2_X1 U8361 ( .A1(n9447), .A2(n9459), .ZN(n9510) );
  NAND2_X1 U8362 ( .A1(n12542), .A2(n6696), .ZN(n7347) );
  NAND2_X1 U8363 ( .A1(n6803), .A2(n6801), .ZN(n10144) );
  NAND2_X1 U8364 ( .A1(n7662), .A2(n9378), .ZN(n6803) );
  NAND2_X1 U8365 ( .A1(n9347), .A2(n6802), .ZN(n6801) );
  OAI21_X1 U8366 ( .B1(n6497), .B2(n7663), .A(n9377), .ZN(n7662) );
  OR2_X1 U8367 ( .A1(n13685), .A2(n12028), .ZN(n12388) );
  INV_X1 U8368 ( .A(n12582), .ZN(n9490) );
  INV_X1 U8369 ( .A(n9364), .ZN(n7535) );
  INV_X1 U8370 ( .A(n7558), .ZN(n7557) );
  INV_X1 U8371 ( .A(n7556), .ZN(n7555) );
  OAI21_X1 U8372 ( .B1(n7559), .B2(n7557), .A(n9319), .ZN(n7556) );
  NOR2_X1 U8373 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n6686) );
  INV_X1 U8374 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9181) );
  AOI21_X1 U8375 ( .B1(n9161), .B2(n7541), .A(n6633), .ZN(n7540) );
  INV_X1 U8376 ( .A(n9161), .ZN(n7542) );
  INV_X1 U8377 ( .A(n9106), .ZN(n7546) );
  AND2_X1 U8378 ( .A1(n10314), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9125) );
  INV_X1 U8379 ( .A(n8973), .ZN(n6821) );
  AND2_X1 U8380 ( .A1(n8938), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8963) );
  INV_X1 U8381 ( .A(n8514), .ZN(n7189) );
  OR4_X1 U8382 ( .A1(n12882), .A2(n12881), .A3(n12880), .A4(n12879), .ZN(
        n12883) );
  AND2_X1 U8383 ( .A1(n12874), .A2(n6515), .ZN(n12877) );
  OAI21_X1 U8384 ( .B1(n7057), .B2(n6499), .A(n7058), .ZN(n12806) );
  NAND2_X1 U8385 ( .A1(n12802), .A2(n12804), .ZN(n7058) );
  INV_X1 U8386 ( .A(n13838), .ZN(n12828) );
  NOR2_X1 U8387 ( .A1(n13970), .A2(n14119), .ZN(n7409) );
  NAND2_X1 U8388 ( .A1(n7412), .A2(n14126), .ZN(n7411) );
  INV_X1 U8389 ( .A(n8866), .ZN(n7578) );
  NOR2_X1 U8390 ( .A1(n7197), .A2(n7196), .ZN(n7195) );
  INV_X1 U8391 ( .A(n8714), .ZN(n8408) );
  NOR2_X1 U8392 ( .A1(n8660), .A2(n8645), .ZN(n7190) );
  INV_X1 U8393 ( .A(n8646), .ZN(n8407) );
  NAND2_X1 U8394 ( .A1(n8847), .A2(n12886), .ZN(n6944) );
  INV_X1 U8395 ( .A(n11869), .ZN(n6947) );
  NOR2_X1 U8396 ( .A1(n12733), .A2(n7405), .ZN(n7404) );
  INV_X1 U8397 ( .A(n7406), .ZN(n7405) );
  NOR2_X1 U8398 ( .A1(n11270), .A2(n7192), .ZN(n7191) );
  INV_X1 U8399 ( .A(n8582), .ZN(n8406) );
  NOR2_X1 U8400 ( .A1(n12711), .A2(n14212), .ZN(n7406) );
  INV_X1 U8401 ( .A(n8839), .ZN(n6933) );
  INV_X1 U8402 ( .A(n7568), .ZN(n7567) );
  NOR2_X1 U8403 ( .A1(n7571), .A2(n8842), .ZN(n7570) );
  INV_X1 U8404 ( .A(n8840), .ZN(n7571) );
  NAND2_X1 U8405 ( .A1(n13859), .A2(n11582), .ZN(n7568) );
  NAND2_X1 U8406 ( .A1(n11346), .A2(n8839), .ZN(n8841) );
  NAND2_X1 U8407 ( .A1(n11404), .A2(n12906), .ZN(n6994) );
  NOR2_X1 U8408 ( .A1(n14081), .A2(n7401), .ZN(n14047) );
  NAND2_X1 U8409 ( .A1(n8841), .A2(n8840), .ZN(n11566) );
  NAND2_X1 U8410 ( .A1(n6931), .A2(n8837), .ZN(n11239) );
  NOR2_X1 U8411 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6741) );
  NOR2_X1 U8412 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6742) );
  NOR2_X1 U8413 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6743) );
  NOR2_X1 U8414 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6744) );
  INV_X1 U8415 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8415) );
  INV_X1 U8416 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8414) );
  INV_X1 U8417 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8413) );
  INV_X1 U8418 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n11996) );
  INV_X1 U8419 ( .A(n14302), .ZN(n6728) );
  AND2_X1 U8420 ( .A1(n14367), .A2(n14366), .ZN(n14368) );
  XNOR2_X1 U8421 ( .A(n6721), .B(n11660), .ZN(n10788) );
  NAND2_X1 U8422 ( .A1(n10531), .A2(n10532), .ZN(n6721) );
  INV_X1 U8423 ( .A(n14265), .ZN(n6715) );
  NAND2_X1 U8424 ( .A1(n7497), .A2(n7496), .ZN(n10127) );
  INV_X1 U8425 ( .A(n10107), .ZN(n7497) );
  INV_X1 U8426 ( .A(n10106), .ZN(n7496) );
  NAND2_X1 U8427 ( .A1(n7501), .A2(n7500), .ZN(n10105) );
  NAND2_X1 U8428 ( .A1(n10096), .A2(n10095), .ZN(n7500) );
  NAND2_X1 U8429 ( .A1(n10124), .A2(n10127), .ZN(n10116) );
  INV_X1 U8430 ( .A(n8220), .ZN(n7722) );
  AND2_X1 U8431 ( .A1(n6513), .A2(n14867), .ZN(n7693) );
  INV_X1 U8432 ( .A(n9965), .ZN(n6787) );
  NOR2_X1 U8433 ( .A1(n8110), .A2(n6870), .ZN(n8134) );
  NAND2_X1 U8434 ( .A1(n14989), .A2(n8115), .ZN(n8117) );
  NOR2_X1 U8435 ( .A1(n15112), .A2(n14573), .ZN(n8115) );
  NAND2_X1 U8436 ( .A1(n8088), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8110) );
  INV_X1 U8437 ( .A(n8090), .ZN(n8088) );
  OR2_X1 U8438 ( .A1(n15107), .A2(n14966), .ZN(n9977) );
  INV_X1 U8439 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8064) );
  OR2_X1 U8440 ( .A1(n8065), .A2(n8064), .ZN(n8090) );
  NOR2_X1 U8441 ( .A1(n15112), .A2(n7695), .ZN(n7694) );
  INV_X1 U8442 ( .A(n7696), .ZN(n7695) );
  NOR2_X1 U8443 ( .A1(n12236), .A2(n12205), .ZN(n7696) );
  OAI21_X1 U8444 ( .B1(n11460), .B2(n7420), .A(n7418), .ZN(n11738) );
  NOR2_X1 U8445 ( .A1(n11723), .A2(n7699), .ZN(n7697) );
  NAND2_X1 U8446 ( .A1(n11747), .A2(n7700), .ZN(n7699) );
  INV_X1 U8447 ( .A(n10075), .ZN(n11099) );
  AND2_X1 U8448 ( .A1(n14918), .A2(n15082), .ZN(n14907) );
  INV_X1 U8449 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7015) );
  AND2_X1 U8450 ( .A1(n7482), .A2(n7481), .ZN(n7480) );
  OR2_X1 U8451 ( .A1(n10058), .A2(n10059), .ZN(n7481) );
  NAND2_X1 U8452 ( .A1(n7486), .A2(n7483), .ZN(n7482) );
  NAND2_X1 U8453 ( .A1(n7486), .A2(n7485), .ZN(n7484) );
  INV_X1 U8454 ( .A(n7489), .ZN(n7485) );
  AOI21_X1 U8455 ( .B1(n7466), .B2(n6465), .A(n6630), .ZN(n7465) );
  NAND2_X1 U8456 ( .A1(n6965), .A2(n6962), .ZN(n7790) );
  NAND4_X1 U8457 ( .A1(n6964), .A2(n6963), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6962) );
  INV_X1 U8458 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U8459 ( .A1(n8194), .A2(SI_21_), .ZN(n8222) );
  INV_X1 U8460 ( .A(n6766), .ZN(n6765) );
  OAI21_X1 U8461 ( .B1(n7460), .B2(n6488), .A(n8197), .ZN(n6766) );
  NAND2_X1 U8462 ( .A1(n7139), .A2(n6558), .ZN(n7138) );
  INV_X1 U8463 ( .A(n8119), .ZN(n7139) );
  OR2_X1 U8464 ( .A1(n8024), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8025) );
  NAND2_X1 U8465 ( .A1(n7470), .A2(n7471), .ZN(n7469) );
  OAI21_X1 U8466 ( .B1(n6439), .B2(n7817), .A(n7816), .ZN(n7839) );
  NAND2_X1 U8467 ( .A1(n6439), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U8468 ( .A1(n10206), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10295) );
  INV_X1 U8469 ( .A(n10205), .ZN(n10206) );
  AOI21_X1 U8470 ( .B1(n10970), .B2(n10969), .A(n10968), .ZN(n10972) );
  OAI21_X1 U8471 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n11625), .A(n11624), .ZN(
        n11850) );
  NAND2_X1 U8472 ( .A1(n12336), .A2(n12335), .ZN(n15182) );
  OR2_X1 U8473 ( .A1(n12334), .A2(n12333), .ZN(n12336) );
  NAND2_X1 U8474 ( .A1(n6831), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n6830) );
  AND2_X1 U8475 ( .A1(n7304), .A2(n6830), .ZN(n6828) );
  OR2_X1 U8476 ( .A1(n15228), .A2(n15227), .ZN(n15229) );
  NAND2_X1 U8477 ( .A1(n13046), .A2(n13045), .ZN(n7331) );
  INV_X1 U8478 ( .A(n7327), .ZN(n7324) );
  XNOR2_X1 U8479 ( .A(n13072), .B(n13071), .ZN(n13073) );
  NAND2_X1 U8480 ( .A1(n7321), .A2(n7326), .ZN(n7320) );
  NAND2_X1 U8481 ( .A1(n13073), .A2(n7329), .ZN(n7326) );
  INV_X1 U8482 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10944) );
  NAND2_X1 U8483 ( .A1(n12020), .A2(n12019), .ZN(n12173) );
  AND2_X1 U8484 ( .A1(n7378), .A2(n6601), .ZN(n7376) );
  NAND2_X1 U8485 ( .A1(n7366), .A2(n7370), .ZN(n13126) );
  NAND2_X1 U8486 ( .A1(n7368), .A2(n7367), .ZN(n7366) );
  INV_X1 U8487 ( .A(n13137), .ZN(n7368) );
  NAND3_X1 U8488 ( .A1(n11075), .A2(n11079), .A3(n7349), .ZN(n11181) );
  AND2_X1 U8489 ( .A1(n11180), .A2(n11074), .ZN(n7349) );
  NOR2_X1 U8490 ( .A1(n7359), .A2(n7356), .ZN(n7355) );
  INV_X1 U8491 ( .A(n13171), .ZN(n7356) );
  INV_X1 U8492 ( .A(n13060), .ZN(n7359) );
  AND2_X1 U8493 ( .A1(n6912), .A2(n6707), .ZN(n9276) );
  INV_X1 U8494 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n6707) );
  AOI21_X1 U8495 ( .B1(n10879), .B2(P3_D_REG_0__SCAN_IN), .A(n7362), .ZN(n7361) );
  INV_X1 U8496 ( .A(n10881), .ZN(n7362) );
  AND4_X1 U8497 ( .A1(n12371), .A2(n12370), .A3(n12369), .A4(n12368), .ZN(
        n13363) );
  OR2_X1 U8498 ( .A1(n9425), .A2(n9830), .ZN(n12371) );
  NAND2_X1 U8499 ( .A1(n6444), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8960) );
  OR2_X1 U8500 ( .A1(n9425), .A2(n15554), .ZN(n8936) );
  OR2_X1 U8501 ( .A1(n12365), .A2(n15558), .ZN(n8934) );
  OR2_X1 U8502 ( .A1(n12366), .A2(n10627), .ZN(n8937) );
  OAI21_X1 U8503 ( .B1(n7198), .B2(n9568), .A(n9571), .ZN(n10621) );
  AOI21_X1 U8504 ( .B1(n10628), .B2(P3_REG1_REG_1__SCAN_IN), .A(n9617), .ZN(
        n10567) );
  INV_X1 U8505 ( .A(n7093), .ZN(n10566) );
  OAI211_X1 U8506 ( .C1(n10451), .C2(n7086), .A(n7083), .B(n7082), .ZN(n7246)
         );
  INV_X1 U8507 ( .A(n10781), .ZN(n7083) );
  OR2_X1 U8508 ( .A1(n7084), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7082) );
  NAND2_X1 U8509 ( .A1(n10451), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7244) );
  AND2_X1 U8510 ( .A1(n9541), .A2(n9542), .ZN(n7285) );
  XNOR2_X1 U8511 ( .A(n9619), .B(n10746), .ZN(n10741) );
  NAND2_X1 U8512 ( .A1(n9540), .A2(n10746), .ZN(n9542) );
  AND2_X1 U8513 ( .A1(n7098), .A2(n6522), .ZN(n9621) );
  NOR2_X1 U8514 ( .A1(n10836), .A2(n10837), .ZN(n10835) );
  OAI21_X1 U8515 ( .B1(n10836), .B2(n7287), .A(n7286), .ZN(n10942) );
  NAND2_X1 U8516 ( .A1(n7288), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7287) );
  NAND2_X1 U8517 ( .A1(n9548), .A2(n7288), .ZN(n7286) );
  INV_X1 U8518 ( .A(n10943), .ZN(n7288) );
  NOR2_X1 U8519 ( .A1(n7215), .A2(n7217), .ZN(n7211) );
  OR2_X1 U8520 ( .A1(n7218), .A2(n7217), .ZN(n7216) );
  INV_X1 U8521 ( .A(n10940), .ZN(n7219) );
  NOR2_X1 U8522 ( .A1(n9553), .A2(n7281), .ZN(n13225) );
  NOR2_X1 U8523 ( .A1(n11413), .A2(n11307), .ZN(n7275) );
  NAND2_X1 U8524 ( .A1(n7278), .A2(n9624), .ZN(n7274) );
  NAND2_X1 U8525 ( .A1(n13225), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n13232) );
  AND2_X1 U8526 ( .A1(n10291), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7295) );
  INV_X1 U8527 ( .A(n7293), .ZN(n13275) );
  NAND2_X1 U8528 ( .A1(n13279), .A2(n13280), .ZN(n13278) );
  NAND2_X1 U8529 ( .A1(n13261), .A2(n9629), .ZN(n13279) );
  XNOR2_X1 U8530 ( .A(n9631), .B(n13304), .ZN(n13292) );
  OR2_X1 U8531 ( .A1(n13300), .A2(n13299), .ZN(n7234) );
  NAND2_X1 U8532 ( .A1(n9605), .A2(n13304), .ZN(n7233) );
  INV_X1 U8533 ( .A(n7080), .ZN(n7079) );
  OAI21_X1 U8534 ( .B1(n9629), .B2(n7081), .A(n9630), .ZN(n7080) );
  INV_X1 U8535 ( .A(n13280), .ZN(n7081) );
  OR2_X1 U8536 ( .A1(n13334), .A2(n7203), .ZN(n7202) );
  NOR2_X1 U8537 ( .A1(n7204), .A2(n13338), .ZN(n7203) );
  AOI21_X1 U8538 ( .B1(n7175), .B2(n6697), .A(n6696), .ZN(n6695) );
  INV_X1 U8539 ( .A(n7175), .ZN(n6698) );
  INV_X1 U8540 ( .A(n7176), .ZN(n6697) );
  NAND2_X1 U8541 ( .A1(n9647), .A2(n9363), .ZN(n13390) );
  INV_X1 U8542 ( .A(n12510), .ZN(n12566) );
  INV_X1 U8543 ( .A(n9347), .ZN(n13413) );
  OR2_X1 U8544 ( .A1(n9310), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9322) );
  AND2_X1 U8545 ( .A1(n9276), .A2(n9275), .ZN(n9292) );
  NAND2_X1 U8546 ( .A1(n9292), .A2(n9291), .ZN(n9310) );
  INV_X1 U8547 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13120) );
  NAND2_X1 U8548 ( .A1(n9219), .A2(n13120), .ZN(n9263) );
  AND2_X1 U8549 ( .A1(n9203), .A2(n13110), .ZN(n9219) );
  INV_X1 U8550 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9153) );
  NAND2_X1 U8551 ( .A1(n9154), .A2(n9153), .ZN(n9171) );
  NAND2_X1 U8552 ( .A1(n6706), .A2(n6705), .ZN(n9136) );
  INV_X1 U8553 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U8554 ( .A1(n9077), .A2(n9076), .ZN(n9095) );
  INV_X1 U8555 ( .A(n6706), .ZN(n9116) );
  AND2_X1 U8556 ( .A1(n12439), .A2(n12440), .ZN(n15506) );
  AND4_X1 U8557 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(n15509)
         );
  INV_X1 U8558 ( .A(n12555), .ZN(n11785) );
  OR2_X1 U8559 ( .A1(n11448), .A2(n12552), .ZN(n11676) );
  NAND2_X1 U8560 ( .A1(n6704), .A2(n6929), .ZN(n9031) );
  INV_X1 U8561 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n6929) );
  INV_X1 U8562 ( .A(n9013), .ZN(n6704) );
  NAND2_X1 U8563 ( .A1(n11325), .A2(n9473), .ZN(n7332) );
  OR2_X1 U8564 ( .A1(n12551), .A2(n12414), .ZN(n7333) );
  NOR2_X2 U8565 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8996) );
  NAND2_X1 U8566 ( .A1(n9024), .A2(n10580), .ZN(n6701) );
  OAI22_X1 U8567 ( .A1(n10181), .A2(n9149), .B1(n12376), .B2(SI_2_), .ZN(n6666) );
  INV_X1 U8568 ( .A(n12393), .ZN(n15542) );
  AND2_X1 U8569 ( .A1(n12527), .A2(n9810), .ZN(n12570) );
  NAND2_X1 U8570 ( .A1(n12568), .A2(n10147), .ZN(n6799) );
  AND2_X1 U8571 ( .A1(n12502), .A2(n12497), .ZN(n13443) );
  AOI21_X1 U8572 ( .B1(n7180), .B2(n7182), .A(n7178), .ZN(n7177) );
  NAND2_X1 U8573 ( .A1(n7352), .A2(n7180), .ZN(n7179) );
  INV_X1 U8574 ( .A(n12493), .ZN(n7178) );
  INV_X1 U8575 ( .A(n15541), .ZN(n13595) );
  AND2_X1 U8576 ( .A1(n9270), .A2(n9269), .ZN(n13490) );
  NAND2_X1 U8577 ( .A1(n6655), .A2(n7641), .ZN(n6654) );
  AND2_X1 U8578 ( .A1(n13521), .A2(n7642), .ZN(n7641) );
  NAND2_X1 U8579 ( .A1(n6664), .A2(n7183), .ZN(n13532) );
  AOI21_X1 U8580 ( .B1(n6457), .B2(n7392), .A(n7184), .ZN(n7183) );
  NAND2_X1 U8581 ( .A1(n13532), .A2(n13534), .ZN(n13531) );
  INV_X1 U8582 ( .A(n7649), .ZN(n7001) );
  AOI21_X1 U8583 ( .B1(n7338), .B2(n7339), .A(n7335), .ZN(n7334) );
  NAND2_X1 U8584 ( .A1(n15505), .A2(n7338), .ZN(n7336) );
  INV_X1 U8585 ( .A(n12443), .ZN(n7335) );
  AND2_X1 U8586 ( .A1(n10853), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10310) );
  NAND2_X1 U8587 ( .A1(n7394), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8931) );
  AND2_X1 U8588 ( .A1(n9438), .A2(n7666), .ZN(n7393) );
  NOR2_X1 U8589 ( .A1(n9395), .A2(n7563), .ZN(n7562) );
  INV_X1 U8590 ( .A(n9381), .ZN(n7563) );
  OR2_X1 U8591 ( .A1(n8927), .A2(n6677), .ZN(n6676) );
  NAND2_X1 U8592 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), 
        .ZN(n6677) );
  INV_X1 U8593 ( .A(n7390), .ZN(n7388) );
  AND2_X1 U8594 ( .A1(n9238), .A2(n9237), .ZN(n9254) );
  OR2_X1 U8595 ( .A1(n9088), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9109) );
  AND2_X1 U8596 ( .A1(n9056), .A2(n9088), .ZN(n10945) );
  XNOR2_X1 U8597 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n9048) );
  AOI21_X1 U8598 ( .B1(n7524), .B2(n7526), .A(n6579), .ZN(n7522) );
  XNOR2_X1 U8599 ( .A(n8898), .B(n8897), .ZN(n11730) );
  OR2_X1 U8600 ( .A1(n8896), .A2(n8895), .ZN(n8898) );
  INV_X1 U8601 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8528) );
  INV_X1 U8602 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8634) );
  OR2_X1 U8603 ( .A1(n8635), .A2(n8634), .ZN(n8646) );
  NAND2_X1 U8604 ( .A1(n11049), .A2(n11048), .ZN(n6984) );
  NAND2_X1 U8605 ( .A1(n8408), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8725) );
  AND2_X1 U8606 ( .A1(n9708), .A2(n6989), .ZN(n6988) );
  OR2_X1 U8607 ( .A1(n12590), .A2(n6990), .ZN(n6989) );
  INV_X1 U8608 ( .A(n9702), .ZN(n6990) );
  INV_X1 U8609 ( .A(n7252), .ZN(n6987) );
  AOI21_X1 U8610 ( .B1(n12191), .B2(n9708), .A(n6572), .ZN(n7252) );
  AND2_X1 U8611 ( .A1(n7262), .A2(n9763), .ZN(n7261) );
  NAND2_X1 U8612 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8514) );
  INV_X1 U8613 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11994) );
  NAND2_X1 U8614 ( .A1(n7254), .A2(n7253), .ZN(n11581) );
  AOI21_X1 U8615 ( .B1(n7255), .B2(n7257), .A(n6582), .ZN(n7253) );
  NAND2_X1 U8616 ( .A1(n9688), .A2(n7255), .ZN(n7254) );
  OR2_X1 U8617 ( .A1(n8621), .A2(n13777), .ZN(n8635) );
  NAND2_X1 U8618 ( .A1(n9757), .A2(n9756), .ZN(n13726) );
  OR2_X1 U8619 ( .A1(n12190), .A2(n12191), .ZN(n12189) );
  NAND2_X1 U8620 ( .A1(n9688), .A2(n9687), .ZN(n11553) );
  NAND2_X1 U8621 ( .A1(n7189), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U8622 ( .A1(n7187), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U8623 ( .A1(n12832), .A2(n12805), .ZN(n7439) );
  INV_X1 U8624 ( .A(n12858), .ZN(n7144) );
  AND2_X1 U8625 ( .A1(n8732), .A2(n8731), .ZN(n13787) );
  OR2_X1 U8626 ( .A1(n14011), .A2(n8690), .ZN(n8732) );
  AND4_X1 U8627 ( .A1(n8578), .A2(n8577), .A3(n8576), .A4(n8575), .ZN(n11761)
         );
  NAND2_X1 U8628 ( .A1(n8440), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U8629 ( .A1(n7166), .A2(n7164), .ZN(n7162) );
  AND2_X1 U8630 ( .A1(n7170), .A2(n7164), .ZN(n7163) );
  OR2_X1 U8631 ( .A1(n11267), .A2(n11266), .ZN(n11363) );
  NAND2_X1 U8632 ( .A1(n7148), .A2(n7147), .ZN(n11355) );
  NAND2_X1 U8633 ( .A1(n7150), .A2(n7158), .ZN(n7147) );
  XNOR2_X1 U8634 ( .A(n12319), .B(n15407), .ZN(n15411) );
  NOR2_X1 U8635 ( .A1(n15391), .A2(n6617), .ZN(n15404) );
  XNOR2_X1 U8636 ( .A(n13876), .B(n7145), .ZN(n13874) );
  OR2_X1 U8637 ( .A1(n13909), .A2(n15422), .ZN(n13911) );
  AOI21_X1 U8638 ( .B1(n14252), .B2(n8496), .A(n6629), .ZN(n12968) );
  NAND2_X1 U8639 ( .A1(n12969), .A2(n12968), .ZN(n12967) );
  INV_X1 U8640 ( .A(n12968), .ZN(n14100) );
  AND2_X1 U8641 ( .A1(n8774), .A2(n8773), .ZN(n13955) );
  NOR3_X1 U8642 ( .A1(n13992), .A2(n13970), .A3(n14138), .ZN(n13965) );
  NOR2_X1 U8643 ( .A1(n13992), .A2(n14138), .ZN(n13975) );
  NAND2_X1 U8644 ( .A1(n8408), .A2(n7195), .ZN(n8740) );
  INV_X1 U8645 ( .A(n14151), .ZN(n14010) );
  OR2_X1 U8646 ( .A1(n14023), .A2(n8722), .ZN(n7661) );
  OR2_X1 U8647 ( .A1(n14163), .A2(n7401), .ZN(n7400) );
  OR2_X1 U8648 ( .A1(n8688), .A2(n8687), .ZN(n8705) );
  INV_X1 U8649 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n11975) );
  NAND2_X1 U8650 ( .A1(n7603), .A2(n7601), .ZN(n14001) );
  NAND2_X1 U8651 ( .A1(n14044), .A2(n14045), .ZN(n6751) );
  NAND2_X1 U8652 ( .A1(n6940), .A2(n6493), .ZN(n6939) );
  NOR2_X1 U8653 ( .A1(n14188), .A2(n13850), .ZN(n6938) );
  NAND2_X1 U8654 ( .A1(n8407), .A2(n7190), .ZN(n8673) );
  NAND2_X1 U8655 ( .A1(n8407), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U8656 ( .A1(n6936), .A2(n6940), .ZN(n14074) );
  NAND2_X1 U8657 ( .A1(n11869), .A2(n6943), .ZN(n6936) );
  NAND2_X1 U8658 ( .A1(n7647), .A2(n7646), .ZN(n14071) );
  OR2_X1 U8659 ( .A1(n12308), .A2(n12885), .ZN(n7647) );
  OR2_X1 U8660 ( .A1(n6458), .A2(n7669), .ZN(n7668) );
  OR2_X1 U8661 ( .A1(n8628), .A2(n7670), .ZN(n7669) );
  NAND2_X1 U8662 ( .A1(n11698), .A2(n7404), .ZN(n12282) );
  OR2_X1 U8663 ( .A1(n12141), .A2(n12884), .ZN(n12276) );
  NAND2_X1 U8664 ( .A1(n8406), .A2(n7191), .ZN(n8610) );
  OR2_X1 U8665 ( .A1(n11869), .A2(n12882), .ZN(n12140) );
  NAND2_X1 U8666 ( .A1(n11698), .A2(n8885), .ZN(n11873) );
  NAND2_X1 U8667 ( .A1(n7569), .A2(n7568), .ZN(n11701) );
  NAND2_X1 U8668 ( .A1(n8841), .A2(n7570), .ZN(n7569) );
  INV_X1 U8669 ( .A(n11698), .ZN(n11757) );
  NOR2_X1 U8670 ( .A1(n15458), .A2(n9781), .ZN(n10990) );
  OR2_X1 U8671 ( .A1(n8539), .A2(n8528), .ZN(n8562) );
  INV_X1 U8672 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8561) );
  OR2_X1 U8673 ( .A1(n8562), .A2(n8561), .ZN(n8573) );
  OR2_X1 U8674 ( .A1(n12692), .A2(n13861), .ZN(n11341) );
  NOR2_X1 U8675 ( .A1(n12700), .A2(n7398), .ZN(n7397) );
  INV_X1 U8676 ( .A(n15444), .ZN(n7399) );
  NOR2_X1 U8677 ( .A1(n15444), .A2(n7398), .ZN(n11344) );
  NAND2_X1 U8678 ( .A1(n6876), .A2(n6875), .ZN(n8521) );
  NOR2_X1 U8679 ( .A1(n11194), .A2(n15471), .ZN(n15441) );
  NAND2_X1 U8680 ( .A1(n7395), .A2(n11397), .ZN(n11194) );
  INV_X1 U8681 ( .A(n11172), .ZN(n7395) );
  NAND2_X1 U8682 ( .A1(n10694), .A2(n12663), .ZN(n6930) );
  AND2_X1 U8683 ( .A1(n10413), .A2(n8879), .ZN(n13801) );
  INV_X1 U8684 ( .A(n15456), .ZN(n9782) );
  INV_X1 U8685 ( .A(n13930), .ZN(n6956) );
  AND2_X1 U8686 ( .A1(n14115), .A2(n15472), .ZN(n6961) );
  NAND2_X1 U8687 ( .A1(n7586), .A2(n7585), .ZN(n7584) );
  INV_X1 U8688 ( .A(n12864), .ZN(n7585) );
  NAND2_X1 U8689 ( .A1(n8870), .A2(n7588), .ZN(n7587) );
  NOR2_X1 U8690 ( .A1(n12863), .A2(n7589), .ZN(n7588) );
  INV_X1 U8691 ( .A(n8869), .ZN(n7589) );
  NAND2_X1 U8692 ( .A1(n6589), .A2(n7683), .ZN(n7680) );
  NAND2_X1 U8693 ( .A1(n13945), .A2(n12830), .ZN(n7684) );
  NAND2_X1 U8694 ( .A1(n7683), .A2(n7682), .ZN(n7681) );
  INV_X1 U8695 ( .A(n8781), .ZN(n7682) );
  INV_X1 U8696 ( .A(n15443), .ZN(n14166) );
  INV_X1 U8697 ( .A(n13831), .ZN(n14195) );
  AND2_X1 U8698 ( .A1(n12905), .A2(n9784), .ZN(n15472) );
  INV_X1 U8699 ( .A(n15472), .ZN(n15490) );
  NAND2_X1 U8700 ( .A1(n11381), .A2(n8822), .ZN(n8823) );
  AND2_X1 U8701 ( .A1(n10160), .A2(n11730), .ZN(n9796) );
  INV_X1 U8702 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U8703 ( .A1(n8818), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8701) );
  INV_X1 U8704 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8655) );
  NOR2_X1 U8705 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6749) );
  NOR2_X1 U8706 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6748) );
  OR2_X1 U8707 ( .A1(n8555), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8557) );
  OR2_X1 U8708 ( .A1(n8557), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8579) );
  INV_X1 U8709 ( .A(n8605), .ZN(n8501) );
  INV_X1 U8710 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8938) );
  AND2_X1 U8711 ( .A1(n14482), .A2(n14334), .ZN(n14392) );
  INV_X1 U8712 ( .A(n14310), .ZN(n7627) );
  NAND2_X1 U8713 ( .A1(n14494), .A2(n14495), .ZN(n7628) );
  INV_X1 U8714 ( .A(n10802), .ZN(n6735) );
  INV_X1 U8715 ( .A(n11656), .ZN(n7614) );
  XNOR2_X1 U8716 ( .A(n7009), .B(n14359), .ZN(n12213) );
  NAND2_X1 U8717 ( .A1(n7010), .A2(n12036), .ZN(n7009) );
  NAND2_X1 U8718 ( .A1(n12044), .A2(n14346), .ZN(n7010) );
  NAND2_X1 U8719 ( .A1(n8043), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8065) );
  INV_X1 U8720 ( .A(n8045), .ZN(n8043) );
  AND2_X1 U8721 ( .A1(n14390), .A2(n14325), .ZN(n14503) );
  NAND2_X1 U8722 ( .A1(n10475), .A2(n10476), .ZN(n6879) );
  OR2_X1 U8723 ( .A1(n15292), .A2(n14414), .ZN(n10475) );
  AOI21_X1 U8724 ( .B1(n10474), .B2(n10794), .A(n10477), .ZN(n10536) );
  XNOR2_X1 U8725 ( .A(n10788), .B(n6720), .ZN(n6722) );
  INV_X1 U8726 ( .A(n6531), .ZN(n6720) );
  NAND2_X1 U8727 ( .A1(n14770), .A2(n6516), .ZN(n10091) );
  NOR2_X1 U8728 ( .A1(n10094), .A2(n6907), .ZN(n6906) );
  AND2_X1 U8729 ( .A1(n8162), .A2(n8161), .ZN(n14407) );
  INV_X1 U8730 ( .A(n7836), .ZN(n7811) );
  AND2_X1 U8731 ( .A1(n14624), .A2(n10327), .ZN(n14632) );
  NAND2_X1 U8732 ( .A1(n10607), .A2(n10606), .ZN(n14674) );
  NAND2_X1 U8733 ( .A1(n10610), .A2(n10611), .ZN(n10647) );
  OR2_X1 U8734 ( .A1(n10724), .A2(n10725), .ZN(n11002) );
  OR2_X1 U8735 ( .A1(n11005), .A2(n11004), .ZN(n14701) );
  NAND2_X1 U8736 ( .A1(n11010), .A2(n11007), .ZN(n14692) );
  NOR3_X1 U8737 ( .A1(n11644), .A2(n11517), .A3(n11516), .ZN(n12086) );
  NAND2_X1 U8738 ( .A1(n6501), .A2(n9838), .ZN(n6972) );
  AND2_X1 U8739 ( .A1(n8293), .A2(n8306), .ZN(n14794) );
  AND2_X1 U8740 ( .A1(n8352), .A2(n8351), .ZN(n8353) );
  NOR2_X1 U8741 ( .A1(n14824), .A2(n7730), .ZN(n7729) );
  INV_X1 U8742 ( .A(n8250), .ZN(n7730) );
  NAND2_X1 U8743 ( .A1(n8350), .A2(n8347), .ZN(n14817) );
  AND2_X1 U8744 ( .A1(n14918), .A2(n6513), .ZN(n14885) );
  NAND2_X1 U8745 ( .A1(n14918), .A2(n7693), .ZN(n14862) );
  NAND2_X1 U8746 ( .A1(n14931), .A2(n6974), .ZN(n6975) );
  NAND2_X1 U8747 ( .A1(n14915), .A2(n9991), .ZN(n14897) );
  INV_X1 U8748 ( .A(n14911), .ZN(n14896) );
  NAND2_X1 U8749 ( .A1(n14930), .A2(n7436), .ZN(n14915) );
  NAND2_X1 U8750 ( .A1(n14931), .A2(n6905), .ZN(n14930) );
  NAND2_X1 U8751 ( .A1(n6788), .A2(n9972), .ZN(n7702) );
  INV_X1 U8752 ( .A(n14990), .ZN(n7431) );
  INV_X1 U8753 ( .A(n15009), .ZN(n14966) );
  AND3_X1 U8754 ( .A1(n8140), .A2(n8139), .A3(n8138), .ZN(n14967) );
  NAND2_X1 U8755 ( .A1(n9977), .A2(n9954), .ZN(n14989) );
  NAND2_X1 U8756 ( .A1(n7704), .A2(n7703), .ZN(n14985) );
  AOI21_X1 U8757 ( .B1(n7706), .B2(n7708), .A(n6546), .ZN(n7703) );
  NAND2_X1 U8758 ( .A1(n7694), .A2(n12072), .ZN(n15013) );
  NAND2_X1 U8759 ( .A1(n12072), .A2(n7696), .ZN(n15016) );
  NAND2_X1 U8760 ( .A1(n6869), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8029) );
  INV_X1 U8761 ( .A(n8012), .ZN(n6869) );
  AND2_X1 U8762 ( .A1(n7417), .A2(n8329), .ZN(n7416) );
  AND2_X1 U8763 ( .A1(n12072), .A2(n14449), .ZN(n11841) );
  INV_X1 U8764 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7996) );
  OR2_X1 U8765 ( .A1(n7997), .A2(n7996), .ZN(n8012) );
  NAND2_X1 U8766 ( .A1(n12097), .A2(n12098), .ZN(n12096) );
  NAND2_X1 U8767 ( .A1(n6925), .A2(n7986), .ZN(n12097) );
  NAND2_X1 U8768 ( .A1(n7976), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7997) );
  INV_X1 U8769 ( .A(n7978), .ZN(n7976) );
  NAND2_X1 U8770 ( .A1(n7698), .A2(n7697), .ZN(n12102) );
  INV_X1 U8771 ( .A(n7925), .ZN(n7923) );
  INV_X1 U8772 ( .A(n6432), .ZN(n15015) );
  INV_X1 U8773 ( .A(n10548), .ZN(n10546) );
  OAI22_X1 U8774 ( .A1(n10517), .A2(n7810), .B1(n10474), .B2(n10521), .ZN(
        n10545) );
  AND2_X1 U8775 ( .A1(n10511), .A2(n15292), .ZN(n10556) );
  NAND2_X1 U8776 ( .A1(n12943), .A2(n10556), .ZN(n10713) );
  INV_X1 U8777 ( .A(n14587), .ZN(n10509) );
  INV_X1 U8778 ( .A(n15008), .ZN(n14993) );
  NAND2_X1 U8779 ( .A1(n6790), .A2(n10088), .ZN(n6789) );
  NAND2_X1 U8780 ( .A1(n6797), .A2(n6795), .ZN(n6794) );
  NAND2_X1 U8781 ( .A1(n6793), .A2(n6795), .ZN(n6792) );
  NAND2_X1 U8782 ( .A1(n8275), .A2(n8274), .ZN(n15050) );
  OR2_X1 U8783 ( .A1(n7008), .A2(n12156), .ZN(n8274) );
  INV_X1 U8784 ( .A(n14867), .ZN(n15068) );
  NAND2_X1 U8785 ( .A1(n14359), .A2(n7769), .ZN(n15314) );
  XNOR2_X1 U8786 ( .A(n10037), .B(n10036), .ZN(n14252) );
  OAI21_X1 U8787 ( .B1(n9849), .B2(n9848), .A(n9847), .ZN(n10037) );
  XNOR2_X1 U8788 ( .A(n7140), .B(n8798), .ZN(n12944) );
  NAND2_X1 U8789 ( .A1(n8374), .A2(n6451), .ZN(n8377) );
  NAND2_X1 U8790 ( .A1(n7504), .A2(n7503), .ZN(n8395) );
  INV_X1 U8791 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7503) );
  OR2_X1 U8792 ( .A1(n8078), .A2(n8079), .ZN(n6883) );
  NAND2_X1 U8793 ( .A1(n6886), .A2(n6885), .ZN(n6884) );
  XNOR2_X1 U8794 ( .A(n8060), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14698) );
  NAND2_X1 U8795 ( .A1(n6763), .A2(n6529), .ZN(n8052) );
  XNOR2_X1 U8796 ( .A(n8023), .B(n8022), .ZN(n10313) );
  INV_X1 U8797 ( .A(n7470), .ZN(n7473) );
  OR2_X1 U8798 ( .A1(n7992), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n8007) );
  XNOR2_X1 U8799 ( .A(n7941), .B(n7957), .ZN(n10265) );
  AND2_X1 U8800 ( .A1(n7940), .A2(n7958), .ZN(n7941) );
  OR2_X1 U8801 ( .A1(n7846), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n7858) );
  INV_X1 U8802 ( .A(n10162), .ZN(n10220) );
  NAND2_X1 U8803 ( .A1(n10198), .A2(n7297), .ZN(n10221) );
  OR2_X1 U8804 ( .A1(n10202), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n7316) );
  NAND2_X1 U8805 ( .A1(n10202), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10203) );
  NAND2_X1 U8806 ( .A1(n7310), .A2(n10957), .ZN(n10962) );
  NAND2_X1 U8807 ( .A1(n10960), .A2(n10959), .ZN(n10970) );
  AOI21_X1 U8808 ( .B1(n10986), .B2(n6838), .A(n6462), .ZN(n11617) );
  OR2_X1 U8809 ( .A1(n10985), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8810 ( .A1(n6829), .A2(n6826), .ZN(n15232) );
  AOI21_X1 U8811 ( .B1(n15204), .B2(n6828), .A(n6827), .ZN(n6826) );
  NAND2_X1 U8812 ( .A1(n6448), .A2(n6830), .ZN(n6829) );
  NOR2_X1 U8813 ( .A1(n6831), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n6827) );
  AND2_X1 U8814 ( .A1(n9400), .A2(n9389), .ZN(n13371) );
  AND2_X1 U8815 ( .A1(n9331), .A2(n9330), .ZN(n13417) );
  NAND2_X1 U8816 ( .A1(n9321), .A2(n9320), .ZN(n13582) );
  NAND2_X1 U8817 ( .A1(n11604), .A2(n11603), .ZN(n12020) );
  NAND2_X1 U8818 ( .A1(n13061), .A2(n13060), .ZN(n13059) );
  NAND2_X1 U8819 ( .A1(n13170), .A2(n13031), .ZN(n13061) );
  NAND2_X1 U8820 ( .A1(n7377), .A2(n7378), .ZN(n13109) );
  NAND2_X1 U8821 ( .A1(n13024), .A2(n7379), .ZN(n7377) );
  NAND2_X1 U8822 ( .A1(n11181), .A2(n11180), .ZN(n11182) );
  NAND2_X1 U8823 ( .A1(n7385), .A2(n7387), .ZN(n7383) );
  OR2_X1 U8824 ( .A1(n13028), .A2(n13027), .ZN(n13029) );
  NAND2_X1 U8825 ( .A1(n13172), .A2(n13171), .ZN(n13170) );
  INV_X1 U8826 ( .A(n13190), .ZN(n13151) );
  NAND2_X1 U8827 ( .A1(n10873), .A2(n10889), .ZN(n13193) );
  AOI21_X1 U8828 ( .B1(n13024), .B2(n13023), .A(n7382), .ZN(n13189) );
  NAND2_X1 U8829 ( .A1(n10861), .A2(n10860), .ZN(n13195) );
  AND2_X1 U8830 ( .A1(n10870), .A2(n10869), .ZN(n13196) );
  INV_X1 U8831 ( .A(n13387), .ZN(n13204) );
  INV_X1 U8832 ( .A(n15509), .ZN(n13209) );
  OR2_X1 U8833 ( .A1(n12365), .A2(n9570), .ZN(n8946) );
  XNOR2_X1 U8834 ( .A(n9618), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10565) );
  OAI22_X1 U8835 ( .A1(n7223), .A2(n7222), .B1(n6464), .B2(n7221), .ZN(n10740)
         );
  INV_X1 U8836 ( .A(n7229), .ZN(n7221) );
  NAND2_X1 U8837 ( .A1(n7227), .A2(n7229), .ZN(n7222) );
  NAND2_X1 U8838 ( .A1(n9583), .A2(n10785), .ZN(n7229) );
  AND2_X1 U8839 ( .A1(n7097), .A2(n7099), .ZN(n10824) );
  OAI21_X1 U8840 ( .B1(n10832), .B2(n7240), .A(n7239), .ZN(n7242) );
  AOI21_X1 U8841 ( .B1(n10832), .B2(P3_REG1_REG_7__SCAN_IN), .A(n7240), .ZN(
        n10938) );
  AND2_X1 U8842 ( .A1(n7208), .A2(n7205), .ZN(n11299) );
  INV_X1 U8843 ( .A(n7209), .ZN(n7205) );
  NAND2_X1 U8844 ( .A1(n11413), .A2(n11306), .ZN(n7277) );
  NAND2_X1 U8845 ( .A1(n7100), .A2(n6480), .ZN(n11296) );
  NAND2_X1 U8846 ( .A1(n13255), .A2(n6619), .ZN(n13269) );
  NAND2_X1 U8847 ( .A1(n7658), .A2(n10150), .ZN(n13370) );
  OAI21_X1 U8848 ( .B1(n10143), .B2(n12542), .A(n10142), .ZN(n13369) );
  AND2_X1 U8849 ( .A1(n9388), .A2(n9372), .ZN(n13394) );
  XNOR2_X1 U8850 ( .A(n13384), .B(n13389), .ZN(n13573) );
  AND2_X1 U8851 ( .A1(n9371), .A2(n9358), .ZN(n13400) );
  AND2_X1 U8852 ( .A1(n9341), .A2(n9357), .ZN(n13420) );
  NAND2_X1 U8853 ( .A1(n7634), .A2(n9318), .ZN(n13432) );
  NAND2_X1 U8854 ( .A1(n7340), .A2(n12440), .ZN(n11687) );
  OR2_X1 U8855 ( .A1(n15505), .A2(n9477), .ZN(n7340) );
  INV_X1 U8856 ( .A(n15555), .ZN(n13440) );
  NAND2_X1 U8857 ( .A1(n10869), .A2(n15526), .ZN(n15553) );
  OR2_X1 U8858 ( .A1(n6435), .A2(n10177), .ZN(n8955) );
  INV_X1 U8859 ( .A(n15553), .ZN(n15518) );
  NAND2_X1 U8860 ( .A1(n12364), .A2(n12363), .ZN(n13361) );
  NAND2_X1 U8861 ( .A1(n12378), .A2(n12377), .ZN(n13624) );
  AND2_X1 U8862 ( .A1(n7004), .A2(n7005), .ZN(n13456) );
  AND2_X1 U8863 ( .A1(n7352), .A2(n12481), .ZN(n13464) );
  NAND2_X1 U8864 ( .A1(n13499), .A2(n12478), .ZN(n13481) );
  NOR2_X1 U8865 ( .A1(n6674), .A2(n6673), .ZN(n7732) );
  INV_X1 U8866 ( .A(n12473), .ZN(n6673) );
  INV_X1 U8867 ( .A(n13511), .ZN(n6674) );
  NAND2_X1 U8868 ( .A1(n9218), .A2(n9217), .ZN(n13667) );
  INV_X1 U8869 ( .A(n7640), .ZN(n13524) );
  AOI21_X1 U8870 ( .B1(n13535), .B2(n12561), .A(n7643), .ZN(n7640) );
  NAND2_X1 U8871 ( .A1(n9188), .A2(n9187), .ZN(n13679) );
  OR2_X1 U8872 ( .A1(n13554), .A2(n7392), .ZN(n7185) );
  INV_X1 U8873 ( .A(n12029), .ZN(n13692) );
  NAND2_X1 U8874 ( .A1(n7648), .A2(n7650), .ZN(n13557) );
  OR2_X1 U8875 ( .A1(n9123), .A2(n7653), .ZN(n7648) );
  NAND2_X1 U8876 ( .A1(n7654), .A2(n7652), .ZN(n12112) );
  NAND2_X1 U8877 ( .A1(n7337), .A2(n7341), .ZN(n11810) );
  NAND2_X1 U8878 ( .A1(n15505), .A2(n7343), .ZN(n7337) );
  INV_X1 U8879 ( .A(n11019), .ZN(n10936) );
  OR2_X1 U8880 ( .A1(n9447), .A2(P3_D_REG_0__SCAN_IN), .ZN(n10880) );
  AND2_X1 U8881 ( .A1(n7666), .A2(n7665), .ZN(n7664) );
  INV_X1 U8882 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7665) );
  CLKBUF_X1 U8883 ( .A(n9422), .Z(n9423) );
  INV_X1 U8884 ( .A(n8927), .ZN(n9442) );
  INV_X1 U8885 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9435) );
  OAI21_X1 U8886 ( .B1(n9434), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U8887 ( .A1(n7537), .A2(n7536), .ZN(n9365) );
  NAND2_X1 U8888 ( .A1(n9351), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7536) );
  INV_X1 U8889 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U8890 ( .A1(n9434), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U8891 ( .A1(n9272), .A2(n7559), .ZN(n7554) );
  AOI21_X1 U8892 ( .B1(n9286), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n9285), .ZN(
        n9288) );
  XNOR2_X1 U8893 ( .A(n9418), .B(n9417), .ZN(n11640) );
  XNOR2_X1 U8894 ( .A(n9286), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11637) );
  INV_X1 U8895 ( .A(SI_19_), .ZN(n11152) );
  NAND2_X1 U8896 ( .A1(n9253), .A2(n9233), .ZN(n9236) );
  INV_X1 U8897 ( .A(SI_18_), .ZN(n11090) );
  NAND2_X1 U8898 ( .A1(n7549), .A2(n9229), .ZN(n9251) );
  INV_X1 U8899 ( .A(SI_17_), .ZN(n10932) );
  NAND2_X1 U8900 ( .A1(n6810), .A2(n9197), .ZN(n9210) );
  NAND2_X1 U8901 ( .A1(n9196), .A2(n9195), .ZN(n6810) );
  INV_X1 U8902 ( .A(SI_14_), .ZN(n10469) );
  NAND2_X1 U8903 ( .A1(n9161), .A2(n9162), .ZN(n9178) );
  INV_X1 U8904 ( .A(SI_13_), .ZN(n10402) );
  INV_X1 U8905 ( .A(SI_12_), .ZN(n10290) );
  NAND2_X1 U8906 ( .A1(n7545), .A2(n9124), .ZN(n9129) );
  INV_X1 U8907 ( .A(SI_11_), .ZN(n10248) );
  OAI21_X1 U8908 ( .B1(n9069), .B2(n6819), .A(n6817), .ZN(n9107) );
  NAND2_X1 U8909 ( .A1(n6816), .A2(n7527), .ZN(n9104) );
  NAND2_X1 U8910 ( .A1(n9069), .A2(n7529), .ZN(n6816) );
  NAND2_X1 U8911 ( .A1(n7528), .A2(n9071), .ZN(n9086) );
  NAND2_X1 U8912 ( .A1(n9069), .A2(n9068), .ZN(n7528) );
  INV_X1 U8913 ( .A(n10945), .ZN(n10188) );
  XNOR2_X1 U8914 ( .A(n9045), .B(n9044), .ZN(n10840) );
  NAND2_X1 U8915 ( .A1(n9007), .A2(n9006), .ZN(n7523) );
  NAND2_X1 U8916 ( .A1(n8974), .A2(n8973), .ZN(n6823) );
  NAND2_X1 U8917 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8940) );
  OAI21_X1 U8918 ( .B1(n9688), .B2(n7257), .A(n7255), .ZN(n11576) );
  NAND2_X1 U8919 ( .A1(n12596), .A2(n9702), .ZN(n12190) );
  NAND2_X1 U8920 ( .A1(n6984), .A2(n9668), .ZN(n15329) );
  NAND2_X1 U8921 ( .A1(n6991), .A2(n7263), .ZN(n12651) );
  AND2_X1 U8922 ( .A1(n9744), .A2(n7264), .ZN(n7263) );
  NAND2_X1 U8923 ( .A1(n12189), .A2(n9708), .ZN(n12636) );
  NAND2_X1 U8924 ( .A1(n9764), .A2(n7261), .ZN(n13740) );
  NAND2_X1 U8925 ( .A1(n9678), .A2(n12928), .ZN(n12935) );
  NAND2_X1 U8926 ( .A1(n9698), .A2(n12590), .ZN(n12596) );
  NAND2_X1 U8927 ( .A1(n8571), .A2(n8570), .ZN(n12706) );
  NAND2_X1 U8928 ( .A1(n8827), .A2(n11173), .ZN(n12661) );
  NAND2_X1 U8929 ( .A1(n8497), .A2(n14259), .ZN(n6913) );
  AOI21_X1 U8930 ( .B1(n13994), .B2(n8787), .A(n8745), .ZN(n13791) );
  OR2_X1 U8931 ( .A1(n11510), .A2(n8757), .ZN(n8738) );
  AND4_X1 U8932 ( .A1(n8588), .A2(n8587), .A3(n8586), .A4(n8585), .ZN(n12262)
         );
  INV_X1 U8933 ( .A(n13821), .ZN(n13790) );
  NAND2_X1 U8934 ( .A1(n7268), .A2(n7266), .ZN(n13799) );
  NAND2_X1 U8935 ( .A1(n7268), .A2(n7269), .ZN(n13798) );
  AND2_X1 U8936 ( .A1(n7259), .A2(n6519), .ZN(n13810) );
  NAND2_X1 U8937 ( .A1(n8793), .A2(n8792), .ZN(n13839) );
  INV_X1 U8938 ( .A(n13787), .ZN(n13845) );
  OAI21_X1 U8939 ( .B1(n14034), .B2(n8690), .A(n8710), .ZN(n13847) );
  OR2_X1 U8940 ( .A1(n14059), .A2(n8690), .ZN(n8679) );
  NAND2_X1 U8941 ( .A1(n8440), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U8942 ( .A1(n15341), .A2(n6542), .ZN(n15340) );
  AOI21_X1 U8943 ( .B1(n10425), .B2(n15340), .A(n10426), .ZN(n10483) );
  NAND2_X1 U8944 ( .A1(n7167), .A2(n7168), .ZN(n10588) );
  NAND2_X1 U8945 ( .A1(n10502), .A2(n10501), .ZN(n10586) );
  NAND2_X1 U8946 ( .A1(n7152), .A2(n7154), .ZN(n11143) );
  NOR2_X1 U8947 ( .A1(n11356), .A2(n11357), .ZN(n15390) );
  AND2_X1 U8948 ( .A1(n12317), .A2(n12316), .ZN(n15400) );
  OR2_X1 U8949 ( .A1(n15415), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n15417) );
  NAND2_X1 U8950 ( .A1(n12826), .A2(n12825), .ZN(n14093) );
  INV_X1 U8951 ( .A(n13000), .ZN(n12993) );
  NAND2_X1 U8952 ( .A1(n8870), .A2(n8869), .ZN(n13947) );
  XNOR2_X1 U8953 ( .A(n6878), .B(n6877), .ZN(n14123) );
  INV_X1 U8954 ( .A(n13948), .ZN(n6877) );
  NAND2_X1 U8955 ( .A1(n7576), .A2(n8866), .ZN(n13964) );
  NAND2_X1 U8956 ( .A1(n13987), .A2(n7579), .ZN(n7576) );
  NAND2_X1 U8957 ( .A1(n13987), .A2(n8864), .ZN(n13980) );
  NAND2_X1 U8958 ( .A1(n7603), .A2(n12721), .ZN(n14046) );
  NAND2_X1 U8959 ( .A1(n7594), .A2(n8851), .ZN(n12309) );
  NAND2_X1 U8960 ( .A1(n8850), .A2(n7595), .ZN(n7594) );
  NAND2_X1 U8961 ( .A1(n7667), .A2(n8616), .ZN(n12285) );
  NAND2_X1 U8962 ( .A1(n6458), .A2(n7671), .ZN(n7667) );
  NAND2_X1 U8963 ( .A1(n7671), .A2(n7672), .ZN(n12138) );
  OR2_X1 U8964 ( .A1(n6438), .A2(n13916), .ZN(n14089) );
  NAND2_X1 U8965 ( .A1(n7573), .A2(n8835), .ZN(n11058) );
  INV_X1 U8966 ( .A(n14070), .ZN(n14054) );
  OR2_X1 U8967 ( .A1(n6438), .A2(n10994), .ZN(n12149) );
  OAI21_X1 U8968 ( .B1(n14110), .B2(n6752), .A(n6551), .ZN(n14226) );
  NOR2_X1 U8969 ( .A1(n14109), .A2(n14108), .ZN(n6752) );
  INV_X1 U8970 ( .A(n15459), .ZN(n15461) );
  OR2_X1 U8971 ( .A1(n9790), .A2(n15461), .ZN(n15456) );
  NAND2_X1 U8972 ( .A1(n8433), .A2(n7064), .ZN(n7063) );
  INV_X1 U8973 ( .A(n7067), .ZN(n7064) );
  INV_X1 U8974 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8431) );
  XNOR2_X1 U8975 ( .A(n8892), .B(P2_IR_REG_26__SCAN_IN), .ZN(n12351) );
  OAI21_X1 U8976 ( .B1(n8891), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8892) );
  XNOR2_X1 U8977 ( .A(n8887), .B(P2_IR_REG_25__SCAN_IN), .ZN(n12151) );
  INV_X1 U8978 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8889) );
  INV_X1 U8979 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11511) );
  INV_X1 U8980 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11976) );
  INV_X1 U8981 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10767) );
  INV_X1 U8982 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10406) );
  INV_X1 U8983 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10316) );
  INV_X1 U8984 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10275) );
  INV_X1 U8985 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10289) );
  INV_X1 U8986 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10277) );
  INV_X1 U8987 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U8988 ( .A1(n7146), .A2(n8470), .ZN(n10482) );
  INV_X1 U8989 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10172) );
  XNOR2_X1 U8990 ( .A(n8456), .B(n8457), .ZN(n15335) );
  OR2_X1 U8991 ( .A1(n10261), .A2(P1_U3086), .ZN(n10161) );
  NAND2_X1 U8992 ( .A1(n6732), .A2(n6731), .ZN(n14382) );
  NAND2_X1 U8993 ( .A1(n14266), .A2(n14265), .ZN(n6732) );
  CLKBUF_X1 U8994 ( .A(n14393), .Z(n14394) );
  NOR2_X1 U8995 ( .A1(n14403), .A2(n7622), .ZN(n7621) );
  INV_X1 U8996 ( .A(n14293), .ZN(n7622) );
  NAND2_X1 U8997 ( .A1(n14527), .A2(n14293), .ZN(n14404) );
  NOR2_X1 U8998 ( .A1(n7026), .A2(n6711), .ZN(n6710) );
  NAND2_X1 U8999 ( .A1(n7028), .A2(n7027), .ZN(n7026) );
  NAND2_X1 U9000 ( .A1(n7609), .A2(n7607), .ZN(n11666) );
  INV_X1 U9001 ( .A(n7611), .ZN(n7607) );
  OR2_X1 U9002 ( .A1(n10471), .A2(n11660), .ZN(n10472) );
  CLKBUF_X1 U9003 ( .A(n10534), .Z(n10478) );
  NAND2_X1 U9004 ( .A1(n7628), .A2(n14310), .ZN(n14428) );
  INV_X1 U9005 ( .A(n14278), .ZN(n7025) );
  OR2_X1 U9006 ( .A1(n14462), .A2(n7620), .ZN(n7020) );
  AND2_X1 U9007 ( .A1(n8133), .A2(n8132), .ZN(n14955) );
  OR2_X1 U9008 ( .A1(n14462), .A2(n7023), .ZN(n7017) );
  NAND2_X1 U9009 ( .A1(n11023), .A2(n10802), .ZN(n11118) );
  AND2_X1 U9010 ( .A1(n8178), .A2(n8177), .ZN(n14932) );
  INV_X1 U9011 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14509) );
  INV_X1 U9012 ( .A(n6722), .ZN(n6723) );
  NAND2_X1 U9013 ( .A1(n11218), .A2(n11219), .ZN(n6718) );
  NAND2_X1 U9014 ( .A1(n10809), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14556) );
  INV_X1 U9015 ( .A(n14420), .ZN(n14547) );
  NAND2_X1 U9016 ( .A1(n14538), .A2(n14539), .ZN(n14537) );
  AOI21_X1 U9017 ( .B1(n14452), .B2(n6730), .A(n7618), .ZN(n6729) );
  NOR2_X2 U9018 ( .A1(n10392), .A2(n10391), .ZN(n14540) );
  INV_X1 U9019 ( .A(n14540), .ZN(n14561) );
  INV_X1 U9020 ( .A(n10028), .ZN(n14565) );
  INV_X1 U9021 ( .A(n15033), .ZN(n14566) );
  INV_X1 U9022 ( .A(n14543), .ZN(n14567) );
  INV_X1 U9023 ( .A(n14455), .ZN(n14568) );
  NAND2_X1 U9024 ( .A1(n8271), .A2(n8270), .ZN(n14570) );
  OR2_X1 U9025 ( .A1(n14831), .A2(n9851), .ZN(n8271) );
  NAND2_X1 U9026 ( .A1(n8248), .A2(n8247), .ZN(n14571) );
  OR2_X1 U9027 ( .A1(n14843), .A2(n9851), .ZN(n8248) );
  INV_X1 U9028 ( .A(n14932), .ZN(n14900) );
  INV_X1 U9029 ( .A(n14407), .ZN(n14950) );
  INV_X1 U9030 ( .A(n14967), .ZN(n14572) );
  NAND4_X1 U9031 ( .A1(n7922), .A2(n7921), .A3(n7920), .A4(n7919), .ZN(n14581)
         );
  CLKBUF_X1 U9032 ( .A(P1_U4016), .Z(n14580) );
  NAND3_X2 U9033 ( .A1(n7837), .A2(n7414), .A3(n7838), .ZN(n14584) );
  AND2_X1 U9034 ( .A1(n7737), .A2(n7415), .ZN(n7414) );
  INV_X1 U9035 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U9036 ( .A1(n14647), .A2(n14646), .ZN(n14661) );
  OR2_X1 U9037 ( .A1(n11530), .A2(n11529), .ZN(n12084) );
  INV_X1 U9038 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7785) );
  XNOR2_X1 U9039 ( .A(n6861), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14740) );
  NAND2_X1 U9040 ( .A1(n6863), .A2(n6862), .ZN(n6861) );
  NAND2_X1 U9041 ( .A1(n14724), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6863) );
  NAND2_X1 U9042 ( .A1(n10044), .A2(n10043), .ZN(n14756) );
  OR2_X1 U9043 ( .A1(n7008), .A2(n12936), .ZN(n10043) );
  OR2_X1 U9044 ( .A1(n14763), .A2(n8372), .ZN(n14783) );
  AND2_X1 U9045 ( .A1(n8290), .A2(n8289), .ZN(n15048) );
  OR2_X1 U9046 ( .A1(n7008), .A2(n12349), .ZN(n8289) );
  NAND2_X1 U9047 ( .A1(n7723), .A2(n8220), .ZN(n14868) );
  NAND2_X1 U9048 ( .A1(n15167), .A2(n7856), .ZN(n14867) );
  AND2_X1 U9049 ( .A1(n14881), .A2(n14880), .ZN(n15073) );
  OR2_X1 U9050 ( .A1(n7008), .A2(n11406), .ZN(n8204) );
  NAND2_X1 U9051 ( .A1(n8109), .A2(n8108), .ZN(n14981) );
  NAND2_X1 U9052 ( .A1(n7425), .A2(n8334), .ZN(n15007) );
  NAND2_X1 U9053 ( .A1(n11832), .A2(n10080), .ZN(n7705) );
  OAI21_X1 U9054 ( .B1(n6925), .B2(n7719), .A(n7715), .ZN(n12076) );
  NAND2_X1 U9055 ( .A1(n7423), .A2(n8326), .ZN(n11718) );
  NAND2_X1 U9056 ( .A1(n11460), .A2(n8325), .ZN(n7423) );
  NAND2_X1 U9057 ( .A1(n10706), .A2(n10707), .ZN(n7713) );
  INV_X1 U9058 ( .A(n15279), .ZN(n14980) );
  INV_X1 U9059 ( .A(n14997), .ZN(n15301) );
  NAND2_X1 U9060 ( .A1(n7887), .A2(n7888), .ZN(n11213) );
  NAND2_X1 U9061 ( .A1(n15044), .A2(n6842), .ZN(n15126) );
  AND2_X1 U9062 ( .A1(n15043), .A2(n15042), .ZN(n6843) );
  OR2_X1 U9063 ( .A1(n15059), .A2(n15058), .ZN(n15129) );
  OR2_X1 U9064 ( .A1(n15066), .A2(n15065), .ZN(n15130) );
  AND2_X1 U9065 ( .A1(n7913), .A2(n7914), .ZN(n11291) );
  NAND2_X1 U9066 ( .A1(n10252), .A2(n10260), .ZN(n15308) );
  NAND4_X1 U9067 ( .A1(n6717), .A2(n6459), .A3(n7903), .A4(n7432), .ZN(n15152)
         );
  INV_X1 U9068 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7432) );
  INV_X1 U9069 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7793) );
  NAND2_X1 U9070 ( .A1(n7492), .A2(n8272), .ZN(n8273) );
  INV_X1 U9071 ( .A(n7493), .ZN(n7492) );
  NOR2_X1 U9072 ( .A1(n7504), .A2(n7763), .ZN(n7764) );
  NOR2_X1 U9073 ( .A1(n7762), .A2(n15151), .ZN(n6724) );
  NAND2_X1 U9074 ( .A1(n8209), .A2(n8208), .ZN(n11382) );
  INV_X1 U9075 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10956) );
  INV_X1 U9076 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10704) );
  INV_X1 U9077 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10766) );
  INV_X1 U9078 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10408) );
  INV_X1 U9079 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10314) );
  INV_X1 U9080 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10245) );
  AND2_X1 U9081 ( .A1(n10303), .A2(n10214), .ZN(n10235) );
  XNOR2_X1 U9082 ( .A(n10962), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n15171) );
  NAND2_X1 U9083 ( .A1(n7311), .A2(n7312), .ZN(n10988) );
  OR2_X1 U9084 ( .A1(n10986), .A2(n10985), .ZN(n7311) );
  NAND2_X1 U9085 ( .A1(n10986), .A2(n10985), .ZN(n7312) );
  NAND2_X1 U9086 ( .A1(n11849), .A2(n11848), .ZN(n11858) );
  OAI21_X1 U9087 ( .B1(n6836), .B2(n6835), .A(n6576), .ZN(n11862) );
  NOR2_X1 U9088 ( .A1(n11627), .A2(n11629), .ZN(n6835) );
  NAND2_X1 U9089 ( .A1(n11627), .A2(n11629), .ZN(n6834) );
  NAND2_X1 U9090 ( .A1(n7313), .A2(n6538), .ZN(n15190) );
  NOR2_X1 U9091 ( .A1(n7319), .A2(n13199), .ZN(n7317) );
  AOI21_X1 U9092 ( .B1(n6682), .B2(n6683), .A(n6481), .ZN(P3_U3296) );
  AOI21_X1 U9093 ( .B1(n6679), .B2(n12578), .A(n6678), .ZN(n6682) );
  NAND2_X1 U9094 ( .A1(n6684), .A2(n12538), .ZN(n6683) );
  AOI21_X1 U9095 ( .B1(n10570), .B2(n10457), .A(n10456), .ZN(n10459) );
  NAND2_X1 U9096 ( .A1(n7225), .A2(n7226), .ZN(n10770) );
  XNOR2_X1 U9097 ( .A(n7104), .B(n9623), .ZN(n11409) );
  NOR2_X1 U9098 ( .A1(n7273), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7272) );
  AOI21_X1 U9099 ( .B1(n7251), .B2(n9642), .A(n7247), .ZN(n13340) );
  NAND2_X1 U9100 ( .A1(n7250), .A2(n7248), .ZN(n7247) );
  NAND2_X1 U9101 ( .A1(n6866), .A2(n13270), .ZN(n6865) );
  AOI21_X1 U9102 ( .B1(n9615), .B2(n13270), .A(n9614), .ZN(n9644) );
  INV_X1 U9103 ( .A(n9507), .ZN(n9508) );
  OAI21_X1 U9104 ( .B1(n9527), .B2(n13566), .A(n9506), .ZN(n9507) );
  NAND2_X1 U9105 ( .A1(n12613), .A2(n12612), .ZN(n6891) );
  INV_X1 U9106 ( .A(n9496), .ZN(n9497) );
  OAI21_X1 U9107 ( .B1(n7657), .B2(n15609), .A(n7656), .ZN(n10158) );
  NAND2_X1 U9108 ( .A1(n15609), .A2(n10155), .ZN(n7656) );
  OAI21_X1 U9109 ( .B1(n13633), .B2(n15609), .A(n7006), .ZN(P3_U3485) );
  INV_X1 U9110 ( .A(n7007), .ZN(n7006) );
  OAI22_X1 U9111 ( .A1(n13634), .A2(n13598), .B1(n15612), .B2(n13576), .ZN(
        n7007) );
  NOR2_X1 U9112 ( .A1(n13399), .A2(n6668), .ZN(n9653) );
  NOR2_X1 U9113 ( .A1(n6524), .A2(n6923), .ZN(n6922) );
  OR2_X1 U9114 ( .A1(n13631), .A2(n13695), .ZN(n6924) );
  OAI211_X1 U9115 ( .C1(n9522), .C2(n15598), .A(n9529), .B(n6618), .ZN(
        P3_U3455) );
  INV_X1 U9116 ( .A(n9528), .ZN(n9529) );
  OAI21_X1 U9117 ( .B1(n9527), .B2(n13695), .A(n9526), .ZN(n9528) );
  NAND2_X1 U9118 ( .A1(n7657), .A2(n15600), .ZN(n10154) );
  OAI21_X1 U9119 ( .B1(n13633), .B2(n15598), .A(n6887), .ZN(P3_U3453) );
  NOR2_X1 U9120 ( .A1(n6889), .A2(n6888), .ZN(n6887) );
  NOR2_X1 U9121 ( .A1(n15600), .A2(n13632), .ZN(n6888) );
  NOR2_X1 U9122 ( .A1(n13634), .A2(n13654), .ZN(n6889) );
  NAND2_X1 U9123 ( .A1(n6671), .A2(n6477), .ZN(n9656) );
  OAI21_X1 U9124 ( .B1(n9802), .B2(n15327), .A(n9801), .ZN(P2_U3186) );
  XNOR2_X1 U9125 ( .A(n9779), .B(n9778), .ZN(n9802) );
  AOI21_X1 U9126 ( .B1(n14138), .B2(n15332), .A(n13729), .ZN(n6998) );
  INV_X1 U9127 ( .A(n7030), .ZN(P2_U3531) );
  AOI21_X1 U9128 ( .B1(n13858), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n7031), .ZN(
        n7030) );
  NOR2_X1 U9129 ( .A1(n13858), .A2(n7032), .ZN(n7031) );
  NAND2_X1 U9130 ( .A1(n7153), .A2(n7160), .ZN(n11142) );
  AOI21_X1 U9131 ( .B1(n7174), .B2(n13916), .A(n7173), .ZN(n7172) );
  NAND2_X1 U9132 ( .A1(n6957), .A2(n13930), .ZN(n14113) );
  NAND2_X1 U9133 ( .A1(n6901), .A2(n6899), .ZN(P2_U3526) );
  OR2_X1 U9134 ( .A1(n15502), .A2(n6900), .ZN(n6899) );
  NAND2_X1 U9135 ( .A1(n14227), .A2(n15502), .ZN(n6901) );
  INV_X1 U9136 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6900) );
  NAND2_X1 U9137 ( .A1(n8826), .A2(n15496), .ZN(n6958) );
  INV_X1 U9138 ( .A(n6951), .ZN(n6950) );
  OAI21_X1 U9139 ( .B1(n13931), .B2(n6479), .A(n6952), .ZN(n6951) );
  OR2_X1 U9140 ( .A1(n10071), .A2(n7109), .ZN(n6770) );
  AOI21_X1 U9141 ( .B1(n15034), .B2(n15273), .A(n9876), .ZN(n9883) );
  NOR2_X1 U9142 ( .A1(n6622), .A2(n6895), .ZN(n6894) );
  NOR2_X1 U9143 ( .A1(n6896), .A2(n8400), .ZN(n6895) );
  NOR2_X1 U9144 ( .A1(n6623), .A2(n6898), .ZN(n6897) );
  NOR2_X1 U9145 ( .A1(n15319), .A2(n8404), .ZN(n6898) );
  NAND2_X1 U9146 ( .A1(n7309), .A2(n10957), .ZN(n10958) );
  INV_X1 U9147 ( .A(n7310), .ZN(n7309) );
  OAI21_X1 U9148 ( .B1(n15208), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n15207), .ZN(
        n15213) );
  OAI21_X1 U9149 ( .B1(n6463), .B2(n6448), .A(n15223), .ZN(n15225) );
  NAND2_X1 U9150 ( .A1(n15241), .A2(n15244), .ZN(n15242) );
  NOR2_X1 U9151 ( .A1(n15246), .A2(n15245), .ZN(n6824) );
  NOR2_X1 U9152 ( .A1(n6456), .A2(n7306), .ZN(n6448) );
  AND2_X1 U9153 ( .A1(n7370), .A2(n7365), .ZN(n6449) );
  INV_X1 U9154 ( .A(n9924), .ZN(n9920) );
  AND2_X1 U9155 ( .A1(n15215), .A2(n15214), .ZN(n6450) );
  NAND2_X1 U9156 ( .A1(n14405), .A2(n14302), .ZN(n14494) );
  INV_X1 U9157 ( .A(n13862), .ZN(n6875) );
  AND3_X1 U9158 ( .A1(n7772), .A2(n7771), .A3(n7770), .ZN(n6451) );
  NAND2_X1 U9159 ( .A1(n9290), .A2(n9289), .ZN(n13645) );
  AND2_X1 U9160 ( .A1(n8419), .A2(n8434), .ZN(n6452) );
  AND2_X1 U9161 ( .A1(n6484), .A2(n14016), .ZN(n6453) );
  AND2_X1 U9162 ( .A1(n12735), .A2(n12734), .ZN(n6454) );
  NAND2_X1 U9163 ( .A1(n6701), .A2(n6665), .ZN(n15524) );
  AND2_X1 U9164 ( .A1(n7462), .A2(n6544), .ZN(n6455) );
  OR2_X1 U9165 ( .A1(n7307), .A2(n6494), .ZN(n6456) );
  AND2_X1 U9166 ( .A1(n13545), .A2(n12458), .ZN(n6457) );
  INV_X1 U9167 ( .A(n14126), .ZN(n13958) );
  AND2_X1 U9168 ( .A1(n8770), .A2(n8769), .ZN(n14126) );
  INV_X1 U9169 ( .A(n7653), .ZN(n7652) );
  NAND2_X1 U9170 ( .A1(n12113), .A2(n6504), .ZN(n7653) );
  AND2_X1 U9171 ( .A1(n7672), .A2(n6590), .ZN(n6458) );
  NOR2_X1 U9172 ( .A1(n7792), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n6459) );
  NOR2_X1 U9173 ( .A1(n13094), .A2(n7372), .ZN(n6461) );
  NAND2_X1 U9174 ( .A1(n8560), .A2(n8559), .ZN(n14217) );
  INV_X1 U9175 ( .A(n13407), .ZN(n13412) );
  NAND2_X1 U9176 ( .A1(n12500), .A2(n12506), .ZN(n13407) );
  OR2_X1 U9177 ( .A1(n13079), .A2(n13048), .ZN(n12523) );
  AND2_X1 U9178 ( .A1(n10985), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6462) );
  AND2_X1 U9179 ( .A1(n15204), .A2(n7304), .ZN(n6463) );
  AND2_X1 U9180 ( .A1(n7226), .A2(n7224), .ZN(n6464) );
  INV_X1 U9181 ( .A(n14358), .ZN(n7618) );
  INV_X1 U9182 ( .A(n13038), .ZN(n7367) );
  AND2_X1 U9183 ( .A1(n8733), .A2(n9307), .ZN(n6465) );
  INV_X1 U9184 ( .A(n12386), .ZN(n7635) );
  AND2_X1 U9185 ( .A1(n15117), .A2(n14575), .ZN(n6466) );
  AND2_X1 U9186 ( .A1(n9964), .A2(n8142), .ZN(n6467) );
  AND2_X1 U9187 ( .A1(n8042), .A2(n8041), .ZN(n12307) );
  INV_X1 U9188 ( .A(n12307), .ZN(n12236) );
  INV_X1 U9189 ( .A(n13045), .ZN(n13205) );
  OR2_X1 U9190 ( .A1(n9284), .A2(n7630), .ZN(n6468) );
  AND2_X1 U9191 ( .A1(n14583), .A2(n6430), .ZN(n6469) );
  OR2_X1 U9192 ( .A1(n9475), .A2(n9474), .ZN(n6470) );
  AND2_X1 U9193 ( .A1(n10008), .A2(n7122), .ZN(n6471) );
  AND2_X1 U9194 ( .A1(n12789), .A2(n12791), .ZN(n6472) );
  INV_X1 U9195 ( .A(n10590), .ZN(n7164) );
  AND2_X1 U9196 ( .A1(n10009), .A2(n10007), .ZN(n6473) );
  NAND2_X1 U9197 ( .A1(n8087), .A2(n8086), .ZN(n15107) );
  OR2_X1 U9198 ( .A1(n7216), .A2(n7212), .ZN(n6474) );
  AND3_X1 U9199 ( .A1(n8114), .A2(n8113), .A3(n8112), .ZN(n14994) );
  INV_X1 U9200 ( .A(n14994), .ZN(n6981) );
  AND2_X1 U9201 ( .A1(n7697), .A2(n7701), .ZN(n6475) );
  AOI21_X1 U9202 ( .B1(n7567), .B2(n11695), .A(n6554), .ZN(n7566) );
  AND2_X1 U9203 ( .A1(n9304), .A2(n9303), .ZN(n6476) );
  OR2_X1 U9204 ( .A1(n15600), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n6477) );
  INV_X1 U9205 ( .A(n11418), .ZN(n9623) );
  OR2_X1 U9206 ( .A1(n10040), .A2(n12616), .ZN(n6478) );
  OR2_X1 U9207 ( .A1(n6954), .A2(n14186), .ZN(n6479) );
  NAND2_X1 U9208 ( .A1(n7185), .A2(n12458), .ZN(n13542) );
  OR2_X1 U9209 ( .A1(n7102), .A2(n6627), .ZN(n6480) );
  AND2_X1 U9210 ( .A1(n12583), .A2(n12584), .ZN(n6481) );
  AND2_X1 U9211 ( .A1(n9364), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6482) );
  AND2_X1 U9212 ( .A1(n13346), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U9213 ( .A1(n7068), .A2(n6452), .ZN(n14245) );
  INV_X1 U9214 ( .A(n9716), .ZN(n11066) );
  INV_X2 U9215 ( .A(n8516), .ZN(n8483) );
  INV_X1 U9216 ( .A(n6659), .ZN(n15540) );
  NAND2_X1 U9217 ( .A1(n14028), .A2(n13734), .ZN(n6484) );
  NOR2_X1 U9218 ( .A1(n8590), .A2(n12881), .ZN(n6485) );
  AND2_X1 U9219 ( .A1(n13209), .A2(n13087), .ZN(n6486) );
  AND3_X1 U9220 ( .A1(n7854), .A2(n7853), .A3(n7852), .ZN(n6487) );
  INV_X1 U9221 ( .A(n13970), .ZN(n14133) );
  NAND2_X1 U9222 ( .A1(n8759), .A2(n8758), .ZN(n13970) );
  AND2_X1 U9223 ( .A1(n8192), .A2(n11152), .ZN(n6488) );
  INV_X1 U9224 ( .A(n10746), .ZN(n6489) );
  INV_X1 U9225 ( .A(n14475), .ZN(n7016) );
  NAND2_X1 U9226 ( .A1(n9385), .A2(n9384), .ZN(n13374) );
  XNOR2_X1 U9227 ( .A(n13594), .B(n13487), .ZN(n13465) );
  OR2_X1 U9228 ( .A1(n9588), .A2(n10840), .ZN(n6490) );
  INV_X1 U9229 ( .A(n7836), .ZN(n8173) );
  NAND2_X1 U9230 ( .A1(n14848), .A2(n8249), .ZN(n14851) );
  NAND2_X1 U9231 ( .A1(n7725), .A2(n8179), .ZN(n14889) );
  AND2_X1 U9232 ( .A1(n7628), .A2(n7626), .ZN(n6491) );
  OR2_X1 U9233 ( .A1(n7400), .A2(n14081), .ZN(n6492) );
  NAND2_X1 U9234 ( .A1(n7661), .A2(n6453), .ZN(n14017) );
  INV_X1 U9235 ( .A(n10794), .ZN(n14411) );
  XNOR2_X1 U9236 ( .A(n7767), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10092) );
  OR2_X1 U9237 ( .A1(n14086), .A2(n12719), .ZN(n6493) );
  XNOR2_X1 U9238 ( .A(n14780), .B(n14567), .ZN(n10090) );
  AND2_X1 U9239 ( .A1(n15216), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U9240 ( .A1(n15204), .A2(n15203), .ZN(n15207) );
  AND2_X1 U9241 ( .A1(n7330), .A2(n13069), .ZN(n7329) );
  XNOR2_X1 U9242 ( .A(n8931), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8929) );
  OR2_X1 U9243 ( .A1(n7593), .A2(n8853), .ZN(n6495) );
  NOR2_X1 U9244 ( .A1(n12794), .A2(n12792), .ZN(n6496) );
  AND2_X1 U9245 ( .A1(n12566), .A2(n9348), .ZN(n6497) );
  AND2_X1 U9246 ( .A1(n7157), .A2(n7160), .ZN(n6498) );
  AND2_X1 U9247 ( .A1(n12796), .A2(n12795), .ZN(n6499) );
  XNOR2_X1 U9248 ( .A(n12665), .B(n13866), .ZN(n10694) );
  OR2_X1 U9249 ( .A1(n14583), .A2(n6430), .ZN(n6500) );
  INV_X1 U9250 ( .A(n13545), .ZN(n13543) );
  AND2_X1 U9251 ( .A1(n12388), .A2(n12463), .ZN(n13545) );
  INV_X1 U9252 ( .A(n7565), .ZN(n7564) );
  AND2_X1 U9253 ( .A1(n11695), .A2(n7570), .ZN(n7565) );
  OR2_X1 U9254 ( .A1(n14768), .A2(n14566), .ZN(n6501) );
  NAND2_X1 U9255 ( .A1(n14264), .A2(n14263), .ZN(n6502) );
  NAND2_X1 U9256 ( .A1(n13463), .A2(n12490), .ZN(n13453) );
  AND2_X1 U9257 ( .A1(n8080), .A2(n7738), .ZN(n6503) );
  NAND2_X1 U9258 ( .A1(n12449), .A2(n13157), .ZN(n6504) );
  NAND2_X1 U9259 ( .A1(n9413), .A2(n7388), .ZN(n6505) );
  AND2_X1 U9260 ( .A1(n12069), .A2(n11741), .ZN(n6506) );
  NAND2_X1 U9261 ( .A1(n15057), .A2(n14454), .ZN(n6507) );
  XNOR2_X1 U9262 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n8964) );
  INV_X1 U9263 ( .A(n15223), .ZN(n6831) );
  INV_X1 U9264 ( .A(n12561), .ZN(n13534) );
  NAND2_X1 U9265 ( .A1(n6845), .A2(n8965), .ZN(n8974) );
  NAND2_X1 U9266 ( .A1(n7523), .A2(n9008), .ZN(n9022) );
  NAND2_X1 U9267 ( .A1(n7702), .A2(n8142), .ZN(n14928) );
  NAND2_X1 U9268 ( .A1(n8549), .A2(n8548), .ZN(n12692) );
  INV_X1 U9269 ( .A(n14451), .ZN(n6730) );
  OAI21_X1 U9270 ( .B1(SI_10_), .B2(n7141), .A(n8004), .ZN(n8005) );
  AND4_X1 U9271 ( .A1(n14066), .A2(n12888), .A3(n12885), .A4(n12886), .ZN(
        n6508) );
  XNOR2_X1 U9272 ( .A(n13861), .B(n15491), .ZN(n12875) );
  INV_X1 U9273 ( .A(n12875), .ZN(n6859) );
  INV_X1 U9274 ( .A(n11596), .ZN(n7700) );
  INV_X1 U9275 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7541) );
  NAND2_X1 U9276 ( .A1(n8620), .A2(n8619), .ZN(n14206) );
  INV_X1 U9277 ( .A(n14206), .ZN(n7407) );
  AND2_X1 U9278 ( .A1(n7554), .A2(n7558), .ZN(n6509) );
  AND3_X1 U9279 ( .A1(n8415), .A2(n8414), .A3(n8413), .ZN(n6510) );
  INV_X1 U9280 ( .A(n10081), .ZN(n11804) );
  INV_X1 U9281 ( .A(n12518), .ZN(n6696) );
  AND2_X1 U9282 ( .A1(n14856), .A2(n8341), .ZN(n6511) );
  INV_X1 U9283 ( .A(n9620), .ZN(n10822) );
  AND4_X1 U9284 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n8523), .ZN(n6512)
         );
  INV_X1 U9285 ( .A(n12463), .ZN(n7184) );
  AOI21_X1 U9286 ( .B1(n12964), .B2(n15479), .A(n12963), .ZN(n14112) );
  AND2_X1 U9287 ( .A1(n15135), .A2(n15082), .ZN(n6513) );
  AND4_X1 U9288 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n6514)
         );
  AND4_X1 U9289 ( .A1(n6859), .A2(n12873), .A3(n12872), .A4(n15429), .ZN(n6515) );
  AND3_X1 U9290 ( .A1(n6906), .A2(n10090), .A3(n6774), .ZN(n6516) );
  NAND2_X1 U9291 ( .A1(n14527), .A2(n7621), .ZN(n14405) );
  OR3_X1 U9292 ( .A1(n13992), .A2(n7411), .A3(n13970), .ZN(n6517) );
  AND2_X1 U9293 ( .A1(n7647), .A2(n8651), .ZN(n6518) );
  INV_X1 U9294 ( .A(n12703), .ZN(n7056) );
  INV_X1 U9295 ( .A(n9940), .ZN(n7511) );
  INV_X1 U9296 ( .A(n9927), .ZN(n7127) );
  OR2_X1 U9297 ( .A1(n13655), .A2(n13504), .ZN(n12481) );
  NAND2_X1 U9298 ( .A1(n9770), .A2(n9769), .ZN(n6519) );
  AND2_X1 U9299 ( .A1(n7956), .A2(n7960), .ZN(n6520) );
  INV_X1 U9300 ( .A(n9938), .ZN(n7514) );
  NOR2_X1 U9301 ( .A1(n14991), .A2(n8336), .ZN(n6521) );
  OR2_X1 U9302 ( .A1(n9620), .A2(n9012), .ZN(n6522) );
  INV_X1 U9303 ( .A(n10027), .ZN(n15036) );
  AOI21_X1 U9304 ( .B1(n14252), .B2(n10061), .A(n9850), .ZN(n10027) );
  INV_X1 U9305 ( .A(n10000), .ZN(n7112) );
  NAND2_X1 U9306 ( .A1(n8527), .A2(n8526), .ZN(n12700) );
  NAND2_X1 U9307 ( .A1(n8609), .A2(n8608), .ZN(n12733) );
  NAND2_X1 U9308 ( .A1(n9530), .A2(n8921), .ZN(n9111) );
  INV_X1 U9309 ( .A(n9111), .ZN(n6854) );
  AND3_X1 U9310 ( .A1(n6651), .A2(n6650), .A3(n9089), .ZN(n6523) );
  INV_X1 U9311 ( .A(n10016), .ZN(n6841) );
  AND2_X1 U9312 ( .A1(n13630), .A2(n13691), .ZN(n6524) );
  AND2_X1 U9313 ( .A1(n12175), .A2(n12021), .ZN(n6525) );
  INV_X1 U9314 ( .A(n7530), .ZN(n7529) );
  OAI21_X1 U9315 ( .B1(n9068), .B2(n7531), .A(n9085), .ZN(n7530) );
  AND2_X1 U9316 ( .A1(n13032), .A2(n13504), .ZN(n6526) );
  AND2_X1 U9317 ( .A1(n7404), .A2(n7407), .ZN(n6527) );
  AND3_X1 U9318 ( .A1(n13925), .A2(n12896), .A3(n12895), .ZN(n6528) );
  INV_X1 U9319 ( .A(n8848), .ZN(n6946) );
  AND2_X1 U9320 ( .A1(n6762), .A2(n6978), .ZN(n6529) );
  NOR2_X1 U9321 ( .A1(n8856), .A2(n7602), .ZN(n7601) );
  NOR2_X1 U9322 ( .A1(n9482), .A2(n7353), .ZN(n6530) );
  AND4_X1 U9323 ( .A1(n8071), .A2(n8070), .A3(n8069), .A4(n8068), .ZN(n14992)
         );
  INV_X1 U9324 ( .A(n14992), .ZN(n14573) );
  AND2_X1 U9325 ( .A1(n10529), .A2(n10528), .ZN(n6531) );
  AND2_X1 U9326 ( .A1(n13068), .A2(n13387), .ZN(n6532) );
  INV_X1 U9327 ( .A(n12696), .ZN(n7444) );
  NAND2_X1 U9328 ( .A1(n8713), .A2(n8712), .ZN(n14159) );
  OR2_X1 U9329 ( .A1(n13037), .A2(n13429), .ZN(n6533) );
  NOR2_X1 U9330 ( .A1(n12687), .A2(n12684), .ZN(n7078) );
  INV_X1 U9331 ( .A(n12205), .ZN(n14449) );
  NAND2_X1 U9332 ( .A1(n8027), .A2(n8026), .ZN(n12205) );
  AND2_X1 U9333 ( .A1(n6942), .A2(n6493), .ZN(n6534) );
  INV_X1 U9334 ( .A(n9363), .ZN(n7663) );
  AND2_X1 U9335 ( .A1(n7314), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n6535) );
  INV_X1 U9336 ( .A(n8420), .ZN(n8438) );
  INV_X1 U9337 ( .A(n13813), .ZN(n13841) );
  AND2_X1 U9338 ( .A1(n8780), .A2(n8779), .ZN(n13813) );
  AND2_X1 U9339 ( .A1(n7428), .A2(n7427), .ZN(n6536) );
  AND2_X1 U9340 ( .A1(n14086), .A2(n13850), .ZN(n6537) );
  AND2_X1 U9341 ( .A1(n15179), .A2(n15186), .ZN(n6538) );
  OR2_X1 U9342 ( .A1(n14812), .A2(n6778), .ZN(n6539) );
  AND2_X1 U9343 ( .A1(n6500), .A2(n7850), .ZN(n6540) );
  INV_X1 U9344 ( .A(n9935), .ZN(n7516) );
  AND2_X1 U9345 ( .A1(n7515), .A2(n7514), .ZN(n6541) );
  AND2_X1 U9346 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n6542) );
  AND2_X1 U9347 ( .A1(n12520), .A2(n9826), .ZN(n12542) );
  AND2_X1 U9348 ( .A1(n7469), .A2(n8021), .ZN(n6543) );
  INV_X1 U9349 ( .A(n7403), .ZN(n14058) );
  NOR2_X1 U9350 ( .A1(n14081), .A2(n14181), .ZN(n7403) );
  OR2_X1 U9351 ( .A1(n8186), .A2(SI_18_), .ZN(n6544) );
  AND2_X1 U9352 ( .A1(n14787), .A2(n6539), .ZN(n6545) );
  AND2_X1 U9353 ( .A1(n12307), .A2(n14386), .ZN(n6546) );
  OR2_X1 U9354 ( .A1(n7625), .A2(n6728), .ZN(n6547) );
  NAND2_X1 U9355 ( .A1(n9880), .A2(n9879), .ZN(n14770) );
  AND2_X1 U9356 ( .A1(n13970), .A2(n8868), .ZN(n6548) );
  INV_X1 U9357 ( .A(n7716), .ZN(n7715) );
  OR2_X1 U9358 ( .A1(n10825), .A2(n6489), .ZN(n6549) );
  AND2_X1 U9359 ( .A1(n15509), .A2(n13087), .ZN(n6550) );
  AND2_X1 U9360 ( .A1(n14112), .A2(n14111), .ZN(n6551) );
  AND2_X1 U9361 ( .A1(n6712), .A2(n6710), .ZN(n6552) );
  OR2_X1 U9362 ( .A1(n8189), .A2(n8188), .ZN(n6553) );
  AND2_X1 U9363 ( .A1(n8304), .A2(n8303), .ZN(n14365) );
  INV_X1 U9364 ( .A(n14365), .ZN(n14780) );
  AND2_X1 U9365 ( .A1(n14358), .A2(n14356), .ZN(n14452) );
  INV_X1 U9366 ( .A(n14452), .ZN(n7616) );
  INV_X1 U9367 ( .A(n7766), .ZN(n7504) );
  OR2_X1 U9368 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7792) );
  NOR2_X1 U9369 ( .A1(n12706), .A2(n11761), .ZN(n6554) );
  NOR2_X1 U9370 ( .A1(n11723), .A2(n12041), .ZN(n6555) );
  NOR2_X1 U9371 ( .A1(n15068), .A2(n14879), .ZN(n6556) );
  NOR2_X1 U9372 ( .A1(n14010), .A2(n13787), .ZN(n6557) );
  OR2_X1 U9373 ( .A1(n8098), .A2(SI_15_), .ZN(n6558) );
  AND2_X1 U9374 ( .A1(n12125), .A2(n13558), .ZN(n6559) );
  OR2_X1 U9375 ( .A1(n7401), .A2(n14159), .ZN(n6560) );
  INV_X1 U9376 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8523) );
  OR2_X1 U9377 ( .A1(n6494), .A2(n7305), .ZN(n6561) );
  NAND2_X1 U9378 ( .A1(n10589), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U9379 ( .A1(n11783), .A2(n11675), .ZN(n6563) );
  NAND2_X1 U9380 ( .A1(n14181), .A2(n8855), .ZN(n6564) );
  INV_X1 U9381 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10657) );
  INV_X1 U9382 ( .A(n8337), .ZN(n10083) );
  XNOR2_X1 U9383 ( .A(n14981), .B(n6981), .ZN(n8337) );
  AND2_X1 U9384 ( .A1(n12029), .A2(n12246), .ZN(n6565) );
  OR2_X1 U9385 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n6566) );
  INV_X1 U9386 ( .A(n7186), .ZN(n8801) );
  NOR2_X1 U9387 ( .A1(n8784), .A2(n8785), .ZN(n7186) );
  AND2_X1 U9388 ( .A1(n8145), .A2(n10932), .ZN(n6567) );
  NAND2_X1 U9389 ( .A1(n6452), .A2(n14246), .ZN(n6568) );
  INV_X1 U9390 ( .A(n7624), .ZN(n7623) );
  OAI21_X1 U9391 ( .B1(n14495), .B2(n7625), .A(n14502), .ZN(n7624) );
  NOR2_X1 U9392 ( .A1(n13025), .A2(n13113), .ZN(n6569) );
  NAND2_X1 U9393 ( .A1(n14851), .A2(n7729), .ZN(n6570) );
  AND2_X1 U9394 ( .A1(n13594), .A2(n13487), .ZN(n6571) );
  AND2_X1 U9395 ( .A1(n12633), .A2(n9710), .ZN(n6572) );
  INV_X1 U9396 ( .A(n12863), .ZN(n7586) );
  AND2_X1 U9397 ( .A1(n8038), .A2(n10290), .ZN(n6573) );
  AND2_X1 U9398 ( .A1(n14357), .A2(n14452), .ZN(n6574) );
  AND2_X1 U9399 ( .A1(n6841), .A2(n7508), .ZN(n6575) );
  AND2_X1 U9400 ( .A1(n11860), .A2(n6834), .ZN(n6576) );
  BUF_X1 U9401 ( .A(n8939), .Z(n9564) );
  NAND2_X1 U9402 ( .A1(n6916), .A2(n6915), .ZN(n7303) );
  AND2_X1 U9403 ( .A1(n9738), .A2(n9737), .ZN(n6577) );
  INV_X1 U9404 ( .A(n13072), .ZN(n12568) );
  OR2_X1 U9405 ( .A1(n6825), .A2(n6463), .ZN(n6578) );
  INV_X1 U9406 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9460) );
  INV_X1 U9407 ( .A(n7369), .ZN(n13145) );
  NAND2_X1 U9408 ( .A1(n13137), .A2(n6461), .ZN(n7369) );
  AND2_X1 U9409 ( .A1(n10281), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U9410 ( .A1(n7290), .A2(n7291), .ZN(n6580) );
  AND2_X1 U9411 ( .A1(n13026), .A2(n13192), .ZN(n6581) );
  NAND2_X1 U9412 ( .A1(n11590), .A2(n9694), .ZN(n6582) );
  AND2_X1 U9413 ( .A1(n9087), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6583) );
  INV_X1 U9414 ( .A(n7344), .ZN(n7343) );
  OR2_X1 U9415 ( .A1(n9478), .A2(n7345), .ZN(n7344) );
  NAND2_X1 U9416 ( .A1(n13041), .A2(n13042), .ZN(n6584) );
  NOR2_X1 U9417 ( .A1(n14272), .A2(n14271), .ZN(n6585) );
  INV_X1 U9418 ( .A(n14929), .ZN(n6905) );
  NOR2_X1 U9419 ( .A1(n13937), .A2(n13815), .ZN(n6586) );
  OR2_X1 U9420 ( .A1(n9125), .A2(n7546), .ZN(n6587) );
  NAND2_X1 U9421 ( .A1(n9828), .A2(n7347), .ZN(n6588) );
  NAND2_X1 U9422 ( .A1(n7685), .A2(n7684), .ZN(n6589) );
  OR2_X1 U9423 ( .A1(n12733), .A2(n13854), .ZN(n6590) );
  INV_X1 U9424 ( .A(n7150), .ZN(n7149) );
  NAND2_X1 U9425 ( .A1(n7154), .A2(n7151), .ZN(n7150) );
  INV_X1 U9426 ( .A(n7166), .ZN(n7165) );
  NAND2_X1 U9427 ( .A1(n7168), .A2(n6562), .ZN(n7166) );
  INV_X1 U9428 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U9429 ( .A1(n12956), .A2(n8808), .ZN(n14104) );
  INV_X1 U9430 ( .A(n14104), .ZN(n7582) );
  XNOR2_X1 U9431 ( .A(n15254), .B(n15253), .ZN(n6591) );
  OR2_X1 U9432 ( .A1(n7324), .A2(n13073), .ZN(n6592) );
  AND2_X1 U9433 ( .A1(n7418), .A2(n6506), .ZN(n6593) );
  AND2_X1 U9434 ( .A1(n7234), .A2(n7233), .ZN(n6594) );
  AND2_X1 U9435 ( .A1(n7191), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6595) );
  NOR2_X1 U9436 ( .A1(n13797), .A2(n7267), .ZN(n7266) );
  AND2_X1 U9437 ( .A1(n6957), .A2(n6955), .ZN(n6596) );
  AND3_X1 U9438 ( .A1(n8924), .A2(n8923), .A3(n8922), .ZN(n9438) );
  AND2_X1 U9439 ( .A1(n8249), .A2(n6507), .ZN(n6597) );
  AND2_X1 U9440 ( .A1(n14930), .A2(n9988), .ZN(n6598) );
  AND2_X1 U9441 ( .A1(n7903), .A2(n6776), .ZN(n6599) );
  AND2_X1 U9442 ( .A1(n6859), .A2(n8837), .ZN(n6600) );
  NAND2_X1 U9443 ( .A1(n13107), .A2(n13536), .ZN(n6601) );
  AND2_X1 U9444 ( .A1(n13415), .A2(n9348), .ZN(n6602) );
  AND2_X1 U9445 ( .A1(n6924), .A2(n6922), .ZN(n6603) );
  INV_X1 U9446 ( .A(n7243), .ZN(n7240) );
  NAND2_X1 U9447 ( .A1(n9622), .A2(n10840), .ZN(n7243) );
  AND2_X1 U9448 ( .A1(n13407), .A2(n9363), .ZN(n6604) );
  INV_X1 U9449 ( .A(n10166), .ZN(n10462) );
  AND2_X1 U9450 ( .A1(n7261), .A2(n7260), .ZN(n6605) );
  OR2_X1 U9451 ( .A1(n9939), .A2(n7511), .ZN(n6606) );
  OAI21_X1 U9452 ( .B1(n6452), .B2(n7067), .A(n7066), .ZN(n7065) );
  AND2_X1 U9453 ( .A1(n6498), .A2(n7158), .ZN(n6607) );
  AND2_X1 U9454 ( .A1(n6890), .A2(n12614), .ZN(n6608) );
  NAND2_X1 U9455 ( .A1(n9530), .A2(n8962), .ZN(n6609) );
  AND2_X1 U9456 ( .A1(n12523), .A2(n12542), .ZN(n6610) );
  INV_X1 U9457 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n11906) );
  AND2_X1 U9458 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .ZN(n6611) );
  AND2_X1 U9459 ( .A1(n9923), .A2(n7518), .ZN(n6612) );
  INV_X1 U9460 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8434) );
  INV_X1 U9461 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U9462 ( .A1(n12570), .A2(n10147), .ZN(n6613) );
  AND2_X1 U9463 ( .A1(n7661), .A2(n6484), .ZN(n6614) );
  AND2_X2 U9464 ( .A1(n8915), .A2(n10992), .ZN(n15496) );
  INV_X1 U9465 ( .A(n15496), .ZN(n6954) );
  NAND2_X1 U9466 ( .A1(n8816), .A2(n8815), .ZN(n11381) );
  INV_X1 U9467 ( .A(n11381), .ZN(n6993) );
  NAND2_X1 U9468 ( .A1(n6649), .A2(n9102), .ZN(n11811) );
  INV_X1 U9469 ( .A(n15327), .ZN(n13822) );
  INV_X1 U9470 ( .A(n11307), .ZN(n7280) );
  XNOR2_X1 U9471 ( .A(n12160), .B(n14521), .ZN(n12098) );
  INV_X1 U9472 ( .A(n12098), .ZN(n7719) );
  AND2_X1 U9473 ( .A1(n11698), .A2(n7406), .ZN(n6615) );
  NOR2_X1 U9474 ( .A1(n7008), .A2(n10060), .ZN(n6616) );
  INV_X1 U9475 ( .A(n14138), .ZN(n7412) );
  XNOR2_X1 U9476 ( .A(n11617), .B(n11618), .ZN(n15174) );
  INV_X1 U9477 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7817) );
  AND2_X1 U9478 ( .A1(n15397), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6617) );
  INV_X1 U9479 ( .A(n9847), .ZN(n7488) );
  AOI21_X1 U9480 ( .B1(n11755), .B2(n8591), .A(n6485), .ZN(n11866) );
  NAND2_X1 U9481 ( .A1(n9084), .A2(n9083), .ZN(n11688) );
  OR2_X1 U9482 ( .A1(n15600), .A2(n9523), .ZN(n6618) );
  NAND2_X1 U9483 ( .A1(n7705), .A2(n8035), .ZN(n11803) );
  INV_X1 U9484 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n6651) );
  AND2_X1 U9485 ( .A1(n13253), .A2(n13254), .ZN(n6619) );
  AND2_X1 U9486 ( .A1(n13236), .A2(n13237), .ZN(n6620) );
  OR2_X1 U9487 ( .A1(n10083), .A2(n8336), .ZN(n7429) );
  INV_X1 U9488 ( .A(n7429), .ZN(n7427) );
  AND2_X1 U9489 ( .A1(n7020), .A2(n7025), .ZN(n6621) );
  NOR2_X1 U9490 ( .A1(n14365), .A2(n15096), .ZN(n6622) );
  NOR2_X1 U9491 ( .A1(n14365), .A2(n15143), .ZN(n6623) );
  INV_X1 U9492 ( .A(n6943), .ZN(n6942) );
  NOR2_X1 U9493 ( .A1(n6495), .A2(n6944), .ZN(n6943) );
  INV_X1 U9494 ( .A(n7428), .ZN(n14991) );
  NAND2_X1 U9495 ( .A1(n7431), .A2(n7430), .ZN(n7428) );
  INV_X1 U9496 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7192) );
  INV_X1 U9497 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7193) );
  AND2_X1 U9498 ( .A1(n7017), .A2(n7021), .ZN(n6624) );
  NAND2_X1 U9499 ( .A1(n9302), .A2(n9301), .ZN(n6625) );
  NOR2_X1 U9500 ( .A1(n15496), .A2(n6959), .ZN(n6626) );
  OR2_X1 U9501 ( .A1(n9623), .A2(n15610), .ZN(n6627) );
  AND2_X1 U9502 ( .A1(n7609), .A2(n7608), .ZN(n6628) );
  NOR2_X1 U9503 ( .A1(n12824), .A2(n14253), .ZN(n6629) );
  NOR2_X1 U9504 ( .A1(n8254), .A2(SI_23_), .ZN(n6630) );
  AND2_X1 U9505 ( .A1(n7152), .A2(n7149), .ZN(n6631) );
  AND2_X1 U9506 ( .A1(n7185), .A2(n6457), .ZN(n6632) );
  AND2_X1 U9507 ( .A1(n10767), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n6633) );
  INV_X1 U9508 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n6689) );
  AND2_X1 U9509 ( .A1(n7332), .A2(n7333), .ZN(n6634) );
  AND2_X1 U9510 ( .A1(n7190), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6635) );
  AND2_X1 U9511 ( .A1(n6732), .A2(n6502), .ZN(n6636) );
  INV_X1 U9512 ( .A(n12552), .ZN(n9029) );
  AND2_X1 U9513 ( .A1(n12425), .A2(n12424), .ZN(n12552) );
  AND2_X1 U9514 ( .A1(n7277), .A2(n7280), .ZN(n6637) );
  INV_X1 U9515 ( .A(n12807), .ZN(n7440) );
  AND2_X2 U9516 ( .A1(n8403), .A2(n8402), .ZN(n15319) );
  NAND2_X1 U9517 ( .A1(n7995), .A2(n7994), .ZN(n12160) );
  INV_X1 U9518 ( .A(n12160), .ZN(n7701) );
  INV_X1 U9519 ( .A(n13875), .ZN(n7145) );
  INV_X1 U9520 ( .A(n13472), .ZN(n10147) );
  INV_X1 U9521 ( .A(n10053), .ZN(n7490) );
  AND2_X2 U9522 ( .A1(n9501), .A2(n9467), .ZN(n15612) );
  OR2_X1 U9523 ( .A1(n15444), .A2(n12933), .ZN(n6638) );
  INV_X1 U9524 ( .A(n12933), .ZN(n6876) );
  NAND2_X1 U9525 ( .A1(n7713), .A2(n7850), .ZN(n10895) );
  INV_X1 U9526 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11380) );
  INV_X1 U9527 ( .A(n7220), .ZN(n7217) );
  NAND2_X1 U9528 ( .A1(n10867), .A2(n10866), .ZN(n13199) );
  AND2_X1 U9529 ( .A1(n7167), .A2(n7165), .ZN(n6639) );
  NOR2_X1 U9530 ( .A1(n10835), .A2(n9548), .ZN(n6640) );
  INV_X1 U9531 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6870) );
  INV_X1 U9532 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U9533 ( .A1(n10797), .A2(n10796), .ZN(n11023) );
  NAND2_X1 U9534 ( .A1(n9592), .A2(n11418), .ZN(n6641) );
  AND2_X1 U9535 ( .A1(n7225), .A2(n6464), .ZN(n6642) );
  AND2_X1 U9536 ( .A1(n12156), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6643) );
  AND2_X1 U9537 ( .A1(n11511), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6644) );
  INV_X1 U9538 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n6691) );
  OR2_X1 U9539 ( .A1(n9804), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6645) );
  AOI21_X1 U9540 ( .B1(n7093), .B2(n7092), .A(n10166), .ZN(n7084) );
  INV_X1 U9541 ( .A(n7086), .ZN(n7085) );
  INV_X1 U9542 ( .A(n8433), .ZN(n7068) );
  AND2_X1 U9543 ( .A1(n6832), .A2(n10957), .ZN(n6646) );
  INV_X1 U9544 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6914) );
  INV_X1 U9545 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n6908) );
  INV_X1 U9546 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7308) );
  MUX2_X1 U9547 ( .A(n12657), .B(n12656), .S(n15322), .Z(n12658) );
  AND2_X1 U9548 ( .A1(n6649), .A2(n6647), .ZN(n7002) );
  NAND2_X1 U9549 ( .A1(n13544), .A2(n13543), .ZN(n9177) );
  NAND2_X1 U9550 ( .A1(n6657), .A2(n8966), .ZN(n11157) );
  AND2_X1 U9551 ( .A1(n6656), .A2(n8994), .ZN(n11253) );
  NAND3_X1 U9552 ( .A1(n6657), .A2(n8966), .A3(n7733), .ZN(n6656) );
  NAND2_X1 U9553 ( .A1(n15529), .A2(n15528), .ZN(n6657) );
  AOI21_X1 U9554 ( .B1(n13415), .B2(n13414), .A(n13472), .ZN(n13419) );
  NAND2_X2 U9555 ( .A1(n8944), .A2(n6658), .ZN(n6659) );
  AND2_X1 U9556 ( .A1(n8943), .A2(n8945), .ZN(n6658) );
  NAND3_X1 U9557 ( .A1(n6659), .A2(n6660), .A3(n6661), .ZN(n9470) );
  AND2_X1 U9558 ( .A1(n8934), .A2(n8936), .ZN(n6660) );
  AND2_X1 U9559 ( .A1(n8937), .A2(n8935), .ZN(n6661) );
  NAND2_X1 U9560 ( .A1(n6663), .A2(n12417), .ZN(n11444) );
  NAND3_X1 U9561 ( .A1(n7332), .A2(n6699), .A3(n7333), .ZN(n6663) );
  NAND2_X1 U9562 ( .A1(n11154), .A2(n11159), .ZN(n11325) );
  NAND2_X1 U9563 ( .A1(n13553), .A2(n6457), .ZN(n6664) );
  INV_X1 U9564 ( .A(n15524), .ZN(n6700) );
  INV_X1 U9565 ( .A(n6666), .ZN(n6665) );
  NAND2_X1 U9566 ( .A1(n8939), .A2(n10193), .ZN(n9149) );
  NAND3_X1 U9567 ( .A1(n6670), .A2(n6667), .A3(n6669), .ZN(n6671) );
  OR2_X2 U9568 ( .A1(n13406), .A2(n15551), .ZN(n6670) );
  XNOR2_X1 U9569 ( .A(n9646), .B(n12566), .ZN(n13406) );
  NAND3_X1 U9570 ( .A1(n6703), .A2(n6566), .A3(n6676), .ZN(n9424) );
  NAND3_X1 U9571 ( .A1(n6681), .A2(n6610), .A3(n7175), .ZN(n6680) );
  NAND2_X1 U9572 ( .A1(n13425), .A2(n7176), .ZN(n6681) );
  NAND2_X2 U9573 ( .A1(n9483), .A2(n12502), .ZN(n13425) );
  NAND4_X1 U9574 ( .A1(n6686), .A2(n6689), .A3(n6688), .A4(n9181), .ZN(n9214)
         );
  NAND3_X1 U9575 ( .A1(n9239), .A2(n6689), .A3(n6688), .ZN(n6687) );
  NAND4_X1 U9576 ( .A1(n6692), .A2(n9237), .A3(n6691), .A4(n9240), .ZN(n6690)
         );
  OAI21_X2 U9577 ( .B1(n11443), .B2(n6694), .A(n6693), .ZN(n15505) );
  OAI21_X1 U9578 ( .B1(n13425), .B2(n6698), .A(n6695), .ZN(n10143) );
  NAND2_X1 U9579 ( .A1(n6702), .A2(n6700), .ZN(n12407) );
  NAND4_X2 U9580 ( .A1(n8957), .A2(n8959), .A3(n8958), .A4(n8960), .ZN(n15544)
         );
  NAND2_X1 U9581 ( .A1(n7029), .A2(n7617), .ZN(n14373) );
  NAND2_X1 U9582 ( .A1(n14426), .A2(n6708), .ZN(P1_U3220) );
  OR2_X1 U9583 ( .A1(n7029), .A2(n6713), .ZN(n6712) );
  OAI21_X2 U9584 ( .B1(n14266), .B2(n6716), .A(n6714), .ZN(n14462) );
  NAND2_X1 U9585 ( .A1(n6717), .A2(n7903), .ZN(n8380) );
  NAND2_X1 U9586 ( .A1(n6856), .A2(n6717), .ZN(n6855) );
  NAND2_X1 U9587 ( .A1(n6599), .A2(n6717), .ZN(n6777) );
  OAI21_X1 U9588 ( .B1(n11218), .B2(n11219), .A(n11217), .ZN(n6719) );
  NAND2_X1 U9589 ( .A1(n14393), .A2(n14390), .ZN(n14335) );
  NAND2_X1 U9590 ( .A1(n10540), .A2(n6722), .ZN(n10790) );
  XNOR2_X1 U9591 ( .A(n10540), .B(n6723), .ZN(n10544) );
  AND2_X2 U9592 ( .A1(n7757), .A2(n7903), .ZN(n8374) );
  NOR2_X1 U9593 ( .A1(n11117), .A2(n6735), .ZN(n6734) );
  NAND2_X2 U9594 ( .A1(n7061), .A2(n7063), .ZN(n12355) );
  AND2_X2 U9595 ( .A1(n6514), .A2(n6745), .ZN(n8809) );
  NOR2_X2 U9596 ( .A1(n8470), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8498) );
  NAND2_X2 U9597 ( .A1(n8467), .A2(n8417), .ZN(n8470) );
  OAI21_X2 U9598 ( .B1(n14067), .B2(n8681), .A(n8680), .ZN(n14044) );
  NAND2_X2 U9599 ( .A1(n11696), .A2(n12880), .ZN(n11755) );
  OR2_X2 U9600 ( .A1(n11561), .A2(n12878), .ZN(n11560) );
  OAI22_X2 U9601 ( .A1(n13962), .A2(n13963), .B1(n8868), .B2(n14133), .ZN(
        n13952) );
  AOI21_X2 U9602 ( .B1(n13974), .B2(n12865), .A(n12866), .ZN(n13962) );
  NAND2_X1 U9603 ( .A1(n6977), .A2(n8036), .ZN(n6762) );
  NAND3_X1 U9604 ( .A1(n7968), .A2(n7471), .A3(n6976), .ZN(n6763) );
  NAND2_X1 U9605 ( .A1(n6977), .A2(n6754), .ZN(n6753) );
  INV_X1 U9606 ( .A(n8036), .ZN(n6755) );
  NAND4_X1 U9607 ( .A1(n7968), .A2(n7471), .A3(n6976), .A4(n6758), .ZN(n6756)
         );
  NOR2_X1 U9608 ( .A1(n8051), .A2(n6760), .ZN(n6759) );
  INV_X1 U9609 ( .A(n8054), .ZN(n6760) );
  NAND2_X1 U9610 ( .A1(n6768), .A2(n6520), .ZN(n7965) );
  NAND2_X1 U9611 ( .A1(n6768), .A2(n7956), .ZN(n7908) );
  NAND2_X1 U9612 ( .A1(n6857), .A2(n7457), .ZN(n6768) );
  NAND3_X1 U9613 ( .A1(n7106), .A2(n6771), .A3(n6770), .ZN(P1_U3242) );
  AND2_X2 U9614 ( .A1(n6773), .A2(n6772), .ZN(n6771) );
  OR2_X2 U9615 ( .A1(n7108), .A2(n10071), .ZN(n6773) );
  NAND2_X1 U9616 ( .A1(n6775), .A2(n8080), .ZN(n7774) );
  AND2_X1 U9617 ( .A1(n7012), .A2(n7015), .ZN(n7014) );
  AND2_X2 U9618 ( .A1(n6451), .A2(n6775), .ZN(n7012) );
  OAI21_X2 U9619 ( .B1(n14813), .B2(n6778), .A(n6545), .ZN(n14785) );
  NAND2_X1 U9620 ( .A1(n6781), .A2(n11743), .ZN(n6780) );
  NAND3_X1 U9621 ( .A1(n6780), .A2(n6779), .A3(n7706), .ZN(n7704) );
  NAND2_X1 U9622 ( .A1(n6782), .A2(n8018), .ZN(n11832) );
  NAND2_X1 U9623 ( .A1(n6784), .A2(n7714), .ZN(n6782) );
  INV_X1 U9624 ( .A(n14946), .ZN(n6788) );
  NAND2_X1 U9625 ( .A1(n6786), .A2(n6785), .ZN(n14923) );
  AOI21_X1 U9626 ( .B1(n6467), .B2(n8141), .A(n6787), .ZN(n6785) );
  NAND2_X1 U9627 ( .A1(n6467), .A2(n14946), .ZN(n6786) );
  NAND4_X1 U9628 ( .A1(n6794), .A2(n6792), .A3(n6791), .A4(n6789), .ZN(n15039)
         );
  NAND3_X1 U9629 ( .A1(n9878), .A2(n10088), .A3(n7709), .ZN(n6791) );
  OAI211_X1 U9630 ( .C1(n15039), .C2(n15314), .A(n15038), .B(n15037), .ZN(
        n15125) );
  AOI21_X1 U9631 ( .B1(n6798), .B2(n9821), .A(n9431), .ZN(n9522) );
  NAND2_X1 U9632 ( .A1(n9069), .A2(n6817), .ZN(n6815) );
  NAND3_X1 U9633 ( .A1(n6845), .A2(n8975), .A3(n8965), .ZN(n6822) );
  NAND3_X1 U9634 ( .A1(n6822), .A2(n6820), .A3(n8985), .ZN(n6873) );
  NAND2_X1 U9635 ( .A1(n6823), .A2(n8975), .ZN(n8986) );
  XNOR2_X1 U9636 ( .A(n6824), .B(n6591), .ZN(SUB_1596_U4) );
  NAND2_X1 U9637 ( .A1(n6837), .A2(n10295), .ZN(n10298) );
  NAND2_X1 U9638 ( .A1(n10210), .A2(n6837), .ZN(n10213) );
  NAND3_X1 U9639 ( .A1(n10207), .A2(n10295), .A3(n10208), .ZN(n6837) );
  NAND3_X1 U9640 ( .A1(n7311), .A2(n7312), .A3(n10987), .ZN(n11612) );
  NAND3_X1 U9641 ( .A1(n7316), .A2(n7314), .A3(n10203), .ZN(n10215) );
  OAI21_X1 U9642 ( .B1(n7002), .B2(n7001), .A(n9160), .ZN(n13544) );
  INV_X1 U9643 ( .A(n7637), .ZN(n7636) );
  AOI21_X2 U9644 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(n10070) );
  NAND2_X1 U9645 ( .A1(n6892), .A2(n7132), .ZN(n7131) );
  NAND2_X1 U9646 ( .A1(n6893), .A2(n7112), .ZN(n10001) );
  NAND2_X1 U9647 ( .A1(n6873), .A2(n8987), .ZN(n9007) );
  NAND2_X1 U9648 ( .A1(n15191), .A2(n15192), .ZN(n15204) );
  AOI21_X2 U9649 ( .B1(n14761), .B2(n14874), .A(n14760), .ZN(n15044) );
  NAND2_X2 U9650 ( .A1(n11283), .A2(n8324), .ZN(n11460) );
  NAND2_X1 U9651 ( .A1(n11800), .A2(n10081), .ZN(n7425) );
  NAND2_X1 U9652 ( .A1(n8335), .A2(n9955), .ZN(n14990) );
  MUX2_X1 U9653 ( .A(n15264), .B(n15168), .S(n7856), .Z(n10511) );
  NAND3_X1 U9654 ( .A1(n7005), .A2(n7004), .A3(n9299), .ZN(n13455) );
  NAND2_X1 U9655 ( .A1(n8963), .A2(n8964), .ZN(n6845) );
  NAND4_X2 U9656 ( .A1(n8949), .A2(n8948), .A3(n8947), .A4(n8946), .ZN(n15545)
         );
  AOI21_X1 U9657 ( .B1(n12381), .B2(n12527), .A(n7348), .ZN(n12384) );
  NAND2_X1 U9658 ( .A1(n6846), .A2(n11397), .ZN(n8482) );
  NAND3_X1 U9659 ( .A1(n8465), .A2(n8478), .A3(n13865), .ZN(n6846) );
  OAI21_X1 U9660 ( .B1(n12626), .B2(n15475), .A(n7749), .ZN(n8916) );
  OAI21_X1 U9661 ( .B1(n13917), .B2(n13916), .A(n7172), .ZN(P2_U3233) );
  OAI22_X2 U9662 ( .A1(n12133), .A2(n8639), .B1(n12727), .B2(n12726), .ZN(
        n12308) );
  NAND3_X1 U9663 ( .A1(n6851), .A2(n6850), .A3(n7044), .ZN(n7042) );
  NAND2_X1 U9664 ( .A1(n12788), .A2(n12787), .ZN(n6850) );
  NAND2_X1 U9665 ( .A1(n12784), .A2(n12783), .ZN(n6851) );
  NAND2_X1 U9666 ( .A1(n6852), .A2(n6927), .ZN(n6872) );
  NAND2_X1 U9667 ( .A1(n12516), .A2(n12515), .ZN(n6852) );
  NAND3_X1 U9668 ( .A1(n12487), .A2(n13465), .A3(n12488), .ZN(n12492) );
  NAND2_X1 U9669 ( .A1(n12462), .A2(n6853), .ZN(n12464) );
  NAND2_X1 U9670 ( .A1(n9413), .A2(n9409), .ZN(n9411) );
  NAND2_X1 U9671 ( .A1(n12716), .A2(n7037), .ZN(n7036) );
  OAI22_X1 U9672 ( .A1(n12782), .A2(n7449), .B1(n7448), .B2(n12781), .ZN(
        n12785) );
  OAI22_X1 U9673 ( .A1(n12708), .A2(n7454), .B1(n12709), .B2(n7453), .ZN(
        n12714) );
  OAI21_X1 U9674 ( .B1(n12702), .B2(n7051), .A(n7046), .ZN(n7054) );
  NAND3_X1 U9675 ( .A1(n12806), .A2(n12807), .A3(n12832), .ZN(n7438) );
  NAND2_X1 U9676 ( .A1(n7955), .A2(n7954), .ZN(n11714) );
  NAND2_X1 U9677 ( .A1(n14923), .A2(n8340), .ZN(n7725) );
  NAND2_X1 U9678 ( .A1(n7985), .A2(n11737), .ZN(n11743) );
  NAND2_X1 U9679 ( .A1(n7645), .A2(n7644), .ZN(n14067) );
  NOR2_X1 U9680 ( .A1(n13465), .A2(n7743), .ZN(n9283) );
  NAND2_X1 U9681 ( .A1(n6891), .A2(n6608), .ZN(P3_U3488) );
  NAND2_X1 U9682 ( .A1(n7931), .A2(n7700), .ZN(n7933) );
  INV_X1 U9684 ( .A(n6860), .ZN(P2_U3328) );
  OAI211_X1 U9685 ( .C1(n12921), .C2(n12922), .A(n12920), .B(n12919), .ZN(
        n6860) );
  NAND4_X1 U9686 ( .A1(n12894), .A2(n7582), .A3(n14101), .A4(n6528), .ZN(
        n12897) );
  NAND4_X1 U9687 ( .A1(n12887), .A2(n14043), .A3(n12889), .A4(n6508), .ZN(
        n12890) );
  NAND2_X1 U9688 ( .A1(n15234), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7302) );
  NAND2_X1 U9689 ( .A1(n14725), .A2(n14727), .ZN(n6862) );
  XNOR2_X2 U9690 ( .A(n7799), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14595) );
  NAND2_X1 U9691 ( .A1(n7336), .A2(n7334), .ZN(n12111) );
  NAND2_X1 U9692 ( .A1(n9479), .A2(n12456), .ZN(n13553) );
  NAND3_X1 U9693 ( .A1(n6867), .A2(n13358), .A3(n6865), .ZN(P3_U3200) );
  OAI21_X1 U9694 ( .B1(n13349), .B2(n6580), .A(n13348), .ZN(n6867) );
  OAI21_X1 U9695 ( .B1(n13275), .B2(n13273), .A(n13274), .ZN(n13272) );
  INV_X1 U9696 ( .A(n7279), .ZN(n7278) );
  INV_X1 U9697 ( .A(n9546), .ZN(n6919) );
  NOR2_X2 U9698 ( .A1(n9551), .A2(n9623), .ZN(n9552) );
  NAND2_X2 U9699 ( .A1(n8292), .A2(n8266), .ZN(n14831) );
  NAND2_X1 U9700 ( .A1(n7915), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7925) );
  NAND2_X1 U9701 ( .A1(n8240), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8265) );
  NOR2_X2 U9702 ( .A1(n8155), .A2(n8154), .ZN(n6871) );
  INV_X1 U9703 ( .A(n7729), .ZN(n7728) );
  NAND2_X1 U9704 ( .A1(n7728), .A2(n6507), .ZN(n7727) );
  NOR2_X1 U9705 ( .A1(n12541), .A2(n12380), .ZN(n12536) );
  NOR2_X1 U9706 ( .A1(n7535), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7534) );
  NAND2_X1 U9707 ( .A1(n6872), .A2(n12521), .ZN(n12522) );
  NAND2_X1 U9708 ( .A1(n7131), .A2(n9911), .ZN(n7129) );
  XNOR2_X1 U9709 ( .A(n6879), .B(n14359), .ZN(n10535) );
  NAND2_X1 U9710 ( .A1(n7606), .A2(n7605), .ZN(n12223) );
  NAND2_X1 U9711 ( .A1(n7113), .A2(n7110), .ZN(n6893) );
  INV_X1 U9712 ( .A(n7469), .ZN(n6977) );
  NAND2_X1 U9713 ( .A1(n7720), .A2(n7725), .ZN(n7723) );
  NAND3_X1 U9714 ( .A1(n8077), .A2(n6884), .A3(n6883), .ZN(n10703) );
  OAI21_X1 U9715 ( .B1(n14968), .B2(n8337), .A(n8118), .ZN(n14946) );
  OAI21_X1 U9716 ( .B1(n9029), .B2(n6563), .A(n9067), .ZN(n7637) );
  NAND2_X1 U9717 ( .A1(n9283), .A2(n6921), .ZN(n7004) );
  OR2_X1 U9718 ( .A1(n13631), .A2(n13620), .ZN(n6890) );
  NAND3_X1 U9719 ( .A1(n9906), .A2(n10896), .A3(n9905), .ZN(n6892) );
  OAI22_X2 U9720 ( .A1(n14784), .A2(n14787), .B1(n15048), .B2(n14568), .ZN(
        n8355) );
  OAI21_X1 U9721 ( .B1(n9953), .B2(n9944), .A(n9943), .ZN(n9950) );
  NAND2_X1 U9722 ( .A1(n7130), .A2(n7129), .ZN(n9914) );
  OAI21_X1 U9723 ( .B1(n8405), .B2(n15320), .A(n6894), .ZN(P1_U3555) );
  OAI21_X1 U9724 ( .B1(n8405), .B2(n15317), .A(n6897), .ZN(P1_U3523) );
  NAND2_X1 U9725 ( .A1(n7474), .A2(n7989), .ZN(n8006) );
  NAND2_X1 U9726 ( .A1(n7717), .A2(n8003), .ZN(n7716) );
  OAI21_X1 U9727 ( .B1(n13952), .B2(n7681), .A(n7680), .ZN(n13926) );
  NAND2_X2 U9728 ( .A1(n13425), .A2(n7635), .ZN(n13427) );
  NAND3_X2 U9729 ( .A1(n8443), .A2(n8442), .A3(n8441), .ZN(n8827) );
  NAND2_X1 U9730 ( .A1(n7179), .A2(n7177), .ZN(n13442) );
  NAND4_X1 U9731 ( .A1(n10086), .A2(n10087), .A3(n14849), .A4(n14802), .ZN(
        n6907) );
  NAND2_X1 U9732 ( .A1(n6910), .A2(n6909), .ZN(P3_U3160) );
  NAND2_X1 U9733 ( .A1(n7317), .A2(n13179), .ZN(n6909) );
  INV_X1 U9734 ( .A(n6911), .ZN(n6910) );
  NOR2_X2 U9735 ( .A1(n12958), .A2(n12957), .ZN(n12959) );
  OAI21_X2 U9736 ( .B1(n8497), .B2(n6914), .A(n6913), .ZN(n11070) );
  NAND2_X1 U9737 ( .A1(n7302), .A2(n7303), .ZN(n7301) );
  INV_X1 U9738 ( .A(n15231), .ZN(n6915) );
  INV_X1 U9739 ( .A(n15232), .ZN(n6916) );
  NAND2_X1 U9740 ( .A1(n12332), .A2(n12331), .ZN(n15178) );
  NAND2_X1 U9741 ( .A1(n10207), .A2(n10295), .ZN(n10209) );
  NAND2_X1 U9742 ( .A1(n10564), .A2(n10565), .ZN(n10563) );
  NAND2_X1 U9743 ( .A1(n7289), .A2(n13338), .ZN(n7292) );
  NAND2_X1 U9744 ( .A1(n6919), .A2(n6918), .ZN(n6917) );
  INV_X1 U9745 ( .A(n10840), .ZN(n6918) );
  NOR2_X2 U9746 ( .A1(n9552), .A2(n6920), .ZN(n11414) );
  NAND2_X1 U9747 ( .A1(n13445), .A2(n9317), .ZN(n7634) );
  OAI21_X1 U9748 ( .B1(n13629), .B2(n15598), .A(n6603), .ZN(P3_U3456) );
  INV_X1 U9749 ( .A(n7953), .ZN(n7954) );
  NAND2_X1 U9750 ( .A1(n13952), .A2(n7678), .ZN(n6926) );
  INV_X1 U9751 ( .A(n8604), .ZN(n7674) );
  OAI211_X2 U9752 ( .C1(n7671), .C2(n7669), .A(n8627), .B(n7668), .ZN(n12133)
         );
  INV_X1 U9753 ( .A(n9323), .ZN(n9340) );
  NAND2_X1 U9754 ( .A1(n6930), .A2(n8828), .ZN(n10697) );
  NAND2_X1 U9755 ( .A1(n6931), .A2(n6600), .ZN(n11241) );
  INV_X1 U9756 ( .A(n13861), .ZN(n11387) );
  OAI211_X1 U9757 ( .C1(n11346), .C2(n7564), .A(n6932), .B(n7566), .ZN(n11759)
         );
  NAND2_X1 U9758 ( .A1(n11759), .A2(n11760), .ZN(n8844) );
  NAND2_X1 U9759 ( .A1(n6934), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6935) );
  NAND4_X1 U9760 ( .A1(n8809), .A2(n8418), .A3(n8434), .A4(n8498), .ZN(n6934)
         );
  XNOR2_X2 U9761 ( .A(n6935), .B(n8419), .ZN(n8420) );
  OAI21_X2 U9762 ( .B1(n11869), .B2(n6939), .A(n6937), .ZN(n14057) );
  OAI21_X1 U9763 ( .B1(n14116), .B2(n6958), .A(n6950), .ZN(P2_U3494) );
  OAI21_X1 U9764 ( .B1(n14116), .B2(n15475), .A(n6596), .ZN(n14227) );
  INV_X2 U9765 ( .A(n7790), .ZN(n7818) );
  NAND4_X1 U9766 ( .A1(n7785), .A2(n6967), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n6966), .ZN(n6965) );
  INV_X1 U9767 ( .A(n6968), .ZN(n14758) );
  AOI21_X2 U9768 ( .B1(n8355), .B2(n10090), .A(n6969), .ZN(n6968) );
  OAI21_X1 U9769 ( .B1(n8355), .B2(n6972), .A(n6970), .ZN(n6973) );
  NAND2_X2 U9770 ( .A1(n14947), .A2(n8339), .ZN(n14931) );
  NAND2_X1 U9771 ( .A1(n7968), .A2(n7475), .ZN(n7474) );
  NAND3_X1 U9772 ( .A1(n7968), .A2(n7471), .A3(n7475), .ZN(n6980) );
  NAND2_X1 U9773 ( .A1(n6980), .A2(n6543), .ZN(n8037) );
  NAND2_X1 U9774 ( .A1(n9698), .A2(n6988), .ZN(n6985) );
  NAND2_X1 U9775 ( .A1(n6985), .A2(n6986), .ZN(n9711) );
  NAND3_X1 U9776 ( .A1(n13016), .A2(n9725), .A3(n7266), .ZN(n6991) );
  NAND2_X2 U9777 ( .A1(n9657), .A2(n6445), .ZN(n9716) );
  NAND3_X1 U9778 ( .A1(n13731), .A2(n6998), .A3(n6995), .ZN(P2_U3188) );
  NOR2_X4 U9779 ( .A1(n8470), .A2(n8427), .ZN(n8605) );
  NAND2_X1 U9780 ( .A1(n8809), .A2(n8605), .ZN(n8819) );
  NAND2_X1 U9781 ( .A1(n7000), .A2(n6999), .ZN(n15507) );
  NAND3_X1 U9782 ( .A1(n11252), .A2(n9011), .A3(n7636), .ZN(n6999) );
  AND4_X2 U9783 ( .A1(n9112), .A2(n9438), .A3(n9407), .A4(n8925), .ZN(n8927)
         );
  CLKBUF_X1 U9784 ( .A(n7868), .Z(n7008) );
  NAND3_X1 U9785 ( .A1(n7825), .A2(n7756), .A3(n7755), .ZN(n7909) );
  NAND3_X1 U9786 ( .A1(n7903), .A2(n6503), .A3(n7014), .ZN(n7013) );
  NAND3_X1 U9787 ( .A1(n7019), .A2(n7018), .A3(n14287), .ZN(n14528) );
  NAND2_X1 U9788 ( .A1(n13801), .A2(n8827), .ZN(n11169) );
  INV_X1 U9789 ( .A(n8827), .ZN(n7032) );
  NAND2_X1 U9790 ( .A1(n8440), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8519) );
  NAND3_X1 U9791 ( .A1(n7035), .A2(n7034), .A3(n7033), .ZN(n12673) );
  NAND3_X1 U9792 ( .A1(n7437), .A2(n12667), .A3(n12664), .ZN(n7033) );
  NAND2_X1 U9793 ( .A1(n12669), .A2(n12667), .ZN(n7034) );
  NAND3_X1 U9794 ( .A1(n12669), .A2(n7437), .A3(n12664), .ZN(n7035) );
  NAND2_X1 U9795 ( .A1(n12713), .A2(n7039), .ZN(n7038) );
  NAND3_X1 U9796 ( .A1(n7041), .A2(n7038), .A3(n7036), .ZN(n12771) );
  AND2_X1 U9797 ( .A1(n12768), .A2(n12738), .ZN(n7041) );
  NAND2_X1 U9798 ( .A1(n7042), .A2(n7043), .ZN(n7451) );
  INV_X1 U9799 ( .A(n12789), .ZN(n7045) );
  NAND2_X1 U9800 ( .A1(n7054), .A2(n7053), .ZN(n12708) );
  NAND2_X1 U9801 ( .A1(n12801), .A2(n7059), .ZN(n7057) );
  INV_X1 U9802 ( .A(n12802), .ZN(n7060) );
  NOR2_X1 U9803 ( .A1(n7062), .A2(n7065), .ZN(n7061) );
  INV_X1 U9804 ( .A(n12685), .ZN(n7076) );
  OR2_X1 U9805 ( .A1(n12685), .A2(n7078), .ZN(n7075) );
  AOI21_X1 U9806 ( .B1(n7093), .B2(n7092), .A(n10166), .ZN(n7086) );
  NAND3_X1 U9807 ( .A1(n10462), .A2(n7093), .A3(n7092), .ZN(n7087) );
  INV_X1 U9808 ( .A(n10568), .ZN(n7090) );
  INV_X1 U9809 ( .A(n7098), .ZN(n10823) );
  NAND3_X1 U9810 ( .A1(n7236), .A2(n7235), .A3(n7101), .ZN(n7100) );
  AND2_X1 U9811 ( .A1(n11303), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7103) );
  NOR2_X4 U9812 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n9530) );
  NAND2_X4 U9813 ( .A1(n10033), .A2(n7105), .ZN(n9924) );
  NAND2_X1 U9814 ( .A1(n9884), .A2(n9885), .ZN(n9887) );
  NAND2_X2 U9815 ( .A1(n10048), .A2(n9886), .ZN(n10033) );
  NAND3_X1 U9816 ( .A1(n7108), .A2(n7109), .A3(n7107), .ZN(n7106) );
  NAND2_X1 U9817 ( .A1(n10070), .A2(n10069), .ZN(n7108) );
  NAND2_X1 U9818 ( .A1(n9994), .A2(n7115), .ZN(n7113) );
  NAND2_X1 U9819 ( .A1(n7113), .A2(n7111), .ZN(n9999) );
  NAND2_X1 U9820 ( .A1(n10004), .A2(n7120), .ZN(n7119) );
  NAND2_X1 U9821 ( .A1(n7119), .A2(n7118), .ZN(n10011) );
  NAND2_X1 U9822 ( .A1(n7125), .A2(n7123), .ZN(n9929) );
  NAND2_X1 U9823 ( .A1(n9926), .A2(n7126), .ZN(n7125) );
  OAI21_X1 U9824 ( .B1(n9911), .B2(n7131), .A(n9910), .ZN(n7130) );
  NAND2_X1 U9825 ( .A1(n9909), .A2(n9908), .ZN(n7132) );
  NAND2_X1 U9826 ( .A1(n7133), .A2(n7510), .ZN(n9953) );
  NAND3_X1 U9827 ( .A1(n7135), .A2(n7134), .A3(n6606), .ZN(n7133) );
  NAND2_X1 U9828 ( .A1(n9937), .A2(n9936), .ZN(n7134) );
  OAI21_X2 U9829 ( .B1(n8120), .B2(n7138), .A(n8124), .ZN(n8129) );
  MUX2_X1 U9830 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n10193), .Z(n7141) );
  NAND3_X1 U9831 ( .A1(n7143), .A2(n7142), .A3(n12862), .ZN(n12922) );
  NAND3_X1 U9832 ( .A1(n7144), .A2(n12808), .A3(n7440), .ZN(n7142) );
  NAND3_X1 U9833 ( .A1(n7438), .A2(n7144), .A3(n7439), .ZN(n7143) );
  MUX2_X1 U9834 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n8460), .S(n10482), .Z(n10426) );
  MUX2_X1 U9835 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8469), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n7146) );
  MUX2_X1 U9836 ( .A(n10423), .B(P2_REG1_REG_1__SCAN_IN), .S(n15335), .Z(
        n15341) );
  NAND2_X1 U9837 ( .A1(n10922), .A2(n6607), .ZN(n7148) );
  OR2_X1 U9838 ( .A1(n11140), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7159) );
  NAND2_X1 U9839 ( .A1(n7163), .A2(n15364), .ZN(n7161) );
  NAND2_X1 U9840 ( .A1(n7162), .A2(n7161), .ZN(n10674) );
  NAND3_X1 U9841 ( .A1(n8955), .A2(n8953), .A3(n8954), .ZN(n11019) );
  NAND2_X1 U9842 ( .A1(n7189), .A2(n6611), .ZN(n8539) );
  NAND2_X1 U9843 ( .A1(n8407), .A2(n6635), .ZN(n8688) );
  NAND2_X1 U9844 ( .A1(n8406), .A2(n6595), .ZN(n8621) );
  INV_X1 U9845 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7197) );
  NAND3_X1 U9846 ( .A1(n10150), .A2(n7658), .A3(n7655), .ZN(n7657) );
  OAI21_X2 U9847 ( .B1(n12997), .B2(n8690), .A(n8807), .ZN(n13838) );
  NAND2_X1 U9848 ( .A1(n12971), .A2(n8802), .ZN(n12997) );
  NOR2_X1 U9849 ( .A1(n7202), .A2(n13354), .ZN(n7201) );
  NOR2_X1 U9850 ( .A1(n13344), .A2(n13345), .ZN(n13343) );
  INV_X1 U9851 ( .A(n9607), .ZN(n7204) );
  NAND2_X1 U9852 ( .A1(n10834), .A2(n7213), .ZN(n7208) );
  OAI21_X1 U9853 ( .B1(n10834), .B2(n10833), .A(n6490), .ZN(n10941) );
  AOI21_X1 U9854 ( .B1(n10833), .B2(n6490), .A(n7219), .ZN(n7218) );
  NAND2_X1 U9855 ( .A1(n9590), .A2(n10945), .ZN(n7220) );
  INV_X1 U9856 ( .A(n10570), .ZN(n7223) );
  INV_X1 U9857 ( .A(n7234), .ZN(n13298) );
  XNOR2_X1 U9858 ( .A(n9604), .B(n10672), .ZN(n13300) );
  NAND3_X1 U9859 ( .A1(n7237), .A2(n7241), .A3(n7243), .ZN(n7236) );
  INV_X1 U9860 ( .A(n10832), .ZN(n7237) );
  INV_X1 U9861 ( .A(n7242), .ZN(n10937) );
  INV_X1 U9862 ( .A(n7246), .ZN(n10779) );
  NOR2_X1 U9863 ( .A1(n8501), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U9864 ( .A1(n9764), .A2(n6605), .ZN(n7259) );
  OR2_X1 U9865 ( .A1(n9766), .A2(n9765), .ZN(n7262) );
  OAI21_X1 U9866 ( .B1(n12599), .B2(n9735), .A(n9734), .ZN(n12610) );
  NAND2_X1 U9867 ( .A1(n7270), .A2(n13304), .ZN(n7271) );
  INV_X1 U9868 ( .A(n9555), .ZN(n7270) );
  AND3_X2 U9869 ( .A1(n7271), .A2(n9556), .A3(P3_REG2_REG_15__SCAN_IN), .ZN(
        n13321) );
  NOR2_X1 U9870 ( .A1(n13321), .A2(n7272), .ZN(n13306) );
  NOR2_X1 U9871 ( .A1(n7275), .A2(n7274), .ZN(n7281) );
  NAND2_X1 U9872 ( .A1(n11303), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7282) );
  NAND3_X1 U9873 ( .A1(n9541), .A2(P3_REG2_REG_5__SCAN_IN), .A3(n9542), .ZN(
        n10742) );
  OAI21_X1 U9874 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n7285), .A(n10742), .ZN(
        n10743) );
  INV_X1 U9875 ( .A(n9558), .ZN(n7289) );
  NAND2_X1 U9876 ( .A1(n7292), .A2(n9559), .ZN(n13329) );
  NAND3_X1 U9877 ( .A1(n7290), .A2(n7291), .A3(n9561), .ZN(n9562) );
  NAND3_X1 U9878 ( .A1(n7292), .A2(n9559), .A3(n6483), .ZN(n7291) );
  NAND3_X1 U9879 ( .A1(n10299), .A2(n10300), .A3(n10959), .ZN(n10960) );
  INV_X1 U9880 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7296) );
  NAND3_X1 U9881 ( .A1(n7302), .A2(n7303), .A3(n15240), .ZN(n15244) );
  NAND2_X1 U9882 ( .A1(n7301), .A2(n7300), .ZN(n15241) );
  INV_X1 U9883 ( .A(n15240), .ZN(n7300) );
  NAND2_X1 U9884 ( .A1(n15175), .A2(n11984), .ZN(n7313) );
  NAND2_X1 U9885 ( .A1(n7313), .A2(n15179), .ZN(n15188) );
  NAND2_X1 U9886 ( .A1(n7316), .A2(n10203), .ZN(n7315) );
  INV_X1 U9887 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7314) );
  NAND2_X1 U9888 ( .A1(n7315), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U9889 ( .A1(n9539), .A2(n6489), .ZN(n9541) );
  INV_X1 U9890 ( .A(n10298), .ZN(n10297) );
  NAND2_X1 U9891 ( .A1(n9711), .A2(n12632), .ZN(n12639) );
  OAI21_X1 U9892 ( .B1(n13179), .B2(n13180), .A(n7331), .ZN(n13070) );
  NAND2_X1 U9893 ( .A1(n9471), .A2(n12407), .ZN(n11154) );
  NAND2_X1 U9894 ( .A1(n11079), .A2(n11180), .ZN(n11081) );
  NAND2_X1 U9895 ( .A1(n11075), .A2(n11074), .ZN(n11082) );
  NAND2_X1 U9896 ( .A1(n7350), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9131) );
  NOR2_X1 U9897 ( .A1(n7350), .A2(n9214), .ZN(n9238) );
  NOR2_X1 U9898 ( .A1(n7350), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U9899 ( .A1(n9113), .A2(n7350), .ZN(n13222) );
  NAND2_X1 U9900 ( .A1(n7354), .A2(n7357), .ZN(n13139) );
  NAND2_X1 U9901 ( .A1(n13172), .A2(n7355), .ZN(n7354) );
  NAND2_X1 U9902 ( .A1(n9447), .A2(n10879), .ZN(n7360) );
  NAND2_X1 U9903 ( .A1(n13137), .A2(n6449), .ZN(n7364) );
  NAND2_X1 U9904 ( .A1(n13137), .A2(n13034), .ZN(n13093) );
  INV_X1 U9905 ( .A(n13034), .ZN(n7372) );
  NAND2_X1 U9906 ( .A1(n11604), .A2(n7385), .ZN(n7384) );
  NAND3_X1 U9907 ( .A1(n7384), .A2(n12025), .A3(n7383), .ZN(n12249) );
  NAND4_X1 U9908 ( .A1(n9407), .A2(n9112), .A3(n8925), .A4(n7393), .ZN(n7394)
         );
  INV_X2 U9909 ( .A(n11397), .ZN(n12670) );
  AND3_X2 U9910 ( .A1(n8475), .A2(n8476), .A3(n8477), .ZN(n15466) );
  OAI211_X1 U9911 ( .C1(n12969), .C2(n12968), .A(n15443), .B(n12967), .ZN(
        n14099) );
  NAND2_X1 U9912 ( .A1(n15491), .A2(n6876), .ZN(n7398) );
  AND2_X2 U9913 ( .A1(n7399), .A2(n7397), .ZN(n11345) );
  INV_X1 U9914 ( .A(n11344), .ZN(n8884) );
  NOR3_X2 U9915 ( .A1(n14081), .A2(n14163), .A3(n6560), .ZN(n14008) );
  NOR2_X2 U9916 ( .A1(n13992), .A2(n7408), .ZN(n7413) );
  INV_X1 U9917 ( .A(n7413), .ZN(n13940) );
  NAND2_X1 U9918 ( .A1(n10708), .A2(n10073), .ZN(n8320) );
  NAND3_X1 U9919 ( .A1(n7418), .A2(n7420), .A3(n6506), .ZN(n7417) );
  NAND2_X1 U9920 ( .A1(n7425), .A2(n7424), .ZN(n8335) );
  INV_X1 U9921 ( .A(n8355), .ZN(n9839) );
  AOI21_X1 U9922 ( .B1(n14990), .B2(n7427), .A(n7426), .ZN(n14949) );
  OAI22_X1 U9923 ( .A1(n12680), .A2(n7442), .B1(n12681), .B2(n7441), .ZN(
        n12685) );
  NAND2_X1 U9924 ( .A1(n7445), .A2(n7443), .ZN(n12694) );
  NAND2_X1 U9925 ( .A1(n12689), .A2(n7446), .ZN(n7445) );
  NAND2_X1 U9926 ( .A1(n12785), .A2(n12786), .ZN(n12784) );
  NAND2_X1 U9927 ( .A1(n7451), .A2(n7452), .ZN(n12797) );
  NAND2_X1 U9928 ( .A1(n12714), .A2(n12715), .ZN(n12713) );
  OAI21_X1 U9929 ( .B1(n7865), .B2(n7864), .A(n7863), .ZN(n7458) );
  NAND2_X1 U9930 ( .A1(n7864), .A2(n7863), .ZN(n7456) );
  NAND2_X1 U9931 ( .A1(n7865), .A2(n7863), .ZN(n7457) );
  NAND2_X1 U9932 ( .A1(n7458), .A2(n7881), .ZN(n7882) );
  XNOR2_X1 U9933 ( .A(n7458), .B(n7880), .ZN(n10197) );
  INV_X1 U9934 ( .A(n8252), .ZN(n7466) );
  INV_X1 U9935 ( .A(n8005), .ZN(n7467) );
  NAND2_X1 U9936 ( .A1(n7468), .A2(n8004), .ZN(n8023) );
  NAND2_X1 U9937 ( .A1(n7474), .A2(n7473), .ZN(n7468) );
  INV_X1 U9938 ( .A(n8004), .ZN(n7472) );
  NAND2_X1 U9939 ( .A1(n7968), .A2(n7967), .ZN(n7991) );
  NOR2_X1 U9940 ( .A1(n7990), .A2(n7476), .ZN(n7475) );
  INV_X1 U9941 ( .A(n7967), .ZN(n7476) );
  NAND2_X1 U9942 ( .A1(n9849), .A2(n9847), .ZN(n7477) );
  NAND2_X1 U9943 ( .A1(n7477), .A2(n7486), .ZN(n10056) );
  NAND2_X1 U9944 ( .A1(n10057), .A2(n7478), .ZN(n14244) );
  OAI21_X1 U9945 ( .B1(n9849), .B2(n7484), .A(n7480), .ZN(n7479) );
  INV_X1 U9946 ( .A(n9848), .ZN(n7491) );
  NAND2_X1 U9947 ( .A1(n10097), .A2(n9920), .ZN(n7501) );
  XNOR2_X2 U9948 ( .A(n7502), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8371) );
  INV_X1 U9949 ( .A(n9887), .ZN(n7505) );
  NAND2_X1 U9950 ( .A1(n7507), .A2(n7506), .ZN(n10015) );
  NAND2_X1 U9951 ( .A1(n10011), .A2(n7508), .ZN(n7507) );
  NAND2_X1 U9952 ( .A1(n9934), .A2(n7515), .ZN(n7512) );
  NAND2_X1 U9953 ( .A1(n7512), .A2(n7513), .ZN(n9937) );
  AOI21_X1 U9954 ( .B1(n7517), .B2(n7515), .A(n7514), .ZN(n7513) );
  OAI22_X1 U9955 ( .A1(n9922), .A2(n6612), .B1(n9923), .B2(n7518), .ZN(n9926)
         );
  NAND2_X1 U9956 ( .A1(n7521), .A2(n7522), .ZN(n9040) );
  NAND2_X1 U9957 ( .A1(n9007), .A2(n7524), .ZN(n7521) );
  NAND2_X1 U9958 ( .A1(n9349), .A2(n7534), .ZN(n7533) );
  NAND2_X1 U9959 ( .A1(n7533), .A2(n7532), .ZN(n9380) );
  NAND2_X1 U9960 ( .A1(n7540), .A2(n7542), .ZN(n7538) );
  NAND2_X1 U9961 ( .A1(n9146), .A2(n7540), .ZN(n7539) );
  NAND2_X1 U9962 ( .A1(n9107), .A2(n9106), .ZN(n9126) );
  NAND2_X1 U9963 ( .A1(n9212), .A2(n9211), .ZN(n9231) );
  NAND2_X1 U9964 ( .A1(n9272), .A2(n7555), .ZN(n7552) );
  NAND2_X1 U9965 ( .A1(n7552), .A2(n7553), .ZN(n9334) );
  NAND2_X1 U9966 ( .A1(n9382), .A2(n7562), .ZN(n7561) );
  NAND2_X1 U9967 ( .A1(n7561), .A2(n9396), .ZN(n9803) );
  NAND2_X1 U9968 ( .A1(n7561), .A2(n7560), .ZN(n9806) );
  NAND2_X2 U9969 ( .A1(n8450), .A2(n8420), .ZN(n8516) );
  NAND3_X1 U9970 ( .A1(n8450), .A2(n8420), .A3(P2_REG2_REG_2__SCAN_IN), .ZN(
        n8464) );
  NAND2_X1 U9971 ( .A1(n13987), .A2(n6460), .ZN(n7574) );
  NAND2_X1 U9972 ( .A1(n7574), .A2(n7575), .ZN(n13954) );
  OR2_X1 U9973 ( .A1(n7579), .A2(n7578), .ZN(n7577) );
  NAND2_X1 U9974 ( .A1(n7587), .A2(n7581), .ZN(n7583) );
  INV_X1 U9975 ( .A(n7583), .ZN(n13927) );
  NAND2_X1 U9976 ( .A1(n7587), .A2(n7584), .ZN(n13929) );
  NAND2_X1 U9977 ( .A1(n8850), .A2(n8849), .ZN(n12129) );
  NOR2_X1 U9978 ( .A1(n8852), .A2(n7596), .ZN(n7595) );
  INV_X1 U9979 ( .A(n8849), .ZN(n7596) );
  INV_X1 U9980 ( .A(n14057), .ZN(n7604) );
  NAND2_X1 U9981 ( .A1(n7597), .A2(n7598), .ZN(n8863) );
  NAND2_X1 U9982 ( .A1(n10539), .A2(n10538), .ZN(n10540) );
  NAND3_X1 U9983 ( .A1(n11476), .A2(n7613), .A3(n12034), .ZN(n7606) );
  NOR2_X1 U9984 ( .A1(n7611), .A2(n11665), .ZN(n7608) );
  OAI22_X1 U9985 ( .A1(n11656), .A2(n7612), .B1(n11654), .B2(n11655), .ZN(
        n7611) );
  AND2_X1 U9986 ( .A1(n11475), .A2(n7614), .ZN(n7613) );
  NAND2_X1 U9987 ( .A1(n7631), .A2(n9228), .ZN(n13466) );
  INV_X1 U9988 ( .A(n9228), .ZN(n7630) );
  NAND2_X1 U9989 ( .A1(n7634), .A2(n7632), .ZN(n13430) );
  NAND2_X1 U9990 ( .A1(n12308), .A2(n7646), .ZN(n7645) );
  NAND2_X1 U9991 ( .A1(n13369), .A2(n15596), .ZN(n7655) );
  NAND2_X1 U9992 ( .A1(n7659), .A2(n7660), .ZN(n13984) );
  NAND2_X1 U9993 ( .A1(n14023), .A2(n6453), .ZN(n7659) );
  NAND2_X1 U9994 ( .A1(n8927), .A2(n7664), .ZN(n13697) );
  NAND2_X2 U9995 ( .A1(n11755), .A2(n7675), .ZN(n7671) );
  NAND3_X2 U9996 ( .A1(n7830), .A2(n7829), .A3(n7828), .ZN(n10530) );
  NAND3_X1 U9997 ( .A1(n12943), .A2(n10556), .A3(n7686), .ZN(n10901) );
  INV_X2 U9998 ( .A(n10530), .ZN(n12943) );
  NAND2_X1 U9999 ( .A1(n14793), .A2(n7687), .ZN(n7689) );
  INV_X1 U10000 ( .A(n7689), .ZN(n14752) );
  AOI21_X1 U10001 ( .B1(n14762), .B2(n15036), .A(n15015), .ZN(n7690) );
  NAND2_X1 U10002 ( .A1(n7691), .A2(n14918), .ZN(n14844) );
  NAND3_X1 U10003 ( .A1(n7694), .A2(n15003), .A3(n12072), .ZN(n15000) );
  NAND2_X1 U10004 ( .A1(n7698), .A2(n6475), .ZN(n7740) );
  NAND3_X1 U10005 ( .A1(n7832), .A2(n7831), .A3(n6540), .ZN(n7711) );
  NAND2_X1 U10006 ( .A1(n7712), .A2(n7711), .ZN(n11100) );
  NAND2_X1 U10007 ( .A1(n14848), .A2(n6597), .ZN(n7726) );
  NAND2_X1 U10008 ( .A1(n7726), .A2(n7727), .ZN(n14813) );
  CLKBUF_X1 U10009 ( .A(n14008), .Z(n14024) );
  INV_X1 U10010 ( .A(n14163), .ZN(n14033) );
  OR3_X1 U10011 ( .A1(n12260), .A2(n9446), .A3(n13720), .ZN(n10854) );
  AND2_X1 U10012 ( .A1(n8605), .A2(n6510), .ZN(n8428) );
  NAND2_X1 U10013 ( .A1(n12249), .A2(n12248), .ZN(n12252) );
  OAI21_X2 U10014 ( .B1(n13321), .B2(n13320), .A(n13319), .ZN(n13323) );
  OR2_X1 U10015 ( .A1(n11738), .A2(n11737), .ZN(n12067) );
  OR2_X1 U10016 ( .A1(n14222), .A2(n12899), .ZN(n9792) );
  INV_X1 U10017 ( .A(n12899), .ZN(n11404) );
  AND2_X1 U10018 ( .A1(n6437), .A2(n12899), .ZN(n10413) );
  NAND2_X1 U10019 ( .A1(n12310), .A2(n14195), .ZN(n14080) );
  NAND2_X1 U10020 ( .A1(n10417), .A2(n10420), .ZN(n8447) );
  OR2_X1 U10021 ( .A1(n13000), .A2(n12828), .ZN(n12956) );
  NAND2_X1 U10022 ( .A1(n13629), .A2(n15612), .ZN(n12613) );
  AND2_X1 U10023 ( .A1(n12540), .A2(n12533), .ZN(n12534) );
  INV_X1 U10024 ( .A(n15039), .ZN(n9881) );
  INV_X1 U10025 ( .A(n14756), .ZN(n15124) );
  OR2_X1 U10026 ( .A1(n10423), .A2(n8420), .ZN(n8451) );
  OR2_X1 U10027 ( .A1(n8253), .A2(SI_22_), .ZN(n8224) );
  NAND2_X1 U10028 ( .A1(n9881), .A2(n15282), .ZN(n9882) );
  INV_X1 U10029 ( .A(n13624), .ZN(n13571) );
  OR2_X1 U10030 ( .A1(n8516), .A2(n8448), .ZN(n8455) );
  INV_X1 U10031 ( .A(n12391), .ZN(n12546) );
  INV_X1 U10032 ( .A(n14910), .ZN(n15082) );
  AOI22_X2 U10033 ( .A1(n13100), .A2(n13101), .B1(n13416), .B2(n13044), .ZN(
        n13179) );
  NOR2_X2 U10034 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n7825) );
  AOI21_X1 U10035 ( .B1(n12536), .B2(n12384), .A(n12383), .ZN(n12385) );
  INV_X1 U10036 ( .A(n7779), .ZN(n15160) );
  OAI211_X2 U10037 ( .C1(n12223), .C2(n12222), .A(n14441), .B(n12221), .ZN(
        n14440) );
  AND2_X1 U10038 ( .A1(n10371), .A2(n8401), .ZN(n15311) );
  AND3_X1 U10039 ( .A1(n8429), .A2(n6510), .A3(n8416), .ZN(n8418) );
  NAND2_X1 U10040 ( .A1(n7890), .A2(n10075), .ZN(n11098) );
  NAND2_X1 U10041 ( .A1(n10474), .A2(n15292), .ZN(n9893) );
  AND2_X1 U10042 ( .A1(n12659), .A2(n14563), .ZN(n10096) );
  INV_X1 U10043 ( .A(n12659), .ZN(n14748) );
  INV_X1 U10044 ( .A(n7780), .ZN(n7778) );
  AND2_X1 U10045 ( .A1(n12548), .A2(n8993), .ZN(n7733) );
  NAND2_X1 U10046 ( .A1(n14335), .A2(n14392), .ZN(n14395) );
  INV_X1 U10047 ( .A(n13333), .ZN(n9642) );
  INV_X2 U10048 ( .A(n15561), .ZN(n15559) );
  OR2_X1 U10049 ( .A1(n9655), .A2(n13654), .ZN(n7734) );
  INV_X2 U10050 ( .A(n15598), .ZN(n15600) );
  AND2_X1 U10051 ( .A1(n9895), .A2(n9894), .ZN(n7735) );
  AND2_X1 U10052 ( .A1(n12933), .A2(n13862), .ZN(n7736) );
  INV_X1 U10053 ( .A(n10090), .ZN(n8313) );
  NAND2_X1 U10054 ( .A1(n8063), .A2(n7834), .ZN(n7737) );
  AND2_X1 U10055 ( .A1(n11953), .A2(n7773), .ZN(n7738) );
  NAND2_X1 U10056 ( .A1(n9643), .A2(n9642), .ZN(n7739) );
  AND2_X1 U10057 ( .A1(n11785), .A2(n9476), .ZN(n7741) );
  OR2_X1 U10058 ( .A1(n13997), .A2(n13791), .ZN(n7742) );
  INV_X1 U10059 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15151) );
  INV_X1 U10060 ( .A(n15552), .ZN(n15526) );
  XNOR2_X1 U10061 ( .A(n14100), .B(n13837), .ZN(n14101) );
  INV_X1 U10062 ( .A(SI_24_), .ZN(n12296) );
  INV_X1 U10063 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8895) );
  INV_X1 U10064 ( .A(n12711), .ZN(n8885) );
  AND2_X1 U10065 ( .A1(n13467), .A2(n13468), .ZN(n7743) );
  OR2_X1 U10066 ( .A1(n12449), .A2(n13157), .ZN(n7744) );
  AND3_X1 U10067 ( .A1(n12977), .A2(n12981), .A3(n12984), .ZN(n7745) );
  OR2_X1 U10068 ( .A1(n9655), .A2(n13598), .ZN(n7746) );
  NAND2_X1 U10069 ( .A1(n15612), .A2(n13595), .ZN(n13598) );
  INV_X1 U10070 ( .A(n13504), .ZN(n13473) );
  AND2_X1 U10071 ( .A1(n15050), .A2(n14542), .ZN(n7747) );
  OR2_X1 U10072 ( .A1(n15037), .A2(n15307), .ZN(n7748) );
  AND2_X1 U10073 ( .A1(n12621), .A2(n8886), .ZN(n7749) );
  AND2_X1 U10074 ( .A1(n9886), .A2(n9885), .ZN(n14988) );
  AND3_X2 U10075 ( .A1(n9782), .A2(n8914), .A3(n9794), .ZN(n15502) );
  INV_X1 U10076 ( .A(n15475), .ZN(n8826) );
  INV_X1 U10077 ( .A(n10066), .ZN(n9947) );
  NAND2_X1 U10078 ( .A1(n9948), .A2(n9947), .ZN(n9949) );
  AND2_X1 U10079 ( .A1(n9982), .A2(n9981), .ZN(n9983) );
  OR2_X1 U10080 ( .A1(n13213), .A2(n11328), .ZN(n8993) );
  OR2_X1 U10081 ( .A1(n13315), .A2(n13607), .ZN(n9633) );
  INV_X1 U10082 ( .A(n12542), .ZN(n9394) );
  INV_X1 U10083 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9409) );
  INV_X1 U10084 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8660) );
  NOR2_X1 U10085 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8820) );
  NAND2_X1 U10086 ( .A1(n14801), .A2(n14569), .ZN(n8351) );
  NOR2_X1 U10087 ( .A1(n7747), .A2(n8348), .ZN(n8349) );
  NAND2_X1 U10088 ( .A1(n10297), .A2(n10296), .ZN(n10299) );
  INV_X1 U10089 ( .A(n13546), .ZN(n12246) );
  INV_X1 U10090 ( .A(n13338), .ZN(n9634) );
  XNOR2_X1 U10091 ( .A(n13213), .B(n11328), .ZN(n12551) );
  OAI21_X1 U10092 ( .B1(n14108), .B2(n14104), .A(n14103), .ZN(n14105) );
  NOR2_X1 U10093 ( .A1(n8821), .A2(n8820), .ZN(n8822) );
  INV_X1 U10094 ( .A(n15466), .ZN(n12665) );
  INV_X1 U10095 ( .A(n14290), .ZN(n14291) );
  NAND2_X1 U10096 ( .A1(n14583), .A2(n14295), .ZN(n10804) );
  AOI211_X1 U10097 ( .C1(n10120), .C2(n10119), .A(n10118), .B(n10117), .ZN(
        n10134) );
  NAND2_X1 U10098 ( .A1(n14780), .A2(n14543), .ZN(n9838) );
  INV_X1 U10099 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n11921) );
  INV_X1 U10100 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7867) );
  OR2_X1 U10101 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14644), .ZN(n10969) );
  INV_X1 U10102 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9076) );
  INV_X1 U10103 ( .A(n11502), .ZN(n11499) );
  OR2_X1 U10104 ( .A1(n13315), .A2(n13527), .ZN(n9557) );
  INV_X1 U10105 ( .A(n13465), .ZN(n13470) );
  INV_X1 U10106 ( .A(SI_22_), .ZN(n9307) );
  INV_X1 U10107 ( .A(n9510), .ZN(n9517) );
  INV_X1 U10108 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9165) );
  INV_X1 U10109 ( .A(n11556), .ZN(n9687) );
  INV_X1 U10110 ( .A(n12979), .ZN(n12987) );
  INV_X1 U10111 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13110) );
  INV_X1 U10112 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U10113 ( .A1(n14292), .A2(n14291), .ZN(n14293) );
  NAND2_X1 U10114 ( .A1(n8305), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U10115 ( .A1(n7897), .A2(SI_4_), .ZN(n7895) );
  INV_X1 U10116 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U10117 ( .A1(n12250), .A2(n13546), .ZN(n12251) );
  OR2_X1 U10118 ( .A1(n13033), .A2(n13064), .ZN(n13034) );
  INV_X1 U10119 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8995) );
  NAND2_X1 U10120 ( .A1(n10911), .A2(n10910), .ZN(n10912) );
  NOR2_X1 U10121 ( .A1(n9563), .A2(n10846), .ZN(n12580) );
  INV_X1 U10122 ( .A(n9015), .ZN(n9075) );
  NAND2_X1 U10123 ( .A1(n9558), .A2(n9634), .ZN(n9559) );
  NAND2_X1 U10124 ( .A1(n11637), .A2(n12375), .ZN(n9274) );
  INV_X1 U10125 ( .A(n11153), .ZN(n12573) );
  OR2_X1 U10126 ( .A1(n9504), .A2(n15526), .ZN(n11782) );
  AND2_X1 U10127 ( .A1(n9514), .A2(n9419), .ZN(n13472) );
  INV_X1 U10128 ( .A(n12548), .ZN(n11159) );
  NAND2_X1 U10129 ( .A1(n13808), .A2(n7745), .ZN(n12991) );
  INV_X1 U10130 ( .A(n13855), .ZN(n12718) );
  INV_X1 U10131 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11270) );
  NOR3_X1 U10132 ( .A1(n15390), .A2(n15389), .A3(n15394), .ZN(n15391) );
  INV_X1 U10133 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n13777) );
  INV_X1 U10134 ( .A(n14101), .ZN(n12965) );
  INV_X1 U10135 ( .A(n14159), .ZN(n14028) );
  AND2_X1 U10136 ( .A1(n10420), .A2(n10413), .ZN(n13802) );
  INV_X1 U10137 ( .A(n13802), .ZN(n13814) );
  INV_X2 U10138 ( .A(n10193), .ZN(n10171) );
  XNOR2_X1 U10139 ( .A(n10805), .B(n14359), .ZN(n11113) );
  OR2_X1 U10140 ( .A1(n10395), .A2(n10389), .ZN(n10392) );
  OR2_X1 U10141 ( .A1(n14778), .A2(n9851), .ZN(n8312) );
  INV_X1 U10142 ( .A(n10087), .ZN(n14787) );
  INV_X1 U10143 ( .A(n15107), .ZN(n15003) );
  INV_X1 U10144 ( .A(n14579), .ZN(n11667) );
  OR2_X1 U10145 ( .A1(n14985), .A2(n15020), .ZN(n15022) );
  NAND2_X1 U10146 ( .A1(n10339), .A2(n10390), .ZN(n15032) );
  INV_X1 U10147 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7775) );
  OR2_X1 U10148 ( .A1(n8106), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n8130) );
  XNOR2_X1 U10149 ( .A(n8053), .B(SI_13_), .ZN(n8051) );
  NAND2_X1 U10150 ( .A1(n10965), .A2(n10964), .ZN(n10975) );
  INV_X1 U10151 ( .A(n11628), .ZN(n11627) );
  INV_X1 U10152 ( .A(n13193), .ZN(n13181) );
  INV_X1 U10153 ( .A(n13199), .ZN(n13169) );
  AND4_X1 U10154 ( .A1(n12371), .A2(n9817), .A3(n9816), .A4(n9815), .ZN(n12382) );
  AND2_X1 U10155 ( .A1(n9316), .A2(n9315), .ZN(n13429) );
  INV_X1 U10156 ( .A(n13157), .ZN(n12448) );
  INV_X1 U10157 ( .A(n13355), .ZN(n13339) );
  INV_X1 U10158 ( .A(n13629), .ZN(n9825) );
  NAND2_X1 U10159 ( .A1(n12573), .A2(n11640), .ZN(n15552) );
  NAND2_X1 U10160 ( .A1(n15609), .A2(n12611), .ZN(n12612) );
  INV_X1 U10161 ( .A(n13598), .ZN(n13617) );
  AND3_X1 U10162 ( .A1(n9511), .A2(n9462), .A3(n9518), .ZN(n9501) );
  INV_X1 U10163 ( .A(n12559), .ZN(n12113) );
  OR2_X1 U10164 ( .A1(n10872), .A2(n9519), .ZN(n9520) );
  INV_X1 U10165 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9417) );
  OR2_X1 U10166 ( .A1(n9184), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n9199) );
  OR2_X1 U10167 ( .A1(n9728), .A2(n9727), .ZN(n9735) );
  OR2_X1 U10168 ( .A1(n15472), .A2(n10413), .ZN(n9783) );
  INV_X1 U10169 ( .A(n15392), .ZN(n15419) );
  AND2_X1 U10170 ( .A1(n10418), .A2(n12903), .ZN(n15423) );
  INV_X1 U10171 ( .A(n13017), .ZN(n13916) );
  AND2_X1 U10172 ( .A1(n11560), .A2(n11562), .ZN(n11565) );
  NAND2_X1 U10173 ( .A1(n10993), .A2(n15434), .ZN(n14064) );
  NAND2_X1 U10174 ( .A1(n12905), .A2(n10413), .ZN(n9794) );
  AND2_X1 U10175 ( .A1(n8871), .A2(n12913), .ZN(n14186) );
  AND2_X1 U10176 ( .A1(n14072), .A2(n14222), .ZN(n15475) );
  AND2_X1 U10177 ( .A1(n9794), .A2(n9790), .ZN(n10992) );
  INV_X1 U10178 ( .A(n14555), .ZN(n14534) );
  INV_X1 U10179 ( .A(n14719), .ZN(n14737) );
  INV_X1 U10180 ( .A(n11646), .ZN(n14739) );
  INV_X1 U10181 ( .A(n14735), .ZN(n14733) );
  INV_X1 U10182 ( .A(n15032), .ZN(n15010) );
  NAND2_X1 U10183 ( .A1(n9862), .A2(n10260), .ZN(n14997) );
  INV_X1 U10184 ( .A(n15096), .ZN(n11749) );
  AND2_X1 U10185 ( .A1(n9861), .A2(n10374), .ZN(n8402) );
  AND3_X1 U10186 ( .A1(n9860), .A2(n10375), .A3(n10394), .ZN(n8403) );
  NAND2_X1 U10187 ( .A1(n10305), .A2(n10306), .ZN(n10957) );
  AND2_X1 U10188 ( .A1(n9612), .A2(n9611), .ZN(n15503) );
  INV_X1 U10189 ( .A(n13196), .ZN(n13177) );
  AND4_X1 U10190 ( .A1(n12371), .A2(n9429), .A3(n9428), .A4(n9427), .ZN(n13077) );
  INV_X1 U10191 ( .A(n13417), .ZN(n13447) );
  INV_X1 U10192 ( .A(n13192), .ZN(n13536) );
  OR2_X1 U10193 ( .A1(n9641), .A2(n9640), .ZN(n13333) );
  INV_X1 U10194 ( .A(n13270), .ZN(n13359) );
  AOI21_X1 U10195 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9836) );
  OR2_X1 U10196 ( .A1(n15561), .A2(n9503), .ZN(n13566) );
  OR2_X1 U10197 ( .A1(n15561), .A2(n11155), .ZN(n15555) );
  AND2_X1 U10198 ( .A1(n9504), .A2(n15553), .ZN(n15561) );
  NAND2_X1 U10199 ( .A1(n15612), .A2(n9524), .ZN(n13620) );
  INV_X1 U10200 ( .A(n15612), .ZN(n15609) );
  INV_X1 U10201 ( .A(n10152), .ZN(n10153) );
  OR2_X1 U10202 ( .A1(n15598), .A2(n9525), .ZN(n13695) );
  AND2_X1 U10203 ( .A1(n9521), .A2(n9520), .ZN(n15598) );
  NAND2_X1 U10204 ( .A1(n9447), .A2(n10310), .ZN(n10311) );
  INV_X1 U10205 ( .A(n10310), .ZN(n10270) );
  XNOR2_X1 U10206 ( .A(n9436), .B(n9435), .ZN(n12260) );
  INV_X1 U10207 ( .A(SI_9_), .ZN(n10191) );
  NAND2_X1 U10208 ( .A1(n9798), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15334) );
  OR2_X2 U10209 ( .A1(n9783), .A2(n9787), .ZN(n15327) );
  INV_X1 U10210 ( .A(n15332), .ZN(n13820) );
  INV_X1 U10211 ( .A(n12719), .ZN(n13850) );
  OR2_X1 U10212 ( .A1(n15361), .A2(P2_U3088), .ZN(n15408) );
  OR2_X1 U10213 ( .A1(n10428), .A2(P2_U3088), .ZN(n15427) );
  AND3_X1 U10214 ( .A1(n14078), .A2(n14077), .A3(n14076), .ZN(n14192) );
  INV_X1 U10215 ( .A(n15446), .ZN(n14056) );
  NAND2_X1 U10216 ( .A1(n8916), .A2(n15502), .ZN(n8913) );
  INV_X1 U10217 ( .A(n15502), .ZN(n15500) );
  NAND2_X1 U10218 ( .A1(n15459), .A2(n15449), .ZN(n15455) );
  AND2_X1 U10219 ( .A1(n9796), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15459) );
  XNOR2_X1 U10220 ( .A(n8890), .B(n8889), .ZN(n11795) );
  INV_X1 U10221 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11977) );
  INV_X1 U10222 ( .A(n15050), .ZN(n14810) );
  INV_X1 U10223 ( .A(n10393), .ZN(n14550) );
  OR2_X1 U10224 ( .A1(n15272), .A2(n15261), .ZN(n11646) );
  OR2_X1 U10225 ( .A1(n15272), .A2(n10339), .ZN(n14719) );
  OR2_X1 U10226 ( .A1(n15272), .A2(n10341), .ZN(n14735) );
  OR2_X1 U10227 ( .A1(n14965), .A2(n14964), .ZN(n15102) );
  INV_X1 U10228 ( .A(n15273), .ZN(n14984) );
  AND2_X1 U10229 ( .A1(n8403), .A2(n8399), .ZN(n15322) );
  INV_X1 U10230 ( .A(n14888), .ZN(n15135) );
  INV_X1 U10231 ( .A(n15319), .ZN(n15317) );
  INV_X1 U10232 ( .A(n10161), .ZN(n10257) );
  NAND2_X1 U10233 ( .A1(n8380), .A2(n8376), .ZN(n12154) );
  INV_X1 U10234 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11974) );
  INV_X1 U10235 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10466) );
  INV_X1 U10236 ( .A(n13214), .ZN(P3_U3897) );
  AND2_X1 U10237 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10415), .ZN(P2_U3947) );
  NOR2_X1 U10238 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n7752) );
  NOR2_X1 U10239 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n7754) );
  NOR2_X1 U10240 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7753) );
  INV_X1 U10241 ( .A(n7774), .ZN(n7757) );
  NAND2_X1 U10242 ( .A1(n7772), .A2(n11988), .ZN(n7759) );
  NAND2_X1 U10243 ( .A1(n7760), .A2(n7903), .ZN(n7766) );
  AND2_X1 U10244 ( .A1(n8398), .A2(n8371), .ZN(n7768) );
  NAND2_X2 U10245 ( .A1(n7765), .A2(n7764), .ZN(n15297) );
  NAND2_X1 U10246 ( .A1(n7766), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U10247 ( .A1(n10380), .A2(n8371), .ZN(n7769) );
  NOR2_X1 U10248 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n7771) );
  NOR2_X1 U10249 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n7770) );
  NAND2_X1 U10250 ( .A1(n7811), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U10251 ( .A1(n7835), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7783) );
  NAND2_X1 U10252 ( .A1(n7851), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7781) );
  INV_X1 U10253 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10194) );
  MUX2_X1 U10254 ( .A(n10194), .B(n10172), .S(n6439), .Z(n7789) );
  AND2_X1 U10255 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U10256 ( .A1(n10193), .A2(n7786), .ZN(n7808) );
  AND2_X1 U10257 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U10258 ( .A1(n7818), .A2(n7787), .ZN(n8445) );
  NAND2_X1 U10259 ( .A1(n7808), .A2(n8445), .ZN(n7821) );
  XNOR2_X1 U10260 ( .A(n7821), .B(SI_1_), .ZN(n7788) );
  XNOR2_X1 U10261 ( .A(n7789), .B(n7788), .ZN(n10195) );
  NAND2_X1 U10262 ( .A1(n10171), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7791) );
  OAI21_X1 U10263 ( .B1(n10195), .B2(n10171), .A(n7791), .ZN(n7795) );
  XNOR2_X2 U10264 ( .A(n7794), .B(n7793), .ZN(n7809) );
  INV_X1 U10265 ( .A(n7809), .ZN(n10339) );
  NAND2_X1 U10266 ( .A1(n7795), .A2(n10339), .ZN(n7802) );
  NAND2_X1 U10267 ( .A1(n10195), .A2(n10193), .ZN(n7798) );
  XNOR2_X2 U10268 ( .A(n7797), .B(n7796), .ZN(n10433) );
  INV_X1 U10269 ( .A(n10433), .ZN(n15261) );
  OAI211_X1 U10270 ( .C1(n10193), .C2(P2_DATAO_REG_1__SCAN_IN), .A(n7798), .B(
        n15261), .ZN(n7801) );
  INV_X1 U10271 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15264) );
  NAND2_X1 U10272 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n7799) );
  NAND3_X1 U10273 ( .A1(n7809), .A2(n14595), .A3(n10433), .ZN(n7800) );
  OR2_X1 U10274 ( .A1(n10474), .A2(n15292), .ZN(n8316) );
  NAND2_X1 U10275 ( .A1(n7811), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U10276 ( .A1(n7835), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7804) );
  NAND2_X1 U10277 ( .A1(n7833), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7803) );
  INV_X1 U10278 ( .A(SI_0_), .ZN(n10177) );
  INV_X1 U10279 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8950) );
  OAI21_X1 U10280 ( .B1(n10171), .B2(n10177), .A(n8950), .ZN(n7807) );
  NAND2_X1 U10281 ( .A1(n7808), .A2(n7807), .ZN(n15168) );
  INV_X1 U10282 ( .A(n10511), .ZN(n10399) );
  NAND2_X1 U10283 ( .A1(n14587), .A2(n10399), .ZN(n10516) );
  INV_X1 U10284 ( .A(n10516), .ZN(n7810) );
  INV_X1 U10285 ( .A(n15292), .ZN(n10521) );
  NAND2_X1 U10286 ( .A1(n7851), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U10287 ( .A1(n8063), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U10288 ( .A1(n7835), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U10289 ( .A1(n7811), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7812) );
  NAND4_X4 U10290 ( .A1(n7815), .A2(n7814), .A3(n7813), .A4(n7812), .ZN(n14585) );
  INV_X1 U10291 ( .A(SI_2_), .ZN(n10182) );
  XNOR2_X1 U10292 ( .A(n7839), .B(n10182), .ZN(n7843) );
  NAND2_X1 U10293 ( .A1(n7818), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7819) );
  INV_X1 U10294 ( .A(SI_1_), .ZN(n10176) );
  OAI211_X1 U10295 ( .C1(n6439), .C2(n10194), .A(n7819), .B(n10176), .ZN(n7820) );
  NAND2_X1 U10296 ( .A1(n7821), .A2(n7820), .ZN(n7824) );
  NAND2_X1 U10297 ( .A1(n6439), .A2(n10172), .ZN(n7822) );
  OAI211_X1 U10298 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n6439), .A(n7822), .B(
        SI_1_), .ZN(n7823) );
  NAND2_X1 U10299 ( .A1(n7824), .A2(n7823), .ZN(n7842) );
  XNOR2_X1 U10300 ( .A(n7843), .B(n7842), .ZN(n10278) );
  OR2_X1 U10301 ( .A1(n8262), .A2(n10278), .ZN(n7830) );
  INV_X1 U10302 ( .A(n7825), .ZN(n7826) );
  NAND2_X1 U10303 ( .A1(n7826), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7827) );
  INV_X1 U10304 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7844) );
  XNOR2_X1 U10305 ( .A(n7827), .B(n7844), .ZN(n10436) );
  OR2_X1 U10306 ( .A1(n7856), .A2(n10436), .ZN(n7829) );
  NAND2_X1 U10307 ( .A1(n7856), .A2(n10171), .ZN(n7868) );
  OR2_X1 U10308 ( .A1(n7868), .A2(n7817), .ZN(n7828) );
  XNOR2_X2 U10309 ( .A(n14585), .B(n10530), .ZN(n10548) );
  NAND2_X1 U10310 ( .A1(n10545), .A2(n10546), .ZN(n7832) );
  OR2_X1 U10311 ( .A1(n14585), .A2(n10530), .ZN(n7831) );
  BUF_X2 U10312 ( .A(n7833), .Z(n8063) );
  INV_X1 U10313 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U10314 ( .A1(n9866), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10315 ( .A1(n8173), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n7837) );
  INV_X1 U10316 ( .A(n7839), .ZN(n7840) );
  NOR2_X1 U10317 ( .A1(n7840), .A2(n10182), .ZN(n7841) );
  MUX2_X1 U10318 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7818), .Z(n7862) );
  XNOR2_X1 U10319 ( .A(n7862), .B(SI_3_), .ZN(n7864) );
  XNOR2_X1 U10320 ( .A(n7864), .B(n7865), .ZN(n10276) );
  NAND2_X1 U10321 ( .A1(n7825), .A2(n7844), .ZN(n7846) );
  NAND2_X1 U10322 ( .A1(n7846), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7845) );
  MUX2_X1 U10323 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7845), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n7847) );
  NAND2_X1 U10324 ( .A1(n7847), .A2(n7858), .ZN(n14606) );
  OR2_X1 U10325 ( .A1(n7856), .A2(n14606), .ZN(n7849) );
  INV_X1 U10326 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10250) );
  INV_X1 U10327 ( .A(n14584), .ZN(n10810) );
  NAND2_X1 U10328 ( .A1(n10810), .A2(n7686), .ZN(n7850) );
  NAND2_X1 U10329 ( .A1(n8173), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7854) );
  NAND2_X1 U10330 ( .A1(n7835), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7853) );
  NAND2_X1 U10331 ( .A1(n7851), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7852) );
  XNOR2_X1 U10332 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10902) );
  OR2_X1 U10333 ( .A1(n9851), .A2(n10902), .ZN(n7855) );
  NAND2_X1 U10334 ( .A1(n7858), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7857) );
  MUX2_X1 U10335 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7857), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n7861) );
  INV_X1 U10336 ( .A(n7858), .ZN(n7860) );
  INV_X1 U10337 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10338 ( .A1(n7860), .A2(n7859), .ZN(n7885) );
  NAND2_X1 U10339 ( .A1(n7861), .A2(n7885), .ZN(n14619) );
  NAND2_X1 U10340 ( .A1(n7862), .A2(SI_3_), .ZN(n7863) );
  NAND2_X1 U10341 ( .A1(n6439), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7866) );
  XNOR2_X1 U10342 ( .A(n7897), .B(SI_4_), .ZN(n7880) );
  NAND2_X1 U10343 ( .A1(n10197), .A2(n10061), .ZN(n7870) );
  INV_X1 U10344 ( .A(n11100), .ZN(n7890) );
  NAND2_X1 U10345 ( .A1(n8173), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7879) );
  INV_X1 U10346 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7872) );
  OR2_X1 U10347 ( .A1(n7871), .A2(n7872), .ZN(n7878) );
  NAND3_X2 U10348 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n7917) );
  INV_X1 U10349 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U10350 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7873) );
  NAND2_X1 U10351 ( .A1(n7874), .A2(n7873), .ZN(n7875) );
  NAND2_X1 U10352 ( .A1(n7917), .A2(n7875), .ZN(n11123) );
  OR2_X1 U10353 ( .A1(n9851), .A2(n11123), .ZN(n7877) );
  INV_X1 U10354 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10351) );
  OR2_X1 U10355 ( .A1(n10032), .A2(n10351), .ZN(n7876) );
  INV_X1 U10356 ( .A(n7880), .ZN(n7881) );
  NAND2_X1 U10357 ( .A1(n7882), .A2(n7895), .ZN(n7884) );
  MUX2_X1 U10358 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6439), .Z(n7898) );
  XNOR2_X1 U10359 ( .A(n7898), .B(SI_5_), .ZN(n7883) );
  NAND2_X1 U10360 ( .A1(n10238), .A2(n10061), .ZN(n7888) );
  NAND2_X1 U10361 ( .A1(n7885), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7886) );
  XNOR2_X1 U10362 ( .A(n7886), .B(P1_IR_REG_5__SCAN_IN), .ZN(n14635) );
  AOI22_X1 U10363 ( .A1(n8167), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8166), .B2(
        n14635), .ZN(n7887) );
  NAND2_X1 U10364 ( .A1(n11284), .A2(n11213), .ZN(n11280) );
  INV_X1 U10365 ( .A(n11284), .ZN(n14582) );
  NAND2_X1 U10366 ( .A1(n11120), .A2(n14582), .ZN(n7889) );
  NAND2_X1 U10367 ( .A1(n11280), .A2(n7889), .ZN(n10075) );
  INV_X1 U10368 ( .A(SI_4_), .ZN(n11991) );
  INV_X1 U10369 ( .A(n7897), .ZN(n7892) );
  INV_X1 U10370 ( .A(n7898), .ZN(n7891) );
  INV_X1 U10371 ( .A(SI_5_), .ZN(n7894) );
  AOI22_X1 U10372 ( .A1(n11991), .A2(n7892), .B1(n7891), .B2(n7894), .ZN(n7893) );
  NAND2_X1 U10373 ( .A1(n7895), .A2(n7894), .ZN(n7899) );
  AND2_X1 U10374 ( .A1(SI_4_), .A2(SI_5_), .ZN(n7896) );
  AOI22_X1 U10375 ( .A1(n7899), .A2(n7898), .B1(n7897), .B2(n7896), .ZN(n7956)
         );
  MUX2_X1 U10376 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n7818), .Z(n7900) );
  INV_X1 U10377 ( .A(n7907), .ZN(n7961) );
  NAND2_X1 U10378 ( .A1(n7908), .A2(n7961), .ZN(n7937) );
  NAND2_X1 U10379 ( .A1(n7900), .A2(SI_6_), .ZN(n7936) );
  NAND2_X1 U10380 ( .A1(n10246), .A2(n10061), .ZN(n7906) );
  INV_X1 U10381 ( .A(n7903), .ZN(n7911) );
  NAND2_X1 U10382 ( .A1(n7911), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7904) );
  XNOR2_X1 U10383 ( .A(n7904), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14664) );
  AOI22_X1 U10384 ( .A1(n8167), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8166), .B2(
        n14664), .ZN(n7905) );
  NAND2_X1 U10385 ( .A1(n10243), .A2(n10061), .ZN(n7914) );
  NAND2_X1 U10386 ( .A1(n7909), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7910) );
  MUX2_X1 U10387 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7910), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n7912) );
  AND2_X1 U10388 ( .A1(n7912), .A2(n7911), .ZN(n14648) );
  AOI22_X1 U10389 ( .A1(n8167), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8166), .B2(
        n14648), .ZN(n7913) );
  NAND2_X1 U10390 ( .A1(n8173), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7922) );
  INV_X1 U10391 ( .A(n7917), .ZN(n7915) );
  INV_X1 U10392 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10393 ( .A1(n7917), .A2(n7916), .ZN(n7918) );
  NAND2_X1 U10394 ( .A1(n7925), .A2(n7918), .ZN(n11427) );
  OR2_X1 U10395 ( .A1(n9851), .A2(n11427), .ZN(n7921) );
  NAND2_X1 U10396 ( .A1(n9866), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10397 ( .A1(n7835), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7919) );
  INV_X1 U10398 ( .A(n14581), .ZN(n11220) );
  NAND2_X1 U10399 ( .A1(n8173), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7930) );
  INV_X1 U10400 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U10401 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  NAND2_X1 U10402 ( .A1(n7947), .A2(n7926), .ZN(n11594) );
  OR2_X1 U10403 ( .A1(n9851), .A2(n11594), .ZN(n7929) );
  NAND2_X1 U10404 ( .A1(n9866), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7928) );
  NAND2_X1 U10405 ( .A1(n7835), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7927) );
  NAND4_X1 U10406 ( .A1(n7930), .A2(n7929), .A3(n7928), .A4(n7927), .ZN(n14579) );
  NAND3_X1 U10407 ( .A1(n11291), .A2(n11220), .A3(n11667), .ZN(n7932) );
  NAND2_X1 U10408 ( .A1(n7933), .A2(n7932), .ZN(n11710) );
  AND2_X1 U10409 ( .A1(n11284), .A2(n11120), .ZN(n11276) );
  NOR2_X1 U10410 ( .A1(n11710), .A2(n11276), .ZN(n7934) );
  NAND2_X1 U10411 ( .A1(n11098), .A2(n7934), .ZN(n7955) );
  AOI22_X1 U10412 ( .A1(n11596), .A2(n14579), .B1(n11429), .B2(n14581), .ZN(
        n11709) );
  NAND2_X1 U10413 ( .A1(n7935), .A2(SI_7_), .ZN(n7938) );
  NAND2_X1 U10414 ( .A1(n7937), .A2(n7960), .ZN(n7940) );
  MUX2_X1 U10415 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6439), .Z(n7966) );
  XNOR2_X1 U10416 ( .A(n7966), .B(SI_8_), .ZN(n7957) );
  NAND2_X1 U10417 ( .A1(n10265), .A2(n10061), .ZN(n7944) );
  NAND2_X1 U10418 ( .A1(n7903), .A2(n11921), .ZN(n7970) );
  NAND2_X1 U10419 ( .A1(n7970), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7942) );
  XNOR2_X1 U10420 ( .A(n7942), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U10421 ( .A1(n8167), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8166), .B2(
        n10605), .ZN(n7943) );
  NAND2_X2 U10422 ( .A1(n7944), .A2(n7943), .ZN(n11723) );
  INV_X1 U10423 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7946) );
  NAND2_X1 U10424 ( .A1(n7947), .A2(n7946), .ZN(n7948) );
  NAND2_X1 U10425 ( .A1(n7978), .A2(n7948), .ZN(n15275) );
  OR2_X1 U10426 ( .A1(n9851), .A2(n15275), .ZN(n7952) );
  NAND2_X1 U10427 ( .A1(n9866), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U10428 ( .A1(n7835), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10429 ( .A1(n8173), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7949) );
  NAND4_X1 U10430 ( .A1(n7952), .A2(n7951), .A3(n7950), .A4(n7949), .ZN(n14578) );
  OAI21_X1 U10431 ( .B1(n11710), .B2(n11709), .A(n11719), .ZN(n7953) );
  OR2_X1 U10432 ( .A1(n11723), .A2(n14578), .ZN(n11740) );
  NAND2_X1 U10433 ( .A1(n11714), .A2(n11740), .ZN(n7985) );
  INV_X1 U10434 ( .A(n7957), .ZN(n7959) );
  AND2_X1 U10435 ( .A1(n7959), .A2(n7958), .ZN(n7964) );
  OR2_X1 U10436 ( .A1(n7962), .A2(n7961), .ZN(n7963) );
  NAND2_X1 U10437 ( .A1(n7966), .A2(SI_8_), .ZN(n7967) );
  MUX2_X1 U10438 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10039), .Z(n7987) );
  XNOR2_X1 U10439 ( .A(n7987), .B(SI_9_), .ZN(n7969) );
  XNOR2_X1 U10440 ( .A(n7991), .B(n7969), .ZN(n10241) );
  NAND2_X1 U10441 ( .A1(n10241), .A2(n10061), .ZN(n7975) );
  INV_X1 U10442 ( .A(n7970), .ZN(n7972) );
  INV_X1 U10443 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n7971) );
  NAND2_X1 U10444 ( .A1(n7972), .A2(n7971), .ZN(n7992) );
  NAND2_X1 U10445 ( .A1(n7992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7973) );
  XNOR2_X1 U10446 ( .A(n7973), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14680) );
  AOI22_X1 U10447 ( .A1(n8167), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8166), .B2(
        n14680), .ZN(n7974) );
  NAND2_X1 U10448 ( .A1(n8173), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7983) );
  INV_X1 U10449 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U10450 ( .A1(n7978), .A2(n7977), .ZN(n7979) );
  NAND2_X1 U10451 ( .A1(n7997), .A2(n7979), .ZN(n12040) );
  OR2_X1 U10452 ( .A1(n9851), .A2(n12040), .ZN(n7982) );
  NAND2_X1 U10453 ( .A1(n9866), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7981) );
  NAND2_X1 U10454 ( .A1(n7835), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7980) );
  NAND4_X1 U10455 ( .A1(n7983), .A2(n7982), .A3(n7981), .A4(n7980), .ZN(n14577) );
  OR2_X1 U10456 ( .A1(n12044), .A2(n14577), .ZN(n7986) );
  NAND2_X1 U10457 ( .A1(n12044), .A2(n14577), .ZN(n7984) );
  NAND2_X1 U10458 ( .A1(n7986), .A2(n7984), .ZN(n11741) );
  INV_X1 U10459 ( .A(n11741), .ZN(n11737) );
  NOR2_X1 U10460 ( .A1(n7988), .A2(n10191), .ZN(n7990) );
  NAND2_X1 U10461 ( .A1(n7988), .A2(n10191), .ZN(n7989) );
  XNOR2_X1 U10462 ( .A(n8006), .B(n7467), .ZN(n10272) );
  NAND2_X1 U10463 ( .A1(n10272), .A2(n10061), .ZN(n7995) );
  NAND2_X1 U10464 ( .A1(n8007), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7993) );
  XNOR2_X1 U10465 ( .A(n7993), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U10466 ( .A1(n8167), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8166), 
        .B2(n10649), .ZN(n7994) );
  NAND2_X1 U10467 ( .A1(n9866), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U10468 ( .A1(n7997), .A2(n7996), .ZN(n7998) );
  NAND2_X1 U10469 ( .A1(n8012), .A2(n7998), .ZN(n12289) );
  OR2_X1 U10470 ( .A1(n9851), .A2(n12289), .ZN(n8001) );
  NAND2_X1 U10471 ( .A1(n8173), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10472 ( .A1(n7835), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7999) );
  NAND4_X1 U10473 ( .A1(n8002), .A2(n8001), .A3(n8000), .A4(n7999), .ZN(n14576) );
  OR2_X1 U10474 ( .A1(n12160), .A2(n14576), .ZN(n8003) );
  MUX2_X1 U10475 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10039), .Z(n8019) );
  NAND2_X1 U10476 ( .A1(n10313), .A2(n10061), .ZN(n8011) );
  INV_X1 U10477 ( .A(n8007), .ZN(n8008) );
  NAND2_X1 U10478 ( .A1(n8008), .A2(n11911), .ZN(n8024) );
  NAND2_X1 U10479 ( .A1(n8024), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8009) );
  XNOR2_X1 U10480 ( .A(n8009), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U10481 ( .A1(n8167), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8166), 
        .B2(n10720), .ZN(n8010) );
  NAND2_X1 U10482 ( .A1(n9866), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8017) );
  NAND2_X1 U10483 ( .A1(n8012), .A2(n10657), .ZN(n8013) );
  NAND2_X1 U10484 ( .A1(n8029), .A2(n8013), .ZN(n14520) );
  OR2_X1 U10485 ( .A1(n9851), .A2(n14520), .ZN(n8016) );
  NAND2_X1 U10486 ( .A1(n7835), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U10487 ( .A1(n10029), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8014) );
  NAND4_X1 U10488 ( .A1(n8017), .A2(n8016), .A3(n8015), .A4(n8014), .ZN(n14575) );
  OR2_X1 U10489 ( .A1(n15117), .A2(n14575), .ZN(n8018) );
  INV_X1 U10490 ( .A(n8019), .ZN(n8020) );
  NAND2_X1 U10491 ( .A1(n8020), .A2(n10248), .ZN(n8021) );
  MUX2_X1 U10492 ( .A(n10408), .B(n10406), .S(n10039), .Z(n8038) );
  XNOR2_X1 U10493 ( .A(n8038), .B(SI_12_), .ZN(n8036) );
  XNOR2_X1 U10494 ( .A(n8037), .B(n8036), .ZN(n10405) );
  NAND2_X1 U10495 ( .A1(n10405), .A2(n10061), .ZN(n8027) );
  NAND2_X1 U10496 ( .A1(n8025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8039) );
  XNOR2_X1 U10497 ( .A(n8039), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U10498 ( .A1(n8167), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11006), 
        .B2(n8166), .ZN(n8026) );
  INV_X1 U10499 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U10500 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  NAND2_X1 U10501 ( .A1(n8045), .A2(n8030), .ZN(n14443) );
  OR2_X1 U10502 ( .A1(n9851), .A2(n14443), .ZN(n8034) );
  INV_X1 U10503 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11843) );
  OR2_X1 U10504 ( .A1(n10032), .A2(n11843), .ZN(n8033) );
  NAND2_X1 U10505 ( .A1(n9866), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10506 ( .A1(n10029), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8031) );
  NAND4_X1 U10507 ( .A1(n8034), .A2(n8033), .A3(n8032), .A4(n8031), .ZN(n14574) );
  INV_X1 U10508 ( .A(n14574), .ZN(n8331) );
  XNOR2_X1 U10509 ( .A(n12205), .B(n8331), .ZN(n10080) );
  OR2_X1 U10510 ( .A1(n12205), .A2(n14574), .ZN(n8035) );
  MUX2_X1 U10511 ( .A(n10466), .B(n7541), .S(n10039), .Z(n8053) );
  XNOR2_X1 U10512 ( .A(n8052), .B(n8051), .ZN(n10463) );
  NAND2_X1 U10513 ( .A1(n10463), .A2(n10061), .ZN(n8042) );
  NAND2_X1 U10514 ( .A1(n8039), .A2(n11887), .ZN(n8040) );
  NAND2_X1 U10515 ( .A1(n8040), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8058) );
  XNOR2_X1 U10516 ( .A(n8058), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U10517 ( .A1(n11520), .A2(n8166), .B1(n8167), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8041) );
  NAND2_X1 U10518 ( .A1(n9866), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8050) );
  INV_X1 U10519 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11805) );
  OR2_X1 U10520 ( .A1(n10032), .A2(n11805), .ZN(n8049) );
  INV_X1 U10521 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8044) );
  NAND2_X1 U10522 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  NAND2_X1 U10523 ( .A1(n8065), .A2(n8046), .ZN(n12234) );
  OR2_X1 U10524 ( .A1(n9851), .A2(n12234), .ZN(n8048) );
  INV_X1 U10525 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n12302) );
  OR2_X1 U10526 ( .A1(n7836), .A2(n12302), .ZN(n8047) );
  XNOR2_X1 U10527 ( .A(n12236), .B(n15011), .ZN(n10081) );
  NAND2_X1 U10528 ( .A1(n8053), .A2(n10402), .ZN(n8054) );
  NAND2_X1 U10529 ( .A1(n8120), .A2(n10469), .ZN(n8055) );
  OAI21_X1 U10530 ( .B1(n8120), .B2(n10469), .A(n8055), .ZN(n8056) );
  MUX2_X1 U10531 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10039), .Z(n8072) );
  XNOR2_X1 U10532 ( .A(n8056), .B(n8072), .ZN(n10765) );
  NAND2_X1 U10533 ( .A1(n10765), .A2(n10061), .ZN(n8062) );
  INV_X1 U10534 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10535 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  NAND2_X1 U10536 ( .A1(n8059), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8060) );
  AOI22_X1 U10537 ( .A1(n14698), .A2(n8166), .B1(n8167), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U10538 ( .A1(n8065), .A2(n8064), .ZN(n8066) );
  AND2_X1 U10539 ( .A1(n8090), .A2(n8066), .ZN(n15017) );
  NAND2_X1 U10540 ( .A1(n8063), .A2(n15017), .ZN(n8071) );
  INV_X1 U10541 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8067) );
  OR2_X1 U10542 ( .A1(n7836), .A2(n8067), .ZN(n8070) );
  INV_X1 U10543 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11512) );
  OR2_X1 U10544 ( .A1(n7871), .A2(n11512), .ZN(n8069) );
  INV_X1 U10545 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11521) );
  OR2_X1 U10546 ( .A1(n10032), .A2(n11521), .ZN(n8068) );
  NAND2_X1 U10547 ( .A1(n15112), .A2(n14573), .ZN(n14986) );
  MUX2_X1 U10548 ( .A(n10704), .B(n11976), .S(n10171), .Z(n8097) );
  XNOR2_X1 U10549 ( .A(n8097), .B(SI_15_), .ZN(n8074) );
  NOR2_X1 U10550 ( .A1(n8076), .A2(n8119), .ZN(n8079) );
  INV_X1 U10551 ( .A(n8072), .ZN(n8073) );
  NOR2_X1 U10552 ( .A1(n8074), .A2(n8075), .ZN(n8078) );
  NAND2_X1 U10553 ( .A1(n8120), .A2(n8121), .ZN(n8077) );
  NAND2_X1 U10554 ( .A1(n10703), .A2(n10061), .ZN(n8087) );
  INV_X1 U10555 ( .A(n8080), .ZN(n8083) );
  INV_X1 U10556 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8081) );
  NAND4_X1 U10557 ( .A1(n11887), .A2(n11911), .A3(n8081), .A4(n11921), .ZN(
        n8082) );
  NOR2_X1 U10558 ( .A1(n8083), .A2(n8082), .ZN(n8084) );
  NAND2_X1 U10559 ( .A1(n7903), .A2(n8084), .ZN(n8102) );
  NAND2_X1 U10560 ( .A1(n8102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8085) );
  XNOR2_X1 U10561 ( .A(n8085), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U10562 ( .A1(n8167), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8166), 
        .B2(n11525), .ZN(n8086) );
  INV_X1 U10563 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U10564 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  NAND2_X1 U10565 ( .A1(n8110), .A2(n8091), .ZN(n14998) );
  OR2_X1 U10566 ( .A1(n14998), .A2(n9851), .ZN(n8095) );
  NAND2_X1 U10567 ( .A1(n8173), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10568 ( .A1(n9866), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U10569 ( .A1(n7835), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8092) );
  NAND4_X1 U10570 ( .A1(n8095), .A2(n8094), .A3(n8093), .A4(n8092), .ZN(n15009) );
  NAND2_X1 U10571 ( .A1(n15107), .A2(n14966), .ZN(n9954) );
  AND2_X1 U10572 ( .A1(n14986), .A2(n14989), .ZN(n8096) );
  NAND2_X1 U10573 ( .A1(n14985), .A2(n8096), .ZN(n14968) );
  OAI21_X1 U10574 ( .B1(n8120), .B2(n8119), .A(n8121), .ZN(n8099) );
  INV_X1 U10575 ( .A(n8097), .ZN(n8098) );
  NAND2_X1 U10576 ( .A1(n8099), .A2(n6558), .ZN(n8101) );
  MUX2_X1 U10577 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n10171), .Z(n8125) );
  XNOR2_X1 U10578 ( .A(n8125), .B(SI_16_), .ZN(n8122) );
  INV_X1 U10579 ( .A(n8122), .ZN(n8100) );
  NAND2_X1 U10580 ( .A1(n10751), .A2(n10061), .ZN(n8109) );
  INV_X1 U10581 ( .A(n8102), .ZN(n8104) );
  INV_X1 U10582 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U10583 ( .A1(n8104), .A2(n8103), .ZN(n8106) );
  NAND2_X1 U10584 ( .A1(n8106), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8105) );
  MUX2_X1 U10585 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8105), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8107) );
  AOI22_X1 U10586 ( .A1(n8167), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8166), 
        .B2(n12087), .ZN(n8108) );
  INV_X1 U10587 ( .A(n8134), .ZN(n8136) );
  NAND2_X1 U10588 ( .A1(n8110), .A2(n6870), .ZN(n8111) );
  AND2_X1 U10589 ( .A1(n8136), .A2(n8111), .ZN(n14469) );
  NAND2_X1 U10590 ( .A1(n14469), .A2(n8063), .ZN(n8114) );
  AOI22_X1 U10591 ( .A1(n9866), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8173), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10592 ( .A1(n7835), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8112) );
  INV_X1 U10593 ( .A(n15112), .ZN(n15019) );
  NAND2_X1 U10594 ( .A1(n15003), .A2(n14966), .ZN(n8116) );
  NAND2_X1 U10595 ( .A1(n8117), .A2(n8116), .ZN(n14969) );
  AOI22_X1 U10596 ( .A1(n10083), .A2(n14969), .B1(n15105), .B2(n14994), .ZN(
        n8118) );
  INV_X1 U10597 ( .A(n8121), .ZN(n8123) );
  INV_X1 U10598 ( .A(n8125), .ZN(n8127) );
  INV_X1 U10599 ( .A(SI_16_), .ZN(n8126) );
  NAND2_X1 U10600 ( .A1(n8127), .A2(n8126), .ZN(n8128) );
  MUX2_X1 U10601 ( .A(n10956), .B(n11977), .S(n10171), .Z(n8145) );
  XNOR2_X1 U10602 ( .A(n8144), .B(n8143), .ZN(n10953) );
  NAND2_X1 U10603 ( .A1(n10953), .A2(n10061), .ZN(n8133) );
  NAND2_X1 U10604 ( .A1(n8130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8131) );
  XNOR2_X1 U10605 ( .A(n8131), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14707) );
  AOI22_X1 U10606 ( .A1(n8167), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8166), 
        .B2(n14707), .ZN(n8132) );
  INV_X1 U10607 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U10608 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  NAND2_X1 U10609 ( .A1(n8155), .A2(n8137), .ZN(n14956) );
  OR2_X1 U10610 ( .A1(n14956), .A2(n9851), .ZN(n8140) );
  AOI22_X1 U10611 ( .A1(n7835), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9866), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n8139) );
  NAND2_X1 U10612 ( .A1(n10029), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8138) );
  OR2_X1 U10613 ( .A1(n15099), .A2(n14572), .ZN(n9972) );
  INV_X1 U10614 ( .A(n9972), .ZN(n8141) );
  AND2_X1 U10615 ( .A1(n15099), .A2(n14572), .ZN(n9966) );
  INV_X1 U10616 ( .A(n9966), .ZN(n8142) );
  OR2_X1 U10617 ( .A1(n8190), .A2(n11090), .ZN(n8163) );
  NAND2_X1 U10618 ( .A1(n8190), .A2(n11090), .ZN(n8146) );
  MUX2_X1 U10619 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10039), .Z(n8186) );
  NAND2_X1 U10620 ( .A1(n8147), .A2(n8186), .ZN(n8164) );
  INV_X1 U10621 ( .A(n8147), .ZN(n8148) );
  INV_X1 U10622 ( .A(n8186), .ZN(n8187) );
  NAND2_X1 U10623 ( .A1(n8148), .A2(n8187), .ZN(n8149) );
  NAND2_X1 U10624 ( .A1(n8164), .A2(n8149), .ZN(n11131) );
  OR2_X1 U10625 ( .A1(n11131), .A2(n8262), .ZN(n8153) );
  INV_X1 U10626 ( .A(n8374), .ZN(n8150) );
  NAND2_X1 U10627 ( .A1(n8150), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8151) );
  XNOR2_X1 U10628 ( .A(n8151), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14727) );
  AOI22_X1 U10629 ( .A1(n8167), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8166), 
        .B2(n14727), .ZN(n8152) );
  INV_X1 U10630 ( .A(n15144), .ZN(n14940) );
  INV_X1 U10631 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U10632 ( .A1(n8155), .A2(n8154), .ZN(n8156) );
  AND2_X1 U10633 ( .A1(n8171), .A2(n8156), .ZN(n14941) );
  NAND2_X1 U10634 ( .A1(n14941), .A2(n8063), .ZN(n8162) );
  INV_X1 U10635 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10636 ( .A1(n8173), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U10637 ( .A1(n9866), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8157) );
  OAI211_X1 U10638 ( .C1(n8159), .C2(n10032), .A(n8158), .B(n8157), .ZN(n8160)
         );
  INV_X1 U10639 ( .A(n8160), .ZN(n8161) );
  NAND2_X1 U10640 ( .A1(n14940), .A2(n14950), .ZN(n9964) );
  NAND2_X1 U10641 ( .A1(n15144), .A2(n14407), .ZN(n9965) );
  NAND2_X1 U10642 ( .A1(n8164), .A2(n8163), .ZN(n8165) );
  MUX2_X1 U10643 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10039), .Z(n8191) );
  XNOR2_X1 U10644 ( .A(n8191), .B(SI_19_), .ZN(n8189) );
  XNOR2_X1 U10645 ( .A(n8165), .B(n8189), .ZN(n11423) );
  NAND2_X1 U10646 ( .A1(n11423), .A2(n10061), .ZN(n8169) );
  AOI22_X1 U10647 ( .A1(n8167), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8166), 
        .B2(n15296), .ZN(n8168) );
  INV_X1 U10648 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U10649 ( .A1(n8171), .A2(n8170), .ZN(n8172) );
  NAND2_X1 U10650 ( .A1(n8212), .A2(n8172), .ZN(n14919) );
  OR2_X1 U10651 ( .A1(n14919), .A2(n9851), .ZN(n8178) );
  INV_X1 U10652 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n12006) );
  NAND2_X1 U10653 ( .A1(n7835), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U10654 ( .A1(n8173), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8174) );
  OAI211_X1 U10655 ( .C1(n7871), .C2(n12006), .A(n8175), .B(n8174), .ZN(n8176)
         );
  INV_X1 U10656 ( .A(n8176), .ZN(n8177) );
  XNOR2_X1 U10657 ( .A(n15088), .B(n14900), .ZN(n14924) );
  INV_X1 U10658 ( .A(n14924), .ZN(n8340) );
  OR2_X1 U10659 ( .A1(n15088), .A2(n14900), .ZN(n8179) );
  INV_X1 U10660 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14496) );
  INV_X1 U10661 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14429) );
  OAI21_X1 U10662 ( .B1(n8212), .B2(n14496), .A(n14429), .ZN(n8180) );
  OR3_X2 U10663 ( .A1(n8212), .A2(n14496), .A3(n14429), .ZN(n8226) );
  NAND2_X1 U10664 ( .A1(n8180), .A2(n8226), .ZN(n14883) );
  OR2_X1 U10665 ( .A1(n14883), .A2(n9851), .ZN(n8185) );
  INV_X1 U10666 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14882) );
  NAND2_X1 U10667 ( .A1(n10029), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U10668 ( .A1(n9866), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8181) );
  OAI211_X1 U10669 ( .C1(n14882), .C2(n10032), .A(n8182), .B(n8181), .ZN(n8183) );
  INV_X1 U10670 ( .A(n8183), .ZN(n8184) );
  NOR2_X1 U10671 ( .A1(n8187), .A2(n11090), .ZN(n8188) );
  INV_X1 U10672 ( .A(n8191), .ZN(n8192) );
  INV_X1 U10673 ( .A(SI_20_), .ZN(n11639) );
  OR2_X1 U10674 ( .A1(n8198), .A2(n11639), .ZN(n8195) );
  NAND2_X1 U10675 ( .A1(n8198), .A2(n11639), .ZN(n8193) );
  NAND2_X1 U10676 ( .A1(n8195), .A2(n8193), .ZN(n8207) );
  MUX2_X1 U10677 ( .A(n11380), .B(n11383), .S(n10039), .Z(n8206) );
  OR2_X1 U10678 ( .A1(n8207), .A2(n8206), .ZN(n8209) );
  MUX2_X1 U10679 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10171), .Z(n8194) );
  OAI21_X1 U10680 ( .B1(n8194), .B2(SI_21_), .A(n8222), .ZN(n8201) );
  AND2_X1 U10681 ( .A1(n8195), .A2(n8201), .ZN(n8196) );
  NAND2_X1 U10682 ( .A1(n8209), .A2(n8196), .ZN(n8203) );
  NAND2_X1 U10683 ( .A1(n8199), .A2(SI_20_), .ZN(n8197) );
  NOR2_X1 U10684 ( .A1(n8199), .A2(SI_20_), .ZN(n8200) );
  NOR2_X1 U10685 ( .A1(n8201), .A2(n8200), .ZN(n8202) );
  NAND2_X1 U10686 ( .A1(n8203), .A2(n8223), .ZN(n11407) );
  OR2_X1 U10687 ( .A1(n11407), .A2(n8262), .ZN(n8205) );
  INV_X1 U10688 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11406) );
  NAND2_X1 U10689 ( .A1(n8207), .A2(n8206), .ZN(n8208) );
  OR2_X1 U10690 ( .A1(n11382), .A2(n8262), .ZN(n8211) );
  XNOR2_X1 U10691 ( .A(n8212), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n14497) );
  NAND2_X1 U10692 ( .A1(n14497), .A2(n8063), .ZN(n8217) );
  INV_X1 U10693 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14904) );
  NAND2_X1 U10694 ( .A1(n10029), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U10695 ( .A1(n9866), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8213) );
  OAI211_X1 U10696 ( .C1(n14904), .C2(n10032), .A(n8214), .B(n8213), .ZN(n8215) );
  INV_X1 U10697 ( .A(n8215), .ZN(n8216) );
  NAND2_X1 U10698 ( .A1(n8217), .A2(n8216), .ZN(n14878) );
  NAND2_X1 U10699 ( .A1(n15082), .A2(n14878), .ZN(n14873) );
  INV_X1 U10700 ( .A(n14878), .ZN(n14431) );
  NAND2_X1 U10701 ( .A1(n14910), .A2(n14431), .ZN(n8341) );
  OAI21_X1 U10702 ( .B1(n14901), .B2(n14888), .A(n14896), .ZN(n8221) );
  NAND2_X1 U10703 ( .A1(n14910), .A2(n14878), .ZN(n14891) );
  INV_X1 U10704 ( .A(n14901), .ZN(n14507) );
  NAND2_X1 U10705 ( .A1(n14891), .A2(n14507), .ZN(n8219) );
  INV_X1 U10706 ( .A(n14891), .ZN(n8218) );
  AOI22_X1 U10707 ( .A1(n14888), .A2(n8219), .B1(n8218), .B2(n14901), .ZN(
        n8220) );
  NAND2_X1 U10708 ( .A1(n8253), .A2(SI_22_), .ZN(n8235) );
  NAND2_X1 U10709 ( .A1(n8235), .A2(n8224), .ZN(n8734) );
  OR2_X1 U10710 ( .A1(n8734), .A2(n10039), .ZN(n8225) );
  XNOR2_X1 U10711 ( .A(n8225), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15167) );
  OR2_X2 U10712 ( .A1(n8226), .A2(n14509), .ZN(n8242) );
  NAND2_X1 U10713 ( .A1(n8226), .A2(n14509), .ZN(n8227) );
  AND2_X1 U10714 ( .A1(n8242), .A2(n8227), .ZN(n14865) );
  NAND2_X1 U10715 ( .A1(n14865), .A2(n8063), .ZN(n8233) );
  INV_X1 U10716 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8230) );
  NAND2_X1 U10717 ( .A1(n10029), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8229) );
  NAND2_X1 U10718 ( .A1(n9866), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8228) );
  OAI211_X1 U10719 ( .C1(n8230), .C2(n10032), .A(n8229), .B(n8228), .ZN(n8231)
         );
  INV_X1 U10720 ( .A(n8231), .ZN(n8232) );
  XNOR2_X1 U10721 ( .A(n14867), .B(n14879), .ZN(n14869) );
  INV_X1 U10722 ( .A(n14869), .ZN(n8234) );
  MUX2_X1 U10723 ( .A(n11951), .B(n11511), .S(n10171), .Z(n8733) );
  OR2_X1 U10724 ( .A1(n8734), .A2(n8733), .ZN(n8736) );
  NAND2_X1 U10725 ( .A1(n8736), .A2(n8235), .ZN(n8237) );
  MUX2_X1 U10726 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10039), .Z(n8254) );
  XNOR2_X1 U10727 ( .A(n8254), .B(SI_23_), .ZN(n8236) );
  NAND2_X1 U10728 ( .A1(n11733), .A2(n10061), .ZN(n8239) );
  INV_X1 U10729 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11736) );
  INV_X1 U10730 ( .A(n8242), .ZN(n8240) );
  INV_X1 U10731 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U10732 ( .A1(n8242), .A2(n8241), .ZN(n8243) );
  NAND2_X1 U10733 ( .A1(n8265), .A2(n8243), .ZN(n14843) );
  INV_X1 U10734 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14842) );
  NAND2_X1 U10735 ( .A1(n10029), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U10736 ( .A1(n9866), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8244) );
  OAI211_X1 U10737 ( .C1(n14842), .C2(n10032), .A(n8245), .B(n8244), .ZN(n8246) );
  INV_X1 U10738 ( .A(n8246), .ZN(n8247) );
  XNOR2_X1 U10739 ( .A(n15061), .B(n14571), .ZN(n14849) );
  INV_X1 U10740 ( .A(n14849), .ZN(n8249) );
  NAND2_X1 U10741 ( .A1(n15061), .A2(n14571), .ZN(n8250) );
  INV_X1 U10742 ( .A(n8254), .ZN(n8251) );
  INV_X1 U10743 ( .A(SI_23_), .ZN(n11636) );
  OAI22_X1 U10744 ( .A1(n8733), .A2(n9307), .B1(n8251), .B2(n11636), .ZN(n8252) );
  INV_X1 U10745 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11797) );
  INV_X1 U10746 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11794) );
  MUX2_X1 U10747 ( .A(n11797), .B(n11794), .S(n10171), .Z(n8259) );
  NAND2_X1 U10748 ( .A1(n8260), .A2(n8259), .ZN(n8261) );
  NAND2_X1 U10749 ( .A1(n8273), .A2(n8261), .ZN(n11798) );
  OR2_X1 U10750 ( .A1(n11798), .A2(n8262), .ZN(n8264) );
  INV_X1 U10751 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14489) );
  OR2_X2 U10752 ( .A1(n8265), .A2(n14489), .ZN(n8292) );
  NAND2_X1 U10753 ( .A1(n8265), .A2(n14489), .ZN(n8266) );
  INV_X1 U10754 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n14830) );
  NAND2_X1 U10755 ( .A1(n10029), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U10756 ( .A1(n9866), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8267) );
  OAI211_X1 U10757 ( .C1(n14830), .C2(n10032), .A(n8268), .B(n8267), .ZN(n8269) );
  INV_X1 U10758 ( .A(n8269), .ZN(n8270) );
  NAND2_X1 U10759 ( .A1(n15057), .A2(n14570), .ZN(n8350) );
  INV_X1 U10760 ( .A(n14570), .ZN(n14454) );
  NAND2_X1 U10761 ( .A1(n14833), .A2(n14454), .ZN(n8347) );
  INV_X1 U10762 ( .A(n14817), .ZN(n14824) );
  MUX2_X1 U10763 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10171), .Z(n8283) );
  XNOR2_X1 U10764 ( .A(n8283), .B(SI_25_), .ZN(n8286) );
  XNOR2_X1 U10765 ( .A(n8287), .B(n8286), .ZN(n12150) );
  NAND2_X1 U10766 ( .A1(n12150), .A2(n10061), .ZN(n8275) );
  INV_X1 U10767 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12156) );
  XNOR2_X1 U10768 ( .A(n8292), .B(P1_REG3_REG_25__SCAN_IN), .ZN(n14808) );
  NAND2_X1 U10769 ( .A1(n14808), .A2(n8063), .ZN(n8281) );
  INV_X1 U10770 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8278) );
  NAND2_X1 U10771 ( .A1(n9866), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U10772 ( .A1(n10029), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8276) );
  OAI211_X1 U10773 ( .C1(n8278), .C2(n10032), .A(n8277), .B(n8276), .ZN(n8279)
         );
  INV_X1 U10774 ( .A(n8279), .ZN(n8280) );
  NAND2_X2 U10775 ( .A1(n8281), .A2(n8280), .ZN(n14569) );
  XNOR2_X1 U10776 ( .A(n15050), .B(n14569), .ZN(n14802) );
  INV_X1 U10777 ( .A(n14802), .ZN(n14812) );
  NAND2_X1 U10778 ( .A1(n15050), .A2(n14569), .ZN(n8282) );
  INV_X1 U10779 ( .A(n8283), .ZN(n8284) );
  INV_X1 U10780 ( .A(SI_25_), .ZN(n12259) );
  NAND2_X1 U10781 ( .A1(n8284), .A2(n12259), .ZN(n8285) );
  INV_X1 U10782 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12349) );
  INV_X1 U10783 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12352) );
  MUX2_X1 U10784 ( .A(n12349), .B(n12352), .S(n10171), .Z(n8300) );
  XNOR2_X1 U10785 ( .A(n8300), .B(SI_26_), .ZN(n8288) );
  NAND2_X1 U10786 ( .A1(n12348), .A2(n10061), .ZN(n8290) );
  INV_X1 U10787 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14456) );
  INV_X1 U10788 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14544) );
  OAI21_X1 U10789 ( .B1(n8292), .B2(n14456), .A(n14544), .ZN(n8293) );
  NAND2_X1 U10790 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n8291) );
  NAND2_X1 U10791 ( .A1(n14794), .A2(n8063), .ZN(n8298) );
  INV_X1 U10792 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11898) );
  NAND2_X1 U10793 ( .A1(n7835), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U10794 ( .A1(n9866), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8294) );
  OAI211_X1 U10795 ( .C1(n7836), .C2(n11898), .A(n8295), .B(n8294), .ZN(n8296)
         );
  INV_X1 U10796 ( .A(n8296), .ZN(n8297) );
  AND2_X2 U10797 ( .A1(n8298), .A2(n8297), .ZN(n14455) );
  XNOR2_X1 U10798 ( .A(n9888), .B(n14568), .ZN(n10087) );
  OR2_X1 U10799 ( .A1(n15048), .A2(n14455), .ZN(n8299) );
  INV_X1 U10800 ( .A(n8356), .ZN(n8314) );
  INV_X1 U10801 ( .A(SI_26_), .ZN(n13718) );
  INV_X1 U10802 ( .A(n8300), .ZN(n8301) );
  MUX2_X1 U10803 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10171), .Z(n9843) );
  NAND2_X1 U10804 ( .A1(n15162), .A2(n10061), .ZN(n8304) );
  INV_X1 U10805 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15166) );
  INV_X1 U10806 ( .A(n8306), .ZN(n8305) );
  INV_X1 U10807 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U10808 ( .A1(n8306), .A2(n14375), .ZN(n8307) );
  NAND2_X1 U10809 ( .A1(n8361), .A2(n8307), .ZN(n14778) );
  INV_X1 U10810 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n14777) );
  NAND2_X1 U10811 ( .A1(n10029), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U10812 ( .A1(n9866), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8308) );
  OAI211_X1 U10813 ( .C1(n14777), .C2(n10032), .A(n8309), .B(n8308), .ZN(n8310) );
  INV_X1 U10814 ( .A(n8310), .ZN(n8311) );
  INV_X1 U10815 ( .A(n6430), .ZN(n10903) );
  NOR2_X1 U10816 ( .A1(n14583), .A2(n10903), .ZN(n8322) );
  NAND2_X1 U10817 ( .A1(n10509), .A2(n10399), .ZN(n9890) );
  INV_X1 U10818 ( .A(n9890), .ZN(n8315) );
  NAND2_X1 U10819 ( .A1(n9892), .A2(n8316), .ZN(n10549) );
  NAND2_X1 U10820 ( .A1(n10549), .A2(n10548), .ZN(n8318) );
  OR2_X1 U10821 ( .A1(n14585), .A2(n12943), .ZN(n8317) );
  NAND2_X1 U10822 ( .A1(n8318), .A2(n8317), .ZN(n10708) );
  NAND2_X1 U10823 ( .A1(n10810), .A2(n6434), .ZN(n8319) );
  NAND2_X1 U10824 ( .A1(n8320), .A2(n8319), .ZN(n10897) );
  NAND2_X1 U10825 ( .A1(n14583), .A2(n10903), .ZN(n8321) );
  OAI21_X1 U10826 ( .B1(n8322), .B2(n10897), .A(n8321), .ZN(n8323) );
  XNOR2_X1 U10827 ( .A(n11429), .B(n14581), .ZN(n11279) );
  NAND2_X1 U10828 ( .A1(n11220), .A2(n11429), .ZN(n8324) );
  OR2_X1 U10829 ( .A1(n11667), .A2(n11596), .ZN(n8325) );
  NAND2_X1 U10830 ( .A1(n11596), .A2(n11667), .ZN(n8326) );
  OR2_X1 U10831 ( .A1(n12160), .A2(n14521), .ZN(n12069) );
  INV_X1 U10832 ( .A(n14577), .ZN(n12167) );
  AND2_X1 U10833 ( .A1(n12044), .A2(n12167), .ZN(n12065) );
  AOI22_X1 U10834 ( .A1(n12069), .A2(n12065), .B1(n14521), .B2(n12160), .ZN(
        n8328) );
  INV_X1 U10835 ( .A(n14575), .ZN(n14444) );
  NAND2_X1 U10836 ( .A1(n15117), .A2(n14444), .ZN(n8327) );
  AND2_X1 U10837 ( .A1(n8328), .A2(n8327), .ZN(n8329) );
  OR2_X1 U10838 ( .A1(n15117), .A2(n14444), .ZN(n8330) );
  INV_X1 U10839 ( .A(n10080), .ZN(n11836) );
  OR2_X1 U10840 ( .A1(n12205), .A2(n8331), .ZN(n8332) );
  NAND2_X1 U10841 ( .A1(n8333), .A2(n8332), .ZN(n11800) );
  NAND2_X1 U10842 ( .A1(n12307), .A2(n15011), .ZN(n8334) );
  OR2_X1 U10843 ( .A1(n15112), .A2(n14992), .ZN(n9978) );
  NAND2_X1 U10844 ( .A1(n15112), .A2(n14992), .ZN(n9955) );
  INV_X1 U10845 ( .A(n9977), .ZN(n8336) );
  OR2_X1 U10846 ( .A1(n15105), .A2(n6981), .ZN(n8338) );
  XNOR2_X1 U10847 ( .A(n15099), .B(n14572), .ZN(n14948) );
  NAND2_X1 U10848 ( .A1(n14949), .A2(n14948), .ZN(n14947) );
  NAND2_X1 U10849 ( .A1(n14955), .A2(n14572), .ZN(n8339) );
  NAND2_X1 U10850 ( .A1(n15144), .A2(n14950), .ZN(n9988) );
  NAND2_X1 U10851 ( .A1(n14940), .A2(n14407), .ZN(n9986) );
  NAND2_X1 U10852 ( .A1(n9988), .A2(n9986), .ZN(n14929) );
  NAND2_X1 U10853 ( .A1(n15088), .A2(n14932), .ZN(n9991) );
  XNOR2_X1 U10854 ( .A(n14888), .B(n14901), .ZN(n14856) );
  INV_X1 U10855 ( .A(n14873), .ZN(n8342) );
  NAND2_X1 U10856 ( .A1(n14856), .A2(n8342), .ZN(n8343) );
  NAND2_X1 U10857 ( .A1(n15135), .A2(n14901), .ZN(n14857) );
  NAND2_X1 U10858 ( .A1(n8343), .A2(n14857), .ZN(n8344) );
  NOR2_X1 U10859 ( .A1(n14869), .A2(n8344), .ZN(n8345) );
  INV_X1 U10860 ( .A(n14879), .ZN(n14430) );
  NAND2_X1 U10861 ( .A1(n15068), .A2(n14430), .ZN(n8346) );
  NAND2_X1 U10862 ( .A1(n14838), .A2(n14849), .ZN(n14800) );
  INV_X1 U10863 ( .A(n14569), .ZN(n14542) );
  INV_X1 U10864 ( .A(n14571), .ZN(n14508) );
  NAND2_X1 U10865 ( .A1(n15061), .A2(n14508), .ZN(n14799) );
  NAND2_X1 U10866 ( .A1(n8347), .A2(n14799), .ZN(n8348) );
  NAND2_X1 U10867 ( .A1(n14800), .A2(n8349), .ZN(n8354) );
  INV_X1 U10868 ( .A(n8350), .ZN(n14801) );
  OAI21_X1 U10869 ( .B1(n14801), .B2(n14569), .A(n14810), .ZN(n8352) );
  INV_X1 U10870 ( .A(n10092), .ZN(n11408) );
  OR2_X1 U10871 ( .A1(n15297), .A2(n11408), .ZN(n9886) );
  NAND2_X1 U10872 ( .A1(n8371), .A2(n15296), .ZN(n9885) );
  INV_X2 U10873 ( .A(n14988), .ZN(n14874) );
  NAND2_X1 U10874 ( .A1(n9839), .A2(n14874), .ZN(n8358) );
  AOI22_X1 U10875 ( .A1(n15078), .A2(n8356), .B1(n8355), .B2(n14874), .ZN(
        n8357) );
  INV_X1 U10876 ( .A(n8361), .ZN(n8359) );
  NAND2_X1 U10877 ( .A1(n8359), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9865) );
  INV_X1 U10878 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U10879 ( .A1(n8361), .A2(n8360), .ZN(n8362) );
  NAND2_X1 U10880 ( .A1(n14766), .A2(n8063), .ZN(n8367) );
  INV_X1 U10881 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14764) );
  NAND2_X1 U10882 ( .A1(n10029), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U10883 ( .A1(n9866), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8363) );
  OAI211_X1 U10884 ( .C1(n14764), .C2(n10032), .A(n8364), .B(n8363), .ZN(n8365) );
  INV_X1 U10885 ( .A(n8365), .ZN(n8366) );
  NAND2_X1 U10886 ( .A1(n8371), .A2(n10092), .ZN(n10262) );
  OAI22_X1 U10887 ( .A1(n15033), .A2(n14993), .B1(n14455), .B2(n15032), .ZN(
        n8368) );
  INV_X1 U10888 ( .A(n8368), .ZN(n8369) );
  OAI211_X1 U10889 ( .C1(n15314), .C2(n9878), .A(n8370), .B(n8369), .ZN(n14776) );
  NOR2_X2 U10890 ( .A1(n10901), .A2(n6430), .ZN(n11105) );
  NAND2_X1 U10891 ( .A1(n11105), .A2(n11120), .ZN(n11288) );
  OR2_X2 U10892 ( .A1(n11288), .A2(n11429), .ZN(n11465) );
  INV_X1 U10893 ( .A(n11723), .ZN(n15280) );
  INV_X1 U10894 ( .A(n12044), .ZN(n11747) );
  NAND2_X1 U10895 ( .A1(n14953), .A2(n15144), .ZN(n14937) );
  NOR2_X2 U10896 ( .A1(n14937), .A2(n15088), .ZN(n14918) );
  NOR2_X2 U10897 ( .A1(n14844), .A2(n14833), .ZN(n14828) );
  OAI21_X1 U10898 ( .B1(n14365), .B2(n14793), .A(n6432), .ZN(n8372) );
  INV_X1 U10899 ( .A(n14783), .ZN(n8373) );
  NOR2_X1 U10900 ( .A1(n14776), .A2(n8373), .ZN(n8405) );
  INV_X1 U10901 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8400) );
  OAI21_X1 U10902 ( .B1(n8377), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10903 ( .A1(n12154), .A2(P1_B_REG_SCAN_IN), .ZN(n8379) );
  NAND2_X1 U10904 ( .A1(n8377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8378) );
  MUX2_X1 U10905 ( .A(n8379), .B(P1_B_REG_SCAN_IN), .S(n11796), .Z(n8382) );
  NAND2_X1 U10906 ( .A1(n8380), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8381) );
  INV_X1 U10907 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U10908 ( .A1(n10251), .A2(n10255), .ZN(n8383) );
  INV_X1 U10909 ( .A(n8397), .ZN(n12350) );
  NAND2_X1 U10910 ( .A1(n12154), .A2(n12350), .ZN(n10253) );
  NAND2_X1 U10911 ( .A1(n8383), .A2(n10253), .ZN(n9860) );
  NOR4_X1 U10912 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n8392) );
  NOR4_X1 U10913 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n8391) );
  OR4_X1 U10914 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n8389) );
  NOR4_X1 U10915 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n8387) );
  NOR4_X1 U10916 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n8386) );
  NOR4_X1 U10917 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8385) );
  NOR4_X1 U10918 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8384) );
  NAND4_X1 U10919 ( .A1(n8387), .A2(n8386), .A3(n8385), .A4(n8384), .ZN(n8388)
         );
  NOR4_X1 U10920 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n8389), .A4(n8388), .ZN(n8390) );
  NAND3_X1 U10921 ( .A1(n8392), .A2(n8391), .A3(n8390), .ZN(n8393) );
  NAND2_X1 U10922 ( .A1(n10251), .A2(n8393), .ZN(n10375) );
  NAND2_X1 U10923 ( .A1(n6432), .A2(n15296), .ZN(n10394) );
  INV_X1 U10924 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U10925 ( .A1(n10251), .A2(n10259), .ZN(n8394) );
  OR2_X1 U10926 ( .A1(n8397), .A2(n11796), .ZN(n10256) );
  NAND2_X1 U10927 ( .A1(n8394), .A2(n10256), .ZN(n10374) );
  OAI21_X1 U10928 ( .B1(n8395), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8396) );
  XNOR2_X1 U10929 ( .A(n8396), .B(P1_IR_REG_23__SCAN_IN), .ZN(n10261) );
  AND2_X1 U10930 ( .A1(n10257), .A2(n10383), .ZN(n10260) );
  NAND2_X1 U10931 ( .A1(n15297), .A2(n8398), .ZN(n8401) );
  NAND2_X1 U10932 ( .A1(n8401), .A2(n10390), .ZN(n10111) );
  NAND2_X1 U10933 ( .A1(n10260), .A2(n10111), .ZN(n10378) );
  NOR2_X1 U10934 ( .A1(n10374), .A2(n10378), .ZN(n8399) );
  INV_X2 U10935 ( .A(n15322), .ZN(n15320) );
  NAND2_X1 U10936 ( .A1(n15322), .A2(n15311), .ZN(n15096) );
  INV_X1 U10937 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8404) );
  INV_X1 U10938 ( .A(n10378), .ZN(n9861) );
  INV_X1 U10939 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8687) );
  INV_X1 U10940 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8739) );
  INV_X1 U10941 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8760) );
  INV_X1 U10942 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8771) );
  INV_X1 U10943 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13816) );
  NAND2_X1 U10944 ( .A1(n8774), .A2(n13816), .ZN(n8410) );
  NAND2_X1 U10945 ( .A1(n8785), .A2(n8410), .ZN(n13941) );
  NOR2_X1 U10946 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n8412) );
  NOR2_X1 U10947 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8411) );
  NOR2_X1 U10948 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n8416) );
  OR2_X4 U10949 ( .A1(n12355), .A2(n8420), .ZN(n8690) );
  INV_X1 U10950 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U10951 ( .A1(n12816), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8422) );
  NAND2_X1 U10952 ( .A1(n8483), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8421) );
  OAI211_X1 U10953 ( .C1(n8423), .C2(n12820), .A(n8422), .B(n8421), .ZN(n8424)
         );
  INV_X1 U10954 ( .A(n8424), .ZN(n8425) );
  NAND2_X1 U10955 ( .A1(n8809), .A2(n8428), .ZN(n8811) );
  INV_X1 U10956 ( .A(n8429), .ZN(n8430) );
  OAI21_X2 U10957 ( .B1(n8811), .B2(n8430), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8432) );
  NAND2_X1 U10958 ( .A1(n8433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8435) );
  INV_X2 U10959 ( .A(n8757), .ZN(n8496) );
  NAND2_X1 U10960 ( .A1(n12348), .A2(n8496), .ZN(n8437) );
  NAND2_X1 U10961 ( .A1(n8447), .A2(n10193), .ZN(n8471) );
  OR2_X1 U10962 ( .A1(n8471), .A2(n12352), .ZN(n8436) );
  INV_X1 U10963 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10636) );
  INV_X1 U10964 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8439) );
  INV_X1 U10965 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11067) );
  NAND2_X1 U10966 ( .A1(n8440), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10967 ( .A1(n10171), .A2(SI_0_), .ZN(n8444) );
  NAND2_X1 U10968 ( .A1(n8444), .A2(n8938), .ZN(n8446) );
  AND2_X1 U10969 ( .A1(n8446), .A2(n8445), .ZN(n14259) );
  INV_X1 U10970 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8448) );
  INV_X1 U10971 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8449) );
  OR2_X1 U10972 ( .A1(n8485), .A2(n8449), .ZN(n8454) );
  INV_X1 U10973 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11170) );
  INV_X1 U10974 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10423) );
  OR2_X1 U10975 ( .A1(n8451), .A2(n8450), .ZN(n8452) );
  NAND2_X1 U10976 ( .A1(n11176), .A2(n13866), .ZN(n8479) );
  INV_X1 U10977 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10978 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8456) );
  OR2_X1 U10979 ( .A1(n8757), .A2(n10195), .ZN(n8476) );
  OR2_X1 U10980 ( .A1(n8471), .A2(n10172), .ZN(n8477) );
  NAND2_X1 U10981 ( .A1(n8479), .A2(n15466), .ZN(n8465) );
  INV_X1 U10982 ( .A(n11176), .ZN(n8459) );
  NAND2_X1 U10983 ( .A1(n8459), .A2(n8458), .ZN(n8478) );
  INV_X1 U10984 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11973) );
  OR2_X1 U10985 ( .A1(n8485), .A2(n11973), .ZN(n8463) );
  INV_X1 U10986 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8460) );
  INV_X1 U10987 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11394) );
  OR2_X1 U10988 ( .A1(n8690), .A2(n11394), .ZN(n8461) );
  INV_X1 U10989 ( .A(n10278), .ZN(n8466) );
  NAND2_X1 U10990 ( .A1(n8496), .A2(n8466), .ZN(n8474) );
  INV_X1 U10991 ( .A(n8467), .ZN(n8468) );
  NAND2_X1 U10992 ( .A1(n8468), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8469) );
  OR2_X1 U10993 ( .A1(n8497), .A2(n10482), .ZN(n8473) );
  OR2_X1 U10994 ( .A1(n8471), .A2(n10279), .ZN(n8472) );
  NAND3_X1 U10995 ( .A1(n8477), .A2(n8476), .A3(n8475), .ZN(n12666) );
  NAND2_X1 U10996 ( .A1(n8478), .A2(n12666), .ZN(n8480) );
  INV_X1 U10997 ( .A(n13865), .ZN(n8829) );
  NAND3_X1 U10998 ( .A1(n8480), .A2(n8829), .A3(n8479), .ZN(n8481) );
  NAND2_X1 U10999 ( .A1(n8482), .A2(n8481), .ZN(n11190) );
  NAND2_X1 U11000 ( .A1(n8483), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8489) );
  INV_X1 U11001 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8484) );
  OR2_X1 U11002 ( .A1(n8485), .A2(n8484), .ZN(n8488) );
  INV_X1 U11003 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10484) );
  OR2_X1 U11004 ( .A1(n8690), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8486) );
  NOR2_X1 U11005 ( .A1(n10276), .A2(n8757), .ZN(n8493) );
  NAND2_X1 U11006 ( .A1(n8470), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8491) );
  INV_X1 U11007 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8490) );
  OAI22_X1 U11008 ( .A1(n8471), .A2(n10277), .B1(n8497), .B2(n15348), .ZN(
        n8492) );
  OR2_X2 U11009 ( .A1(n8493), .A2(n8492), .ZN(n15471) );
  XNOR2_X1 U11010 ( .A(n11316), .B(n15471), .ZN(n8832) );
  NAND2_X1 U11011 ( .A1(n11190), .A2(n8832), .ZN(n8495) );
  INV_X1 U11012 ( .A(n15471), .ZN(n11197) );
  NAND2_X1 U11013 ( .A1(n11197), .A2(n11316), .ZN(n8494) );
  NAND2_X1 U11014 ( .A1(n8495), .A2(n8494), .ZN(n15439) );
  NAND2_X1 U11015 ( .A1(n10197), .A2(n8496), .ZN(n8504) );
  INV_X2 U11016 ( .A(n8497), .ZN(n10412) );
  INV_X1 U11017 ( .A(n8498), .ZN(n8499) );
  NAND2_X1 U11018 ( .A1(n8499), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8500) );
  MUX2_X1 U11019 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8500), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8502) );
  NAND2_X1 U11020 ( .A1(n8502), .A2(n8501), .ZN(n15360) );
  INV_X1 U11021 ( .A(n15360), .ZN(n10499) );
  NAND2_X1 U11022 ( .A1(n12816), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8508) );
  INV_X1 U11023 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10491) );
  OR2_X1 U11024 ( .A1(n8516), .A2(n10491), .ZN(n8507) );
  OAI21_X1 U11025 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8514), .ZN(n15433) );
  OR2_X1 U11026 ( .A1(n8690), .A2(n15433), .ZN(n8506) );
  INV_X1 U11027 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10485) );
  XNOR2_X1 U11028 ( .A(n12683), .B(n11191), .ZN(n15440) );
  NAND2_X1 U11029 ( .A1(n10238), .A2(n8496), .ZN(n8511) );
  NAND2_X1 U11030 ( .A1(n8501), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8509) );
  XNOR2_X1 U11031 ( .A(n8509), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U11032 ( .A1(n8702), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10412), 
        .B2(n10589), .ZN(n8510) );
  NAND2_X1 U11033 ( .A1(n12816), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8520) );
  INV_X1 U11034 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8512) );
  INV_X1 U11035 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U11036 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  NAND2_X1 U11037 ( .A1(n8537), .A2(n8515), .ZN(n12926) );
  OR2_X1 U11038 ( .A1(n8690), .A2(n12926), .ZN(n8518) );
  INV_X1 U11039 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10500) );
  OR2_X1 U11040 ( .A1(n8516), .A2(n10500), .ZN(n8517) );
  NAND4_X1 U11041 ( .A1(n8520), .A2(n8519), .A3(n8518), .A4(n8517), .ZN(n13862) );
  INV_X1 U11042 ( .A(n11191), .ZN(n13863) );
  OR2_X1 U11043 ( .A1(n13863), .A2(n12683), .ZN(n11054) );
  AND2_X1 U11044 ( .A1(n8521), .A2(n11054), .ZN(n8522) );
  NAND2_X1 U11045 ( .A1(n10246), .A2(n8496), .ZN(n8527) );
  INV_X1 U11046 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U11047 ( .A1(n8545), .A2(n8524), .ZN(n8555) );
  NAND2_X1 U11048 ( .A1(n8555), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8525) );
  XNOR2_X1 U11049 ( .A(n8525), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U11050 ( .A1(n8702), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10412), 
        .B2(n10680), .ZN(n8526) );
  NAND2_X1 U11051 ( .A1(n12816), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8534) );
  INV_X1 U11052 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10679) );
  OR2_X1 U11053 ( .A1(n8516), .A2(n10679), .ZN(n8533) );
  NAND2_X1 U11054 ( .A1(n8539), .A2(n8528), .ZN(n8529) );
  NAND2_X1 U11055 ( .A1(n8562), .A2(n8529), .ZN(n11433) );
  OR2_X1 U11056 ( .A1(n8690), .A2(n11433), .ZN(n8532) );
  INV_X1 U11057 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8530) );
  OR2_X1 U11058 ( .A1(n12820), .A2(n8530), .ZN(n8531) );
  NAND4_X1 U11059 ( .A1(n8534), .A2(n8533), .A3(n8532), .A4(n8531), .ZN(n13860) );
  NAND2_X1 U11060 ( .A1(n8483), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8544) );
  INV_X1 U11061 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8535) );
  OR2_X1 U11062 ( .A1(n8485), .A2(n8535), .ZN(n8543) );
  INV_X1 U11063 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U11064 ( .A1(n8537), .A2(n8536), .ZN(n8538) );
  NAND2_X1 U11065 ( .A1(n8539), .A2(n8538), .ZN(n11552) );
  OR2_X1 U11066 ( .A1(n8690), .A2(n11552), .ZN(n8542) );
  INV_X1 U11067 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8540) );
  OR2_X1 U11068 ( .A1(n12820), .A2(n8540), .ZN(n8541) );
  NAND4_X1 U11069 ( .A1(n8544), .A2(n8543), .A3(n8542), .A4(n8541), .ZN(n13861) );
  NAND2_X1 U11070 ( .A1(n10243), .A2(n8496), .ZN(n8549) );
  INV_X1 U11071 ( .A(n8545), .ZN(n8546) );
  NAND2_X1 U11072 ( .A1(n8546), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8547) );
  XNOR2_X1 U11073 ( .A(n8547), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U11074 ( .A1(n8702), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10412), 
        .B2(n10676), .ZN(n8548) );
  AOI22_X1 U11075 ( .A1(n12700), .A2(n13860), .B1(n13861), .B2(n12692), .ZN(
        n8550) );
  NAND2_X1 U11076 ( .A1(n11237), .A2(n8550), .ZN(n8554) );
  INV_X1 U11077 ( .A(n12700), .ZN(n11436) );
  NAND2_X1 U11078 ( .A1(n11341), .A2(n13860), .ZN(n8552) );
  NOR2_X1 U11079 ( .A1(n13861), .A2(n13860), .ZN(n8551) );
  AOI22_X1 U11080 ( .A1(n11436), .A2(n8552), .B1(n15491), .B2(n8551), .ZN(
        n8553) );
  NAND2_X1 U11081 ( .A1(n8554), .A2(n8553), .ZN(n11561) );
  NAND2_X1 U11082 ( .A1(n10265), .A2(n8496), .ZN(n8560) );
  NAND2_X1 U11083 ( .A1(n8557), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8556) );
  MUX2_X1 U11084 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8556), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8558) );
  NAND2_X1 U11085 ( .A1(n8558), .A2(n8579), .ZN(n10929) );
  INV_X1 U11086 ( .A(n10929), .ZN(n10683) );
  AOI22_X1 U11087 ( .A1(n10412), .A2(n10683), .B1(n8702), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U11088 ( .A1(n12816), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8567) );
  INV_X1 U11089 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10675) );
  OR2_X1 U11090 ( .A1(n12820), .A2(n10675), .ZN(n8566) );
  NAND2_X1 U11091 ( .A1(n8562), .A2(n8561), .ZN(n8563) );
  NAND2_X1 U11092 ( .A1(n8573), .A2(n8563), .ZN(n11586) );
  OR2_X1 U11093 ( .A1(n8690), .A2(n11586), .ZN(n8565) );
  INV_X1 U11094 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10682) );
  OR2_X1 U11095 ( .A1(n8516), .A2(n10682), .ZN(n8564) );
  NAND4_X1 U11096 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n13859) );
  XNOR2_X1 U11097 ( .A(n14217), .B(n13859), .ZN(n12878) );
  NAND2_X1 U11098 ( .A1(n14217), .A2(n13859), .ZN(n8568) );
  NAND2_X1 U11099 ( .A1(n10241), .A2(n8496), .ZN(n8571) );
  NAND2_X1 U11100 ( .A1(n8579), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8569) );
  XNOR2_X1 U11101 ( .A(n8569), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11140) );
  AOI22_X1 U11102 ( .A1(n10412), .A2(n11140), .B1(n8702), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U11103 ( .A1(n12816), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8578) );
  INV_X1 U11104 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8572) );
  OR2_X1 U11105 ( .A1(n12820), .A2(n8572), .ZN(n8577) );
  NAND2_X1 U11106 ( .A1(n8573), .A2(n11994), .ZN(n8574) );
  NAND2_X1 U11107 ( .A1(n8582), .A2(n8574), .ZN(n12588) );
  OR2_X1 U11108 ( .A1(n8690), .A2(n12588), .ZN(n8576) );
  INV_X1 U11109 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11133) );
  OR2_X1 U11110 ( .A1(n8516), .A2(n11133), .ZN(n8575) );
  XNOR2_X1 U11111 ( .A(n12706), .B(n11761), .ZN(n12880) );
  INV_X1 U11112 ( .A(n11761), .ZN(n13857) );
  NAND2_X1 U11113 ( .A1(n12706), .A2(n13857), .ZN(n11754) );
  NAND2_X1 U11114 ( .A1(n10272), .A2(n8496), .ZN(n8581) );
  OAI21_X1 U11115 ( .B1(n8579), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8593) );
  XNOR2_X1 U11116 ( .A(n8593), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U11117 ( .A1(n11268), .A2(n10412), .B1(n8702), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U11118 ( .A1(n8483), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8588) );
  INV_X1 U11119 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11912) );
  OR2_X1 U11120 ( .A1(n8485), .A2(n11912), .ZN(n8587) );
  NAND2_X1 U11121 ( .A1(n8582), .A2(n7192), .ZN(n8583) );
  NAND2_X1 U11122 ( .A1(n8598), .A2(n8583), .ZN(n12188) );
  OR2_X1 U11123 ( .A1(n8690), .A2(n12188), .ZN(n8586) );
  INV_X1 U11124 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8584) );
  OR2_X1 U11125 ( .A1(n12820), .A2(n8584), .ZN(n8585) );
  INV_X1 U11126 ( .A(n12262), .ZN(n13856) );
  NAND2_X1 U11127 ( .A1(n12711), .A2(n13856), .ZN(n8589) );
  AND2_X1 U11128 ( .A1(n11754), .A2(n8589), .ZN(n8591) );
  INV_X1 U11129 ( .A(n8589), .ZN(n8590) );
  NAND2_X1 U11130 ( .A1(n10313), .A2(n8496), .ZN(n8597) );
  INV_X1 U11131 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U11132 ( .A1(n8593), .A2(n8592), .ZN(n8594) );
  NAND2_X1 U11133 ( .A1(n8594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8595) );
  XNOR2_X1 U11134 ( .A(n8595), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U11135 ( .A1(n11359), .A2(n10412), .B1(n8702), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8596) );
  NAND2_X2 U11136 ( .A1(n8597), .A2(n8596), .ZN(n14212) );
  NAND2_X1 U11137 ( .A1(n12816), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8603) );
  INV_X1 U11138 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11353) );
  OR2_X1 U11139 ( .A1(n12820), .A2(n11353), .ZN(n8602) );
  NAND2_X1 U11140 ( .A1(n8598), .A2(n11270), .ZN(n8599) );
  NAND2_X1 U11141 ( .A1(n8610), .A2(n8599), .ZN(n12269) );
  OR2_X1 U11142 ( .A1(n8690), .A2(n12269), .ZN(n8601) );
  INV_X1 U11143 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11874) );
  OR2_X1 U11144 ( .A1(n8516), .A2(n11874), .ZN(n8600) );
  NAND4_X1 U11145 ( .A1(n8603), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n13855) );
  AND2_X1 U11146 ( .A1(n14212), .A2(n13855), .ZN(n8604) );
  NAND2_X1 U11147 ( .A1(n10405), .A2(n8496), .ZN(n8609) );
  INV_X1 U11148 ( .A(n8617), .ZN(n8606) );
  NAND2_X1 U11149 ( .A1(n8606), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U11150 ( .A(n8607), .B(P2_IR_REG_12__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U11151 ( .A1(n8702), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10412), 
        .B2(n12322), .ZN(n8608) );
  NAND2_X1 U11152 ( .A1(n8610), .A2(n7193), .ZN(n8611) );
  NAND2_X1 U11153 ( .A1(n8621), .A2(n8611), .ZN(n12627) );
  OR2_X1 U11154 ( .A1(n8690), .A2(n12627), .ZN(n8615) );
  INV_X1 U11155 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n12144) );
  OR2_X1 U11156 ( .A1(n8516), .A2(n12144), .ZN(n8614) );
  INV_X1 U11157 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n12346) );
  OR2_X1 U11158 ( .A1(n8485), .A2(n12346), .ZN(n8613) );
  INV_X1 U11159 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n12343) );
  OR2_X1 U11160 ( .A1(n12820), .A2(n12343), .ZN(n8612) );
  NAND4_X1 U11161 ( .A1(n8615), .A2(n8614), .A3(n8613), .A4(n8612), .ZN(n13854) );
  NAND2_X1 U11162 ( .A1(n12733), .A2(n13854), .ZN(n8616) );
  NAND2_X1 U11163 ( .A1(n10463), .A2(n8496), .ZN(n8620) );
  NAND2_X1 U11164 ( .A1(n8617), .A2(n11996), .ZN(n8629) );
  NAND2_X1 U11165 ( .A1(n8629), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8618) );
  XNOR2_X1 U11166 ( .A(n8618), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15397) );
  AOI22_X1 U11167 ( .A1(n8702), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10412), 
        .B2(n15397), .ZN(n8619) );
  NAND2_X1 U11168 ( .A1(n8621), .A2(n13777), .ZN(n8622) );
  NAND2_X1 U11169 ( .A1(n8635), .A2(n8622), .ZN(n13780) );
  NAND2_X1 U11170 ( .A1(n12816), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U11171 ( .A1(n8440), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8623) );
  AND2_X1 U11172 ( .A1(n8624), .A2(n8623), .ZN(n8626) );
  NAND2_X1 U11173 ( .A1(n8483), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8625) );
  OAI211_X1 U11174 ( .C1(n8690), .C2(n13780), .A(n8626), .B(n8625), .ZN(n13853) );
  AND2_X1 U11175 ( .A1(n14206), .A2(n13853), .ZN(n8628) );
  OR2_X1 U11176 ( .A1(n14206), .A2(n13853), .ZN(n8627) );
  NAND2_X1 U11177 ( .A1(n10765), .A2(n8496), .ZN(n8633) );
  NOR2_X2 U11178 ( .A1(n8629), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8641) );
  INV_X1 U11179 ( .A(n8641), .ZN(n8630) );
  NAND2_X1 U11180 ( .A1(n8630), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8631) );
  XNOR2_X1 U11181 ( .A(n8631), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U11182 ( .A1(n8702), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10412), 
        .B2(n12323), .ZN(n8632) );
  NAND2_X1 U11183 ( .A1(n8635), .A2(n8634), .ZN(n8636) );
  NAND2_X1 U11184 ( .A1(n8646), .A2(n8636), .ZN(n13006) );
  AOI22_X1 U11185 ( .A1(n8483), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12816), 
        .B2(P2_REG0_REG_14__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U11186 ( .A1(n8440), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8637) );
  OAI211_X1 U11187 ( .C1(n13006), .C2(n8690), .A(n8638), .B(n8637), .ZN(n13852) );
  NOR2_X1 U11188 ( .A1(n14201), .A2(n13852), .ZN(n8639) );
  INV_X1 U11189 ( .A(n13852), .ZN(n12727) );
  INV_X1 U11190 ( .A(n14201), .ZN(n12726) );
  NAND2_X1 U11191 ( .A1(n10703), .A2(n8496), .ZN(n8644) );
  NAND2_X1 U11192 ( .A1(n8641), .A2(n8640), .ZN(n8652) );
  NAND2_X1 U11193 ( .A1(n8652), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8642) );
  XNOR2_X1 U11194 ( .A(n8642), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U11195 ( .A1(n10412), .A2(n13875), .B1(n8702), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n8643) );
  INV_X1 U11196 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8650) );
  INV_X1 U11197 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U11198 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  NAND2_X1 U11199 ( .A1(n8661), .A2(n8647), .ZN(n13829) );
  OR2_X1 U11200 ( .A1(n13829), .A2(n8690), .ZN(n8649) );
  AOI22_X1 U11201 ( .A1(n8483), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12816), 
        .B2(P2_REG0_REG_15__SCAN_IN), .ZN(n8648) );
  OAI211_X1 U11202 ( .C1(n12820), .C2(n8650), .A(n8649), .B(n8648), .ZN(n13851) );
  XNOR2_X1 U11203 ( .A(n13831), .B(n13851), .ZN(n12885) );
  OR2_X1 U11204 ( .A1(n13831), .A2(n13851), .ZN(n8651) );
  NAND2_X1 U11205 ( .A1(n10751), .A2(n8496), .ZN(n8659) );
  INV_X1 U11206 ( .A(n8656), .ZN(n8653) );
  NAND2_X1 U11207 ( .A1(n8653), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8654) );
  MUX2_X1 U11208 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8654), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8657) );
  NAND2_X1 U11209 ( .A1(n8656), .A2(n8655), .ZN(n8682) );
  AND2_X1 U11210 ( .A1(n8657), .A2(n8682), .ZN(n13891) );
  AOI22_X1 U11211 ( .A1(n13891), .A2(n10412), .B1(n8702), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U11212 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  AND2_X1 U11213 ( .A1(n8673), .A2(n8662), .ZN(n14084) );
  NAND2_X1 U11214 ( .A1(n14084), .A2(n8787), .ZN(n8667) );
  INV_X1 U11215 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13867) );
  NAND2_X1 U11216 ( .A1(n12816), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U11217 ( .A1(n8440), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8663) );
  OAI211_X1 U11218 ( .C1(n13867), .C2(n8516), .A(n8664), .B(n8663), .ZN(n8665)
         );
  INV_X1 U11219 ( .A(n8665), .ZN(n8666) );
  XNOR2_X1 U11220 ( .A(n14086), .B(n12719), .ZN(n14073) );
  NAND2_X1 U11221 ( .A1(n10953), .A2(n8496), .ZN(n8671) );
  NAND2_X1 U11222 ( .A1(n8682), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8668) );
  XNOR2_X1 U11223 ( .A(n8668), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13906) );
  NOR2_X1 U11224 ( .A1(n12824), .A2(n11977), .ZN(n8669) );
  AOI21_X1 U11225 ( .B1(n13906), .B2(n10412), .A(n8669), .ZN(n8670) );
  NAND2_X2 U11226 ( .A1(n8671), .A2(n8670), .ZN(n14181) );
  INV_X1 U11227 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8672) );
  NAND2_X1 U11228 ( .A1(n8673), .A2(n8672), .ZN(n8674) );
  NAND2_X1 U11229 ( .A1(n8688), .A2(n8674), .ZN(n14059) );
  INV_X1 U11230 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14063) );
  NAND2_X1 U11231 ( .A1(n12816), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U11232 ( .A1(n8440), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8675) );
  OAI211_X1 U11233 ( .C1(n8516), .C2(n14063), .A(n8676), .B(n8675), .ZN(n8677)
         );
  INV_X1 U11234 ( .A(n8677), .ZN(n8678) );
  NAND2_X1 U11235 ( .A1(n8679), .A2(n8678), .ZN(n13849) );
  AND2_X1 U11236 ( .A1(n14181), .A2(n13849), .ZN(n8681) );
  OR2_X1 U11237 ( .A1(n14181), .A2(n13849), .ZN(n8680) );
  OR2_X1 U11238 ( .A1(n11131), .A2(n8757), .ZN(n8686) );
  NOR2_X2 U11239 ( .A1(n8682), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8699) );
  INV_X1 U11240 ( .A(n8699), .ZN(n8683) );
  NAND2_X1 U11241 ( .A1(n8683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8684) );
  XNOR2_X1 U11242 ( .A(n8684), .B(P2_IR_REG_18__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U11243 ( .A1(n15422), .A2(n10412), .B1(n8702), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U11244 ( .A1(n8688), .A2(n8687), .ZN(n8689) );
  NAND2_X1 U11245 ( .A1(n8705), .A2(n8689), .ZN(n14049) );
  OR2_X1 U11246 ( .A1(n14049), .A2(n8690), .ZN(n8696) );
  INV_X1 U11247 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U11248 ( .A1(n8483), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U11249 ( .A1(n12816), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8691) );
  OAI211_X1 U11250 ( .C1(n8693), .C2(n12820), .A(n8692), .B(n8691), .ZN(n8694)
         );
  INV_X1 U11251 ( .A(n8694), .ZN(n8695) );
  XNOR2_X1 U11252 ( .A(n14048), .B(n12645), .ZN(n14045) );
  NAND2_X1 U11253 ( .A1(n14173), .A2(n12645), .ZN(n8697) );
  NAND2_X1 U11254 ( .A1(n11423), .A2(n8496), .ZN(n8704) );
  INV_X1 U11255 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8698) );
  XNOR2_X2 U11256 ( .A(n8701), .B(n8700), .ZN(n9657) );
  AOI22_X1 U11257 ( .A1(n13916), .A2(n10412), .B1(n8702), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U11258 ( .A1(n8705), .A2(n11975), .ZN(n8706) );
  NAND2_X1 U11259 ( .A1(n8714), .A2(n8706), .ZN(n14034) );
  INV_X1 U11260 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14035) );
  NAND2_X1 U11261 ( .A1(n8440), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11262 ( .A1(n12816), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8707) );
  OAI211_X1 U11263 ( .C1(n8516), .C2(n14035), .A(n8708), .B(n8707), .ZN(n8709)
         );
  INV_X1 U11264 ( .A(n8709), .ZN(n8710) );
  NOR2_X1 U11265 ( .A1(n14163), .A2(n13847), .ZN(n8711) );
  INV_X1 U11266 ( .A(n13847), .ZN(n13771) );
  OR2_X1 U11267 ( .A1(n12824), .A2(n11383), .ZN(n8712) );
  NAND2_X1 U11268 ( .A1(n8714), .A2(n7196), .ZN(n8715) );
  AND2_X1 U11269 ( .A1(n8725), .A2(n8715), .ZN(n14025) );
  NAND2_X1 U11270 ( .A1(n14025), .A2(n8787), .ZN(n8721) );
  INV_X1 U11271 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U11272 ( .A1(n8483), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U11273 ( .A1(n12816), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8716) );
  OAI211_X1 U11274 ( .C1(n8718), .C2(n12820), .A(n8717), .B(n8716), .ZN(n8719)
         );
  INV_X1 U11275 ( .A(n8719), .ZN(n8720) );
  NAND2_X1 U11276 ( .A1(n8721), .A2(n8720), .ZN(n13846) );
  AND2_X1 U11277 ( .A1(n14159), .A2(n13846), .ZN(n8722) );
  INV_X1 U11278 ( .A(n13846), .ZN(n13734) );
  OR2_X1 U11279 ( .A1(n11407), .A2(n8757), .ZN(n8724) );
  INV_X1 U11280 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11405) );
  OR2_X1 U11281 ( .A1(n12824), .A2(n11405), .ZN(n8723) );
  NAND2_X1 U11282 ( .A1(n8725), .A2(n7197), .ZN(n8726) );
  NAND2_X1 U11283 ( .A1(n8740), .A2(n8726), .ZN(n14011) );
  INV_X1 U11284 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U11285 ( .A1(n8483), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U11286 ( .A1(n12816), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8727) );
  OAI211_X1 U11287 ( .C1(n8729), .C2(n12820), .A(n8728), .B(n8727), .ZN(n8730)
         );
  INV_X1 U11288 ( .A(n8730), .ZN(n8731) );
  XNOR2_X1 U11289 ( .A(n14151), .B(n13787), .ZN(n14016) );
  NAND2_X1 U11290 ( .A1(n8734), .A2(n8733), .ZN(n8735) );
  NAND2_X1 U11291 ( .A1(n8736), .A2(n8735), .ZN(n11510) );
  OR2_X1 U11292 ( .A1(n12824), .A2(n11511), .ZN(n8737) );
  NAND2_X1 U11293 ( .A1(n8740), .A2(n8739), .ZN(n8741) );
  AND2_X1 U11294 ( .A1(n8749), .A2(n8741), .ZN(n13994) );
  INV_X1 U11295 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11296 ( .A1(n8483), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11297 ( .A1(n12816), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8742) );
  OAI211_X1 U11298 ( .C1(n8744), .C2(n12820), .A(n8743), .B(n8742), .ZN(n8745)
         );
  XNOR2_X1 U11299 ( .A(n14147), .B(n13791), .ZN(n13986) );
  INV_X1 U11300 ( .A(n14147), .ZN(n13997) );
  NAND2_X1 U11301 ( .A1(n11733), .A2(n8496), .ZN(n8747) );
  INV_X1 U11302 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11732) );
  OR2_X1 U11303 ( .A1(n12824), .A2(n11732), .ZN(n8746) );
  INV_X1 U11304 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11305 ( .A1(n8749), .A2(n8748), .ZN(n8750) );
  NAND2_X1 U11306 ( .A1(n8761), .A2(n8750), .ZN(n13721) );
  INV_X1 U11307 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11308 ( .A1(n8483), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U11309 ( .A1(n12816), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8751) );
  OAI211_X1 U11310 ( .C1(n8753), .C2(n12820), .A(n8752), .B(n8751), .ZN(n8754)
         );
  INV_X1 U11311 ( .A(n8754), .ZN(n8755) );
  OR2_X1 U11312 ( .A1(n14138), .A2(n13843), .ZN(n12865) );
  AND2_X1 U11313 ( .A1(n14138), .A2(n13843), .ZN(n12866) );
  OR2_X1 U11314 ( .A1(n11798), .A2(n8757), .ZN(n8759) );
  OR2_X1 U11315 ( .A1(n8471), .A2(n11794), .ZN(n8758) );
  NAND2_X1 U11316 ( .A1(n8761), .A2(n8760), .ZN(n8762) );
  AND2_X1 U11317 ( .A1(n8772), .A2(n8762), .ZN(n13967) );
  NAND2_X1 U11318 ( .A1(n13967), .A2(n8787), .ZN(n8768) );
  INV_X1 U11319 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U11320 ( .A1(n8483), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11321 ( .A1(n12816), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8763) );
  OAI211_X1 U11322 ( .C1(n8765), .C2(n12820), .A(n8764), .B(n8763), .ZN(n8766)
         );
  INV_X1 U11323 ( .A(n8766), .ZN(n8767) );
  INV_X1 U11324 ( .A(n13842), .ZN(n8868) );
  NAND2_X1 U11325 ( .A1(n12150), .A2(n8496), .ZN(n8770) );
  INV_X1 U11326 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12153) );
  OR2_X1 U11327 ( .A1(n12824), .A2(n12153), .ZN(n8769) );
  NAND2_X1 U11328 ( .A1(n8772), .A2(n8771), .ZN(n8773) );
  NAND2_X1 U11329 ( .A1(n13955), .A2(n8787), .ZN(n8780) );
  INV_X1 U11330 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U11331 ( .A1(n12816), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11332 ( .A1(n8483), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8775) );
  OAI211_X1 U11333 ( .C1(n12820), .C2(n8777), .A(n8776), .B(n8775), .ZN(n8778)
         );
  INV_X1 U11334 ( .A(n8778), .ZN(n8779) );
  NOR2_X1 U11335 ( .A1(n14126), .A2(n13813), .ZN(n8781) );
  NAND2_X1 U11336 ( .A1(n15162), .A2(n8496), .ZN(n8783) );
  INV_X1 U11337 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12955) );
  OR2_X1 U11338 ( .A1(n12824), .A2(n12955), .ZN(n8782) );
  INV_X1 U11339 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U11340 ( .A1(n8785), .A2(n8784), .ZN(n8786) );
  NAND2_X1 U11341 ( .A1(n13934), .A2(n8787), .ZN(n8793) );
  INV_X1 U11342 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U11343 ( .A1(n8440), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U11344 ( .A1(n12816), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8788) );
  OAI211_X1 U11345 ( .C1(n8516), .C2(n8790), .A(n8789), .B(n8788), .ZN(n8791)
         );
  INV_X1 U11346 ( .A(n8791), .ZN(n8792) );
  INV_X1 U11347 ( .A(n13839), .ZN(n13815) );
  INV_X1 U11348 ( .A(n14115), .ZN(n13937) );
  NAND2_X1 U11349 ( .A1(n9849), .A2(n9843), .ZN(n8795) );
  MUX2_X1 U11350 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n10171), .Z(n8796) );
  NAND2_X1 U11351 ( .A1(n8796), .A2(SI_28_), .ZN(n9845) );
  NOR2_X1 U11352 ( .A1(n8796), .A2(SI_28_), .ZN(n9844) );
  INV_X1 U11353 ( .A(n9844), .ZN(n8797) );
  NAND2_X1 U11354 ( .A1(n9845), .A2(n8797), .ZN(n8798) );
  NAND2_X1 U11355 ( .A1(n12944), .A2(n8496), .ZN(n8800) );
  INV_X1 U11356 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9804) );
  OR2_X1 U11357 ( .A1(n12824), .A2(n9804), .ZN(n8799) );
  NAND2_X2 U11358 ( .A1(n8800), .A2(n8799), .ZN(n13000) );
  NAND2_X1 U11359 ( .A1(n7186), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12971) );
  INV_X1 U11360 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U11361 ( .A1(n8801), .A2(n12996), .ZN(n8802) );
  INV_X1 U11362 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U11363 ( .A1(n8483), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8804) );
  NAND2_X1 U11364 ( .A1(n12816), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8803) );
  OAI211_X1 U11365 ( .C1(n8805), .C2(n12820), .A(n8804), .B(n8803), .ZN(n8806)
         );
  INV_X1 U11366 ( .A(n8806), .ZN(n8807) );
  NAND2_X1 U11367 ( .A1(n13000), .A2(n12828), .ZN(n8808) );
  XNOR2_X1 U11368 ( .A(n14109), .B(n14104), .ZN(n12626) );
  OAI21_X1 U11369 ( .B1(n8815), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8810) );
  NAND2_X1 U11370 ( .A1(n8819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8814) );
  MUX2_X1 U11371 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8814), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8816) );
  NAND2_X1 U11372 ( .A1(n12899), .A2(n11381), .ZN(n12901) );
  XNOR2_X1 U11373 ( .A(n6437), .B(n12901), .ZN(n8817) );
  NAND3_X1 U11374 ( .A1(n8818), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_19__SCAN_IN), .ZN(n8825) );
  INV_X1 U11375 ( .A(n8819), .ZN(n8821) );
  NOR2_X1 U11376 ( .A1(n6437), .A2(n8823), .ZN(n8824) );
  NAND2_X1 U11377 ( .A1(n8458), .A2(n12665), .ZN(n8828) );
  XNOR2_X1 U11378 ( .A(n13865), .B(n12670), .ZN(n12870) );
  NAND2_X1 U11379 ( .A1(n10697), .A2(n12870), .ZN(n8831) );
  NAND2_X1 U11380 ( .A1(n8829), .A2(n12670), .ZN(n8830) );
  NAND2_X1 U11381 ( .A1(n8831), .A2(n8830), .ZN(n11200) );
  INV_X1 U11382 ( .A(n8832), .ZN(n12873) );
  NAND2_X1 U11383 ( .A1(n11200), .A2(n12873), .ZN(n8834) );
  NAND2_X1 U11384 ( .A1(n11316), .A2(n15471), .ZN(n8833) );
  NAND2_X1 U11385 ( .A1(n8834), .A2(n8833), .ZN(n15430) );
  INV_X1 U11386 ( .A(n15440), .ZN(n15429) );
  NAND2_X1 U11387 ( .A1(n12683), .A2(n11191), .ZN(n8835) );
  OR2_X1 U11388 ( .A1(n12933), .A2(n6875), .ZN(n8837) );
  NAND2_X1 U11389 ( .A1(n12692), .A2(n11387), .ZN(n8838) );
  NAND2_X1 U11390 ( .A1(n11241), .A2(n8838), .ZN(n11346) );
  INV_X1 U11391 ( .A(n13860), .ZN(n11578) );
  OR2_X1 U11392 ( .A1(n12700), .A2(n11578), .ZN(n8839) );
  NAND2_X1 U11393 ( .A1(n12700), .A2(n11578), .ZN(n8840) );
  INV_X1 U11394 ( .A(n13859), .ZN(n11347) );
  AND2_X1 U11395 ( .A1(n14217), .A2(n11347), .ZN(n8842) );
  INV_X1 U11396 ( .A(n12880), .ZN(n11695) );
  INV_X1 U11397 ( .A(n12881), .ZN(n11760) );
  OR2_X1 U11398 ( .A1(n12711), .A2(n12262), .ZN(n8843) );
  NAND2_X1 U11399 ( .A1(n8844), .A2(n8843), .ZN(n11869) );
  INV_X1 U11400 ( .A(n13854), .ZN(n12732) );
  OR2_X1 U11401 ( .A1(n12733), .A2(n12732), .ZN(n12275) );
  OAI21_X1 U11402 ( .B1(n12718), .B2(n14212), .A(n12275), .ZN(n8848) );
  NAND2_X1 U11403 ( .A1(n14212), .A2(n12718), .ZN(n12139) );
  NAND2_X1 U11404 ( .A1(n12139), .A2(n13854), .ZN(n8846) );
  NOR2_X1 U11405 ( .A1(n13854), .A2(n13855), .ZN(n8845) );
  AOI22_X1 U11406 ( .A1(n12733), .A2(n8846), .B1(n8845), .B2(n14212), .ZN(
        n8847) );
  XNOR2_X1 U11407 ( .A(n14206), .B(n13853), .ZN(n12886) );
  INV_X1 U11408 ( .A(n13853), .ZN(n13008) );
  OR2_X1 U11409 ( .A1(n14206), .A2(n13008), .ZN(n8849) );
  NOR2_X1 U11410 ( .A1(n14201), .A2(n12727), .ZN(n8852) );
  NAND2_X1 U11411 ( .A1(n14201), .A2(n12727), .ZN(n8851) );
  INV_X1 U11412 ( .A(n13851), .ZN(n12724) );
  AND2_X1 U11413 ( .A1(n13831), .A2(n12724), .ZN(n8853) );
  OR2_X1 U11414 ( .A1(n13831), .A2(n12724), .ZN(n8854) );
  INV_X1 U11415 ( .A(n14086), .ZN(n14188) );
  INV_X1 U11416 ( .A(n13849), .ZN(n8855) );
  OR2_X1 U11417 ( .A1(n14181), .A2(n8855), .ZN(n12721) );
  NOR2_X1 U11418 ( .A1(n14048), .A2(n12645), .ZN(n8856) );
  NAND2_X1 U11419 ( .A1(n14151), .A2(n13787), .ZN(n8860) );
  NAND2_X1 U11420 ( .A1(n14159), .A2(n13734), .ZN(n12868) );
  NAND2_X1 U11421 ( .A1(n14163), .A2(n13771), .ZN(n8857) );
  NAND2_X1 U11422 ( .A1(n14048), .A2(n12645), .ZN(n14000) );
  AND4_X1 U11423 ( .A1(n8860), .A2(n12868), .A3(n8857), .A4(n14000), .ZN(n8858) );
  INV_X1 U11424 ( .A(n12868), .ZN(n14004) );
  OR2_X1 U11425 ( .A1(n14163), .A2(n13771), .ZN(n14002) );
  NAND2_X1 U11426 ( .A1(n14028), .A2(n13846), .ZN(n12869) );
  NAND2_X1 U11427 ( .A1(n14010), .A2(n13845), .ZN(n8859) );
  OAI211_X1 U11428 ( .C1(n14004), .C2(n14002), .A(n12869), .B(n8859), .ZN(
        n8861) );
  NAND2_X1 U11429 ( .A1(n8861), .A2(n8860), .ZN(n8862) );
  NAND2_X1 U11430 ( .A1(n8863), .A2(n8862), .ZN(n13989) );
  INV_X1 U11431 ( .A(n13986), .ZN(n13988) );
  NAND2_X1 U11432 ( .A1(n13989), .A2(n13988), .ZN(n13987) );
  INV_X1 U11433 ( .A(n13791), .ZN(n13844) );
  NAND2_X1 U11434 ( .A1(n13997), .A2(n13844), .ZN(n8864) );
  INV_X1 U11435 ( .A(n13843), .ZN(n8865) );
  NOR2_X1 U11436 ( .A1(n14138), .A2(n8865), .ZN(n8867) );
  NAND2_X1 U11437 ( .A1(n14138), .A2(n8865), .ZN(n8866) );
  XNOR2_X1 U11438 ( .A(n13958), .B(n13841), .ZN(n13953) );
  NAND2_X1 U11439 ( .A1(n13954), .A2(n13953), .ZN(n8870) );
  NAND2_X1 U11440 ( .A1(n13958), .A2(n13813), .ZN(n8869) );
  OR2_X1 U11441 ( .A1(n14119), .A2(n12830), .ZN(n12864) );
  AND2_X1 U11442 ( .A1(n14119), .A2(n12830), .ZN(n12863) );
  INV_X1 U11443 ( .A(n13925), .ZN(n13928) );
  NOR2_X1 U11444 ( .A1(n13937), .A2(n13839), .ZN(n8872) );
  NAND2_X1 U11445 ( .A1(n13916), .A2(n6437), .ZN(n8871) );
  NAND2_X1 U11446 ( .A1(n12899), .A2(n6993), .ZN(n12913) );
  NOR2_X1 U11447 ( .A1(n12958), .A2(n14186), .ZN(n8883) );
  OAI21_X1 U11448 ( .B1(n13927), .B2(n8872), .A(n14104), .ZN(n8882) );
  OR2_X1 U11449 ( .A1(n12971), .A2(n8690), .ZN(n8878) );
  INV_X1 U11450 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U11451 ( .A1(n8483), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11452 ( .A1(n12816), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8873) );
  OAI211_X1 U11453 ( .C1(n12820), .C2(n8875), .A(n8874), .B(n8873), .ZN(n8876)
         );
  INV_X1 U11454 ( .A(n8876), .ZN(n8877) );
  NAND2_X1 U11455 ( .A1(n8878), .A2(n8877), .ZN(n13837) );
  NAND2_X1 U11456 ( .A1(n13837), .A2(n13802), .ZN(n8881) );
  INV_X1 U11457 ( .A(n10420), .ZN(n8879) );
  NAND2_X1 U11458 ( .A1(n13839), .A2(n13801), .ZN(n8880) );
  NAND2_X1 U11459 ( .A1(n8881), .A2(n8880), .ZN(n12999) );
  AOI21_X1 U11460 ( .B1(n8883), .B2(n8882), .A(n12999), .ZN(n12621) );
  INV_X1 U11461 ( .A(n12683), .ZN(n15482) );
  NAND2_X1 U11462 ( .A1(n15441), .A2(n15482), .ZN(n15444) );
  INV_X1 U11463 ( .A(n14217), .ZN(n11582) );
  NOR2_X4 U11464 ( .A1(n11697), .A2(n12706), .ZN(n11698) );
  INV_X1 U11465 ( .A(n12733), .ZN(n12731) );
  NOR2_X2 U11466 ( .A1(n7731), .A2(n14201), .ZN(n12310) );
  OR2_X2 U11467 ( .A1(n14080), .A2(n14086), .ZN(n14081) );
  NAND2_X1 U11468 ( .A1(n14008), .A2(n14010), .ZN(n14009) );
  OR2_X2 U11469 ( .A1(n14009), .A2(n14147), .ZN(n13992) );
  OR2_X2 U11470 ( .A1(n14115), .A2(n13940), .ZN(n13932) );
  NOR2_X2 U11471 ( .A1(n13932), .A2(n13000), .ZN(n12969) );
  AOI211_X1 U11472 ( .C1(n13000), .C2(n13932), .A(n14166), .B(n12969), .ZN(
        n12624) );
  AOI21_X1 U11473 ( .B1(n15472), .B2(n13000), .A(n12624), .ZN(n8886) );
  NAND2_X1 U11474 ( .A1(n8891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8887) );
  INV_X1 U11475 ( .A(P2_B_REG_SCAN_IN), .ZN(n12949) );
  NAND2_X1 U11476 ( .A1(n8888), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8890) );
  XNOR2_X1 U11477 ( .A(n12949), .B(n11795), .ZN(n8893) );
  OAI22_X1 U11478 ( .A1(n15449), .A2(P2_D_REG_0__SCAN_IN), .B1(n8894), .B2(
        n12351), .ZN(n9790) );
  NAND3_X1 U11479 ( .A1(n12351), .A2(n8894), .A3(n12151), .ZN(n10160) );
  NOR4_X1 U11480 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8902) );
  NOR4_X1 U11481 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8901) );
  NOR4_X1 U11482 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8900) );
  NOR4_X1 U11483 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8899) );
  NAND4_X1 U11484 ( .A1(n8902), .A2(n8901), .A3(n8900), .A4(n8899), .ZN(n8909)
         );
  NOR2_X1 U11485 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .ZN(
        n8906) );
  NOR4_X1 U11486 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8905) );
  NOR4_X1 U11487 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n8904) );
  NOR4_X1 U11488 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8903) );
  NAND4_X1 U11489 ( .A1(n8906), .A2(n8905), .A3(n8904), .A4(n8903), .ZN(n8908)
         );
  INV_X1 U11490 ( .A(n15449), .ZN(n8907) );
  OAI21_X1 U11491 ( .B1(n8909), .B2(n8908), .A(n8907), .ZN(n9780) );
  OR2_X1 U11492 ( .A1(n15449), .A2(P2_D_REG_1__SCAN_IN), .ZN(n8911) );
  OR2_X1 U11493 ( .A1(n12351), .A2(n12151), .ZN(n8910) );
  NAND2_X1 U11494 ( .A1(n8911), .A2(n8910), .ZN(n15458) );
  AND3_X1 U11495 ( .A1(n9792), .A2(n9780), .A3(n15458), .ZN(n8914) );
  NAND2_X1 U11496 ( .A1(n15500), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U11497 ( .A1(n8913), .A2(n8912), .ZN(P2_U3527) );
  AND2_X1 U11498 ( .A1(n8914), .A2(n15459), .ZN(n8915) );
  NAND2_X1 U11499 ( .A1(n8916), .A2(n15496), .ZN(n8919) );
  INV_X1 U11500 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8917) );
  OR2_X1 U11501 ( .A1(n15496), .A2(n8917), .ZN(n8918) );
  NAND2_X1 U11502 ( .A1(n8919), .A2(n8918), .ZN(P2_U3495) );
  INV_X1 U11503 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9468) );
  INV_X1 U11504 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8920) );
  NOR2_X1 U11505 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), 
        .ZN(n8924) );
  NOR2_X1 U11506 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), 
        .ZN(n8923) );
  NOR2_X1 U11507 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8922) );
  INV_X1 U11508 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8926) );
  XNOR2_X2 U11509 ( .A(n8928), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8933) );
  NAND2_X4 U11510 ( .A1(n12617), .A2(n8929), .ZN(n12366) );
  INV_X1 U11511 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10627) );
  INV_X1 U11512 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15554) );
  INV_X1 U11513 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8930) );
  OR2_X1 U11514 ( .A1(n9015), .A2(n8930), .ZN(n8935) );
  XOR2_X1 U11515 ( .A(n8931), .B(P3_IR_REG_29__SCAN_IN), .Z(n8932) );
  NAND2_X2 U11516 ( .A1(n8933), .A2(n8932), .ZN(n12365) );
  INV_X1 U11517 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15558) );
  OR2_X1 U11518 ( .A1(n12376), .A2(n10176), .ZN(n8945) );
  INV_X1 U11519 ( .A(n8963), .ZN(n8952) );
  XNOR2_X1 U11520 ( .A(n8964), .B(n8952), .ZN(n10175) );
  OR2_X1 U11521 ( .A1(n9149), .A2(n10175), .ZN(n8944) );
  INV_X2 U11522 ( .A(n9564), .ZN(n9024) );
  INV_X1 U11523 ( .A(n9530), .ZN(n8941) );
  NAND2_X2 U11524 ( .A1(n8942), .A2(n8941), .ZN(n10634) );
  INV_X1 U11525 ( .A(n10634), .ZN(n9568) );
  NAND2_X1 U11526 ( .A1(n9024), .A2(n9568), .ZN(n8943) );
  INV_X1 U11527 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n9569) );
  OR2_X1 U11528 ( .A1(n12366), .A2(n9569), .ZN(n8949) );
  NAND2_X1 U11529 ( .A1(n9075), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8948) );
  INV_X1 U11530 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10876) );
  OR2_X1 U11531 ( .A1(n9425), .A2(n10876), .ZN(n8947) );
  INV_X1 U11532 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U11533 ( .A1(n8950), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8951) );
  AND2_X1 U11534 ( .A1(n8952), .A2(n8951), .ZN(n10178) );
  OR2_X1 U11535 ( .A1(n9149), .A2(n10178), .ZN(n8954) );
  NAND2_X1 U11536 ( .A1(n9024), .A2(n6864), .ZN(n8953) );
  AND2_X1 U11537 ( .A1(n15545), .A2(n11019), .ZN(n15547) );
  INV_X1 U11538 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15527) );
  OR2_X1 U11539 ( .A1(n9425), .A2(n15527), .ZN(n8959) );
  INV_X1 U11540 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8956) );
  OR2_X1 U11541 ( .A1(n9015), .A2(n8956), .ZN(n8958) );
  INV_X1 U11542 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n9573) );
  OR2_X1 U11543 ( .A1(n12365), .A2(n9573), .ZN(n8957) );
  NOR2_X1 U11544 ( .A1(n9530), .A2(n9165), .ZN(n8961) );
  INV_X1 U11545 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11546 ( .A1(n10172), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8965) );
  XNOR2_X1 U11547 ( .A(n8974), .B(n8973), .ZN(n10181) );
  NAND2_X1 U11548 ( .A1(n15544), .A2(n15524), .ZN(n12402) );
  OR2_X1 U11549 ( .A1(n15544), .A2(n6700), .ZN(n8966) );
  NAND2_X1 U11550 ( .A1(n9093), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8970) );
  OR2_X1 U11551 ( .A1(n9425), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8969) );
  INV_X1 U11552 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n11995) );
  OR2_X1 U11553 ( .A1(n9015), .A2(n11995), .ZN(n8968) );
  INV_X1 U11554 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11162) );
  OR2_X1 U11555 ( .A1(n12365), .A2(n11162), .ZN(n8967) );
  NAND4_X2 U11556 ( .A1(n8970), .A2(n8969), .A3(n8968), .A4(n8967), .ZN(n15532) );
  NAND2_X1 U11557 ( .A1(n6609), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8971) );
  MUX2_X1 U11558 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8971), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n8972) );
  AND2_X1 U11559 ( .A1(n8972), .A2(n9111), .ZN(n10166) );
  NAND2_X1 U11560 ( .A1(n10279), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8975) );
  XNOR2_X1 U11561 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8985) );
  XNOR2_X1 U11562 ( .A(n8986), .B(n8985), .ZN(n10167) );
  OR2_X1 U11563 ( .A1(n9149), .A2(n10167), .ZN(n8977) );
  OR2_X1 U11564 ( .A1(n6435), .A2(SI_3_), .ZN(n8976) );
  OAI211_X1 U11565 ( .C1(n10166), .C2(n9564), .A(n8977), .B(n8976), .ZN(n11163) );
  NAND2_X1 U11566 ( .A1(n15532), .A2(n11163), .ZN(n12409) );
  NAND2_X1 U11567 ( .A1(n9813), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8984) );
  INV_X1 U11568 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n8978) );
  OR2_X1 U11569 ( .A1(n12366), .A2(n8978), .ZN(n8983) );
  AND2_X1 U11570 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8979) );
  NOR2_X1 U11571 ( .A1(n8996), .A2(n8979), .ZN(n11329) );
  OR2_X1 U11572 ( .A1(n9425), .A2(n11329), .ZN(n8982) );
  INV_X1 U11573 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8980) );
  OR2_X1 U11574 ( .A1(n9015), .A2(n8980), .ZN(n8981) );
  OR2_X1 U11575 ( .A1(n6435), .A2(SI_4_), .ZN(n8992) );
  NAND2_X1 U11576 ( .A1(n10277), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8987) );
  XNOR2_X1 U11577 ( .A(n9007), .B(n9006), .ZN(n10184) );
  OR2_X1 U11578 ( .A1(n9149), .A2(n10184), .ZN(n8991) );
  NAND2_X1 U11579 ( .A1(n9111), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8988) );
  MUX2_X1 U11580 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8988), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8989) );
  NAND2_X1 U11581 ( .A1(n8989), .A2(n9004), .ZN(n10186) );
  NAND2_X1 U11582 ( .A1(n9024), .A2(n10186), .ZN(n8990) );
  INV_X1 U11583 ( .A(n11163), .ZN(n11037) );
  AND2_X1 U11584 ( .A1(n15532), .A2(n11037), .ZN(n11330) );
  AOI22_X1 U11585 ( .A1(n11330), .A2(n8993), .B1(n11328), .B2(n13213), .ZN(
        n8994) );
  NAND2_X1 U11586 ( .A1(n9813), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9002) );
  INV_X1 U11587 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9584) );
  OR2_X1 U11588 ( .A1(n12366), .A2(n9584), .ZN(n9001) );
  NAND2_X1 U11589 ( .A1(n8996), .A2(n8995), .ZN(n9013) );
  OR2_X1 U11590 ( .A1(n8996), .A2(n8995), .ZN(n8997) );
  AND2_X1 U11591 ( .A1(n9013), .A2(n8997), .ZN(n11260) );
  OR2_X1 U11592 ( .A1(n9425), .A2(n11260), .ZN(n9000) );
  INV_X1 U11593 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8998) );
  OR2_X1 U11594 ( .A1(n9015), .A2(n8998), .ZN(n8999) );
  NAND4_X1 U11595 ( .A1(n9002), .A2(n9001), .A3(n9000), .A4(n8999), .ZN(n13212) );
  NAND2_X1 U11596 ( .A1(n9004), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9003) );
  MUX2_X1 U11597 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9003), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n9005) );
  NAND2_X1 U11598 ( .A1(n9005), .A2(n9041), .ZN(n10746) );
  OR2_X1 U11599 ( .A1(n6435), .A2(SI_5_), .ZN(n9010) );
  NAND2_X1 U11600 ( .A1(n10289), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9008) );
  XNOR2_X1 U11601 ( .A(n9022), .B(n9021), .ZN(n10169) );
  OR2_X1 U11602 ( .A1(n9149), .A2(n10169), .ZN(n9009) );
  OAI211_X1 U11603 ( .C1(n6489), .C2(n9564), .A(n9010), .B(n9009), .ZN(n11259)
         );
  OR2_X1 U11604 ( .A1(n13212), .A2(n11259), .ZN(n12417) );
  NAND2_X1 U11605 ( .A1(n13212), .A2(n11259), .ZN(n12418) );
  NAND2_X1 U11606 ( .A1(n11253), .A2(n12547), .ZN(n11252) );
  INV_X1 U11607 ( .A(n11259), .ZN(n11187) );
  OR2_X1 U11608 ( .A1(n13212), .A2(n11187), .ZN(n9011) );
  NAND2_X1 U11609 ( .A1(n9813), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9020) );
  INV_X1 U11610 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n9012) );
  OR2_X1 U11611 ( .A1(n12366), .A2(n9012), .ZN(n9019) );
  NAND2_X1 U11612 ( .A1(n9013), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9014) );
  AND2_X1 U11613 ( .A1(n9031), .A2(n9014), .ZN(n11447) );
  OR2_X1 U11614 ( .A1(n9425), .A2(n11447), .ZN(n9018) );
  INV_X1 U11615 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9016) );
  OR2_X1 U11616 ( .A1(n12367), .A2(n9016), .ZN(n9017) );
  INV_X1 U11617 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10281) );
  XNOR2_X1 U11618 ( .A(n10275), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n9023) );
  XNOR2_X1 U11619 ( .A(n9040), .B(n9023), .ZN(n10180) );
  OR2_X1 U11620 ( .A1(n10180), .A2(n9149), .ZN(n9028) );
  NAND2_X1 U11621 ( .A1(n9041), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U11622 ( .A1(n9259), .A2(n9620), .ZN(n9027) );
  INV_X1 U11623 ( .A(SI_6_), .ZN(n10179) );
  OR2_X1 U11624 ( .A1(n6435), .A2(n10179), .ZN(n9026) );
  NAND2_X1 U11625 ( .A1(n13211), .A2(n11372), .ZN(n12424) );
  NAND2_X1 U11626 ( .A1(n9813), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9037) );
  INV_X1 U11627 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9030) );
  OR2_X1 U11628 ( .A1(n12366), .A2(n9030), .ZN(n9036) );
  AND2_X1 U11629 ( .A1(n9031), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9032) );
  NOR2_X1 U11630 ( .A1(n9060), .A2(n9032), .ZN(n11674) );
  OR2_X1 U11631 ( .A1(n9425), .A2(n11674), .ZN(n9035) );
  INV_X1 U11632 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n9033) );
  OR2_X1 U11633 ( .A1(n9015), .A2(n9033), .ZN(n9034) );
  NAND4_X1 U11634 ( .A1(n9037), .A2(n9036), .A3(n9035), .A4(n9034), .ZN(n13210) );
  NAND2_X1 U11635 ( .A1(n10245), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9038) );
  OAI21_X1 U11636 ( .B1(n9040), .B2(n9039), .A(n9038), .ZN(n9049) );
  XNOR2_X1 U11637 ( .A(n9049), .B(n9048), .ZN(n10174) );
  INV_X2 U11638 ( .A(n9149), .ZN(n12375) );
  NAND2_X1 U11639 ( .A1(n10174), .A2(n12375), .ZN(n9047) );
  INV_X1 U11640 ( .A(SI_7_), .ZN(n10173) );
  INV_X1 U11641 ( .A(n9041), .ZN(n9043) );
  INV_X1 U11642 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U11643 ( .A1(n9043), .A2(n9042), .ZN(n9053) );
  NAND2_X1 U11644 ( .A1(n9053), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9045) );
  INV_X1 U11645 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9044) );
  AOI22_X1 U11646 ( .A1(n9260), .A2(n10173), .B1(n9259), .B2(n10840), .ZN(
        n9046) );
  NAND2_X1 U11647 ( .A1(n13210), .A2(n11673), .ZN(n11783) );
  INV_X1 U11648 ( .A(n11372), .ZN(n11446) );
  NAND2_X1 U11649 ( .A1(n13211), .A2(n11446), .ZN(n11675) );
  NAND2_X1 U11650 ( .A1(n9049), .A2(n9048), .ZN(n9051) );
  NAND2_X1 U11651 ( .A1(n7902), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U11652 ( .A1(n9051), .A2(n9050), .ZN(n9069) );
  INV_X1 U11653 ( .A(n9068), .ZN(n9052) );
  XNOR2_X1 U11654 ( .A(n9069), .B(n9052), .ZN(n10187) );
  NAND2_X1 U11655 ( .A1(n10187), .A2(n12375), .ZN(n9058) );
  OAI21_X1 U11656 ( .B1(n9053), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9054) );
  MUX2_X1 U11657 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9054), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n9056) );
  NAND2_X1 U11658 ( .A1(n6854), .A2(n9055), .ZN(n9088) );
  AOI22_X1 U11659 ( .A1(n9260), .A2(SI_8_), .B1(n9259), .B2(n10945), .ZN(n9057) );
  NAND2_X1 U11660 ( .A1(n9058), .A2(n9057), .ZN(n13087) );
  INV_X1 U11661 ( .A(n13087), .ZN(n11486) );
  NAND2_X1 U11662 ( .A1(n9813), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9066) );
  INV_X1 U11663 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n9059) );
  OR2_X1 U11664 ( .A1(n12366), .A2(n9059), .ZN(n9065) );
  NOR2_X1 U11665 ( .A1(n9060), .A2(n10944), .ZN(n9061) );
  OR2_X1 U11666 ( .A1(n9077), .A2(n9061), .ZN(n13088) );
  INV_X1 U11667 ( .A(n13088), .ZN(n11781) );
  OR2_X1 U11668 ( .A1(n9425), .A2(n11781), .ZN(n9064) );
  INV_X1 U11669 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n9062) );
  OR2_X1 U11670 ( .A1(n12367), .A2(n9062), .ZN(n9063) );
  INV_X1 U11671 ( .A(n13210), .ZN(n11491) );
  AOI22_X1 U11672 ( .A1(n11486), .A2(n15509), .B1(n11491), .B2(n12428), .ZN(
        n9067) );
  NAND2_X1 U11673 ( .A1(n9070), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9071) );
  XNOR2_X1 U11674 ( .A(n9086), .B(n9085), .ZN(n10192) );
  NAND2_X1 U11675 ( .A1(n10192), .A2(n12375), .ZN(n9074) );
  NAND2_X1 U11676 ( .A1(n9088), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9072) );
  XNOR2_X1 U11677 ( .A(n9072), .B(n6651), .ZN(n11418) );
  AOI22_X1 U11678 ( .A1(n9260), .A2(n10191), .B1(n9259), .B2(n11418), .ZN(
        n9073) );
  NAND2_X1 U11679 ( .A1(n9074), .A2(n9073), .ZN(n15516) );
  NAND2_X1 U11680 ( .A1(n9814), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9082) );
  INV_X1 U11681 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15610) );
  OR2_X1 U11682 ( .A1(n12366), .A2(n15610), .ZN(n9081) );
  OR2_X1 U11683 ( .A1(n9077), .A2(n9076), .ZN(n9078) );
  AND2_X1 U11684 ( .A1(n9095), .A2(n9078), .ZN(n11506) );
  OR2_X1 U11685 ( .A1(n9425), .A2(n11506), .ZN(n9080) );
  INV_X1 U11686 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15521) );
  OR2_X1 U11687 ( .A1(n12365), .A2(n15521), .ZN(n9079) );
  NAND4_X1 U11688 ( .A1(n9082), .A2(n9081), .A3(n9080), .A4(n9079), .ZN(n13208) );
  OR2_X1 U11689 ( .A1(n15516), .A2(n13208), .ZN(n12439) );
  NAND2_X1 U11690 ( .A1(n15516), .A2(n13208), .ZN(n12440) );
  NAND2_X1 U11691 ( .A1(n15507), .A2(n15504), .ZN(n9084) );
  INV_X1 U11692 ( .A(n13208), .ZN(n11607) );
  OR2_X1 U11693 ( .A1(n15516), .A2(n11607), .ZN(n9083) );
  XNOR2_X1 U11694 ( .A(n9104), .B(n9103), .ZN(n10237) );
  NAND2_X1 U11695 ( .A1(n10237), .A2(n12375), .ZN(n9092) );
  INV_X1 U11696 ( .A(SI_10_), .ZN(n10236) );
  NAND2_X1 U11697 ( .A1(n9109), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9090) );
  INV_X1 U11698 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9089) );
  XNOR2_X1 U11699 ( .A(n9090), .B(n9089), .ZN(n11303) );
  AOI22_X1 U11700 ( .A1(n9260), .A2(n10236), .B1(n9259), .B2(n11303), .ZN(
        n9091) );
  NAND2_X1 U11701 ( .A1(n9092), .A2(n9091), .ZN(n12064) );
  NAND2_X1 U11702 ( .A1(n9093), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9101) );
  INV_X1 U11703 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n9094) );
  OR2_X1 U11704 ( .A1(n12365), .A2(n9094), .ZN(n9100) );
  NAND2_X1 U11705 ( .A1(n9095), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9096) );
  AND2_X1 U11706 ( .A1(n9116), .A2(n9096), .ZN(n12055) );
  OR2_X1 U11707 ( .A1(n9425), .A2(n12055), .ZN(n9099) );
  INV_X1 U11708 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n9097) );
  OR2_X1 U11709 ( .A1(n12367), .A2(n9097), .ZN(n9098) );
  NAND4_X1 U11710 ( .A1(n9101), .A2(n9100), .A3(n9099), .A4(n9098), .ZN(n13207) );
  OR2_X1 U11711 ( .A1(n12064), .A2(n13207), .ZN(n12444) );
  NAND2_X1 U11712 ( .A1(n12064), .A2(n13207), .ZN(n12451) );
  INV_X1 U11713 ( .A(n13207), .ZN(n15511) );
  OR2_X1 U11714 ( .A1(n12064), .A2(n15511), .ZN(n9102) );
  NAND2_X1 U11715 ( .A1(n9105), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9106) );
  XNOR2_X1 U11716 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9108) );
  XNOR2_X1 U11717 ( .A(n9126), .B(n9108), .ZN(n10249) );
  NAND2_X1 U11718 ( .A1(n10249), .A2(n12375), .ZN(n9115) );
  OAI21_X1 U11719 ( .B1(n9109), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9110) );
  MUX2_X1 U11720 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9110), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n9113) );
  AOI22_X1 U11721 ( .A1(n9260), .A2(n10248), .B1(n9259), .B2(n13222), .ZN(
        n9114) );
  NAND2_X1 U11722 ( .A1(n9115), .A2(n9114), .ZN(n12449) );
  NAND2_X1 U11723 ( .A1(n9813), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9122) );
  INV_X1 U11724 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11820) );
  OR2_X1 U11725 ( .A1(n12366), .A2(n11820), .ZN(n9121) );
  NAND2_X1 U11726 ( .A1(n9116), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U11727 ( .A1(n9136), .A2(n9117), .ZN(n13163) );
  INV_X1 U11728 ( .A(n13163), .ZN(n9118) );
  OR2_X1 U11729 ( .A1(n9425), .A2(n9118), .ZN(n9120) );
  INV_X1 U11730 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n11813) );
  OR2_X1 U11731 ( .A1(n12367), .A2(n11813), .ZN(n9119) );
  NAND2_X1 U11732 ( .A1(n10316), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U11733 ( .A1(n10408), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9142) );
  NAND2_X1 U11734 ( .A1(n10406), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9127) );
  NAND2_X1 U11735 ( .A1(n9142), .A2(n9127), .ZN(n9128) );
  NAND2_X1 U11736 ( .A1(n9129), .A2(n9128), .ZN(n9130) );
  NAND2_X1 U11737 ( .A1(n9143), .A2(n9130), .ZN(n10292) );
  MUX2_X1 U11738 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9131), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9133) );
  INV_X1 U11739 ( .A(n9164), .ZN(n9132) );
  NAND2_X1 U11740 ( .A1(n9133), .A2(n9132), .ZN(n10291) );
  INV_X1 U11741 ( .A(n10291), .ZN(n13243) );
  AOI22_X1 U11742 ( .A1(n9260), .A2(SI_12_), .B1(n9259), .B2(n13243), .ZN(
        n9134) );
  INV_X1 U11743 ( .A(n12125), .ZN(n12179) );
  AND2_X1 U11744 ( .A1(n9136), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9137) );
  OR2_X1 U11745 ( .A1(n9137), .A2(n9154), .ZN(n12182) );
  NAND2_X1 U11746 ( .A1(n9325), .A2(n12182), .ZN(n9141) );
  INV_X1 U11747 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12123) );
  OR2_X1 U11748 ( .A1(n12365), .A2(n12123), .ZN(n9140) );
  INV_X1 U11749 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12120) );
  OR2_X1 U11750 ( .A1(n12366), .A2(n12120), .ZN(n9139) );
  INV_X1 U11751 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n12117) );
  OR2_X1 U11752 ( .A1(n12367), .A2(n12117), .ZN(n9138) );
  NAND2_X1 U11753 ( .A1(n12179), .A2(n13558), .ZN(n12454) );
  NAND2_X1 U11754 ( .A1(n12125), .A2(n13161), .ZN(n12456) );
  INV_X1 U11755 ( .A(n9146), .ZN(n9147) );
  NAND2_X1 U11756 ( .A1(n9147), .A2(n7541), .ZN(n9148) );
  NAND2_X1 U11757 ( .A1(n9162), .A2(n9148), .ZN(n10404) );
  OR2_X1 U11758 ( .A1(n9164), .A2(n9165), .ZN(n9150) );
  XNOR2_X1 U11759 ( .A(n9150), .B(P3_IR_REG_13__SCAN_IN), .ZN(n13260) );
  AOI22_X1 U11760 ( .A1(n9260), .A2(SI_13_), .B1(n9259), .B2(n13260), .ZN(
        n9151) );
  OR2_X1 U11761 ( .A1(n9154), .A2(n9153), .ZN(n9155) );
  NAND2_X1 U11762 ( .A1(n9171), .A2(n9155), .ZN(n13562) );
  NAND2_X1 U11763 ( .A1(n13562), .A2(n9325), .ZN(n9159) );
  NAND2_X1 U11764 ( .A1(n9813), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9158) );
  INV_X1 U11765 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13616) );
  OR2_X1 U11766 ( .A1(n12366), .A2(n13616), .ZN(n9157) );
  INV_X1 U11767 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13690) );
  OR2_X1 U11768 ( .A1(n12367), .A2(n13690), .ZN(n9156) );
  NAND4_X1 U11769 ( .A1(n9159), .A2(n9158), .A3(n9157), .A4(n9156), .ZN(n13546) );
  NAND2_X1 U11770 ( .A1(n13692), .A2(n13546), .ZN(n9160) );
  XNOR2_X1 U11771 ( .A(n10767), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n9163) );
  XNOR2_X1 U11772 ( .A(n9178), .B(n9163), .ZN(n10467) );
  NAND2_X1 U11773 ( .A1(n10467), .A2(n12375), .ZN(n9168) );
  AND2_X1 U11774 ( .A1(n9164), .A2(n6689), .ZN(n9182) );
  OR2_X1 U11775 ( .A1(n9182), .A2(n9165), .ZN(n9166) );
  XNOR2_X1 U11776 ( .A(n9166), .B(P3_IR_REG_14__SCAN_IN), .ZN(n13286) );
  AOI22_X1 U11777 ( .A1(n9260), .A2(SI_14_), .B1(n13286), .B2(n9259), .ZN(
        n9167) );
  NAND2_X1 U11778 ( .A1(n9813), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U11779 ( .A1(n9093), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9169) );
  AND2_X1 U11780 ( .A1(n9170), .A2(n9169), .ZN(n9175) );
  NAND2_X1 U11781 ( .A1(n9171), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U11782 ( .A1(n9189), .A2(n9172), .ZN(n13550) );
  NAND2_X1 U11783 ( .A1(n13550), .A2(n9325), .ZN(n9174) );
  NAND2_X1 U11784 ( .A1(n9814), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U11785 ( .A1(n13685), .A2(n12028), .ZN(n12463) );
  NAND2_X1 U11786 ( .A1(n13685), .A2(n13559), .ZN(n9176) );
  NAND2_X1 U11787 ( .A1(n10766), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9179) );
  XNOR2_X1 U11788 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9195) );
  INV_X1 U11789 ( .A(n9195), .ZN(n9180) );
  XNOR2_X1 U11790 ( .A(n9196), .B(n9180), .ZN(n10670) );
  NAND2_X1 U11791 ( .A1(n10670), .A2(n12375), .ZN(n9188) );
  NAND2_X1 U11792 ( .A1(n9182), .A2(n9181), .ZN(n9184) );
  NAND2_X1 U11793 ( .A1(n9184), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9183) );
  MUX2_X1 U11794 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9183), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n9185) );
  NAND2_X1 U11795 ( .A1(n9185), .A2(n9199), .ZN(n10672) );
  INV_X1 U11796 ( .A(SI_15_), .ZN(n10671) );
  OAI22_X1 U11797 ( .A1(n10672), .A2(n9564), .B1(n6435), .B2(n10671), .ZN(
        n9186) );
  INV_X1 U11798 ( .A(n9186), .ZN(n9187) );
  AND2_X1 U11799 ( .A1(n9189), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9190) );
  OR2_X1 U11800 ( .A1(n9190), .A2(n9203), .ZN(n13539) );
  NAND2_X1 U11801 ( .A1(n13539), .A2(n9325), .ZN(n9193) );
  AOI22_X1 U11802 ( .A1(n9813), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n9093), .B2(
        P3_REG1_REG_15__SCAN_IN), .ZN(n9192) );
  NAND2_X1 U11803 ( .A1(n9814), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9191) );
  OR2_X1 U11804 ( .A1(n13679), .A2(n13113), .ZN(n12387) );
  NAND2_X1 U11805 ( .A1(n13679), .A2(n13113), .ZN(n12468) );
  NAND2_X1 U11806 ( .A1(n12387), .A2(n12468), .ZN(n12561) );
  INV_X1 U11807 ( .A(n13113), .ZN(n13547) );
  NAND2_X1 U11808 ( .A1(n13679), .A2(n13547), .ZN(n9194) );
  NAND2_X1 U11809 ( .A1(n10704), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9197) );
  XNOR2_X1 U11810 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9209) );
  INV_X1 U11811 ( .A(n9209), .ZN(n9198) );
  XNOR2_X1 U11812 ( .A(n9210), .B(n9198), .ZN(n10763) );
  NAND2_X1 U11813 ( .A1(n10763), .A2(n12375), .ZN(n9202) );
  NAND2_X1 U11814 ( .A1(n9199), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9200) );
  XNOR2_X1 U11815 ( .A(n9200), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13315) );
  AOI22_X1 U11816 ( .A1(n13315), .A2(n9259), .B1(n9260), .B2(SI_16_), .ZN(
        n9201) );
  NOR2_X1 U11817 ( .A1(n9203), .A2(n13110), .ZN(n9204) );
  OR2_X1 U11818 ( .A1(n9219), .A2(n9204), .ZN(n13528) );
  NAND2_X1 U11819 ( .A1(n13528), .A2(n9325), .ZN(n9207) );
  AOI22_X1 U11820 ( .A1(n9813), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n9093), .B2(
        P3_REG1_REG_16__SCAN_IN), .ZN(n9206) );
  NAND2_X1 U11821 ( .A1(n9814), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9205) );
  OR2_X1 U11822 ( .A1(n13673), .A2(n13192), .ZN(n12470) );
  INV_X1 U11823 ( .A(n13523), .ZN(n13521) );
  NAND2_X1 U11824 ( .A1(n13673), .A2(n13536), .ZN(n9208) );
  INV_X1 U11825 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10754) );
  NAND2_X1 U11826 ( .A1(n10754), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9211) );
  XNOR2_X1 U11827 ( .A(n11977), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9213) );
  XNOR2_X1 U11828 ( .A(n9231), .B(n9213), .ZN(n10930) );
  NAND2_X1 U11829 ( .A1(n10930), .A2(n12375), .ZN(n9218) );
  INV_X1 U11830 ( .A(n9238), .ZN(n9215) );
  NAND2_X1 U11831 ( .A1(n9215), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9216) );
  XNOR2_X1 U11832 ( .A(n9216), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U11833 ( .A1(n9260), .A2(SI_17_), .B1(n9259), .B2(n13338), .ZN(
        n9217) );
  OR2_X1 U11834 ( .A1(n9219), .A2(n13120), .ZN(n9220) );
  NAND2_X1 U11835 ( .A1(n9263), .A2(n9220), .ZN(n13518) );
  NAND2_X1 U11836 ( .A1(n13518), .A2(n9325), .ZN(n9225) );
  INV_X1 U11837 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13517) );
  NAND2_X1 U11838 ( .A1(n9814), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U11839 ( .A1(n9093), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9221) );
  OAI211_X1 U11840 ( .C1(n12365), .C2(n13517), .A(n9222), .B(n9221), .ZN(n9223) );
  INV_X1 U11841 ( .A(n9223), .ZN(n9224) );
  NOR2_X1 U11842 ( .A1(n13667), .A2(n13027), .ZN(n12476) );
  INV_X1 U11843 ( .A(n12476), .ZN(n9226) );
  NAND2_X1 U11844 ( .A1(n13667), .A2(n13027), .ZN(n12473) );
  INV_X1 U11845 ( .A(n13513), .ZN(n9227) );
  NAND2_X1 U11846 ( .A1(n13667), .A2(n13525), .ZN(n9228) );
  AND2_X1 U11847 ( .A1(n10956), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U11848 ( .A1(n11977), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U11849 ( .A1(n11974), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9233) );
  INV_X1 U11850 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11130) );
  NAND2_X1 U11851 ( .A1(n11130), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11852 ( .A1(n9233), .A2(n9232), .ZN(n9250) );
  INV_X1 U11853 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11424) );
  NAND2_X1 U11854 ( .A1(n11424), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9271) );
  INV_X1 U11855 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13020) );
  NAND2_X1 U11856 ( .A1(n13020), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9234) );
  OAI21_X1 U11857 ( .B1(n9236), .B2(n9235), .A(n9272), .ZN(n11151) );
  NAND2_X1 U11858 ( .A1(n11151), .A2(n12375), .ZN(n9243) );
  NAND2_X1 U11859 ( .A1(n9254), .A2(n9239), .ZN(n9257) );
  NAND2_X1 U11860 ( .A1(n9257), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9241) );
  AOI22_X1 U11861 ( .A1(n9260), .A2(n11152), .B1(n11153), .B2(n9259), .ZN(
        n9242) );
  AND2_X1 U11862 ( .A1(n9265), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9244) );
  OR2_X1 U11863 ( .A1(n9244), .A2(n9276), .ZN(n13493) );
  NAND2_X1 U11864 ( .A1(n13493), .A2(n9325), .ZN(n9249) );
  INV_X1 U11865 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13492) );
  NAND2_X1 U11866 ( .A1(n9093), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U11867 ( .A1(n9814), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9245) );
  OAI211_X1 U11868 ( .C1(n13492), .C2(n12365), .A(n9246), .B(n9245), .ZN(n9247) );
  INV_X1 U11869 ( .A(n9247), .ZN(n9248) );
  NAND2_X1 U11870 ( .A1(n9249), .A2(n9248), .ZN(n13504) );
  OR2_X1 U11871 ( .A1(n13655), .A2(n13473), .ZN(n13468) );
  NAND2_X1 U11872 ( .A1(n9251), .A2(n9250), .ZN(n9252) );
  AND2_X1 U11873 ( .A1(n9253), .A2(n9252), .ZN(n11089) );
  NAND2_X1 U11874 ( .A1(n11089), .A2(n12375), .ZN(n9262) );
  INV_X1 U11875 ( .A(n9254), .ZN(n9255) );
  NAND2_X1 U11876 ( .A1(n9255), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9256) );
  MUX2_X1 U11877 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9256), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n9258) );
  NAND2_X1 U11878 ( .A1(n9258), .A2(n9257), .ZN(n13354) );
  INV_X1 U11879 ( .A(n13354), .ZN(n9637) );
  AOI22_X1 U11880 ( .A1(n9260), .A2(SI_18_), .B1(n9637), .B2(n9259), .ZN(n9261) );
  INV_X1 U11881 ( .A(n13661), .ZN(n13178) );
  NAND2_X1 U11882 ( .A1(n9263), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U11883 ( .A1(n9265), .A2(n9264), .ZN(n13507) );
  NAND2_X1 U11884 ( .A1(n13507), .A2(n9325), .ZN(n9270) );
  INV_X1 U11885 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13506) );
  NAND2_X1 U11886 ( .A1(n9093), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U11887 ( .A1(n9814), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9266) );
  OAI211_X1 U11888 ( .C1(n12365), .C2(n13506), .A(n9267), .B(n9266), .ZN(n9268) );
  INV_X1 U11889 ( .A(n9268), .ZN(n9269) );
  NAND2_X1 U11890 ( .A1(n13178), .A2(n13515), .ZN(n12478) );
  NAND2_X1 U11891 ( .A1(n13661), .A2(n13490), .ZN(n12480) );
  NAND2_X1 U11892 ( .A1(n12478), .A2(n12480), .ZN(n13502) );
  NAND2_X1 U11893 ( .A1(n13468), .A2(n13502), .ZN(n9284) );
  OR2_X1 U11894 ( .A1(n6435), .A2(n11639), .ZN(n9273) );
  INV_X1 U11895 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n9275) );
  NOR2_X1 U11896 ( .A1(n9276), .A2(n9275), .ZN(n9277) );
  OR2_X1 U11897 ( .A1(n9292), .A2(n9277), .ZN(n13475) );
  NAND2_X1 U11898 ( .A1(n13475), .A2(n9325), .ZN(n9282) );
  INV_X1 U11899 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13477) );
  NAND2_X1 U11900 ( .A1(n9093), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U11901 ( .A1(n9814), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9278) );
  OAI211_X1 U11902 ( .C1(n12365), .C2(n13477), .A(n9279), .B(n9278), .ZN(n9280) );
  INV_X1 U11903 ( .A(n9280), .ZN(n9281) );
  NAND2_X1 U11904 ( .A1(n13655), .A2(n13504), .ZN(n12479) );
  NAND2_X1 U11905 ( .A1(n12481), .A2(n12479), .ZN(n13485) );
  OR2_X1 U11906 ( .A1(n13661), .A2(n13515), .ZN(n13482) );
  NAND2_X1 U11907 ( .A1(n13485), .A2(n13482), .ZN(n13467) );
  NOR2_X1 U11908 ( .A1(n9305), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U11909 ( .A1(n11405), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U11910 ( .A1(n11406), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U11911 ( .A1(n9302), .A2(n9303), .ZN(n9287) );
  XNOR2_X1 U11912 ( .A(n9288), .B(n9287), .ZN(n11684) );
  NAND2_X1 U11913 ( .A1(n11684), .A2(n12375), .ZN(n9290) );
  INV_X1 U11914 ( .A(SI_21_), .ZN(n11686) );
  OR2_X1 U11915 ( .A1(n6435), .A2(n11686), .ZN(n9289) );
  INV_X1 U11916 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9291) );
  OR2_X1 U11917 ( .A1(n9292), .A2(n9291), .ZN(n9293) );
  NAND2_X1 U11918 ( .A1(n9310), .A2(n9293), .ZN(n13460) );
  NAND2_X1 U11919 ( .A1(n13460), .A2(n9325), .ZN(n9298) );
  INV_X1 U11920 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U11921 ( .A1(n9813), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9295) );
  NAND2_X1 U11922 ( .A1(n9814), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9294) );
  OAI211_X1 U11923 ( .C1(n12366), .C2(n13590), .A(n9295), .B(n9294), .ZN(n9296) );
  INV_X1 U11924 ( .A(n9296), .ZN(n9297) );
  NAND2_X1 U11925 ( .A1(n13645), .A2(n13474), .ZN(n12494) );
  INV_X1 U11926 ( .A(n13474), .ZN(n13446) );
  OR2_X1 U11927 ( .A1(n13645), .A2(n13446), .ZN(n9300) );
  NAND2_X1 U11928 ( .A1(n11383), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9301) );
  NAND3_X1 U11929 ( .A1(n9302), .A2(P1_DATAO_REG_20__SCAN_IN), .A3(n11380), 
        .ZN(n9304) );
  XNOR2_X1 U11930 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .ZN(n9319) );
  INV_X1 U11931 ( .A(n9319), .ZN(n9306) );
  XNOR2_X1 U11932 ( .A(n6509), .B(n9306), .ZN(n11546) );
  NAND2_X1 U11933 ( .A1(n11546), .A2(n12375), .ZN(n9309) );
  OR2_X1 U11934 ( .A1(n6435), .A2(n9307), .ZN(n9308) );
  NAND2_X1 U11935 ( .A1(n9310), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11936 ( .A1(n9322), .A2(n9311), .ZN(n13450) );
  NAND2_X1 U11937 ( .A1(n13450), .A2(n9325), .ZN(n9316) );
  INV_X1 U11938 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U11939 ( .A1(n9814), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U11940 ( .A1(n9093), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9312) );
  OAI211_X1 U11941 ( .C1(n12365), .C2(n13449), .A(n9313), .B(n9312), .ZN(n9314) );
  INV_X1 U11942 ( .A(n9314), .ZN(n9315) );
  NAND2_X1 U11943 ( .A1(n13639), .A2(n13457), .ZN(n9317) );
  OR2_X1 U11944 ( .A1(n13639), .A2(n13457), .ZN(n9318) );
  XNOR2_X1 U11945 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9333) );
  XNOR2_X1 U11946 ( .A(n9334), .B(n9333), .ZN(n11634) );
  NAND2_X1 U11947 ( .A1(n11634), .A2(n12375), .ZN(n9321) );
  OR2_X1 U11948 ( .A1(n6435), .A2(n11636), .ZN(n9320) );
  NAND2_X1 U11949 ( .A1(n9322), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9324) );
  NOR2_X2 U11950 ( .A1(n9322), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U11951 ( .A1(n9324), .A2(n9340), .ZN(n13436) );
  NAND2_X1 U11952 ( .A1(n13436), .A2(n9325), .ZN(n9331) );
  INV_X1 U11953 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U11954 ( .A1(n9814), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U11955 ( .A1(n9093), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9326) );
  OAI211_X1 U11956 ( .C1(n12365), .C2(n9328), .A(n9327), .B(n9326), .ZN(n9329)
         );
  INV_X1 U11957 ( .A(n9329), .ZN(n9330) );
  NAND2_X1 U11958 ( .A1(n13582), .A2(n13417), .ZN(n12504) );
  NAND2_X1 U11959 ( .A1(n12498), .A2(n12504), .ZN(n12386) );
  NAND2_X1 U11960 ( .A1(n13582), .A2(n13447), .ZN(n9332) );
  NAND2_X1 U11961 ( .A1(n9334), .A2(n9333), .ZN(n9336) );
  NAND2_X1 U11962 ( .A1(n11732), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9335) );
  XNOR2_X1 U11963 ( .A(n9349), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n12295) );
  NAND2_X1 U11964 ( .A1(n12295), .A2(n12375), .ZN(n9338) );
  OR2_X1 U11965 ( .A1(n6435), .A2(n12296), .ZN(n9337) );
  NAND2_X1 U11966 ( .A1(n9813), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9346) );
  INV_X1 U11967 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n9339) );
  OR2_X1 U11968 ( .A1(n12366), .A2(n9339), .ZN(n9345) );
  NAND2_X1 U11969 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n9340), .ZN(n9341) );
  INV_X1 U11970 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n9342) );
  OR2_X1 U11971 ( .A1(n12367), .A2(n9342), .ZN(n9343) );
  AND4_X2 U11972 ( .A1(n9346), .A2(n9345), .A3(n9344), .A4(n9343), .ZN(n13428)
         );
  INV_X1 U11973 ( .A(n13428), .ZN(n13206) );
  OR2_X1 U11974 ( .A1(n13577), .A2(n13206), .ZN(n9348) );
  INV_X1 U11975 ( .A(n9350), .ZN(n9351) );
  XNOR2_X1 U11976 ( .A(n12153), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9352) );
  XNOR2_X1 U11977 ( .A(n9365), .B(n9352), .ZN(n12258) );
  NAND2_X1 U11978 ( .A1(n12258), .A2(n12375), .ZN(n9354) );
  OR2_X1 U11979 ( .A1(n6435), .A2(n12259), .ZN(n9353) );
  NAND2_X1 U11980 ( .A1(n9813), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9362) );
  INV_X1 U11981 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n9651) );
  OR2_X1 U11982 ( .A1(n12366), .A2(n9651), .ZN(n9361) );
  INV_X1 U11983 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9355) );
  AND2_X2 U11984 ( .A1(n9356), .A2(n9355), .ZN(n9370) );
  INV_X1 U11985 ( .A(n9370), .ZN(n9371) );
  NAND2_X1 U11986 ( .A1(n9357), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9358) );
  INV_X1 U11987 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n9654) );
  OR2_X1 U11988 ( .A1(n12367), .A2(n9654), .ZN(n9359) );
  NAND2_X1 U11989 ( .A1(n13403), .A2(n13385), .ZN(n9363) );
  NAND2_X1 U11990 ( .A1(n12153), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9364) );
  XNOR2_X1 U11991 ( .A(n12352), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9366) );
  XNOR2_X1 U11992 ( .A(n9380), .B(n9366), .ZN(n13715) );
  NAND2_X1 U11993 ( .A1(n13715), .A2(n12375), .ZN(n9368) );
  OR2_X1 U11994 ( .A1(n6435), .A2(n13718), .ZN(n9367) );
  NAND2_X1 U11995 ( .A1(n9093), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9376) );
  INV_X1 U11996 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13632) );
  OR2_X1 U11997 ( .A1(n12367), .A2(n13632), .ZN(n9375) );
  INV_X1 U11998 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n9369) );
  AND2_X2 U11999 ( .A1(n9370), .A2(n9369), .ZN(n9387) );
  INV_X1 U12000 ( .A(n9387), .ZN(n9388) );
  NAND2_X1 U12001 ( .A1(n9371), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9372) );
  INV_X1 U12002 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n13395) );
  OR2_X1 U12003 ( .A1(n12365), .A2(n13395), .ZN(n9373) );
  AND4_X2 U12004 ( .A1(n9376), .A2(n9375), .A3(n9374), .A4(n9373), .ZN(n13045)
         );
  OR2_X1 U12005 ( .A1(n13572), .A2(n13205), .ZN(n9377) );
  NAND2_X1 U12006 ( .A1(n13572), .A2(n13205), .ZN(n9378) );
  AND2_X1 U12007 ( .A1(n12349), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9379) );
  NAND2_X1 U12008 ( .A1(n12352), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9381) );
  XNOR2_X1 U12009 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9383) );
  NAND2_X1 U12010 ( .A1(n13711), .A2(n12375), .ZN(n9385) );
  INV_X1 U12011 ( .A(SI_27_), .ZN(n13712) );
  OR2_X1 U12012 ( .A1(n6435), .A2(n13712), .ZN(n9384) );
  NAND2_X1 U12013 ( .A1(n9093), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9393) );
  INV_X1 U12014 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n13372) );
  OR2_X1 U12015 ( .A1(n12365), .A2(n13372), .ZN(n9392) );
  INV_X1 U12016 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U12017 ( .A1(n9388), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9389) );
  INV_X1 U12018 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n10151) );
  OR2_X1 U12019 ( .A1(n12367), .A2(n10151), .ZN(n9390) );
  AND4_X2 U12020 ( .A1(n9393), .A2(n9392), .A3(n9391), .A4(n9390), .ZN(n13387)
         );
  NAND2_X1 U12021 ( .A1(n13374), .A2(n13387), .ZN(n9826) );
  NOR2_X1 U12022 ( .A1(n15166), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9395) );
  NAND2_X1 U12023 ( .A1(n15166), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9396) );
  XNOR2_X1 U12024 ( .A(n9804), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9397) );
  XNOR2_X1 U12025 ( .A(n9803), .B(n9397), .ZN(n13708) );
  NAND2_X1 U12026 ( .A1(n13708), .A2(n12375), .ZN(n9399) );
  INV_X1 U12027 ( .A(SI_28_), .ZN(n13710) );
  OR2_X1 U12028 ( .A1(n6435), .A2(n13710), .ZN(n9398) );
  NAND2_X1 U12029 ( .A1(n9093), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9405) );
  INV_X1 U12030 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n9523) );
  OR2_X1 U12031 ( .A1(n12367), .A2(n9523), .ZN(n9404) );
  OR2_X2 U12032 ( .A1(n9400), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U12033 ( .A1(n9400), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9401) );
  INV_X1 U12034 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n9502) );
  OR2_X1 U12035 ( .A1(n12365), .A2(n9502), .ZN(n9402) );
  NAND2_X1 U12036 ( .A1(n13079), .A2(n13048), .ZN(n9827) );
  AND2_X2 U12037 ( .A1(n12523), .A2(n9827), .ZN(n13072) );
  NOR2_X1 U12038 ( .A1(n13374), .A2(n13204), .ZN(n9420) );
  NOR2_X1 U12039 ( .A1(n13072), .A2(n9420), .ZN(n9406) );
  INV_X1 U12040 ( .A(n9407), .ZN(n9408) );
  NAND2_X1 U12041 ( .A1(n9411), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9410) );
  MUX2_X1 U12042 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9410), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9412) );
  NAND2_X1 U12043 ( .A1(n12573), .A2(n12582), .ZN(n9514) );
  INV_X1 U12044 ( .A(n9413), .ZN(n9414) );
  NAND2_X1 U12045 ( .A1(n9414), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9415) );
  INV_X1 U12047 ( .A(n9416), .ZN(n9440) );
  NAND2_X1 U12048 ( .A1(n9440), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9418) );
  AND2_X1 U12049 ( .A1(n12394), .A2(n9513), .ZN(n12578) );
  INV_X1 U12050 ( .A(n12578), .ZN(n9419) );
  INV_X1 U12051 ( .A(n10146), .ZN(n9421) );
  OR2_X1 U12052 ( .A1(n9423), .A2(n13714), .ZN(n9567) );
  NAND2_X1 U12053 ( .A1(n9567), .A2(n9564), .ZN(n10889) );
  INV_X1 U12054 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n9426) );
  OR2_X1 U12055 ( .A1(n12365), .A2(n9426), .ZN(n9429) );
  INV_X1 U12056 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n12611) );
  OR2_X1 U12057 ( .A1(n12366), .A2(n12611), .ZN(n9428) );
  INV_X1 U12058 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n13628) );
  OR2_X1 U12059 ( .A1(n12367), .A2(n13628), .ZN(n9427) );
  INV_X1 U12060 ( .A(n10889), .ZN(n9430) );
  INV_X1 U12061 ( .A(n15543), .ZN(n15510) );
  OAI22_X1 U12062 ( .A1(n13387), .A2(n15508), .B1(n13077), .B2(n15510), .ZN(
        n9431) );
  XNOR2_X1 U12063 ( .A(n9446), .B(P3_B_REG_SCAN_IN), .ZN(n9437) );
  NAND2_X1 U12064 ( .A1(n9437), .A2(n12260), .ZN(n9445) );
  INV_X1 U12065 ( .A(n9438), .ZN(n9439) );
  OAI21_X1 U12066 ( .B1(n9440), .B2(n9439), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9441) );
  MUX2_X1 U12067 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9441), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9443) );
  NAND2_X1 U12068 ( .A1(n9443), .A2(n9442), .ZN(n13720) );
  INV_X1 U12069 ( .A(n13720), .ZN(n9444) );
  NAND2_X1 U12070 ( .A1(n9445), .A2(n9444), .ZN(n9447) );
  NAND2_X1 U12071 ( .A1(n9446), .A2(n13720), .ZN(n10878) );
  NAND2_X1 U12072 ( .A1(n10880), .A2(n10878), .ZN(n10271) );
  NAND2_X1 U12073 ( .A1(n12260), .A2(n13720), .ZN(n9448) );
  NOR2_X1 U12074 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .ZN(
        n12004) );
  NOR4_X1 U12075 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n9452) );
  NOR4_X1 U12076 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9451) );
  NOR4_X1 U12077 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9450) );
  NAND4_X1 U12078 ( .A1(n12004), .A2(n9452), .A3(n9451), .A4(n9450), .ZN(n9458) );
  NOR4_X1 U12079 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9456) );
  NOR4_X1 U12080 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9455) );
  NOR4_X1 U12081 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9454) );
  NOR4_X1 U12082 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n9453) );
  NAND4_X1 U12083 ( .A1(n9456), .A2(n9455), .A3(n9454), .A4(n9453), .ZN(n9457)
         );
  NOR2_X1 U12084 ( .A1(n9458), .A2(n9457), .ZN(n9459) );
  NAND2_X1 U12085 ( .A1(n6505), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9461) );
  INV_X1 U12086 ( .A(n9563), .ZN(n10866) );
  AND2_X1 U12087 ( .A1(n9510), .A2(n10866), .ZN(n9462) );
  NAND2_X1 U12088 ( .A1(n10271), .A2(n10268), .ZN(n9518) );
  NAND2_X1 U12089 ( .A1(n11153), .A2(n11640), .ZN(n12537) );
  NAND2_X1 U12090 ( .A1(n12529), .A2(n12537), .ZN(n10852) );
  AND2_X1 U12091 ( .A1(n11153), .A2(n9513), .ZN(n9463) );
  NAND2_X1 U12092 ( .A1(n9463), .A2(n12582), .ZN(n9493) );
  NAND2_X1 U12093 ( .A1(n9493), .A2(n12524), .ZN(n9499) );
  AND2_X1 U12094 ( .A1(n10852), .A2(n9499), .ZN(n9466) );
  OAI22_X1 U12095 ( .A1(n15541), .A2(n9513), .B1(n12573), .B2(n9490), .ZN(
        n9464) );
  AOI21_X1 U12096 ( .B1(n9464), .B2(n12537), .A(n12529), .ZN(n9465) );
  MUX2_X1 U12097 ( .A(n9466), .B(n9465), .S(n10268), .Z(n9467) );
  MUX2_X1 U12098 ( .A(n9468), .B(n9522), .S(n15612), .Z(n9498) );
  INV_X1 U12099 ( .A(n15545), .ZN(n9469) );
  NAND2_X1 U12100 ( .A1(n15523), .A2(n12400), .ZN(n9471) );
  INV_X1 U12101 ( .A(n11328), .ZN(n12413) );
  NOR2_X1 U12102 ( .A1(n13213), .A2(n12413), .ZN(n12414) );
  INV_X1 U12103 ( .A(n12414), .ZN(n9472) );
  AND2_X1 U12104 ( .A1(n12408), .A2(n9472), .ZN(n9473) );
  NAND2_X1 U12105 ( .A1(n11444), .A2(n12552), .ZN(n11443) );
  OR2_X1 U12106 ( .A1(n13210), .A2(n12428), .ZN(n11778) );
  INV_X1 U12107 ( .A(n11778), .ZN(n9475) );
  INV_X1 U12108 ( .A(n12425), .ZN(n9474) );
  XNOR2_X1 U12109 ( .A(n15509), .B(n13087), .ZN(n12555) );
  NAND2_X1 U12110 ( .A1(n13210), .A2(n12428), .ZN(n9476) );
  INV_X1 U12111 ( .A(n12439), .ZN(n9477) );
  INV_X1 U12112 ( .A(n12451), .ZN(n9478) );
  XNOR2_X1 U12113 ( .A(n12449), .B(n13157), .ZN(n12558) );
  OR2_X1 U12114 ( .A1(n12449), .A2(n12448), .ZN(n12443) );
  NAND2_X1 U12115 ( .A1(n12111), .A2(n12559), .ZN(n9479) );
  NAND2_X1 U12116 ( .A1(n13692), .A2(n12246), .ZN(n12457) );
  NAND2_X1 U12117 ( .A1(n12029), .A2(n13546), .ZN(n12458) );
  NAND2_X1 U12118 ( .A1(n9480), .A2(n12469), .ZN(n13510) );
  INV_X1 U12119 ( .A(n12479), .ZN(n9482) );
  OR2_X1 U12120 ( .A1(n13594), .A2(n13064), .ZN(n12490) );
  NAND2_X1 U12121 ( .A1(n13639), .A2(n13429), .ZN(n12497) );
  NAND2_X1 U12122 ( .A1(n13442), .A2(n12497), .ZN(n9483) );
  AND2_X1 U12123 ( .A1(n12506), .A2(n12504), .ZN(n13378) );
  NAND2_X1 U12124 ( .A1(n12500), .A2(n12498), .ZN(n9484) );
  NAND2_X1 U12125 ( .A1(n9484), .A2(n12506), .ZN(n9485) );
  NAND2_X1 U12126 ( .A1(n12510), .A2(n9485), .ZN(n13379) );
  NAND2_X1 U12127 ( .A1(n13379), .A2(n13382), .ZN(n9486) );
  NAND2_X1 U12128 ( .A1(n13572), .A2(n13045), .ZN(n12518) );
  NAND2_X1 U12129 ( .A1(n10142), .A2(n9826), .ZN(n9487) );
  NAND2_X1 U12130 ( .A1(n12582), .A2(n11640), .ZN(n9488) );
  NAND2_X1 U12131 ( .A1(n9488), .A2(n12573), .ZN(n9489) );
  NAND2_X1 U12132 ( .A1(n9489), .A2(n12392), .ZN(n9492) );
  OAI21_X1 U12133 ( .B1(n12394), .B2(n9513), .A(n9490), .ZN(n9491) );
  NAND2_X1 U12134 ( .A1(n9492), .A2(n9491), .ZN(n10862) );
  INV_X1 U12135 ( .A(n12537), .ZN(n9512) );
  NAND3_X1 U12136 ( .A1(n10862), .A2(n9512), .A3(n15541), .ZN(n9494) );
  NOR2_X2 U12137 ( .A1(n15552), .A2(n12582), .ZN(n15596) );
  OR2_X1 U12138 ( .A1(n13435), .A2(n15596), .ZN(n9524) );
  NAND2_X1 U12139 ( .A1(n13079), .A2(n13617), .ZN(n9495) );
  NAND2_X1 U12140 ( .A1(n9498), .A2(n9497), .ZN(P3_U3487) );
  XNOR2_X1 U12141 ( .A(n10268), .B(n9499), .ZN(n9500) );
  NAND3_X1 U12142 ( .A1(n9501), .A2(n10852), .A3(n9500), .ZN(n9504) );
  MUX2_X1 U12143 ( .A(n9502), .B(n9522), .S(n15559), .Z(n9509) );
  NOR2_X1 U12144 ( .A1(n15552), .A2(n12392), .ZN(n15538) );
  NOR2_X1 U12145 ( .A1(n13435), .A2(n15538), .ZN(n9503) );
  INV_X1 U12146 ( .A(n9505), .ZN(n13074) );
  AOI22_X1 U12147 ( .A1(n13079), .A2(n6428), .B1(n15518), .B2(n13074), .ZN(
        n9506) );
  NAND2_X1 U12148 ( .A1(n9509), .A2(n9508), .ZN(P3_U3205) );
  NAND2_X1 U12149 ( .A1(n12529), .A2(n9512), .ZN(n10846) );
  NAND2_X1 U12150 ( .A1(n12392), .A2(n9513), .ZN(n12575) );
  OR2_X1 U12151 ( .A1(n9514), .A2(n12575), .ZN(n10863) );
  NOR2_X1 U12152 ( .A1(n9563), .A2(n10863), .ZN(n9515) );
  OR2_X1 U12153 ( .A1(n12580), .A2(n9515), .ZN(n9516) );
  NAND2_X1 U12154 ( .A1(n10868), .A2(n9516), .ZN(n9521) );
  INV_X1 U12155 ( .A(n10862), .ZN(n10858) );
  OR2_X1 U12156 ( .A1(n9563), .A2(n10858), .ZN(n9519) );
  INV_X1 U12157 ( .A(n9524), .ZN(n9525) );
  NAND2_X1 U12158 ( .A1(n13079), .A2(n13691), .ZN(n9526) );
  NOR2_X1 U12159 ( .A1(n9570), .A2(n6864), .ZN(n9531) );
  NAND2_X1 U12160 ( .A1(n9530), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9532) );
  OAI21_X1 U12161 ( .B1(n10634), .B2(n9531), .A(n9532), .ZN(n10617) );
  OR2_X2 U12162 ( .A1(n10617), .A2(n15558), .ZN(n10619) );
  OR2_X1 U12163 ( .A1(n9618), .A2(n9573), .ZN(n9533) );
  NAND2_X1 U12164 ( .A1(n10563), .A2(n9533), .ZN(n9534) );
  NAND2_X1 U12165 ( .A1(n9534), .A2(n10462), .ZN(n10772) );
  NAND2_X1 U12166 ( .A1(n10774), .A2(n10772), .ZN(n9537) );
  INV_X1 U12167 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9536) );
  XNOR2_X1 U12168 ( .A(n10186), .B(n9536), .ZN(n10771) );
  NAND2_X1 U12169 ( .A1(n9537), .A2(n10771), .ZN(n10776) );
  NAND2_X1 U12170 ( .A1(n10186), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U12171 ( .A1(n10776), .A2(n9538), .ZN(n9540) );
  INV_X1 U12172 ( .A(n9540), .ZN(n9539) );
  NAND2_X1 U12173 ( .A1(n10742), .A2(n9542), .ZN(n10818) );
  NAND2_X1 U12174 ( .A1(n10822), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9545) );
  INV_X1 U12175 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U12176 ( .A1(n9620), .A2(n9543), .ZN(n9544) );
  AND2_X1 U12177 ( .A1(n9545), .A2(n9544), .ZN(n10819) );
  NAND2_X1 U12178 ( .A1(n10818), .A2(n10819), .ZN(n10817) );
  NAND2_X1 U12179 ( .A1(n10817), .A2(n9545), .ZN(n9546) );
  NAND2_X1 U12180 ( .A1(n9546), .A2(n10840), .ZN(n9547) );
  INV_X1 U12181 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10837) );
  INV_X1 U12182 ( .A(n9547), .ZN(n9548) );
  NAND2_X1 U12183 ( .A1(n10188), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9549) );
  OAI21_X1 U12184 ( .B1(n10188), .B2(P3_REG2_REG_8__SCAN_IN), .A(n9549), .ZN(
        n10943) );
  INV_X1 U12185 ( .A(n9549), .ZN(n9550) );
  INV_X1 U12186 ( .A(n9552), .ZN(n11306) );
  XNOR2_X1 U12187 ( .A(n11303), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n11307) );
  INV_X1 U12188 ( .A(n13222), .ZN(n9624) );
  INV_X1 U12189 ( .A(n9553), .ZN(n13230) );
  XNOR2_X1 U12190 ( .A(n10291), .B(P3_REG2_REG_12__SCAN_IN), .ZN(n13231) );
  INV_X1 U12191 ( .A(n13260), .ZN(n10403) );
  INV_X1 U12192 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13561) );
  INV_X1 U12193 ( .A(n13286), .ZN(n10468) );
  NAND2_X1 U12194 ( .A1(n10468), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9602) );
  INV_X1 U12195 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13549) );
  NAND2_X1 U12196 ( .A1(n13286), .A2(n13549), .ZN(n9554) );
  AND2_X1 U12197 ( .A1(n9602), .A2(n9554), .ZN(n13274) );
  NAND2_X1 U12198 ( .A1(n13272), .A2(n9602), .ZN(n9555) );
  NAND2_X1 U12199 ( .A1(n9555), .A2(n10672), .ZN(n9556) );
  INV_X1 U12200 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13538) );
  INV_X1 U12201 ( .A(n9556), .ZN(n13320) );
  XNOR2_X1 U12202 ( .A(n13315), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13319) );
  INV_X1 U12203 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U12204 ( .A1(n13323), .A2(n9557), .ZN(n9558) );
  INV_X1 U12205 ( .A(n9559), .ZN(n13347) );
  NAND2_X1 U12206 ( .A1(n13354), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9561) );
  OAI21_X1 U12207 ( .B1(n13354), .B2(P3_REG2_REG_18__SCAN_IN), .A(n9561), .ZN(
        n9560) );
  INV_X1 U12208 ( .A(n9560), .ZN(n13346) );
  XNOR2_X1 U12209 ( .A(n11153), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n9608) );
  XNOR2_X1 U12210 ( .A(n9562), .B(n9608), .ZN(n9645) );
  INV_X1 U12211 ( .A(n10853), .ZN(n9565) );
  NAND2_X1 U12212 ( .A1(n9565), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12584) );
  NAND2_X1 U12213 ( .A1(n9563), .A2(n12584), .ZN(n9612) );
  OAI21_X1 U12214 ( .B1(n9565), .B2(n12524), .A(n9564), .ZN(n9611) );
  INV_X1 U12215 ( .A(n9611), .ZN(n9566) );
  NAND2_X1 U12216 ( .A1(n9612), .A2(n9566), .ZN(n9641) );
  MUX2_X1 U12217 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13714), .Z(n9607) );
  INV_X1 U12218 ( .A(n10186), .ZN(n10785) );
  MUX2_X1 U12219 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13714), .Z(n9582) );
  INV_X1 U12220 ( .A(n9582), .ZN(n9583) );
  MUX2_X1 U12221 ( .A(n9570), .B(n9569), .S(n13714), .Z(n10664) );
  NAND2_X1 U12222 ( .A1(n10664), .A2(n6864), .ZN(n10663) );
  INV_X1 U12223 ( .A(n9571), .ZN(n10572) );
  INV_X1 U12224 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9572) );
  MUX2_X1 U12225 ( .A(n9573), .B(n9572), .S(n13714), .Z(n9574) );
  NAND2_X1 U12226 ( .A1(n9574), .A2(n9618), .ZN(n10457) );
  INV_X1 U12227 ( .A(n9574), .ZN(n9575) );
  INV_X1 U12228 ( .A(n9618), .ZN(n10580) );
  NAND2_X1 U12229 ( .A1(n9575), .A2(n10580), .ZN(n9576) );
  AND2_X1 U12230 ( .A1(n10457), .A2(n9576), .ZN(n10571) );
  OAI21_X1 U12231 ( .B1(n10620), .B2(n10572), .A(n10571), .ZN(n10570) );
  INV_X1 U12232 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10450) );
  MUX2_X1 U12233 ( .A(n11162), .B(n10450), .S(n13714), .Z(n9577) );
  NAND2_X1 U12234 ( .A1(n9577), .A2(n10166), .ZN(n9580) );
  INV_X1 U12235 ( .A(n9577), .ZN(n9578) );
  NAND2_X1 U12236 ( .A1(n9578), .A2(n10462), .ZN(n9579) );
  NAND2_X1 U12237 ( .A1(n9580), .A2(n9579), .ZN(n10456) );
  INV_X1 U12238 ( .A(n9580), .ZN(n9581) );
  XNOR2_X1 U12239 ( .A(n9582), .B(n10186), .ZN(n10769) );
  INV_X1 U12240 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11258) );
  MUX2_X1 U12241 ( .A(n11258), .B(n9584), .S(n13714), .Z(n9585) );
  NOR2_X1 U12242 ( .A1(n9585), .A2(n6489), .ZN(n10738) );
  NAND2_X1 U12243 ( .A1(n9585), .A2(n6489), .ZN(n10736) );
  OAI21_X1 U12244 ( .B1(n10740), .B2(n10738), .A(n10736), .ZN(n10815) );
  MUX2_X1 U12245 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13714), .Z(n9586) );
  XNOR2_X1 U12246 ( .A(n9586), .B(n9620), .ZN(n10816) );
  INV_X1 U12247 ( .A(n9586), .ZN(n9587) );
  AOI22_X1 U12248 ( .A1(n10815), .A2(n10816), .B1(n9620), .B2(n9587), .ZN(
        n10834) );
  MUX2_X1 U12249 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13714), .Z(n9588) );
  XNOR2_X1 U12250 ( .A(n9588), .B(n10840), .ZN(n10833) );
  MUX2_X1 U12251 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13714), .Z(n9589) );
  XNOR2_X1 U12252 ( .A(n9589), .B(n10945), .ZN(n10940) );
  INV_X1 U12253 ( .A(n9589), .ZN(n9590) );
  MUX2_X1 U12254 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13714), .Z(n9592) );
  INV_X1 U12255 ( .A(n9592), .ZN(n9591) );
  NAND2_X1 U12256 ( .A1(n9591), .A2(n9623), .ZN(n11410) );
  MUX2_X1 U12257 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13714), .Z(n9593) );
  NOR2_X1 U12258 ( .A1(n9593), .A2(n11303), .ZN(n9594) );
  AOI21_X1 U12259 ( .B1(n9593), .B2(n11303), .A(n9594), .ZN(n11300) );
  INV_X1 U12260 ( .A(n9594), .ZN(n9595) );
  NAND2_X1 U12261 ( .A1(n11298), .A2(n9595), .ZN(n13219) );
  MUX2_X1 U12262 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13714), .Z(n9596) );
  XOR2_X1 U12263 ( .A(n13222), .B(n9596), .Z(n13218) );
  INV_X1 U12264 ( .A(n9596), .ZN(n9597) );
  NAND2_X1 U12265 ( .A1(n9597), .A2(n9624), .ZN(n13237) );
  MUX2_X1 U12266 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13714), .Z(n9598) );
  XNOR2_X1 U12267 ( .A(n9598), .B(n13243), .ZN(n13236) );
  NAND2_X1 U12268 ( .A1(n9598), .A2(n10291), .ZN(n13254) );
  MUX2_X1 U12269 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13714), .Z(n9599) );
  XNOR2_X1 U12270 ( .A(n9599), .B(n13260), .ZN(n13253) );
  INV_X1 U12271 ( .A(n9599), .ZN(n9600) );
  NAND2_X1 U12272 ( .A1(n9600), .A2(n13260), .ZN(n13268) );
  NAND2_X1 U12273 ( .A1(n10468), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9630) );
  INV_X1 U12274 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U12275 ( .A1(n13286), .A2(n13613), .ZN(n9601) );
  AND2_X1 U12276 ( .A1(n9630), .A2(n9601), .ZN(n13280) );
  MUX2_X1 U12277 ( .A(n13274), .B(n13280), .S(n13714), .Z(n13267) );
  MUX2_X1 U12278 ( .A(n9602), .B(n9630), .S(n13714), .Z(n9603) );
  NAND2_X1 U12279 ( .A1(n13271), .A2(n9603), .ZN(n9604) );
  INV_X1 U12280 ( .A(n9604), .ZN(n9605) );
  INV_X1 U12281 ( .A(n10672), .ZN(n13304) );
  MUX2_X1 U12282 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13714), .Z(n13299) );
  INV_X1 U12283 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13607) );
  MUX2_X1 U12284 ( .A(n13527), .B(n13607), .S(n13714), .Z(n9606) );
  NOR2_X1 U12285 ( .A1(n13315), .A2(n9606), .ZN(n13312) );
  NAND2_X1 U12286 ( .A1(n13315), .A2(n9606), .ZN(n13310) );
  XOR2_X1 U12287 ( .A(n13338), .B(n9607), .Z(n13336) );
  NOR2_X1 U12288 ( .A1(n13335), .A2(n13336), .ZN(n13334) );
  MUX2_X1 U12289 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13714), .Z(n13345) );
  XNOR2_X1 U12290 ( .A(n11153), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n9638) );
  MUX2_X1 U12291 ( .A(n9608), .B(n9638), .S(n13714), .Z(n9609) );
  XNOR2_X1 U12292 ( .A(n9610), .B(n9609), .ZN(n9615) );
  INV_X1 U12293 ( .A(n9423), .ZN(n12579) );
  MUX2_X1 U12294 ( .A(n13214), .B(n9641), .S(n9423), .Z(n13355) );
  NAND2_X1 U12295 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13062)
         );
  NAND2_X1 U12296 ( .A1(n15503), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n9613) );
  OAI211_X1 U12297 ( .C1(n13355), .C2(n11153), .A(n13062), .B(n9613), .ZN(
        n9614) );
  XNOR2_X1 U12298 ( .A(n13315), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13308) );
  INV_X1 U12299 ( .A(n6864), .ZN(n10669) );
  AOI21_X1 U12300 ( .B1(P3_REG1_REG_0__SCAN_IN), .B2(n10669), .A(n10634), .ZN(
        n9616) );
  NOR3_X1 U12301 ( .A1(n9569), .A2(P3_IR_REG_1__SCAN_IN), .A3(n6864), .ZN(
        n9617) );
  NOR2_X1 U12302 ( .A1(n9616), .A2(n9617), .ZN(n10628) );
  MUX2_X1 U12303 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n9572), .S(n9618), .Z(n10568) );
  MUX2_X1 U12304 ( .A(n8978), .B(P3_REG1_REG_4__SCAN_IN), .S(n10186), .Z(
        n10781) );
  MUX2_X1 U12305 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n9012), .S(n9620), .Z(n10825) );
  XNOR2_X1 U12306 ( .A(n9621), .B(n10840), .ZN(n10832) );
  INV_X1 U12307 ( .A(n9621), .ZN(n9622) );
  MUX2_X1 U12308 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n9059), .S(n10945), .Z(
        n10939) );
  XOR2_X1 U12309 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n11303), .Z(n11297) );
  OR2_X1 U12310 ( .A1(n9625), .A2(n9624), .ZN(n9626) );
  XNOR2_X1 U12311 ( .A(n9625), .B(n13222), .ZN(n13216) );
  NAND2_X1 U12312 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n13216), .ZN(n13215) );
  NAND2_X1 U12313 ( .A1(n9626), .A2(n13215), .ZN(n13245) );
  AOI22_X1 U12314 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10291), .B1(n13243), 
        .B2(n12120), .ZN(n13246) );
  NAND2_X1 U12315 ( .A1(n13245), .A2(n13246), .ZN(n13244) );
  NAND2_X1 U12316 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10291), .ZN(n9627) );
  NAND2_X1 U12317 ( .A1(n9628), .A2(n10403), .ZN(n9629) );
  XNOR2_X1 U12318 ( .A(n9628), .B(n13260), .ZN(n13262) );
  NAND2_X1 U12319 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n13262), .ZN(n13261) );
  NAND2_X1 U12320 ( .A1(n10672), .A2(n9631), .ZN(n9632) );
  NAND2_X1 U12321 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n13292), .ZN(n13291) );
  NAND2_X1 U12322 ( .A1(n9632), .A2(n13291), .ZN(n13309) );
  NAND2_X1 U12323 ( .A1(n13308), .A2(n13309), .ZN(n13307) );
  INV_X1 U12324 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13604) );
  INV_X1 U12325 ( .A(n9635), .ZN(n9636) );
  OAI22_X1 U12326 ( .A1(n13330), .A2(n13604), .B1(n13338), .B2(n9636), .ZN(
        n13351) );
  XNOR2_X1 U12327 ( .A(n9637), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U12328 ( .A1(n13351), .A2(n13350), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n13354), .ZN(n9639) );
  XNOR2_X1 U12329 ( .A(n9639), .B(n9638), .ZN(n9643) );
  INV_X1 U12330 ( .A(n13714), .ZN(n9640) );
  OAI211_X1 U12331 ( .C1(n9645), .C2(n13341), .A(n9644), .B(n7739), .ZN(
        P3_U3201) );
  NAND3_X1 U12332 ( .A1(n13427), .A2(n13412), .A3(n12498), .ZN(n13411) );
  NAND2_X1 U12333 ( .A1(n13411), .A2(n12506), .ZN(n9646) );
  INV_X1 U12334 ( .A(n13406), .ZN(n9650) );
  INV_X1 U12335 ( .A(n13435), .ZN(n15551) );
  AOI22_X1 U12336 ( .A1(n15546), .A2(n13206), .B1(n13205), .B2(n15543), .ZN(
        n9649) );
  OAI211_X1 U12337 ( .C1(n6602), .C2(n12566), .A(n9647), .B(n10147), .ZN(n9648) );
  MUX2_X1 U12338 ( .A(n9651), .B(n9653), .S(n15612), .Z(n9652) );
  INV_X1 U12339 ( .A(n13403), .ZN(n9655) );
  NAND2_X1 U12340 ( .A1(n9652), .A2(n7746), .ZN(P3_U3484) );
  NAND2_X1 U12341 ( .A1(n9656), .A2(n7734), .ZN(P3_U3452) );
  XNOR2_X1 U12342 ( .A(n13970), .B(n9771), .ZN(n9760) );
  AND2_X1 U12343 ( .A1(n13842), .A2(n9716), .ZN(n13758) );
  NAND2_X1 U12344 ( .A1(n9760), .A2(n13758), .ZN(n9658) );
  XNOR2_X1 U12345 ( .A(n14138), .B(n12992), .ZN(n13754) );
  AND2_X1 U12346 ( .A1(n13843), .A2(n9716), .ZN(n13755) );
  NAND2_X1 U12347 ( .A1(n13754), .A2(n13755), .ZN(n13756) );
  AND2_X1 U12348 ( .A1(n9658), .A2(n13756), .ZN(n9758) );
  INV_X1 U12349 ( .A(n9758), .ZN(n9766) );
  XNOR2_X1 U12350 ( .A(n14147), .B(n9777), .ZN(n13724) );
  OR2_X1 U12351 ( .A1(n13791), .A2(n11066), .ZN(n13723) );
  NAND2_X1 U12352 ( .A1(n13724), .A2(n13723), .ZN(n9765) );
  XNOR2_X1 U12353 ( .A(n9726), .B(n12666), .ZN(n9660) );
  NAND2_X1 U12354 ( .A1(n9716), .A2(n13866), .ZN(n9661) );
  XNOR2_X1 U12355 ( .A(n9660), .B(n9661), .ZN(n11203) );
  NAND2_X1 U12356 ( .A1(n9726), .A2(n11173), .ZN(n9659) );
  AND2_X1 U12357 ( .A1(n11070), .A2(n9784), .ZN(n10997) );
  NOR2_X1 U12358 ( .A1(n12663), .A2(n10997), .ZN(n11064) );
  NAND2_X1 U12359 ( .A1(n9659), .A2(n11064), .ZN(n11204) );
  NAND2_X1 U12360 ( .A1(n11203), .A2(n11204), .ZN(n9664) );
  INV_X1 U12361 ( .A(n9660), .ZN(n9662) );
  NAND2_X1 U12362 ( .A1(n9662), .A2(n9661), .ZN(n9663) );
  NAND2_X1 U12363 ( .A1(n9664), .A2(n9663), .ZN(n11049) );
  XNOR2_X1 U12364 ( .A(n9726), .B(n12670), .ZN(n9665) );
  NAND2_X1 U12365 ( .A1(n9716), .A2(n13865), .ZN(n9666) );
  XNOR2_X1 U12366 ( .A(n9665), .B(n9666), .ZN(n11048) );
  INV_X1 U12367 ( .A(n9665), .ZN(n9667) );
  NAND2_X1 U12368 ( .A1(n9667), .A2(n9666), .ZN(n9668) );
  XNOR2_X1 U12369 ( .A(n9726), .B(n15471), .ZN(n9669) );
  INV_X1 U12370 ( .A(n11316), .ZN(n13864) );
  AND2_X1 U12371 ( .A1(n9716), .A2(n13864), .ZN(n9670) );
  NAND2_X1 U12372 ( .A1(n9669), .A2(n9670), .ZN(n9673) );
  INV_X1 U12373 ( .A(n9669), .ZN(n11313) );
  INV_X1 U12374 ( .A(n9670), .ZN(n9671) );
  NAND2_X1 U12375 ( .A1(n11313), .A2(n9671), .ZN(n9672) );
  NAND2_X1 U12376 ( .A1(n9673), .A2(n9672), .ZN(n15328) );
  NAND2_X1 U12377 ( .A1(n9716), .A2(n13863), .ZN(n9675) );
  XNOR2_X1 U12378 ( .A(n12927), .B(n9675), .ZN(n11323) );
  AND2_X1 U12379 ( .A1(n11323), .A2(n9673), .ZN(n9674) );
  INV_X1 U12380 ( .A(n12927), .ZN(n9676) );
  NAND2_X1 U12381 ( .A1(n9676), .A2(n9675), .ZN(n9677) );
  NAND2_X1 U12382 ( .A1(n11315), .A2(n9677), .ZN(n9678) );
  XNOR2_X1 U12383 ( .A(n9771), .B(n12933), .ZN(n9679) );
  NAND2_X1 U12384 ( .A1(n9716), .A2(n13862), .ZN(n9680) );
  XNOR2_X1 U12385 ( .A(n9679), .B(n9680), .ZN(n12928) );
  INV_X1 U12386 ( .A(n9679), .ZN(n9681) );
  NAND2_X1 U12387 ( .A1(n9681), .A2(n9680), .ZN(n9682) );
  NAND2_X1 U12388 ( .A1(n12935), .A2(n9682), .ZN(n11555) );
  XNOR2_X1 U12389 ( .A(n12992), .B(n12692), .ZN(n9683) );
  AND2_X1 U12390 ( .A1(n9716), .A2(n13861), .ZN(n9684) );
  NAND2_X1 U12391 ( .A1(n9683), .A2(n9684), .ZN(n9689) );
  INV_X1 U12392 ( .A(n9683), .ZN(n11386) );
  INV_X1 U12393 ( .A(n9684), .ZN(n9685) );
  NAND2_X1 U12394 ( .A1(n11386), .A2(n9685), .ZN(n9686) );
  NAND2_X1 U12395 ( .A1(n9689), .A2(n9686), .ZN(n11556) );
  XNOR2_X1 U12396 ( .A(n9771), .B(n12700), .ZN(n9690) );
  AND2_X1 U12397 ( .A1(n9716), .A2(n13860), .ZN(n9691) );
  NAND2_X1 U12398 ( .A1(n9690), .A2(n9691), .ZN(n9694) );
  INV_X1 U12399 ( .A(n9690), .ZN(n11577) );
  INV_X1 U12400 ( .A(n9691), .ZN(n9692) );
  NAND2_X1 U12401 ( .A1(n11577), .A2(n9692), .ZN(n9693) );
  AND2_X1 U12402 ( .A1(n9694), .A2(n9693), .ZN(n11384) );
  XNOR2_X1 U12403 ( .A(n14217), .B(n12992), .ZN(n12589) );
  NAND2_X1 U12404 ( .A1(n9716), .A2(n13859), .ZN(n9695) );
  XNOR2_X1 U12405 ( .A(n12589), .B(n9695), .ZN(n11590) );
  INV_X1 U12406 ( .A(n12589), .ZN(n9696) );
  NAND2_X1 U12407 ( .A1(n9696), .A2(n9695), .ZN(n9697) );
  NAND2_X1 U12408 ( .A1(n11581), .A2(n9697), .ZN(n9698) );
  XNOR2_X1 U12409 ( .A(n12706), .B(n9771), .ZN(n9699) );
  NAND2_X1 U12410 ( .A1(n9716), .A2(n13857), .ZN(n9700) );
  XNOR2_X1 U12411 ( .A(n9699), .B(n9700), .ZN(n12590) );
  INV_X1 U12412 ( .A(n9699), .ZN(n9701) );
  NAND2_X1 U12413 ( .A1(n9701), .A2(n9700), .ZN(n9702) );
  XNOR2_X1 U12414 ( .A(n12711), .B(n9771), .ZN(n9703) );
  AND2_X1 U12415 ( .A1(n9716), .A2(n13856), .ZN(n9704) );
  NAND2_X1 U12416 ( .A1(n9703), .A2(n9704), .ZN(n9707) );
  INV_X1 U12417 ( .A(n9703), .ZN(n12263) );
  INV_X1 U12418 ( .A(n9704), .ZN(n9705) );
  NAND2_X1 U12419 ( .A1(n12263), .A2(n9705), .ZN(n9706) );
  NAND2_X1 U12420 ( .A1(n9707), .A2(n9706), .ZN(n12191) );
  XNOR2_X1 U12421 ( .A(n14212), .B(n9771), .ZN(n9709) );
  NAND2_X1 U12422 ( .A1(n9716), .A2(n13855), .ZN(n9710) );
  XNOR2_X1 U12423 ( .A(n9709), .B(n9710), .ZN(n12273) );
  AND2_X1 U12424 ( .A1(n12273), .A2(n9707), .ZN(n9708) );
  INV_X1 U12425 ( .A(n9709), .ZN(n12633) );
  XNOR2_X1 U12426 ( .A(n12733), .B(n9771), .ZN(n9712) );
  NAND2_X1 U12427 ( .A1(n9716), .A2(n13854), .ZN(n9713) );
  XNOR2_X1 U12428 ( .A(n9712), .B(n9713), .ZN(n12632) );
  INV_X1 U12429 ( .A(n9712), .ZN(n9714) );
  NAND2_X1 U12430 ( .A1(n9714), .A2(n9713), .ZN(n9715) );
  NAND2_X1 U12431 ( .A1(n12639), .A2(n9715), .ZN(n13782) );
  XNOR2_X1 U12432 ( .A(n14206), .B(n12992), .ZN(n9717) );
  AND2_X1 U12433 ( .A1(n9716), .A2(n13853), .ZN(n9718) );
  NAND2_X1 U12434 ( .A1(n9717), .A2(n9718), .ZN(n9721) );
  INV_X1 U12435 ( .A(n9717), .ZN(n13009) );
  INV_X1 U12436 ( .A(n9718), .ZN(n9719) );
  NAND2_X1 U12437 ( .A1(n13009), .A2(n9719), .ZN(n9720) );
  NAND2_X1 U12438 ( .A1(n9721), .A2(n9720), .ZN(n13783) );
  OR2_X2 U12439 ( .A1(n13782), .A2(n13783), .ZN(n13007) );
  XNOR2_X1 U12440 ( .A(n14201), .B(n9771), .ZN(n9722) );
  NAND2_X1 U12441 ( .A1(n9716), .A2(n13852), .ZN(n9723) );
  XNOR2_X1 U12442 ( .A(n9722), .B(n9723), .ZN(n13011) );
  INV_X1 U12443 ( .A(n9722), .ZN(n9724) );
  NAND2_X1 U12444 ( .A1(n9724), .A2(n9723), .ZN(n9725) );
  XNOR2_X1 U12445 ( .A(n14086), .B(n9777), .ZN(n12602) );
  NAND2_X1 U12446 ( .A1(n13850), .A2(n9716), .ZN(n12601) );
  AND2_X1 U12447 ( .A1(n12602), .A2(n12601), .ZN(n9728) );
  XNOR2_X1 U12448 ( .A(n13831), .B(n9777), .ZN(n12600) );
  NAND2_X1 U12449 ( .A1(n9716), .A2(n13851), .ZN(n9729) );
  AND2_X1 U12450 ( .A1(n12600), .A2(n9729), .ZN(n9727) );
  XNOR2_X1 U12451 ( .A(n14181), .B(n12992), .ZN(n9736) );
  NAND2_X1 U12452 ( .A1(n13849), .A2(n9716), .ZN(n9737) );
  XNOR2_X1 U12453 ( .A(n9736), .B(n9737), .ZN(n12604) );
  INV_X1 U12454 ( .A(n9728), .ZN(n9730) );
  INV_X1 U12455 ( .A(n9729), .ZN(n12598) );
  INV_X1 U12456 ( .A(n12600), .ZN(n12597) );
  NAND3_X1 U12457 ( .A1(n9730), .A2(n12598), .A3(n12597), .ZN(n9733) );
  INV_X1 U12458 ( .A(n12602), .ZN(n12603) );
  INV_X1 U12459 ( .A(n12601), .ZN(n9731) );
  NAND2_X1 U12460 ( .A1(n12603), .A2(n9731), .ZN(n9732) );
  AND3_X1 U12461 ( .A1(n12604), .A2(n9733), .A3(n9732), .ZN(n9734) );
  INV_X1 U12462 ( .A(n9736), .ZN(n9738) );
  XNOR2_X1 U12463 ( .A(n14048), .B(n9771), .ZN(n12640) );
  NOR2_X1 U12464 ( .A1(n12645), .A2(n11066), .ZN(n9739) );
  NAND2_X1 U12465 ( .A1(n12640), .A2(n9739), .ZN(n9743) );
  INV_X1 U12466 ( .A(n12640), .ZN(n9741) );
  INV_X1 U12467 ( .A(n9739), .ZN(n9740) );
  NAND2_X1 U12468 ( .A1(n9741), .A2(n9740), .ZN(n9742) );
  NAND2_X1 U12469 ( .A1(n9743), .A2(n9742), .ZN(n13797) );
  XNOR2_X1 U12470 ( .A(n14163), .B(n9771), .ZN(n9745) );
  NAND2_X1 U12471 ( .A1(n13847), .A2(n9716), .ZN(n9746) );
  XNOR2_X1 U12472 ( .A(n9745), .B(n9746), .ZN(n12642) );
  AND2_X1 U12473 ( .A1(n12642), .A2(n9743), .ZN(n9744) );
  INV_X1 U12474 ( .A(n9745), .ZN(n9747) );
  NAND2_X1 U12475 ( .A1(n9747), .A2(n9746), .ZN(n9748) );
  XNOR2_X1 U12476 ( .A(n14159), .B(n9777), .ZN(n9749) );
  NAND2_X1 U12477 ( .A1(n13846), .A2(n9716), .ZN(n9750) );
  AND2_X1 U12478 ( .A1(n9749), .A2(n9750), .ZN(n13766) );
  INV_X1 U12479 ( .A(n9749), .ZN(n9752) );
  INV_X1 U12480 ( .A(n9750), .ZN(n9751) );
  NAND2_X1 U12481 ( .A1(n9752), .A2(n9751), .ZN(n13767) );
  XNOR2_X1 U12482 ( .A(n14151), .B(n9771), .ZN(n9755) );
  NAND2_X1 U12483 ( .A1(n13845), .A2(n9716), .ZN(n9753) );
  XNOR2_X1 U12484 ( .A(n9755), .B(n9753), .ZN(n13732) );
  NAND2_X1 U12485 ( .A1(n13733), .A2(n13732), .ZN(n9757) );
  INV_X1 U12486 ( .A(n9753), .ZN(n9754) );
  NAND2_X1 U12487 ( .A1(n9755), .A2(n9754), .ZN(n9756) );
  OAI21_X1 U12488 ( .B1(n13724), .B2(n13723), .A(n9758), .ZN(n9759) );
  OAI21_X1 U12489 ( .B1(n13754), .B2(n13843), .A(n13758), .ZN(n9762) );
  INV_X1 U12490 ( .A(n9760), .ZN(n13759) );
  INV_X1 U12491 ( .A(n13754), .ZN(n13727) );
  OAI21_X1 U12492 ( .B1(n13842), .B2(n13843), .A(n9716), .ZN(n9761) );
  AOI22_X1 U12493 ( .A1(n9762), .A2(n13759), .B1(n13727), .B2(n9761), .ZN(
        n9763) );
  XNOR2_X1 U12494 ( .A(n14126), .B(n12992), .ZN(n9767) );
  NAND2_X1 U12495 ( .A1(n13841), .A2(n9716), .ZN(n9768) );
  XNOR2_X1 U12496 ( .A(n9767), .B(n9768), .ZN(n13739) );
  INV_X1 U12497 ( .A(n9767), .ZN(n9770) );
  INV_X1 U12498 ( .A(n9768), .ZN(n9769) );
  XNOR2_X1 U12499 ( .A(n13945), .B(n9771), .ZN(n9772) );
  NAND2_X1 U12500 ( .A1(n13840), .A2(n9716), .ZN(n9773) );
  NAND2_X1 U12501 ( .A1(n9772), .A2(n9773), .ZN(n12981) );
  INV_X1 U12502 ( .A(n9772), .ZN(n9775) );
  INV_X1 U12503 ( .A(n9773), .ZN(n9774) );
  NAND2_X1 U12504 ( .A1(n9775), .A2(n9774), .ZN(n9776) );
  AND2_X1 U12505 ( .A1(n12981), .A2(n9776), .ZN(n13809) );
  NAND2_X1 U12506 ( .A1(n13808), .A2(n12981), .ZN(n9779) );
  XNOR2_X1 U12507 ( .A(n14115), .B(n9777), .ZN(n12979) );
  NAND2_X1 U12508 ( .A1(n13839), .A2(n9716), .ZN(n12983) );
  XNOR2_X1 U12509 ( .A(n12987), .B(n12983), .ZN(n12977) );
  INV_X1 U12510 ( .A(n9780), .ZN(n9781) );
  NAND2_X1 U12511 ( .A1(n9782), .A2(n10990), .ZN(n9787) );
  NAND2_X1 U12512 ( .A1(n9784), .A2(n6993), .ZN(n11171) );
  OR2_X1 U12513 ( .A1(n9787), .A2(n11171), .ZN(n9786) );
  AOI22_X1 U12514 ( .A1(n13838), .A2(n13802), .B1(n13801), .B2(n13840), .ZN(
        n13930) );
  INV_X1 U12515 ( .A(n9787), .ZN(n9789) );
  INV_X1 U12516 ( .A(n12905), .ZN(n9788) );
  INV_X1 U12517 ( .A(n9790), .ZN(n9791) );
  NAND2_X1 U12518 ( .A1(n10990), .A2(n9791), .ZN(n9793) );
  NAND2_X1 U12519 ( .A1(n9793), .A2(n9792), .ZN(n9795) );
  NAND2_X1 U12520 ( .A1(n9795), .A2(n9794), .ZN(n11047) );
  INV_X1 U12521 ( .A(n9796), .ZN(n9797) );
  OR2_X1 U12522 ( .A1(n11047), .A2(n9797), .ZN(n9798) );
  INV_X1 U12523 ( .A(n15334), .ZN(n13804) );
  AOI22_X1 U12524 ( .A1(n13934), .A2(n13804), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9799) );
  OAI21_X1 U12525 ( .B1(n13930), .B2(n15325), .A(n9799), .ZN(n9800) );
  AOI21_X1 U12526 ( .B1(n14115), .B2(n15332), .A(n9800), .ZN(n9801) );
  INV_X1 U12527 ( .A(n13048), .ZN(n13203) );
  AOI21_X1 U12528 ( .B1(n13079), .B2(n13203), .A(n13472), .ZN(n9811) );
  NAND2_X1 U12529 ( .A1(n9804), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U12530 ( .A1(n9806), .A2(n9805), .ZN(n12358) );
  INV_X1 U12531 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14253) );
  XNOR2_X1 U12532 ( .A(n14253), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n12357) );
  INV_X1 U12533 ( .A(n12357), .ZN(n9807) );
  XNOR2_X1 U12534 ( .A(n12358), .B(n9807), .ZN(n13705) );
  NAND2_X1 U12535 ( .A1(n13705), .A2(n12375), .ZN(n9809) );
  INV_X1 U12536 ( .A(SI_29_), .ZN(n13707) );
  OR2_X1 U12537 ( .A1(n6435), .A2(n13707), .ZN(n9808) );
  INV_X1 U12538 ( .A(n12380), .ZN(n9810) );
  NAND3_X1 U12539 ( .A1(n9821), .A2(n9811), .A3(n9829), .ZN(n9824) );
  NOR2_X1 U12540 ( .A1(n13048), .A2(n13472), .ZN(n9812) );
  AND2_X1 U12541 ( .A1(n13079), .A2(n9812), .ZN(n9820) );
  NAND2_X1 U12542 ( .A1(n9813), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U12543 ( .A1(n9093), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9816) );
  NAND2_X1 U12544 ( .A1(n9814), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9815) );
  NAND2_X1 U12545 ( .A1(n12579), .A2(P3_B_REG_SCAN_IN), .ZN(n9818) );
  NAND2_X1 U12546 ( .A1(n15531), .A2(n9818), .ZN(n13362) );
  OAI22_X1 U12547 ( .A1(n12382), .A2(n13362), .B1(n13048), .B2(n15508), .ZN(
        n9819) );
  AOI21_X1 U12548 ( .B1(n12570), .B2(n9820), .A(n9819), .ZN(n9823) );
  NAND2_X1 U12549 ( .A1(n9825), .A2(n15559), .ZN(n9837) );
  NAND2_X1 U12550 ( .A1(n9827), .A2(n9826), .ZN(n12525) );
  INV_X1 U12551 ( .A(n12525), .ZN(n9828) );
  XNOR2_X1 U12552 ( .A(n12381), .B(n9829), .ZN(n13631) );
  INV_X1 U12553 ( .A(n13631), .ZN(n9835) );
  INV_X1 U12554 ( .A(n13566), .ZN(n9834) );
  NOR2_X1 U12555 ( .A1(n15553), .A2(n9830), .ZN(n13364) );
  AOI21_X1 U12556 ( .B1(n13630), .B2(n6428), .A(n13364), .ZN(n9832) );
  NAND2_X1 U12557 ( .A1(n15561), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U12558 ( .A1(n9832), .A2(n9831), .ZN(n9833) );
  NAND2_X1 U12559 ( .A1(n9837), .A2(n9836), .ZN(P3_U3204) );
  NAND2_X1 U12560 ( .A1(n12944), .A2(n10061), .ZN(n9841) );
  INV_X1 U12561 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12945) );
  INV_X1 U12562 ( .A(n9843), .ZN(n9842) );
  OAI21_X1 U12563 ( .B1(n9842), .B2(n13712), .A(n9845), .ZN(n9848) );
  NOR2_X1 U12564 ( .A1(n9843), .A2(SI_27_), .ZN(n9846) );
  AOI21_X1 U12565 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9847) );
  INV_X1 U12566 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15157) );
  MUX2_X1 U12567 ( .A(n15157), .B(n14253), .S(n10171), .Z(n10038) );
  XNOR2_X1 U12568 ( .A(n10038), .B(SI_29_), .ZN(n10036) );
  OR2_X1 U12569 ( .A1(n9865), .A2(n9851), .ZN(n9858) );
  INV_X1 U12570 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U12571 ( .A1(n7835), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U12572 ( .A1(n10029), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9853) );
  OAI211_X1 U12573 ( .C1(n9855), .C2(n7871), .A(n9854), .B(n9853), .ZN(n9856)
         );
  INV_X1 U12574 ( .A(n9856), .ZN(n9857) );
  INV_X1 U12575 ( .A(n9860), .ZN(n10376) );
  NAND4_X1 U12576 ( .A1(n10376), .A2(n9861), .A3(n10374), .A4(n10375), .ZN(
        n9871) );
  INV_X1 U12577 ( .A(n10394), .ZN(n9862) );
  NAND2_X2 U12578 ( .A1(n9871), .A2(n14997), .ZN(n15305) );
  INV_X1 U12579 ( .A(n15297), .ZN(n9863) );
  NAND2_X1 U12580 ( .A1(n10371), .A2(n9863), .ZN(n15291) );
  INV_X1 U12581 ( .A(n15291), .ZN(n9864) );
  INV_X1 U12582 ( .A(n9865), .ZN(n9874) );
  INV_X1 U12583 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14753) );
  NAND2_X1 U12584 ( .A1(n9866), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U12585 ( .A1(n10029), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9867) );
  OAI211_X1 U12586 ( .C1(n10032), .C2(n14753), .A(n9868), .B(n9867), .ZN(
        n14564) );
  NAND2_X1 U12587 ( .A1(n15261), .A2(P1_B_REG_SCAN_IN), .ZN(n9869) );
  AND2_X1 U12588 ( .A1(n15008), .A2(n9869), .ZN(n12653) );
  NAND2_X1 U12589 ( .A1(n14564), .A2(n12653), .ZN(n15031) );
  NAND3_X1 U12590 ( .A1(n9871), .A2(P1_REG2_REG_29__SCAN_IN), .A3(n14997), 
        .ZN(n9870) );
  OAI21_X1 U12591 ( .B1(n9871), .B2(n15031), .A(n9870), .ZN(n9873) );
  NOR3_X1 U12592 ( .A1(n15033), .A2(n15307), .A3(n15032), .ZN(n9872) );
  AOI211_X1 U12593 ( .C1(n15301), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9875)
         );
  OAI21_X1 U12594 ( .B1(n10027), .B2(n15279), .A(n9875), .ZN(n9876) );
  NAND2_X1 U12595 ( .A1(n14365), .A2(n14543), .ZN(n9877) );
  NAND2_X1 U12596 ( .A1(n15041), .A2(n14566), .ZN(n9880) );
  OR2_X1 U12597 ( .A1(n15041), .A2(n14566), .ZN(n9879) );
  NAND2_X1 U12598 ( .A1(n15305), .A2(n15078), .ZN(n15023) );
  NAND3_X1 U12599 ( .A1(n7748), .A2(n9883), .A3(n9882), .ZN(P1_U3356) );
  INV_X1 U12600 ( .A(n8371), .ZN(n10113) );
  INV_X2 U12601 ( .A(n9920), .ZN(n10095) );
  MUX2_X1 U12602 ( .A(n14568), .B(n9888), .S(n10095), .Z(n10020) );
  INV_X1 U12603 ( .A(n10020), .ZN(n10024) );
  OR2_X1 U12604 ( .A1(n14587), .A2(n10399), .ZN(n9889) );
  NAND2_X1 U12605 ( .A1(n10516), .A2(n9889), .ZN(n10369) );
  NAND2_X1 U12606 ( .A1(n10369), .A2(n10380), .ZN(n9897) );
  NAND3_X1 U12607 ( .A1(n8316), .A2(n9890), .A3(n9924), .ZN(n9891) );
  OAI21_X1 U12608 ( .B1(n9892), .B2(n9924), .A(n9891), .ZN(n9896) );
  NAND2_X1 U12609 ( .A1(n8316), .A2(n9898), .ZN(n9895) );
  NAND2_X1 U12610 ( .A1(n9893), .A2(n9924), .ZN(n9894) );
  NAND2_X1 U12611 ( .A1(n10530), .A2(n9898), .ZN(n9900) );
  NAND2_X1 U12612 ( .A1(n12943), .A2(n9924), .ZN(n9899) );
  MUX2_X1 U12613 ( .A(n9900), .B(n9899), .S(n14585), .Z(n9901) );
  OAI211_X1 U12614 ( .C1(n9902), .C2(n10546), .A(n10073), .B(n9901), .ZN(n9906) );
  XNOR2_X1 U12615 ( .A(n14583), .B(n15310), .ZN(n10896) );
  NAND2_X1 U12616 ( .A1(n6434), .A2(n9924), .ZN(n9904) );
  OR2_X1 U12617 ( .A1(n6434), .A2(n9924), .ZN(n9903) );
  MUX2_X1 U12618 ( .A(n9904), .B(n9903), .S(n14584), .Z(n9905) );
  OAI21_X1 U12619 ( .B1(n14583), .B2(n10095), .A(n6430), .ZN(n9909) );
  NAND2_X1 U12620 ( .A1(n14583), .A2(n9924), .ZN(n9907) );
  NAND2_X1 U12621 ( .A1(n9907), .A2(n10903), .ZN(n9908) );
  MUX2_X1 U12622 ( .A(n11284), .B(n11120), .S(n9947), .Z(n9911) );
  MUX2_X1 U12623 ( .A(n11213), .B(n14582), .S(n10095), .Z(n9910) );
  MUX2_X1 U12624 ( .A(n11429), .B(n14581), .S(n9947), .Z(n9915) );
  NAND2_X1 U12625 ( .A1(n9914), .A2(n9915), .ZN(n9913) );
  MUX2_X1 U12626 ( .A(n14581), .B(n11429), .S(n9947), .Z(n9912) );
  NAND2_X1 U12627 ( .A1(n9913), .A2(n9912), .ZN(n9919) );
  INV_X1 U12628 ( .A(n9914), .ZN(n9917) );
  INV_X1 U12629 ( .A(n9915), .ZN(n9916) );
  NAND2_X1 U12630 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  NAND2_X1 U12631 ( .A1(n9919), .A2(n9918), .ZN(n9922) );
  MUX2_X1 U12632 ( .A(n14579), .B(n11596), .S(n10095), .Z(n9923) );
  MUX2_X1 U12633 ( .A(n14579), .B(n11596), .S(n9920), .Z(n9921) );
  INV_X2 U12634 ( .A(n9924), .ZN(n10066) );
  MUX2_X1 U12635 ( .A(n14578), .B(n11723), .S(n10066), .Z(n9927) );
  MUX2_X1 U12636 ( .A(n14578), .B(n11723), .S(n9947), .Z(n9925) );
  MUX2_X1 U12637 ( .A(n14577), .B(n12044), .S(n9924), .Z(n9930) );
  MUX2_X1 U12638 ( .A(n14577), .B(n12044), .S(n10066), .Z(n9928) );
  NAND2_X1 U12639 ( .A1(n9929), .A2(n9928), .ZN(n9932) );
  MUX2_X1 U12640 ( .A(n14576), .B(n12160), .S(n10066), .Z(n9935) );
  MUX2_X1 U12641 ( .A(n14576), .B(n12160), .S(n9924), .Z(n9933) );
  MUX2_X1 U12642 ( .A(n14575), .B(n15117), .S(n10095), .Z(n9938) );
  MUX2_X1 U12643 ( .A(n14575), .B(n15117), .S(n10066), .Z(n9936) );
  MUX2_X1 U12644 ( .A(n14574), .B(n12205), .S(n10066), .Z(n9940) );
  MUX2_X1 U12645 ( .A(n14574), .B(n12205), .S(n9924), .Z(n9939) );
  XNOR2_X1 U12646 ( .A(n15112), .B(n14573), .ZN(n15020) );
  MUX2_X1 U12647 ( .A(n14386), .B(n12307), .S(n9924), .Z(n9951) );
  NAND3_X1 U12648 ( .A1(n15020), .A2(n9951), .A3(n9977), .ZN(n9944) );
  OAI21_X1 U12649 ( .B1(n9955), .B2(n15009), .A(n15003), .ZN(n9942) );
  NAND2_X1 U12650 ( .A1(n9955), .A2(n15009), .ZN(n9941) );
  NAND3_X1 U12651 ( .A1(n9942), .A2(n10066), .A3(n9941), .ZN(n9943) );
  MUX2_X1 U12652 ( .A(n14967), .B(n14955), .S(n10066), .Z(n9967) );
  NAND2_X1 U12653 ( .A1(n9967), .A2(n9972), .ZN(n9946) );
  MUX2_X1 U12654 ( .A(n14994), .B(n15105), .S(n10066), .Z(n9961) );
  MUX2_X1 U12655 ( .A(n6981), .B(n14981), .S(n9924), .Z(n9960) );
  NAND2_X1 U12656 ( .A1(n9961), .A2(n9960), .ZN(n9945) );
  AND2_X1 U12657 ( .A1(n9946), .A2(n9945), .ZN(n9980) );
  INV_X1 U12658 ( .A(n9954), .ZN(n9948) );
  NAND3_X1 U12659 ( .A1(n9950), .A2(n9980), .A3(n9949), .ZN(n9985) );
  INV_X1 U12660 ( .A(n9951), .ZN(n9952) );
  NAND2_X1 U12661 ( .A1(n9953), .A2(n9952), .ZN(n9959) );
  NAND4_X1 U12662 ( .A1(n15020), .A2(n10066), .A3(n12236), .A4(n9977), .ZN(
        n9957) );
  AND2_X1 U12663 ( .A1(n9954), .A2(n9924), .ZN(n9975) );
  NAND3_X1 U12664 ( .A1(n9955), .A2(n9975), .A3(n15011), .ZN(n9956) );
  NAND2_X1 U12665 ( .A1(n9957), .A2(n9956), .ZN(n9958) );
  NAND3_X1 U12666 ( .A1(n9959), .A2(n9980), .A3(n9958), .ZN(n9984) );
  INV_X1 U12667 ( .A(n9960), .ZN(n9963) );
  INV_X1 U12668 ( .A(n9961), .ZN(n9962) );
  NAND2_X1 U12669 ( .A1(n9963), .A2(n9962), .ZN(n9973) );
  NAND2_X1 U12670 ( .A1(n9965), .A2(n9964), .ZN(n9971) );
  NAND2_X1 U12671 ( .A1(n9973), .A2(n9966), .ZN(n9969) );
  INV_X1 U12672 ( .A(n9967), .ZN(n9968) );
  NAND2_X1 U12673 ( .A1(n9969), .A2(n9968), .ZN(n9970) );
  OAI211_X1 U12674 ( .C1(n9973), .C2(n9972), .A(n9971), .B(n9970), .ZN(n9974)
         );
  INV_X1 U12675 ( .A(n9974), .ZN(n9982) );
  INV_X1 U12676 ( .A(n9975), .ZN(n9976) );
  AOI21_X1 U12677 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n9979) );
  NAND2_X1 U12678 ( .A1(n9980), .A2(n9979), .ZN(n9981) );
  NAND3_X1 U12679 ( .A1(n9985), .A2(n9984), .A3(n9983), .ZN(n9990) );
  AND2_X1 U12680 ( .A1(n9991), .A2(n9986), .ZN(n9987) );
  MUX2_X1 U12681 ( .A(n9988), .B(n9987), .S(n10095), .Z(n9989) );
  OR2_X1 U12682 ( .A1(n15088), .A2(n14932), .ZN(n9992) );
  NAND3_X1 U12683 ( .A1(n9990), .A2(n9989), .A3(n9992), .ZN(n9994) );
  MUX2_X1 U12684 ( .A(n9992), .B(n9991), .S(n10066), .Z(n9993) );
  MUX2_X1 U12685 ( .A(n14878), .B(n14910), .S(n9924), .Z(n9995) );
  INV_X1 U12686 ( .A(n9995), .ZN(n9997) );
  MUX2_X1 U12687 ( .A(n14910), .B(n14878), .S(n9924), .Z(n9996) );
  MUX2_X1 U12688 ( .A(n14888), .B(n14901), .S(n9924), .Z(n10000) );
  MUX2_X1 U12689 ( .A(n14888), .B(n14901), .S(n10066), .Z(n9998) );
  NAND2_X1 U12690 ( .A1(n9999), .A2(n9998), .ZN(n10002) );
  NAND2_X1 U12691 ( .A1(n10002), .A2(n10001), .ZN(n10004) );
  MUX2_X1 U12692 ( .A(n14879), .B(n15068), .S(n10095), .Z(n10005) );
  MUX2_X1 U12693 ( .A(n14879), .B(n15068), .S(n10066), .Z(n10003) );
  INV_X1 U12694 ( .A(n10005), .ZN(n10006) );
  MUX2_X1 U12695 ( .A(n14571), .B(n15061), .S(n10066), .Z(n10008) );
  MUX2_X1 U12696 ( .A(n14571), .B(n15061), .S(n10095), .Z(n10007) );
  INV_X1 U12697 ( .A(n10008), .ZN(n10009) );
  MUX2_X1 U12698 ( .A(n14570), .B(n14833), .S(n10095), .Z(n10012) );
  MUX2_X1 U12699 ( .A(n14833), .B(n14570), .S(n10095), .Z(n10010) );
  INV_X1 U12700 ( .A(n10012), .ZN(n10013) );
  MUX2_X1 U12701 ( .A(n14569), .B(n15050), .S(n10066), .Z(n10016) );
  MUX2_X1 U12702 ( .A(n14569), .B(n15050), .S(n10095), .Z(n10014) );
  NAND2_X1 U12703 ( .A1(n10015), .A2(n10014), .ZN(n10018) );
  NAND2_X1 U12704 ( .A1(n10018), .A2(n10017), .ZN(n10021) );
  INV_X1 U12705 ( .A(n10021), .ZN(n10023) );
  MUX2_X1 U12706 ( .A(n15048), .B(n14455), .S(n10095), .Z(n10019) );
  AOI21_X1 U12707 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10022) );
  MUX2_X1 U12708 ( .A(n14365), .B(n14543), .S(n10095), .Z(n10069) );
  MUX2_X1 U12709 ( .A(n14543), .B(n14365), .S(n10095), .Z(n10025) );
  INV_X1 U12710 ( .A(n10025), .ZN(n10026) );
  MUX2_X1 U12711 ( .A(n14565), .B(n15036), .S(n10095), .Z(n10114) );
  INV_X1 U12712 ( .A(n10114), .ZN(n10123) );
  MUX2_X1 U12713 ( .A(n10028), .B(n10027), .S(n10066), .Z(n10115) );
  INV_X1 U12714 ( .A(n10115), .ZN(n10122) );
  NAND2_X1 U12715 ( .A1(n10261), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11734) );
  INV_X1 U12716 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n14746) );
  NAND2_X1 U12717 ( .A1(n9866), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U12718 ( .A1(n10029), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n10030) );
  OAI211_X1 U12719 ( .C1(n10032), .C2(n14746), .A(n10031), .B(n10030), .ZN(
        n14563) );
  INV_X1 U12720 ( .A(n10033), .ZN(n10034) );
  OAI21_X1 U12721 ( .B1(n14563), .B2(n10034), .A(n14564), .ZN(n10035) );
  INV_X1 U12722 ( .A(n10035), .ZN(n10045) );
  NAND2_X1 U12723 ( .A1(n10038), .A2(n13707), .ZN(n10050) );
  NAND2_X1 U12724 ( .A1(n10056), .A2(n10050), .ZN(n10042) );
  INV_X1 U12725 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12936) );
  INV_X1 U12726 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12810) );
  MUX2_X1 U12727 ( .A(n12936), .B(n12810), .S(n10039), .Z(n10040) );
  INV_X1 U12728 ( .A(SI_30_), .ZN(n12616) );
  NAND2_X1 U12729 ( .A1(n10040), .A2(n12616), .ZN(n10051) );
  AND2_X1 U12730 ( .A1(n6478), .A2(n10051), .ZN(n10041) );
  NAND2_X1 U12731 ( .A1(n12809), .A2(n10061), .ZN(n10044) );
  NAND2_X1 U12732 ( .A1(n14563), .A2(n10066), .ZN(n10047) );
  INV_X1 U12733 ( .A(n14564), .ZN(n10046) );
  AOI21_X1 U12734 ( .B1(n10048), .B2(n10047), .A(n10046), .ZN(n10049) );
  AOI21_X1 U12735 ( .B1(n14756), .B2(n10095), .A(n10049), .ZN(n10106) );
  NAND2_X1 U12736 ( .A1(n10107), .A2(n10106), .ZN(n10129) );
  NAND2_X1 U12737 ( .A1(n10051), .A2(n10050), .ZN(n10054) );
  MUX2_X1 U12738 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10171), .Z(n10052) );
  XNOR2_X1 U12739 ( .A(n10052), .B(SI_31_), .ZN(n10053) );
  NOR2_X1 U12740 ( .A1(n10054), .A2(n10053), .ZN(n10059) );
  XNOR2_X1 U12741 ( .A(n10053), .B(n6478), .ZN(n10058) );
  NOR2_X1 U12742 ( .A1(n10054), .A2(n7490), .ZN(n10055) );
  NAND2_X1 U12743 ( .A1(n10056), .A2(n10055), .ZN(n10057) );
  INV_X1 U12744 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10060) );
  XNOR2_X1 U12745 ( .A(n14748), .B(n14563), .ZN(n10072) );
  OR2_X1 U12746 ( .A1(n10379), .A2(n8398), .ZN(n10064) );
  NAND2_X1 U12747 ( .A1(n15297), .A2(n10113), .ZN(n10062) );
  NAND2_X1 U12748 ( .A1(n10062), .A2(n10262), .ZN(n10063) );
  NAND2_X1 U12749 ( .A1(n10064), .A2(n10063), .ZN(n10100) );
  INV_X1 U12750 ( .A(n10100), .ZN(n10065) );
  AND2_X1 U12751 ( .A1(n10072), .A2(n10065), .ZN(n10125) );
  NAND2_X1 U12752 ( .A1(n10129), .A2(n10125), .ZN(n10121) );
  AOI211_X1 U12753 ( .C1(n10123), .C2(n10122), .A(n11734), .B(n10121), .ZN(
        n10119) );
  MUX2_X1 U12754 ( .A(n14566), .B(n15041), .S(n10095), .Z(n10108) );
  INV_X1 U12755 ( .A(n10108), .ZN(n10068) );
  MUX2_X1 U12756 ( .A(n15033), .B(n14768), .S(n10066), .Z(n10109) );
  INV_X1 U12757 ( .A(n10109), .ZN(n10067) );
  NAND2_X1 U12758 ( .A1(n10068), .A2(n10067), .ZN(n10136) );
  NAND2_X1 U12759 ( .A1(n10119), .A2(n10136), .ZN(n10071) );
  INV_X1 U12760 ( .A(n11734), .ZN(n10139) );
  XOR2_X1 U12761 ( .A(n14564), .B(n14756), .Z(n10089) );
  INV_X1 U12762 ( .A(n10072), .ZN(n10094) );
  XNOR2_X1 U12763 ( .A(n15117), .B(n14444), .ZN(n12075) );
  NAND4_X1 U12764 ( .A1(n10073), .A2(n10548), .A3(n10517), .A4(n10369), .ZN(
        n10076) );
  INV_X1 U12765 ( .A(n10896), .ZN(n10074) );
  NOR3_X1 U12766 ( .A1(n10076), .A2(n10075), .A3(n10074), .ZN(n10077) );
  XNOR2_X1 U12767 ( .A(n11596), .B(n14579), .ZN(n11459) );
  NAND4_X1 U12768 ( .A1(n11741), .A2(n10077), .A3(n11279), .A4(n11459), .ZN(
        n10078) );
  NOR3_X1 U12769 ( .A1(n14989), .A2(n10080), .A3(n10079), .ZN(n10082) );
  NAND4_X1 U12770 ( .A1(n14911), .A2(n14856), .A3(n10084), .A4(n14924), .ZN(
        n10085) );
  NOR3_X1 U12771 ( .A1(n14817), .A2(n14869), .A3(n10085), .ZN(n10086) );
  XOR2_X1 U12772 ( .A(n15296), .B(n10091), .Z(n10103) );
  OR2_X1 U12773 ( .A1(n15297), .A2(n10092), .ZN(n10102) );
  NAND2_X1 U12774 ( .A1(n10100), .A2(n10102), .ZN(n10104) );
  INV_X1 U12775 ( .A(n10104), .ZN(n10093) );
  NAND2_X1 U12776 ( .A1(n10094), .A2(n10093), .ZN(n10099) );
  NOR2_X1 U12777 ( .A1(n12659), .A2(n14563), .ZN(n10097) );
  INV_X1 U12778 ( .A(n10105), .ZN(n10098) );
  MUX2_X1 U12779 ( .A(n10100), .B(n10099), .S(n10098), .Z(n10101) );
  OAI21_X1 U12780 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(n10138) );
  INV_X1 U12781 ( .A(n10141), .ZN(n10135) );
  NAND2_X1 U12782 ( .A1(n10109), .A2(n10108), .ZN(n10140) );
  INV_X1 U12783 ( .A(n10140), .ZN(n10120) );
  INV_X1 U12784 ( .A(P1_B_REG_SCAN_IN), .ZN(n12001) );
  INV_X1 U12785 ( .A(n10261), .ZN(n10110) );
  NAND3_X1 U12786 ( .A1(n10111), .A2(n10383), .A3(n10110), .ZN(n10396) );
  NAND2_X1 U12787 ( .A1(n15261), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15163) );
  NOR3_X1 U12788 ( .A1(n10396), .A2(n15032), .A3(n15163), .ZN(n10112) );
  AOI211_X1 U12789 ( .C1(n10139), .C2(n10113), .A(n12001), .B(n10112), .ZN(
        n10118) );
  NOR4_X1 U12790 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n11734), .ZN(
        n10117) );
  INV_X1 U12791 ( .A(n10121), .ZN(n10132) );
  NOR3_X1 U12792 ( .A1(n10123), .A2(n10122), .A3(n11734), .ZN(n10131) );
  INV_X1 U12793 ( .A(n10124), .ZN(n10128) );
  INV_X1 U12794 ( .A(n10125), .ZN(n10126) );
  OAI22_X1 U12795 ( .A1(n10129), .A2(n10128), .B1(n10127), .B2(n10126), .ZN(
        n10130) );
  AOI22_X1 U12796 ( .A1(n10132), .A2(n10131), .B1(n10139), .B2(n10130), .ZN(
        n10133) );
  OAI211_X1 U12797 ( .C1(n10136), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        n10137) );
  NAND2_X1 U12798 ( .A1(n10146), .A2(n10145), .ZN(n10148) );
  OAI22_X1 U12799 ( .A1(n13045), .A2(n15508), .B1(n13048), .B2(n15510), .ZN(
        n10149) );
  AOI21_X1 U12800 ( .B1(n13369), .B2(n13435), .A(n10149), .ZN(n10150) );
  INV_X1 U12801 ( .A(n13374), .ZN(n10156) );
  OAI22_X1 U12802 ( .A1(n10156), .A2(n13654), .B1(n15600), .B2(n10151), .ZN(
        n10152) );
  NAND2_X1 U12803 ( .A1(n10154), .A2(n10153), .ZN(P3_U3454) );
  INV_X1 U12804 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n10155) );
  NAND2_X1 U12805 ( .A1(n13374), .A2(n13617), .ZN(n10157) );
  NAND2_X1 U12806 ( .A1(n10158), .A2(n10157), .ZN(P3_U3486) );
  INV_X1 U12807 ( .A(n11730), .ZN(n10159) );
  NOR2_X1 U12808 ( .A1(n10160), .A2(n10159), .ZN(n10415) );
  NOR2_X2 U12809 ( .A1(n10161), .A2(n10383), .ZN(P1_U4016) );
  INV_X1 U12810 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10163) );
  AOI21_X1 U12811 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n10163), .A(n10162), .ZN(
        n10165) );
  INV_X1 U12812 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10164) );
  NOR2_X1 U12813 ( .A1(n10165), .A2(n10164), .ZN(n15617) );
  AOI21_X1 U12814 ( .B1(n10165), .B2(n10164), .A(n15617), .ZN(SUB_1596_U53) );
  NOR2_X1 U12815 ( .A1(n10039), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13702) );
  AND2_X1 U12816 ( .A1(n10171), .A2(P3_U3151), .ZN(n10762) );
  AOI222_X1 U12817 ( .A1(n10167), .A2(n13702), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10166), .C1(SI_3_), .C2(n10762), .ZN(n10168) );
  INV_X1 U12818 ( .A(n10168), .ZN(P3_U3292) );
  AOI222_X1 U12819 ( .A1(n10169), .A2(n13702), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n6489), .C1(SI_5_), .C2(n10762), .ZN(n10170) );
  INV_X1 U12820 ( .A(n10170), .ZN(P3_U3290) );
  NAND2_X1 U12821 ( .A1(n10171), .A2(P2_U3088), .ZN(n13019) );
  NOR2_X1 U12822 ( .A1(n10171), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14255) );
  INV_X2 U12823 ( .A(n14255), .ZN(n14247) );
  OAI222_X1 U12824 ( .A1(n15335), .A2(P2_U3088), .B1(n13019), .B2(n10195), 
        .C1(n10172), .C2(n14247), .ZN(P2_U3326) );
  INV_X2 U12825 ( .A(n10762), .ZN(n13719) );
  OAI222_X1 U12826 ( .A1(n13717), .A2(n10174), .B1(n13719), .B2(n10173), .C1(
        n10840), .C2(P3_U3151), .ZN(P3_U3288) );
  OAI222_X1 U12827 ( .A1(n10669), .A2(P3_U3151), .B1(n13717), .B2(n10178), 
        .C1(n10177), .C2(n13719), .ZN(P3_U3295) );
  OAI222_X1 U12828 ( .A1(n10822), .A2(P3_U3151), .B1(n13717), .B2(n10180), 
        .C1(n10179), .C2(n13719), .ZN(P3_U3289) );
  INV_X1 U12829 ( .A(n10181), .ZN(n10183) );
  OAI222_X1 U12830 ( .A1(n10580), .A2(P3_U3151), .B1(n13717), .B2(n10183), 
        .C1(n10182), .C2(n13719), .ZN(P3_U3293) );
  INV_X1 U12831 ( .A(n10184), .ZN(n10185) );
  OAI222_X1 U12832 ( .A1(n10186), .A2(P3_U3151), .B1(n13717), .B2(n10185), 
        .C1(n11991), .C2(n13719), .ZN(P3_U3291) );
  INV_X1 U12833 ( .A(n10187), .ZN(n10190) );
  INV_X1 U12834 ( .A(SI_8_), .ZN(n10189) );
  OAI222_X1 U12835 ( .A1(n13717), .A2(n10190), .B1(n13719), .B2(n10189), .C1(
        n10188), .C2(P3_U3151), .ZN(P3_U3287) );
  OAI222_X1 U12836 ( .A1(n13717), .A2(n10192), .B1(n13719), .B2(n10191), .C1(
        n11418), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U12837 ( .A(n14595), .ZN(n10196) );
  AND2_X1 U12838 ( .A1(n10193), .A2(P1_U3086), .ZN(n15161) );
  INV_X2 U12839 ( .A(n15161), .ZN(n15159) );
  OAI222_X1 U12840 ( .A1(n10196), .A2(P1_U3086), .B1(n15159), .B2(n10195), 
        .C1(n10194), .C2(n15165), .ZN(P1_U3354) );
  OAI222_X1 U12841 ( .A1(n15165), .A2(n7817), .B1(n15159), .B2(n10278), .C1(
        P1_U3086), .C2(n10436), .ZN(P1_U3353) );
  INV_X1 U12842 ( .A(n10197), .ZN(n10288) );
  OAI222_X1 U12843 ( .A1(n15165), .A2(n7867), .B1(n15159), .B2(n10288), .C1(
        P1_U3086), .C2(n14619), .ZN(P1_U3351) );
  NAND2_X1 U12844 ( .A1(n10223), .A2(n10198), .ZN(n10219) );
  INV_X1 U12845 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U12846 ( .A1(n10199), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10200) );
  AND2_X1 U12847 ( .A1(n10201), .A2(n10200), .ZN(n10218) );
  NAND2_X1 U12848 ( .A1(n10219), .A2(n10218), .ZN(n10217) );
  NAND2_X1 U12849 ( .A1(n10217), .A2(n10201), .ZN(n10202) );
  INV_X1 U12850 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U12851 ( .A1(n10205), .A2(n10204), .ZN(n10207) );
  INV_X1 U12852 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U12853 ( .A1(n10209), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10210) );
  INV_X1 U12854 ( .A(n10213), .ZN(n10212) );
  INV_X1 U12855 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U12856 ( .A1(n10212), .A2(n10211), .ZN(n10303) );
  NAND2_X1 U12857 ( .A1(n10213), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10214) );
  NAND2_X1 U12858 ( .A1(n10215), .A2(n10216), .ZN(n15614) );
  OAI21_X1 U12859 ( .B1(n10219), .B2(n10218), .A(n10217), .ZN(n10227) );
  NAND2_X1 U12860 ( .A1(n10221), .A2(n10220), .ZN(n10222) );
  NAND2_X1 U12861 ( .A1(n10223), .A2(n10222), .ZN(n10224) );
  NAND2_X1 U12862 ( .A1(n10224), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10226) );
  XOR2_X1 U12863 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10224), .Z(n15616) );
  NAND2_X1 U12864 ( .A1(n15617), .A2(n15616), .ZN(n10225) );
  NAND2_X1 U12865 ( .A1(n10226), .A2(n10225), .ZN(n10228) );
  NAND2_X1 U12866 ( .A1(n10227), .A2(n10228), .ZN(n15257) );
  INV_X1 U12867 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15259) );
  NAND2_X1 U12868 ( .A1(n15257), .A2(n15259), .ZN(n10231) );
  INV_X1 U12869 ( .A(n10227), .ZN(n10230) );
  INV_X1 U12870 ( .A(n10228), .ZN(n10229) );
  NAND2_X1 U12871 ( .A1(n10230), .A2(n10229), .ZN(n15258) );
  AND2_X1 U12872 ( .A1(n10231), .A2(n15258), .ZN(n15613) );
  OAI21_X1 U12873 ( .B1(n15614), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n15613), .ZN(
        n10233) );
  NAND2_X1 U12874 ( .A1(n15614), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n10232) );
  AND2_X1 U12875 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  NAND2_X1 U12876 ( .A1(n10235), .A2(n10234), .ZN(n10304) );
  OAI21_X1 U12877 ( .B1(n10235), .B2(n10234), .A(n10304), .ZN(SUB_1596_U59) );
  OAI222_X1 U12878 ( .A1(n13717), .A2(n10237), .B1(n13719), .B2(n10236), .C1(
        n11303), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12879 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10240) );
  INV_X1 U12880 ( .A(n10238), .ZN(n10280) );
  INV_X1 U12881 ( .A(n14635), .ZN(n10239) );
  OAI222_X1 U12882 ( .A1(n15165), .A2(n10240), .B1(n15159), .B2(n10280), .C1(
        P1_U3086), .C2(n10239), .ZN(P1_U3350) );
  INV_X1 U12883 ( .A(n10241), .ZN(n10282) );
  INV_X1 U12884 ( .A(n15165), .ZN(n15154) );
  AOI22_X1 U12885 ( .A1(n14680), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n15154), .ZN(n10242) );
  OAI21_X1 U12886 ( .B1(n10282), .B2(n15159), .A(n10242), .ZN(P1_U3346) );
  INV_X1 U12887 ( .A(n10243), .ZN(n10274) );
  INV_X1 U12888 ( .A(n14648), .ZN(n10244) );
  OAI222_X1 U12889 ( .A1(n15165), .A2(n10245), .B1(n15159), .B2(n10274), .C1(
        P1_U3086), .C2(n10244), .ZN(P1_U3349) );
  INV_X1 U12890 ( .A(n10246), .ZN(n10286) );
  AOI22_X1 U12891 ( .A1(n14664), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n15154), .ZN(n10247) );
  OAI21_X1 U12892 ( .B1(n10286), .B2(n15159), .A(n10247), .ZN(P1_U3348) );
  OAI222_X1 U12893 ( .A1(n13717), .A2(n10249), .B1(n13719), .B2(n10248), .C1(
        n13222), .C2(P3_U3151), .ZN(P3_U3284) );
  OAI222_X1 U12894 ( .A1(n15165), .A2(n10250), .B1(n15159), .B2(n10276), .C1(
        P1_U3086), .C2(n14606), .ZN(P1_U3352) );
  INV_X1 U12895 ( .A(n10251), .ZN(n10252) );
  INV_X1 U12896 ( .A(n10253), .ZN(n10254) );
  AOI22_X1 U12897 ( .A1(n15308), .A2(n10255), .B1(n10257), .B2(n10254), .ZN(
        P1_U3446) );
  INV_X1 U12898 ( .A(n10256), .ZN(n10258) );
  AOI22_X1 U12899 ( .A1(n15308), .A2(n10259), .B1(n10258), .B2(n10257), .ZN(
        P1_U3445) );
  INV_X1 U12900 ( .A(n10260), .ZN(n10389) );
  NAND2_X1 U12901 ( .A1(n10389), .A2(n11734), .ZN(n10338) );
  OR2_X1 U12902 ( .A1(n10262), .A2(n10261), .ZN(n10263) );
  AND2_X1 U12903 ( .A1(n7856), .A2(n10263), .ZN(n10337) );
  INV_X1 U12904 ( .A(n10337), .ZN(n10264) );
  AND2_X1 U12905 ( .A1(n10338), .A2(n10264), .ZN(n15269) );
  NOR2_X1 U12906 ( .A1(n15269), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12907 ( .A(n10265), .ZN(n10284) );
  AOI22_X1 U12908 ( .A1(n10605), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n15154), .ZN(n10266) );
  OAI21_X1 U12909 ( .B1(n10284), .B2(n15159), .A(n10266), .ZN(P1_U3347) );
  NAND2_X1 U12910 ( .A1(n10270), .A2(P3_D_REG_1__SCAN_IN), .ZN(n10267) );
  OAI21_X1 U12911 ( .B1(n10268), .B2(n10270), .A(n10267), .ZN(P3_U3377) );
  NAND2_X1 U12912 ( .A1(n10270), .A2(P3_D_REG_0__SCAN_IN), .ZN(n10269) );
  OAI21_X1 U12913 ( .B1(n10271), .B2(n10270), .A(n10269), .ZN(P3_U3376) );
  INV_X1 U12914 ( .A(n10272), .ZN(n10294) );
  AOI22_X1 U12915 ( .A1(n10649), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n15154), .ZN(n10273) );
  OAI21_X1 U12916 ( .B1(n10294), .B2(n15159), .A(n10273), .ZN(P1_U3345) );
  INV_X1 U12917 ( .A(n13019), .ZN(n11729) );
  INV_X1 U12918 ( .A(n11729), .ZN(n14257) );
  INV_X1 U12919 ( .A(n10676), .ZN(n10596) );
  OAI222_X1 U12920 ( .A1(n14247), .A2(n10275), .B1(n14257), .B2(n10274), .C1(
        P2_U3088), .C2(n10596), .ZN(P2_U3321) );
  OAI222_X1 U12921 ( .A1(n14247), .A2(n10277), .B1(n14257), .B2(n10276), .C1(
        P2_U3088), .C2(n15348), .ZN(P2_U3324) );
  OAI222_X1 U12922 ( .A1(n14247), .A2(n10279), .B1(n14257), .B2(n10278), .C1(
        P2_U3088), .C2(n10482), .ZN(P2_U3325) );
  INV_X1 U12923 ( .A(n10589), .ZN(n10508) );
  OAI222_X1 U12924 ( .A1(n14247), .A2(n10281), .B1(n14257), .B2(n10280), .C1(
        P2_U3088), .C2(n10508), .ZN(P2_U3322) );
  INV_X1 U12925 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10283) );
  INV_X1 U12926 ( .A(n11140), .ZN(n11134) );
  OAI222_X1 U12927 ( .A1(n14247), .A2(n10283), .B1(n14257), .B2(n10282), .C1(
        P2_U3088), .C2(n11134), .ZN(P2_U3318) );
  INV_X1 U12928 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10285) );
  OAI222_X1 U12929 ( .A1(n14247), .A2(n10285), .B1(n14257), .B2(n10284), .C1(
        P2_U3088), .C2(n10929), .ZN(P2_U3319) );
  INV_X1 U12930 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10287) );
  INV_X1 U12931 ( .A(n10680), .ZN(n15377) );
  OAI222_X1 U12932 ( .A1(n14247), .A2(n10287), .B1(n14257), .B2(n10286), .C1(
        P2_U3088), .C2(n15377), .ZN(P2_U3320) );
  OAI222_X1 U12933 ( .A1(n14247), .A2(n10289), .B1(n14257), .B2(n10288), .C1(
        P2_U3088), .C2(n15360), .ZN(P2_U3323) );
  OAI222_X1 U12934 ( .A1(n13717), .A2(n10292), .B1(n10291), .B2(P3_U3151), 
        .C1(n10290), .C2(n13719), .ZN(P3_U3283) );
  INV_X1 U12935 ( .A(n11268), .ZN(n11150) );
  INV_X1 U12936 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10293) );
  OAI222_X1 U12937 ( .A1(P2_U3088), .A2(n11150), .B1(n14257), .B2(n10294), 
        .C1(n10293), .C2(n14247), .ZN(P2_U3317) );
  INV_X1 U12938 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n10296) );
  NAND2_X1 U12939 ( .A1(n10298), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10959) );
  NAND2_X1 U12940 ( .A1(n10301), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10302) );
  INV_X1 U12941 ( .A(n10307), .ZN(n10305) );
  NAND2_X1 U12942 ( .A1(n10304), .A2(n10303), .ZN(n10306) );
  INV_X1 U12943 ( .A(n10306), .ZN(n10308) );
  INV_X1 U12944 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10309) );
  OAI21_X1 U12945 ( .B1(n6646), .B2(n10309), .A(n10958), .ZN(SUB_1596_U58) );
  AND2_X1 U12946 ( .A1(n10311), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12947 ( .A1(n10311), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12948 ( .A1(n10311), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12949 ( .A1(n10311), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12950 ( .A1(n10311), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12951 ( .A1(n10311), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12952 ( .A1(n10311), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12953 ( .A1(n10311), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12954 ( .A1(n10311), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12955 ( .A1(n10311), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12956 ( .A1(n10311), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12957 ( .A1(n10311), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12958 ( .A1(n10311), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12959 ( .A1(n10311), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12960 ( .A1(n10311), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12961 ( .A1(n10311), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12962 ( .A1(n10311), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12963 ( .A1(n10311), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12964 ( .A1(n10311), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12965 ( .A1(n10311), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12966 ( .A1(n10311), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12967 ( .A1(n10311), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12968 ( .A1(n10311), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12969 ( .A1(n10311), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12970 ( .A1(n10311), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12971 ( .A1(n10311), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12972 ( .A1(n10311), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12973 ( .A1(n10311), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  INV_X1 U12974 ( .A(n10311), .ZN(n10312) );
  INV_X1 U12975 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n11885) );
  NOR2_X1 U12976 ( .A1(n10312), .A2(n11885), .ZN(P3_U3250) );
  INV_X1 U12977 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n11886) );
  NOR2_X1 U12978 ( .A1(n10312), .A2(n11886), .ZN(P3_U3262) );
  INV_X1 U12979 ( .A(n10313), .ZN(n10315) );
  INV_X1 U12980 ( .A(n10720), .ZN(n10660) );
  OAI222_X1 U12981 ( .A1(n15165), .A2(n10314), .B1(n15159), .B2(n10315), .C1(
        P1_U3086), .C2(n10660), .ZN(P1_U3344) );
  INV_X1 U12982 ( .A(n11359), .ZN(n11352) );
  OAI222_X1 U12983 ( .A1(n14247), .A2(n10316), .B1(n14257), .B2(n10315), .C1(
        P2_U3088), .C2(n11352), .ZN(P2_U3316) );
  INV_X1 U12984 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10317) );
  MUX2_X1 U12985 ( .A(n10317), .B(P1_REG1_REG_8__SCAN_IN), .S(n10605), .Z(
        n10336) );
  INV_X1 U12986 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10318) );
  MUX2_X1 U12987 ( .A(n10318), .B(P1_REG1_REG_4__SCAN_IN), .S(n14619), .Z(
        n10326) );
  INV_X1 U12988 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10319) );
  MUX2_X1 U12989 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10319), .S(n14595), .Z(
        n14593) );
  AND2_X1 U12990 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14594) );
  NAND2_X1 U12991 ( .A1(n14593), .A2(n14594), .ZN(n14592) );
  NAND2_X1 U12992 ( .A1(n14595), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U12993 ( .A1(n14592), .A2(n10320), .ZN(n10439) );
  XNOR2_X1 U12994 ( .A(n10436), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10440) );
  NAND2_X1 U12995 ( .A1(n10439), .A2(n10440), .ZN(n10323) );
  INV_X1 U12996 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10321) );
  OR2_X1 U12997 ( .A1(n10436), .A2(n10321), .ZN(n10322) );
  NAND2_X1 U12998 ( .A1(n10323), .A2(n10322), .ZN(n14600) );
  INV_X1 U12999 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10324) );
  MUX2_X1 U13000 ( .A(n10324), .B(P1_REG1_REG_3__SCAN_IN), .S(n14606), .Z(
        n14601) );
  NAND2_X1 U13001 ( .A1(n14600), .A2(n14601), .ZN(n14621) );
  OR2_X1 U13002 ( .A1(n14606), .A2(n10324), .ZN(n14620) );
  NAND2_X1 U13003 ( .A1(n14621), .A2(n14620), .ZN(n10325) );
  NAND2_X1 U13004 ( .A1(n10326), .A2(n10325), .ZN(n14624) );
  INV_X1 U13005 ( .A(n14619), .ZN(n10350) );
  NAND2_X1 U13006 ( .A1(n10350), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10327) );
  MUX2_X1 U13007 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7872), .S(n14635), .Z(
        n14633) );
  NAND2_X1 U13008 ( .A1(n14632), .A2(n14633), .ZN(n14631) );
  OR2_X1 U13009 ( .A1(n14635), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10328) );
  AND2_X1 U13010 ( .A1(n14631), .A2(n10328), .ZN(n14647) );
  INV_X1 U13011 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10329) );
  MUX2_X1 U13012 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10329), .S(n14648), .Z(
        n14646) );
  NAND2_X1 U13013 ( .A1(n14648), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n14660) );
  NAND2_X1 U13014 ( .A1(n14661), .A2(n14660), .ZN(n10332) );
  INV_X1 U13015 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10330) );
  MUX2_X1 U13016 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10330), .S(n14664), .Z(
        n10331) );
  NAND2_X1 U13017 ( .A1(n10332), .A2(n10331), .ZN(n14663) );
  NAND2_X1 U13018 ( .A1(n14664), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10333) );
  NAND2_X1 U13019 ( .A1(n14663), .A2(n10333), .ZN(n10335) );
  INV_X1 U13020 ( .A(n10607), .ZN(n10334) );
  AOI21_X1 U13021 ( .B1(n10336), .B2(n10335), .A(n10334), .ZN(n10366) );
  NAND2_X1 U13022 ( .A1(n10338), .A2(n10337), .ZN(n15272) );
  INV_X1 U13023 ( .A(n15269), .ZN(n14745) );
  INV_X1 U13024 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U13025 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11668) );
  OAI21_X1 U13026 ( .B1(n14745), .B2(n10982), .A(n11668), .ZN(n10340) );
  AOI21_X1 U13027 ( .B1(n10605), .B2(n14737), .A(n10340), .ZN(n10365) );
  OR2_X1 U13028 ( .A1(n7809), .A2(n10433), .ZN(n10341) );
  INV_X1 U13029 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10900) );
  MUX2_X1 U13030 ( .A(n10900), .B(P1_REG2_REG_4__SCAN_IN), .S(n14619), .Z(
        n10349) );
  INV_X1 U13031 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10342) );
  MUX2_X1 U13032 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10342), .S(n14595), .Z(
        n14590) );
  AND2_X1 U13033 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10343) );
  NAND2_X1 U13034 ( .A1(n14590), .A2(n10343), .ZN(n14589) );
  NAND2_X1 U13035 ( .A1(n14595), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U13036 ( .A1(n14589), .A2(n10344), .ZN(n10441) );
  INV_X1 U13037 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10345) );
  MUX2_X1 U13038 ( .A(n10345), .B(P1_REG2_REG_2__SCAN_IN), .S(n10436), .Z(
        n10442) );
  NAND2_X1 U13039 ( .A1(n10441), .A2(n10442), .ZN(n14603) );
  OR2_X1 U13040 ( .A1(n10436), .A2(n10345), .ZN(n14602) );
  NAND2_X1 U13041 ( .A1(n14603), .A2(n14602), .ZN(n10347) );
  INV_X1 U13042 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11031) );
  MUX2_X1 U13043 ( .A(n11031), .B(P1_REG2_REG_3__SCAN_IN), .S(n14606), .Z(
        n10346) );
  NAND2_X1 U13044 ( .A1(n10347), .A2(n10346), .ZN(n14616) );
  OR2_X1 U13045 ( .A1(n14606), .A2(n11031), .ZN(n14615) );
  NAND2_X1 U13046 ( .A1(n14616), .A2(n14615), .ZN(n10348) );
  NAND2_X1 U13047 ( .A1(n10349), .A2(n10348), .ZN(n14638) );
  NAND2_X1 U13048 ( .A1(n10350), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14637) );
  NAND2_X1 U13049 ( .A1(n14638), .A2(n14637), .ZN(n10353) );
  MUX2_X1 U13050 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10351), .S(n14635), .Z(
        n10352) );
  NAND2_X1 U13051 ( .A1(n10353), .A2(n10352), .ZN(n14651) );
  NAND2_X1 U13052 ( .A1(n14635), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14650) );
  NAND2_X1 U13053 ( .A1(n14651), .A2(n14650), .ZN(n10355) );
  INV_X1 U13054 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11426) );
  MUX2_X1 U13055 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11426), .S(n14648), .Z(
        n10354) );
  NAND2_X1 U13056 ( .A1(n10355), .A2(n10354), .ZN(n14667) );
  NAND2_X1 U13057 ( .A1(n14648), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14666) );
  NAND2_X1 U13058 ( .A1(n14667), .A2(n14666), .ZN(n10357) );
  INV_X1 U13059 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11592) );
  MUX2_X1 U13060 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11592), .S(n14664), .Z(
        n10356) );
  NAND2_X1 U13061 ( .A1(n10357), .A2(n10356), .ZN(n14669) );
  NAND2_X1 U13062 ( .A1(n14664), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10362) );
  NAND2_X1 U13063 ( .A1(n14669), .A2(n10362), .ZN(n10360) );
  INV_X1 U13064 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10358) );
  MUX2_X1 U13065 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10358), .S(n10605), .Z(
        n10359) );
  NAND2_X1 U13066 ( .A1(n10360), .A2(n10359), .ZN(n14683) );
  MUX2_X1 U13067 ( .A(n10358), .B(P1_REG2_REG_8__SCAN_IN), .S(n10605), .Z(
        n10361) );
  NAND3_X1 U13068 ( .A1(n14669), .A2(n10362), .A3(n10361), .ZN(n10363) );
  NAND3_X1 U13069 ( .A1(n14733), .A2(n14683), .A3(n10363), .ZN(n10364) );
  OAI211_X1 U13070 ( .C1(n10366), .C2(n11646), .A(n10365), .B(n10364), .ZN(
        P1_U3251) );
  INV_X1 U13071 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n11981) );
  NAND2_X1 U13072 ( .A1(P3_U3897), .A2(n12448), .ZN(n10367) );
  OAI21_X1 U13073 ( .B1(P3_U3897), .B2(n11981), .A(n10367), .ZN(P3_U3502) );
  AND2_X1 U13074 ( .A1(n15314), .A2(n14988), .ZN(n10368) );
  NOR2_X1 U13075 ( .A1(n10369), .A2(n10368), .ZN(n15302) );
  INV_X1 U13076 ( .A(n10474), .ZN(n10370) );
  NOR2_X1 U13077 ( .A1(n10370), .A2(n14993), .ZN(n15298) );
  INV_X1 U13078 ( .A(n10371), .ZN(n10372) );
  NOR2_X1 U13079 ( .A1(n10511), .A2(n10372), .ZN(n15300) );
  NOR3_X1 U13080 ( .A1(n15302), .A2(n15298), .A3(n15300), .ZN(n10410) );
  NAND2_X1 U13081 ( .A1(n15320), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10373) );
  OAI21_X1 U13082 ( .B1(n10410), .B2(n15320), .A(n10373), .ZN(P1_U3528) );
  INV_X1 U13083 ( .A(n10374), .ZN(n10377) );
  NAND3_X1 U13084 ( .A1(n10377), .A2(n10376), .A3(n10375), .ZN(n10395) );
  OR2_X1 U13085 ( .A1(n10395), .A2(n10378), .ZN(n14420) );
  NAND2_X1 U13086 ( .A1(n14547), .A2(n15008), .ZN(n14555) );
  OAI22_X1 U13087 ( .A1(n10511), .A2(n10527), .B1(n15264), .B2(n10383), .ZN(
        n10381) );
  INV_X1 U13088 ( .A(n10381), .ZN(n10382) );
  INV_X2 U13089 ( .A(n10527), .ZN(n14351) );
  NAND2_X1 U13090 ( .A1(n14587), .A2(n14351), .ZN(n10387) );
  INV_X1 U13091 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10384) );
  OAI22_X1 U13092 ( .A1(n10511), .A2(n14414), .B1(n10384), .B2(n10383), .ZN(
        n10385) );
  INV_X1 U13093 ( .A(n10385), .ZN(n10386) );
  NAND2_X1 U13094 ( .A1(n10387), .A2(n10386), .ZN(n10471) );
  OAI21_X1 U13095 ( .B1(n10388), .B2(n10471), .A(n10473), .ZN(n10432) );
  OR2_X1 U13096 ( .A1(n15311), .A2(n10390), .ZN(n10391) );
  AOI22_X1 U13097 ( .A1(n14534), .A2(n10474), .B1(n10432), .B2(n14540), .ZN(
        n10401) );
  NAND2_X1 U13098 ( .A1(n10395), .A2(n10394), .ZN(n10398) );
  INV_X1 U13099 ( .A(n10396), .ZN(n10397) );
  NAND2_X1 U13100 ( .A1(n10398), .A2(n10397), .ZN(n10809) );
  OR2_X1 U13101 ( .A1(n10809), .A2(P1_U3086), .ZN(n10541) );
  AOI22_X1 U13102 ( .A1(n10393), .A2(n10399), .B1(n10541), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10400) );
  NAND2_X1 U13103 ( .A1(n10401), .A2(n10400), .ZN(P1_U3232) );
  OAI222_X1 U13104 ( .A1(n13717), .A2(n10404), .B1(n10403), .B2(P3_U3151), 
        .C1(n10402), .C2(n13719), .ZN(P3_U3282) );
  INV_X1 U13105 ( .A(n12322), .ZN(n10407) );
  INV_X1 U13106 ( .A(n10405), .ZN(n10409) );
  OAI222_X1 U13107 ( .A1(P2_U3088), .A2(n10407), .B1(n14257), .B2(n10409), 
        .C1(n10406), .C2(n14247), .ZN(P2_U3315) );
  INV_X1 U13108 ( .A(n11006), .ZN(n10726) );
  OAI222_X1 U13109 ( .A1(P1_U3086), .A2(n10726), .B1(n15159), .B2(n10409), 
        .C1(n10408), .C2(n15165), .ZN(P1_U3343) );
  INV_X1 U13110 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n11922) );
  OR2_X1 U13111 ( .A1(n10410), .A2(n15317), .ZN(n10411) );
  OAI21_X1 U13112 ( .B1(n15319), .B2(n11922), .A(n10411), .ZN(P1_U3459) );
  AOI21_X1 U13113 ( .B1(n10413), .B2(n11730), .A(n10412), .ZN(n10414) );
  OR2_X1 U13114 ( .A1(n10415), .A2(n10414), .ZN(n10428) );
  NOR2_X1 U13115 ( .A1(n10420), .A2(P2_U3088), .ZN(n14254) );
  NAND2_X1 U13116 ( .A1(n10428), .A2(n14254), .ZN(n10422) );
  INV_X1 U13117 ( .A(n10422), .ZN(n10418) );
  INV_X1 U13118 ( .A(n10417), .ZN(n12903) );
  INV_X1 U13119 ( .A(n15423), .ZN(n12329) );
  XNOR2_X1 U13120 ( .A(n15335), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n15339) );
  AND2_X1 U13121 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15338) );
  NAND2_X1 U13122 ( .A1(n15339), .A2(n15338), .ZN(n15337) );
  INV_X1 U13123 ( .A(n15335), .ZN(n10424) );
  NAND2_X1 U13124 ( .A1(n10424), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10419) );
  NAND2_X1 U13125 ( .A1(n15337), .A2(n10419), .ZN(n10493) );
  XNOR2_X1 U13126 ( .A(n10482), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n10492) );
  XNOR2_X1 U13127 ( .A(n10493), .B(n10492), .ZN(n10421) );
  NAND2_X1 U13128 ( .A1(n10428), .A2(n10420), .ZN(n15361) );
  OAI22_X1 U13129 ( .A1(n12329), .A2(n10421), .B1(n10482), .B2(n15408), .ZN(
        n10431) );
  NAND2_X1 U13130 ( .A1(n10424), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10425) );
  AND3_X1 U13131 ( .A1(n10426), .A2(n15340), .A3(n10425), .ZN(n10427) );
  NOR3_X1 U13132 ( .A1(n15392), .A2(n10483), .A3(n10427), .ZN(n10430) );
  OAI22_X1 U13133 ( .A1(n15427), .A2(n15259), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11394), .ZN(n10429) );
  OR3_X1 U13134 ( .A1(n10431), .A2(n10430), .A3(n10429), .ZN(P2_U3216) );
  NAND2_X1 U13135 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14588) );
  MUX2_X1 U13136 ( .A(n14588), .B(n10432), .S(n10433), .Z(n10435) );
  NOR2_X1 U13137 ( .A1(n10433), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10434) );
  OR2_X1 U13138 ( .A1(n7809), .A2(n10434), .ZN(n15262) );
  NAND2_X1 U13139 ( .A1(n15262), .A2(n15264), .ZN(n15267) );
  OAI211_X1 U13140 ( .C1(n10435), .C2(n7809), .A(n14580), .B(n15267), .ZN(
        n14628) );
  INV_X1 U13141 ( .A(n10436), .ZN(n10447) );
  INV_X1 U13142 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10437) );
  OAI22_X1 U13143 ( .A1(n14745), .A2(n10438), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10437), .ZN(n10446) );
  XNOR2_X1 U13144 ( .A(n10439), .B(n10440), .ZN(n10444) );
  OAI211_X1 U13145 ( .C1(n10442), .C2(n10441), .A(n14733), .B(n14603), .ZN(
        n10443) );
  OAI21_X1 U13146 ( .B1(n10444), .B2(n11646), .A(n10443), .ZN(n10445) );
  AOI211_X1 U13147 ( .C1(n10447), .C2(n14737), .A(n10446), .B(n10445), .ZN(
        n10448) );
  NAND2_X1 U13148 ( .A1(n14628), .A2(n10448), .ZN(P1_U3245) );
  OAI21_X1 U13149 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n10449), .A(n10774), .ZN(
        n10455) );
  XNOR2_X1 U13150 ( .A(n10451), .B(n10450), .ZN(n10453) );
  AOI22_X1 U13151 ( .A1(n15503), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n10452) );
  OAI21_X1 U13152 ( .B1(n10453), .B2(n13333), .A(n10452), .ZN(n10454) );
  AOI21_X1 U13153 ( .B1(n13348), .B2(n10455), .A(n10454), .ZN(n10461) );
  AND3_X1 U13154 ( .A1(n10570), .A2(n10457), .A3(n10456), .ZN(n10458) );
  OAI21_X1 U13155 ( .B1(n10459), .B2(n10458), .A(n13270), .ZN(n10460) );
  OAI211_X1 U13156 ( .C1(n13355), .C2(n10462), .A(n10461), .B(n10460), .ZN(
        P3_U3185) );
  INV_X1 U13157 ( .A(n15397), .ZN(n10464) );
  INV_X1 U13158 ( .A(n10463), .ZN(n10465) );
  OAI222_X1 U13159 ( .A1(P2_U3088), .A2(n10464), .B1(n13019), .B2(n10465), 
        .C1(n7541), .C2(n14247), .ZN(P2_U3314) );
  INV_X1 U13160 ( .A(n11520), .ZN(n11014) );
  OAI222_X1 U13161 ( .A1(n15165), .A2(n10466), .B1(n15159), .B2(n10465), .C1(
        n11014), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U13162 ( .A(n10467), .ZN(n10470) );
  OAI222_X1 U13163 ( .A1(n13717), .A2(n10470), .B1(n13719), .B2(n10469), .C1(
        n10468), .C2(P3_U3151), .ZN(P3_U3281) );
  NAND2_X1 U13164 ( .A1(n10473), .A2(n10472), .ZN(n10533) );
  NAND2_X1 U13165 ( .A1(n10474), .A2(n14351), .ZN(n10476) );
  NOR2_X1 U13166 ( .A1(n15292), .A2(n10527), .ZN(n10477) );
  XNOR2_X1 U13167 ( .A(n10535), .B(n10536), .ZN(n10534) );
  XOR2_X1 U13168 ( .A(n10533), .B(n10478), .Z(n10481) );
  NOR2_X1 U13169 ( .A1(n14420), .A2(n15032), .ZN(n14377) );
  AOI22_X1 U13170 ( .A1(n14534), .A2(n14585), .B1(n14377), .B2(n14587), .ZN(
        n10480) );
  AOI22_X1 U13171 ( .A1(n10393), .A2(n10521), .B1(n10541), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10479) );
  OAI211_X1 U13172 ( .C1(n10481), .C2(n14561), .A(n10480), .B(n10479), .ZN(
        P1_U3222) );
  INV_X1 U13173 ( .A(n15427), .ZN(n15373) );
  NAND2_X1 U13174 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n12925) );
  INV_X1 U13175 ( .A(n12925), .ZN(n10490) );
  INV_X1 U13176 ( .A(n10482), .ZN(n10494) );
  AOI21_X1 U13177 ( .B1(n10494), .B2(P2_REG1_REG_2__SCAN_IN), .A(n10483), .ZN(
        n15354) );
  MUX2_X1 U13178 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10484), .S(n15348), .Z(
        n15353) );
  OR2_X1 U13179 ( .A1(n15354), .A2(n15353), .ZN(n15356) );
  OAI21_X1 U13180 ( .B1(n15348), .B2(n10484), .A(n15356), .ZN(n15364) );
  MUX2_X1 U13181 ( .A(n10485), .B(P2_REG1_REG_4__SCAN_IN), .S(n15360), .Z(
        n15365) );
  NAND2_X1 U13182 ( .A1(n10499), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10487) );
  MUX2_X1 U13183 ( .A(n8512), .B(P2_REG1_REG_5__SCAN_IN), .S(n10589), .Z(
        n10486) );
  AND3_X1 U13184 ( .A1(n15363), .A2(n10487), .A3(n10486), .ZN(n10488) );
  NOR3_X1 U13185 ( .A1(n15392), .A2(n10588), .A3(n10488), .ZN(n10489) );
  AOI211_X1 U13186 ( .C1(n15373), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10490), .B(
        n10489), .ZN(n10507) );
  MUX2_X1 U13187 ( .A(n10491), .B(P2_REG2_REG_4__SCAN_IN), .S(n15360), .Z(
        n15368) );
  NAND2_X1 U13188 ( .A1(n10493), .A2(n10492), .ZN(n10496) );
  NAND2_X1 U13189 ( .A1(n10494), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10495) );
  NAND2_X1 U13190 ( .A1(n10496), .A2(n10495), .ZN(n15351) );
  INV_X1 U13191 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10497) );
  MUX2_X1 U13192 ( .A(n10497), .B(P2_REG2_REG_3__SCAN_IN), .S(n15348), .Z(
        n15352) );
  NAND2_X1 U13193 ( .A1(n15351), .A2(n15352), .ZN(n15350) );
  OR2_X1 U13194 ( .A1(n15348), .A2(n10497), .ZN(n10498) );
  NAND2_X1 U13195 ( .A1(n15350), .A2(n10498), .ZN(n15367) );
  NAND2_X1 U13196 ( .A1(n15368), .A2(n15367), .ZN(n15366) );
  NAND2_X1 U13197 ( .A1(n10499), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10504) );
  NAND2_X1 U13198 ( .A1(n15366), .A2(n10504), .ZN(n10502) );
  MUX2_X1 U13199 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10500), .S(n10589), .Z(
        n10501) );
  MUX2_X1 U13200 ( .A(n10500), .B(P2_REG2_REG_5__SCAN_IN), .S(n10589), .Z(
        n10503) );
  NAND3_X1 U13201 ( .A1(n15366), .A2(n10504), .A3(n10503), .ZN(n10505) );
  NAND3_X1 U13202 ( .A1(n15423), .A2(n10586), .A3(n10505), .ZN(n10506) );
  OAI211_X1 U13203 ( .C1(n15408), .C2(n10508), .A(n10507), .B(n10506), .ZN(
        P2_U3219) );
  INV_X1 U13204 ( .A(n10517), .ZN(n10510) );
  OAI21_X1 U13205 ( .B1(n10510), .B2(n10509), .A(n14874), .ZN(n10515) );
  NOR2_X1 U13206 ( .A1(n10511), .A2(n15292), .ZN(n10512) );
  OR2_X1 U13207 ( .A1(n10556), .A2(n10512), .ZN(n10520) );
  XNOR2_X1 U13208 ( .A(n10520), .B(n10474), .ZN(n10513) );
  AOI21_X1 U13209 ( .B1(n10513), .B2(n14874), .A(n14587), .ZN(n10514) );
  AOI21_X1 U13210 ( .B1(n10515), .B2(n15032), .A(n10514), .ZN(n15286) );
  XNOR2_X1 U13211 ( .A(n10517), .B(n10516), .ZN(n10519) );
  INV_X1 U13212 ( .A(n14585), .ZN(n10518) );
  OAI22_X1 U13213 ( .A1(n10519), .A2(n15314), .B1(n10518), .B2(n14993), .ZN(
        n15287) );
  NOR2_X1 U13214 ( .A1(n10520), .A2(n15015), .ZN(n15288) );
  NOR3_X1 U13215 ( .A1(n15286), .A2(n15287), .A3(n15288), .ZN(n10526) );
  AOI22_X1 U13216 ( .A1(n11749), .A2(n10521), .B1(n15320), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n10522) );
  OAI21_X1 U13217 ( .B1(n10526), .B2(n15320), .A(n10522), .ZN(P1_U3529) );
  INV_X1 U13218 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10523) );
  OAI22_X1 U13219 ( .A1(n15143), .A2(n15292), .B1(n15319), .B2(n10523), .ZN(
        n10524) );
  INV_X1 U13220 ( .A(n10524), .ZN(n10525) );
  OAI21_X1 U13221 ( .B1(n10526), .B2(n15317), .A(n10525), .ZN(P1_U3462) );
  NAND2_X1 U13222 ( .A1(n14585), .A2(n10794), .ZN(n10529) );
  NAND2_X1 U13223 ( .A1(n10530), .A2(n14351), .ZN(n10528) );
  NAND2_X1 U13224 ( .A1(n10530), .A2(n14346), .ZN(n10532) );
  NAND2_X1 U13225 ( .A1(n14585), .A2(n14351), .ZN(n10531) );
  NAND2_X1 U13226 ( .A1(n10534), .A2(n10533), .ZN(n10539) );
  INV_X1 U13227 ( .A(n10535), .ZN(n10537) );
  NAND2_X1 U13228 ( .A1(n10537), .A2(n10536), .ZN(n10538) );
  AOI22_X1 U13229 ( .A1(n14534), .A2(n14584), .B1(n14377), .B2(n10474), .ZN(
        n10543) );
  AOI22_X1 U13230 ( .A1(n10393), .A2(n10530), .B1(n10541), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10542) );
  OAI211_X1 U13231 ( .C1(n10544), .C2(n14561), .A(n10543), .B(n10542), .ZN(
        P1_U3237) );
  XNOR2_X1 U13232 ( .A(n10545), .B(n10546), .ZN(n10547) );
  NAND2_X1 U13233 ( .A1(n10547), .A2(n15078), .ZN(n10555) );
  XNOR2_X1 U13234 ( .A(n10549), .B(n10548), .ZN(n10553) );
  NAND2_X1 U13235 ( .A1(n10474), .A2(n15010), .ZN(n10551) );
  NAND2_X1 U13236 ( .A1(n14584), .A2(n15008), .ZN(n10550) );
  NAND2_X1 U13237 ( .A1(n10551), .A2(n10550), .ZN(n10552) );
  AOI21_X1 U13238 ( .B1(n10553), .B2(n14874), .A(n10552), .ZN(n10554) );
  NAND2_X1 U13239 ( .A1(n10555), .A2(n10554), .ZN(n12938) );
  OR2_X1 U13240 ( .A1(n12943), .A2(n10556), .ZN(n10557) );
  AND3_X1 U13241 ( .A1(n10713), .A2(n10557), .A3(n6432), .ZN(n12940) );
  NOR2_X1 U13242 ( .A1(n12938), .A2(n12940), .ZN(n10562) );
  INV_X1 U13243 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10558) );
  OAI22_X1 U13244 ( .A1(n15143), .A2(n12943), .B1(n15319), .B2(n10558), .ZN(
        n10559) );
  INV_X1 U13245 ( .A(n10559), .ZN(n10560) );
  OAI21_X1 U13246 ( .B1(n10562), .B2(n15317), .A(n10560), .ZN(P1_U3465) );
  AOI22_X1 U13247 ( .A1(n11749), .A2(n10530), .B1(P1_REG1_REG_2__SCAN_IN), 
        .B2(n15320), .ZN(n10561) );
  OAI21_X1 U13248 ( .B1(n10562), .B2(n15320), .A(n10561), .ZN(P1_U3530) );
  OAI21_X1 U13249 ( .B1(n10565), .B2(n10564), .A(n10563), .ZN(n10578) );
  AOI21_X1 U13250 ( .B1(n10568), .B2(n10567), .A(n10566), .ZN(n10569) );
  NOR2_X1 U13251 ( .A1(n13333), .A2(n10569), .ZN(n10577) );
  AOI22_X1 U13252 ( .A1(n15503), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10575) );
  NOR3_X1 U13253 ( .A1(n10620), .A2(n10572), .A3(n10571), .ZN(n10573) );
  OAI21_X1 U13254 ( .B1(n7223), .B2(n10573), .A(n13270), .ZN(n10574) );
  NAND2_X1 U13255 ( .A1(n10575), .A2(n10574), .ZN(n10576) );
  AOI211_X1 U13256 ( .C1(n13348), .C2(n10578), .A(n10577), .B(n10576), .ZN(
        n10579) );
  OAI21_X1 U13257 ( .B1(n10580), .B2(n13355), .A(n10579), .ZN(P3_U3184) );
  NAND2_X1 U13258 ( .A1(n10589), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13259 ( .A1(n10586), .A2(n10585), .ZN(n10583) );
  INV_X1 U13260 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10581) );
  MUX2_X1 U13261 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10581), .S(n10676), .Z(
        n10582) );
  NAND2_X1 U13262 ( .A1(n10583), .A2(n10582), .ZN(n10678) );
  MUX2_X1 U13263 ( .A(n10581), .B(P2_REG2_REG_6__SCAN_IN), .S(n10676), .Z(
        n10584) );
  NAND3_X1 U13264 ( .A1(n10586), .A2(n10585), .A3(n10584), .ZN(n10587) );
  NAND3_X1 U13265 ( .A1(n15423), .A2(n10678), .A3(n10587), .ZN(n10595) );
  NAND2_X1 U13266 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n11551) );
  MUX2_X1 U13267 ( .A(n8540), .B(P2_REG1_REG_6__SCAN_IN), .S(n10676), .Z(
        n10590) );
  AOI211_X1 U13268 ( .C1(n10590), .C2(n6639), .A(n10674), .B(n15392), .ZN(
        n10591) );
  INV_X1 U13269 ( .A(n10591), .ZN(n10592) );
  NAND2_X1 U13270 ( .A1(n11551), .A2(n10592), .ZN(n10593) );
  AOI21_X1 U13271 ( .B1(n15373), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10593), .ZN(
        n10594) );
  OAI211_X1 U13272 ( .C1(n15408), .C2(n10596), .A(n10595), .B(n10594), .ZN(
        P2_U3220) );
  INV_X1 U13273 ( .A(n10649), .ZN(n10616) );
  NAND2_X1 U13274 ( .A1(n10605), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n14682) );
  NAND2_X1 U13275 ( .A1(n14683), .A2(n14682), .ZN(n10598) );
  INV_X1 U13276 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11771) );
  MUX2_X1 U13277 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n11771), .S(n14680), .Z(
        n10597) );
  NAND2_X1 U13278 ( .A1(n10598), .A2(n10597), .ZN(n14685) );
  NAND2_X1 U13279 ( .A1(n14680), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10603) );
  NAND2_X1 U13280 ( .A1(n14685), .A2(n10603), .ZN(n10601) );
  INV_X1 U13281 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10599) );
  MUX2_X1 U13282 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10599), .S(n10649), .Z(
        n10600) );
  NAND2_X1 U13283 ( .A1(n10601), .A2(n10600), .ZN(n10655) );
  MUX2_X1 U13284 ( .A(n10599), .B(P1_REG2_REG_10__SCAN_IN), .S(n10649), .Z(
        n10602) );
  NAND3_X1 U13285 ( .A1(n14685), .A2(n10603), .A3(n10602), .ZN(n10604) );
  NAND3_X1 U13286 ( .A1(n10655), .A2(n14733), .A3(n10604), .ZN(n10615) );
  NAND2_X1 U13287 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12166)
         );
  INV_X1 U13288 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n12109) );
  XNOR2_X1 U13289 ( .A(n10649), .B(n12109), .ZN(n10611) );
  OR2_X1 U13290 ( .A1(n10605), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10606) );
  INV_X1 U13291 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10608) );
  XNOR2_X1 U13292 ( .A(n14680), .B(n10608), .ZN(n14675) );
  NAND2_X1 U13293 ( .A1(n14674), .A2(n14675), .ZN(n14673) );
  OR2_X1 U13294 ( .A1(n14680), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10609) );
  AND2_X1 U13295 ( .A1(n14673), .A2(n10609), .ZN(n10610) );
  OAI211_X1 U13296 ( .C1(n10611), .C2(n10610), .A(n14739), .B(n10647), .ZN(
        n10612) );
  NAND2_X1 U13297 ( .A1(n12166), .A2(n10612), .ZN(n10613) );
  AOI21_X1 U13298 ( .B1(n15269), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10613), 
        .ZN(n10614) );
  OAI211_X1 U13299 ( .C1(n14719), .C2(n10616), .A(n10615), .B(n10614), .ZN(
        P1_U3253) );
  NAND2_X1 U13300 ( .A1(n10617), .A2(n15558), .ZN(n10618) );
  NAND2_X1 U13301 ( .A1(n10619), .A2(n10618), .ZN(n10632) );
  NAND2_X1 U13302 ( .A1(n15503), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10626) );
  INV_X1 U13303 ( .A(n10620), .ZN(n10623) );
  NAND2_X1 U13304 ( .A1(n10621), .A2(n10663), .ZN(n10622) );
  NAND2_X1 U13305 ( .A1(n10623), .A2(n10622), .ZN(n10624) );
  NAND2_X1 U13306 ( .A1(n13270), .A2(n10624), .ZN(n10625) );
  OAI211_X1 U13307 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n15554), .A(n10626), .B(
        n10625), .ZN(n10631) );
  XNOR2_X1 U13308 ( .A(n10628), .B(n10627), .ZN(n10629) );
  NOR2_X1 U13309 ( .A1(n13333), .A2(n10629), .ZN(n10630) );
  AOI211_X1 U13310 ( .C1(n13348), .C2(n10632), .A(n10631), .B(n10630), .ZN(
        n10633) );
  OAI21_X1 U13311 ( .B1(n10634), .B2(n13355), .A(n10633), .ZN(P3_U3183) );
  INV_X1 U13312 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10635) );
  OAI22_X1 U13313 ( .A1(n12329), .A2(n10636), .B1(n10635), .B2(n15392), .ZN(
        n10639) );
  NAND2_X1 U13314 ( .A1(n15423), .A2(n10636), .ZN(n10637) );
  OAI211_X1 U13315 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15392), .A(n10637), .B(
        n15408), .ZN(n10638) );
  MUX2_X1 U13316 ( .A(n10639), .B(n10638), .S(P2_IR_REG_0__SCAN_IN), .Z(n10641) );
  OAI22_X1 U13317 ( .A1(n15427), .A2(n10164), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11067), .ZN(n10640) );
  OR2_X1 U13318 ( .A1(n10641), .A2(n10640), .ZN(P2_U3214) );
  INV_X1 U13319 ( .A(n10647), .ZN(n10643) );
  AND2_X1 U13320 ( .A1(n10649), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10644) );
  OR2_X1 U13321 ( .A1(n10720), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10728) );
  NAND2_X1 U13322 ( .A1(n10720), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13323 ( .A1(n10728), .A2(n10642), .ZN(n10645) );
  OAI21_X1 U13324 ( .B1(n10643), .B2(n10644), .A(n10645), .ZN(n10648) );
  NOR2_X1 U13325 ( .A1(n10645), .A2(n10644), .ZN(n10646) );
  NAND2_X1 U13326 ( .A1(n10647), .A2(n10646), .ZN(n10729) );
  AOI21_X1 U13327 ( .B1(n10648), .B2(n10729), .A(n11646), .ZN(n10662) );
  NAND2_X1 U13328 ( .A1(n10649), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10654) );
  NAND2_X1 U13329 ( .A1(n10655), .A2(n10654), .ZN(n10652) );
  INV_X1 U13330 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10650) );
  MUX2_X1 U13331 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10650), .S(n10720), .Z(
        n10651) );
  NAND2_X1 U13332 ( .A1(n10652), .A2(n10651), .ZN(n10722) );
  MUX2_X1 U13333 ( .A(n10650), .B(P1_REG2_REG_11__SCAN_IN), .S(n10720), .Z(
        n10653) );
  NAND3_X1 U13334 ( .A1(n10655), .A2(n10654), .A3(n10653), .ZN(n10656) );
  NAND3_X1 U13335 ( .A1(n10722), .A2(n14733), .A3(n10656), .ZN(n10659) );
  NOR2_X1 U13336 ( .A1(n10657), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14523) );
  AOI21_X1 U13337 ( .B1(n15269), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n14523), 
        .ZN(n10658) );
  OAI211_X1 U13338 ( .C1(n14719), .C2(n10660), .A(n10659), .B(n10658), .ZN(
        n10661) );
  OR2_X1 U13339 ( .A1(n10662), .A2(n10661), .ZN(P1_U3254) );
  NAND3_X1 U13340 ( .A1(n13359), .A2(n13341), .A3(n13333), .ZN(n10666) );
  OAI21_X1 U13341 ( .B1(n6864), .B2(n10664), .A(n10663), .ZN(n10665) );
  NAND2_X1 U13342 ( .A1(n10666), .A2(n10665), .ZN(n10668) );
  AOI22_X1 U13343 ( .A1(n15503), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10667) );
  OAI211_X1 U13344 ( .C1(n13355), .C2(n10669), .A(n10668), .B(n10667), .ZN(
        P3_U3182) );
  INV_X1 U13345 ( .A(n10670), .ZN(n10673) );
  OAI222_X1 U13346 ( .A1(n13717), .A2(n10673), .B1(n10672), .B2(P3_U3151), 
        .C1(n10671), .C2(n13719), .ZN(P3_U3280) );
  XNOR2_X1 U13347 ( .A(n11140), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n11141) );
  AOI21_X1 U13348 ( .B1(n10676), .B2(P2_REG1_REG_6__SCAN_IN), .A(n10674), .ZN(
        n15380) );
  MUX2_X1 U13349 ( .A(n8530), .B(P2_REG1_REG_7__SCAN_IN), .S(n10680), .Z(
        n15381) );
  NOR2_X1 U13350 ( .A1(n15380), .A2(n15381), .ZN(n15379) );
  AOI21_X1 U13351 ( .B1(n10680), .B2(P2_REG1_REG_7__SCAN_IN), .A(n15379), .ZN(
        n10922) );
  XNOR2_X1 U13352 ( .A(n10929), .B(n10675), .ZN(n10921) );
  XOR2_X1 U13353 ( .A(n11141), .B(n11142), .Z(n10693) );
  NAND2_X1 U13354 ( .A1(n10676), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10677) );
  NAND2_X1 U13355 ( .A1(n10678), .A2(n10677), .ZN(n15384) );
  MUX2_X1 U13356 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10679), .S(n10680), .Z(
        n15385) );
  NAND2_X1 U13357 ( .A1(n15384), .A2(n15385), .ZN(n15383) );
  NAND2_X1 U13358 ( .A1(n10680), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10681) );
  NAND2_X1 U13359 ( .A1(n15383), .A2(n10681), .ZN(n10919) );
  MUX2_X1 U13360 ( .A(n10682), .B(P2_REG2_REG_8__SCAN_IN), .S(n10929), .Z(
        n10920) );
  NAND2_X1 U13361 ( .A1(n10919), .A2(n10920), .ZN(n10918) );
  NAND2_X1 U13362 ( .A1(n10683), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10684) );
  NAND2_X1 U13363 ( .A1(n10918), .A2(n10684), .ZN(n10686) );
  INV_X1 U13364 ( .A(n10686), .ZN(n10688) );
  MUX2_X1 U13365 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11133), .S(n11140), .Z(
        n10687) );
  MUX2_X1 U13366 ( .A(n11133), .B(P2_REG2_REG_9__SCAN_IN), .S(n11140), .Z(
        n10685) );
  OAI21_X1 U13367 ( .B1(n10688), .B2(n10687), .A(n11136), .ZN(n10691) );
  NOR2_X1 U13368 ( .A1(n11994), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12585) );
  AOI21_X1 U13369 ( .B1(n15373), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n12585), .ZN(
        n10689) );
  OAI21_X1 U13370 ( .B1(n11134), .B2(n15408), .A(n10689), .ZN(n10690) );
  AOI21_X1 U13371 ( .B1(n15423), .B2(n10691), .A(n10690), .ZN(n10692) );
  OAI21_X1 U13372 ( .B1(n10693), .B2(n15392), .A(n10692), .ZN(P2_U3223) );
  OAI22_X1 U13373 ( .A1(n10694), .A2(n11176), .B1(n12665), .B2(n13866), .ZN(
        n10695) );
  XNOR2_X1 U13374 ( .A(n10695), .B(n12870), .ZN(n11398) );
  INV_X1 U13375 ( .A(n11194), .ZN(n10696) );
  AOI211_X1 U13376 ( .C1(n12670), .C2(n11172), .A(n14166), .B(n10696), .ZN(
        n11401) );
  AOI21_X1 U13377 ( .B1(n15472), .B2(n12670), .A(n11401), .ZN(n10699) );
  XNOR2_X1 U13378 ( .A(n10697), .B(n12870), .ZN(n10698) );
  OAI22_X1 U13379 ( .A1(n8458), .A2(n13812), .B1(n11316), .B2(n13814), .ZN(
        n11051) );
  AOI21_X1 U13380 ( .B1(n15479), .B2(n10698), .A(n11051), .ZN(n11403) );
  OAI211_X1 U13381 ( .C1(n15475), .C2(n11398), .A(n10699), .B(n11403), .ZN(
        n10701) );
  NAND2_X1 U13382 ( .A1(n10701), .A2(n15502), .ZN(n10700) );
  OAI21_X1 U13383 ( .B1(n15502), .B2(n8460), .A(n10700), .ZN(P2_U3501) );
  NAND2_X1 U13384 ( .A1(n10701), .A2(n15496), .ZN(n10702) );
  OAI21_X1 U13385 ( .B1(n15496), .B2(n11973), .A(n10702), .ZN(P2_U3436) );
  INV_X1 U13386 ( .A(n10703), .ZN(n10705) );
  INV_X1 U13387 ( .A(n11525), .ZN(n11643) );
  OAI222_X1 U13388 ( .A1(n15165), .A2(n10704), .B1(n15159), .B2(n10705), .C1(
        P1_U3086), .C2(n11643), .ZN(P1_U3340) );
  OAI222_X1 U13389 ( .A1(n14247), .A2(n11976), .B1(n13019), .B2(n10705), .C1(
        P2_U3088), .C2(n7145), .ZN(P2_U3312) );
  XNOR2_X1 U13390 ( .A(n10706), .B(n10707), .ZN(n10712) );
  XNOR2_X1 U13391 ( .A(n10708), .B(n10707), .ZN(n10710) );
  AOI22_X1 U13392 ( .A1(n15010), .A2(n14585), .B1(n14583), .B2(n15008), .ZN(
        n10709) );
  OAI21_X1 U13393 ( .B1(n10710), .B2(n14988), .A(n10709), .ZN(n10711) );
  AOI21_X1 U13394 ( .B1(n15078), .B2(n10712), .A(n10711), .ZN(n11030) );
  INV_X1 U13395 ( .A(n10713), .ZN(n10714) );
  OAI211_X1 U13396 ( .C1(n10714), .C2(n7686), .A(n6432), .B(n10901), .ZN(
        n11035) );
  AND2_X1 U13397 ( .A1(n11030), .A2(n11035), .ZN(n10719) );
  AOI22_X1 U13398 ( .A1(n11749), .A2(n6434), .B1(n15320), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n10715) );
  OAI21_X1 U13399 ( .B1(n10719), .B2(n15320), .A(n10715), .ZN(P1_U3531) );
  INV_X1 U13400 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10716) );
  OAI22_X1 U13401 ( .A1(n15143), .A2(n7686), .B1(n15319), .B2(n10716), .ZN(
        n10717) );
  INV_X1 U13402 ( .A(n10717), .ZN(n10718) );
  OAI21_X1 U13403 ( .B1(n10719), .B2(n15317), .A(n10718), .ZN(P1_U3468) );
  MUX2_X1 U13404 ( .A(n11843), .B(P1_REG2_REG_12__SCAN_IN), .S(n11006), .Z(
        n10725) );
  NAND2_X1 U13405 ( .A1(n10720), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10721) );
  NAND2_X1 U13406 ( .A1(n10722), .A2(n10721), .ZN(n10724) );
  INV_X1 U13407 ( .A(n11002), .ZN(n10723) );
  AOI21_X1 U13408 ( .B1(n10725), .B2(n10724), .A(n10723), .ZN(n10735) );
  AND2_X1 U13409 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14446) );
  NOR2_X1 U13410 ( .A1(n14719), .A2(n10726), .ZN(n10727) );
  AOI211_X1 U13411 ( .C1(n15269), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n14446), 
        .B(n10727), .ZN(n10734) );
  INV_X1 U13412 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n12244) );
  XNOR2_X1 U13413 ( .A(n11006), .B(n12244), .ZN(n10731) );
  NAND2_X1 U13414 ( .A1(n10729), .A2(n10728), .ZN(n10730) );
  NAND2_X1 U13415 ( .A1(n10730), .A2(n10731), .ZN(n11010) );
  OAI21_X1 U13416 ( .B1(n10731), .B2(n10730), .A(n11010), .ZN(n10732) );
  NAND2_X1 U13417 ( .A1(n10732), .A2(n14739), .ZN(n10733) );
  OAI211_X1 U13418 ( .C1(n10735), .C2(n14735), .A(n10734), .B(n10733), .ZN(
        P1_U3255) );
  INV_X1 U13419 ( .A(n10736), .ZN(n10737) );
  NOR2_X1 U13420 ( .A1(n10738), .A2(n10737), .ZN(n10739) );
  XNOR2_X1 U13421 ( .A(n10740), .B(n10739), .ZN(n10750) );
  XNOR2_X1 U13422 ( .A(n10741), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n10748) );
  NOR2_X1 U13423 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8995), .ZN(n11186) );
  AOI21_X1 U13424 ( .B1(n15503), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11186), .ZN(
        n10745) );
  NAND2_X1 U13425 ( .A1(n13348), .A2(n10743), .ZN(n10744) );
  OAI211_X1 U13426 ( .C1(n13355), .C2(n10746), .A(n10745), .B(n10744), .ZN(
        n10747) );
  AOI21_X1 U13427 ( .B1(n10748), .B2(n9642), .A(n10747), .ZN(n10749) );
  OAI21_X1 U13428 ( .B1(n13359), .B2(n10750), .A(n10749), .ZN(P3_U3187) );
  INV_X1 U13429 ( .A(n13891), .ZN(n13883) );
  INV_X1 U13430 ( .A(n10751), .ZN(n10753) );
  INV_X1 U13431 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10752) );
  OAI222_X1 U13432 ( .A1(P2_U3088), .A2(n13883), .B1(n13019), .B2(n10753), 
        .C1(n10752), .C2(n14247), .ZN(P2_U3311) );
  INV_X1 U13433 ( .A(n12087), .ZN(n11536) );
  OAI222_X1 U13434 ( .A1(n15165), .A2(n10754), .B1(n15159), .B2(n10753), .C1(
        n11536), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13435 ( .A(n12661), .ZN(n10755) );
  NOR2_X1 U13436 ( .A1(n12663), .A2(n10755), .ZN(n12871) );
  INV_X1 U13437 ( .A(n14072), .ZN(n11872) );
  NOR2_X1 U13438 ( .A1(n15479), .A2(n11872), .ZN(n10756) );
  NAND2_X1 U13439 ( .A1(n13866), .A2(n13802), .ZN(n11065) );
  OAI21_X1 U13440 ( .B1(n10756), .B2(n12871), .A(n11065), .ZN(n10995) );
  INV_X1 U13441 ( .A(n10995), .ZN(n10758) );
  INV_X1 U13442 ( .A(n10997), .ZN(n10757) );
  OAI211_X1 U13443 ( .C1(n12871), .C2(n14222), .A(n10758), .B(n10757), .ZN(
        n10760) );
  NAND2_X1 U13444 ( .A1(n10760), .A2(n15502), .ZN(n10759) );
  OAI21_X1 U13445 ( .B1(n15502), .B2(n10635), .A(n10759), .ZN(P2_U3499) );
  NAND2_X1 U13446 ( .A1(n10760), .A2(n15496), .ZN(n10761) );
  OAI21_X1 U13447 ( .B1(n15496), .B2(n8439), .A(n10761), .ZN(P2_U3430) );
  AOI222_X1 U13448 ( .A1(n10763), .A2(n13702), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13315), .C1(SI_16_), .C2(n10762), .ZN(n10764) );
  INV_X1 U13449 ( .A(n10764), .ZN(P3_U3279) );
  INV_X1 U13450 ( .A(n10765), .ZN(n10768) );
  INV_X1 U13451 ( .A(n14698), .ZN(n14695) );
  OAI222_X1 U13452 ( .A1(n15165), .A2(n10766), .B1(n15159), .B2(n10768), .C1(
        n14695), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U13453 ( .A(n12323), .ZN(n15407) );
  OAI222_X1 U13454 ( .A1(P2_U3088), .A2(n15407), .B1(n13019), .B2(n10768), 
        .C1(n10767), .C2(n14247), .ZN(P2_U3313) );
  AOI21_X1 U13455 ( .B1(n10770), .B2(n10769), .A(n6642), .ZN(n10787) );
  INV_X1 U13456 ( .A(n10771), .ZN(n10773) );
  NAND3_X1 U13457 ( .A1(n10774), .A2(n10773), .A3(n10772), .ZN(n10775) );
  AND2_X1 U13458 ( .A1(n10776), .A2(n10775), .ZN(n10778) );
  NAND2_X1 U13459 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U13460 ( .A1(n15503), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10777) );
  OAI211_X1 U13461 ( .C1(n13341), .C2(n10778), .A(n11083), .B(n10777), .ZN(
        n10784) );
  AOI21_X1 U13462 ( .B1(n10781), .B2(n10780), .A(n10779), .ZN(n10782) );
  NOR2_X1 U13463 ( .A1(n10782), .A2(n13333), .ZN(n10783) );
  AOI211_X1 U13464 ( .C1(n13339), .C2(n10785), .A(n10784), .B(n10783), .ZN(
        n10786) );
  OAI21_X1 U13465 ( .B1(n10787), .B2(n13359), .A(n10786), .ZN(P3_U3186) );
  NAND2_X1 U13466 ( .A1(n10788), .A2(n6531), .ZN(n10789) );
  NAND2_X1 U13467 ( .A1(n10790), .A2(n10789), .ZN(n11022) );
  INV_X1 U13468 ( .A(n11022), .ZN(n10797) );
  NAND2_X1 U13469 ( .A1(n14584), .A2(n14351), .ZN(n10792) );
  NAND2_X1 U13470 ( .A1(n6434), .A2(n14346), .ZN(n10791) );
  NAND2_X1 U13471 ( .A1(n10792), .A2(n10791), .ZN(n10793) );
  XNOR2_X1 U13472 ( .A(n10793), .B(n11660), .ZN(n10798) );
  AND2_X1 U13473 ( .A1(n6434), .A2(n14351), .ZN(n10795) );
  AOI21_X1 U13474 ( .B1(n14584), .B2(n10794), .A(n10795), .ZN(n10799) );
  XNOR2_X1 U13475 ( .A(n10798), .B(n10799), .ZN(n11025) );
  INV_X1 U13476 ( .A(n11025), .ZN(n10796) );
  INV_X1 U13477 ( .A(n10798), .ZN(n10801) );
  INV_X1 U13478 ( .A(n10799), .ZN(n10800) );
  NAND2_X1 U13479 ( .A1(n10801), .A2(n10800), .ZN(n10802) );
  NAND2_X1 U13480 ( .A1(n6430), .A2(n14346), .ZN(n10803) );
  NAND2_X1 U13481 ( .A1(n10804), .A2(n10803), .ZN(n10805) );
  NAND2_X1 U13482 ( .A1(n14583), .A2(n10794), .ZN(n10807) );
  NAND2_X1 U13483 ( .A1(n6430), .A2(n14351), .ZN(n10806) );
  NAND2_X1 U13484 ( .A1(n10807), .A2(n10806), .ZN(n11112) );
  INV_X1 U13485 ( .A(n11112), .ZN(n11114) );
  XNOR2_X1 U13486 ( .A(n11113), .B(n11114), .ZN(n10808) );
  XNOR2_X1 U13487 ( .A(n11118), .B(n10808), .ZN(n10814) );
  OAI22_X1 U13488 ( .A1(n10810), .A2(n15032), .B1(n11284), .B2(n14993), .ZN(
        n10898) );
  NAND2_X1 U13489 ( .A1(n10898), .A2(n14547), .ZN(n10811) );
  NAND2_X1 U13490 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14613) );
  OAI211_X1 U13491 ( .C1(n14556), .C2(n10902), .A(n10811), .B(n14613), .ZN(
        n10812) );
  AOI21_X1 U13492 ( .B1(n6430), .B2(n10393), .A(n10812), .ZN(n10813) );
  OAI21_X1 U13493 ( .B1(n10814), .B2(n14561), .A(n10813), .ZN(P1_U3230) );
  XOR2_X1 U13494 ( .A(n10816), .B(n10815), .Z(n10831) );
  OAI21_X1 U13495 ( .B1(n10819), .B2(n10818), .A(n10817), .ZN(n10829) );
  AND2_X1 U13496 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11377) );
  AOI21_X1 U13497 ( .B1(n15503), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11377), .ZN(
        n10821) );
  OAI21_X1 U13498 ( .B1(n13355), .B2(n10822), .A(n10821), .ZN(n10828) );
  AOI21_X1 U13499 ( .B1(n10825), .B2(n10824), .A(n10823), .ZN(n10826) );
  NOR2_X1 U13500 ( .A1(n10826), .A2(n13333), .ZN(n10827) );
  AOI211_X1 U13501 ( .C1(n13348), .C2(n10829), .A(n10828), .B(n10827), .ZN(
        n10830) );
  OAI21_X1 U13502 ( .B1(n10831), .B2(n13359), .A(n10830), .ZN(P3_U3188) );
  XOR2_X1 U13503 ( .A(P3_REG1_REG_7__SCAN_IN), .B(n10832), .Z(n10845) );
  XNOR2_X1 U13504 ( .A(n10834), .B(n10833), .ZN(n10843) );
  AOI21_X1 U13505 ( .B1(n10837), .B2(n10836), .A(n10835), .ZN(n10838) );
  NOR2_X1 U13506 ( .A1(n10838), .A2(n13341), .ZN(n10842) );
  INV_X1 U13507 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n12005) );
  NOR2_X1 U13508 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12005), .ZN(n11543) );
  AOI21_X1 U13509 ( .B1(n15503), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11543), .ZN(
        n10839) );
  OAI21_X1 U13510 ( .B1(n13355), .B2(n10840), .A(n10839), .ZN(n10841) );
  AOI211_X1 U13511 ( .C1(n10843), .C2(n13270), .A(n10842), .B(n10841), .ZN(
        n10844) );
  OAI21_X1 U13512 ( .B1(n10845), .B2(n13333), .A(n10844), .ZN(P3_U3189) );
  NAND2_X1 U13513 ( .A1(n15545), .A2(n10936), .ZN(n12395) );
  NAND2_X1 U13514 ( .A1(n15542), .A2(n12395), .ZN(n12545) );
  AND2_X1 U13515 ( .A1(n10846), .A2(n15541), .ZN(n10847) );
  NAND2_X1 U13516 ( .A1(n12545), .A2(n10847), .ZN(n10849) );
  NAND2_X1 U13517 ( .A1(n15533), .A2(n15531), .ZN(n10848) );
  NAND2_X1 U13518 ( .A1(n10849), .A2(n10848), .ZN(n11018) );
  NOR2_X1 U13519 ( .A1(n15612), .A2(n9569), .ZN(n10850) );
  AOI21_X1 U13520 ( .B1(n15612), .B2(n11018), .A(n10850), .ZN(n10851) );
  OAI21_X1 U13521 ( .B1(n10936), .B2(n13598), .A(n10851), .ZN(P3_U3459) );
  INV_X1 U13522 ( .A(n10863), .ZN(n10856) );
  NAND3_X1 U13523 ( .A1(n10854), .A2(n10853), .A3(n10852), .ZN(n10855) );
  AOI21_X1 U13524 ( .B1(n10872), .B2(n10856), .A(n10855), .ZN(n10857) );
  OAI21_X1 U13525 ( .B1(n10868), .B2(n10858), .A(n10857), .ZN(n10859) );
  NAND2_X1 U13526 ( .A1(n10859), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10861) );
  NAND2_X1 U13527 ( .A1(n10872), .A2(n12580), .ZN(n10860) );
  NOR2_X1 U13528 ( .A1(n13195), .A2(P3_U3151), .ZN(n10917) );
  NAND3_X1 U13529 ( .A1(n10868), .A2(n15541), .A3(n10862), .ZN(n10865) );
  OR2_X1 U13530 ( .A1(n10872), .A2(n10863), .ZN(n10864) );
  NAND2_X1 U13531 ( .A1(n10865), .A2(n10864), .ZN(n10867) );
  OR2_X1 U13532 ( .A1(n10868), .A2(n15526), .ZN(n10870) );
  INV_X1 U13533 ( .A(n15533), .ZN(n10908) );
  INV_X1 U13534 ( .A(n12580), .ZN(n10871) );
  INV_X1 U13535 ( .A(n10890), .ZN(n10873) );
  OAI22_X1 U13536 ( .A1(n13177), .A2(n10936), .B1(n10908), .B2(n13193), .ZN(
        n10874) );
  AOI21_X1 U13537 ( .B1(n13169), .B2(n12545), .A(n10874), .ZN(n10875) );
  OAI21_X1 U13538 ( .B1(n10917), .B2(n10876), .A(n10875), .ZN(P3_U3172) );
  INV_X1 U13539 ( .A(n12575), .ZN(n10877) );
  AND2_X1 U13540 ( .A1(n10878), .A2(n10877), .ZN(n10879) );
  OAI21_X1 U13541 ( .B1(n11153), .B2(n12394), .A(n11640), .ZN(n10881) );
  NAND2_X1 U13542 ( .A1(n12546), .A2(n13035), .ZN(n10883) );
  NAND2_X1 U13543 ( .A1(n6431), .A2(n9470), .ZN(n10882) );
  NAND2_X1 U13544 ( .A1(n10883), .A2(n10882), .ZN(n10888) );
  INV_X1 U13545 ( .A(n15547), .ZN(n10887) );
  OAI21_X1 U13546 ( .B1(n6431), .B2(n15547), .A(n10884), .ZN(n10885) );
  NAND2_X1 U13547 ( .A1(n10888), .A2(n10885), .ZN(n10911) );
  NAND3_X1 U13548 ( .A1(n6431), .A2(n15542), .A3(n12546), .ZN(n10886) );
  OAI211_X1 U13549 ( .C1(n10888), .C2(n10887), .A(n10911), .B(n10886), .ZN(
        n10893) );
  INV_X1 U13550 ( .A(n15544), .ZN(n11156) );
  NOR2_X2 U13551 ( .A1(n10890), .A2(n10889), .ZN(n13190) );
  AOI22_X1 U13552 ( .A1(n13196), .A2(n6659), .B1(n13190), .B2(n15545), .ZN(
        n10891) );
  OAI21_X1 U13553 ( .B1(n11156), .B2(n13193), .A(n10891), .ZN(n10892) );
  AOI21_X1 U13554 ( .B1(n13169), .B2(n10893), .A(n10892), .ZN(n10894) );
  OAI21_X1 U13555 ( .B1(n10917), .B2(n15554), .A(n10894), .ZN(P3_U3162) );
  XNOR2_X1 U13556 ( .A(n10895), .B(n10896), .ZN(n15315) );
  XNOR2_X1 U13557 ( .A(n10897), .B(n10896), .ZN(n10899) );
  AOI21_X1 U13558 ( .B1(n10899), .B2(n14874), .A(n10898), .ZN(n15313) );
  MUX2_X1 U13559 ( .A(n10900), .B(n15313), .S(n15305), .Z(n10906) );
  AOI211_X1 U13560 ( .C1(n6430), .C2(n10901), .A(n15015), .B(n11105), .ZN(
        n15309) );
  OAI22_X1 U13561 ( .A1(n15279), .A2(n10903), .B1(n10902), .B2(n14997), .ZN(
        n10904) );
  AOI21_X1 U13562 ( .B1(n15309), .B2(n15273), .A(n10904), .ZN(n10905) );
  OAI211_X1 U13563 ( .C1(n15023), .C2(n15315), .A(n10906), .B(n10905), .ZN(
        P1_U3289) );
  OAI22_X1 U13564 ( .A1(n15524), .A2(n13177), .B1(n13151), .B2(n10908), .ZN(
        n10907) );
  AOI21_X1 U13565 ( .B1(n13181), .B2(n15532), .A(n10907), .ZN(n10916) );
  XNOR2_X1 U13566 ( .A(n11036), .B(n15544), .ZN(n10913) );
  XNOR2_X1 U13567 ( .A(n6431), .B(n6659), .ZN(n10909) );
  NAND2_X1 U13568 ( .A1(n10909), .A2(n10908), .ZN(n10910) );
  NAND2_X1 U13569 ( .A1(n10912), .A2(n10913), .ZN(n11041) );
  OAI21_X1 U13570 ( .B1(n10913), .B2(n10912), .A(n11041), .ZN(n10914) );
  NAND2_X1 U13571 ( .A1(n10914), .A2(n13169), .ZN(n10915) );
  OAI211_X1 U13572 ( .C1(n10917), .C2(n15527), .A(n10916), .B(n10915), .ZN(
        P3_U3177) );
  OAI211_X1 U13573 ( .C1(n10920), .C2(n10919), .A(n15423), .B(n10918), .ZN(
        n10925) );
  XOR2_X1 U13574 ( .A(n10922), .B(n10921), .Z(n10923) );
  NAND2_X1 U13575 ( .A1(n15419), .A2(n10923), .ZN(n10924) );
  NAND2_X1 U13576 ( .A1(n10925), .A2(n10924), .ZN(n10927) );
  NAND2_X1 U13577 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11585) );
  INV_X1 U13578 ( .A(n11585), .ZN(n10926) );
  AOI211_X1 U13579 ( .C1(n15373), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n10927), .B(
        n10926), .ZN(n10928) );
  OAI21_X1 U13580 ( .B1(n10929), .B2(n15408), .A(n10928), .ZN(P2_U3222) );
  INV_X1 U13581 ( .A(n10930), .ZN(n10931) );
  OAI222_X1 U13582 ( .A1(n13719), .A2(n10932), .B1(n9634), .B2(P3_U3151), .C1(
        n13717), .C2(n10931), .ZN(P3_U3278) );
  INV_X1 U13583 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10933) );
  NOR2_X1 U13584 ( .A1(n15600), .A2(n10933), .ZN(n10934) );
  AOI21_X1 U13585 ( .B1(n15600), .B2(n11018), .A(n10934), .ZN(n10935) );
  OAI21_X1 U13586 ( .B1(n10936), .B2(n13654), .A(n10935), .ZN(P3_U3390) );
  AOI21_X1 U13587 ( .B1(n10939), .B2(n10938), .A(n10937), .ZN(n10952) );
  XNOR2_X1 U13588 ( .A(n10941), .B(n10940), .ZN(n10950) );
  AOI21_X1 U13589 ( .B1(n6640), .B2(n10943), .A(n10942), .ZN(n10948) );
  NOR2_X1 U13590 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10944), .ZN(n13086) );
  AOI21_X1 U13591 ( .B1(n15503), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n13086), .ZN(
        n10947) );
  NAND2_X1 U13592 ( .A1(n13339), .A2(n10945), .ZN(n10946) );
  OAI211_X1 U13593 ( .C1(n10948), .C2(n13341), .A(n10947), .B(n10946), .ZN(
        n10949) );
  AOI21_X1 U13594 ( .B1(n10950), .B2(n13270), .A(n10949), .ZN(n10951) );
  OAI21_X1 U13595 ( .B1(n10952), .B2(n13333), .A(n10951), .ZN(P3_U3190) );
  INV_X1 U13596 ( .A(n13906), .ZN(n10954) );
  INV_X1 U13597 ( .A(n10953), .ZN(n10955) );
  OAI222_X1 U13598 ( .A1(P2_U3088), .A2(n10954), .B1(n13019), .B2(n10955), 
        .C1(n11977), .C2(n14247), .ZN(P2_U3310) );
  INV_X1 U13599 ( .A(n14707), .ZN(n14710) );
  OAI222_X1 U13600 ( .A1(n15165), .A2(n10956), .B1(n15159), .B2(n10955), .C1(
        n14710), .C2(P1_U3086), .ZN(P1_U3338) );
  XNOR2_X1 U13601 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n10961) );
  XNOR2_X1 U13602 ( .A(n10970), .B(n10961), .ZN(n15170) );
  NAND2_X1 U13603 ( .A1(n15171), .A2(n15170), .ZN(n10965) );
  INV_X1 U13604 ( .A(n10962), .ZN(n10963) );
  NAND2_X1 U13605 ( .A1(n10963), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10964) );
  INV_X1 U13606 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10966) );
  XNOR2_X1 U13607 ( .A(n10975), .B(n10966), .ZN(n15172) );
  INV_X1 U13608 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14644) );
  INV_X1 U13609 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10967) );
  NOR2_X1 U13610 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10967), .ZN(n10968) );
  INV_X1 U13611 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10971) );
  NAND2_X1 U13612 ( .A1(n10972), .A2(n10971), .ZN(n10979) );
  INV_X1 U13613 ( .A(n10972), .ZN(n10973) );
  NAND2_X1 U13614 ( .A1(n10973), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U13615 ( .A1(n10979), .A2(n10974), .ZN(n10978) );
  XNOR2_X1 U13616 ( .A(n10978), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15173) );
  NAND2_X1 U13617 ( .A1(n15172), .A2(n15173), .ZN(n10977) );
  NAND2_X1 U13618 ( .A1(n10975), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U13619 ( .A1(n10977), .A2(n10976), .ZN(n10986) );
  INV_X1 U13620 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14657) );
  INV_X1 U13621 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10981) );
  NAND2_X1 U13622 ( .A1(n10981), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n11613) );
  NAND2_X1 U13623 ( .A1(n10982), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n10983) );
  AND2_X1 U13624 ( .A1(n11613), .A2(n10983), .ZN(n11615) );
  INV_X1 U13625 ( .A(n11615), .ZN(n10984) );
  XNOR2_X1 U13626 ( .A(n11616), .B(n10984), .ZN(n10985) );
  INV_X1 U13627 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U13628 ( .A1(n10988), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10989) );
  NAND2_X1 U13629 ( .A1(n11612), .A2(n10989), .ZN(SUB_1596_U55) );
  AND2_X1 U13630 ( .A1(n10990), .A2(n15459), .ZN(n10991) );
  NAND2_X1 U13631 ( .A1(n10992), .A2(n10991), .ZN(n10993) );
  OR2_X1 U13632 ( .A1(n13017), .A2(n6993), .ZN(n10996) );
  INV_X1 U13633 ( .A(n10996), .ZN(n12911) );
  NAND2_X1 U13634 ( .A1(n12911), .A2(n12899), .ZN(n10994) );
  AOI21_X1 U13635 ( .B1(n10997), .B2(n10996), .A(n10995), .ZN(n10998) );
  OAI22_X1 U13636 ( .A1(n10998), .A2(n6438), .B1(n11067), .B2(n15434), .ZN(
        n10999) );
  AOI21_X1 U13637 ( .B1(n6438), .B2(P2_REG2_REG_0__SCAN_IN), .A(n10999), .ZN(
        n11000) );
  OAI21_X1 U13638 ( .B1(n12871), .B2(n12149), .A(n11000), .ZN(P2_U3265) );
  OR2_X1 U13639 ( .A1(n11006), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11001) );
  NAND2_X1 U13640 ( .A1(n11002), .A2(n11001), .ZN(n11005) );
  MUX2_X1 U13641 ( .A(n11805), .B(P1_REG2_REG_13__SCAN_IN), .S(n11520), .Z(
        n11004) );
  INV_X1 U13642 ( .A(n14701), .ZN(n11003) );
  AOI211_X1 U13643 ( .C1(n11005), .C2(n11004), .A(n14735), .B(n11003), .ZN(
        n11017) );
  INV_X1 U13644 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n12305) );
  XNOR2_X1 U13645 ( .A(n11520), .B(n12305), .ZN(n11008) );
  OR2_X1 U13646 ( .A1(n11006), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11009) );
  AND2_X1 U13647 ( .A1(n11008), .A2(n11009), .ZN(n11007) );
  INV_X1 U13648 ( .A(n14692), .ZN(n11012) );
  AOI21_X1 U13649 ( .B1(n11010), .B2(n11009), .A(n11008), .ZN(n11011) );
  NOR3_X1 U13650 ( .A1(n11012), .A2(n11011), .A3(n11646), .ZN(n11016) );
  NAND2_X1 U13651 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12233)
         );
  NAND2_X1 U13652 ( .A1(n15269), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11013) );
  OAI211_X1 U13653 ( .C1(n14719), .C2(n11014), .A(n12233), .B(n11013), .ZN(
        n11015) );
  OR3_X1 U13654 ( .A1(n11017), .A2(n11016), .A3(n11015), .ZN(P1_U3256) );
  AOI22_X1 U13655 ( .A1(n15559), .A2(n11018), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n15518), .ZN(n11021) );
  NAND2_X1 U13656 ( .A1(n6428), .A2(n11019), .ZN(n11020) );
  OAI211_X1 U13657 ( .C1(n9570), .C2(n15559), .A(n11021), .B(n11020), .ZN(
        P3_U3233) );
  INV_X1 U13658 ( .A(n11023), .ZN(n11024) );
  AOI211_X1 U13659 ( .C1(n11025), .C2(n11022), .A(n14561), .B(n11024), .ZN(
        n11029) );
  AOI22_X1 U13660 ( .A1(n14534), .A2(n14583), .B1(n14377), .B2(n14585), .ZN(
        n11027) );
  MUX2_X1 U13661 ( .A(n14556), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n11026) );
  OAI211_X1 U13662 ( .C1(n7686), .C2(n14550), .A(n11027), .B(n11026), .ZN(
        n11028) );
  OR2_X1 U13663 ( .A1(n11029), .A2(n11028), .ZN(P1_U3218) );
  MUX2_X1 U13664 ( .A(n11031), .B(n11030), .S(n15305), .Z(n11034) );
  AOI22_X1 U13665 ( .A1(n14980), .A2(n6434), .B1(n15301), .B2(n7834), .ZN(
        n11033) );
  OAI211_X1 U13666 ( .C1(n14984), .C2(n11035), .A(n11034), .B(n11033), .ZN(
        P1_U3290) );
  NAND2_X1 U13667 ( .A1(n11036), .A2(n11156), .ZN(n11038) );
  XNOR2_X1 U13668 ( .A(n11072), .B(n15532), .ZN(n11039) );
  AOI21_X1 U13669 ( .B1(n11041), .B2(n11038), .A(n11039), .ZN(n11046) );
  AND2_X1 U13670 ( .A1(n11039), .A2(n11038), .ZN(n11040) );
  NAND2_X1 U13671 ( .A1(n11041), .A2(n11040), .ZN(n11075) );
  NAND2_X1 U13672 ( .A1(n11075), .A2(n13169), .ZN(n11045) );
  INV_X1 U13673 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11164) );
  MUX2_X1 U13674 ( .A(P3_U3151), .B(n13195), .S(n11164), .Z(n11043) );
  OAI22_X1 U13675 ( .A1(n11163), .A2(n13177), .B1(n13151), .B2(n11156), .ZN(
        n11042) );
  AOI211_X1 U13676 ( .C1(n13181), .C2(n13213), .A(n11043), .B(n11042), .ZN(
        n11044) );
  OAI21_X1 U13677 ( .B1(n11046), .B2(n11045), .A(n11044), .ZN(P3_U3158) );
  NOR2_X1 U13678 ( .A1(n11047), .A2(n15461), .ZN(n11205) );
  XNOR2_X1 U13679 ( .A(n11049), .B(n11048), .ZN(n11050) );
  NAND2_X1 U13680 ( .A1(n11050), .A2(n13822), .ZN(n11053) );
  AOI22_X1 U13681 ( .A1(n13826), .A2(n11051), .B1(n15332), .B2(n12670), .ZN(
        n11052) );
  OAI211_X1 U13682 ( .C1(n11205), .C2(n11394), .A(n11053), .B(n11052), .ZN(
        P2_U3209) );
  INV_X1 U13683 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11968) );
  NAND2_X1 U13684 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  XNOR2_X1 U13685 ( .A(n12933), .B(n13862), .ZN(n12872) );
  XNOR2_X1 U13686 ( .A(n11056), .B(n12872), .ZN(n11236) );
  OAI22_X1 U13687 ( .A1(n11191), .A2(n13812), .B1(n11387), .B2(n13814), .ZN(
        n12923) );
  AOI21_X1 U13688 ( .B1(n15444), .B2(n12933), .A(n14166), .ZN(n11057) );
  AND2_X1 U13689 ( .A1(n11057), .A2(n6638), .ZN(n11232) );
  AOI211_X1 U13690 ( .C1(n15472), .C2(n12933), .A(n12923), .B(n11232), .ZN(
        n11060) );
  XNOR2_X1 U13691 ( .A(n11058), .B(n12872), .ZN(n11233) );
  NAND2_X1 U13692 ( .A1(n11233), .A2(n15479), .ZN(n11059) );
  OAI211_X1 U13693 ( .C1(n11236), .C2(n15475), .A(n11060), .B(n11059), .ZN(
        n11062) );
  NAND2_X1 U13694 ( .A1(n11062), .A2(n15496), .ZN(n11061) );
  OAI21_X1 U13695 ( .B1(n15496), .B2(n11968), .A(n11061), .ZN(P2_U3445) );
  NAND2_X1 U13696 ( .A1(n11062), .A2(n15502), .ZN(n11063) );
  OAI21_X1 U13697 ( .B1(n15502), .B2(n8512), .A(n11063), .ZN(P2_U3504) );
  OAI22_X1 U13698 ( .A1(n15325), .A2(n11065), .B1(n11064), .B2(n15327), .ZN(
        n11069) );
  OAI22_X1 U13699 ( .A1(n13790), .A2(n12661), .B1(n11205), .B2(n11067), .ZN(
        n11068) );
  AOI211_X1 U13700 ( .C1(n11070), .C2(n15332), .A(n11069), .B(n11068), .ZN(
        n11071) );
  INV_X1 U13701 ( .A(n11071), .ZN(P2_U3204) );
  INV_X1 U13702 ( .A(n11072), .ZN(n11073) );
  NAND2_X1 U13703 ( .A1(n11073), .A2(n15532), .ZN(n11074) );
  XNOR2_X1 U13704 ( .A(n11076), .B(n11328), .ZN(n11077) );
  INV_X1 U13705 ( .A(n13213), .ZN(n11254) );
  NAND2_X1 U13706 ( .A1(n11077), .A2(n11254), .ZN(n11180) );
  INV_X1 U13707 ( .A(n11077), .ZN(n11078) );
  NAND2_X1 U13708 ( .A1(n11078), .A2(n13213), .ZN(n11079) );
  INV_X1 U13709 ( .A(n11181), .ZN(n11080) );
  AOI21_X1 U13710 ( .B1(n11082), .B2(n11081), .A(n11080), .ZN(n11088) );
  INV_X1 U13711 ( .A(n11329), .ZN(n11086) );
  AOI22_X1 U13712 ( .A1(n13181), .A2(n13212), .B1(n13190), .B2(n15532), .ZN(
        n11084) );
  OAI211_X1 U13713 ( .C1(n13177), .C2(n12413), .A(n11084), .B(n11083), .ZN(
        n11085) );
  AOI21_X1 U13714 ( .B1(n11086), .B2(n13195), .A(n11085), .ZN(n11087) );
  OAI21_X1 U13715 ( .B1(n11088), .B2(n13199), .A(n11087), .ZN(P3_U3170) );
  INV_X1 U13716 ( .A(n11089), .ZN(n11091) );
  OAI222_X1 U13717 ( .A1(n13717), .A2(n11091), .B1(n13719), .B2(n11090), .C1(
        n13354), .C2(P3_U3151), .ZN(P3_U3277) );
  OAI21_X1 U13718 ( .B1(n11099), .B2(n11093), .A(n11092), .ZN(n11097) );
  NAND2_X1 U13719 ( .A1(n14583), .A2(n15010), .ZN(n11095) );
  NAND2_X1 U13720 ( .A1(n14581), .A2(n15008), .ZN(n11094) );
  NAND2_X1 U13721 ( .A1(n11095), .A2(n11094), .ZN(n11096) );
  AOI21_X1 U13722 ( .B1(n11097), .B2(n14874), .A(n11096), .ZN(n11104) );
  NAND2_X1 U13723 ( .A1(n11100), .A2(n11099), .ZN(n11101) );
  NAND2_X1 U13724 ( .A1(n11098), .A2(n11101), .ZN(n11102) );
  NAND2_X1 U13725 ( .A1(n11102), .A2(n15078), .ZN(n11103) );
  NAND2_X1 U13726 ( .A1(n11104), .A2(n11103), .ZN(n11210) );
  OAI211_X1 U13727 ( .C1(n11105), .C2(n11120), .A(n6432), .B(n11288), .ZN(
        n11216) );
  INV_X1 U13728 ( .A(n11216), .ZN(n11106) );
  NOR2_X1 U13729 ( .A1(n11210), .A2(n11106), .ZN(n11111) );
  AOI22_X1 U13730 ( .A1(n11749), .A2(n11213), .B1(n15320), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n11107) );
  OAI21_X1 U13731 ( .B1(n11111), .B2(n15320), .A(n11107), .ZN(P1_U3533) );
  INV_X1 U13732 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11108) );
  OAI22_X1 U13733 ( .A1(n15143), .A2(n11120), .B1(n15319), .B2(n11108), .ZN(
        n11109) );
  INV_X1 U13734 ( .A(n11109), .ZN(n11110) );
  OAI21_X1 U13735 ( .B1(n11111), .B2(n15317), .A(n11110), .ZN(P1_U3474) );
  AND2_X1 U13736 ( .A1(n11113), .A2(n11112), .ZN(n11117) );
  INV_X1 U13737 ( .A(n11113), .ZN(n11115) );
  NAND2_X1 U13738 ( .A1(n11115), .A2(n11114), .ZN(n11116) );
  OAI22_X1 U13739 ( .A1(n11284), .A2(n14413), .B1(n11120), .B2(n14414), .ZN(
        n11119) );
  XNOR2_X1 U13740 ( .A(n11119), .B(n14359), .ZN(n11217) );
  OR2_X1 U13741 ( .A1(n11120), .A2(n14413), .ZN(n11121) );
  OAI21_X1 U13742 ( .B1(n11284), .B2(n14411), .A(n11121), .ZN(n11219) );
  XNOR2_X1 U13743 ( .A(n11217), .B(n11219), .ZN(n11122) );
  XNOR2_X1 U13744 ( .A(n11218), .B(n11122), .ZN(n11128) );
  INV_X1 U13745 ( .A(n14556), .ZN(n14418) );
  INV_X1 U13746 ( .A(n11123), .ZN(n11212) );
  AOI22_X1 U13747 ( .A1(n14418), .A2(n11212), .B1(n14377), .B2(n14583), .ZN(
        n11126) );
  NAND2_X1 U13748 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14629) );
  NAND2_X1 U13749 ( .A1(n10393), .A2(n11213), .ZN(n11125) );
  NAND2_X1 U13750 ( .A1(n14534), .A2(n14581), .ZN(n11124) );
  NAND4_X1 U13751 ( .A1(n11126), .A2(n14629), .A3(n11125), .A4(n11124), .ZN(
        n11127) );
  AOI21_X1 U13752 ( .B1(n11128), .B2(n14540), .A(n11127), .ZN(n11129) );
  INV_X1 U13753 ( .A(n11129), .ZN(P1_U3227) );
  INV_X1 U13754 ( .A(n14727), .ZN(n14718) );
  OAI222_X1 U13755 ( .A1(n15165), .A2(n11974), .B1(n15159), .B2(n11131), .C1(
        n14718), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13756 ( .A(n15422), .ZN(n11132) );
  OAI222_X1 U13757 ( .A1(P2_U3088), .A2(n11132), .B1(n13019), .B2(n11131), 
        .C1(n11130), .C2(n14247), .ZN(P2_U3309) );
  NAND2_X1 U13758 ( .A1(n11134), .A2(n11133), .ZN(n11135) );
  AND2_X1 U13759 ( .A1(n11136), .A2(n11135), .ZN(n11139) );
  INV_X1 U13760 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11137) );
  MUX2_X1 U13761 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n11137), .S(n11268), .Z(
        n11138) );
  NAND2_X1 U13762 ( .A1(n11139), .A2(n11138), .ZN(n11265) );
  OAI211_X1 U13763 ( .C1(n11139), .C2(n11138), .A(n11265), .B(n15423), .ZN(
        n11149) );
  NAND2_X1 U13764 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n12187)
         );
  XNOR2_X1 U13765 ( .A(n11268), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n11144) );
  AOI211_X1 U13766 ( .C1(n11144), .C2(n11143), .A(n6631), .B(n15392), .ZN(
        n11145) );
  INV_X1 U13767 ( .A(n11145), .ZN(n11146) );
  NAND2_X1 U13768 ( .A1(n12187), .A2(n11146), .ZN(n11147) );
  AOI21_X1 U13769 ( .B1(n15373), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n11147), 
        .ZN(n11148) );
  OAI211_X1 U13770 ( .C1(n15408), .C2(n11150), .A(n11149), .B(n11148), .ZN(
        P2_U3224) );
  OAI222_X1 U13771 ( .A1(P3_U3151), .A2(n11153), .B1(n13719), .B2(n11152), 
        .C1(n13717), .C2(n11151), .ZN(P3_U3276) );
  XNOR2_X1 U13772 ( .A(n11154), .B(n11159), .ZN(n15572) );
  INV_X1 U13773 ( .A(n15572), .ZN(n11167) );
  INV_X1 U13774 ( .A(n15538), .ZN(n11155) );
  OAI22_X1 U13775 ( .A1(n11156), .A2(n15508), .B1(n11254), .B2(n15510), .ZN(
        n11161) );
  OR2_X1 U13776 ( .A1(n11157), .A2(n11159), .ZN(n11332) );
  INV_X1 U13777 ( .A(n11332), .ZN(n11158) );
  AOI211_X1 U13778 ( .C1(n11159), .C2(n11157), .A(n13472), .B(n11158), .ZN(
        n11160) );
  AOI211_X1 U13779 ( .C1(n15572), .C2(n13435), .A(n11161), .B(n11160), .ZN(
        n15569) );
  MUX2_X1 U13780 ( .A(n11162), .B(n15569), .S(n15559), .Z(n11166) );
  INV_X1 U13781 ( .A(n11782), .ZN(n15519) );
  NOR2_X1 U13782 ( .A1(n15541), .A2(n11163), .ZN(n15571) );
  AOI22_X1 U13783 ( .A1(n15519), .A2(n15571), .B1(n15518), .B2(n11164), .ZN(
        n11165) );
  OAI211_X1 U13784 ( .C1(n11167), .C2(n15555), .A(n11166), .B(n11165), .ZN(
        P3_U3230) );
  NAND2_X1 U13785 ( .A1(n13865), .A2(n13802), .ZN(n11168) );
  AND2_X1 U13786 ( .A1(n11169), .A2(n11168), .ZN(n15465) );
  OAI22_X1 U13787 ( .A1(n6438), .A2(n15465), .B1(n11170), .B2(n15434), .ZN(
        n11175) );
  OAI211_X1 U13788 ( .C1(n11173), .C2(n15466), .A(n15443), .B(n11172), .ZN(
        n15464) );
  OAI22_X1 U13789 ( .A1(n15466), .A2(n15437), .B1(n14089), .B2(n15464), .ZN(
        n11174) );
  AOI211_X1 U13790 ( .C1(P2_REG2_REG_1__SCAN_IN), .C2(n6438), .A(n11175), .B(
        n11174), .ZN(n11179) );
  XNOR2_X1 U13791 ( .A(n11176), .B(n10694), .ZN(n15463) );
  OR2_X1 U13792 ( .A1(n6438), .A2(n14072), .ZN(n11177) );
  OR2_X1 U13793 ( .A1(n6438), .A2(n14186), .ZN(n14070) );
  XNOR2_X1 U13794 ( .A(n10694), .B(n12663), .ZN(n15469) );
  AOI22_X1 U13795 ( .A1(n15463), .A2(n15446), .B1(n14054), .B2(n15469), .ZN(
        n11178) );
  NAND2_X1 U13796 ( .A1(n11179), .A2(n11178), .ZN(P2_U3264) );
  XNOR2_X1 U13797 ( .A(n13071), .B(n11187), .ZN(n11371) );
  XNOR2_X1 U13798 ( .A(n11371), .B(n13212), .ZN(n11183) );
  NAND2_X1 U13799 ( .A1(n11182), .A2(n11183), .ZN(n11490) );
  OAI21_X1 U13800 ( .B1(n11183), .B2(n11182), .A(n11490), .ZN(n11184) );
  NAND2_X1 U13801 ( .A1(n11184), .A2(n13169), .ZN(n11189) );
  INV_X1 U13802 ( .A(n13211), .ZN(n11541) );
  OAI22_X1 U13803 ( .A1(n13151), .A2(n11254), .B1(n11541), .B2(n13193), .ZN(
        n11185) );
  AOI211_X1 U13804 ( .C1(n13196), .C2(n11187), .A(n11186), .B(n11185), .ZN(
        n11188) );
  OAI211_X1 U13805 ( .C1(n11260), .C2(n13184), .A(n11189), .B(n11188), .ZN(
        P3_U3167) );
  XNOR2_X1 U13806 ( .A(n11190), .B(n12873), .ZN(n15476) );
  OR2_X1 U13807 ( .A1(n13814), .A2(n11191), .ZN(n11193) );
  NAND2_X1 U13808 ( .A1(n13865), .A2(n13801), .ZN(n11192) );
  NAND2_X1 U13809 ( .A1(n11193), .A2(n11192), .ZN(n15470) );
  INV_X1 U13810 ( .A(n15470), .ZN(n15324) );
  INV_X1 U13811 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15323) );
  OAI22_X1 U13812 ( .A1(n6438), .A2(n15324), .B1(n15434), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n11199) );
  NAND2_X1 U13813 ( .A1(n11194), .A2(n15471), .ZN(n11195) );
  NAND2_X1 U13814 ( .A1(n11195), .A2(n15443), .ZN(n11196) );
  OR2_X1 U13815 ( .A1(n11196), .A2(n15441), .ZN(n15473) );
  OAI22_X1 U13816 ( .A1(n11197), .A2(n15437), .B1(n14089), .B2(n15473), .ZN(
        n11198) );
  AOI211_X1 U13817 ( .C1(n6438), .C2(P2_REG2_REG_3__SCAN_IN), .A(n11199), .B(
        n11198), .ZN(n11202) );
  XNOR2_X1 U13818 ( .A(n11200), .B(n12873), .ZN(n15478) );
  NAND2_X1 U13819 ( .A1(n14054), .A2(n15478), .ZN(n11201) );
  OAI211_X1 U13820 ( .C1(n14056), .C2(n15476), .A(n11202), .B(n11201), .ZN(
        P2_U3262) );
  XOR2_X1 U13821 ( .A(n11204), .B(n11203), .Z(n11209) );
  INV_X1 U13822 ( .A(n11205), .ZN(n11207) );
  OAI22_X1 U13823 ( .A1(n15465), .A2(n15325), .B1(n13820), .B2(n15466), .ZN(
        n11206) );
  AOI21_X1 U13824 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n11207), .A(n11206), .ZN(
        n11208) );
  OAI21_X1 U13825 ( .B1(n11209), .B2(n15327), .A(n11208), .ZN(P2_U3194) );
  MUX2_X1 U13826 ( .A(n11210), .B(P1_REG2_REG_5__SCAN_IN), .S(n15307), .Z(
        n11211) );
  INV_X1 U13827 ( .A(n11211), .ZN(n11215) );
  AOI22_X1 U13828 ( .A1(n14980), .A2(n11213), .B1(n15301), .B2(n11212), .ZN(
        n11214) );
  OAI211_X1 U13829 ( .C1(n14984), .C2(n11216), .A(n11215), .B(n11214), .ZN(
        P1_U3288) );
  OAI22_X1 U13830 ( .A1(n11291), .A2(n14413), .B1(n11220), .B2(n14411), .ZN(
        n11474) );
  NAND2_X1 U13831 ( .A1(n11429), .A2(n14346), .ZN(n11222) );
  NAND2_X1 U13832 ( .A1(n14581), .A2(n14295), .ZN(n11221) );
  NAND2_X1 U13833 ( .A1(n11222), .A2(n11221), .ZN(n11223) );
  XNOR2_X1 U13834 ( .A(n11223), .B(n14359), .ZN(n11473) );
  XOR2_X1 U13835 ( .A(n11474), .B(n11473), .Z(n11475) );
  XNOR2_X1 U13836 ( .A(n11476), .B(n11475), .ZN(n11229) );
  NAND2_X1 U13837 ( .A1(n14377), .A2(n14582), .ZN(n11224) );
  OAI21_X1 U13838 ( .B1(n14556), .B2(n11427), .A(n11224), .ZN(n11226) );
  NAND2_X1 U13839 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14643) );
  OAI21_X1 U13840 ( .B1(n14555), .B2(n11667), .A(n14643), .ZN(n11225) );
  NOR2_X1 U13841 ( .A1(n11226), .A2(n11225), .ZN(n11228) );
  NAND2_X1 U13842 ( .A1(n10393), .A2(n11429), .ZN(n11227) );
  OAI211_X1 U13843 ( .C1(n11229), .C2(n14561), .A(n11228), .B(n11227), .ZN(
        P1_U3239) );
  MUX2_X1 U13844 ( .A(n12923), .B(P2_REG2_REG_5__SCAN_IN), .S(n6438), .Z(
        n11231) );
  OAI22_X1 U13845 ( .A1(n15437), .A2(n6876), .B1(n12926), .B2(n15434), .ZN(
        n11230) );
  AOI211_X1 U13846 ( .C1(n11232), .C2(n15445), .A(n11231), .B(n11230), .ZN(
        n11235) );
  NAND2_X1 U13847 ( .A1(n14054), .A2(n11233), .ZN(n11234) );
  OAI211_X1 U13848 ( .C1(n14056), .C2(n11236), .A(n11235), .B(n11234), .ZN(
        P2_U3260) );
  NAND2_X1 U13849 ( .A1(n11237), .A2(n12875), .ZN(n11342) );
  OR2_X1 U13850 ( .A1(n11237), .A2(n12875), .ZN(n11238) );
  NAND2_X1 U13851 ( .A1(n11342), .A2(n11238), .ZN(n15494) );
  INV_X1 U13852 ( .A(n15494), .ZN(n11251) );
  NAND2_X1 U13853 ( .A1(n11239), .A2(n12875), .ZN(n11240) );
  NAND2_X1 U13854 ( .A1(n11241), .A2(n11240), .ZN(n11244) );
  NAND2_X1 U13855 ( .A1(n13860), .A2(n13802), .ZN(n11243) );
  NAND2_X1 U13856 ( .A1(n13862), .A2(n13801), .ZN(n11242) );
  NAND2_X1 U13857 ( .A1(n11243), .A2(n11242), .ZN(n11549) );
  AOI21_X1 U13858 ( .B1(n11244), .B2(n15479), .A(n11549), .ZN(n11246) );
  NAND2_X1 U13859 ( .A1(n15494), .A2(n11872), .ZN(n11245) );
  NAND2_X1 U13860 ( .A1(n11246), .A2(n11245), .ZN(n15493) );
  MUX2_X1 U13861 ( .A(n15493), .B(P2_REG2_REG_6__SCAN_IN), .S(n6438), .Z(
        n11247) );
  INV_X1 U13862 ( .A(n11247), .ZN(n11250) );
  AOI211_X1 U13863 ( .C1(n12692), .C2(n6638), .A(n14166), .B(n11344), .ZN(
        n15488) );
  OAI22_X1 U13864 ( .A1(n15437), .A2(n15491), .B1(n11552), .B2(n15434), .ZN(
        n11248) );
  AOI21_X1 U13865 ( .B1(n15488), .B2(n15445), .A(n11248), .ZN(n11249) );
  OAI211_X1 U13866 ( .C1(n11251), .C2(n12149), .A(n11250), .B(n11249), .ZN(
        P2_U3259) );
  XNOR2_X1 U13867 ( .A(n6634), .B(n12547), .ZN(n15577) );
  OAI21_X1 U13868 ( .B1(n11253), .B2(n12547), .A(n11252), .ZN(n11257) );
  OAI22_X1 U13869 ( .A1(n11254), .A2(n15508), .B1(n11541), .B2(n15510), .ZN(
        n11256) );
  NOR2_X1 U13870 ( .A1(n15577), .A2(n15551), .ZN(n11255) );
  AOI211_X1 U13871 ( .C1(n10147), .C2(n11257), .A(n11256), .B(n11255), .ZN(
        n15578) );
  MUX2_X1 U13872 ( .A(n11258), .B(n15578), .S(n15559), .Z(n11263) );
  NOR2_X1 U13873 ( .A1(n15541), .A2(n11259), .ZN(n15580) );
  INV_X1 U13874 ( .A(n11260), .ZN(n11261) );
  AOI22_X1 U13875 ( .A1(n15519), .A2(n15580), .B1(n15518), .B2(n11261), .ZN(
        n11262) );
  OAI211_X1 U13876 ( .C1(n15577), .C2(n15555), .A(n11263), .B(n11262), .ZN(
        P3_U3228) );
  NAND2_X1 U13877 ( .A1(n11268), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11264) );
  NAND2_X1 U13878 ( .A1(n11265), .A2(n11264), .ZN(n11267) );
  MUX2_X1 U13879 ( .A(n11874), .B(P2_REG2_REG_11__SCAN_IN), .S(n11359), .Z(
        n11266) );
  INV_X1 U13880 ( .A(n11363), .ZN(n11361) );
  AOI21_X1 U13881 ( .B1(n11267), .B2(n11266), .A(n11361), .ZN(n11274) );
  XNOR2_X1 U13882 ( .A(n11359), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n11354) );
  XOR2_X1 U13883 ( .A(n11354), .B(n11355), .Z(n11269) );
  NAND2_X1 U13884 ( .A1(n11269), .A2(n15419), .ZN(n11273) );
  NOR2_X1 U13885 ( .A1(n11270), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12266) );
  NOR2_X1 U13886 ( .A1(n15408), .A2(n11352), .ZN(n11271) );
  AOI211_X1 U13887 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n15373), .A(n12266), 
        .B(n11271), .ZN(n11272) );
  OAI211_X1 U13888 ( .C1(n11274), .C2(n12329), .A(n11273), .B(n11272), .ZN(
        P2_U3225) );
  INV_X1 U13889 ( .A(n11098), .ZN(n11275) );
  NOR2_X1 U13890 ( .A1(n11275), .A2(n11276), .ZN(n11713) );
  OR2_X1 U13891 ( .A1(n11713), .A2(n11279), .ZN(n11457) );
  INV_X1 U13892 ( .A(n11276), .ZN(n11277) );
  NAND3_X1 U13893 ( .A1(n11098), .A2(n11277), .A3(n11279), .ZN(n11278) );
  AOI21_X1 U13894 ( .B1(n11457), .B2(n11278), .A(n15314), .ZN(n11287) );
  INV_X1 U13895 ( .A(n11279), .ZN(n11281) );
  NAND3_X1 U13896 ( .A1(n11092), .A2(n11281), .A3(n11280), .ZN(n11282) );
  AOI21_X1 U13897 ( .B1(n11283), .B2(n11282), .A(n14988), .ZN(n11286) );
  OAI22_X1 U13898 ( .A1(n11667), .A2(n14993), .B1(n11284), .B2(n15032), .ZN(
        n11285) );
  NOR3_X1 U13899 ( .A1(n11287), .A2(n11286), .A3(n11285), .ZN(n11425) );
  INV_X1 U13900 ( .A(n11288), .ZN(n11289) );
  OAI211_X1 U13901 ( .C1(n11289), .C2(n11291), .A(n6432), .B(n11465), .ZN(
        n11432) );
  AND2_X1 U13902 ( .A1(n11425), .A2(n11432), .ZN(n11295) );
  INV_X1 U13903 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11290) );
  OAI22_X1 U13904 ( .A1(n15143), .A2(n11291), .B1(n15319), .B2(n11290), .ZN(
        n11292) );
  INV_X1 U13905 ( .A(n11292), .ZN(n11293) );
  OAI21_X1 U13906 ( .B1(n11295), .B2(n15317), .A(n11293), .ZN(P1_U3477) );
  AOI22_X1 U13907 ( .A1(n11749), .A2(n11429), .B1(n15320), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n11294) );
  OAI21_X1 U13908 ( .B1(n11295), .B2(n15320), .A(n11294), .ZN(P1_U3534) );
  XOR2_X1 U13909 ( .A(n11297), .B(n11296), .Z(n11311) );
  OAI21_X1 U13910 ( .B1(n11300), .B2(n11299), .A(n11298), .ZN(n11305) );
  INV_X1 U13911 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11301) );
  NOR2_X1 U13912 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11301), .ZN(n11609) );
  AOI21_X1 U13913 ( .B1(n15503), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11609), 
        .ZN(n11302) );
  OAI21_X1 U13914 ( .B1(n13355), .B2(n11303), .A(n11302), .ZN(n11304) );
  AOI21_X1 U13915 ( .B1(n11305), .B2(n13270), .A(n11304), .ZN(n11310) );
  AND3_X1 U13916 ( .A1(n11413), .A2(n11307), .A3(n11306), .ZN(n11308) );
  OAI21_X1 U13917 ( .B1(n6637), .B2(n11308), .A(n13348), .ZN(n11309) );
  OAI211_X1 U13918 ( .C1(n11311), .C2(n13333), .A(n11310), .B(n11309), .ZN(
        P3_U3192) );
  INV_X1 U13919 ( .A(n11312), .ZN(n15326) );
  NOR3_X1 U13920 ( .A1(n13790), .A2(n11316), .A3(n11313), .ZN(n11314) );
  AOI21_X1 U13921 ( .B1(n15326), .B2(n13822), .A(n11314), .ZN(n11324) );
  INV_X1 U13922 ( .A(n11315), .ZN(n12930) );
  OR2_X1 U13923 ( .A1(n13812), .A2(n11316), .ZN(n11318) );
  NAND2_X1 U13924 ( .A1(n13862), .A2(n13802), .ZN(n11317) );
  NAND2_X1 U13925 ( .A1(n11318), .A2(n11317), .ZN(n15431) );
  AOI22_X1 U13926 ( .A1(n13826), .A2(n15431), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11320) );
  NAND2_X1 U13927 ( .A1(n15332), .A2(n12683), .ZN(n11319) );
  OAI211_X1 U13928 ( .C1(n15334), .C2(n15433), .A(n11320), .B(n11319), .ZN(
        n11321) );
  AOI21_X1 U13929 ( .B1(n12930), .B2(n13822), .A(n11321), .ZN(n11322) );
  OAI21_X1 U13930 ( .B1(n11324), .B2(n11323), .A(n11322), .ZN(P2_U3202) );
  NAND2_X1 U13931 ( .A1(n11325), .A2(n12408), .ZN(n11327) );
  INV_X1 U13932 ( .A(n12551), .ZN(n11326) );
  XNOR2_X1 U13933 ( .A(n11327), .B(n11326), .ZN(n11337) );
  INV_X1 U13934 ( .A(n11337), .ZN(n15576) );
  NAND2_X1 U13935 ( .A1(n13595), .A2(n11328), .ZN(n15573) );
  OAI22_X1 U13936 ( .A1(n11782), .A2(n15573), .B1(n11329), .B2(n15553), .ZN(
        n11339) );
  INV_X1 U13937 ( .A(n11330), .ZN(n11331) );
  NAND2_X1 U13938 ( .A1(n11332), .A2(n11331), .ZN(n11333) );
  XNOR2_X1 U13939 ( .A(n11333), .B(n12551), .ZN(n11334) );
  NAND2_X1 U13940 ( .A1(n11334), .A2(n10147), .ZN(n11336) );
  AOI22_X1 U13941 ( .A1(n15546), .A2(n15532), .B1(n13212), .B2(n15531), .ZN(
        n11335) );
  OAI211_X1 U13942 ( .C1(n11337), .C2(n15551), .A(n11336), .B(n11335), .ZN(
        n15574) );
  MUX2_X1 U13943 ( .A(n15574), .B(P3_REG2_REG_4__SCAN_IN), .S(n15561), .Z(
        n11338) );
  AOI211_X1 U13944 ( .C1(n15576), .C2(n13440), .A(n11339), .B(n11338), .ZN(
        n11340) );
  INV_X1 U13945 ( .A(n11340), .ZN(P3_U3229) );
  INV_X1 U13946 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n11351) );
  NAND2_X1 U13947 ( .A1(n11342), .A2(n11341), .ZN(n11343) );
  XNOR2_X1 U13948 ( .A(n12700), .B(n13860), .ZN(n12876) );
  XNOR2_X1 U13949 ( .A(n11343), .B(n12876), .ZN(n11437) );
  AOI211_X1 U13950 ( .C1(n12700), .C2(n8884), .A(n14166), .B(n11345), .ZN(
        n11440) );
  AOI21_X1 U13951 ( .B1(n15472), .B2(n12700), .A(n11440), .ZN(n11349) );
  XNOR2_X1 U13952 ( .A(n11346), .B(n12876), .ZN(n11348) );
  OAI22_X1 U13953 ( .A1(n11387), .A2(n13812), .B1(n11347), .B2(n13814), .ZN(
        n11391) );
  AOI21_X1 U13954 ( .B1(n11348), .B2(n15479), .A(n11391), .ZN(n11442) );
  OAI211_X1 U13955 ( .C1(n15475), .C2(n11437), .A(n11349), .B(n11442), .ZN(
        n14223) );
  NAND2_X1 U13956 ( .A1(n14223), .A2(n15496), .ZN(n11350) );
  OAI21_X1 U13957 ( .B1(n15496), .B2(n11351), .A(n11350), .ZN(P2_U3451) );
  XNOR2_X1 U13958 ( .A(n12322), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n11357) );
  OAI22_X1 U13959 ( .A1(n11355), .A2(n11354), .B1(n11353), .B2(n11352), .ZN(
        n11356) );
  AOI21_X1 U13960 ( .B1(n11357), .B2(n11356), .A(n15390), .ZN(n11370) );
  INV_X1 U13961 ( .A(n15408), .ZN(n15421) );
  INV_X1 U13962 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n11984) );
  NAND2_X1 U13963 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n12628)
         );
  OAI21_X1 U13964 ( .B1(n15427), .B2(n11984), .A(n12628), .ZN(n11358) );
  AOI21_X1 U13965 ( .B1(n12322), .B2(n15421), .A(n11358), .ZN(n11369) );
  MUX2_X1 U13966 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n12144), .S(n12322), .Z(
        n11364) );
  OR2_X1 U13967 ( .A1(n11359), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11362) );
  INV_X1 U13968 ( .A(n11362), .ZN(n11360) );
  NOR3_X1 U13969 ( .A1(n11361), .A2(n11364), .A3(n11360), .ZN(n11367) );
  NAND2_X1 U13970 ( .A1(n11363), .A2(n11362), .ZN(n11365) );
  NAND2_X1 U13971 ( .A1(n11365), .A2(n11364), .ZN(n12317) );
  INV_X1 U13972 ( .A(n12317), .ZN(n11366) );
  OAI21_X1 U13973 ( .B1(n11367), .B2(n11366), .A(n15423), .ZN(n11368) );
  OAI211_X1 U13974 ( .C1(n11370), .C2(n15392), .A(n11369), .B(n11368), .ZN(
        P2_U3226) );
  INV_X1 U13975 ( .A(n13212), .ZN(n11375) );
  NAND2_X1 U13976 ( .A1(n11371), .A2(n11375), .ZN(n11487) );
  AND2_X1 U13977 ( .A1(n11490), .A2(n11487), .ZN(n11374) );
  XNOR2_X1 U13978 ( .A(n13071), .B(n11372), .ZN(n11492) );
  XOR2_X1 U13979 ( .A(n13211), .B(n11492), .Z(n11373) );
  NAND2_X1 U13980 ( .A1(n11374), .A2(n11373), .ZN(n11538) );
  OAI211_X1 U13981 ( .C1(n11374), .C2(n11373), .A(n11538), .B(n13169), .ZN(
        n11379) );
  OAI22_X1 U13982 ( .A1(n13151), .A2(n11375), .B1(n11491), .B2(n13193), .ZN(
        n11376) );
  AOI211_X1 U13983 ( .C1(n13196), .C2(n11446), .A(n11377), .B(n11376), .ZN(
        n11378) );
  OAI211_X1 U13984 ( .C1(n11447), .C2(n13184), .A(n11379), .B(n11378), .ZN(
        P3_U3179) );
  OAI222_X1 U13985 ( .A1(P1_U3086), .A2(n15297), .B1(n15159), .B2(n11382), 
        .C1(n11380), .C2(n15165), .ZN(P1_U3335) );
  OAI222_X1 U13986 ( .A1(n14247), .A2(n11383), .B1(n13019), .B2(n11382), .C1(
        n11381), .C2(P2_U3088), .ZN(P2_U3307) );
  INV_X1 U13987 ( .A(n11384), .ZN(n11385) );
  AOI21_X1 U13988 ( .B1(n11553), .B2(n11385), .A(n15327), .ZN(n11389) );
  NOR3_X1 U13989 ( .A1(n13790), .A2(n11387), .A3(n11386), .ZN(n11388) );
  OAI21_X1 U13990 ( .B1(n11389), .B2(n11388), .A(n11576), .ZN(n11393) );
  AND2_X1 U13991 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15374) );
  NOR2_X1 U13992 ( .A1(n15334), .A2(n11433), .ZN(n11390) );
  AOI211_X1 U13993 ( .C1(n13826), .C2(n11391), .A(n15374), .B(n11390), .ZN(
        n11392) );
  OAI211_X1 U13994 ( .C1(n11436), .C2(n13820), .A(n11393), .B(n11392), .ZN(
        P2_U3185) );
  NOR2_X1 U13995 ( .A1(n15434), .A2(n11394), .ZN(n11395) );
  AOI21_X1 U13996 ( .B1(n6438), .B2(P2_REG2_REG_2__SCAN_IN), .A(n11395), .ZN(
        n11396) );
  OAI21_X1 U13997 ( .B1(n15437), .B2(n11397), .A(n11396), .ZN(n11400) );
  NOR2_X1 U13998 ( .A1(n14056), .A2(n11398), .ZN(n11399) );
  AOI211_X1 U13999 ( .C1(n11401), .C2(n15445), .A(n11400), .B(n11399), .ZN(
        n11402) );
  OAI21_X1 U14000 ( .B1(n6438), .B2(n11403), .A(n11402), .ZN(P2_U3263) );
  OAI222_X1 U14001 ( .A1(n14247), .A2(n11405), .B1(n13019), .B2(n11407), .C1(
        n11404), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U14002 ( .A1(P1_U3086), .A2(n11408), .B1(n15159), .B2(n11407), 
        .C1(n11406), .C2(n15165), .ZN(P1_U3334) );
  XNOR2_X1 U14003 ( .A(n11409), .B(P3_REG1_REG_9__SCAN_IN), .ZN(n11422) );
  NAND2_X1 U14004 ( .A1(n6641), .A2(n11410), .ZN(n11411) );
  XNOR2_X1 U14005 ( .A(n11412), .B(n11411), .ZN(n11420) );
  OAI21_X1 U14006 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11414), .A(n11413), .ZN(
        n11415) );
  NAND2_X1 U14007 ( .A1(n11415), .A2(n13348), .ZN(n11417) );
  NOR2_X1 U14008 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9076), .ZN(n11504) );
  AOI21_X1 U14009 ( .B1(n15503), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11504), .ZN(
        n11416) );
  OAI211_X1 U14010 ( .C1(n13355), .C2(n11418), .A(n11417), .B(n11416), .ZN(
        n11419) );
  AOI21_X1 U14011 ( .B1(n13270), .B2(n11420), .A(n11419), .ZN(n11421) );
  OAI21_X1 U14012 ( .B1(n11422), .B2(n13333), .A(n11421), .ZN(P3_U3191) );
  INV_X1 U14013 ( .A(n11423), .ZN(n13018) );
  OAI222_X1 U14014 ( .A1(n15165), .A2(n11424), .B1(n15159), .B2(n13018), .C1(
        P1_U3086), .C2(n8398), .ZN(P1_U3336) );
  MUX2_X1 U14015 ( .A(n11426), .B(n11425), .S(n15305), .Z(n11431) );
  INV_X1 U14016 ( .A(n11427), .ZN(n11428) );
  AOI22_X1 U14017 ( .A1(n14980), .A2(n11429), .B1(n15301), .B2(n11428), .ZN(
        n11430) );
  OAI211_X1 U14018 ( .C1(n14984), .C2(n11432), .A(n11431), .B(n11430), .ZN(
        P1_U3287) );
  INV_X1 U14019 ( .A(n11433), .ZN(n11434) );
  INV_X1 U14020 ( .A(n15434), .ZN(n14083) );
  AOI22_X1 U14021 ( .A1(n6438), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n11434), .B2(
        n14083), .ZN(n11435) );
  OAI21_X1 U14022 ( .B1(n15437), .B2(n11436), .A(n11435), .ZN(n11439) );
  NOR2_X1 U14023 ( .A1(n11437), .A2(n14056), .ZN(n11438) );
  AOI211_X1 U14024 ( .C1(n11440), .C2(n15445), .A(n11439), .B(n11438), .ZN(
        n11441) );
  OAI21_X1 U14025 ( .B1(n6438), .B2(n11442), .A(n11441), .ZN(P2_U3258) );
  OR2_X1 U14026 ( .A1(n11444), .A2(n12552), .ZN(n11445) );
  NAND2_X1 U14027 ( .A1(n11443), .A2(n11445), .ZN(n15585) );
  NAND2_X1 U14028 ( .A1(n13595), .A2(n11446), .ZN(n15582) );
  OAI22_X1 U14029 ( .A1(n11782), .A2(n15582), .B1(n11447), .B2(n15553), .ZN(
        n11454) );
  NAND2_X1 U14030 ( .A1(n15585), .A2(n13435), .ZN(n11452) );
  AOI21_X1 U14031 ( .B1(n11448), .B2(n12552), .A(n13472), .ZN(n11449) );
  NAND2_X1 U14032 ( .A1(n11449), .A2(n11676), .ZN(n11451) );
  AOI22_X1 U14033 ( .A1(n15531), .A2(n13210), .B1(n13212), .B2(n15546), .ZN(
        n11450) );
  NAND3_X1 U14034 ( .A1(n11452), .A2(n11451), .A3(n11450), .ZN(n15583) );
  MUX2_X1 U14035 ( .A(n15583), .B(P3_REG2_REG_6__SCAN_IN), .S(n15561), .Z(
        n11453) );
  AOI211_X1 U14036 ( .C1(n13440), .C2(n15585), .A(n11454), .B(n11453), .ZN(
        n11455) );
  INV_X1 U14037 ( .A(n11455), .ZN(P3_U3227) );
  NAND2_X1 U14038 ( .A1(n11457), .A2(n11456), .ZN(n11458) );
  XOR2_X1 U14039 ( .A(n11458), .B(n11459), .Z(n11464) );
  XOR2_X1 U14040 ( .A(n11460), .B(n11459), .Z(n11462) );
  AOI22_X1 U14041 ( .A1(n15010), .A2(n14581), .B1(n14578), .B2(n15008), .ZN(
        n11461) );
  OAI21_X1 U14042 ( .B1(n11462), .B2(n14988), .A(n11461), .ZN(n11463) );
  AOI21_X1 U14043 ( .B1(n11464), .B2(n15078), .A(n11463), .ZN(n11593) );
  NAND2_X1 U14044 ( .A1(n11465), .A2(n11596), .ZN(n11466) );
  NAND2_X1 U14045 ( .A1(n11466), .A2(n6432), .ZN(n11467) );
  OR2_X1 U14046 ( .A1(n11467), .A2(n11716), .ZN(n11599) );
  AND2_X1 U14047 ( .A1(n11593), .A2(n11599), .ZN(n11472) );
  AOI22_X1 U14048 ( .A1(n11749), .A2(n11596), .B1(n15320), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n11468) );
  OAI21_X1 U14049 ( .B1(n11472), .B2(n15320), .A(n11468), .ZN(P1_U3535) );
  INV_X1 U14050 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11469) );
  OAI22_X1 U14051 ( .A1(n7700), .A2(n15143), .B1(n15319), .B2(n11469), .ZN(
        n11470) );
  INV_X1 U14052 ( .A(n11470), .ZN(n11471) );
  OAI21_X1 U14053 ( .B1(n11472), .B2(n15317), .A(n11471), .ZN(P1_U3480) );
  NAND2_X1 U14054 ( .A1(n11596), .A2(n14346), .ZN(n11478) );
  NAND2_X1 U14055 ( .A1(n14579), .A2(n14295), .ZN(n11477) );
  NAND2_X1 U14056 ( .A1(n11478), .A2(n11477), .ZN(n11479) );
  XNOR2_X1 U14057 ( .A(n11479), .B(n14359), .ZN(n11653) );
  OAI22_X1 U14058 ( .A1(n7700), .A2(n14413), .B1(n11667), .B2(n14411), .ZN(
        n11652) );
  XNOR2_X1 U14059 ( .A(n11653), .B(n11652), .ZN(n11656) );
  XNOR2_X1 U14060 ( .A(n11657), .B(n11656), .ZN(n11485) );
  NAND2_X1 U14061 ( .A1(n14377), .A2(n14581), .ZN(n11480) );
  OAI21_X1 U14062 ( .B1(n14556), .B2(n11594), .A(n11480), .ZN(n11482) );
  NAND2_X1 U14063 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14656) );
  OAI21_X1 U14064 ( .B1(n14555), .B2(n12041), .A(n14656), .ZN(n11481) );
  NOR2_X1 U14065 ( .A1(n11482), .A2(n11481), .ZN(n11484) );
  NAND2_X1 U14066 ( .A1(n10393), .A2(n11596), .ZN(n11483) );
  OAI211_X1 U14067 ( .C1(n11485), .C2(n14561), .A(n11484), .B(n11483), .ZN(
        P1_U3213) );
  XNOR2_X1 U14068 ( .A(n13071), .B(n15516), .ZN(n11600) );
  XNOR2_X1 U14069 ( .A(n11600), .B(n13208), .ZN(n11502) );
  XNOR2_X1 U14070 ( .A(n6431), .B(n11486), .ZN(n11493) );
  XNOR2_X1 U14071 ( .A(n11493), .B(n13209), .ZN(n13083) );
  XNOR2_X1 U14072 ( .A(n13210), .B(n11673), .ZN(n12426) );
  OAI211_X1 U14073 ( .C1(n11492), .C2(n13211), .A(n11487), .B(n13081), .ZN(
        n11488) );
  NOR2_X1 U14074 ( .A1(n13083), .A2(n11488), .ZN(n11489) );
  NAND2_X1 U14075 ( .A1(n11490), .A2(n11489), .ZN(n11497) );
  INV_X1 U14076 ( .A(n13081), .ZN(n11539) );
  OAI21_X1 U14077 ( .B1(n13083), .B2(n11491), .A(n11539), .ZN(n11495) );
  NAND2_X1 U14078 ( .A1(n11492), .A2(n13211), .ZN(n11537) );
  OAI21_X1 U14079 ( .B1(n13083), .B2(n11537), .A(n13081), .ZN(n11494) );
  AOI22_X1 U14080 ( .A1(n11495), .A2(n11494), .B1(n11493), .B2(n13209), .ZN(
        n11496) );
  NAND2_X1 U14081 ( .A1(n11497), .A2(n11496), .ZN(n11498) );
  INV_X1 U14082 ( .A(n11498), .ZN(n11500) );
  INV_X1 U14083 ( .A(n11604), .ZN(n11501) );
  AOI21_X1 U14084 ( .B1(n11502), .B2(n11498), .A(n11501), .ZN(n11509) );
  INV_X1 U14085 ( .A(n15516), .ZN(n11505) );
  OAI22_X1 U14086 ( .A1(n13151), .A2(n15509), .B1(n15511), .B2(n13193), .ZN(
        n11503) );
  AOI211_X1 U14087 ( .C1(n13196), .C2(n11505), .A(n11504), .B(n11503), .ZN(
        n11508) );
  INV_X1 U14088 ( .A(n11506), .ZN(n15517) );
  NAND2_X1 U14089 ( .A1(n13195), .A2(n15517), .ZN(n11507) );
  OAI211_X1 U14090 ( .C1(n11509), .C2(n13199), .A(n11508), .B(n11507), .ZN(
        P3_U3171) );
  OAI222_X1 U14091 ( .A1(n14247), .A2(n11511), .B1(P2_U3088), .B2(n12906), 
        .C1(n13019), .C2(n11510), .ZN(P2_U3305) );
  XNOR2_X1 U14092 ( .A(n14698), .B(n11512), .ZN(n14690) );
  NAND2_X1 U14093 ( .A1(n11520), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n14691) );
  AND2_X1 U14094 ( .A1(n14690), .A2(n14691), .ZN(n11513) );
  NAND2_X1 U14095 ( .A1(n14692), .A2(n11513), .ZN(n14689) );
  OAI21_X1 U14096 ( .B1(n14698), .B2(P1_REG1_REG_14__SCAN_IN), .A(n14689), 
        .ZN(n11514) );
  XOR2_X1 U14097 ( .A(n11525), .B(n11514), .Z(n11645) );
  NOR2_X1 U14098 ( .A1(n11645), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11644) );
  INV_X1 U14099 ( .A(n11514), .ZN(n11515) );
  NOR2_X1 U14100 ( .A1(n11515), .A2(n11525), .ZN(n11517) );
  XNOR2_X1 U14101 ( .A(n12087), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11516) );
  INV_X1 U14102 ( .A(n12086), .ZN(n11519) );
  OAI21_X1 U14103 ( .B1(n11644), .B2(n11517), .A(n11516), .ZN(n11518) );
  NAND3_X1 U14104 ( .A1(n11519), .A2(n14739), .A3(n11518), .ZN(n11535) );
  NAND2_X1 U14105 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14468)
         );
  XNOR2_X1 U14106 ( .A(n12087), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n11529) );
  NAND2_X1 U14107 ( .A1(n11520), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n14700) );
  NAND2_X1 U14108 ( .A1(n14701), .A2(n14700), .ZN(n11523) );
  MUX2_X1 U14109 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11521), .S(n14698), .Z(
        n11522) );
  NAND2_X1 U14110 ( .A1(n11523), .A2(n11522), .ZN(n14703) );
  NAND2_X1 U14111 ( .A1(n14698), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14112 ( .A1(n14703), .A2(n11524), .ZN(n11526) );
  XNOR2_X1 U14113 ( .A(n11526), .B(n11643), .ZN(n11641) );
  INV_X1 U14114 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15002) );
  NAND2_X1 U14115 ( .A1(n11641), .A2(n15002), .ZN(n11528) );
  OR2_X1 U14116 ( .A1(n11526), .A2(n11525), .ZN(n11527) );
  NAND2_X1 U14117 ( .A1(n11528), .A2(n11527), .ZN(n11530) );
  AOI21_X1 U14118 ( .B1(n11529), .B2(n11530), .A(n14735), .ZN(n11531) );
  NAND2_X1 U14119 ( .A1(n11531), .A2(n12084), .ZN(n11532) );
  NAND2_X1 U14120 ( .A1(n14468), .A2(n11532), .ZN(n11533) );
  AOI21_X1 U14121 ( .B1(n15269), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11533), 
        .ZN(n11534) );
  OAI211_X1 U14122 ( .C1(n14719), .C2(n11536), .A(n11535), .B(n11534), .ZN(
        P1_U3259) );
  NAND2_X1 U14123 ( .A1(n11538), .A2(n11537), .ZN(n13082) );
  XNOR2_X1 U14124 ( .A(n13082), .B(n11539), .ZN(n11540) );
  NAND2_X1 U14125 ( .A1(n11540), .A2(n13169), .ZN(n11545) );
  OAI22_X1 U14126 ( .A1(n13151), .A2(n11541), .B1(n15509), .B2(n13193), .ZN(
        n11542) );
  AOI211_X1 U14127 ( .C1(n13196), .C2(n11673), .A(n11543), .B(n11542), .ZN(
        n11544) );
  OAI211_X1 U14128 ( .C1(n11674), .C2(n13184), .A(n11545), .B(n11544), .ZN(
        P3_U3153) );
  INV_X1 U14129 ( .A(n11546), .ZN(n11548) );
  OAI22_X1 U14130 ( .A1(n12582), .A2(P3_U3151), .B1(SI_22_), .B2(n13719), .ZN(
        n11547) );
  AOI21_X1 U14131 ( .B1(n11548), .B2(n13702), .A(n11547), .ZN(P3_U3273) );
  NAND2_X1 U14132 ( .A1(n13826), .A2(n11549), .ZN(n11550) );
  OAI211_X1 U14133 ( .C1(n15334), .C2(n11552), .A(n11551), .B(n11550), .ZN(
        n11558) );
  INV_X1 U14134 ( .A(n11553), .ZN(n11554) );
  AOI211_X1 U14135 ( .C1(n11556), .C2(n11555), .A(n15327), .B(n11554), .ZN(
        n11557) );
  AOI211_X1 U14136 ( .C1(n12692), .C2(n15332), .A(n11558), .B(n11557), .ZN(
        n11559) );
  INV_X1 U14137 ( .A(n11559), .ZN(P2_U3211) );
  NAND2_X1 U14138 ( .A1(n11561), .A2(n12878), .ZN(n11562) );
  INV_X1 U14139 ( .A(n11565), .ZN(n14221) );
  OR2_X1 U14140 ( .A1(n13814), .A2(n11761), .ZN(n11564) );
  NAND2_X1 U14141 ( .A1(n13860), .A2(n13801), .ZN(n11563) );
  NAND2_X1 U14142 ( .A1(n11564), .A2(n11563), .ZN(n11583) );
  AOI21_X1 U14143 ( .B1(n11565), .B2(n11872), .A(n11583), .ZN(n11569) );
  XNOR2_X1 U14144 ( .A(n11566), .B(n12878), .ZN(n11567) );
  NAND2_X1 U14145 ( .A1(n11567), .A2(n15479), .ZN(n11568) );
  NAND2_X1 U14146 ( .A1(n11569), .A2(n11568), .ZN(n14218) );
  MUX2_X1 U14147 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n14218), .S(n14064), .Z(
        n11570) );
  INV_X1 U14148 ( .A(n11570), .ZN(n11575) );
  INV_X1 U14149 ( .A(n11345), .ZN(n11572) );
  INV_X1 U14150 ( .A(n11697), .ZN(n11571) );
  AOI211_X1 U14151 ( .C1(n14217), .C2(n11572), .A(n14166), .B(n11571), .ZN(
        n14216) );
  OAI22_X1 U14152 ( .A1(n15437), .A2(n11582), .B1(n11586), .B2(n15434), .ZN(
        n11573) );
  AOI21_X1 U14153 ( .B1(n14216), .B2(n15445), .A(n11573), .ZN(n11574) );
  OAI211_X1 U14154 ( .C1(n14221), .C2(n12149), .A(n11575), .B(n11574), .ZN(
        P2_U3257) );
  INV_X1 U14155 ( .A(n11576), .ZN(n11580) );
  NOR3_X1 U14156 ( .A1(n13790), .A2(n11578), .A3(n11577), .ZN(n11579) );
  AOI21_X1 U14157 ( .B1(n11580), .B2(n13822), .A(n11579), .ZN(n11591) );
  INV_X1 U14158 ( .A(n11581), .ZN(n12592) );
  NOR2_X1 U14159 ( .A1(n13820), .A2(n11582), .ZN(n11588) );
  NAND2_X1 U14160 ( .A1(n13826), .A2(n11583), .ZN(n11584) );
  OAI211_X1 U14161 ( .C1(n15334), .C2(n11586), .A(n11585), .B(n11584), .ZN(
        n11587) );
  AOI211_X1 U14162 ( .C1(n12592), .C2(n13822), .A(n11588), .B(n11587), .ZN(
        n11589) );
  OAI21_X1 U14163 ( .B1(n11591), .B2(n11590), .A(n11589), .ZN(P2_U3193) );
  MUX2_X1 U14164 ( .A(n11593), .B(n11592), .S(n15307), .Z(n11598) );
  INV_X1 U14165 ( .A(n11594), .ZN(n11595) );
  AOI22_X1 U14166 ( .A1(n14980), .A2(n11596), .B1(n11595), .B2(n15301), .ZN(
        n11597) );
  OAI211_X1 U14167 ( .C1(n14984), .C2(n11599), .A(n11598), .B(n11597), .ZN(
        P1_U3286) );
  INV_X1 U14168 ( .A(n11600), .ZN(n11601) );
  NAND2_X1 U14169 ( .A1(n11601), .A2(n11607), .ZN(n11602) );
  AND2_X1 U14170 ( .A1(n11604), .A2(n11602), .ZN(n11606) );
  XNOR2_X1 U14171 ( .A(n13071), .B(n12064), .ZN(n12018) );
  XNOR2_X1 U14172 ( .A(n12018), .B(n15511), .ZN(n11605) );
  AND2_X1 U14173 ( .A1(n11605), .A2(n11602), .ZN(n11603) );
  OAI211_X1 U14174 ( .C1(n11606), .C2(n11605), .A(n13169), .B(n12020), .ZN(
        n11611) );
  INV_X1 U14175 ( .A(n12064), .ZN(n11693) );
  OAI22_X1 U14176 ( .A1(n13151), .A2(n11607), .B1(n13157), .B2(n13193), .ZN(
        n11608) );
  AOI211_X1 U14177 ( .C1(n13196), .C2(n11693), .A(n11609), .B(n11608), .ZN(
        n11610) );
  OAI211_X1 U14178 ( .C1(n12055), .C2(n13184), .A(n11611), .B(n11610), .ZN(
        P3_U3157) );
  INV_X1 U14179 ( .A(n11613), .ZN(n11614) );
  XNOR2_X1 U14180 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), 
        .ZN(n11623) );
  XNOR2_X1 U14181 ( .A(n11622), .B(n11623), .ZN(n11618) );
  NAND2_X1 U14182 ( .A1(n15174), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11621) );
  INV_X1 U14183 ( .A(n11617), .ZN(n11619) );
  NAND2_X1 U14184 ( .A1(n11619), .A2(n11618), .ZN(n11620) );
  INV_X1 U14185 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U14186 ( .A1(n11623), .A2(n11622), .ZN(n11624) );
  XNOR2_X1 U14187 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n11626) );
  XNOR2_X1 U14188 ( .A(n11850), .B(n11626), .ZN(n11628) );
  INV_X1 U14189 ( .A(n11848), .ZN(n11633) );
  INV_X1 U14190 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n11629) );
  INV_X1 U14191 ( .A(n11630), .ZN(n11631) );
  OAI21_X1 U14192 ( .B1(n11633), .B2(n11631), .A(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n11632) );
  OAI21_X1 U14193 ( .B1(n11633), .B2(n11849), .A(n11632), .ZN(SUB_1596_U70) );
  NAND2_X1 U14194 ( .A1(n11634), .A2(n13702), .ZN(n11635) );
  OAI211_X1 U14195 ( .C1(n11636), .C2(n13719), .A(n11635), .B(n12584), .ZN(
        P3_U3272) );
  INV_X1 U14196 ( .A(n11637), .ZN(n11638) );
  OAI222_X1 U14197 ( .A1(P3_U3151), .A2(n11640), .B1(n13719), .B2(n11639), 
        .C1(n13717), .C2(n11638), .ZN(P3_U3275) );
  XNOR2_X1 U14198 ( .A(n11641), .B(n15002), .ZN(n11650) );
  NAND2_X1 U14199 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14554)
         );
  NAND2_X1 U14200 ( .A1(n15269), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n11642) );
  OAI211_X1 U14201 ( .C1(n14719), .C2(n11643), .A(n14554), .B(n11642), .ZN(
        n11649) );
  AOI21_X1 U14202 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n11645), .A(n11644), 
        .ZN(n11647) );
  NOR2_X1 U14203 ( .A1(n11647), .A2(n11646), .ZN(n11648) );
  AOI211_X1 U14204 ( .C1(n14733), .C2(n11650), .A(n11649), .B(n11648), .ZN(
        n11651) );
  INV_X1 U14205 ( .A(n11651), .ZN(P1_U3258) );
  INV_X1 U14206 ( .A(n11652), .ZN(n11655) );
  INV_X1 U14207 ( .A(n11653), .ZN(n11654) );
  NAND2_X1 U14208 ( .A1(n11723), .A2(n14346), .ZN(n11659) );
  NAND2_X1 U14209 ( .A1(n14578), .A2(n14295), .ZN(n11658) );
  NAND2_X1 U14210 ( .A1(n11659), .A2(n11658), .ZN(n11661) );
  XNOR2_X1 U14211 ( .A(n11661), .B(n11660), .ZN(n11664) );
  AND2_X1 U14212 ( .A1(n14578), .A2(n10794), .ZN(n11662) );
  AOI21_X1 U14213 ( .B1(n11723), .B2(n14295), .A(n11662), .ZN(n11663) );
  NAND2_X1 U14214 ( .A1(n11664), .A2(n11663), .ZN(n12034) );
  OAI21_X1 U14215 ( .B1(n11664), .B2(n11663), .A(n12034), .ZN(n11665) );
  AOI21_X1 U14216 ( .B1(n11666), .B2(n11665), .A(n6628), .ZN(n11672) );
  OAI22_X1 U14217 ( .A1(n11667), .A2(n15032), .B1(n12167), .B2(n14993), .ZN(
        n11720) );
  NAND2_X1 U14218 ( .A1(n11720), .A2(n14547), .ZN(n11669) );
  OAI211_X1 U14219 ( .C1(n14556), .C2(n15275), .A(n11669), .B(n11668), .ZN(
        n11670) );
  AOI21_X1 U14220 ( .B1(n11723), .B2(n10393), .A(n11670), .ZN(n11671) );
  OAI21_X1 U14221 ( .B1(n11672), .B2(n14561), .A(n11671), .ZN(P1_U3221) );
  NAND2_X1 U14222 ( .A1(n11443), .A2(n12425), .ZN(n11777) );
  XNOR2_X1 U14223 ( .A(n11777), .B(n12426), .ZN(n15589) );
  NAND2_X1 U14224 ( .A1(n11673), .A2(n13595), .ZN(n15586) );
  OAI22_X1 U14225 ( .A1(n11782), .A2(n15586), .B1(n11674), .B2(n15553), .ZN(
        n11682) );
  NAND2_X1 U14226 ( .A1(n15589), .A2(n13435), .ZN(n11680) );
  AOI22_X1 U14227 ( .A1(n13209), .A2(n15543), .B1(n15546), .B2(n13211), .ZN(
        n11679) );
  NAND2_X1 U14228 ( .A1(n11676), .A2(n11675), .ZN(n11677) );
  INV_X1 U14229 ( .A(n12426), .ZN(n12553) );
  NAND2_X1 U14230 ( .A1(n11677), .A2(n12553), .ZN(n11784) );
  OAI211_X1 U14231 ( .C1(n11677), .C2(n12553), .A(n11784), .B(n10147), .ZN(
        n11678) );
  NAND3_X1 U14232 ( .A1(n11680), .A2(n11679), .A3(n11678), .ZN(n15587) );
  MUX2_X1 U14233 ( .A(n15587), .B(P3_REG2_REG_7__SCAN_IN), .S(n15561), .Z(
        n11681) );
  AOI211_X1 U14234 ( .C1(n15589), .C2(n13440), .A(n11682), .B(n11681), .ZN(
        n11683) );
  INV_X1 U14235 ( .A(n11683), .ZN(P3_U3226) );
  INV_X1 U14236 ( .A(n11684), .ZN(n11685) );
  OAI222_X1 U14237 ( .A1(P3_U3151), .A2(n12392), .B1(n13719), .B2(n11686), 
        .C1(n13717), .C2(n11685), .ZN(P3_U3274) );
  XNOR2_X1 U14238 ( .A(n11687), .B(n11689), .ZN(n12059) );
  XNOR2_X1 U14239 ( .A(n11688), .B(n11689), .ZN(n11692) );
  NAND2_X1 U14240 ( .A1(n12059), .A2(n13435), .ZN(n11691) );
  AOI22_X1 U14241 ( .A1(n12448), .A2(n15531), .B1(n15546), .B2(n13208), .ZN(
        n11690) );
  OAI211_X1 U14242 ( .C1(n11692), .C2(n13472), .A(n11691), .B(n11690), .ZN(
        n12056) );
  AOI21_X1 U14243 ( .B1(n15596), .B2(n12059), .A(n12056), .ZN(n12061) );
  AOI22_X1 U14244 ( .A1(n13691), .A2(n11693), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n15598), .ZN(n11694) );
  OAI21_X1 U14245 ( .B1(n12061), .B2(n15598), .A(n11694), .ZN(P3_U3420) );
  INV_X1 U14246 ( .A(n14222), .ZN(n15495) );
  XNOR2_X1 U14247 ( .A(n11696), .B(n11695), .ZN(n11830) );
  INV_X1 U14248 ( .A(n12706), .ZN(n11700) );
  AOI21_X1 U14249 ( .B1(n11697), .B2(n12706), .A(n14166), .ZN(n11699) );
  NAND2_X1 U14250 ( .A1(n11699), .A2(n11757), .ZN(n11826) );
  OAI21_X1 U14251 ( .B1(n11700), .B2(n15490), .A(n11826), .ZN(n11707) );
  XNOR2_X1 U14252 ( .A(n11701), .B(n12880), .ZN(n11702) );
  NAND2_X1 U14253 ( .A1(n11702), .A2(n15479), .ZN(n11706) );
  OR2_X1 U14254 ( .A1(n13814), .A2(n12262), .ZN(n11704) );
  NAND2_X1 U14255 ( .A1(n13859), .A2(n13801), .ZN(n11703) );
  NAND2_X1 U14256 ( .A1(n11704), .A2(n11703), .ZN(n12586) );
  AOI21_X1 U14257 ( .B1(n11830), .B2(n11872), .A(n12586), .ZN(n11705) );
  NAND2_X1 U14258 ( .A1(n11706), .A2(n11705), .ZN(n11827) );
  AOI211_X1 U14259 ( .C1(n15495), .C2(n11830), .A(n11707), .B(n11827), .ZN(
        n11880) );
  NAND2_X1 U14260 ( .A1(n15500), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11708) );
  OAI21_X1 U14261 ( .B1(n11880), .B2(n15500), .A(n11708), .ZN(P2_U3508) );
  INV_X1 U14262 ( .A(n11709), .ZN(n11712) );
  INV_X1 U14263 ( .A(n11710), .ZN(n11711) );
  OAI21_X1 U14264 ( .B1(n11713), .B2(n11712), .A(n11711), .ZN(n11715) );
  OAI21_X1 U14265 ( .B1(n11715), .B2(n11719), .A(n11714), .ZN(n15283) );
  XNOR2_X1 U14266 ( .A(n11716), .B(n15280), .ZN(n11717) );
  NOR2_X1 U14267 ( .A1(n11717), .A2(n15015), .ZN(n15274) );
  XOR2_X1 U14268 ( .A(n11719), .B(n11718), .Z(n11721) );
  AOI21_X1 U14269 ( .B1(n11721), .B2(n14874), .A(n11720), .ZN(n15285) );
  INV_X1 U14270 ( .A(n15285), .ZN(n11722) );
  AOI211_X1 U14271 ( .C1(n15078), .C2(n15283), .A(n15274), .B(n11722), .ZN(
        n11728) );
  AOI22_X1 U14272 ( .A1(n11749), .A2(n11723), .B1(n15320), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n11724) );
  OAI21_X1 U14273 ( .B1(n11728), .B2(n15320), .A(n11724), .ZN(P1_U3536) );
  INV_X1 U14274 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11725) );
  OAI22_X1 U14275 ( .A1(n15280), .A2(n15143), .B1(n15319), .B2(n11725), .ZN(
        n11726) );
  INV_X1 U14276 ( .A(n11726), .ZN(n11727) );
  OAI21_X1 U14277 ( .B1(n11728), .B2(n15317), .A(n11727), .ZN(P1_U3483) );
  NAND2_X1 U14278 ( .A1(n11733), .A2(n11729), .ZN(n11731) );
  NOR2_X1 U14279 ( .A1(n11730), .A2(P2_U3088), .ZN(n12907) );
  INV_X1 U14280 ( .A(n12907), .ZN(n12917) );
  OAI211_X1 U14281 ( .C1(n11732), .C2(n14247), .A(n11731), .B(n12917), .ZN(
        P2_U3304) );
  NAND2_X1 U14282 ( .A1(n11733), .A2(n15161), .ZN(n11735) );
  OAI211_X1 U14283 ( .C1(n11736), .C2(n15165), .A(n11735), .B(n11734), .ZN(
        P1_U3332) );
  INV_X1 U14284 ( .A(n11738), .ZN(n11739) );
  OAI21_X1 U14285 ( .B1(n11739), .B2(n11741), .A(n12067), .ZN(n11746) );
  NAND3_X1 U14286 ( .A1(n11714), .A2(n11741), .A3(n11740), .ZN(n11742) );
  AOI21_X1 U14287 ( .B1(n6925), .B2(n11742), .A(n15314), .ZN(n11745) );
  OAI22_X1 U14288 ( .A1(n12041), .A2(n15032), .B1(n14521), .B2(n14993), .ZN(
        n11744) );
  AOI211_X1 U14289 ( .C1(n11746), .C2(n14874), .A(n11745), .B(n11744), .ZN(
        n11772) );
  OAI211_X1 U14290 ( .C1(n11748), .C2(n11747), .A(n6432), .B(n12102), .ZN(
        n11776) );
  AND2_X1 U14291 ( .A1(n11772), .A2(n11776), .ZN(n11753) );
  AOI22_X1 U14292 ( .A1(n12044), .A2(n11749), .B1(P1_REG1_REG_9__SCAN_IN), 
        .B2(n15320), .ZN(n11750) );
  OAI21_X1 U14293 ( .B1(n11753), .B2(n15320), .A(n11750), .ZN(P1_U3537) );
  INV_X1 U14294 ( .A(n15143), .ZN(n11751) );
  AOI22_X1 U14295 ( .A1(n12044), .A2(n11751), .B1(P1_REG0_REG_9__SCAN_IN), 
        .B2(n15317), .ZN(n11752) );
  OAI21_X1 U14296 ( .B1(n11753), .B2(n15317), .A(n11752), .ZN(P1_U3486) );
  NAND2_X1 U14297 ( .A1(n11755), .A2(n11754), .ZN(n11756) );
  XNOR2_X1 U14298 ( .A(n11756), .B(n11760), .ZN(n12053) );
  AOI21_X1 U14299 ( .B1(n11757), .B2(n12711), .A(n14166), .ZN(n11758) );
  NAND2_X1 U14300 ( .A1(n11758), .A2(n11873), .ZN(n12049) );
  OAI21_X1 U14301 ( .B1(n8885), .B2(n15490), .A(n12049), .ZN(n11766) );
  XNOR2_X1 U14302 ( .A(n11759), .B(n11760), .ZN(n11765) );
  OR2_X1 U14303 ( .A1(n13812), .A2(n11761), .ZN(n11763) );
  NAND2_X1 U14304 ( .A1(n13855), .A2(n13802), .ZN(n11762) );
  NAND2_X1 U14305 ( .A1(n11763), .A2(n11762), .ZN(n12185) );
  AOI21_X1 U14306 ( .B1(n12053), .B2(n11872), .A(n12185), .ZN(n11764) );
  OAI21_X1 U14307 ( .B1(n11765), .B2(n14186), .A(n11764), .ZN(n12050) );
  AOI211_X1 U14308 ( .C1(n15495), .C2(n12053), .A(n11766), .B(n12050), .ZN(
        n11769) );
  NAND2_X1 U14309 ( .A1(n6954), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n11767) );
  OAI21_X1 U14310 ( .B1(n11769), .B2(n6954), .A(n11767), .ZN(P2_U3460) );
  NAND2_X1 U14311 ( .A1(n15500), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11768) );
  OAI21_X1 U14312 ( .B1(n11769), .B2(n15500), .A(n11768), .ZN(P2_U3509) );
  NAND2_X1 U14313 ( .A1(n13214), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11770) );
  OAI21_X1 U14314 ( .B1(n13214), .B2(n13077), .A(n11770), .ZN(P3_U3520) );
  MUX2_X1 U14315 ( .A(n11772), .B(n11771), .S(n15307), .Z(n11775) );
  INV_X1 U14316 ( .A(n12040), .ZN(n11773) );
  AOI22_X1 U14317 ( .A1(n12044), .A2(n14980), .B1(n15301), .B2(n11773), .ZN(
        n11774) );
  OAI211_X1 U14318 ( .C1(n14984), .C2(n11776), .A(n11775), .B(n11774), .ZN(
        P1_U3284) );
  NAND2_X1 U14319 ( .A1(n11777), .A2(n12426), .ZN(n11779) );
  NAND2_X1 U14320 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  XNOR2_X1 U14321 ( .A(n11780), .B(n11785), .ZN(n15593) );
  NAND2_X1 U14322 ( .A1(n13087), .A2(n13595), .ZN(n15590) );
  OAI22_X1 U14323 ( .A1(n11782), .A2(n15590), .B1(n11781), .B2(n15553), .ZN(
        n11792) );
  NAND2_X1 U14324 ( .A1(n11784), .A2(n11783), .ZN(n11786) );
  XNOR2_X1 U14325 ( .A(n11786), .B(n11785), .ZN(n11787) );
  NAND2_X1 U14326 ( .A1(n11787), .A2(n10147), .ZN(n11790) );
  NAND2_X1 U14327 ( .A1(n15593), .A2(n13435), .ZN(n11789) );
  AOI22_X1 U14328 ( .A1(n15546), .A2(n13210), .B1(n13208), .B2(n15543), .ZN(
        n11788) );
  NAND3_X1 U14329 ( .A1(n11790), .A2(n11789), .A3(n11788), .ZN(n15591) );
  MUX2_X1 U14330 ( .A(n15591), .B(P3_REG2_REG_8__SCAN_IN), .S(n15561), .Z(
        n11791) );
  AOI211_X1 U14331 ( .C1(n13440), .C2(n15593), .A(n11792), .B(n11791), .ZN(
        n11793) );
  INV_X1 U14332 ( .A(n11793), .ZN(P3_U3225) );
  OAI222_X1 U14333 ( .A1(P2_U3088), .A2(n11795), .B1(n13019), .B2(n11798), 
        .C1(n11794), .C2(n14247), .ZN(P2_U3303) );
  INV_X1 U14334 ( .A(n11796), .ZN(n11799) );
  OAI222_X1 U14335 ( .A1(P1_U3086), .A2(n11799), .B1(n15159), .B2(n11798), 
        .C1(n11797), .C2(n15165), .ZN(P1_U3331) );
  XNOR2_X1 U14336 ( .A(n11800), .B(n11804), .ZN(n11802) );
  NAND2_X1 U14337 ( .A1(n14574), .A2(n15010), .ZN(n11801) );
  OAI21_X1 U14338 ( .B1(n14992), .B2(n14993), .A(n11801), .ZN(n12231) );
  AOI21_X1 U14339 ( .B1(n11802), .B2(n14874), .A(n12231), .ZN(n12301) );
  XNOR2_X1 U14340 ( .A(n11803), .B(n11804), .ZN(n12298) );
  INV_X1 U14341 ( .A(n15023), .ZN(n15282) );
  OAI211_X1 U14342 ( .C1(n11841), .C2(n12307), .A(n6432), .B(n15016), .ZN(
        n12299) );
  OAI22_X1 U14343 ( .A1(n15305), .A2(n11805), .B1(n12234), .B2(n14997), .ZN(
        n11806) );
  AOI21_X1 U14344 ( .B1(n12236), .B2(n14980), .A(n11806), .ZN(n11807) );
  OAI21_X1 U14345 ( .B1(n12299), .B2(n14984), .A(n11807), .ZN(n11808) );
  AOI21_X1 U14346 ( .B1(n12298), .B2(n15282), .A(n11808), .ZN(n11809) );
  OAI21_X1 U14347 ( .B1(n12301), .B2(n15307), .A(n11809), .ZN(P1_U3280) );
  INV_X1 U14348 ( .A(n12558), .ZN(n12452) );
  XNOR2_X1 U14349 ( .A(n11810), .B(n12452), .ZN(n11823) );
  XNOR2_X1 U14350 ( .A(n11811), .B(n12558), .ZN(n11812) );
  AOI222_X1 U14351 ( .A1(n10147), .A2(n11812), .B1(n13558), .B2(n15531), .C1(
        n13207), .C2(n15546), .ZN(n11819) );
  MUX2_X1 U14352 ( .A(n11813), .B(n11819), .S(n15600), .Z(n11815) );
  INV_X1 U14353 ( .A(n12449), .ZN(n13164) );
  NAND2_X1 U14354 ( .A1(n13691), .A2(n13164), .ZN(n11814) );
  OAI211_X1 U14355 ( .C1(n11823), .C2(n13695), .A(n11815), .B(n11814), .ZN(
        P3_U3423) );
  INV_X1 U14356 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11816) );
  MUX2_X1 U14357 ( .A(n11816), .B(n11819), .S(n15559), .Z(n11818) );
  AOI22_X1 U14358 ( .A1(n6428), .A2(n13164), .B1(n15518), .B2(n13163), .ZN(
        n11817) );
  OAI211_X1 U14359 ( .C1(n11823), .C2(n13566), .A(n11818), .B(n11817), .ZN(
        P3_U3222) );
  MUX2_X1 U14360 ( .A(n11820), .B(n11819), .S(n15612), .Z(n11822) );
  NAND2_X1 U14361 ( .A1(n13617), .A2(n13164), .ZN(n11821) );
  OAI211_X1 U14362 ( .C1(n13620), .C2(n11823), .A(n11822), .B(n11821), .ZN(
        P3_U3470) );
  INV_X1 U14363 ( .A(n12149), .ZN(n14091) );
  INV_X1 U14364 ( .A(n12588), .ZN(n11824) );
  AOI22_X1 U14365 ( .A1(n14085), .A2(n12706), .B1(n11824), .B2(n14083), .ZN(
        n11825) );
  OAI21_X1 U14366 ( .B1(n11826), .B2(n14089), .A(n11825), .ZN(n11829) );
  MUX2_X1 U14367 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11827), .S(n14064), .Z(
        n11828) );
  AOI211_X1 U14368 ( .C1(n14091), .C2(n11830), .A(n11829), .B(n11828), .ZN(
        n11831) );
  INV_X1 U14369 ( .A(n11831), .ZN(P2_U3256) );
  AOI22_X1 U14370 ( .A1(n11832), .A2(n15078), .B1(n11833), .B2(n14874), .ZN(
        n11838) );
  INV_X1 U14371 ( .A(n11832), .ZN(n11835) );
  INV_X1 U14372 ( .A(n11833), .ZN(n11834) );
  AOI22_X1 U14373 ( .A1(n11835), .A2(n15078), .B1(n11834), .B2(n14874), .ZN(
        n11837) );
  MUX2_X1 U14374 ( .A(n11838), .B(n11837), .S(n11836), .Z(n11840) );
  AOI22_X1 U14375 ( .A1(n15011), .A2(n15008), .B1(n15010), .B2(n14575), .ZN(
        n11839) );
  NAND2_X1 U14376 ( .A1(n11840), .A2(n11839), .ZN(n12240) );
  INV_X1 U14377 ( .A(n12240), .ZN(n11847) );
  INV_X1 U14378 ( .A(n12072), .ZN(n11842) );
  AOI211_X1 U14379 ( .C1(n12205), .C2(n11842), .A(n15015), .B(n11841), .ZN(
        n12239) );
  NOR2_X1 U14380 ( .A1(n14449), .A2(n15279), .ZN(n11845) );
  OAI22_X1 U14381 ( .A1(n15305), .A2(n11843), .B1(n14443), .B2(n14997), .ZN(
        n11844) );
  AOI211_X1 U14382 ( .C1(n12239), .C2(n15273), .A(n11845), .B(n11844), .ZN(
        n11846) );
  OAI21_X1 U14383 ( .B1(n11847), .B2(n15307), .A(n11846), .ZN(P1_U3281) );
  INV_X1 U14384 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11854) );
  INV_X1 U14385 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n11851) );
  NAND2_X1 U14386 ( .A1(n11851), .A2(n11850), .ZN(n11853) );
  NOR2_X1 U14387 ( .A1(n11851), .A2(n11850), .ZN(n11852) );
  INV_X1 U14388 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11855) );
  NAND2_X1 U14389 ( .A1(n11855), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n12335) );
  INV_X1 U14390 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n11856) );
  NAND2_X1 U14391 ( .A1(n11856), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11857) );
  NAND2_X1 U14392 ( .A1(n12335), .A2(n11857), .ZN(n12334) );
  XNOR2_X1 U14393 ( .A(n12333), .B(n12334), .ZN(n11859) );
  NAND2_X1 U14394 ( .A1(n11858), .A2(n11859), .ZN(n12331) );
  INV_X1 U14395 ( .A(n12331), .ZN(n11865) );
  INV_X1 U14396 ( .A(n11859), .ZN(n11860) );
  INV_X1 U14397 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n11861) );
  NAND2_X1 U14398 ( .A1(n11862), .A2(n11861), .ZN(n12332) );
  INV_X1 U14399 ( .A(n11862), .ZN(n11863) );
  OAI21_X1 U14400 ( .B1(n11863), .B2(n11865), .A(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n11864) );
  OAI21_X1 U14401 ( .B1(n11865), .B2(n12332), .A(n11864), .ZN(SUB_1596_U69) );
  XNOR2_X1 U14402 ( .A(n14212), .B(n12718), .ZN(n12882) );
  XOR2_X1 U14403 ( .A(n11866), .B(n12882), .Z(n14210) );
  OR2_X1 U14404 ( .A1(n13812), .A2(n12262), .ZN(n11868) );
  NAND2_X1 U14405 ( .A1(n13854), .A2(n13802), .ZN(n11867) );
  NAND2_X1 U14406 ( .A1(n11868), .A2(n11867), .ZN(n12267) );
  NAND2_X1 U14407 ( .A1(n11869), .A2(n12882), .ZN(n11870) );
  AOI21_X1 U14408 ( .B1(n12140), .B2(n11870), .A(n14186), .ZN(n11871) );
  AOI211_X1 U14409 ( .C1(n11872), .C2(n14210), .A(n12267), .B(n11871), .ZN(
        n14214) );
  AOI211_X1 U14410 ( .C1(n14212), .C2(n11873), .A(n14166), .B(n6615), .ZN(
        n14211) );
  INV_X1 U14411 ( .A(n14212), .ZN(n12717) );
  NOR2_X1 U14412 ( .A1(n12717), .A2(n15437), .ZN(n11876) );
  OAI22_X1 U14413 ( .A1(n14064), .A2(n11874), .B1(n12269), .B2(n15434), .ZN(
        n11875) );
  AOI211_X1 U14414 ( .C1(n14211), .C2(n15445), .A(n11876), .B(n11875), .ZN(
        n11878) );
  NAND2_X1 U14415 ( .A1(n14210), .A2(n14091), .ZN(n11877) );
  OAI211_X1 U14416 ( .C1(n14214), .C2(n6438), .A(n11878), .B(n11877), .ZN(
        P2_U3254) );
  NAND2_X1 U14417 ( .A1(n6954), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n11879) );
  OAI21_X1 U14418 ( .B1(n11880), .B2(n6954), .A(n11879), .ZN(n12017) );
  INV_X1 U14419 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U14420 ( .A1(n11984), .A2(keyinput5), .B1(n11882), .B2(keyinput35), 
        .ZN(n11881) );
  OAI221_X1 U14421 ( .B1(n11984), .B2(keyinput5), .C1(n11882), .C2(keyinput35), 
        .A(n11881), .ZN(n11892) );
  AOI22_X1 U14422 ( .A1(n13590), .A2(keyinput1), .B1(keyinput51), .B2(n11995), 
        .ZN(n11883) );
  OAI221_X1 U14423 ( .B1(n13590), .B2(keyinput1), .C1(n11995), .C2(keyinput51), 
        .A(n11883), .ZN(n11891) );
  AOI22_X1 U14424 ( .A1(n11886), .A2(keyinput52), .B1(keyinput18), .B2(n11885), 
        .ZN(n11884) );
  OAI221_X1 U14425 ( .B1(n11886), .B2(keyinput52), .C1(n11885), .C2(keyinput18), .A(n11884), .ZN(n11890) );
  AOI22_X1 U14426 ( .A1(n11887), .A2(keyinput11), .B1(n12005), .B2(keyinput25), 
        .ZN(n11888) );
  OAI221_X1 U14427 ( .B1(n11887), .B2(keyinput11), .C1(n12005), .C2(keyinput25), .A(n11888), .ZN(n11889) );
  OR4_X1 U14428 ( .A1(n11892), .A2(n11891), .A3(n11890), .A4(n11889), .ZN(
        n11905) );
  INV_X1 U14429 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U14430 ( .A1(n15451), .A2(keyinput62), .B1(keyinput50), .B2(n11981), 
        .ZN(n11893) );
  OAI221_X1 U14431 ( .B1(n15451), .B2(keyinput62), .C1(n11981), .C2(keyinput50), .A(n11893), .ZN(n11904) );
  AOI22_X1 U14432 ( .A1(n11592), .A2(keyinput33), .B1(n10679), .B2(keyinput22), 
        .ZN(n11894) );
  OAI221_X1 U14433 ( .B1(n11592), .B2(keyinput33), .C1(n10679), .C2(keyinput22), .A(n11894), .ZN(n11903) );
  INV_X1 U14434 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15453) );
  AOI22_X1 U14435 ( .A1(n15453), .A2(keyinput42), .B1(keyinput15), .B2(n11973), 
        .ZN(n11895) );
  OAI221_X1 U14436 ( .B1(n15453), .B2(keyinput42), .C1(n11973), .C2(keyinput15), .A(n11895), .ZN(n11901) );
  INV_X1 U14437 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U14438 ( .A1(n12815), .A2(keyinput20), .B1(keyinput6), .B2(n14375), 
        .ZN(n11896) );
  OAI221_X1 U14439 ( .B1(n12815), .B2(keyinput20), .C1(n14375), .C2(keyinput6), 
        .A(n11896), .ZN(n11900) );
  AOI22_X1 U14440 ( .A1(n12936), .A2(keyinput7), .B1(keyinput36), .B2(n11898), 
        .ZN(n11897) );
  OAI221_X1 U14441 ( .B1(n12936), .B2(keyinput7), .C1(n11898), .C2(keyinput36), 
        .A(n11897), .ZN(n11899) );
  OR3_X1 U14442 ( .A1(n11901), .A2(n11900), .A3(n11899), .ZN(n11902) );
  NOR4_X1 U14443 ( .A1(n11905), .A2(n11904), .A3(n11903), .A4(n11902), .ZN(
        n12015) );
  XOR2_X1 U14444 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput24), .Z(n11910) );
  XOR2_X1 U14445 ( .A(P1_REG3_REG_0__SCAN_IN), .B(keyinput16), .Z(n11909) );
  XOR2_X1 U14446 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput23), .Z(n11908) );
  XNOR2_X1 U14447 ( .A(n11906), .B(keyinput10), .ZN(n11907) );
  NOR4_X1 U14448 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n11930) );
  XNOR2_X1 U14449 ( .A(n11974), .B(keyinput47), .ZN(n11916) );
  XNOR2_X1 U14450 ( .A(n11911), .B(keyinput40), .ZN(n11915) );
  XNOR2_X1 U14451 ( .A(n11912), .B(keyinput61), .ZN(n11914) );
  XNOR2_X1 U14452 ( .A(n6691), .B(keyinput54), .ZN(n11913) );
  NOR4_X1 U14453 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n11929) );
  XNOR2_X1 U14454 ( .A(n11988), .B(keyinput58), .ZN(n11920) );
  XNOR2_X1 U14455 ( .A(n15264), .B(keyinput43), .ZN(n11919) );
  XNOR2_X1 U14456 ( .A(n11991), .B(keyinput27), .ZN(n11918) );
  XNOR2_X1 U14457 ( .A(n11996), .B(keyinput34), .ZN(n11917) );
  NOR4_X1 U14458 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(
        n11928) );
  XNOR2_X1 U14459 ( .A(n11921), .B(keyinput0), .ZN(n11926) );
  XNOR2_X1 U14460 ( .A(n11994), .B(keyinput2), .ZN(n11925) );
  XNOR2_X1 U14461 ( .A(keyinput45), .B(n8790), .ZN(n11924) );
  XNOR2_X1 U14462 ( .A(keyinput49), .B(n11922), .ZN(n11923) );
  NOR4_X1 U14463 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11927) );
  NAND4_X1 U14464 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11927), .ZN(
        n11948) );
  INV_X1 U14465 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15450) );
  AOI22_X1 U14466 ( .A1(n12001), .A2(keyinput48), .B1(n15450), .B2(keyinput12), 
        .ZN(n11931) );
  OAI221_X1 U14467 ( .B1(n12001), .B2(keyinput48), .C1(n15450), .C2(keyinput12), .A(n11931), .ZN(n11947) );
  XNOR2_X1 U14468 ( .A(keyinput41), .B(P3_DATAO_REG_4__SCAN_IN), .ZN(n11935)
         );
  XNOR2_X1 U14469 ( .A(keyinput29), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n11934)
         );
  XNOR2_X1 U14470 ( .A(keyinput31), .B(P2_D_REG_7__SCAN_IN), .ZN(n11933) );
  XNOR2_X1 U14471 ( .A(keyinput14), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n11932)
         );
  NAND4_X1 U14472 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11946) );
  AOI22_X1 U14473 ( .A1(n13372), .A2(keyinput21), .B1(keyinput56), .B2(n8417), 
        .ZN(n11936) );
  OAI221_X1 U14474 ( .B1(n13372), .B2(keyinput21), .C1(n8417), .C2(keyinput56), 
        .A(n11936), .ZN(n11937) );
  INV_X1 U14475 ( .A(n11937), .ZN(n11944) );
  XNOR2_X1 U14476 ( .A(keyinput19), .B(n9076), .ZN(n11939) );
  XNOR2_X1 U14477 ( .A(keyinput55), .B(n8995), .ZN(n11938) );
  NOR2_X1 U14478 ( .A1(n11939), .A2(n11938), .ZN(n11943) );
  AOI22_X1 U14479 ( .A1(n11975), .A2(keyinput26), .B1(n11976), .B2(keyinput13), 
        .ZN(n11940) );
  OAI221_X1 U14480 ( .B1(n11975), .B2(keyinput26), .C1(n11976), .C2(keyinput13), .A(n11940), .ZN(n11941) );
  INV_X1 U14481 ( .A(n11941), .ZN(n11942) );
  NAND3_X1 U14482 ( .A1(n11944), .A2(n11943), .A3(n11942), .ZN(n11945) );
  NOR4_X1 U14483 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n12014) );
  AOI22_X1 U14484 ( .A1(n13110), .A2(keyinput4), .B1(keyinput28), .B2(n10627), 
        .ZN(n11949) );
  OAI221_X1 U14485 ( .B1(n13110), .B2(keyinput4), .C1(n10627), .C2(keyinput28), 
        .A(n11949), .ZN(n11972) );
  AOI22_X1 U14486 ( .A1(n14035), .A2(keyinput44), .B1(n11951), .B2(keyinput63), 
        .ZN(n11950) );
  OAI221_X1 U14487 ( .B1(n14035), .B2(keyinput44), .C1(n11951), .C2(keyinput63), .A(n11950), .ZN(n11965) );
  AOI22_X1 U14488 ( .A1(n8592), .A2(keyinput3), .B1(keyinput32), .B2(n12006), 
        .ZN(n11952) );
  OAI221_X1 U14489 ( .B1(n8592), .B2(keyinput3), .C1(n12006), .C2(keyinput32), 
        .A(n11952), .ZN(n11964) );
  XOR2_X1 U14490 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput17), .Z(n11955) );
  XNOR2_X1 U14491 ( .A(n11953), .B(keyinput59), .ZN(n11954) );
  NOR2_X1 U14492 ( .A1(n11955), .A2(n11954), .ZN(n11957) );
  XNOR2_X1 U14493 ( .A(SI_21_), .B(keyinput8), .ZN(n11956) );
  OAI211_X1 U14494 ( .C1(n10319), .C2(keyinput57), .A(n11957), .B(n11956), 
        .ZN(n11963) );
  XNOR2_X1 U14495 ( .A(P1_REG3_REG_15__SCAN_IN), .B(keyinput38), .ZN(n11961)
         );
  XNOR2_X1 U14496 ( .A(SI_7_), .B(keyinput9), .ZN(n11960) );
  XNOR2_X1 U14497 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput30), .ZN(n11959) );
  XNOR2_X1 U14498 ( .A(SI_2_), .B(keyinput60), .ZN(n11958) );
  NAND4_X1 U14499 ( .A1(n11961), .A2(n11960), .A3(n11959), .A4(n11958), .ZN(
        n11962) );
  OR4_X1 U14500 ( .A1(n11965), .A2(n11964), .A3(n11963), .A4(n11962), .ZN(
        n11971) );
  INV_X1 U14501 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U14502 ( .A1(n12002), .A2(keyinput37), .B1(n11977), .B2(keyinput53), 
        .ZN(n11966) );
  OAI221_X1 U14503 ( .B1(n12002), .B2(keyinput37), .C1(n11977), .C2(keyinput53), .A(n11966), .ZN(n11970) );
  AOI22_X1 U14504 ( .A1(n11968), .A2(keyinput46), .B1(keyinput39), .B2(n14509), 
        .ZN(n11967) );
  OAI221_X1 U14505 ( .B1(n11968), .B2(keyinput46), .C1(n14509), .C2(keyinput39), .A(n11967), .ZN(n11969) );
  NOR4_X1 U14506 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n12013) );
  NOR4_X1 U14507 ( .A1(n11973), .A2(P2_REG0_REG_10__SCAN_IN), .A3(
        P3_DATAO_REG_4__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n11990) );
  NAND3_X1 U14508 ( .A1(P3_REG1_REG_21__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .A3(n11974), .ZN(n11980) );
  NAND4_X1 U14509 ( .A1(SI_7_), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  NAND4_X1 U14510 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_2_), .A3(
        P2_IR_REG_2__SCAN_IN), .A4(P2_REG2_REG_27__SCAN_IN), .ZN(n11978) );
  NOR4_X1 U14511 ( .A1(n11980), .A2(n11979), .A3(n11978), .A4(n13372), .ZN(
        n11986) );
  NAND4_X1 U14512 ( .A1(SI_21_), .A2(P3_IR_REG_9__SCAN_IN), .A3(
        P1_IR_REG_25__SCAN_IN), .A4(n10679), .ZN(n11983) );
  NAND4_X1 U14513 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P1_REG1_REG_2__SCAN_IN), 
        .A3(n12936), .A4(n11981), .ZN(n11982) );
  NOR2_X1 U14514 ( .A1(n11983), .A2(n11982), .ZN(n11985) );
  NAND4_X1 U14515 ( .A1(n11986), .A2(n11985), .A3(n11984), .A4(n14035), .ZN(
        n11987) );
  NOR4_X1 U14516 ( .A1(n11988), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_IR_REG_7__SCAN_IN), .A4(n11987), .ZN(n11989) );
  NAND4_X1 U14517 ( .A1(n11990), .A2(P2_D_REG_19__SCAN_IN), .A3(n11989), .A4(
        P2_D_REG_15__SCAN_IN), .ZN(n12000) );
  NOR4_X1 U14518 ( .A1(n11991), .A2(P1_REG3_REG_22__SCAN_IN), .A3(
        P2_DATAO_REG_22__SCAN_IN), .A4(P1_REG3_REG_4__SCAN_IN), .ZN(n11993) );
  NOR2_X1 U14519 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(P1_REG3_REG_1__SCAN_IN), 
        .ZN(n11992) );
  NAND4_X1 U14520 ( .A1(n11993), .A2(P1_REG2_REG_19__SCAN_IN), .A3(
        P1_REG0_REG_0__SCAN_IN), .A4(n11992), .ZN(n11999) );
  NAND4_X1 U14521 ( .A1(n6691), .A2(P1_REG2_REG_7__SCAN_IN), .A3(
        P3_IR_REG_28__SCAN_IN), .A4(P3_REG3_REG_5__SCAN_IN), .ZN(n11998) );
  NAND4_X1 U14522 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(
        P2_REG2_REG_13__SCAN_IN), .ZN(n11997) );
  OR4_X1 U14523 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12010) );
  NOR4_X1 U14524 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_15__SCAN_IN), 
        .A3(n12815), .A4(n15453), .ZN(n12003) );
  NAND4_X1 U14525 ( .A1(n12004), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12009) );
  NAND4_X1 U14526 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), 
        .A3(n10627), .A4(n12005), .ZN(n12008) );
  NAND4_X1 U14527 ( .A1(P2_REG0_REG_5__SCAN_IN), .A2(P1_REG0_REG_26__SCAN_IN), 
        .A3(n8592), .A4(n12006), .ZN(n12007) );
  NOR4_X1 U14528 ( .A1(n12010), .A2(n12009), .A3(n12008), .A4(n12007), .ZN(
        n12011) );
  OAI21_X1 U14529 ( .B1(n12011), .B2(keyinput57), .A(n10319), .ZN(n12012) );
  NAND4_X1 U14530 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12016) );
  XNOR2_X1 U14531 ( .A(n12017), .B(n12016), .ZN(P2_U3457) );
  NAND2_X1 U14532 ( .A1(n12018), .A2(n13207), .ZN(n12019) );
  INV_X2 U14533 ( .A(n13035), .ZN(n13071) );
  XNOR2_X1 U14534 ( .A(n12125), .B(n13071), .ZN(n12022) );
  NAND2_X1 U14535 ( .A1(n12022), .A2(n13161), .ZN(n12175) );
  XNOR2_X1 U14536 ( .A(n12449), .B(n13071), .ZN(n12172) );
  NAND3_X1 U14537 ( .A1(n12175), .A2(n12448), .A3(n12172), .ZN(n12024) );
  INV_X1 U14538 ( .A(n12022), .ZN(n12023) );
  NAND2_X1 U14539 ( .A1(n12023), .A2(n13558), .ZN(n12174) );
  AND2_X1 U14540 ( .A1(n12024), .A2(n12174), .ZN(n12025) );
  XNOR2_X1 U14541 ( .A(n12029), .B(n13071), .ZN(n12250) );
  XNOR2_X1 U14542 ( .A(n12250), .B(n12246), .ZN(n12026) );
  XNOR2_X1 U14543 ( .A(n12249), .B(n12026), .ZN(n12033) );
  NAND2_X1 U14544 ( .A1(n13190), .A2(n13558), .ZN(n12027) );
  NAND2_X1 U14545 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13252)
         );
  OAI211_X1 U14546 ( .C1(n13193), .C2(n12028), .A(n12027), .B(n13252), .ZN(
        n12031) );
  NOR2_X1 U14547 ( .A1(n12029), .A2(n13177), .ZN(n12030) );
  AOI211_X1 U14548 ( .C1(n13562), .C2(n13195), .A(n12031), .B(n12030), .ZN(
        n12032) );
  OAI21_X1 U14549 ( .B1(n12033), .B2(n13199), .A(n12032), .ZN(P3_U3174) );
  INV_X1 U14550 ( .A(n12034), .ZN(n12035) );
  NAND2_X1 U14551 ( .A1(n14577), .A2(n14351), .ZN(n12036) );
  NAND2_X1 U14552 ( .A1(n12044), .A2(n14295), .ZN(n12038) );
  NAND2_X1 U14553 ( .A1(n14577), .A2(n10794), .ZN(n12037) );
  NAND2_X1 U14554 ( .A1(n12038), .A2(n12037), .ZN(n12208) );
  XNOR2_X1 U14555 ( .A(n12213), .B(n12208), .ZN(n12039) );
  NOR2_X1 U14556 ( .A1(n12223), .A2(n12039), .ZN(n12164) );
  AOI21_X1 U14557 ( .B1(n12223), .B2(n12039), .A(n12164), .ZN(n12046) );
  NAND2_X1 U14558 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n14677) );
  OAI21_X1 U14559 ( .B1(n14555), .B2(n14521), .A(n14677), .ZN(n12043) );
  INV_X1 U14560 ( .A(n14377), .ZN(n14557) );
  OAI22_X1 U14561 ( .A1(n14557), .A2(n12041), .B1(n12040), .B2(n14556), .ZN(
        n12042) );
  AOI211_X1 U14562 ( .C1(n12044), .C2(n10393), .A(n12043), .B(n12042), .ZN(
        n12045) );
  OAI21_X1 U14563 ( .B1(n12046), .B2(n14561), .A(n12045), .ZN(P1_U3231) );
  INV_X1 U14564 ( .A(n12188), .ZN(n12047) );
  AOI22_X1 U14565 ( .A1(n14085), .A2(n12711), .B1(n12047), .B2(n14083), .ZN(
        n12048) );
  OAI21_X1 U14566 ( .B1(n12049), .B2(n14089), .A(n12048), .ZN(n12052) );
  MUX2_X1 U14567 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n12050), .S(n14064), .Z(
        n12051) );
  AOI211_X1 U14568 ( .C1(n14091), .C2(n12053), .A(n12052), .B(n12051), .ZN(
        n12054) );
  INV_X1 U14569 ( .A(n12054), .ZN(P2_U3255) );
  INV_X1 U14570 ( .A(n6428), .ZN(n13495) );
  OAI22_X1 U14571 ( .A1(n13495), .A2(n12064), .B1(n12055), .B2(n15553), .ZN(
        n12058) );
  MUX2_X1 U14572 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n12056), .S(n15559), .Z(
        n12057) );
  AOI211_X1 U14573 ( .C1(n13440), .C2(n12059), .A(n12058), .B(n12057), .ZN(
        n12060) );
  INV_X1 U14574 ( .A(n12060), .ZN(P3_U3223) );
  INV_X1 U14575 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12062) );
  MUX2_X1 U14576 ( .A(n12062), .B(n12061), .S(n15612), .Z(n12063) );
  OAI21_X1 U14577 ( .B1(n13598), .B2(n12064), .A(n12063), .ZN(P3_U3469) );
  INV_X1 U14578 ( .A(n12065), .ZN(n12066) );
  NAND2_X1 U14579 ( .A1(n12067), .A2(n12066), .ZN(n12093) );
  INV_X1 U14580 ( .A(n12093), .ZN(n12068) );
  NAND2_X1 U14581 ( .A1(n12068), .A2(n7719), .ZN(n12094) );
  NAND2_X1 U14582 ( .A1(n12094), .A2(n12069), .ZN(n12070) );
  XNOR2_X1 U14583 ( .A(n12070), .B(n12075), .ZN(n12071) );
  AOI222_X1 U14584 ( .A1(n14874), .A2(n12071), .B1(n14574), .B2(n15008), .C1(
        n14576), .C2(n15010), .ZN(n15119) );
  AOI211_X1 U14585 ( .C1(n15117), .C2(n7740), .A(n15015), .B(n12072), .ZN(
        n15116) );
  INV_X1 U14586 ( .A(n15117), .ZN(n14526) );
  INV_X1 U14587 ( .A(n14520), .ZN(n12073) );
  AOI22_X1 U14588 ( .A1(n15307), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12073), 
        .B2(n15301), .ZN(n12074) );
  OAI21_X1 U14589 ( .B1(n14526), .B2(n15279), .A(n12074), .ZN(n12078) );
  XOR2_X1 U14590 ( .A(n12076), .B(n12075), .Z(n15120) );
  NOR2_X1 U14591 ( .A1(n15120), .A2(n15023), .ZN(n12077) );
  AOI211_X1 U14592 ( .C1(n15116), .C2(n15273), .A(n12078), .B(n12077), .ZN(
        n12079) );
  OAI21_X1 U14593 ( .B1(n15119), .B2(n15307), .A(n12079), .ZN(P1_U3282) );
  NAND2_X1 U14594 ( .A1(n12087), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12083) );
  NAND2_X1 U14595 ( .A1(n12084), .A2(n12083), .ZN(n12081) );
  INV_X1 U14596 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14957) );
  MUX2_X1 U14597 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n14957), .S(n14707), .Z(
        n12080) );
  NAND2_X1 U14598 ( .A1(n12081), .A2(n12080), .ZN(n14709) );
  MUX2_X1 U14599 ( .A(n14957), .B(P1_REG2_REG_17__SCAN_IN), .S(n14707), .Z(
        n12082) );
  NAND3_X1 U14600 ( .A1(n12084), .A2(n12083), .A3(n12082), .ZN(n12085) );
  NAND3_X1 U14601 ( .A1(n14709), .A2(n14733), .A3(n12085), .ZN(n12092) );
  NAND2_X1 U14602 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14477)
         );
  AOI21_X1 U14603 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n12087), .A(n12086), 
        .ZN(n14713) );
  XNOR2_X1 U14604 ( .A(n14707), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n14712) );
  XOR2_X1 U14605 ( .A(n14713), .B(n14712), .Z(n12088) );
  NAND2_X1 U14606 ( .A1(n14739), .A2(n12088), .ZN(n12089) );
  NAND2_X1 U14607 ( .A1(n14477), .A2(n12089), .ZN(n12090) );
  AOI21_X1 U14608 ( .B1(n15269), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n12090), 
        .ZN(n12091) );
  OAI211_X1 U14609 ( .C1(n14719), .C2(n14710), .A(n12092), .B(n12091), .ZN(
        P1_U3260) );
  AOI21_X1 U14610 ( .B1(n12093), .B2(n12098), .A(n14988), .ZN(n12095) );
  NAND2_X1 U14611 ( .A1(n12095), .A2(n12094), .ZN(n12101) );
  OAI21_X1 U14612 ( .B1(n12098), .B2(n12097), .A(n12096), .ZN(n12099) );
  NAND2_X1 U14613 ( .A1(n12099), .A2(n15078), .ZN(n12100) );
  NAND2_X1 U14614 ( .A1(n12101), .A2(n12100), .ZN(n12290) );
  XNOR2_X1 U14615 ( .A(n12102), .B(n7701), .ZN(n12103) );
  NAND2_X1 U14616 ( .A1(n12103), .A2(n6432), .ZN(n12105) );
  AOI22_X1 U14617 ( .A1(n15008), .A2(n14575), .B1(n14577), .B2(n15010), .ZN(
        n12104) );
  NAND2_X1 U14618 ( .A1(n12105), .A2(n12104), .ZN(n12293) );
  NOR2_X1 U14619 ( .A1(n12290), .A2(n12293), .ZN(n12108) );
  INV_X1 U14620 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n12106) );
  MUX2_X1 U14621 ( .A(n12108), .B(n12106), .S(n15317), .Z(n12107) );
  OAI21_X1 U14622 ( .B1(n7701), .B2(n15143), .A(n12107), .ZN(P1_U3489) );
  MUX2_X1 U14623 ( .A(n12109), .B(n12108), .S(n15322), .Z(n12110) );
  OAI21_X1 U14624 ( .B1(n7701), .B2(n15096), .A(n12110), .ZN(P1_U3538) );
  XNOR2_X1 U14625 ( .A(n12111), .B(n12113), .ZN(n12128) );
  OAI211_X1 U14626 ( .C1(n12114), .C2(n12113), .A(n12112), .B(n10147), .ZN(
        n12116) );
  AOI22_X1 U14627 ( .A1(n12448), .A2(n15546), .B1(n15531), .B2(n13546), .ZN(
        n12115) );
  AND2_X1 U14628 ( .A1(n12116), .A2(n12115), .ZN(n12124) );
  MUX2_X1 U14629 ( .A(n12124), .B(n12117), .S(n15598), .Z(n12119) );
  NAND2_X1 U14630 ( .A1(n13691), .A2(n12125), .ZN(n12118) );
  OAI211_X1 U14631 ( .C1(n12128), .C2(n13695), .A(n12119), .B(n12118), .ZN(
        P3_U3426) );
  MUX2_X1 U14632 ( .A(n12124), .B(n12120), .S(n15609), .Z(n12122) );
  NAND2_X1 U14633 ( .A1(n13617), .A2(n12125), .ZN(n12121) );
  OAI211_X1 U14634 ( .C1(n13620), .C2(n12128), .A(n12122), .B(n12121), .ZN(
        P3_U3471) );
  MUX2_X1 U14635 ( .A(n12124), .B(n12123), .S(n15561), .Z(n12127) );
  AOI22_X1 U14636 ( .A1(n6428), .A2(n12125), .B1(n15518), .B2(n12182), .ZN(
        n12126) );
  OAI211_X1 U14637 ( .C1(n12128), .C2(n13566), .A(n12127), .B(n12126), .ZN(
        P3_U3221) );
  XNOR2_X1 U14638 ( .A(n14201), .B(n13852), .ZN(n12888) );
  XOR2_X1 U14639 ( .A(n12129), .B(n12888), .Z(n12130) );
  OAI22_X1 U14640 ( .A1(n12724), .A2(n13814), .B1(n13008), .B2(n13812), .ZN(
        n13004) );
  AOI21_X1 U14641 ( .B1(n12130), .B2(n15479), .A(n13004), .ZN(n14202) );
  AOI211_X1 U14642 ( .C1(n14201), .C2(n7731), .A(n14166), .B(n12310), .ZN(
        n14200) );
  INV_X1 U14643 ( .A(n13006), .ZN(n12131) );
  AOI22_X1 U14644 ( .A1(n6438), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12131), 
        .B2(n14083), .ZN(n12132) );
  OAI21_X1 U14645 ( .B1(n12726), .B2(n15437), .A(n12132), .ZN(n12135) );
  XNOR2_X1 U14646 ( .A(n12133), .B(n12888), .ZN(n14204) );
  NOR2_X1 U14647 ( .A1(n14204), .A2(n14056), .ZN(n12134) );
  AOI211_X1 U14648 ( .C1(n14200), .C2(n15445), .A(n12135), .B(n12134), .ZN(
        n12136) );
  OAI21_X1 U14649 ( .B1(n6438), .B2(n14202), .A(n12136), .ZN(P2_U3251) );
  XNOR2_X1 U14650 ( .A(n12733), .B(n12732), .ZN(n12884) );
  INV_X1 U14651 ( .A(n12884), .ZN(n12137) );
  XNOR2_X1 U14652 ( .A(n12138), .B(n12137), .ZN(n12337) );
  NAND2_X1 U14653 ( .A1(n12140), .A2(n12139), .ZN(n12141) );
  NAND2_X1 U14654 ( .A1(n12141), .A2(n12884), .ZN(n12142) );
  NAND3_X1 U14655 ( .A1(n12276), .A2(n15479), .A3(n12142), .ZN(n12143) );
  AOI22_X1 U14656 ( .A1(n13853), .A2(n13802), .B1(n13801), .B2(n13855), .ZN(
        n12629) );
  OAI211_X1 U14657 ( .C1(n12337), .C2(n14072), .A(n12143), .B(n12629), .ZN(
        n12342) );
  NAND2_X1 U14658 ( .A1(n12342), .A2(n14064), .ZN(n12148) );
  OAI22_X1 U14659 ( .A1(n14064), .A2(n12144), .B1(n12627), .B2(n15434), .ZN(
        n12146) );
  OAI211_X1 U14660 ( .C1(n6615), .C2(n12731), .A(n15443), .B(n12282), .ZN(
        n12339) );
  NOR2_X1 U14661 ( .A1(n12339), .A2(n14089), .ZN(n12145) );
  AOI211_X1 U14662 ( .C1(n14085), .C2(n12733), .A(n12146), .B(n12145), .ZN(
        n12147) );
  OAI211_X1 U14663 ( .C1(n12337), .C2(n12149), .A(n12148), .B(n12147), .ZN(
        P2_U3253) );
  INV_X1 U14664 ( .A(n12150), .ZN(n12155) );
  INV_X1 U14665 ( .A(n12151), .ZN(n12152) );
  OAI222_X1 U14666 ( .A1(n14247), .A2(n12153), .B1(n13019), .B2(n12155), .C1(
        n12152), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U14667 ( .A1(n15165), .A2(n12156), .B1(n15159), .B2(n12155), .C1(
        P1_U3086), .C2(n12154), .ZN(P1_U3330) );
  NOR2_X1 U14668 ( .A1(n12213), .A2(n12208), .ZN(n12207) );
  NAND2_X1 U14669 ( .A1(n12160), .A2(n14346), .ZN(n12158) );
  NAND2_X1 U14670 ( .A1(n14576), .A2(n14295), .ZN(n12157) );
  NAND2_X1 U14671 ( .A1(n12158), .A2(n12157), .ZN(n12159) );
  XNOR2_X1 U14672 ( .A(n12159), .B(n14359), .ZN(n12216) );
  NAND2_X1 U14673 ( .A1(n12160), .A2(n14351), .ZN(n12162) );
  NAND2_X1 U14674 ( .A1(n14576), .A2(n10794), .ZN(n12161) );
  AND2_X1 U14675 ( .A1(n12162), .A2(n12161), .ZN(n12206) );
  INV_X1 U14676 ( .A(n12206), .ZN(n12209) );
  XNOR2_X1 U14677 ( .A(n12216), .B(n12209), .ZN(n12163) );
  NOR3_X1 U14678 ( .A1(n12164), .A2(n12207), .A3(n12163), .ZN(n14437) );
  INV_X1 U14679 ( .A(n14437), .ZN(n14517) );
  OAI21_X1 U14680 ( .B1(n12164), .B2(n12207), .A(n12163), .ZN(n12165) );
  NAND3_X1 U14681 ( .A1(n14517), .A2(n14540), .A3(n12165), .ZN(n12171) );
  INV_X1 U14682 ( .A(n12166), .ZN(n12169) );
  OAI22_X1 U14683 ( .A1(n14557), .A2(n12167), .B1(n12289), .B2(n14556), .ZN(
        n12168) );
  AOI211_X1 U14684 ( .C1(n14534), .C2(n14575), .A(n12169), .B(n12168), .ZN(
        n12170) );
  OAI211_X1 U14685 ( .C1(n7701), .C2(n14550), .A(n12171), .B(n12170), .ZN(
        P1_U3217) );
  XOR2_X1 U14686 ( .A(n12173), .B(n12172), .Z(n13158) );
  AOI22_X1 U14687 ( .A1(n13158), .A2(n12448), .B1(n12173), .B2(n12172), .ZN(
        n12177) );
  NAND2_X1 U14688 ( .A1(n12175), .A2(n12174), .ZN(n12176) );
  XNOR2_X1 U14689 ( .A(n12177), .B(n12176), .ZN(n12184) );
  NAND2_X1 U14690 ( .A1(n13190), .A2(n12448), .ZN(n12178) );
  NAND2_X1 U14691 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13235)
         );
  OAI211_X1 U14692 ( .C1(n13193), .C2(n12246), .A(n12178), .B(n13235), .ZN(
        n12181) );
  NOR2_X1 U14693 ( .A1(n13177), .A2(n12179), .ZN(n12180) );
  AOI211_X1 U14694 ( .C1(n12182), .C2(n13195), .A(n12181), .B(n12180), .ZN(
        n12183) );
  OAI21_X1 U14695 ( .B1(n12184), .B2(n13199), .A(n12183), .ZN(P3_U3164) );
  NAND2_X1 U14696 ( .A1(n13826), .A2(n12185), .ZN(n12186) );
  OAI211_X1 U14697 ( .C1(n15334), .C2(n12188), .A(n12187), .B(n12186), .ZN(
        n12193) );
  INV_X1 U14698 ( .A(n12189), .ZN(n12265) );
  AOI211_X1 U14699 ( .C1(n12191), .C2(n12190), .A(n15327), .B(n12265), .ZN(
        n12192) );
  AOI211_X1 U14700 ( .C1(n12711), .C2(n15332), .A(n12193), .B(n12192), .ZN(
        n12194) );
  INV_X1 U14701 ( .A(n12194), .ZN(P2_U3189) );
  NAND2_X1 U14702 ( .A1(n15117), .A2(n14346), .ZN(n12196) );
  NAND2_X1 U14703 ( .A1(n14575), .A2(n14295), .ZN(n12195) );
  NAND2_X1 U14704 ( .A1(n12196), .A2(n12195), .ZN(n12197) );
  XNOR2_X1 U14705 ( .A(n12197), .B(n11660), .ZN(n14439) );
  NAND2_X1 U14706 ( .A1(n15117), .A2(n14295), .ZN(n12199) );
  NAND2_X1 U14707 ( .A1(n14575), .A2(n10794), .ZN(n12198) );
  NAND2_X1 U14708 ( .A1(n12199), .A2(n12198), .ZN(n12215) );
  INV_X1 U14709 ( .A(n12215), .ZN(n14438) );
  NAND2_X1 U14710 ( .A1(n12216), .A2(n12209), .ZN(n14516) );
  NAND2_X1 U14711 ( .A1(n12213), .A2(n12208), .ZN(n12200) );
  OAI211_X1 U14712 ( .C1(n14439), .C2(n14438), .A(n14516), .B(n12200), .ZN(
        n12222) );
  NAND2_X1 U14713 ( .A1(n12205), .A2(n14346), .ZN(n12202) );
  NAND2_X1 U14714 ( .A1(n14574), .A2(n14295), .ZN(n12201) );
  NAND2_X1 U14715 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  XNOR2_X1 U14716 ( .A(n12203), .B(n14359), .ZN(n12224) );
  AND2_X1 U14717 ( .A1(n14574), .A2(n10794), .ZN(n12204) );
  AOI21_X1 U14718 ( .B1(n12205), .B2(n14351), .A(n12204), .ZN(n12225) );
  XNOR2_X1 U14719 ( .A(n12224), .B(n12225), .ZN(n14441) );
  NOR2_X1 U14720 ( .A1(n12207), .A2(n12206), .ZN(n12217) );
  NOR2_X1 U14721 ( .A1(n12209), .A2(n12208), .ZN(n12212) );
  INV_X1 U14722 ( .A(n12213), .ZN(n12210) );
  NAND2_X1 U14723 ( .A1(n12212), .A2(n12210), .ZN(n12211) );
  OAI211_X1 U14724 ( .C1(n12217), .C2(n12216), .A(n12215), .B(n12211), .ZN(
        n12220) );
  INV_X1 U14725 ( .A(n12212), .ZN(n12214) );
  NOR3_X1 U14726 ( .A1(n12215), .A2(n12214), .A3(n12213), .ZN(n12219) );
  NOR3_X1 U14727 ( .A1(n12217), .A2(n12216), .A3(n12215), .ZN(n12218) );
  AOI211_X1 U14728 ( .C1(n14439), .C2(n12220), .A(n12219), .B(n12218), .ZN(
        n12221) );
  INV_X1 U14729 ( .A(n12225), .ZN(n12226) );
  NAND2_X1 U14730 ( .A1(n12224), .A2(n12226), .ZN(n12227) );
  NAND2_X1 U14731 ( .A1(n14440), .A2(n12227), .ZN(n14266) );
  OR2_X1 U14732 ( .A1(n12307), .A2(n14413), .ZN(n12229) );
  NAND2_X1 U14733 ( .A1(n15011), .A2(n10794), .ZN(n12228) );
  NAND2_X1 U14734 ( .A1(n12229), .A2(n12228), .ZN(n14263) );
  OAI22_X1 U14735 ( .A1(n12307), .A2(n14414), .B1(n14386), .B2(n14413), .ZN(
        n12230) );
  XNOR2_X1 U14736 ( .A(n12230), .B(n14359), .ZN(n14264) );
  XOR2_X1 U14737 ( .A(n14263), .B(n14264), .Z(n14265) );
  XNOR2_X1 U14738 ( .A(n14266), .B(n14265), .ZN(n12238) );
  NAND2_X1 U14739 ( .A1(n12231), .A2(n14547), .ZN(n12232) );
  OAI211_X1 U14740 ( .C1(n14556), .C2(n12234), .A(n12233), .B(n12232), .ZN(
        n12235) );
  AOI21_X1 U14741 ( .B1(n12236), .B2(n10393), .A(n12235), .ZN(n12237) );
  OAI21_X1 U14742 ( .B1(n12238), .B2(n14561), .A(n12237), .ZN(P1_U3234) );
  INV_X1 U14743 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12241) );
  NOR2_X1 U14744 ( .A1(n12240), .A2(n12239), .ZN(n12243) );
  MUX2_X1 U14745 ( .A(n12241), .B(n12243), .S(n15319), .Z(n12242) );
  OAI21_X1 U14746 ( .B1(n14449), .B2(n15143), .A(n12242), .ZN(P1_U3495) );
  MUX2_X1 U14747 ( .A(n12244), .B(n12243), .S(n15322), .Z(n12245) );
  OAI21_X1 U14748 ( .B1(n14449), .B2(n15096), .A(n12245), .ZN(P1_U3540) );
  INV_X1 U14749 ( .A(n12250), .ZN(n12247) );
  NAND2_X1 U14750 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  XNOR2_X1 U14751 ( .A(n13685), .B(n13071), .ZN(n13021) );
  XNOR2_X1 U14752 ( .A(n13021), .B(n13559), .ZN(n13023) );
  XNOR2_X1 U14753 ( .A(n13024), .B(n13023), .ZN(n12257) );
  NAND2_X1 U14754 ( .A1(n13190), .A2(n13546), .ZN(n12253) );
  NAND2_X1 U14755 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13283)
         );
  OAI211_X1 U14756 ( .C1(n13193), .C2(n13113), .A(n12253), .B(n13283), .ZN(
        n12254) );
  AOI21_X1 U14757 ( .B1(n13550), .B2(n13195), .A(n12254), .ZN(n12256) );
  NAND2_X1 U14758 ( .A1(n13685), .A2(n13196), .ZN(n12255) );
  OAI211_X1 U14759 ( .C1(n12257), .C2(n13199), .A(n12256), .B(n12255), .ZN(
        P3_U3155) );
  INV_X1 U14760 ( .A(n12258), .ZN(n12261) );
  OAI222_X1 U14761 ( .A1(n13717), .A2(n12261), .B1(P3_U3151), .B2(n12260), 
        .C1(n12259), .C2(n13719), .ZN(P3_U3270) );
  NOR3_X1 U14762 ( .A1(n12263), .A2(n12262), .A3(n13790), .ZN(n12264) );
  AOI21_X1 U14763 ( .B1(n12265), .B2(n13822), .A(n12264), .ZN(n12274) );
  AOI21_X1 U14764 ( .B1(n13826), .B2(n12267), .A(n12266), .ZN(n12268) );
  OAI21_X1 U14765 ( .B1(n12269), .B2(n15334), .A(n12268), .ZN(n12271) );
  NOR2_X1 U14766 ( .A1(n12636), .A2(n15327), .ZN(n12270) );
  AOI211_X1 U14767 ( .C1(n14212), .C2(n15332), .A(n12271), .B(n12270), .ZN(
        n12272) );
  OAI21_X1 U14768 ( .B1(n12274), .B2(n12273), .A(n12272), .ZN(P2_U3208) );
  NAND2_X1 U14769 ( .A1(n12276), .A2(n12275), .ZN(n12277) );
  XOR2_X1 U14770 ( .A(n12277), .B(n12886), .Z(n12280) );
  NAND2_X1 U14771 ( .A1(n13852), .A2(n13802), .ZN(n12279) );
  NAND2_X1 U14772 ( .A1(n13854), .A2(n13801), .ZN(n12278) );
  NAND2_X1 U14773 ( .A1(n12279), .A2(n12278), .ZN(n13778) );
  AOI21_X1 U14774 ( .B1(n12280), .B2(n15479), .A(n13778), .ZN(n14208) );
  INV_X1 U14775 ( .A(n7731), .ZN(n12281) );
  AOI211_X1 U14776 ( .C1(n14206), .C2(n12282), .A(n14166), .B(n12281), .ZN(
        n14205) );
  INV_X1 U14777 ( .A(n13780), .ZN(n12283) );
  AOI22_X1 U14778 ( .A1(n6438), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12283), 
        .B2(n14083), .ZN(n12284) );
  OAI21_X1 U14779 ( .B1(n7407), .B2(n15437), .A(n12284), .ZN(n12287) );
  XOR2_X1 U14780 ( .A(n12285), .B(n12886), .Z(n14209) );
  NOR2_X1 U14781 ( .A1(n14209), .A2(n14056), .ZN(n12286) );
  AOI211_X1 U14782 ( .C1(n14205), .C2(n15445), .A(n12287), .B(n12286), .ZN(
        n12288) );
  OAI21_X1 U14783 ( .B1(n6438), .B2(n14208), .A(n12288), .ZN(P2_U3252) );
  OAI22_X1 U14784 ( .A1(n7701), .A2(n15279), .B1(n12289), .B2(n14997), .ZN(
        n12292) );
  MUX2_X1 U14785 ( .A(n12290), .B(P1_REG2_REG_10__SCAN_IN), .S(n15307), .Z(
        n12291) );
  AOI211_X1 U14786 ( .C1(n15273), .C2(n12293), .A(n12292), .B(n12291), .ZN(
        n12294) );
  INV_X1 U14787 ( .A(n12294), .ZN(P1_U3283) );
  INV_X1 U14788 ( .A(n12295), .ZN(n12297) );
  OAI222_X1 U14789 ( .A1(P3_U3151), .A2(n9446), .B1(n13717), .B2(n12297), .C1(
        n12296), .C2(n13719), .ZN(P3_U3271) );
  NAND2_X1 U14790 ( .A1(n12298), .A2(n15078), .ZN(n12300) );
  AND3_X1 U14791 ( .A1(n12301), .A2(n12300), .A3(n12299), .ZN(n12304) );
  MUX2_X1 U14792 ( .A(n12302), .B(n12304), .S(n15319), .Z(n12303) );
  OAI21_X1 U14793 ( .B1(n12307), .B2(n15143), .A(n12303), .ZN(P1_U3498) );
  MUX2_X1 U14794 ( .A(n12305), .B(n12304), .S(n15322), .Z(n12306) );
  OAI21_X1 U14795 ( .B1(n12307), .B2(n15096), .A(n12306), .ZN(P1_U3541) );
  XOR2_X1 U14796 ( .A(n12308), .B(n12885), .Z(n14199) );
  XNOR2_X1 U14797 ( .A(n12309), .B(n12885), .ZN(n14197) );
  OAI211_X1 U14798 ( .C1(n12310), .C2(n14195), .A(n14080), .B(n15443), .ZN(
        n14194) );
  OAI22_X1 U14799 ( .A1(n12719), .A2(n13814), .B1(n12727), .B2(n13812), .ZN(
        n13825) );
  INV_X1 U14800 ( .A(n13825), .ZN(n14193) );
  OAI22_X1 U14801 ( .A1(n6438), .A2(n14193), .B1(n13829), .B2(n15434), .ZN(
        n12312) );
  NOR2_X1 U14802 ( .A1(n14195), .A2(n15437), .ZN(n12311) );
  AOI211_X1 U14803 ( .C1(n6438), .C2(P2_REG2_REG_15__SCAN_IN), .A(n12312), .B(
        n12311), .ZN(n12313) );
  OAI21_X1 U14804 ( .B1(n14194), .B2(n14089), .A(n12313), .ZN(n12314) );
  AOI21_X1 U14805 ( .B1(n14197), .B2(n14054), .A(n12314), .ZN(n12315) );
  OAI21_X1 U14806 ( .B1(n14199), .B2(n14056), .A(n12315), .ZN(P2_U3250) );
  OR2_X1 U14807 ( .A1(n12322), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n12316) );
  MUX2_X1 U14808 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11882), .S(n15397), .Z(
        n15399) );
  NAND2_X1 U14809 ( .A1(n15400), .A2(n15399), .ZN(n15398) );
  NAND2_X1 U14810 ( .A1(n15397), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U14811 ( .A1(n15398), .A2(n12318), .ZN(n12319) );
  NAND2_X1 U14812 ( .A1(n15411), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n12321) );
  NAND2_X1 U14813 ( .A1(n12319), .A2(n12323), .ZN(n12320) );
  NAND2_X1 U14814 ( .A1(n12321), .A2(n12320), .ZN(n13869) );
  XNOR2_X1 U14815 ( .A(n13869), .B(n7145), .ZN(n13868) );
  XNOR2_X1 U14816 ( .A(n13868), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n12330) );
  NOR2_X1 U14817 ( .A1(n12322), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n15389) );
  XNOR2_X1 U14818 ( .A(n15397), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15394) );
  XNOR2_X1 U14819 ( .A(n12323), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n15405) );
  INV_X1 U14820 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12324) );
  XOR2_X1 U14821 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13874), .Z(n12327) );
  NAND2_X1 U14822 ( .A1(n15373), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U14823 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13828)
         );
  OAI211_X1 U14824 ( .C1(n15408), .C2(n7145), .A(n12325), .B(n13828), .ZN(
        n12326) );
  AOI21_X1 U14825 ( .B1(n12327), .B2(n15419), .A(n12326), .ZN(n12328) );
  OAI21_X1 U14826 ( .B1(n12330), .B2(n12329), .A(n12328), .ZN(P2_U3229) );
  INV_X1 U14827 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15180) );
  XNOR2_X1 U14828 ( .A(n15180), .B(P1_ADDR_REG_12__SCAN_IN), .ZN(n15181) );
  XNOR2_X1 U14829 ( .A(n15182), .B(n15181), .ZN(n15176) );
  XNOR2_X1 U14830 ( .A(n15175), .B(n11984), .ZN(SUB_1596_U68) );
  INV_X1 U14831 ( .A(n12337), .ZN(n12338) );
  NAND2_X1 U14832 ( .A1(n12338), .A2(n15495), .ZN(n12340) );
  OAI211_X1 U14833 ( .C1(n12731), .C2(n15490), .A(n12340), .B(n12339), .ZN(
        n12341) );
  NOR2_X1 U14834 ( .A1(n12342), .A2(n12341), .ZN(n12345) );
  MUX2_X1 U14835 ( .A(n12343), .B(n12345), .S(n15502), .Z(n12344) );
  INV_X1 U14836 ( .A(n12344), .ZN(P2_U3511) );
  MUX2_X1 U14837 ( .A(n12346), .B(n12345), .S(n15496), .Z(n12347) );
  INV_X1 U14838 ( .A(n12347), .ZN(P2_U3466) );
  INV_X1 U14839 ( .A(n12348), .ZN(n12353) );
  OAI222_X1 U14840 ( .A1(P1_U3086), .A2(n12350), .B1(n15159), .B2(n12353), 
        .C1(n12349), .C2(n15165), .ZN(P1_U3329) );
  INV_X1 U14841 ( .A(n12351), .ZN(n12354) );
  OAI222_X1 U14842 ( .A1(P2_U3088), .A2(n12354), .B1(n14257), .B2(n12353), 
        .C1(n12352), .C2(n14247), .ZN(P2_U3301) );
  INV_X1 U14843 ( .A(n12809), .ZN(n12937) );
  OAI222_X1 U14844 ( .A1(n14247), .A2(n12810), .B1(P2_U3088), .B2(n12355), 
        .C1(n14257), .C2(n12937), .ZN(P2_U3297) );
  NAND2_X1 U14845 ( .A1(n15157), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12356) );
  XNOR2_X1 U14846 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n12372) );
  NAND2_X1 U14847 ( .A1(n12374), .A2(n12372), .ZN(n12360) );
  NAND2_X1 U14848 ( .A1(n12936), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12359) );
  NAND2_X1 U14849 ( .A1(n12360), .A2(n12359), .ZN(n12362) );
  INV_X1 U14850 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14248) );
  XNOR2_X1 U14851 ( .A(n14248), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12361) );
  XNOR2_X1 U14852 ( .A(n12362), .B(n12361), .ZN(n13703) );
  NAND2_X1 U14853 ( .A1(n13703), .A2(n12375), .ZN(n12364) );
  INV_X1 U14854 ( .A(SI_31_), .ZN(n13699) );
  OR2_X1 U14855 ( .A1(n6435), .A2(n13699), .ZN(n12363) );
  INV_X1 U14856 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13366) );
  OR2_X1 U14857 ( .A1(n12365), .A2(n13366), .ZN(n12370) );
  INV_X1 U14858 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13568) );
  OR2_X1 U14859 ( .A1(n12366), .A2(n13568), .ZN(n12369) );
  INV_X1 U14860 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13623) );
  OR2_X1 U14861 ( .A1(n12367), .A2(n13623), .ZN(n12368) );
  INV_X1 U14862 ( .A(n12372), .ZN(n12373) );
  XNOR2_X1 U14863 ( .A(n12374), .B(n12373), .ZN(n12615) );
  NAND2_X1 U14864 ( .A1(n12615), .A2(n12375), .ZN(n12378) );
  OR2_X1 U14865 ( .A1(n6435), .A2(n12616), .ZN(n12377) );
  NAND2_X1 U14866 ( .A1(n13624), .A2(n12382), .ZN(n12379) );
  NAND2_X1 U14867 ( .A1(n12533), .A2(n12379), .ZN(n12541) );
  INV_X1 U14868 ( .A(n13363), .ZN(n13201) );
  INV_X1 U14869 ( .A(n12382), .ZN(n13202) );
  NAND2_X1 U14870 ( .A1(n13571), .A2(n13202), .ZN(n12531) );
  INV_X1 U14871 ( .A(n13361), .ZN(n12532) );
  AOI21_X1 U14872 ( .B1(n13201), .B2(n12531), .A(n12532), .ZN(n12383) );
  MUX2_X1 U14873 ( .A(n12481), .B(n12479), .S(n12524), .Z(n12488) );
  OAI211_X1 U14874 ( .C1(n12561), .C2(n12388), .A(n12470), .B(n12387), .ZN(
        n12389) );
  NAND2_X1 U14875 ( .A1(n12389), .A2(n12524), .ZN(n12467) );
  MUX2_X1 U14876 ( .A(n9470), .B(n12390), .S(n12524), .Z(n12401) );
  NAND2_X1 U14877 ( .A1(n12393), .A2(n12392), .ZN(n12397) );
  NAND4_X1 U14878 ( .A1(n12391), .A2(n12397), .A3(n12582), .A4(n12395), .ZN(
        n12399) );
  NAND2_X1 U14879 ( .A1(n12395), .A2(n12394), .ZN(n12396) );
  NAND4_X1 U14880 ( .A1(n12397), .A2(n12524), .A3(n9470), .A4(n12396), .ZN(
        n12398) );
  NAND4_X1 U14881 ( .A1(n12400), .A2(n12401), .A3(n12399), .A4(n12398), .ZN(
        n12406) );
  NAND2_X1 U14882 ( .A1(n12409), .A2(n12402), .ZN(n12403) );
  NAND2_X1 U14883 ( .A1(n12403), .A2(n12529), .ZN(n12405) );
  INV_X1 U14884 ( .A(n12408), .ZN(n12404) );
  AOI21_X1 U14885 ( .B1(n12406), .B2(n12405), .A(n12404), .ZN(n12412) );
  AOI21_X1 U14886 ( .B1(n12408), .B2(n12407), .A(n12529), .ZN(n12411) );
  OR2_X1 U14887 ( .A1(n12409), .A2(n12529), .ZN(n12410) );
  OAI211_X1 U14888 ( .C1(n12412), .C2(n12411), .A(n12551), .B(n12410), .ZN(
        n12423) );
  AND2_X1 U14889 ( .A1(n13213), .A2(n12413), .ZN(n12415) );
  MUX2_X1 U14890 ( .A(n12415), .B(n12414), .S(n12524), .Z(n12416) );
  NOR2_X1 U14891 ( .A1(n12416), .A2(n12547), .ZN(n12422) );
  NAND2_X1 U14892 ( .A1(n12425), .A2(n12417), .ZN(n12420) );
  NAND2_X1 U14893 ( .A1(n12424), .A2(n12418), .ZN(n12419) );
  MUX2_X1 U14894 ( .A(n12420), .B(n12419), .S(n12524), .Z(n12421) );
  AOI21_X1 U14895 ( .B1(n12423), .B2(n12422), .A(n12421), .ZN(n12434) );
  MUX2_X1 U14896 ( .A(n12425), .B(n12424), .S(n12529), .Z(n12427) );
  NAND2_X1 U14897 ( .A1(n12427), .A2(n12426), .ZN(n12433) );
  NOR2_X1 U14898 ( .A1(n13210), .A2(n12524), .ZN(n12430) );
  AND2_X1 U14899 ( .A1(n13210), .A2(n12524), .ZN(n12429) );
  MUX2_X1 U14900 ( .A(n12430), .B(n12429), .S(n12428), .Z(n12431) );
  NOR2_X1 U14901 ( .A1(n12555), .A2(n12431), .ZN(n12432) );
  OAI21_X1 U14902 ( .B1(n12434), .B2(n12433), .A(n12432), .ZN(n12438) );
  NAND2_X1 U14903 ( .A1(n13087), .A2(n12524), .ZN(n12436) );
  OR2_X1 U14904 ( .A1(n13087), .A2(n12524), .ZN(n12435) );
  MUX2_X1 U14905 ( .A(n12436), .B(n12435), .S(n13209), .Z(n12437) );
  NAND3_X1 U14906 ( .A1(n12438), .A2(n15506), .A3(n12437), .ZN(n12442) );
  MUX2_X1 U14907 ( .A(n12440), .B(n12439), .S(n12529), .Z(n12441) );
  NAND4_X1 U14908 ( .A1(n12442), .A2(n12557), .A3(n12558), .A4(n12441), .ZN(
        n12447) );
  OAI211_X1 U14909 ( .C1(n12452), .C2(n12444), .A(n12456), .B(n12443), .ZN(
        n12445) );
  NAND2_X1 U14910 ( .A1(n12445), .A2(n12524), .ZN(n12446) );
  NAND2_X1 U14911 ( .A1(n12447), .A2(n12446), .ZN(n12455) );
  NAND2_X1 U14912 ( .A1(n12449), .A2(n12448), .ZN(n12450) );
  OAI211_X1 U14913 ( .C1(n12452), .C2(n12451), .A(n12454), .B(n12450), .ZN(
        n12453) );
  AOI22_X1 U14914 ( .A1(n12455), .A2(n12454), .B1(n12529), .B2(n12453), .ZN(
        n12461) );
  OAI21_X1 U14915 ( .B1(n12524), .B2(n12456), .A(n13556), .ZN(n12460) );
  MUX2_X1 U14916 ( .A(n12458), .B(n12457), .S(n12524), .Z(n12459) );
  OAI211_X1 U14917 ( .C1(n12461), .C2(n12460), .A(n13545), .B(n12459), .ZN(
        n12462) );
  NAND2_X1 U14918 ( .A1(n12464), .A2(n13534), .ZN(n12466) );
  AOI21_X1 U14919 ( .B1(n12467), .B2(n12466), .A(n12465), .ZN(n12472) );
  AOI21_X1 U14920 ( .B1(n12469), .B2(n12468), .A(n12524), .ZN(n12471) );
  OAI22_X1 U14921 ( .A1(n12472), .A2(n12471), .B1(n12524), .B2(n12470), .ZN(
        n12475) );
  NOR2_X1 U14922 ( .A1(n12473), .A2(n12529), .ZN(n12474) );
  AOI21_X1 U14923 ( .B1(n12475), .B2(n13513), .A(n12474), .ZN(n12486) );
  NAND2_X1 U14924 ( .A1(n12480), .A2(n12476), .ZN(n12477) );
  NAND3_X1 U14925 ( .A1(n12479), .A2(n12478), .A3(n12477), .ZN(n12483) );
  NAND2_X1 U14926 ( .A1(n12481), .A2(n12480), .ZN(n12482) );
  MUX2_X1 U14927 ( .A(n12483), .B(n12482), .S(n12524), .Z(n12484) );
  INV_X1 U14928 ( .A(n12484), .ZN(n12485) );
  OAI21_X1 U14929 ( .B1(n12486), .B2(n13502), .A(n12485), .ZN(n12487) );
  NAND2_X1 U14930 ( .A1(n13594), .A2(n13064), .ZN(n12489) );
  MUX2_X1 U14931 ( .A(n12490), .B(n12489), .S(n12524), .Z(n12491) );
  NAND3_X1 U14932 ( .A1(n13454), .A2(n12492), .A3(n12491), .ZN(n12496) );
  MUX2_X1 U14933 ( .A(n12494), .B(n12493), .S(n12524), .Z(n12495) );
  NAND3_X1 U14934 ( .A1(n12496), .A2(n13443), .A3(n12495), .ZN(n12503) );
  NAND2_X1 U14935 ( .A1(n12503), .A2(n12497), .ZN(n12501) );
  INV_X1 U14936 ( .A(n12498), .ZN(n13408) );
  NAND2_X1 U14937 ( .A1(n12506), .A2(n13408), .ZN(n12499) );
  OAI211_X1 U14938 ( .C1(n12544), .C2(n12501), .A(n12500), .B(n12499), .ZN(
        n12509) );
  NAND2_X1 U14939 ( .A1(n12503), .A2(n12502), .ZN(n12507) );
  OR2_X1 U14940 ( .A1(n13407), .A2(n12504), .ZN(n12505) );
  OAI211_X1 U14941 ( .C1(n12544), .C2(n12507), .A(n12506), .B(n12505), .ZN(
        n12508) );
  MUX2_X1 U14942 ( .A(n12509), .B(n12508), .S(n12529), .Z(n12511) );
  NAND2_X1 U14943 ( .A1(n12511), .A2(n12510), .ZN(n12516) );
  NAND2_X1 U14944 ( .A1(n12517), .A2(n12518), .ZN(n12543) );
  NOR2_X1 U14945 ( .A1(n13403), .A2(n13416), .ZN(n12513) );
  MUX2_X1 U14946 ( .A(n12513), .B(n12512), .S(n12529), .Z(n12514) );
  NOR2_X1 U14947 ( .A1(n12543), .A2(n12514), .ZN(n12515) );
  MUX2_X1 U14948 ( .A(n12518), .B(n12517), .S(n12529), .Z(n12519) );
  OR2_X1 U14949 ( .A1(n12520), .A2(n12529), .ZN(n12521) );
  NAND2_X1 U14950 ( .A1(n12522), .A2(n13072), .ZN(n12530) );
  OAI21_X1 U14951 ( .B1(n12525), .B2(n12524), .A(n12523), .ZN(n12526) );
  NAND2_X1 U14952 ( .A1(n12530), .A2(n12526), .ZN(n12528) );
  OAI211_X1 U14953 ( .C1(n12530), .C2(n12529), .A(n12528), .B(n12527), .ZN(
        n12535) );
  OAI21_X1 U14954 ( .B1(n12532), .B2(n13201), .A(n12531), .ZN(n12540) );
  NAND2_X1 U14955 ( .A1(n12539), .A2(n12537), .ZN(n12538) );
  INV_X1 U14956 ( .A(n12540), .ZN(n12572) );
  INV_X1 U14957 ( .A(n12541), .ZN(n12571) );
  INV_X1 U14958 ( .A(n12544), .ZN(n12565) );
  INV_X1 U14959 ( .A(n13443), .ZN(n13444) );
  INV_X1 U14960 ( .A(n13556), .ZN(n13555) );
  NOR2_X1 U14961 ( .A1(n12546), .A2(n12545), .ZN(n12550) );
  NOR3_X1 U14962 ( .A1(n12548), .A2(n12547), .A3(n15528), .ZN(n12549) );
  NAND4_X1 U14963 ( .A1(n12552), .A2(n12551), .A3(n12550), .A4(n12549), .ZN(
        n12554) );
  NOR4_X1 U14964 ( .A1(n12555), .A2(n12554), .A3(n15504), .A4(n12553), .ZN(
        n12556) );
  NAND4_X1 U14965 ( .A1(n12559), .A2(n12558), .A3(n12557), .A4(n12556), .ZN(
        n12560) );
  NOR4_X1 U14966 ( .A1(n12561), .A2(n13543), .A3(n13555), .A4(n12560), .ZN(
        n12562) );
  NAND4_X1 U14967 ( .A1(n9481), .A2(n13513), .A3(n13523), .A4(n12562), .ZN(
        n12563) );
  NOR4_X1 U14968 ( .A1(n9299), .A2(n13444), .A3(n13485), .A4(n12563), .ZN(
        n12564) );
  NAND4_X1 U14969 ( .A1(n13389), .A2(n12565), .A3(n12564), .A4(n13465), .ZN(
        n12567) );
  NOR4_X1 U14970 ( .A1(n12568), .A2(n9394), .A3(n12567), .A4(n12566), .ZN(
        n12569) );
  NAND4_X1 U14971 ( .A1(n12572), .A2(n12571), .A3(n12570), .A4(n12569), .ZN(
        n12574) );
  XNOR2_X1 U14972 ( .A(n12574), .B(n12573), .ZN(n12576) );
  NAND2_X1 U14973 ( .A1(n12576), .A2(n10877), .ZN(n12577) );
  NAND3_X1 U14974 ( .A1(n12580), .A2(n12579), .A3(n13714), .ZN(n12581) );
  OAI211_X1 U14975 ( .C1(n12582), .C2(n12584), .A(n12581), .B(P3_B_REG_SCAN_IN), .ZN(n12583) );
  AOI21_X1 U14976 ( .B1(n13826), .B2(n12586), .A(n12585), .ZN(n12587) );
  OAI21_X1 U14977 ( .B1(n12588), .B2(n15334), .A(n12587), .ZN(n12594) );
  AOI22_X1 U14978 ( .A1(n13821), .A2(n13859), .B1(n13822), .B2(n12589), .ZN(
        n12591) );
  NOR3_X1 U14979 ( .A1(n12592), .A2(n12591), .A3(n12590), .ZN(n12593) );
  AOI211_X1 U14980 ( .C1(n12706), .C2(n15332), .A(n12594), .B(n12593), .ZN(
        n12595) );
  OAI21_X1 U14981 ( .B1(n12596), .B2(n15327), .A(n12595), .ZN(P2_U3203) );
  XNOR2_X1 U14982 ( .A(n12599), .B(n12597), .ZN(n13823) );
  NAND2_X1 U14983 ( .A1(n13823), .A2(n12598), .ZN(n13824) );
  OAI21_X1 U14984 ( .B1(n12600), .B2(n12599), .A(n13824), .ZN(n13746) );
  XNOR2_X1 U14985 ( .A(n12602), .B(n12601), .ZN(n13747) );
  NOR2_X1 U14986 ( .A1(n13746), .A2(n13747), .ZN(n13745) );
  AOI22_X1 U14987 ( .A1(n12603), .A2(n13822), .B1(n13821), .B2(n13850), .ZN(
        n12605) );
  OR3_X1 U14988 ( .A1(n13745), .A2(n12605), .A3(n12604), .ZN(n12609) );
  OAI22_X1 U14989 ( .A1(n12645), .A2(n13814), .B1(n12719), .B2(n13812), .ZN(
        n14180) );
  NAND2_X1 U14990 ( .A1(n14180), .A2(n13826), .ZN(n12606) );
  NAND2_X1 U14991 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13888)
         );
  OAI211_X1 U14992 ( .C1(n15334), .C2(n14059), .A(n12606), .B(n13888), .ZN(
        n12607) );
  AOI21_X1 U14993 ( .B1(n14181), .B2(n15332), .A(n12607), .ZN(n12608) );
  OAI211_X1 U14994 ( .C1(n15327), .C2(n12610), .A(n12609), .B(n12608), .ZN(
        P2_U3200) );
  NAND2_X1 U14995 ( .A1(n13630), .A2(n13617), .ZN(n12614) );
  INV_X1 U14996 ( .A(n12615), .ZN(n12618) );
  OAI222_X1 U14997 ( .A1(n13717), .A2(n12618), .B1(n12617), .B2(P3_U3151), 
        .C1(n12616), .C2(n13719), .ZN(P3_U3265) );
  INV_X1 U14998 ( .A(n12997), .ZN(n12619) );
  AOI22_X1 U14999 ( .A1(n12619), .A2(n14083), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n6438), .ZN(n12620) );
  OAI21_X1 U15000 ( .B1(n12993), .B2(n15437), .A(n12620), .ZN(n12623) );
  NOR2_X1 U15001 ( .A1(n12621), .A2(n6438), .ZN(n12622) );
  AOI211_X1 U15002 ( .C1(n15445), .C2(n12624), .A(n12623), .B(n12622), .ZN(
        n12625) );
  OAI21_X1 U15003 ( .B1(n12626), .B2(n14056), .A(n12625), .ZN(P2_U3237) );
  NOR2_X1 U15004 ( .A1(n15334), .A2(n12627), .ZN(n12631) );
  OAI21_X1 U15005 ( .B1(n15325), .B2(n12629), .A(n12628), .ZN(n12630) );
  AOI211_X1 U15006 ( .C1(n12733), .C2(n15332), .A(n12631), .B(n12630), .ZN(
        n12638) );
  INV_X1 U15007 ( .A(n12632), .ZN(n12635) );
  OAI22_X1 U15008 ( .A1(n12633), .A2(n15327), .B1(n12718), .B2(n13790), .ZN(
        n12634) );
  NAND3_X1 U15009 ( .A1(n12636), .A2(n12635), .A3(n12634), .ZN(n12637) );
  OAI211_X1 U15010 ( .C1(n12639), .C2(n15327), .A(n12638), .B(n12637), .ZN(
        P2_U3196) );
  INV_X1 U15011 ( .A(n12645), .ZN(n13848) );
  NAND3_X1 U15012 ( .A1(n12640), .A2(n13821), .A3(n13848), .ZN(n12641) );
  OAI21_X1 U15013 ( .B1(n13799), .B2(n15327), .A(n12641), .ZN(n12644) );
  INV_X1 U15014 ( .A(n12642), .ZN(n12643) );
  NAND2_X1 U15015 ( .A1(n12644), .A2(n12643), .ZN(n12650) );
  NOR2_X1 U15016 ( .A1(n15334), .A2(n14034), .ZN(n12648) );
  NOR2_X1 U15017 ( .A1(n12645), .A2(n13812), .ZN(n12646) );
  AOI21_X1 U15018 ( .B1(n13846), .B2(n13802), .A(n12646), .ZN(n14165) );
  NAND2_X1 U15019 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13918)
         );
  OAI21_X1 U15020 ( .B1(n14165), .B2(n15325), .A(n13918), .ZN(n12647) );
  AOI211_X1 U15021 ( .C1(n14163), .C2(n15332), .A(n12648), .B(n12647), .ZN(
        n12649) );
  OAI211_X1 U15022 ( .C1(n15327), .C2(n12651), .A(n12650), .B(n12649), .ZN(
        P2_U3191) );
  INV_X1 U15023 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n12654) );
  NAND2_X1 U15024 ( .A1(n14752), .A2(n15124), .ZN(n14751) );
  XNOR2_X1 U15025 ( .A(n14751), .B(n12659), .ZN(n12652) );
  NAND2_X1 U15026 ( .A1(n12652), .A2(n6432), .ZN(n14750) );
  NAND2_X1 U15027 ( .A1(n14563), .A2(n12653), .ZN(n15027) );
  OAI21_X1 U15028 ( .B1(n12659), .B2(n15143), .A(n12655), .ZN(P1_U3527) );
  INV_X1 U15029 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n12657) );
  OAI21_X1 U15030 ( .B1(n12659), .B2(n15096), .A(n12658), .ZN(P1_U3559) );
  INV_X1 U15031 ( .A(n12901), .ZN(n12660) );
  NAND2_X1 U15032 ( .A1(n14222), .A2(n12660), .ZN(n12662) );
  NAND2_X1 U15033 ( .A1(n6447), .A2(n12663), .ZN(n12664) );
  MUX2_X1 U15034 ( .A(n13866), .B(n12665), .S(n6446), .Z(n12668) );
  MUX2_X1 U15035 ( .A(n12666), .B(n13866), .S(n6447), .Z(n12667) );
  INV_X1 U15036 ( .A(n12668), .ZN(n12669) );
  MUX2_X1 U15037 ( .A(n12670), .B(n13865), .S(n6447), .Z(n12674) );
  NAND2_X1 U15038 ( .A1(n12673), .A2(n12674), .ZN(n12672) );
  MUX2_X1 U15039 ( .A(n13865), .B(n12670), .S(n6447), .Z(n12671) );
  NAND2_X1 U15040 ( .A1(n12672), .A2(n12671), .ZN(n12678) );
  INV_X1 U15041 ( .A(n12673), .ZN(n12676) );
  INV_X1 U15042 ( .A(n12674), .ZN(n12675) );
  NAND2_X1 U15043 ( .A1(n12676), .A2(n12675), .ZN(n12677) );
  NAND2_X1 U15044 ( .A1(n12678), .A2(n12677), .ZN(n12680) );
  MUX2_X1 U15045 ( .A(n13864), .B(n15471), .S(n6447), .Z(n12681) );
  MUX2_X1 U15046 ( .A(n15471), .B(n13864), .S(n6447), .Z(n12679) );
  INV_X1 U15047 ( .A(n12681), .ZN(n12682) );
  MUX2_X1 U15048 ( .A(n12683), .B(n13863), .S(n6447), .Z(n12686) );
  MUX2_X1 U15049 ( .A(n13863), .B(n12683), .S(n6447), .Z(n12684) );
  INV_X1 U15050 ( .A(n12686), .ZN(n12687) );
  MUX2_X1 U15051 ( .A(n13862), .B(n12933), .S(n6447), .Z(n12690) );
  MUX2_X1 U15052 ( .A(n12933), .B(n13862), .S(n6447), .Z(n12688) );
  INV_X1 U15053 ( .A(n12690), .ZN(n12691) );
  MUX2_X1 U15054 ( .A(n12692), .B(n13861), .S(n6446), .Z(n12696) );
  MUX2_X1 U15055 ( .A(n13861), .B(n12692), .S(n6447), .Z(n12693) );
  NAND2_X1 U15056 ( .A1(n12694), .A2(n12693), .ZN(n12699) );
  INV_X1 U15057 ( .A(n12695), .ZN(n12697) );
  NAND2_X1 U15058 ( .A1(n12697), .A2(n7444), .ZN(n12698) );
  NAND2_X1 U15059 ( .A1(n12699), .A2(n12698), .ZN(n12702) );
  MUX2_X1 U15060 ( .A(n13860), .B(n12700), .S(n6447), .Z(n12703) );
  MUX2_X1 U15061 ( .A(n12700), .B(n13860), .S(n6447), .Z(n12701) );
  MUX2_X1 U15062 ( .A(n13859), .B(n14217), .S(n6436), .Z(n12705) );
  MUX2_X1 U15063 ( .A(n13859), .B(n14217), .S(n12728), .Z(n12704) );
  MUX2_X1 U15064 ( .A(n13857), .B(n12706), .S(n12728), .Z(n12709) );
  MUX2_X1 U15065 ( .A(n13857), .B(n12706), .S(n6436), .Z(n12707) );
  INV_X1 U15066 ( .A(n12709), .ZN(n12710) );
  MUX2_X1 U15067 ( .A(n13856), .B(n12711), .S(n6436), .Z(n12715) );
  MUX2_X1 U15068 ( .A(n13856), .B(n12711), .S(n12728), .Z(n12712) );
  INV_X1 U15069 ( .A(n12714), .ZN(n12716) );
  MUX2_X1 U15070 ( .A(n12718), .B(n12717), .S(n12728), .Z(n12735) );
  MUX2_X1 U15071 ( .A(n13855), .B(n14212), .S(n6436), .Z(n12734) );
  NOR2_X1 U15072 ( .A1(n12719), .A2(n6447), .ZN(n12720) );
  AOI21_X1 U15073 ( .B1(n14086), .B2(n6446), .A(n12720), .ZN(n12722) );
  NAND3_X1 U15074 ( .A1(n6564), .A2(n12722), .A3(n12721), .ZN(n12753) );
  MUX2_X1 U15075 ( .A(n13850), .B(n14086), .S(n6436), .Z(n12743) );
  XNOR2_X1 U15076 ( .A(n14181), .B(n13849), .ZN(n14066) );
  NAND2_X1 U15077 ( .A1(n12743), .A2(n14066), .ZN(n12723) );
  NAND2_X1 U15078 ( .A1(n12753), .A2(n12723), .ZN(n12748) );
  MUX2_X1 U15079 ( .A(n12724), .B(n14195), .S(n6436), .Z(n12745) );
  MUX2_X1 U15080 ( .A(n13831), .B(n13851), .S(n6436), .Z(n12744) );
  NAND2_X1 U15081 ( .A1(n12745), .A2(n12744), .ZN(n12725) );
  NAND2_X1 U15082 ( .A1(n12748), .A2(n12725), .ZN(n12758) );
  MUX2_X1 U15083 ( .A(n12727), .B(n12726), .S(n6436), .Z(n12757) );
  MUX2_X1 U15084 ( .A(n13852), .B(n14201), .S(n6447), .Z(n12756) );
  AND2_X1 U15085 ( .A1(n12757), .A2(n12756), .ZN(n12729) );
  OR2_X1 U15086 ( .A1(n12758), .A2(n12729), .ZN(n12762) );
  MUX2_X1 U15087 ( .A(n13008), .B(n7407), .S(n6436), .Z(n12740) );
  MUX2_X1 U15088 ( .A(n13853), .B(n14206), .S(n12728), .Z(n12739) );
  AND2_X1 U15089 ( .A1(n12740), .A2(n12739), .ZN(n12730) );
  NOR2_X1 U15090 ( .A1(n12762), .A2(n12730), .ZN(n12768) );
  MUX2_X1 U15091 ( .A(n12732), .B(n12731), .S(n6436), .Z(n12765) );
  MUX2_X1 U15092 ( .A(n13854), .B(n12733), .S(n12728), .Z(n12764) );
  INV_X1 U15093 ( .A(n12734), .ZN(n12737) );
  INV_X1 U15094 ( .A(n12735), .ZN(n12736) );
  AOI22_X1 U15095 ( .A1(n12765), .A2(n12764), .B1(n12737), .B2(n12736), .ZN(
        n12738) );
  INV_X1 U15096 ( .A(n12739), .ZN(n12742) );
  INV_X1 U15097 ( .A(n12740), .ZN(n12741) );
  NAND2_X1 U15098 ( .A1(n12742), .A2(n12741), .ZN(n12761) );
  INV_X1 U15099 ( .A(n12743), .ZN(n12754) );
  INV_X1 U15100 ( .A(n12744), .ZN(n12747) );
  INV_X1 U15101 ( .A(n12745), .ZN(n12746) );
  NAND3_X1 U15102 ( .A1(n12748), .A2(n12747), .A3(n12746), .ZN(n12752) );
  AND2_X1 U15103 ( .A1(n13849), .A2(n12728), .ZN(n12750) );
  OAI21_X1 U15104 ( .B1(n13849), .B2(n12728), .A(n14181), .ZN(n12749) );
  OAI21_X1 U15105 ( .B1(n12750), .B2(n14181), .A(n12749), .ZN(n12751) );
  OAI211_X1 U15106 ( .C1(n12754), .C2(n12753), .A(n12752), .B(n12751), .ZN(
        n12755) );
  INV_X1 U15107 ( .A(n12755), .ZN(n12760) );
  OR3_X1 U15108 ( .A1(n12758), .A2(n12757), .A3(n12756), .ZN(n12759) );
  OAI211_X1 U15109 ( .C1(n12762), .C2(n12761), .A(n12760), .B(n12759), .ZN(
        n12763) );
  INV_X1 U15110 ( .A(n12763), .ZN(n12770) );
  INV_X1 U15111 ( .A(n12764), .ZN(n12767) );
  INV_X1 U15112 ( .A(n12765), .ZN(n12766) );
  NAND3_X1 U15113 ( .A1(n12768), .A2(n12767), .A3(n12766), .ZN(n12769) );
  NAND3_X1 U15114 ( .A1(n12771), .A2(n12770), .A3(n12769), .ZN(n12774) );
  MUX2_X1 U15115 ( .A(n14048), .B(n13848), .S(n12728), .Z(n12775) );
  NAND2_X1 U15116 ( .A1(n12774), .A2(n12775), .ZN(n12773) );
  MUX2_X1 U15117 ( .A(n13848), .B(n14048), .S(n12728), .Z(n12772) );
  NAND2_X1 U15118 ( .A1(n12773), .A2(n12772), .ZN(n12779) );
  INV_X1 U15119 ( .A(n12774), .ZN(n12777) );
  INV_X1 U15120 ( .A(n12775), .ZN(n12776) );
  NAND2_X1 U15121 ( .A1(n12777), .A2(n12776), .ZN(n12778) );
  NAND2_X1 U15122 ( .A1(n12779), .A2(n12778), .ZN(n12782) );
  MUX2_X1 U15123 ( .A(n13847), .B(n14163), .S(n12728), .Z(n12781) );
  MUX2_X1 U15124 ( .A(n13847), .B(n14163), .S(n6436), .Z(n12780) );
  MUX2_X1 U15125 ( .A(n14159), .B(n13846), .S(n12728), .Z(n12786) );
  MUX2_X1 U15126 ( .A(n13846), .B(n14159), .S(n12728), .Z(n12783) );
  INV_X1 U15127 ( .A(n12785), .ZN(n12788) );
  INV_X1 U15128 ( .A(n12786), .ZN(n12787) );
  MUX2_X1 U15129 ( .A(n14151), .B(n13845), .S(n6436), .Z(n12790) );
  MUX2_X1 U15130 ( .A(n14151), .B(n13845), .S(n12728), .Z(n12789) );
  INV_X1 U15131 ( .A(n12790), .ZN(n12791) );
  MUX2_X1 U15132 ( .A(n14147), .B(n13844), .S(n12728), .Z(n12793) );
  MUX2_X1 U15133 ( .A(n13844), .B(n14147), .S(n12728), .Z(n12792) );
  INV_X1 U15134 ( .A(n12793), .ZN(n12794) );
  MUX2_X1 U15135 ( .A(n13843), .B(n14138), .S(n12728), .Z(n12798) );
  NAND2_X1 U15136 ( .A1(n12797), .A2(n12798), .ZN(n12796) );
  MUX2_X1 U15137 ( .A(n13843), .B(n14138), .S(n6436), .Z(n12795) );
  INV_X1 U15138 ( .A(n12797), .ZN(n12800) );
  INV_X1 U15139 ( .A(n12798), .ZN(n12799) );
  NAND2_X1 U15140 ( .A1(n12800), .A2(n12799), .ZN(n12801) );
  MUX2_X1 U15141 ( .A(n13970), .B(n13842), .S(n12728), .Z(n12803) );
  MUX2_X1 U15142 ( .A(n13842), .B(n13970), .S(n12728), .Z(n12802) );
  INV_X1 U15143 ( .A(n12803), .ZN(n12804) );
  MUX2_X1 U15144 ( .A(n13841), .B(n13958), .S(n12728), .Z(n12807) );
  MUX2_X1 U15145 ( .A(n13813), .B(n14126), .S(n6436), .Z(n12805) );
  INV_X1 U15146 ( .A(n12806), .ZN(n12808) );
  NAND2_X1 U15147 ( .A1(n12809), .A2(n8496), .ZN(n12812) );
  OR2_X1 U15148 ( .A1(n12824), .A2(n12810), .ZN(n12811) );
  NAND2_X1 U15149 ( .A1(n12816), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n12814) );
  INV_X1 U15150 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n12948) );
  OR2_X1 U15151 ( .A1(n8516), .A2(n12948), .ZN(n12813) );
  OAI211_X1 U15152 ( .C1(n12820), .C2(n12815), .A(n12814), .B(n12813), .ZN(
        n13836) );
  NAND2_X1 U15153 ( .A1(n12911), .A2(n6437), .ZN(n12912) );
  INV_X1 U15154 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n12819) );
  NAND2_X1 U15155 ( .A1(n12816), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12818) );
  INV_X1 U15156 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n13921) );
  OR2_X1 U15157 ( .A1(n8516), .A2(n13921), .ZN(n12817) );
  OAI211_X1 U15158 ( .C1(n12820), .C2(n12819), .A(n12818), .B(n12817), .ZN(
        n13835) );
  AOI21_X1 U15159 ( .B1(n12728), .B2(n13835), .A(n11404), .ZN(n12821) );
  NAND3_X1 U15160 ( .A1(n12912), .A2(n12821), .A3(n12905), .ZN(n12822) );
  AOI22_X1 U15161 ( .A1(n12952), .A2(n6436), .B1(n13836), .B2(n12822), .ZN(
        n12848) );
  MUX2_X1 U15162 ( .A(n13836), .B(n12952), .S(n12728), .Z(n12847) );
  INV_X1 U15163 ( .A(n13837), .ZN(n12823) );
  MUX2_X1 U15164 ( .A(n12823), .B(n12968), .S(n6436), .Z(n12839) );
  OAI22_X1 U15165 ( .A1(n12848), .A2(n12847), .B1(n12839), .B2(n12838), .ZN(
        n12827) );
  NAND2_X1 U15166 ( .A1(n14244), .A2(n8496), .ZN(n12826) );
  OR2_X1 U15167 ( .A1(n12824), .A2(n14248), .ZN(n12825) );
  XNOR2_X1 U15168 ( .A(n14093), .B(n13835), .ZN(n12895) );
  NAND2_X1 U15169 ( .A1(n12827), .A2(n12895), .ZN(n12850) );
  MUX2_X1 U15170 ( .A(n13838), .B(n13000), .S(n6436), .Z(n12840) );
  MUX2_X1 U15171 ( .A(n13815), .B(n13937), .S(n12728), .Z(n12852) );
  MUX2_X1 U15172 ( .A(n13839), .B(n14115), .S(n6436), .Z(n12851) );
  AND2_X1 U15173 ( .A1(n12852), .A2(n12851), .ZN(n12829) );
  MUX2_X1 U15174 ( .A(n13840), .B(n14119), .S(n6436), .Z(n12835) );
  MUX2_X1 U15175 ( .A(n12830), .B(n13945), .S(n12728), .Z(n12834) );
  NAND2_X1 U15176 ( .A1(n12835), .A2(n12834), .ZN(n12831) );
  INV_X1 U15177 ( .A(n12833), .ZN(n12857) );
  INV_X1 U15178 ( .A(n12834), .ZN(n12837) );
  INV_X1 U15179 ( .A(n12835), .ZN(n12836) );
  NAND2_X1 U15180 ( .A1(n12837), .A2(n12836), .ZN(n12856) );
  INV_X1 U15181 ( .A(n12838), .ZN(n12846) );
  INV_X1 U15182 ( .A(n12839), .ZN(n12845) );
  INV_X1 U15183 ( .A(n12840), .ZN(n12843) );
  INV_X1 U15184 ( .A(n12841), .ZN(n12842) );
  NAND2_X1 U15185 ( .A1(n12843), .A2(n12842), .ZN(n12844) );
  OAI211_X1 U15186 ( .C1(n12846), .C2(n12845), .A(n12844), .B(n12895), .ZN(
        n12849) );
  AOI22_X1 U15187 ( .A1(n12850), .A2(n12849), .B1(n12848), .B2(n12847), .ZN(
        n12855) );
  OR3_X1 U15188 ( .A1(n12853), .A2(n12852), .A3(n12851), .ZN(n12854) );
  OAI211_X1 U15189 ( .C1(n12857), .C2(n12856), .A(n12855), .B(n12854), .ZN(
        n12858) );
  NAND2_X1 U15190 ( .A1(n6436), .A2(n13835), .ZN(n12861) );
  INV_X1 U15191 ( .A(n13835), .ZN(n12859) );
  NAND2_X1 U15192 ( .A1(n12728), .A2(n12859), .ZN(n12860) );
  MUX2_X1 U15193 ( .A(n12861), .B(n12860), .S(n14093), .Z(n12862) );
  NAND2_X1 U15194 ( .A1(n7586), .A2(n12864), .ZN(n13948) );
  INV_X1 U15195 ( .A(n13953), .ZN(n13951) );
  INV_X1 U15196 ( .A(n13963), .ZN(n12893) );
  INV_X1 U15197 ( .A(n12865), .ZN(n12867) );
  NAND2_X1 U15198 ( .A1(n12869), .A2(n12868), .ZN(n14022) );
  INV_X1 U15199 ( .A(n14045), .ZN(n14043) );
  AND4_X1 U15200 ( .A1(n12871), .A2(n6993), .A3(n12870), .A4(n10694), .ZN(
        n12874) );
  NAND3_X1 U15201 ( .A1(n12878), .A2(n12877), .A3(n12876), .ZN(n12879) );
  NOR2_X1 U15202 ( .A1(n12884), .A2(n12883), .ZN(n12887) );
  INV_X1 U15203 ( .A(n14073), .ZN(n12889) );
  NOR3_X1 U15204 ( .A1(n14016), .A2(n14022), .A3(n12890), .ZN(n12891) );
  XNOR2_X1 U15205 ( .A(n14163), .B(n13847), .ZN(n14039) );
  NAND4_X1 U15206 ( .A1(n13981), .A2(n12891), .A3(n13988), .A4(n14039), .ZN(
        n12892) );
  NOR4_X1 U15207 ( .A1(n13948), .A2(n13951), .A3(n12893), .A4(n12892), .ZN(
        n12894) );
  XNOR2_X1 U15208 ( .A(n12952), .B(n13836), .ZN(n12896) );
  XNOR2_X1 U15209 ( .A(n12897), .B(n13916), .ZN(n12898) );
  NAND2_X1 U15210 ( .A1(n12898), .A2(n11404), .ZN(n12915) );
  NAND2_X1 U15211 ( .A1(n13017), .A2(n12899), .ZN(n12900) );
  OAI211_X1 U15212 ( .C1(n6437), .C2(n12901), .A(n12905), .B(n12900), .ZN(
        n12902) );
  INV_X1 U15213 ( .A(n12902), .ZN(n12910) );
  NAND3_X1 U15214 ( .A1(n15459), .A2(n12903), .A3(n13801), .ZN(n12904) );
  OR2_X1 U15215 ( .A1(n12905), .A2(n12904), .ZN(n12909) );
  AOI21_X1 U15216 ( .B1(n12907), .B2(n12906), .A(n12949), .ZN(n12908) );
  NAND2_X1 U15217 ( .A1(n12909), .A2(n12908), .ZN(n12918) );
  OAI211_X1 U15218 ( .C1(n12915), .C2(n12911), .A(n12910), .B(n12918), .ZN(
        n12921) );
  OAI211_X1 U15219 ( .C1(n13017), .C2(n12913), .A(n12912), .B(n12918), .ZN(
        n12914) );
  INV_X1 U15220 ( .A(n12914), .ZN(n12916) );
  NAND3_X1 U15221 ( .A1(n12922), .A2(n12916), .A3(n12915), .ZN(n12920) );
  NAND2_X1 U15222 ( .A1(n12918), .A2(n12917), .ZN(n12919) );
  NAND2_X1 U15223 ( .A1(n13826), .A2(n12923), .ZN(n12924) );
  OAI211_X1 U15224 ( .C1(n15334), .C2(n12926), .A(n12925), .B(n12924), .ZN(
        n12932) );
  AOI22_X1 U15225 ( .A1(n13821), .A2(n13863), .B1(n13822), .B2(n12927), .ZN(
        n12929) );
  NOR3_X1 U15226 ( .A1(n12930), .A2(n12929), .A3(n12928), .ZN(n12931) );
  AOI211_X1 U15227 ( .C1(n12933), .C2(n15332), .A(n12932), .B(n12931), .ZN(
        n12934) );
  OAI21_X1 U15228 ( .B1(n12935), .B2(n15327), .A(n12934), .ZN(P2_U3199) );
  OAI222_X1 U15229 ( .A1(n15159), .A2(n12937), .B1(P1_U3086), .B2(n7780), .C1(
        n12936), .C2(n15165), .ZN(P1_U3325) );
  MUX2_X1 U15230 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n12938), .S(n15305), .Z(
        n12939) );
  INV_X1 U15231 ( .A(n12939), .ZN(n12942) );
  AOI22_X1 U15232 ( .A1(n15273), .A2(n12940), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n15301), .ZN(n12941) );
  OAI211_X1 U15233 ( .C1(n12943), .C2(n15279), .A(n12942), .B(n12941), .ZN(
        P1_U3291) );
  INV_X1 U15234 ( .A(n12944), .ZN(n14258) );
  OAI222_X1 U15235 ( .A1(n15165), .A2(n12945), .B1(n15159), .B2(n14258), .C1(
        n7809), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U15236 ( .A(n12967), .ZN(n12947) );
  INV_X1 U15237 ( .A(n12952), .ZN(n14098) );
  NOR2_X2 U15238 ( .A1(n12967), .A2(n12952), .ZN(n13919) );
  INV_X1 U15239 ( .A(n13919), .ZN(n12946) );
  OAI211_X1 U15240 ( .C1(n12947), .C2(n14098), .A(n12946), .B(n15443), .ZN(
        n14097) );
  NOR2_X1 U15241 ( .A1(n14064), .A2(n12948), .ZN(n12951) );
  OR2_X1 U15242 ( .A1(n10417), .A2(n12949), .ZN(n12950) );
  AND2_X1 U15243 ( .A1(n13802), .A2(n12950), .ZN(n12960) );
  NAND2_X1 U15244 ( .A1(n12960), .A2(n13835), .ZN(n14096) );
  NOR2_X1 U15245 ( .A1(n6438), .A2(n14096), .ZN(n13922) );
  AOI211_X1 U15246 ( .C1(n12952), .C2(n14085), .A(n12951), .B(n13922), .ZN(
        n12953) );
  OAI21_X1 U15247 ( .B1(n14097), .B2(n14089), .A(n12953), .ZN(P2_U3235) );
  INV_X1 U15248 ( .A(n15162), .ZN(n12954) );
  OAI222_X1 U15249 ( .A1(n14247), .A2(n12955), .B1(n13019), .B2(n12954), .C1(
        P2_U3088), .C2(n10417), .ZN(P2_U3300) );
  INV_X1 U15250 ( .A(n12956), .ZN(n12957) );
  XNOR2_X1 U15251 ( .A(n12959), .B(n14101), .ZN(n12964) );
  NAND2_X1 U15252 ( .A1(n12960), .A2(n13836), .ZN(n12961) );
  AND2_X1 U15253 ( .A1(n13000), .A2(n13838), .ZN(n14102) );
  AOI21_X1 U15254 ( .B1(n14109), .B2(n14104), .A(n14102), .ZN(n12966) );
  XNOR2_X1 U15255 ( .A(n12966), .B(n12965), .ZN(n12975) );
  INV_X1 U15256 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n12970) );
  OAI22_X1 U15257 ( .A1(n12971), .A2(n15434), .B1(n12970), .B2(n14064), .ZN(
        n12972) );
  AOI21_X1 U15258 ( .B1(n14100), .B2(n14085), .A(n12972), .ZN(n12973) );
  OAI21_X1 U15259 ( .B1(n14099), .B2(n14089), .A(n12973), .ZN(n12974) );
  AOI21_X1 U15260 ( .B1(n12975), .B2(n15446), .A(n12974), .ZN(n12976) );
  OAI21_X1 U15261 ( .B1(n14112), .B2(n6438), .A(n12976), .ZN(P2_U3236) );
  NAND2_X1 U15262 ( .A1(n13838), .A2(n9716), .ZN(n12982) );
  INV_X1 U15263 ( .A(n12982), .ZN(n12984) );
  OAI211_X1 U15264 ( .C1(n12979), .C2(n12983), .A(n12978), .B(n12982), .ZN(
        n12990) );
  INV_X1 U15265 ( .A(n12983), .ZN(n12980) );
  AOI21_X1 U15266 ( .B1(n12981), .B2(n12980), .A(n12984), .ZN(n12988) );
  MUX2_X1 U15267 ( .A(n12982), .B(n12981), .S(n12983), .Z(n12985) );
  AOI22_X1 U15268 ( .A1(n12987), .A2(n12985), .B1(n12984), .B2(n12983), .ZN(
        n12986) );
  OAI21_X1 U15269 ( .B1(n12988), .B2(n12987), .A(n12986), .ZN(n12989) );
  NAND3_X1 U15270 ( .A1(n12991), .A2(n12990), .A3(n12989), .ZN(n12995) );
  XNOR2_X1 U15271 ( .A(n12993), .B(n9726), .ZN(n12994) );
  XNOR2_X1 U15272 ( .A(n12995), .B(n12994), .ZN(n13003) );
  OAI22_X1 U15273 ( .A1(n12997), .A2(n15334), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12996), .ZN(n12998) );
  AOI21_X1 U15274 ( .B1(n12999), .B2(n13826), .A(n12998), .ZN(n13002) );
  NAND2_X1 U15275 ( .A1(n13000), .A2(n15332), .ZN(n13001) );
  OAI211_X1 U15276 ( .C1(n13003), .C2(n15327), .A(n13002), .B(n13001), .ZN(
        P2_U3192) );
  NAND2_X1 U15277 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n15406)
         );
  NAND2_X1 U15278 ( .A1(n13826), .A2(n13004), .ZN(n13005) );
  OAI211_X1 U15279 ( .C1(n15334), .C2(n13006), .A(n15406), .B(n13005), .ZN(
        n13014) );
  INV_X1 U15280 ( .A(n13007), .ZN(n13781) );
  NOR3_X1 U15281 ( .A1(n13009), .A2(n13008), .A3(n13790), .ZN(n13010) );
  AOI21_X1 U15282 ( .B1(n13781), .B2(n13822), .A(n13010), .ZN(n13012) );
  NOR2_X1 U15283 ( .A1(n13012), .A2(n13011), .ZN(n13013) );
  AOI211_X1 U15284 ( .C1(n14201), .C2(n15332), .A(n13014), .B(n13013), .ZN(
        n13015) );
  OAI21_X1 U15285 ( .B1(n13016), .B2(n15327), .A(n13015), .ZN(P2_U3187) );
  OAI222_X1 U15286 ( .A1(n14247), .A2(n13020), .B1(n13019), .B2(n13018), .C1(
        P2_U3088), .C2(n13017), .ZN(P2_U3308) );
  XNOR2_X1 U15287 ( .A(n13374), .B(n13071), .ZN(n13068) );
  XNOR2_X1 U15288 ( .A(n13068), .B(n13204), .ZN(n13069) );
  XNOR2_X1 U15289 ( .A(n13673), .B(n13035), .ZN(n13107) );
  INV_X1 U15290 ( .A(n13107), .ZN(n13026) );
  INV_X1 U15291 ( .A(n13021), .ZN(n13022) );
  XNOR2_X1 U15292 ( .A(n13679), .B(n13071), .ZN(n13025) );
  XNOR2_X1 U15293 ( .A(n13025), .B(n13113), .ZN(n13188) );
  XNOR2_X1 U15294 ( .A(n13667), .B(n6431), .ZN(n13028) );
  XNOR2_X1 U15295 ( .A(n13028), .B(n13525), .ZN(n13118) );
  NAND2_X1 U15296 ( .A1(n13119), .A2(n13118), .ZN(n13117) );
  NAND2_X1 U15297 ( .A1(n13117), .A2(n13029), .ZN(n13172) );
  XNOR2_X1 U15298 ( .A(n13661), .B(n13071), .ZN(n13030) );
  XNOR2_X1 U15299 ( .A(n13030), .B(n13515), .ZN(n13171) );
  XNOR2_X1 U15300 ( .A(n13655), .B(n13071), .ZN(n13032) );
  XNOR2_X1 U15301 ( .A(n13032), .B(n13473), .ZN(n13060) );
  XNOR2_X1 U15302 ( .A(n13594), .B(n13071), .ZN(n13033) );
  XNOR2_X1 U15303 ( .A(n13033), .B(n13487), .ZN(n13138) );
  NAND2_X1 U15304 ( .A1(n13139), .A2(n13138), .ZN(n13137) );
  XNOR2_X1 U15305 ( .A(n13645), .B(n13071), .ZN(n13036) );
  XNOR2_X1 U15306 ( .A(n13036), .B(n13474), .ZN(n13094) );
  XNOR2_X1 U15307 ( .A(n13639), .B(n13035), .ZN(n13147) );
  NAND2_X1 U15308 ( .A1(n13036), .A2(n13474), .ZN(n13146) );
  OAI21_X1 U15309 ( .B1(n13147), .B2(n13457), .A(n13146), .ZN(n13038) );
  INV_X1 U15310 ( .A(n13147), .ZN(n13037) );
  XNOR2_X1 U15311 ( .A(n13577), .B(n6431), .ZN(n13129) );
  XNOR2_X1 U15312 ( .A(n13582), .B(n6431), .ZN(n13039) );
  OAI22_X1 U15313 ( .A1(n13129), .A2(n13428), .B1(n13417), .B2(n13039), .ZN(
        n13043) );
  NAND3_X1 U15314 ( .A1(n13039), .A2(n13417), .A3(n13428), .ZN(n13042) );
  INV_X1 U15315 ( .A(n13039), .ZN(n13127) );
  OAI21_X1 U15316 ( .B1(n13127), .B2(n13447), .A(n13206), .ZN(n13040) );
  NAND2_X1 U15317 ( .A1(n13129), .A2(n13040), .ZN(n13041) );
  XNOR2_X1 U15318 ( .A(n13403), .B(n6431), .ZN(n13044) );
  XNOR2_X1 U15319 ( .A(n13044), .B(n13385), .ZN(n13101) );
  XNOR2_X1 U15320 ( .A(n13572), .B(n13071), .ZN(n13046) );
  XNOR2_X1 U15321 ( .A(n13046), .B(n13045), .ZN(n13180) );
  XOR2_X1 U15322 ( .A(n13069), .B(n13070), .Z(n13052) );
  NOR2_X1 U15323 ( .A1(n13184), .A2(n13371), .ZN(n13050) );
  AOI22_X1 U15324 ( .A1(n13190), .A2(n13205), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13047) );
  OAI21_X1 U15325 ( .B1(n13048), .B2(n13193), .A(n13047), .ZN(n13049) );
  AOI211_X1 U15326 ( .C1(n13374), .C2(n13196), .A(n13050), .B(n13049), .ZN(
        n13051) );
  OAI21_X1 U15327 ( .B1(n13052), .B2(n13199), .A(n13051), .ZN(P3_U3154) );
  XNOR2_X1 U15328 ( .A(n13126), .B(n13127), .ZN(n13128) );
  XNOR2_X1 U15329 ( .A(n13128), .B(n13417), .ZN(n13058) );
  INV_X1 U15330 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n13053) );
  OAI22_X1 U15331 ( .A1(n13193), .A2(n13428), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13053), .ZN(n13055) );
  NOR2_X1 U15332 ( .A1(n13429), .A2(n13151), .ZN(n13054) );
  AOI211_X1 U15333 ( .C1(n13436), .C2(n13195), .A(n13055), .B(n13054), .ZN(
        n13057) );
  NAND2_X1 U15334 ( .A1(n13582), .A2(n13196), .ZN(n13056) );
  OAI211_X1 U15335 ( .C1(n13058), .C2(n13199), .A(n13057), .B(n13056), .ZN(
        P3_U3156) );
  OAI211_X1 U15336 ( .C1(n13061), .C2(n13060), .A(n13059), .B(n13169), .ZN(
        n13067) );
  NAND2_X1 U15337 ( .A1(n13190), .A2(n13515), .ZN(n13063) );
  OAI211_X1 U15338 ( .C1(n13064), .C2(n13193), .A(n13063), .B(n13062), .ZN(
        n13065) );
  AOI21_X1 U15339 ( .B1(n13493), .B2(n13195), .A(n13065), .ZN(n13066) );
  OAI211_X1 U15340 ( .C1(n13177), .C2(n13655), .A(n13067), .B(n13066), .ZN(
        P3_U3159) );
  AOI22_X1 U15341 ( .A1(n13190), .A2(n13204), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13076) );
  NAND2_X1 U15342 ( .A1(n13195), .A2(n13074), .ZN(n13075) );
  OAI211_X1 U15343 ( .C1(n13077), .C2(n13193), .A(n13076), .B(n13075), .ZN(
        n13078) );
  AOI21_X1 U15344 ( .B1(n13079), .B2(n13196), .A(n13078), .ZN(n13080) );
  MUX2_X1 U15345 ( .A(n13210), .B(n13082), .S(n13081), .Z(n13084) );
  XNOR2_X1 U15346 ( .A(n13084), .B(n13083), .ZN(n13085) );
  NAND2_X1 U15347 ( .A1(n13085), .A2(n13169), .ZN(n13092) );
  AOI21_X1 U15348 ( .B1(n13196), .B2(n13087), .A(n13086), .ZN(n13091) );
  AOI22_X1 U15349 ( .A1(n13181), .A2(n13208), .B1(n13190), .B2(n13210), .ZN(
        n13090) );
  NAND2_X1 U15350 ( .A1(n13195), .A2(n13088), .ZN(n13089) );
  NAND4_X1 U15351 ( .A1(n13092), .A2(n13091), .A3(n13090), .A4(n13089), .ZN(
        P3_U3161) );
  AOI21_X1 U15352 ( .B1(n13094), .B2(n13093), .A(n13145), .ZN(n13099) );
  AOI22_X1 U15353 ( .A1(n13487), .A2(n13190), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13096) );
  NAND2_X1 U15354 ( .A1(n13195), .A2(n13460), .ZN(n13095) );
  OAI211_X1 U15355 ( .C1(n13429), .C2(n13193), .A(n13096), .B(n13095), .ZN(
        n13097) );
  AOI21_X1 U15356 ( .B1(n13645), .B2(n13196), .A(n13097), .ZN(n13098) );
  OAI21_X1 U15357 ( .B1(n13099), .B2(n13199), .A(n13098), .ZN(P3_U3163) );
  XOR2_X1 U15358 ( .A(n13101), .B(n13100), .Z(n13106) );
  AOI22_X1 U15359 ( .A1(n13181), .A2(n13205), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13103) );
  NAND2_X1 U15360 ( .A1(n13190), .A2(n13206), .ZN(n13102) );
  OAI211_X1 U15361 ( .C1(n13184), .C2(n13400), .A(n13103), .B(n13102), .ZN(
        n13104) );
  AOI21_X1 U15362 ( .B1(n13403), .B2(n13196), .A(n13104), .ZN(n13105) );
  OAI21_X1 U15363 ( .B1(n13106), .B2(n13199), .A(n13105), .ZN(P3_U3165) );
  XNOR2_X1 U15364 ( .A(n13107), .B(n13192), .ZN(n13108) );
  XNOR2_X1 U15365 ( .A(n13109), .B(n13108), .ZN(n13116) );
  NOR2_X1 U15366 ( .A1(n13110), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13314) );
  AOI21_X1 U15367 ( .B1(n13181), .B2(n13525), .A(n13314), .ZN(n13112) );
  NAND2_X1 U15368 ( .A1(n13195), .A2(n13528), .ZN(n13111) );
  OAI211_X1 U15369 ( .C1(n13113), .C2(n13151), .A(n13112), .B(n13111), .ZN(
        n13114) );
  AOI21_X1 U15370 ( .B1(n13673), .B2(n13196), .A(n13114), .ZN(n13115) );
  OAI21_X1 U15371 ( .B1(n13116), .B2(n13199), .A(n13115), .ZN(P3_U3166) );
  INV_X1 U15372 ( .A(n13667), .ZN(n13125) );
  OAI211_X1 U15373 ( .C1(n13119), .C2(n13118), .A(n13117), .B(n13169), .ZN(
        n13124) );
  NOR2_X1 U15374 ( .A1(n13120), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13331) );
  AOI21_X1 U15375 ( .B1(n13181), .B2(n13515), .A(n13331), .ZN(n13121) );
  OAI21_X1 U15376 ( .B1(n13192), .B2(n13151), .A(n13121), .ZN(n13122) );
  AOI21_X1 U15377 ( .B1(n13518), .B2(n13195), .A(n13122), .ZN(n13123) );
  OAI211_X1 U15378 ( .C1(n13125), .C2(n13177), .A(n13124), .B(n13123), .ZN(
        P3_U3168) );
  OAI22_X1 U15379 ( .A1(n13128), .A2(n13447), .B1(n13127), .B2(n13126), .ZN(
        n13131) );
  XNOR2_X1 U15380 ( .A(n13129), .B(n13428), .ZN(n13130) );
  XNOR2_X1 U15381 ( .A(n13131), .B(n13130), .ZN(n13136) );
  OAI22_X1 U15382 ( .A1(n13193), .A2(n13416), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n6908), .ZN(n13132) );
  AOI21_X1 U15383 ( .B1(n13447), .B2(n13190), .A(n13132), .ZN(n13133) );
  OAI21_X1 U15384 ( .B1(n13420), .B2(n13184), .A(n13133), .ZN(n13134) );
  AOI21_X1 U15385 ( .B1(n13577), .B2(n13196), .A(n13134), .ZN(n13135) );
  OAI21_X1 U15386 ( .B1(n13136), .B2(n13199), .A(n13135), .ZN(P3_U3169) );
  INV_X1 U15387 ( .A(n13594), .ZN(n13144) );
  OAI211_X1 U15388 ( .C1(n13139), .C2(n13138), .A(n13137), .B(n13169), .ZN(
        n13143) );
  AOI22_X1 U15389 ( .A1(n13446), .A2(n13181), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13140) );
  OAI21_X1 U15390 ( .B1(n13473), .B2(n13151), .A(n13140), .ZN(n13141) );
  AOI21_X1 U15391 ( .B1(n13475), .B2(n13195), .A(n13141), .ZN(n13142) );
  OAI211_X1 U15392 ( .C1(n13144), .C2(n13177), .A(n13143), .B(n13142), .ZN(
        P3_U3173) );
  NAND2_X1 U15393 ( .A1(n7369), .A2(n13146), .ZN(n13149) );
  XNOR2_X1 U15394 ( .A(n13147), .B(n13457), .ZN(n13148) );
  XNOR2_X1 U15395 ( .A(n13149), .B(n13148), .ZN(n13156) );
  INV_X1 U15396 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13150) );
  OAI22_X1 U15397 ( .A1(n13474), .A2(n13151), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13150), .ZN(n13153) );
  NOR2_X1 U15398 ( .A1(n13417), .A2(n13193), .ZN(n13152) );
  AOI211_X1 U15399 ( .C1(n13450), .C2(n13195), .A(n13153), .B(n13152), .ZN(
        n13155) );
  NAND2_X1 U15400 ( .A1(n13639), .A2(n13196), .ZN(n13154) );
  OAI211_X1 U15401 ( .C1(n13156), .C2(n13199), .A(n13155), .B(n13154), .ZN(
        P3_U3175) );
  XNOR2_X1 U15402 ( .A(n13158), .B(n13157), .ZN(n13159) );
  NAND2_X1 U15403 ( .A1(n13159), .A2(n13169), .ZN(n13168) );
  NAND2_X1 U15404 ( .A1(n13190), .A2(n13207), .ZN(n13160) );
  NAND2_X1 U15405 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n13221)
         );
  OAI211_X1 U15406 ( .C1(n13193), .C2(n13161), .A(n13160), .B(n13221), .ZN(
        n13162) );
  INV_X1 U15407 ( .A(n13162), .ZN(n13167) );
  NAND2_X1 U15408 ( .A1(n13195), .A2(n13163), .ZN(n13166) );
  NAND2_X1 U15409 ( .A1(n13196), .A2(n13164), .ZN(n13165) );
  NAND4_X1 U15410 ( .A1(n13168), .A2(n13167), .A3(n13166), .A4(n13165), .ZN(
        P3_U3176) );
  OAI211_X1 U15411 ( .C1(n13172), .C2(n13171), .A(n13170), .B(n13169), .ZN(
        n13176) );
  NAND2_X1 U15412 ( .A1(n13190), .A2(n13525), .ZN(n13173) );
  NAND2_X1 U15413 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13353)
         );
  OAI211_X1 U15414 ( .C1(n13193), .C2(n13473), .A(n13173), .B(n13353), .ZN(
        n13174) );
  AOI21_X1 U15415 ( .B1(n13507), .B2(n13195), .A(n13174), .ZN(n13175) );
  OAI211_X1 U15416 ( .C1(n13178), .C2(n13177), .A(n13176), .B(n13175), .ZN(
        P3_U3178) );
  XOR2_X1 U15417 ( .A(n13180), .B(n13179), .Z(n13187) );
  AOI22_X1 U15418 ( .A1(n13181), .A2(n13204), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13183) );
  NAND2_X1 U15419 ( .A1(n13190), .A2(n13385), .ZN(n13182) );
  OAI211_X1 U15420 ( .C1(n13184), .C2(n13394), .A(n13183), .B(n13182), .ZN(
        n13185) );
  AOI21_X1 U15421 ( .B1(n13572), .B2(n13196), .A(n13185), .ZN(n13186) );
  OAI21_X1 U15422 ( .B1(n13187), .B2(n13199), .A(n13186), .ZN(P3_U3180) );
  XNOR2_X1 U15423 ( .A(n13189), .B(n13188), .ZN(n13200) );
  NAND2_X1 U15424 ( .A1(n13190), .A2(n13559), .ZN(n13191) );
  NAND2_X1 U15425 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13294)
         );
  OAI211_X1 U15426 ( .C1(n13193), .C2(n13192), .A(n13191), .B(n13294), .ZN(
        n13194) );
  AOI21_X1 U15427 ( .B1(n13539), .B2(n13195), .A(n13194), .ZN(n13198) );
  NAND2_X1 U15428 ( .A1(n13679), .A2(n13196), .ZN(n13197) );
  OAI211_X1 U15429 ( .C1(n13200), .C2(n13199), .A(n13198), .B(n13197), .ZN(
        P3_U3181) );
  MUX2_X1 U15430 ( .A(n13201), .B(P3_DATAO_REG_31__SCAN_IN), .S(n13214), .Z(
        P3_U3522) );
  MUX2_X1 U15431 ( .A(n13202), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13214), .Z(
        P3_U3521) );
  MUX2_X1 U15432 ( .A(n13203), .B(P3_DATAO_REG_28__SCAN_IN), .S(n13214), .Z(
        P3_U3519) );
  MUX2_X1 U15433 ( .A(n13204), .B(P3_DATAO_REG_27__SCAN_IN), .S(n13214), .Z(
        P3_U3518) );
  MUX2_X1 U15434 ( .A(n13205), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13214), .Z(
        P3_U3517) );
  MUX2_X1 U15435 ( .A(n13385), .B(P3_DATAO_REG_25__SCAN_IN), .S(n13214), .Z(
        P3_U3516) );
  MUX2_X1 U15436 ( .A(n13206), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13214), .Z(
        P3_U3515) );
  MUX2_X1 U15437 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13447), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U15438 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13457), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15439 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13446), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15440 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13487), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15441 ( .A(n13504), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13214), .Z(
        P3_U3510) );
  MUX2_X1 U15442 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13515), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15443 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13525), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15444 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13536), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15445 ( .A(n13547), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13214), .Z(
        P3_U3506) );
  MUX2_X1 U15446 ( .A(n13559), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13214), .Z(
        P3_U3505) );
  MUX2_X1 U15447 ( .A(n13546), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13214), .Z(
        P3_U3504) );
  MUX2_X1 U15448 ( .A(n13558), .B(P3_DATAO_REG_12__SCAN_IN), .S(n13214), .Z(
        P3_U3503) );
  MUX2_X1 U15449 ( .A(n13207), .B(P3_DATAO_REG_10__SCAN_IN), .S(n13214), .Z(
        P3_U3501) );
  MUX2_X1 U15450 ( .A(n13208), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13214), .Z(
        P3_U3500) );
  MUX2_X1 U15451 ( .A(n13209), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13214), .Z(
        P3_U3499) );
  MUX2_X1 U15452 ( .A(n13210), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13214), .Z(
        P3_U3498) );
  MUX2_X1 U15453 ( .A(n13211), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13214), .Z(
        P3_U3497) );
  MUX2_X1 U15454 ( .A(n13212), .B(P3_DATAO_REG_5__SCAN_IN), .S(n13214), .Z(
        P3_U3496) );
  MUX2_X1 U15455 ( .A(n13213), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13214), .Z(
        P3_U3495) );
  MUX2_X1 U15456 ( .A(n15532), .B(P3_DATAO_REG_3__SCAN_IN), .S(n13214), .Z(
        P3_U3494) );
  MUX2_X1 U15457 ( .A(n15544), .B(P3_DATAO_REG_2__SCAN_IN), .S(n13214), .Z(
        P3_U3493) );
  MUX2_X1 U15458 ( .A(n15533), .B(P3_DATAO_REG_1__SCAN_IN), .S(n13214), .Z(
        P3_U3492) );
  MUX2_X1 U15459 ( .A(n15545), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13214), .Z(
        P3_U3491) );
  OAI21_X1 U15460 ( .B1(n13216), .B2(P3_REG1_REG_11__SCAN_IN), .A(n13215), 
        .ZN(n13217) );
  NAND2_X1 U15461 ( .A1(n13217), .A2(n9642), .ZN(n13229) );
  OAI21_X1 U15462 ( .B1(n13219), .B2(n13218), .A(n13238), .ZN(n13224) );
  NAND2_X1 U15463 ( .A1(n15503), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n13220) );
  OAI211_X1 U15464 ( .C1(n13355), .C2(n13222), .A(n13221), .B(n13220), .ZN(
        n13223) );
  AOI21_X1 U15465 ( .B1(n13224), .B2(n13270), .A(n13223), .ZN(n13228) );
  OAI21_X1 U15466 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n13225), .A(n13232), 
        .ZN(n13226) );
  NAND2_X1 U15467 ( .A1(n13226), .A2(n13348), .ZN(n13227) );
  NAND3_X1 U15468 ( .A1(n13229), .A2(n13228), .A3(n13227), .ZN(P3_U3193) );
  AND3_X1 U15469 ( .A1(n13232), .A2(n13231), .A3(n13230), .ZN(n13233) );
  OAI21_X1 U15470 ( .B1(n13234), .B2(n13233), .A(n13348), .ZN(n13250) );
  INV_X1 U15471 ( .A(n15503), .ZN(n13297) );
  OAI21_X1 U15472 ( .B1(n13297), .B2(n15180), .A(n13235), .ZN(n13242) );
  INV_X1 U15473 ( .A(n13255), .ZN(n13240) );
  AOI21_X1 U15474 ( .B1(n13238), .B2(n13237), .A(n13236), .ZN(n13239) );
  NOR3_X1 U15475 ( .A1(n13240), .A2(n13239), .A3(n13359), .ZN(n13241) );
  AOI211_X1 U15476 ( .C1(n13339), .C2(n13243), .A(n13242), .B(n13241), .ZN(
        n13249) );
  OAI21_X1 U15477 ( .B1(n13246), .B2(n13245), .A(n13244), .ZN(n13247) );
  NAND2_X1 U15478 ( .A1(n13247), .A2(n9642), .ZN(n13248) );
  NAND3_X1 U15479 ( .A1(n13250), .A2(n13249), .A3(n13248), .ZN(P3_U3194) );
  AOI21_X1 U15480 ( .B1(n13561), .B2(n13251), .A(n13273), .ZN(n13266) );
  INV_X1 U15481 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15184) );
  OAI21_X1 U15482 ( .B1(n13297), .B2(n15184), .A(n13252), .ZN(n13259) );
  AOI21_X1 U15483 ( .B1(n13255), .B2(n13254), .A(n13253), .ZN(n13256) );
  INV_X1 U15484 ( .A(n13256), .ZN(n13257) );
  AOI21_X1 U15485 ( .B1(n13257), .B2(n13269), .A(n13359), .ZN(n13258) );
  AOI211_X1 U15486 ( .C1(n13339), .C2(n13260), .A(n13259), .B(n13258), .ZN(
        n13265) );
  OAI21_X1 U15487 ( .B1(n13262), .B2(P3_REG1_REG_13__SCAN_IN), .A(n13261), 
        .ZN(n13263) );
  NAND2_X1 U15488 ( .A1(n13263), .A2(n9642), .ZN(n13264) );
  OAI211_X1 U15489 ( .C1(n13266), .C2(n13341), .A(n13265), .B(n13264), .ZN(
        P3_U3195) );
  AOI21_X1 U15490 ( .B1(n13269), .B2(n13268), .A(n13267), .ZN(n13290) );
  NAND2_X1 U15491 ( .A1(n13271), .A2(n13270), .ZN(n13289) );
  INV_X1 U15492 ( .A(n13272), .ZN(n13277) );
  NOR3_X1 U15493 ( .A1(n13275), .A2(n13274), .A3(n13273), .ZN(n13276) );
  OAI21_X1 U15494 ( .B1(n13277), .B2(n13276), .A(n13348), .ZN(n13288) );
  OAI21_X1 U15495 ( .B1(n13280), .B2(n13279), .A(n13278), .ZN(n13281) );
  INV_X1 U15496 ( .A(n13281), .ZN(n13284) );
  NAND2_X1 U15497 ( .A1(n15503), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n13282) );
  OAI211_X1 U15498 ( .C1(n13333), .C2(n13284), .A(n13283), .B(n13282), .ZN(
        n13285) );
  AOI21_X1 U15499 ( .B1(n13286), .B2(n13339), .A(n13285), .ZN(n13287) );
  OAI211_X1 U15500 ( .C1(n13290), .C2(n13289), .A(n13288), .B(n13287), .ZN(
        P3_U3196) );
  INV_X1 U15501 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13296) );
  OAI21_X1 U15502 ( .B1(n13292), .B2(P3_REG1_REG_15__SCAN_IN), .A(n13291), 
        .ZN(n13293) );
  NAND2_X1 U15503 ( .A1(n9642), .A2(n13293), .ZN(n13295) );
  OAI211_X1 U15504 ( .C1(n13297), .C2(n13296), .A(n13295), .B(n13294), .ZN(
        n13303) );
  AOI21_X1 U15505 ( .B1(n13300), .B2(n13299), .A(n13298), .ZN(n13301) );
  NOR2_X1 U15506 ( .A1(n13301), .A2(n13359), .ZN(n13302) );
  AOI211_X1 U15507 ( .C1(n13339), .C2(n13304), .A(n13303), .B(n13302), .ZN(
        n13305) );
  OAI21_X1 U15508 ( .B1(n13306), .B2(n13341), .A(n13305), .ZN(P3_U3197) );
  OAI21_X1 U15509 ( .B1(n13309), .B2(n13308), .A(n13307), .ZN(n13326) );
  INV_X1 U15510 ( .A(n13310), .ZN(n13311) );
  NOR2_X1 U15511 ( .A1(n13312), .A2(n13311), .ZN(n13313) );
  XNOR2_X1 U15512 ( .A(n6594), .B(n13313), .ZN(n13318) );
  AOI21_X1 U15513 ( .B1(n15503), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13314), 
        .ZN(n13317) );
  NAND2_X1 U15514 ( .A1(n13339), .A2(n13315), .ZN(n13316) );
  OAI211_X1 U15515 ( .C1(n13318), .C2(n13359), .A(n13317), .B(n13316), .ZN(
        n13325) );
  OR3_X1 U15516 ( .A1(n13321), .A2(n13320), .A3(n13319), .ZN(n13322) );
  AOI21_X1 U15517 ( .B1(n13323), .B2(n13322), .A(n13341), .ZN(n13324) );
  AOI211_X1 U15518 ( .C1(n9642), .C2(n13326), .A(n13325), .B(n13324), .ZN(
        n13327) );
  INV_X1 U15519 ( .A(n13327), .ZN(P3_U3198) );
  AOI21_X1 U15520 ( .B1(n13517), .B2(n13329), .A(n13328), .ZN(n13342) );
  AOI21_X1 U15521 ( .B1(n15503), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13331), 
        .ZN(n13332) );
  AOI211_X1 U15522 ( .C1(n13336), .C2(n13335), .A(n13359), .B(n13334), .ZN(
        n13337) );
  OAI21_X1 U15523 ( .B1(n13342), .B2(n13341), .A(n13340), .ZN(P3_U3199) );
  AOI21_X1 U15524 ( .B1(n13345), .B2(n13344), .A(n13343), .ZN(n13360) );
  NOR3_X1 U15525 ( .A1(n13328), .A2(n13347), .A3(n13346), .ZN(n13349) );
  XNOR2_X1 U15526 ( .A(n13351), .B(n13350), .ZN(n13357) );
  NAND2_X1 U15527 ( .A1(n15503), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13352) );
  OAI211_X1 U15528 ( .C1(n13355), .C2(n13354), .A(n13353), .B(n13352), .ZN(
        n13356) );
  AOI21_X1 U15529 ( .B1(n9642), .B2(n13357), .A(n13356), .ZN(n13358) );
  NAND2_X1 U15530 ( .A1(n13361), .A2(n6428), .ZN(n13365) );
  NOR2_X1 U15531 ( .A1(n13363), .A2(n13362), .ZN(n13621) );
  OAI21_X1 U15532 ( .B1(n13364), .B2(n13621), .A(n15559), .ZN(n13367) );
  OAI211_X1 U15533 ( .C1(n15559), .C2(n13366), .A(n13365), .B(n13367), .ZN(
        P3_U3202) );
  NAND2_X1 U15534 ( .A1(n15561), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13368) );
  OAI211_X1 U15535 ( .C1(n13571), .C2(n13495), .A(n13368), .B(n13367), .ZN(
        P3_U3203) );
  INV_X1 U15536 ( .A(n13369), .ZN(n13377) );
  NAND2_X1 U15537 ( .A1(n13370), .A2(n15559), .ZN(n13376) );
  OAI22_X1 U15538 ( .A1(n15559), .A2(n13372), .B1(n13371), .B2(n15553), .ZN(
        n13373) );
  AOI21_X1 U15539 ( .B1(n13374), .B2(n6428), .A(n13373), .ZN(n13375) );
  OAI211_X1 U15540 ( .C1(n13377), .C2(n15555), .A(n13376), .B(n13375), .ZN(
        P3_U3206) );
  NAND2_X1 U15541 ( .A1(n13425), .A2(n13378), .ZN(n13381) );
  INV_X1 U15542 ( .A(n13379), .ZN(n13380) );
  NAND2_X1 U15543 ( .A1(n13381), .A2(n13380), .ZN(n13383) );
  NAND2_X1 U15544 ( .A1(n13383), .A2(n13382), .ZN(n13384) );
  NAND2_X1 U15545 ( .A1(n13385), .A2(n15546), .ZN(n13386) );
  OAI21_X1 U15546 ( .B1(n13387), .B2(n15510), .A(n13386), .ZN(n13388) );
  AOI21_X1 U15547 ( .B1(n13573), .B2(n13435), .A(n13388), .ZN(n13393) );
  XNOR2_X1 U15548 ( .A(n13390), .B(n13389), .ZN(n13391) );
  NAND2_X1 U15549 ( .A1(n13391), .A2(n10147), .ZN(n13392) );
  OAI22_X1 U15550 ( .A1(n15559), .A2(n13395), .B1(n13394), .B2(n15553), .ZN(
        n13396) );
  AOI21_X1 U15551 ( .B1(n13572), .B2(n6428), .A(n13396), .ZN(n13398) );
  NAND2_X1 U15552 ( .A1(n13573), .A2(n13440), .ZN(n13397) );
  OAI211_X1 U15553 ( .C1(n13575), .C2(n15561), .A(n13398), .B(n13397), .ZN(
        P3_U3207) );
  NAND2_X1 U15554 ( .A1(n13399), .A2(n15559), .ZN(n13405) );
  INV_X1 U15555 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n13401) );
  OAI22_X1 U15556 ( .A1(n15559), .A2(n13401), .B1(n13400), .B2(n15553), .ZN(
        n13402) );
  AOI21_X1 U15557 ( .B1(n13403), .B2(n6428), .A(n13402), .ZN(n13404) );
  OAI211_X1 U15558 ( .C1(n13406), .C2(n15555), .A(n13405), .B(n13404), .ZN(
        P3_U3208) );
  INV_X1 U15559 ( .A(n13427), .ZN(n13409) );
  OAI21_X1 U15560 ( .B1(n13409), .B2(n13408), .A(n13407), .ZN(n13410) );
  NAND2_X1 U15561 ( .A1(n13411), .A2(n13410), .ZN(n13578) );
  NAND2_X1 U15562 ( .A1(n13413), .A2(n13412), .ZN(n13414) );
  OAI22_X1 U15563 ( .A1(n13417), .A2(n15508), .B1(n13416), .B2(n15510), .ZN(
        n13418) );
  AOI211_X1 U15564 ( .C1(n13578), .C2(n13435), .A(n13419), .B(n13418), .ZN(
        n13580) );
  INV_X1 U15565 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n13421) );
  OAI22_X1 U15566 ( .A1(n15559), .A2(n13421), .B1(n13420), .B2(n15553), .ZN(
        n13422) );
  AOI21_X1 U15567 ( .B1(n13577), .B2(n6428), .A(n13422), .ZN(n13424) );
  NAND2_X1 U15568 ( .A1(n13578), .A2(n13440), .ZN(n13423) );
  OAI211_X1 U15569 ( .C1(n13580), .C2(n15561), .A(n13424), .B(n13423), .ZN(
        P3_U3209) );
  OR2_X1 U15570 ( .A1(n13425), .A2(n7635), .ZN(n13426) );
  OAI22_X1 U15571 ( .A1(n13429), .A2(n15508), .B1(n13428), .B2(n15510), .ZN(
        n13434) );
  INV_X1 U15572 ( .A(n13430), .ZN(n13431) );
  AOI211_X1 U15573 ( .C1(n7635), .C2(n13432), .A(n13472), .B(n13431), .ZN(
        n13433) );
  NAND2_X1 U15574 ( .A1(n13582), .A2(n6428), .ZN(n13438) );
  AOI22_X1 U15575 ( .A1(n13436), .A2(n15518), .B1(n15561), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13437) );
  NAND2_X1 U15576 ( .A1(n13438), .A2(n13437), .ZN(n13439) );
  AOI21_X1 U15577 ( .B1(n13581), .B2(n13440), .A(n13439), .ZN(n13441) );
  OAI21_X1 U15578 ( .B1(n13584), .B2(n15561), .A(n13441), .ZN(P3_U3210) );
  XNOR2_X1 U15579 ( .A(n13442), .B(n13443), .ZN(n13642) );
  XNOR2_X1 U15580 ( .A(n13445), .B(n13444), .ZN(n13448) );
  AOI222_X1 U15581 ( .A1(n10147), .A2(n13448), .B1(n13447), .B2(n15543), .C1(
        n13446), .C2(n15546), .ZN(n13637) );
  MUX2_X1 U15582 ( .A(n13449), .B(n13637), .S(n15559), .Z(n13452) );
  AOI22_X1 U15583 ( .A1(n13639), .A2(n6428), .B1(n15518), .B2(n13450), .ZN(
        n13451) );
  OAI211_X1 U15584 ( .C1(n13642), .C2(n13566), .A(n13452), .B(n13451), .ZN(
        P3_U3211) );
  XNOR2_X1 U15585 ( .A(n13454), .B(n13453), .ZN(n13648) );
  INV_X1 U15586 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13459) );
  OAI21_X1 U15587 ( .B1(n13456), .B2(n9299), .A(n13455), .ZN(n13458) );
  AOI222_X1 U15588 ( .A1(n10147), .A2(n13458), .B1(n13457), .B2(n15543), .C1(
        n13487), .C2(n15546), .ZN(n13643) );
  MUX2_X1 U15589 ( .A(n13459), .B(n13643), .S(n15559), .Z(n13462) );
  AOI22_X1 U15590 ( .A1(n13645), .A2(n6428), .B1(n15518), .B2(n13460), .ZN(
        n13461) );
  OAI211_X1 U15591 ( .C1(n13648), .C2(n13566), .A(n13462), .B(n13461), .ZN(
        P3_U3212) );
  OAI21_X1 U15592 ( .B1(n13464), .B2(n13465), .A(n13463), .ZN(n13652) );
  NOR2_X1 U15593 ( .A1(n13466), .A2(n9481), .ZN(n13500) );
  OR2_X1 U15594 ( .A1(n13500), .A2(n13467), .ZN(n13484) );
  NAND2_X1 U15595 ( .A1(n13484), .A2(n13468), .ZN(n13469) );
  XNOR2_X1 U15596 ( .A(n13470), .B(n13469), .ZN(n13471) );
  OAI222_X1 U15597 ( .A1(n15510), .A2(n13474), .B1(n15508), .B2(n13473), .C1(
        n13472), .C2(n13471), .ZN(n13593) );
  NAND2_X1 U15598 ( .A1(n13593), .A2(n15559), .ZN(n13480) );
  INV_X1 U15599 ( .A(n13475), .ZN(n13476) );
  OAI22_X1 U15600 ( .A1(n15559), .A2(n13477), .B1(n13476), .B2(n15553), .ZN(
        n13478) );
  AOI21_X1 U15601 ( .B1(n13594), .B2(n6428), .A(n13478), .ZN(n13479) );
  OAI211_X1 U15602 ( .C1(n13652), .C2(n13566), .A(n13480), .B(n13479), .ZN(
        P3_U3213) );
  XOR2_X1 U15603 ( .A(n13481), .B(n13485), .Z(n13656) );
  INV_X1 U15604 ( .A(n13482), .ZN(n13483) );
  NOR2_X1 U15605 ( .A1(n13500), .A2(n13483), .ZN(n13486) );
  OAI211_X1 U15606 ( .C1(n13486), .C2(n13485), .A(n13484), .B(n10147), .ZN(
        n13489) );
  NAND2_X1 U15607 ( .A1(n13487), .A2(n15531), .ZN(n13488) );
  OAI211_X1 U15608 ( .C1(n13490), .C2(n15508), .A(n13489), .B(n13488), .ZN(
        n13653) );
  INV_X1 U15609 ( .A(n13653), .ZN(n13491) );
  MUX2_X1 U15610 ( .A(n13492), .B(n13491), .S(n15559), .Z(n13498) );
  INV_X1 U15611 ( .A(n13493), .ZN(n13494) );
  OAI22_X1 U15612 ( .A1(n13655), .A2(n13495), .B1(n13494), .B2(n15553), .ZN(
        n13496) );
  INV_X1 U15613 ( .A(n13496), .ZN(n13497) );
  OAI211_X1 U15614 ( .C1(n13656), .C2(n13566), .A(n13498), .B(n13497), .ZN(
        P3_U3214) );
  OAI21_X1 U15615 ( .B1(n7732), .B2(n9481), .A(n13499), .ZN(n13664) );
  INV_X1 U15616 ( .A(n13466), .ZN(n13503) );
  INV_X1 U15617 ( .A(n13500), .ZN(n13501) );
  OAI21_X1 U15618 ( .B1(n13503), .B2(n13502), .A(n13501), .ZN(n13505) );
  AOI222_X1 U15619 ( .A1(n10147), .A2(n13505), .B1(n13504), .B2(n15531), .C1(
        n13525), .C2(n15546), .ZN(n13659) );
  MUX2_X1 U15620 ( .A(n13506), .B(n13659), .S(n15559), .Z(n13509) );
  AOI22_X1 U15621 ( .A1(n13661), .A2(n6428), .B1(n15518), .B2(n13507), .ZN(
        n13508) );
  OAI211_X1 U15622 ( .C1(n13664), .C2(n13566), .A(n13509), .B(n13508), .ZN(
        P3_U3215) );
  OAI21_X1 U15623 ( .B1(n13510), .B2(n13513), .A(n13511), .ZN(n13512) );
  INV_X1 U15624 ( .A(n13512), .ZN(n13670) );
  XNOR2_X1 U15625 ( .A(n13514), .B(n13513), .ZN(n13516) );
  AOI222_X1 U15626 ( .A1(n10147), .A2(n13516), .B1(n13515), .B2(n15543), .C1(
        n13536), .C2(n15546), .ZN(n13665) );
  MUX2_X1 U15627 ( .A(n13517), .B(n13665), .S(n15559), .Z(n13520) );
  AOI22_X1 U15628 ( .A1(n13667), .A2(n6428), .B1(n15518), .B2(n13518), .ZN(
        n13519) );
  OAI211_X1 U15629 ( .C1(n13670), .C2(n13566), .A(n13520), .B(n13519), .ZN(
        P3_U3216) );
  XNOR2_X1 U15630 ( .A(n13522), .B(n13521), .ZN(n13676) );
  XNOR2_X1 U15631 ( .A(n13524), .B(n13523), .ZN(n13526) );
  AOI222_X1 U15632 ( .A1(n10147), .A2(n13526), .B1(n13525), .B2(n15543), .C1(
        n13547), .C2(n15546), .ZN(n13671) );
  MUX2_X1 U15633 ( .A(n13527), .B(n13671), .S(n15559), .Z(n13530) );
  AOI22_X1 U15634 ( .A1(n13673), .A2(n6428), .B1(n15518), .B2(n13528), .ZN(
        n13529) );
  OAI211_X1 U15635 ( .C1(n13676), .C2(n13566), .A(n13530), .B(n13529), .ZN(
        P3_U3217) );
  OAI21_X1 U15636 ( .B1(n13532), .B2(n13534), .A(n13531), .ZN(n13533) );
  INV_X1 U15637 ( .A(n13533), .ZN(n13682) );
  XNOR2_X1 U15638 ( .A(n13535), .B(n13534), .ZN(n13537) );
  AOI222_X1 U15639 ( .A1(n10147), .A2(n13537), .B1(n13536), .B2(n15531), .C1(
        n13559), .C2(n15546), .ZN(n13677) );
  MUX2_X1 U15640 ( .A(n13538), .B(n13677), .S(n15559), .Z(n13541) );
  AOI22_X1 U15641 ( .A1(n13679), .A2(n6428), .B1(n15518), .B2(n13539), .ZN(
        n13540) );
  OAI211_X1 U15642 ( .C1(n13682), .C2(n13566), .A(n13541), .B(n13540), .ZN(
        P3_U3218) );
  AOI21_X1 U15643 ( .B1(n13543), .B2(n13542), .A(n6632), .ZN(n13688) );
  XNOR2_X1 U15644 ( .A(n13544), .B(n13545), .ZN(n13548) );
  AOI222_X1 U15645 ( .A1(n10147), .A2(n13548), .B1(n13547), .B2(n15531), .C1(
        n13546), .C2(n15546), .ZN(n13683) );
  MUX2_X1 U15646 ( .A(n13549), .B(n13683), .S(n15559), .Z(n13552) );
  AOI22_X1 U15647 ( .A1(n13685), .A2(n6428), .B1(n15518), .B2(n13550), .ZN(
        n13551) );
  OAI211_X1 U15648 ( .C1(n13688), .C2(n13566), .A(n13552), .B(n13551), .ZN(
        P3_U3219) );
  XNOR2_X1 U15649 ( .A(n13554), .B(n13555), .ZN(n13696) );
  XNOR2_X1 U15650 ( .A(n13557), .B(n13556), .ZN(n13560) );
  AOI222_X1 U15651 ( .A1(n10147), .A2(n13560), .B1(n13559), .B2(n15531), .C1(
        n13558), .C2(n15546), .ZN(n13689) );
  MUX2_X1 U15652 ( .A(n13561), .B(n13689), .S(n15559), .Z(n13565) );
  AOI22_X1 U15653 ( .A1(n13692), .A2(n6428), .B1(n15518), .B2(n13562), .ZN(
        n13564) );
  OAI211_X1 U15654 ( .C1(n13696), .C2(n13566), .A(n13565), .B(n13564), .ZN(
        P3_U3220) );
  NAND2_X1 U15655 ( .A1(n13361), .A2(n13617), .ZN(n13567) );
  NAND2_X1 U15656 ( .A1(n15612), .A2(n13621), .ZN(n13569) );
  OAI211_X1 U15657 ( .C1(n15612), .C2(n13568), .A(n13567), .B(n13569), .ZN(
        P3_U3490) );
  NAND2_X1 U15658 ( .A1(n15609), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13570) );
  OAI211_X1 U15659 ( .C1(n13571), .C2(n13598), .A(n13570), .B(n13569), .ZN(
        P3_U3489) );
  INV_X1 U15660 ( .A(n13572), .ZN(n13634) );
  INV_X1 U15661 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13576) );
  NAND2_X1 U15662 ( .A1(n13573), .A2(n15596), .ZN(n13574) );
  AOI22_X1 U15663 ( .A1(n13578), .A2(n15596), .B1(n13595), .B2(n13577), .ZN(
        n13579) );
  NAND2_X1 U15664 ( .A1(n13580), .A2(n13579), .ZN(n13635) );
  MUX2_X1 U15665 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13635), .S(n15612), .Z(
        P3_U3483) );
  INV_X1 U15666 ( .A(n13581), .ZN(n13586) );
  INV_X1 U15667 ( .A(n15596), .ZN(n13585) );
  NAND2_X1 U15668 ( .A1(n13582), .A2(n13595), .ZN(n13583) );
  OAI211_X1 U15669 ( .C1(n13586), .C2(n13585), .A(n13584), .B(n13583), .ZN(
        n13636) );
  MUX2_X1 U15670 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13636), .S(n15612), .Z(
        P3_U3482) );
  INV_X1 U15671 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13587) );
  MUX2_X1 U15672 ( .A(n13587), .B(n13637), .S(n15612), .Z(n13589) );
  NAND2_X1 U15673 ( .A1(n13639), .A2(n13617), .ZN(n13588) );
  OAI211_X1 U15674 ( .C1(n13642), .C2(n13620), .A(n13589), .B(n13588), .ZN(
        P3_U3481) );
  MUX2_X1 U15675 ( .A(n13590), .B(n13643), .S(n15612), .Z(n13592) );
  NAND2_X1 U15676 ( .A1(n13645), .A2(n13617), .ZN(n13591) );
  OAI211_X1 U15677 ( .C1(n13648), .C2(n13620), .A(n13592), .B(n13591), .ZN(
        P3_U3480) );
  INV_X1 U15678 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13596) );
  AOI21_X1 U15679 ( .B1(n13595), .B2(n13594), .A(n13593), .ZN(n13649) );
  MUX2_X1 U15680 ( .A(n13596), .B(n13649), .S(n15612), .Z(n13597) );
  OAI21_X1 U15681 ( .B1(n13620), .B2(n13652), .A(n13597), .ZN(P3_U3479) );
  MUX2_X1 U15682 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n13653), .S(n15612), .Z(
        n13600) );
  OAI22_X1 U15683 ( .A1(n13656), .A2(n13620), .B1(n13655), .B2(n13598), .ZN(
        n13599) );
  OR2_X1 U15684 ( .A1(n13600), .A2(n13599), .ZN(P3_U3478) );
  INV_X1 U15685 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13601) );
  MUX2_X1 U15686 ( .A(n13601), .B(n13659), .S(n15612), .Z(n13603) );
  NAND2_X1 U15687 ( .A1(n13661), .A2(n13617), .ZN(n13602) );
  OAI211_X1 U15688 ( .C1(n13620), .C2(n13664), .A(n13603), .B(n13602), .ZN(
        P3_U3477) );
  MUX2_X1 U15689 ( .A(n13604), .B(n13665), .S(n15612), .Z(n13606) );
  NAND2_X1 U15690 ( .A1(n13667), .A2(n13617), .ZN(n13605) );
  OAI211_X1 U15691 ( .C1(n13670), .C2(n13620), .A(n13606), .B(n13605), .ZN(
        P3_U3476) );
  MUX2_X1 U15692 ( .A(n13607), .B(n13671), .S(n15612), .Z(n13609) );
  NAND2_X1 U15693 ( .A1(n13673), .A2(n13617), .ZN(n13608) );
  OAI211_X1 U15694 ( .C1(n13620), .C2(n13676), .A(n13609), .B(n13608), .ZN(
        P3_U3475) );
  INV_X1 U15695 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13610) );
  MUX2_X1 U15696 ( .A(n13610), .B(n13677), .S(n15612), .Z(n13612) );
  NAND2_X1 U15697 ( .A1(n13679), .A2(n13617), .ZN(n13611) );
  OAI211_X1 U15698 ( .C1(n13682), .C2(n13620), .A(n13612), .B(n13611), .ZN(
        P3_U3474) );
  MUX2_X1 U15699 ( .A(n13613), .B(n13683), .S(n15612), .Z(n13615) );
  NAND2_X1 U15700 ( .A1(n13685), .A2(n13617), .ZN(n13614) );
  OAI211_X1 U15701 ( .C1(n13688), .C2(n13620), .A(n13615), .B(n13614), .ZN(
        P3_U3473) );
  MUX2_X1 U15702 ( .A(n13616), .B(n13689), .S(n15612), .Z(n13619) );
  NAND2_X1 U15703 ( .A1(n13692), .A2(n13617), .ZN(n13618) );
  OAI211_X1 U15704 ( .C1(n13620), .C2(n13696), .A(n13619), .B(n13618), .ZN(
        P3_U3472) );
  NAND2_X1 U15705 ( .A1(n13361), .A2(n13691), .ZN(n13622) );
  NAND2_X1 U15706 ( .A1(n15600), .A2(n13621), .ZN(n13625) );
  OAI211_X1 U15707 ( .C1(n15600), .C2(n13623), .A(n13622), .B(n13625), .ZN(
        P3_U3458) );
  INV_X1 U15708 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13627) );
  NAND2_X1 U15709 ( .A1(n13624), .A2(n13691), .ZN(n13626) );
  OAI211_X1 U15710 ( .C1(n13627), .C2(n15600), .A(n13626), .B(n13625), .ZN(
        P3_U3457) );
  MUX2_X1 U15711 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13635), .S(n15600), .Z(
        P3_U3451) );
  MUX2_X1 U15712 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13636), .S(n15600), .Z(
        P3_U3450) );
  INV_X1 U15713 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13638) );
  MUX2_X1 U15714 ( .A(n13638), .B(n13637), .S(n15600), .Z(n13641) );
  NAND2_X1 U15715 ( .A1(n13639), .A2(n13691), .ZN(n13640) );
  OAI211_X1 U15716 ( .C1(n13642), .C2(n13695), .A(n13641), .B(n13640), .ZN(
        P3_U3449) );
  INV_X1 U15717 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13644) );
  MUX2_X1 U15718 ( .A(n13644), .B(n13643), .S(n15600), .Z(n13647) );
  NAND2_X1 U15719 ( .A1(n13645), .A2(n13691), .ZN(n13646) );
  OAI211_X1 U15720 ( .C1(n13648), .C2(n13695), .A(n13647), .B(n13646), .ZN(
        P3_U3448) );
  INV_X1 U15721 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13650) );
  MUX2_X1 U15722 ( .A(n13650), .B(n13649), .S(n15600), .Z(n13651) );
  OAI21_X1 U15723 ( .B1(n13652), .B2(n13695), .A(n13651), .ZN(P3_U3447) );
  MUX2_X1 U15724 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n13653), .S(n15600), .Z(
        n13658) );
  OAI22_X1 U15725 ( .A1(n13656), .A2(n13695), .B1(n13655), .B2(n13654), .ZN(
        n13657) );
  OR2_X1 U15726 ( .A1(n13658), .A2(n13657), .ZN(P3_U3446) );
  INV_X1 U15727 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13660) );
  MUX2_X1 U15728 ( .A(n13660), .B(n13659), .S(n15600), .Z(n13663) );
  NAND2_X1 U15729 ( .A1(n13661), .A2(n13691), .ZN(n13662) );
  OAI211_X1 U15730 ( .C1(n13664), .C2(n13695), .A(n13663), .B(n13662), .ZN(
        P3_U3444) );
  INV_X1 U15731 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13666) );
  MUX2_X1 U15732 ( .A(n13666), .B(n13665), .S(n15600), .Z(n13669) );
  NAND2_X1 U15733 ( .A1(n13667), .A2(n13691), .ZN(n13668) );
  OAI211_X1 U15734 ( .C1(n13670), .C2(n13695), .A(n13669), .B(n13668), .ZN(
        P3_U3441) );
  INV_X1 U15735 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13672) );
  MUX2_X1 U15736 ( .A(n13672), .B(n13671), .S(n15600), .Z(n13675) );
  NAND2_X1 U15737 ( .A1(n13673), .A2(n13691), .ZN(n13674) );
  OAI211_X1 U15738 ( .C1(n13676), .C2(n13695), .A(n13675), .B(n13674), .ZN(
        P3_U3438) );
  INV_X1 U15739 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13678) );
  MUX2_X1 U15740 ( .A(n13678), .B(n13677), .S(n15600), .Z(n13681) );
  NAND2_X1 U15741 ( .A1(n13679), .A2(n13691), .ZN(n13680) );
  OAI211_X1 U15742 ( .C1(n13682), .C2(n13695), .A(n13681), .B(n13680), .ZN(
        P3_U3435) );
  INV_X1 U15743 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13684) );
  MUX2_X1 U15744 ( .A(n13684), .B(n13683), .S(n15600), .Z(n13687) );
  NAND2_X1 U15745 ( .A1(n13685), .A2(n13691), .ZN(n13686) );
  OAI211_X1 U15746 ( .C1(n13688), .C2(n13695), .A(n13687), .B(n13686), .ZN(
        P3_U3432) );
  MUX2_X1 U15747 ( .A(n13690), .B(n13689), .S(n15600), .Z(n13694) );
  NAND2_X1 U15748 ( .A1(n13692), .A2(n13691), .ZN(n13693) );
  OAI211_X1 U15749 ( .C1(n13696), .C2(n13695), .A(n13694), .B(n13693), .ZN(
        P3_U3429) );
  INV_X1 U15750 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13698) );
  NAND3_X1 U15751 ( .A1(n13698), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13700) );
  OAI22_X1 U15752 ( .A1(n13697), .A2(n13700), .B1(n13699), .B2(n13719), .ZN(
        n13701) );
  AOI21_X1 U15753 ( .B1(n13703), .B2(n13702), .A(n13701), .ZN(n13704) );
  INV_X1 U15754 ( .A(n13704), .ZN(P3_U3264) );
  INV_X1 U15755 ( .A(n13705), .ZN(n13706) );
  OAI222_X1 U15756 ( .A1(n13719), .A2(n13707), .B1(n13717), .B2(n13706), .C1(
        P3_U3151), .C2(n8932), .ZN(P3_U3266) );
  INV_X1 U15757 ( .A(n13708), .ZN(n13709) );
  OAI222_X1 U15758 ( .A1(P3_U3151), .A2(n9423), .B1(n13719), .B2(n13710), .C1(
        n13717), .C2(n13709), .ZN(P3_U3267) );
  INV_X1 U15759 ( .A(n13711), .ZN(n13713) );
  OAI222_X1 U15760 ( .A1(n13714), .A2(P3_U3151), .B1(n13717), .B2(n13713), 
        .C1(n13712), .C2(n13719), .ZN(P3_U3268) );
  INV_X1 U15761 ( .A(n13715), .ZN(n13716) );
  OAI222_X1 U15762 ( .A1(n13720), .A2(P3_U3151), .B1(n13719), .B2(n13718), 
        .C1(n13717), .C2(n13716), .ZN(P3_U3269) );
  AOI22_X1 U15763 ( .A1(n13842), .A2(n13802), .B1(n13801), .B2(n13844), .ZN(
        n14139) );
  INV_X1 U15764 ( .A(n13721), .ZN(n13976) );
  AOI22_X1 U15765 ( .A1(n13976), .A2(n13804), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13722) );
  OAI21_X1 U15766 ( .B1(n14139), .B2(n15325), .A(n13722), .ZN(n13729) );
  NAND2_X1 U15767 ( .A1(n13792), .A2(n13723), .ZN(n13796) );
  INV_X1 U15768 ( .A(n13724), .ZN(n13725) );
  OR2_X1 U15769 ( .A1(n13726), .A2(n13725), .ZN(n13753) );
  NAND2_X1 U15770 ( .A1(n13796), .A2(n13753), .ZN(n13728) );
  NAND3_X1 U15771 ( .A1(n13730), .A2(n13821), .A3(n13843), .ZN(n13731) );
  XNOR2_X1 U15772 ( .A(n13733), .B(n13732), .ZN(n13738) );
  OAI22_X1 U15773 ( .A1(n13791), .A2(n13814), .B1(n13734), .B2(n13812), .ZN(
        n14006) );
  AOI22_X1 U15774 ( .A1(n14006), .A2(n13826), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13735) );
  OAI21_X1 U15775 ( .B1(n14011), .B2(n15334), .A(n13735), .ZN(n13736) );
  AOI21_X1 U15776 ( .B1(n14151), .B2(n15332), .A(n13736), .ZN(n13737) );
  OAI21_X1 U15777 ( .B1(n13738), .B2(n15327), .A(n13737), .ZN(P2_U3195) );
  XNOR2_X1 U15778 ( .A(n13740), .B(n13739), .ZN(n13744) );
  AOI22_X1 U15779 ( .A1(n13840), .A2(n13802), .B1(n13801), .B2(n13842), .ZN(
        n14124) );
  AOI22_X1 U15780 ( .A1(n13955), .A2(n13804), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13741) );
  OAI21_X1 U15781 ( .B1(n14124), .B2(n15325), .A(n13741), .ZN(n13742) );
  AOI21_X1 U15782 ( .B1(n13958), .B2(n15332), .A(n13742), .ZN(n13743) );
  OAI21_X1 U15783 ( .B1(n13744), .B2(n15327), .A(n13743), .ZN(P2_U3197) );
  AOI21_X1 U15784 ( .B1(n13747), .B2(n13746), .A(n13745), .ZN(n13752) );
  AND2_X1 U15785 ( .A1(n13851), .A2(n13801), .ZN(n13748) );
  AOI21_X1 U15786 ( .B1(n13849), .B2(n13802), .A(n13748), .ZN(n14077) );
  NAND2_X1 U15787 ( .A1(n13804), .A2(n14084), .ZN(n13749) );
  NAND2_X1 U15788 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13879)
         );
  OAI211_X1 U15789 ( .C1(n14077), .C2(n15325), .A(n13749), .B(n13879), .ZN(
        n13750) );
  AOI21_X1 U15790 ( .B1(n14086), .B2(n15332), .A(n13750), .ZN(n13751) );
  OAI21_X1 U15791 ( .B1(n13752), .B2(n15327), .A(n13751), .ZN(P2_U3198) );
  OAI211_X1 U15792 ( .C1(n13755), .C2(n13754), .A(n13796), .B(n13753), .ZN(
        n13757) );
  NAND2_X1 U15793 ( .A1(n13757), .A2(n13756), .ZN(n13761) );
  XNOR2_X1 U15794 ( .A(n13759), .B(n13758), .ZN(n13760) );
  XNOR2_X1 U15795 ( .A(n13761), .B(n13760), .ZN(n13765) );
  AOI22_X1 U15796 ( .A1(n13841), .A2(n13802), .B1(n13801), .B2(n13843), .ZN(
        n14131) );
  AOI22_X1 U15797 ( .A1(n13967), .A2(n13804), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13762) );
  OAI21_X1 U15798 ( .B1(n14131), .B2(n15325), .A(n13762), .ZN(n13763) );
  AOI21_X1 U15799 ( .B1(n13970), .B2(n15332), .A(n13763), .ZN(n13764) );
  OAI21_X1 U15800 ( .B1(n13765), .B2(n15327), .A(n13764), .ZN(P2_U3201) );
  INV_X1 U15801 ( .A(n13766), .ZN(n13768) );
  NAND2_X1 U15802 ( .A1(n13768), .A2(n13767), .ZN(n13769) );
  XNOR2_X1 U15803 ( .A(n13770), .B(n13769), .ZN(n13776) );
  INV_X1 U15804 ( .A(n14025), .ZN(n13773) );
  OAI22_X1 U15805 ( .A1(n13787), .A2(n13814), .B1(n13771), .B2(n13812), .ZN(
        n14158) );
  AOI22_X1 U15806 ( .A1(n14158), .A2(n13826), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13772) );
  OAI21_X1 U15807 ( .B1(n13773), .B2(n15334), .A(n13772), .ZN(n13774) );
  AOI21_X1 U15808 ( .B1(n14159), .B2(n15332), .A(n13774), .ZN(n13775) );
  OAI21_X1 U15809 ( .B1(n13776), .B2(n15327), .A(n13775), .ZN(P2_U3205) );
  NOR2_X1 U15810 ( .A1(n13777), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15396) );
  AOI21_X1 U15811 ( .B1(n13826), .B2(n13778), .A(n15396), .ZN(n13779) );
  OAI21_X1 U15812 ( .B1(n13780), .B2(n15334), .A(n13779), .ZN(n13785) );
  AOI211_X1 U15813 ( .C1(n13783), .C2(n13782), .A(n15327), .B(n13781), .ZN(
        n13784) );
  AOI211_X1 U15814 ( .C1(n14206), .C2(n15332), .A(n13785), .B(n13784), .ZN(
        n13786) );
  INV_X1 U15815 ( .A(n13786), .ZN(P2_U3206) );
  NOR2_X1 U15816 ( .A1(n13787), .A2(n13812), .ZN(n13788) );
  AOI21_X1 U15817 ( .B1(n13843), .B2(n13802), .A(n13788), .ZN(n13990) );
  AOI22_X1 U15818 ( .A1(n13994), .A2(n13804), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13789) );
  OAI21_X1 U15819 ( .B1(n13990), .B2(n15325), .A(n13789), .ZN(n13794) );
  NOR3_X1 U15820 ( .A1(n13792), .A2(n13791), .A3(n13790), .ZN(n13793) );
  AOI211_X1 U15821 ( .C1(n14147), .C2(n15332), .A(n13794), .B(n13793), .ZN(
        n13795) );
  OAI21_X1 U15822 ( .B1(n15327), .B2(n13796), .A(n13795), .ZN(P2_U3207) );
  AOI21_X1 U15823 ( .B1(n13798), .B2(n13797), .A(n15327), .ZN(n13800) );
  NAND2_X1 U15824 ( .A1(n13800), .A2(n13799), .ZN(n13807) );
  INV_X1 U15825 ( .A(n14049), .ZN(n13805) );
  AOI22_X1 U15826 ( .A1(n13847), .A2(n13802), .B1(n13801), .B2(n13849), .ZN(
        n14172) );
  NAND2_X1 U15827 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n15425)
         );
  OAI21_X1 U15828 ( .B1(n14172), .B2(n15325), .A(n15425), .ZN(n13803) );
  AOI21_X1 U15829 ( .B1(n13805), .B2(n13804), .A(n13803), .ZN(n13806) );
  OAI211_X1 U15830 ( .C1(n14173), .C2(n13820), .A(n13807), .B(n13806), .ZN(
        P2_U3210) );
  OAI21_X1 U15831 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(n13811) );
  NAND2_X1 U15832 ( .A1(n13811), .A2(n13822), .ZN(n13819) );
  OAI22_X1 U15833 ( .A1(n13815), .A2(n13814), .B1(n13813), .B2(n13812), .ZN(
        n14118) );
  OAI22_X1 U15834 ( .A1(n13941), .A2(n15334), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13816), .ZN(n13817) );
  AOI21_X1 U15835 ( .B1(n14118), .B2(n13826), .A(n13817), .ZN(n13818) );
  OAI211_X1 U15836 ( .C1(n13945), .C2(n13820), .A(n13819), .B(n13818), .ZN(
        P2_U3212) );
  AOI22_X1 U15837 ( .A1(n13823), .A2(n13822), .B1(n13821), .B2(n13851), .ZN(
        n13834) );
  INV_X1 U15838 ( .A(n13824), .ZN(n13833) );
  NAND2_X1 U15839 ( .A1(n13826), .A2(n13825), .ZN(n13827) );
  OAI211_X1 U15840 ( .C1(n15334), .C2(n13829), .A(n13828), .B(n13827), .ZN(
        n13830) );
  AOI21_X1 U15841 ( .B1(n13831), .B2(n15332), .A(n13830), .ZN(n13832) );
  OAI21_X1 U15842 ( .B1(n13834), .B2(n13833), .A(n13832), .ZN(P2_U3213) );
  INV_X2 U15843 ( .A(P2_U3947), .ZN(n13858) );
  MUX2_X1 U15844 ( .A(n13835), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13858), .Z(
        P2_U3562) );
  MUX2_X1 U15845 ( .A(n13836), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13858), .Z(
        P2_U3561) );
  MUX2_X1 U15846 ( .A(n13837), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13858), .Z(
        P2_U3560) );
  MUX2_X1 U15847 ( .A(n13838), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13858), .Z(
        P2_U3559) );
  MUX2_X1 U15848 ( .A(n13839), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13858), .Z(
        P2_U3558) );
  MUX2_X1 U15849 ( .A(n13840), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13858), .Z(
        P2_U3557) );
  MUX2_X1 U15850 ( .A(n13841), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13858), .Z(
        P2_U3556) );
  MUX2_X1 U15851 ( .A(n13842), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13858), .Z(
        P2_U3555) );
  MUX2_X1 U15852 ( .A(n13843), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13858), .Z(
        P2_U3554) );
  MUX2_X1 U15853 ( .A(n13844), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13858), .Z(
        P2_U3553) );
  MUX2_X1 U15854 ( .A(n13845), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13858), .Z(
        P2_U3552) );
  MUX2_X1 U15855 ( .A(n13846), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13858), .Z(
        P2_U3551) );
  MUX2_X1 U15856 ( .A(n13847), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13858), .Z(
        P2_U3550) );
  MUX2_X1 U15857 ( .A(n13848), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13858), .Z(
        P2_U3549) );
  MUX2_X1 U15858 ( .A(n13849), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13858), .Z(
        P2_U3548) );
  MUX2_X1 U15859 ( .A(n13850), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13858), .Z(
        P2_U3547) );
  MUX2_X1 U15860 ( .A(n13851), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13858), .Z(
        P2_U3546) );
  MUX2_X1 U15861 ( .A(n13852), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13858), .Z(
        P2_U3545) );
  MUX2_X1 U15862 ( .A(n13853), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13858), .Z(
        P2_U3544) );
  MUX2_X1 U15863 ( .A(n13854), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13858), .Z(
        P2_U3543) );
  MUX2_X1 U15864 ( .A(n13855), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13858), .Z(
        P2_U3542) );
  MUX2_X1 U15865 ( .A(n13856), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13858), .Z(
        P2_U3541) );
  MUX2_X1 U15866 ( .A(n13857), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13858), .Z(
        P2_U3540) );
  MUX2_X1 U15867 ( .A(n13859), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13858), .Z(
        P2_U3539) );
  MUX2_X1 U15868 ( .A(n13860), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13858), .Z(
        P2_U3538) );
  MUX2_X1 U15869 ( .A(n13861), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13858), .Z(
        P2_U3537) );
  MUX2_X1 U15870 ( .A(n13862), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13858), .Z(
        P2_U3536) );
  MUX2_X1 U15871 ( .A(n13863), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13858), .Z(
        P2_U3535) );
  MUX2_X1 U15872 ( .A(n13864), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13858), .Z(
        P2_U3534) );
  MUX2_X1 U15873 ( .A(n13865), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13858), .Z(
        P2_U3533) );
  MUX2_X1 U15874 ( .A(n13866), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13858), .Z(
        P2_U3532) );
  MUX2_X1 U15875 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n13867), .S(n13891), .Z(
        n13873) );
  NAND2_X1 U15876 ( .A1(n13868), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n13871) );
  NAND2_X1 U15877 ( .A1(n13869), .A2(n13875), .ZN(n13870) );
  NAND2_X1 U15878 ( .A1(n13871), .A2(n13870), .ZN(n13872) );
  NAND2_X1 U15879 ( .A1(n13872), .A2(n13873), .ZN(n13896) );
  OAI211_X1 U15880 ( .C1(n13873), .C2(n13872), .A(n13896), .B(n15423), .ZN(
        n13882) );
  AOI22_X1 U15881 ( .A1(n13876), .A2(n13875), .B1(P2_REG1_REG_15__SCAN_IN), 
        .B2(n13874), .ZN(n13886) );
  XNOR2_X1 U15882 ( .A(n13891), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13885) );
  XOR2_X1 U15883 ( .A(n13886), .B(n13885), .Z(n13877) );
  NAND2_X1 U15884 ( .A1(n15419), .A2(n13877), .ZN(n13878) );
  NAND2_X1 U15885 ( .A1(n13879), .A2(n13878), .ZN(n13880) );
  AOI21_X1 U15886 ( .B1(n15373), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n13880), 
        .ZN(n13881) );
  OAI211_X1 U15887 ( .C1(n15408), .C2(n13883), .A(n13882), .B(n13881), .ZN(
        P2_U3230) );
  INV_X1 U15888 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13884) );
  OAI22_X1 U15889 ( .A1(n13886), .A2(n13885), .B1(n13884), .B2(n13883), .ZN(
        n13902) );
  INV_X1 U15890 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13887) );
  XNOR2_X1 U15891 ( .A(n13906), .B(n13887), .ZN(n13901) );
  XNOR2_X1 U15892 ( .A(n13902), .B(n13901), .ZN(n13900) );
  INV_X1 U15893 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n13889) );
  OAI21_X1 U15894 ( .B1(n15427), .B2(n13889), .A(n13888), .ZN(n13890) );
  AOI21_X1 U15895 ( .B1(n13906), .B2(n15421), .A(n13890), .ZN(n13899) );
  NAND2_X1 U15896 ( .A1(n13891), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13895) );
  NAND2_X1 U15897 ( .A1(n13896), .A2(n13895), .ZN(n13893) );
  MUX2_X1 U15898 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n14063), .S(n13906), .Z(
        n13892) );
  NAND2_X1 U15899 ( .A1(n13893), .A2(n13892), .ZN(n13908) );
  MUX2_X1 U15900 ( .A(n14063), .B(P2_REG2_REG_17__SCAN_IN), .S(n13906), .Z(
        n13894) );
  NAND3_X1 U15901 ( .A1(n13896), .A2(n13895), .A3(n13894), .ZN(n13897) );
  NAND3_X1 U15902 ( .A1(n13908), .A2(n15423), .A3(n13897), .ZN(n13898) );
  OAI211_X1 U15903 ( .C1(n13900), .C2(n15392), .A(n13899), .B(n13898), .ZN(
        P2_U3231) );
  AOI22_X1 U15904 ( .A1(n13902), .A2(n13901), .B1(P2_REG1_REG_17__SCAN_IN), 
        .B2(n13906), .ZN(n13903) );
  XNOR2_X1 U15905 ( .A(n13903), .B(n15422), .ZN(n15418) );
  INV_X1 U15906 ( .A(n13903), .ZN(n13904) );
  AOI22_X1 U15907 ( .A1(n15418), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n15422), 
        .B2(n13904), .ZN(n13905) );
  XNOR2_X1 U15908 ( .A(n13905), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13914) );
  NAND2_X1 U15909 ( .A1(n13906), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13907) );
  NAND2_X1 U15910 ( .A1(n13908), .A2(n13907), .ZN(n13909) );
  NAND2_X1 U15911 ( .A1(n13909), .A2(n15422), .ZN(n13910) );
  NAND2_X1 U15912 ( .A1(n13911), .A2(n13910), .ZN(n15415) );
  NAND2_X1 U15913 ( .A1(n15417), .A2(n13911), .ZN(n13912) );
  XNOR2_X1 U15914 ( .A(n13912), .B(n14035), .ZN(n13915) );
  INV_X1 U15915 ( .A(n13915), .ZN(n13913) );
  AOI22_X1 U15916 ( .A1(n13914), .A2(n15419), .B1(n13913), .B2(n15423), .ZN(
        n13917) );
  XNOR2_X1 U15917 ( .A(n13919), .B(n14093), .ZN(n13920) );
  NAND2_X1 U15918 ( .A1(n13920), .A2(n15443), .ZN(n14094) );
  NOR2_X1 U15919 ( .A1(n14064), .A2(n13921), .ZN(n13923) );
  AOI211_X1 U15920 ( .C1(n14093), .C2(n14085), .A(n13923), .B(n13922), .ZN(
        n13924) );
  OAI21_X1 U15921 ( .B1(n14094), .B2(n14089), .A(n13924), .ZN(P2_U3234) );
  XNOR2_X1 U15922 ( .A(n13926), .B(n13925), .ZN(n14116) );
  AOI21_X1 U15923 ( .B1(n13929), .B2(n13928), .A(n13927), .ZN(n13931) );
  INV_X1 U15924 ( .A(n13932), .ZN(n13933) );
  AOI211_X1 U15925 ( .C1(n14115), .C2(n13940), .A(n14166), .B(n13933), .ZN(
        n14114) );
  NAND2_X1 U15926 ( .A1(n14114), .A2(n15445), .ZN(n13936) );
  AOI22_X1 U15927 ( .A1(n13934), .A2(n14083), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n6438), .ZN(n13935) );
  OAI211_X1 U15928 ( .C1(n13937), .C2(n15437), .A(n13936), .B(n13935), .ZN(
        n13938) );
  AOI21_X1 U15929 ( .B1(n14113), .B2(n14064), .A(n13938), .ZN(n13939) );
  OAI21_X1 U15930 ( .B1(n14116), .B2(n14056), .A(n13939), .ZN(P2_U3238) );
  AOI211_X1 U15931 ( .C1(n14119), .C2(n6517), .A(n14166), .B(n7413), .ZN(
        n14117) );
  INV_X1 U15932 ( .A(n13941), .ZN(n13942) );
  AOI22_X1 U15933 ( .A1(n13942), .A2(n14083), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n6438), .ZN(n13944) );
  NAND2_X1 U15934 ( .A1(n14118), .A2(n14064), .ZN(n13943) );
  OAI211_X1 U15935 ( .C1(n13945), .C2(n15437), .A(n13944), .B(n13943), .ZN(
        n13946) );
  AOI21_X1 U15936 ( .B1(n14117), .B2(n15445), .A(n13946), .ZN(n13950) );
  XOR2_X1 U15937 ( .A(n13948), .B(n13947), .Z(n14120) );
  NAND2_X1 U15938 ( .A1(n14120), .A2(n14054), .ZN(n13949) );
  OAI211_X1 U15939 ( .C1(n14123), .C2(n14056), .A(n13950), .B(n13949), .ZN(
        P2_U3239) );
  XNOR2_X1 U15940 ( .A(n13952), .B(n13951), .ZN(n14130) );
  XNOR2_X1 U15941 ( .A(n13954), .B(n13953), .ZN(n14128) );
  OAI211_X1 U15942 ( .C1(n13965), .C2(n14126), .A(n15443), .B(n6517), .ZN(
        n14125) );
  AOI22_X1 U15943 ( .A1(n13955), .A2(n14083), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n6438), .ZN(n13956) );
  OAI21_X1 U15944 ( .B1(n14124), .B2(n6438), .A(n13956), .ZN(n13957) );
  AOI21_X1 U15945 ( .B1(n13958), .B2(n14085), .A(n13957), .ZN(n13959) );
  OAI21_X1 U15946 ( .B1(n14125), .B2(n14089), .A(n13959), .ZN(n13960) );
  AOI21_X1 U15947 ( .B1(n14128), .B2(n14054), .A(n13960), .ZN(n13961) );
  OAI21_X1 U15948 ( .B1(n14130), .B2(n14056), .A(n13961), .ZN(P2_U3240) );
  XNOR2_X1 U15949 ( .A(n13962), .B(n13963), .ZN(n14137) );
  XNOR2_X1 U15950 ( .A(n13964), .B(n13963), .ZN(n14135) );
  INV_X1 U15951 ( .A(n13965), .ZN(n13966) );
  OAI211_X1 U15952 ( .C1(n14133), .C2(n13975), .A(n13966), .B(n15443), .ZN(
        n14132) );
  AOI22_X1 U15953 ( .A1(n13967), .A2(n14083), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n6438), .ZN(n13968) );
  OAI21_X1 U15954 ( .B1(n14131), .B2(n6438), .A(n13968), .ZN(n13969) );
  AOI21_X1 U15955 ( .B1(n13970), .B2(n14085), .A(n13969), .ZN(n13971) );
  OAI21_X1 U15956 ( .B1(n14132), .B2(n14089), .A(n13971), .ZN(n13972) );
  AOI21_X1 U15957 ( .B1(n14135), .B2(n14054), .A(n13972), .ZN(n13973) );
  OAI21_X1 U15958 ( .B1(n14137), .B2(n14056), .A(n13973), .ZN(P2_U3241) );
  XOR2_X1 U15959 ( .A(n13974), .B(n13981), .Z(n14144) );
  AOI211_X1 U15960 ( .C1(n14138), .C2(n13992), .A(n14166), .B(n13975), .ZN(
        n14140) );
  NAND2_X1 U15961 ( .A1(n14138), .A2(n14085), .ZN(n13978) );
  AOI22_X1 U15962 ( .A1(n13976), .A2(n14083), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n6438), .ZN(n13977) );
  OAI211_X1 U15963 ( .C1(n6438), .C2(n14139), .A(n13978), .B(n13977), .ZN(
        n13979) );
  AOI21_X1 U15964 ( .B1(n14140), .B2(n15445), .A(n13979), .ZN(n13983) );
  XOR2_X1 U15965 ( .A(n13981), .B(n13980), .Z(n14142) );
  NAND2_X1 U15966 ( .A1(n14142), .A2(n14054), .ZN(n13982) );
  OAI211_X1 U15967 ( .C1(n14144), .C2(n14056), .A(n13983), .B(n13982), .ZN(
        P2_U3242) );
  OAI21_X1 U15968 ( .B1(n13984), .B2(n13986), .A(n13985), .ZN(n14149) );
  OAI211_X1 U15969 ( .C1(n13989), .C2(n13988), .A(n13987), .B(n15479), .ZN(
        n13991) );
  NAND2_X1 U15970 ( .A1(n13991), .A2(n13990), .ZN(n14146) );
  INV_X1 U15971 ( .A(n13992), .ZN(n13993) );
  AOI211_X1 U15972 ( .C1(n14147), .C2(n14009), .A(n14166), .B(n13993), .ZN(
        n14145) );
  NAND2_X1 U15973 ( .A1(n14145), .A2(n15445), .ZN(n13996) );
  AOI22_X1 U15974 ( .A1(n13994), .A2(n14083), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n6438), .ZN(n13995) );
  OAI211_X1 U15975 ( .C1(n13997), .C2(n15437), .A(n13996), .B(n13995), .ZN(
        n13998) );
  AOI21_X1 U15976 ( .B1(n14064), .B2(n14146), .A(n13998), .ZN(n13999) );
  OAI21_X1 U15977 ( .B1(n14149), .B2(n14056), .A(n13999), .ZN(P2_U3243) );
  NAND2_X1 U15978 ( .A1(n14001), .A2(n14000), .ZN(n14040) );
  INV_X1 U15979 ( .A(n14039), .ZN(n14003) );
  OAI21_X1 U15980 ( .B1(n14040), .B2(n14003), .A(n14002), .ZN(n14021) );
  NOR2_X1 U15981 ( .A1(n14021), .A2(n14022), .ZN(n14020) );
  NOR2_X1 U15982 ( .A1(n14020), .A2(n14004), .ZN(n14005) );
  XNOR2_X1 U15983 ( .A(n14005), .B(n14016), .ZN(n14007) );
  AOI21_X1 U15984 ( .B1(n14007), .B2(n15479), .A(n14006), .ZN(n14154) );
  OAI211_X1 U15985 ( .C1(n14024), .C2(n14010), .A(n15443), .B(n14009), .ZN(
        n14152) );
  INV_X1 U15986 ( .A(n14011), .ZN(n14012) );
  AOI22_X1 U15987 ( .A1(n14012), .A2(n14083), .B1(n6438), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n14014) );
  NAND2_X1 U15988 ( .A1(n14151), .A2(n14085), .ZN(n14013) );
  OAI211_X1 U15989 ( .C1(n14152), .C2(n14089), .A(n14014), .B(n14013), .ZN(
        n14015) );
  INV_X1 U15990 ( .A(n14015), .ZN(n14019) );
  OR2_X1 U15991 ( .A1(n6614), .A2(n14016), .ZN(n14150) );
  NAND3_X1 U15992 ( .A1(n14150), .A2(n14017), .A3(n15446), .ZN(n14018) );
  OAI211_X1 U15993 ( .C1(n14154), .C2(n6438), .A(n14019), .B(n14018), .ZN(
        P2_U3244) );
  AOI21_X1 U15994 ( .B1(n14022), .B2(n14021), .A(n14020), .ZN(n14162) );
  XOR2_X1 U15995 ( .A(n14023), .B(n14022), .Z(n14156) );
  NAND2_X1 U15996 ( .A1(n14156), .A2(n15446), .ZN(n14031) );
  AOI211_X1 U15997 ( .C1(n14159), .C2(n6492), .A(n14166), .B(n14024), .ZN(
        n14157) );
  AOI22_X1 U15998 ( .A1(n6438), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14025), 
        .B2(n14083), .ZN(n14027) );
  NAND2_X1 U15999 ( .A1(n14158), .A2(n14064), .ZN(n14026) );
  OAI211_X1 U16000 ( .C1(n14028), .C2(n15437), .A(n14027), .B(n14026), .ZN(
        n14029) );
  AOI21_X1 U16001 ( .B1(n14157), .B2(n15445), .A(n14029), .ZN(n14030) );
  OAI211_X1 U16002 ( .C1(n14162), .C2(n14070), .A(n14031), .B(n14030), .ZN(
        P2_U3245) );
  XNOR2_X1 U16003 ( .A(n14032), .B(n14039), .ZN(n14171) );
  OAI21_X1 U16004 ( .B1(n14033), .B2(n14047), .A(n6492), .ZN(n14167) );
  OAI21_X1 U16005 ( .B1(n14167), .B2(n9716), .A(n14165), .ZN(n14038) );
  NOR2_X1 U16006 ( .A1(n14033), .A2(n15437), .ZN(n14037) );
  OAI22_X1 U16007 ( .A1(n14064), .A2(n14035), .B1(n14034), .B2(n15434), .ZN(
        n14036) );
  AOI211_X1 U16008 ( .C1(n14038), .C2(n14064), .A(n14037), .B(n14036), .ZN(
        n14042) );
  XNOR2_X1 U16009 ( .A(n14040), .B(n14039), .ZN(n14169) );
  NAND2_X1 U16010 ( .A1(n14169), .A2(n14054), .ZN(n14041) );
  OAI211_X1 U16011 ( .C1(n14171), .C2(n14056), .A(n14042), .B(n14041), .ZN(
        P2_U3246) );
  XNOR2_X1 U16012 ( .A(n14044), .B(n14043), .ZN(n14178) );
  XNOR2_X1 U16013 ( .A(n14046), .B(n14045), .ZN(n14176) );
  AOI211_X1 U16014 ( .C1(n14048), .C2(n14058), .A(n14166), .B(n14047), .ZN(
        n14174) );
  NAND2_X1 U16015 ( .A1(n14174), .A2(n15445), .ZN(n14052) );
  OAI22_X1 U16016 ( .A1(n14172), .A2(n6438), .B1(n14049), .B2(n15434), .ZN(
        n14050) );
  AOI21_X1 U16017 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n6438), .A(n14050), .ZN(
        n14051) );
  OAI211_X1 U16018 ( .C1(n14173), .C2(n15437), .A(n14052), .B(n14051), .ZN(
        n14053) );
  AOI21_X1 U16019 ( .B1(n14054), .B2(n14176), .A(n14053), .ZN(n14055) );
  OAI21_X1 U16020 ( .B1(n14178), .B2(n14056), .A(n14055), .ZN(P2_U3247) );
  XOR2_X1 U16021 ( .A(n14057), .B(n14066), .Z(n14185) );
  AOI211_X1 U16022 ( .C1(n14181), .C2(n14081), .A(n14166), .B(n7403), .ZN(
        n14179) );
  NAND2_X1 U16023 ( .A1(n14181), .A2(n14085), .ZN(n14062) );
  INV_X1 U16024 ( .A(n14059), .ZN(n14060) );
  AOI22_X1 U16025 ( .A1(n14064), .A2(n14180), .B1(n14060), .B2(n14083), .ZN(
        n14061) );
  OAI211_X1 U16026 ( .C1(n14064), .C2(n14063), .A(n14062), .B(n14061), .ZN(
        n14065) );
  AOI21_X1 U16027 ( .B1(n14179), .B2(n15445), .A(n14065), .ZN(n14069) );
  XNOR2_X1 U16028 ( .A(n14067), .B(n14066), .ZN(n14182) );
  NAND2_X1 U16029 ( .A1(n14182), .A2(n15446), .ZN(n14068) );
  OAI211_X1 U16030 ( .C1(n14185), .C2(n14070), .A(n14069), .B(n14068), .ZN(
        P2_U3248) );
  OAI21_X1 U16031 ( .B1(n6518), .B2(n14073), .A(n14071), .ZN(n14079) );
  OR2_X1 U16032 ( .A1(n14079), .A2(n14072), .ZN(n14078) );
  XNOR2_X1 U16033 ( .A(n14074), .B(n14073), .ZN(n14075) );
  NAND2_X1 U16034 ( .A1(n14075), .A2(n15479), .ZN(n14076) );
  INV_X1 U16035 ( .A(n14079), .ZN(n14190) );
  AOI21_X1 U16036 ( .B1(n14080), .B2(n14086), .A(n14166), .ZN(n14082) );
  NAND2_X1 U16037 ( .A1(n14082), .A2(n14081), .ZN(n14187) );
  AOI22_X1 U16038 ( .A1(n6438), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n14084), 
        .B2(n14083), .ZN(n14088) );
  NAND2_X1 U16039 ( .A1(n14086), .A2(n14085), .ZN(n14087) );
  OAI211_X1 U16040 ( .C1(n14187), .C2(n14089), .A(n14088), .B(n14087), .ZN(
        n14090) );
  AOI21_X1 U16041 ( .B1(n14190), .B2(n14091), .A(n14090), .ZN(n14092) );
  OAI21_X1 U16042 ( .B1(n14192), .B2(n6438), .A(n14092), .ZN(P2_U3249) );
  INV_X1 U16043 ( .A(n14093), .ZN(n14095) );
  OAI211_X1 U16044 ( .C1(n14095), .C2(n15490), .A(n14094), .B(n14096), .ZN(
        n14224) );
  MUX2_X1 U16045 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14224), .S(n15502), .Z(
        P2_U3530) );
  OAI211_X1 U16046 ( .C1(n14098), .C2(n15490), .A(n14097), .B(n14096), .ZN(
        n14225) );
  MUX2_X1 U16047 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14225), .S(n15502), .Z(
        P2_U3529) );
  NAND3_X1 U16048 ( .A1(n14109), .A2(n12965), .A3(n14104), .ZN(n14107) );
  AOI21_X1 U16049 ( .B1(n12965), .B2(n14102), .A(n15475), .ZN(n14103) );
  INV_X1 U16050 ( .A(n14105), .ZN(n14106) );
  NAND2_X1 U16051 ( .A1(n14107), .A2(n14106), .ZN(n14110) );
  MUX2_X1 U16052 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14226), .S(n15502), .Z(
        P2_U3528) );
  AOI211_X1 U16053 ( .C1(n15472), .C2(n14119), .A(n14118), .B(n14117), .ZN(
        n14122) );
  NAND2_X1 U16054 ( .A1(n14120), .A2(n15479), .ZN(n14121) );
  OAI211_X1 U16055 ( .C1(n14123), .C2(n15475), .A(n14122), .B(n14121), .ZN(
        n14228) );
  MUX2_X1 U16056 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14228), .S(n15502), .Z(
        P2_U3525) );
  OAI211_X1 U16057 ( .C1(n14126), .C2(n15490), .A(n14125), .B(n14124), .ZN(
        n14127) );
  AOI21_X1 U16058 ( .B1(n14128), .B2(n15479), .A(n14127), .ZN(n14129) );
  OAI21_X1 U16059 ( .B1(n14130), .B2(n15475), .A(n14129), .ZN(n14229) );
  MUX2_X1 U16060 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14229), .S(n15502), .Z(
        P2_U3524) );
  OAI211_X1 U16061 ( .C1(n14133), .C2(n15490), .A(n14132), .B(n14131), .ZN(
        n14134) );
  AOI21_X1 U16062 ( .B1(n14135), .B2(n15479), .A(n14134), .ZN(n14136) );
  OAI21_X1 U16063 ( .B1(n14137), .B2(n15475), .A(n14136), .ZN(n14230) );
  MUX2_X1 U16064 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14230), .S(n15502), .Z(
        P2_U3523) );
  OAI21_X1 U16065 ( .B1(n7412), .B2(n15490), .A(n14139), .ZN(n14141) );
  AOI211_X1 U16066 ( .C1(n14142), .C2(n15479), .A(n14141), .B(n14140), .ZN(
        n14143) );
  OAI21_X1 U16067 ( .B1(n14144), .B2(n15475), .A(n14143), .ZN(n14231) );
  MUX2_X1 U16068 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14231), .S(n15502), .Z(
        P2_U3522) );
  AOI211_X1 U16069 ( .C1(n15472), .C2(n14147), .A(n14146), .B(n14145), .ZN(
        n14148) );
  OAI21_X1 U16070 ( .B1(n14149), .B2(n15475), .A(n14148), .ZN(n14232) );
  MUX2_X1 U16071 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14232), .S(n15502), .Z(
        P2_U3521) );
  NAND3_X1 U16072 ( .A1(n14150), .A2(n14017), .A3(n8826), .ZN(n14155) );
  NAND2_X1 U16073 ( .A1(n14151), .A2(n15472), .ZN(n14153) );
  NAND4_X1 U16074 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        n14233) );
  MUX2_X1 U16075 ( .A(n14233), .B(P2_REG1_REG_21__SCAN_IN), .S(n15500), .Z(
        P2_U3520) );
  NAND2_X1 U16076 ( .A1(n14156), .A2(n8826), .ZN(n14161) );
  AOI211_X1 U16077 ( .C1(n15472), .C2(n14159), .A(n14158), .B(n14157), .ZN(
        n14160) );
  OAI211_X1 U16078 ( .C1(n14162), .C2(n14186), .A(n14161), .B(n14160), .ZN(
        n14234) );
  MUX2_X1 U16079 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14234), .S(n15502), .Z(
        P2_U3519) );
  NAND2_X1 U16080 ( .A1(n14163), .A2(n15472), .ZN(n14164) );
  OAI211_X1 U16081 ( .C1(n14167), .C2(n14166), .A(n14165), .B(n14164), .ZN(
        n14168) );
  AOI21_X1 U16082 ( .B1(n14169), .B2(n15479), .A(n14168), .ZN(n14170) );
  OAI21_X1 U16083 ( .B1(n14171), .B2(n15475), .A(n14170), .ZN(n14235) );
  MUX2_X1 U16084 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14235), .S(n15502), .Z(
        P2_U3518) );
  OAI21_X1 U16085 ( .B1(n14173), .B2(n15490), .A(n14172), .ZN(n14175) );
  AOI211_X1 U16086 ( .C1(n14176), .C2(n15479), .A(n14175), .B(n14174), .ZN(
        n14177) );
  OAI21_X1 U16087 ( .B1(n14178), .B2(n15475), .A(n14177), .ZN(n14236) );
  MUX2_X1 U16088 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14236), .S(n15502), .Z(
        P2_U3517) );
  AOI211_X1 U16089 ( .C1(n15472), .C2(n14181), .A(n14180), .B(n14179), .ZN(
        n14184) );
  NAND2_X1 U16090 ( .A1(n14182), .A2(n8826), .ZN(n14183) );
  OAI211_X1 U16091 ( .C1(n14186), .C2(n14185), .A(n14184), .B(n14183), .ZN(
        n14237) );
  MUX2_X1 U16092 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14237), .S(n15502), .Z(
        P2_U3516) );
  OAI21_X1 U16093 ( .B1(n14188), .B2(n15490), .A(n14187), .ZN(n14189) );
  AOI21_X1 U16094 ( .B1(n14190), .B2(n15495), .A(n14189), .ZN(n14191) );
  NAND2_X1 U16095 ( .A1(n14192), .A2(n14191), .ZN(n14238) );
  MUX2_X1 U16096 ( .A(n14238), .B(P2_REG1_REG_16__SCAN_IN), .S(n15500), .Z(
        P2_U3515) );
  OAI211_X1 U16097 ( .C1(n14195), .C2(n15490), .A(n14194), .B(n14193), .ZN(
        n14196) );
  AOI21_X1 U16098 ( .B1(n14197), .B2(n15479), .A(n14196), .ZN(n14198) );
  OAI21_X1 U16099 ( .B1(n14199), .B2(n15475), .A(n14198), .ZN(n14239) );
  MUX2_X1 U16100 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14239), .S(n15502), .Z(
        P2_U3514) );
  AOI21_X1 U16101 ( .B1(n15472), .B2(n14201), .A(n14200), .ZN(n14203) );
  OAI211_X1 U16102 ( .C1(n15475), .C2(n14204), .A(n14203), .B(n14202), .ZN(
        n14240) );
  MUX2_X1 U16103 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14240), .S(n15502), .Z(
        P2_U3513) );
  AOI21_X1 U16104 ( .B1(n15472), .B2(n14206), .A(n14205), .ZN(n14207) );
  OAI211_X1 U16105 ( .C1(n15475), .C2(n14209), .A(n14208), .B(n14207), .ZN(
        n14241) );
  MUX2_X1 U16106 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14241), .S(n15502), .Z(
        P2_U3512) );
  INV_X1 U16107 ( .A(n14210), .ZN(n14215) );
  AOI21_X1 U16108 ( .B1(n15472), .B2(n14212), .A(n14211), .ZN(n14213) );
  OAI211_X1 U16109 ( .C1(n14215), .C2(n14222), .A(n14214), .B(n14213), .ZN(
        n14242) );
  MUX2_X1 U16110 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n14242), .S(n15502), .Z(
        P2_U3510) );
  AOI21_X1 U16111 ( .B1(n15472), .B2(n14217), .A(n14216), .ZN(n14220) );
  INV_X1 U16112 ( .A(n14218), .ZN(n14219) );
  OAI211_X1 U16113 ( .C1(n14222), .C2(n14221), .A(n14220), .B(n14219), .ZN(
        n14243) );
  MUX2_X1 U16114 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14243), .S(n15502), .Z(
        P2_U3507) );
  MUX2_X1 U16115 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n14223), .S(n15502), .Z(
        P2_U3506) );
  MUX2_X1 U16116 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14224), .S(n15496), .Z(
        P2_U3498) );
  MUX2_X1 U16117 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14225), .S(n15496), .Z(
        P2_U3497) );
  MUX2_X1 U16118 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14226), .S(n15496), .Z(
        P2_U3496) );
  MUX2_X1 U16119 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14228), .S(n15496), .Z(
        P2_U3493) );
  MUX2_X1 U16120 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14229), .S(n15496), .Z(
        P2_U3492) );
  MUX2_X1 U16121 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14230), .S(n15496), .Z(
        P2_U3491) );
  MUX2_X1 U16122 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14231), .S(n15496), .Z(
        P2_U3490) );
  MUX2_X1 U16123 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14232), .S(n15496), .Z(
        P2_U3489) );
  MUX2_X1 U16124 ( .A(n14233), .B(P2_REG0_REG_21__SCAN_IN), .S(n6954), .Z(
        P2_U3488) );
  MUX2_X1 U16125 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14234), .S(n15496), .Z(
        P2_U3487) );
  MUX2_X1 U16126 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14235), .S(n15496), .Z(
        P2_U3486) );
  MUX2_X1 U16127 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14236), .S(n15496), .Z(
        P2_U3484) );
  MUX2_X1 U16128 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14237), .S(n15496), .Z(
        P2_U3481) );
  MUX2_X1 U16129 ( .A(n14238), .B(P2_REG0_REG_16__SCAN_IN), .S(n6954), .Z(
        P2_U3478) );
  MUX2_X1 U16130 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14239), .S(n15496), .Z(
        P2_U3475) );
  MUX2_X1 U16131 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14240), .S(n15496), .Z(
        P2_U3472) );
  MUX2_X1 U16132 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14241), .S(n15496), .Z(
        P2_U3469) );
  MUX2_X1 U16133 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n14242), .S(n15496), .Z(
        P2_U3463) );
  MUX2_X1 U16134 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n14243), .S(n15496), .Z(
        P2_U3454) );
  INV_X1 U16135 ( .A(n14244), .ZN(n15156) );
  NAND3_X1 U16136 ( .A1(n14246), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14249) );
  OAI22_X1 U16137 ( .A1(n14245), .A2(n14249), .B1(n14248), .B2(n14247), .ZN(
        n14250) );
  INV_X1 U16138 ( .A(n14250), .ZN(n14251) );
  OAI21_X1 U16139 ( .B1(n15156), .B2(n14257), .A(n14251), .ZN(P2_U3296) );
  INV_X1 U16140 ( .A(n14252), .ZN(n15158) );
  OAI222_X1 U16141 ( .A1(n14247), .A2(n14253), .B1(n14257), .B2(n15158), .C1(
        n8420), .C2(P2_U3088), .ZN(P2_U3298) );
  AOI21_X1 U16142 ( .B1(n14255), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14254), 
        .ZN(n14256) );
  OAI21_X1 U16143 ( .B1(n14258), .B2(n14257), .A(n14256), .ZN(P2_U3299) );
  MUX2_X1 U16144 ( .A(n14259), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OR2_X1 U16145 ( .A1(n15003), .A2(n14413), .ZN(n14261) );
  NAND2_X1 U16146 ( .A1(n15009), .A2(n10794), .ZN(n14260) );
  OAI22_X1 U16147 ( .A1(n15003), .A2(n14414), .B1(n14966), .B2(n14413), .ZN(
        n14262) );
  XNOR2_X1 U16148 ( .A(n14262), .B(n11660), .ZN(n14461) );
  OAI22_X1 U16149 ( .A1(n15019), .A2(n14413), .B1(n14992), .B2(n14411), .ZN(
        n14271) );
  NAND2_X1 U16150 ( .A1(n15112), .A2(n14346), .ZN(n14269) );
  NAND2_X1 U16151 ( .A1(n14573), .A2(n14295), .ZN(n14267) );
  NAND3_X1 U16152 ( .A1(n14269), .A2(n14359), .A3(n14267), .ZN(n14268) );
  OAI21_X1 U16153 ( .B1(n14269), .B2(n14359), .A(n14268), .ZN(n14270) );
  XNOR2_X1 U16154 ( .A(n14271), .B(n14270), .ZN(n14383) );
  INV_X1 U16155 ( .A(n14270), .ZN(n14272) );
  OAI22_X1 U16156 ( .A1(n15105), .A2(n14414), .B1(n14994), .B2(n14413), .ZN(
        n14273) );
  XNOR2_X1 U16157 ( .A(n14273), .B(n14359), .ZN(n14277) );
  OR2_X1 U16158 ( .A1(n15105), .A2(n14413), .ZN(n14275) );
  NAND2_X1 U16159 ( .A1(n6981), .A2(n10794), .ZN(n14274) );
  NAND2_X1 U16160 ( .A1(n14275), .A2(n14274), .ZN(n14276) );
  NOR2_X1 U16161 ( .A1(n14277), .A2(n14276), .ZN(n14475) );
  AOI21_X1 U16162 ( .B1(n14277), .B2(n14276), .A(n14475), .ZN(n14466) );
  OAI21_X1 U16163 ( .B1(n14461), .B2(n14463), .A(n14466), .ZN(n14278) );
  OAI22_X1 U16164 ( .A1(n14955), .A2(n14414), .B1(n14967), .B2(n14413), .ZN(
        n14279) );
  XNOR2_X1 U16165 ( .A(n14279), .B(n11660), .ZN(n14282) );
  OR2_X1 U16166 ( .A1(n14955), .A2(n14413), .ZN(n14281) );
  NAND2_X1 U16167 ( .A1(n14572), .A2(n10794), .ZN(n14280) );
  AND2_X1 U16168 ( .A1(n14281), .A2(n14280), .ZN(n14283) );
  NAND2_X1 U16169 ( .A1(n14282), .A2(n14283), .ZN(n14287) );
  INV_X1 U16170 ( .A(n14282), .ZN(n14285) );
  INV_X1 U16171 ( .A(n14283), .ZN(n14284) );
  NAND2_X1 U16172 ( .A1(n14285), .A2(n14284), .ZN(n14286) );
  AND2_X1 U16173 ( .A1(n14287), .A2(n14286), .ZN(n14474) );
  OAI22_X1 U16174 ( .A1(n15144), .A2(n14413), .B1(n14407), .B2(n14411), .ZN(
        n14290) );
  OAI22_X1 U16175 ( .A1(n15144), .A2(n14414), .B1(n14407), .B2(n14413), .ZN(
        n14288) );
  XNOR2_X1 U16176 ( .A(n14288), .B(n14359), .ZN(n14289) );
  XOR2_X1 U16177 ( .A(n14290), .B(n14289), .Z(n14529) );
  INV_X1 U16178 ( .A(n14289), .ZN(n14292) );
  NOR2_X1 U16179 ( .A1(n14932), .A2(n14411), .ZN(n14294) );
  AOI21_X1 U16180 ( .B1(n15088), .B2(n14351), .A(n14294), .ZN(n14300) );
  NAND2_X1 U16181 ( .A1(n15088), .A2(n14346), .ZN(n14297) );
  NAND2_X1 U16182 ( .A1(n14900), .A2(n14295), .ZN(n14296) );
  NAND2_X1 U16183 ( .A1(n14297), .A2(n14296), .ZN(n14298) );
  XNOR2_X1 U16184 ( .A(n14298), .B(n14359), .ZN(n14299) );
  XOR2_X1 U16185 ( .A(n14300), .B(n14299), .Z(n14403) );
  INV_X1 U16186 ( .A(n14300), .ZN(n14301) );
  NAND2_X1 U16187 ( .A1(n14299), .A2(n14301), .ZN(n14302) );
  NAND2_X1 U16188 ( .A1(n14910), .A2(n14346), .ZN(n14304) );
  NAND2_X1 U16189 ( .A1(n14878), .A2(n14351), .ZN(n14303) );
  NAND2_X1 U16190 ( .A1(n14304), .A2(n14303), .ZN(n14305) );
  XNOR2_X1 U16191 ( .A(n14305), .B(n14359), .ZN(n14309) );
  AND2_X1 U16192 ( .A1(n14878), .A2(n10794), .ZN(n14306) );
  AOI21_X1 U16193 ( .B1(n14910), .B2(n14351), .A(n14306), .ZN(n14307) );
  XNOR2_X1 U16194 ( .A(n14309), .B(n14307), .ZN(n14495) );
  INV_X1 U16195 ( .A(n14307), .ZN(n14308) );
  NAND2_X1 U16196 ( .A1(n14309), .A2(n14308), .ZN(n14310) );
  NAND2_X1 U16197 ( .A1(n14888), .A2(n14346), .ZN(n14312) );
  NAND2_X1 U16198 ( .A1(n14901), .A2(n14295), .ZN(n14311) );
  NAND2_X1 U16199 ( .A1(n14312), .A2(n14311), .ZN(n14313) );
  XNOR2_X1 U16200 ( .A(n14313), .B(n11660), .ZN(n14316) );
  AND2_X1 U16201 ( .A1(n14901), .A2(n10794), .ZN(n14314) );
  AOI21_X1 U16202 ( .B1(n14888), .B2(n14351), .A(n14314), .ZN(n14315) );
  OAI21_X1 U16203 ( .B1(n14316), .B2(n14315), .A(n14502), .ZN(n14427) );
  NAND2_X1 U16204 ( .A1(n15068), .A2(n14346), .ZN(n14318) );
  NAND2_X1 U16205 ( .A1(n14879), .A2(n14295), .ZN(n14317) );
  NAND2_X1 U16206 ( .A1(n14318), .A2(n14317), .ZN(n14319) );
  XNOR2_X1 U16207 ( .A(n14319), .B(n11660), .ZN(n14321) );
  AND2_X1 U16208 ( .A1(n14879), .A2(n10794), .ZN(n14320) );
  AOI21_X1 U16209 ( .B1(n15068), .B2(n14351), .A(n14320), .ZN(n14322) );
  NAND2_X1 U16210 ( .A1(n14321), .A2(n14322), .ZN(n14390) );
  INV_X1 U16211 ( .A(n14321), .ZN(n14324) );
  INV_X1 U16212 ( .A(n14322), .ZN(n14323) );
  NAND2_X1 U16213 ( .A1(n14324), .A2(n14323), .ZN(n14325) );
  NAND2_X1 U16214 ( .A1(n15061), .A2(n14346), .ZN(n14327) );
  NAND2_X1 U16215 ( .A1(n14571), .A2(n14351), .ZN(n14326) );
  NAND2_X1 U16216 ( .A1(n14327), .A2(n14326), .ZN(n14328) );
  XNOR2_X1 U16217 ( .A(n14328), .B(n11660), .ZN(n14330) );
  AND2_X1 U16218 ( .A1(n14571), .A2(n10794), .ZN(n14329) );
  AOI21_X1 U16219 ( .B1(n15061), .B2(n14351), .A(n14329), .ZN(n14331) );
  NAND2_X1 U16220 ( .A1(n14330), .A2(n14331), .ZN(n14482) );
  INV_X1 U16221 ( .A(n14330), .ZN(n14333) );
  INV_X1 U16222 ( .A(n14331), .ZN(n14332) );
  NAND2_X1 U16223 ( .A1(n14333), .A2(n14332), .ZN(n14334) );
  NAND2_X1 U16224 ( .A1(n14395), .A2(n14482), .ZN(n14345) );
  NAND2_X1 U16225 ( .A1(n14833), .A2(n14346), .ZN(n14337) );
  NAND2_X1 U16226 ( .A1(n14570), .A2(n14351), .ZN(n14336) );
  NAND2_X1 U16227 ( .A1(n14337), .A2(n14336), .ZN(n14338) );
  XNOR2_X1 U16228 ( .A(n14338), .B(n11660), .ZN(n14340) );
  AND2_X1 U16229 ( .A1(n14570), .A2(n10794), .ZN(n14339) );
  AOI21_X1 U16230 ( .B1(n14833), .B2(n14351), .A(n14339), .ZN(n14341) );
  NAND2_X1 U16231 ( .A1(n14340), .A2(n14341), .ZN(n14451) );
  INV_X1 U16232 ( .A(n14340), .ZN(n14343) );
  INV_X1 U16233 ( .A(n14341), .ZN(n14342) );
  NAND2_X1 U16234 ( .A1(n14343), .A2(n14342), .ZN(n14344) );
  NAND2_X1 U16235 ( .A1(n14345), .A2(n14483), .ZN(n14450) );
  NAND2_X1 U16236 ( .A1(n15050), .A2(n14346), .ZN(n14348) );
  NAND2_X1 U16237 ( .A1(n14569), .A2(n14295), .ZN(n14347) );
  NAND2_X1 U16238 ( .A1(n14348), .A2(n14347), .ZN(n14349) );
  XNOR2_X1 U16239 ( .A(n14349), .B(n11660), .ZN(n14352) );
  AND2_X1 U16240 ( .A1(n14569), .A2(n10794), .ZN(n14350) );
  AOI21_X1 U16241 ( .B1(n15050), .B2(n14351), .A(n14350), .ZN(n14353) );
  NAND2_X1 U16242 ( .A1(n14352), .A2(n14353), .ZN(n14358) );
  INV_X1 U16243 ( .A(n14352), .ZN(n14355) );
  INV_X1 U16244 ( .A(n14353), .ZN(n14354) );
  NAND2_X1 U16245 ( .A1(n14355), .A2(n14354), .ZN(n14356) );
  OAI22_X1 U16246 ( .A1(n15048), .A2(n14414), .B1(n14455), .B2(n14413), .ZN(
        n14360) );
  XNOR2_X1 U16247 ( .A(n14360), .B(n14359), .ZN(n14362) );
  OAI22_X1 U16248 ( .A1(n15048), .A2(n14413), .B1(n14455), .B2(n14411), .ZN(
        n14361) );
  NOR2_X1 U16249 ( .A1(n14362), .A2(n14361), .ZN(n14363) );
  AOI21_X1 U16250 ( .B1(n14362), .B2(n14361), .A(n14363), .ZN(n14539) );
  OAI22_X1 U16251 ( .A1(n14365), .A2(n14414), .B1(n14543), .B2(n14413), .ZN(
        n14364) );
  XNOR2_X1 U16252 ( .A(n14364), .B(n11660), .ZN(n14369) );
  INV_X1 U16253 ( .A(n14369), .ZN(n14371) );
  OR2_X1 U16254 ( .A1(n14365), .A2(n14413), .ZN(n14367) );
  NAND2_X1 U16255 ( .A1(n14567), .A2(n10794), .ZN(n14366) );
  INV_X1 U16256 ( .A(n14368), .ZN(n14370) );
  AOI21_X1 U16257 ( .B1(n14371), .B2(n14370), .A(n14422), .ZN(n14372) );
  NOR2_X1 U16258 ( .A1(n14373), .A2(n14372), .ZN(n14374) );
  OAI21_X1 U16259 ( .B1(n14417), .B2(n14374), .A(n14540), .ZN(n14381) );
  OAI22_X1 U16260 ( .A1(n14778), .A2(n14556), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14375), .ZN(n14376) );
  AOI21_X1 U16261 ( .B1(n14568), .B2(n14377), .A(n14376), .ZN(n14378) );
  OAI21_X1 U16262 ( .B1(n15033), .B2(n14555), .A(n14378), .ZN(n14379) );
  AOI21_X1 U16263 ( .B1(n14780), .B2(n10393), .A(n14379), .ZN(n14380) );
  NAND2_X1 U16264 ( .A1(n14381), .A2(n14380), .ZN(P1_U3214) );
  OAI21_X1 U16265 ( .B1(n6636), .B2(n14383), .A(n14382), .ZN(n14384) );
  NAND2_X1 U16266 ( .A1(n14384), .A2(n14540), .ZN(n14389) );
  AND2_X1 U16267 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14697) );
  INV_X1 U16268 ( .A(n15017), .ZN(n14385) );
  OAI22_X1 U16269 ( .A1(n14557), .A2(n14386), .B1(n14556), .B2(n14385), .ZN(
        n14387) );
  AOI211_X1 U16270 ( .C1(n14534), .C2(n15009), .A(n14697), .B(n14387), .ZN(
        n14388) );
  OAI211_X1 U16271 ( .C1(n15019), .C2(n14550), .A(n14389), .B(n14388), .ZN(
        P1_U3215) );
  INV_X1 U16272 ( .A(n14390), .ZN(n14391) );
  NOR2_X1 U16273 ( .A1(n14392), .A2(n14391), .ZN(n14396) );
  INV_X1 U16274 ( .A(n14395), .ZN(n14485) );
  AOI21_X1 U16275 ( .B1(n14396), .B2(n14394), .A(n14485), .ZN(n14402) );
  AND2_X1 U16276 ( .A1(n14879), .A2(n15010), .ZN(n14397) );
  AOI21_X1 U16277 ( .B1(n14570), .B2(n15008), .A(n14397), .ZN(n14840) );
  INV_X1 U16278 ( .A(n14843), .ZN(n14398) );
  AOI22_X1 U16279 ( .A1(n14398), .A2(n14418), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14399) );
  OAI21_X1 U16280 ( .B1(n14840), .B2(n14420), .A(n14399), .ZN(n14400) );
  AOI21_X1 U16281 ( .B1(n15061), .B2(n10393), .A(n14400), .ZN(n14401) );
  OAI21_X1 U16282 ( .B1(n14402), .B2(n14561), .A(n14401), .ZN(P1_U3216) );
  INV_X1 U16283 ( .A(n15088), .ZN(n14922) );
  AOI21_X1 U16284 ( .B1(n14404), .B2(n14403), .A(n14561), .ZN(n14406) );
  NAND2_X1 U16285 ( .A1(n14406), .A2(n14405), .ZN(n14410) );
  OAI22_X1 U16286 ( .A1(n14431), .A2(n14993), .B1(n14407), .B2(n15032), .ZN(
        n14916) );
  NAND2_X1 U16287 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14743)
         );
  OAI21_X1 U16288 ( .B1(n14919), .B2(n14556), .A(n14743), .ZN(n14408) );
  AOI21_X1 U16289 ( .B1(n14916), .B2(n14547), .A(n14408), .ZN(n14409) );
  OAI211_X1 U16290 ( .C1(n14922), .C2(n14550), .A(n14410), .B(n14409), .ZN(
        P1_U3219) );
  OAI22_X1 U16291 ( .A1(n14768), .A2(n14413), .B1(n15033), .B2(n14411), .ZN(
        n14412) );
  XNOR2_X1 U16292 ( .A(n14412), .B(n11660), .ZN(n14416) );
  OAI22_X1 U16293 ( .A1(n14768), .A2(n14414), .B1(n15033), .B2(n14413), .ZN(
        n14415) );
  XNOR2_X1 U16294 ( .A(n14416), .B(n14415), .ZN(n14423) );
  NAND3_X1 U16295 ( .A1(n14417), .A2(n14423), .A3(n14540), .ZN(n14426) );
  AOI22_X1 U16296 ( .A1(n15008), .A2(n14565), .B1(n14567), .B2(n15010), .ZN(
        n14759) );
  AOI22_X1 U16297 ( .A1(n14766), .A2(n14418), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14419) );
  OAI21_X1 U16298 ( .B1(n14759), .B2(n14420), .A(n14419), .ZN(n14421) );
  AOI21_X1 U16299 ( .B1(n15041), .B2(n10393), .A(n14421), .ZN(n14425) );
  NAND3_X1 U16300 ( .A1(n14423), .A2(n14540), .A3(n14422), .ZN(n14424) );
  AOI21_X1 U16301 ( .B1(n14428), .B2(n14427), .A(n6491), .ZN(n14435) );
  OAI22_X1 U16302 ( .A1(n14430), .A2(n14555), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14429), .ZN(n14433) );
  OAI22_X1 U16303 ( .A1(n14431), .A2(n14557), .B1(n14556), .B2(n14883), .ZN(
        n14432) );
  AOI211_X1 U16304 ( .C1(n14888), .C2(n10393), .A(n14433), .B(n14432), .ZN(
        n14434) );
  OAI21_X1 U16305 ( .B1(n14435), .B2(n14561), .A(n14434), .ZN(P1_U3223) );
  INV_X1 U16306 ( .A(n14516), .ZN(n14436) );
  XNOR2_X1 U16307 ( .A(n14439), .B(n14438), .ZN(n14514) );
  NOR3_X1 U16308 ( .A1(n14437), .A2(n14436), .A3(n14514), .ZN(n14519) );
  AOI21_X1 U16309 ( .B1(n14439), .B2(n14438), .A(n14519), .ZN(n14442) );
  OAI211_X1 U16310 ( .C1(n14442), .C2(n14441), .A(n14540), .B(n14440), .ZN(
        n14448) );
  OAI22_X1 U16311 ( .A1(n14557), .A2(n14444), .B1(n14443), .B2(n14556), .ZN(
        n14445) );
  AOI211_X1 U16312 ( .C1(n14534), .C2(n15011), .A(n14446), .B(n14445), .ZN(
        n14447) );
  OAI211_X1 U16313 ( .C1(n14449), .C2(n14550), .A(n14448), .B(n14447), .ZN(
        P1_U3224) );
  INV_X1 U16314 ( .A(n14450), .ZN(n14486) );
  NOR3_X1 U16315 ( .A1(n14486), .A2(n6730), .A3(n14452), .ZN(n14453) );
  OAI21_X1 U16316 ( .B1(n14453), .B2(n6574), .A(n14540), .ZN(n14460) );
  OAI22_X1 U16317 ( .A1(n14455), .A2(n14993), .B1(n14454), .B2(n15032), .ZN(
        n14804) );
  INV_X1 U16318 ( .A(n14808), .ZN(n14457) );
  OAI22_X1 U16319 ( .A1(n14457), .A2(n14556), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14456), .ZN(n14458) );
  AOI21_X1 U16320 ( .B1(n14804), .B2(n14547), .A(n14458), .ZN(n14459) );
  OAI211_X1 U16321 ( .C1(n14810), .C2(n14550), .A(n14460), .B(n14459), .ZN(
        P1_U3225) );
  NAND2_X1 U16322 ( .A1(n14462), .A2(n14461), .ZN(n14464) );
  OAI21_X1 U16323 ( .B1(n14462), .B2(n14461), .A(n14464), .ZN(n14552) );
  INV_X1 U16324 ( .A(n14463), .ZN(n14553) );
  NOR2_X1 U16325 ( .A1(n14552), .A2(n14553), .ZN(n14551) );
  INV_X1 U16326 ( .A(n14464), .ZN(n14465) );
  NOR3_X1 U16327 ( .A1(n14551), .A2(n14466), .A3(n14465), .ZN(n14467) );
  OAI21_X1 U16328 ( .B1(n14467), .B2(n6621), .A(n14540), .ZN(n14473) );
  INV_X1 U16329 ( .A(n14468), .ZN(n14471) );
  INV_X1 U16330 ( .A(n14469), .ZN(n14977) );
  OAI22_X1 U16331 ( .A1(n14557), .A2(n14966), .B1(n14977), .B2(n14556), .ZN(
        n14470) );
  AOI211_X1 U16332 ( .C1(n14534), .C2(n14572), .A(n14471), .B(n14470), .ZN(
        n14472) );
  OAI211_X1 U16333 ( .C1(n15105), .C2(n14550), .A(n14473), .B(n14472), .ZN(
        P1_U3226) );
  NOR3_X1 U16334 ( .A1(n6621), .A2(n14475), .A3(n14474), .ZN(n14476) );
  OAI21_X1 U16335 ( .B1(n6624), .B2(n14476), .A(n14540), .ZN(n14481) );
  INV_X1 U16336 ( .A(n14477), .ZN(n14479) );
  OAI22_X1 U16337 ( .A1(n14557), .A2(n14994), .B1(n14956), .B2(n14556), .ZN(
        n14478) );
  AOI211_X1 U16338 ( .C1(n14534), .C2(n14950), .A(n14479), .B(n14478), .ZN(
        n14480) );
  OAI211_X1 U16339 ( .C1(n14955), .C2(n14550), .A(n14481), .B(n14480), .ZN(
        P1_U3228) );
  INV_X1 U16340 ( .A(n14482), .ZN(n14484) );
  NOR3_X1 U16341 ( .A1(n14485), .A2(n14484), .A3(n14483), .ZN(n14487) );
  OAI21_X1 U16342 ( .B1(n14487), .B2(n14486), .A(n14540), .ZN(n14493) );
  AND2_X1 U16343 ( .A1(n14571), .A2(n15010), .ZN(n14488) );
  AOI21_X1 U16344 ( .B1(n14569), .B2(n15008), .A(n14488), .ZN(n14822) );
  INV_X1 U16345 ( .A(n14822), .ZN(n14491) );
  OAI22_X1 U16346 ( .A1(n14831), .A2(n14556), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14489), .ZN(n14490) );
  AOI21_X1 U16347 ( .B1(n14491), .B2(n14547), .A(n14490), .ZN(n14492) );
  OAI211_X1 U16348 ( .C1(n15057), .C2(n14550), .A(n14493), .B(n14492), .ZN(
        P1_U3229) );
  XNOR2_X1 U16349 ( .A(n14494), .B(n14495), .ZN(n14501) );
  OAI22_X1 U16350 ( .A1(n14507), .A2(n14555), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14496), .ZN(n14499) );
  INV_X1 U16351 ( .A(n14497), .ZN(n14905) );
  OAI22_X1 U16352 ( .A1(n14932), .A2(n14557), .B1(n14905), .B2(n14556), .ZN(
        n14498) );
  AOI211_X1 U16353 ( .C1(n14910), .C2(n10393), .A(n14499), .B(n14498), .ZN(
        n14500) );
  OAI21_X1 U16354 ( .B1(n14501), .B2(n14561), .A(n14500), .ZN(P1_U3233) );
  INV_X1 U16355 ( .A(n14502), .ZN(n14504) );
  NOR3_X1 U16356 ( .A1(n6491), .A2(n14504), .A3(n14503), .ZN(n14506) );
  INV_X1 U16357 ( .A(n14394), .ZN(n14505) );
  OAI21_X1 U16358 ( .B1(n14506), .B2(n14505), .A(n14540), .ZN(n14513) );
  OAI22_X1 U16359 ( .A1(n14508), .A2(n14993), .B1(n14507), .B2(n15032), .ZN(
        n14860) );
  INV_X1 U16360 ( .A(n14865), .ZN(n14510) );
  OAI22_X1 U16361 ( .A1(n14510), .A2(n14556), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14509), .ZN(n14511) );
  AOI21_X1 U16362 ( .B1(n14860), .B2(n14547), .A(n14511), .ZN(n14512) );
  OAI211_X1 U16363 ( .C1(n14550), .C2(n14867), .A(n14513), .B(n14512), .ZN(
        P1_U3235) );
  INV_X1 U16364 ( .A(n14514), .ZN(n14515) );
  AOI21_X1 U16365 ( .B1(n14517), .B2(n14516), .A(n14515), .ZN(n14518) );
  OAI21_X1 U16366 ( .B1(n14519), .B2(n14518), .A(n14540), .ZN(n14525) );
  OAI22_X1 U16367 ( .A1(n14557), .A2(n14521), .B1(n14556), .B2(n14520), .ZN(
        n14522) );
  AOI211_X1 U16368 ( .C1(n14534), .C2(n14574), .A(n14523), .B(n14522), .ZN(
        n14524) );
  OAI211_X1 U16369 ( .C1(n14526), .C2(n14550), .A(n14525), .B(n14524), .ZN(
        P1_U3236) );
  OAI21_X1 U16370 ( .B1(n14529), .B2(n14528), .A(n14527), .ZN(n14530) );
  NAND2_X1 U16371 ( .A1(n14530), .A2(n14540), .ZN(n14536) );
  NAND2_X1 U16372 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14717)
         );
  INV_X1 U16373 ( .A(n14717), .ZN(n14533) );
  INV_X1 U16374 ( .A(n14941), .ZN(n14531) );
  OAI22_X1 U16375 ( .A1(n14557), .A2(n14967), .B1(n14531), .B2(n14556), .ZN(
        n14532) );
  AOI211_X1 U16376 ( .C1(n14534), .C2(n14900), .A(n14533), .B(n14532), .ZN(
        n14535) );
  OAI211_X1 U16377 ( .C1(n15144), .C2(n14550), .A(n14536), .B(n14535), .ZN(
        P1_U3238) );
  OAI21_X1 U16378 ( .B1(n14539), .B2(n14538), .A(n14537), .ZN(n14541) );
  NAND2_X1 U16379 ( .A1(n14541), .A2(n14540), .ZN(n14549) );
  OAI22_X1 U16380 ( .A1(n14543), .A2(n14993), .B1(n14542), .B2(n15032), .ZN(
        n14790) );
  INV_X1 U16381 ( .A(n14794), .ZN(n14545) );
  OAI22_X1 U16382 ( .A1(n14545), .A2(n14556), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14544), .ZN(n14546) );
  AOI21_X1 U16383 ( .B1(n14790), .B2(n14547), .A(n14546), .ZN(n14548) );
  OAI211_X1 U16384 ( .C1(n15048), .C2(n14550), .A(n14549), .B(n14548), .ZN(
        P1_U3240) );
  AOI21_X1 U16385 ( .B1(n14553), .B2(n14552), .A(n14551), .ZN(n14562) );
  OAI21_X1 U16386 ( .B1(n14555), .B2(n14994), .A(n14554), .ZN(n14559) );
  OAI22_X1 U16387 ( .A1(n14557), .A2(n14992), .B1(n14998), .B2(n14556), .ZN(
        n14558) );
  AOI211_X1 U16388 ( .C1(n15107), .C2(n10393), .A(n14559), .B(n14558), .ZN(
        n14560) );
  OAI21_X1 U16389 ( .B1(n14562), .B2(n14561), .A(n14560), .ZN(P1_U3241) );
  MUX2_X1 U16390 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14563), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16391 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14564), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16392 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14565), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16393 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14566), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16394 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14567), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16395 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14568), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16396 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14569), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16397 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14570), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16398 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14571), .S(n14580), .Z(
        P1_U3583) );
  MUX2_X1 U16399 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14879), .S(n14580), .Z(
        P1_U3582) );
  MUX2_X1 U16400 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14901), .S(n14580), .Z(
        P1_U3581) );
  MUX2_X1 U16401 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14878), .S(n14580), .Z(
        P1_U3580) );
  MUX2_X1 U16402 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14900), .S(n14580), .Z(
        P1_U3579) );
  MUX2_X1 U16403 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14950), .S(n14580), .Z(
        P1_U3578) );
  MUX2_X1 U16404 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14572), .S(n14580), .Z(
        P1_U3577) );
  MUX2_X1 U16405 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n6981), .S(n14580), .Z(
        P1_U3576) );
  MUX2_X1 U16406 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15009), .S(n14580), .Z(
        P1_U3575) );
  MUX2_X1 U16407 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14573), .S(n14580), .Z(
        P1_U3574) );
  MUX2_X1 U16408 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15011), .S(n14580), .Z(
        P1_U3573) );
  MUX2_X1 U16409 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14574), .S(n14580), .Z(
        P1_U3572) );
  MUX2_X1 U16410 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14575), .S(n14580), .Z(
        P1_U3571) );
  MUX2_X1 U16411 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14576), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16412 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14577), .S(n14580), .Z(
        P1_U3569) );
  MUX2_X1 U16413 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14578), .S(n14580), .Z(
        P1_U3568) );
  MUX2_X1 U16414 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14579), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16415 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14581), .S(n14580), .Z(
        P1_U3566) );
  MUX2_X1 U16416 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14582), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16417 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14583), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16418 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14584), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16419 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14585), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16420 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10474), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16421 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14587), .S(P1_U4016), .Z(
        P1_U3560) );
  INV_X1 U16422 ( .A(n14588), .ZN(n14591) );
  OAI211_X1 U16423 ( .C1(n14591), .C2(n14590), .A(n14733), .B(n14589), .ZN(
        n14599) );
  OAI211_X1 U16424 ( .C1(n14594), .C2(n14593), .A(n14739), .B(n14592), .ZN(
        n14598) );
  AOI22_X1 U16425 ( .A1(n15269), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14597) );
  NAND2_X1 U16426 ( .A1(n14737), .A2(n14595), .ZN(n14596) );
  NAND4_X1 U16427 ( .A1(n14599), .A2(n14598), .A3(n14597), .A4(n14596), .ZN(
        P1_U3244) );
  OAI211_X1 U16428 ( .C1(n14601), .C2(n14600), .A(n14739), .B(n14621), .ZN(
        n14611) );
  MUX2_X1 U16429 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11031), .S(n14606), .Z(
        n14604) );
  NAND3_X1 U16430 ( .A1(n14604), .A2(n14603), .A3(n14602), .ZN(n14605) );
  NAND3_X1 U16431 ( .A1(n14733), .A2(n14616), .A3(n14605), .ZN(n14610) );
  INV_X1 U16432 ( .A(n14606), .ZN(n14607) );
  NAND2_X1 U16433 ( .A1(n14737), .A2(n14607), .ZN(n14609) );
  AOI22_X1 U16434 ( .A1(n15269), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n14608) );
  NAND4_X1 U16435 ( .A1(n14611), .A2(n14610), .A3(n14609), .A4(n14608), .ZN(
        P1_U3246) );
  NAND2_X1 U16436 ( .A1(n15269), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n14612) );
  OAI211_X1 U16437 ( .C1(n14719), .C2(n14619), .A(n14613), .B(n14612), .ZN(
        n14614) );
  INV_X1 U16438 ( .A(n14614), .ZN(n14627) );
  MUX2_X1 U16439 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10900), .S(n14619), .Z(
        n14617) );
  NAND3_X1 U16440 ( .A1(n14617), .A2(n14616), .A3(n14615), .ZN(n14618) );
  NAND3_X1 U16441 ( .A1(n14733), .A2(n14638), .A3(n14618), .ZN(n14626) );
  MUX2_X1 U16442 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10318), .S(n14619), .Z(
        n14622) );
  NAND3_X1 U16443 ( .A1(n14622), .A2(n14621), .A3(n14620), .ZN(n14623) );
  NAND3_X1 U16444 ( .A1(n14739), .A2(n14624), .A3(n14623), .ZN(n14625) );
  NAND4_X1 U16445 ( .A1(n14628), .A2(n14627), .A3(n14626), .A4(n14625), .ZN(
        P1_U3247) );
  OAI21_X1 U16446 ( .B1(n14745), .B2(n10300), .A(n14629), .ZN(n14630) );
  AOI21_X1 U16447 ( .B1(n14635), .B2(n14737), .A(n14630), .ZN(n14642) );
  OAI21_X1 U16448 ( .B1(n14633), .B2(n14632), .A(n14631), .ZN(n14634) );
  NAND2_X1 U16449 ( .A1(n14739), .A2(n14634), .ZN(n14641) );
  MUX2_X1 U16450 ( .A(n10351), .B(P1_REG2_REG_5__SCAN_IN), .S(n14635), .Z(
        n14636) );
  NAND3_X1 U16451 ( .A1(n14638), .A2(n14637), .A3(n14636), .ZN(n14639) );
  NAND3_X1 U16452 ( .A1(n14733), .A2(n14651), .A3(n14639), .ZN(n14640) );
  NAND3_X1 U16453 ( .A1(n14642), .A2(n14641), .A3(n14640), .ZN(P1_U3248) );
  OAI21_X1 U16454 ( .B1(n14745), .B2(n14644), .A(n14643), .ZN(n14645) );
  AOI21_X1 U16455 ( .B1(n14648), .B2(n14737), .A(n14645), .ZN(n14655) );
  OAI211_X1 U16456 ( .C1(n14647), .C2(n14646), .A(n14739), .B(n14661), .ZN(
        n14654) );
  MUX2_X1 U16457 ( .A(n11426), .B(P1_REG2_REG_6__SCAN_IN), .S(n14648), .Z(
        n14649) );
  NAND3_X1 U16458 ( .A1(n14651), .A2(n14650), .A3(n14649), .ZN(n14652) );
  NAND3_X1 U16459 ( .A1(n14733), .A2(n14667), .A3(n14652), .ZN(n14653) );
  NAND3_X1 U16460 ( .A1(n14655), .A2(n14654), .A3(n14653), .ZN(P1_U3249) );
  OAI21_X1 U16461 ( .B1(n14745), .B2(n14657), .A(n14656), .ZN(n14658) );
  AOI21_X1 U16462 ( .B1(n14664), .B2(n14737), .A(n14658), .ZN(n14672) );
  MUX2_X1 U16463 ( .A(n10330), .B(P1_REG1_REG_7__SCAN_IN), .S(n14664), .Z(
        n14659) );
  NAND3_X1 U16464 ( .A1(n14661), .A2(n14660), .A3(n14659), .ZN(n14662) );
  NAND3_X1 U16465 ( .A1(n14739), .A2(n14663), .A3(n14662), .ZN(n14671) );
  MUX2_X1 U16466 ( .A(n11592), .B(P1_REG2_REG_7__SCAN_IN), .S(n14664), .Z(
        n14665) );
  NAND3_X1 U16467 ( .A1(n14667), .A2(n14666), .A3(n14665), .ZN(n14668) );
  NAND3_X1 U16468 ( .A1(n14733), .A2(n14669), .A3(n14668), .ZN(n14670) );
  NAND3_X1 U16469 ( .A1(n14672), .A2(n14671), .A3(n14670), .ZN(P1_U3250) );
  OAI21_X1 U16470 ( .B1(n14675), .B2(n14674), .A(n14673), .ZN(n14676) );
  NAND2_X1 U16471 ( .A1(n14676), .A2(n14739), .ZN(n14688) );
  INV_X1 U16472 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14678) );
  OAI21_X1 U16473 ( .B1(n14745), .B2(n14678), .A(n14677), .ZN(n14679) );
  AOI21_X1 U16474 ( .B1(n14680), .B2(n14737), .A(n14679), .ZN(n14687) );
  MUX2_X1 U16475 ( .A(n11771), .B(P1_REG2_REG_9__SCAN_IN), .S(n14680), .Z(
        n14681) );
  NAND3_X1 U16476 ( .A1(n14683), .A2(n14682), .A3(n14681), .ZN(n14684) );
  NAND3_X1 U16477 ( .A1(n14685), .A2(n14733), .A3(n14684), .ZN(n14686) );
  NAND3_X1 U16478 ( .A1(n14688), .A2(n14687), .A3(n14686), .ZN(P1_U3252) );
  INV_X1 U16479 ( .A(n14689), .ZN(n14694) );
  AOI21_X1 U16480 ( .B1(n14692), .B2(n14691), .A(n14690), .ZN(n14693) );
  OAI21_X1 U16481 ( .B1(n14694), .B2(n14693), .A(n14739), .ZN(n14706) );
  NOR2_X1 U16482 ( .A1(n14719), .A2(n14695), .ZN(n14696) );
  AOI211_X1 U16483 ( .C1(n15269), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n14697), 
        .B(n14696), .ZN(n14705) );
  MUX2_X1 U16484 ( .A(n11521), .B(P1_REG2_REG_14__SCAN_IN), .S(n14698), .Z(
        n14699) );
  NAND3_X1 U16485 ( .A1(n14701), .A2(n14700), .A3(n14699), .ZN(n14702) );
  NAND3_X1 U16486 ( .A1(n14703), .A2(n14733), .A3(n14702), .ZN(n14704) );
  NAND3_X1 U16487 ( .A1(n14706), .A2(n14705), .A3(n14704), .ZN(P1_U3257) );
  NAND2_X1 U16488 ( .A1(n14707), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14708) );
  NAND2_X1 U16489 ( .A1(n14709), .A2(n14708), .ZN(n14728) );
  XNOR2_X1 U16490 ( .A(n14728), .B(n14718), .ZN(n14726) );
  XNOR2_X1 U16491 ( .A(n14726), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14723) );
  INV_X1 U16492 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15094) );
  INV_X1 U16493 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14711) );
  OAI22_X1 U16494 ( .A1(n14713), .A2(n14712), .B1(n14711), .B2(n14710), .ZN(
        n14725) );
  INV_X1 U16495 ( .A(n14725), .ZN(n14714) );
  XNOR2_X1 U16496 ( .A(n14714), .B(n14727), .ZN(n14724) );
  XNOR2_X1 U16497 ( .A(n15094), .B(n14724), .ZN(n14715) );
  NAND2_X1 U16498 ( .A1(n14739), .A2(n14715), .ZN(n14716) );
  NAND2_X1 U16499 ( .A1(n14717), .A2(n14716), .ZN(n14721) );
  NOR2_X1 U16500 ( .A1(n14719), .A2(n14718), .ZN(n14720) );
  AOI211_X1 U16501 ( .C1(n15269), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n14721), 
        .B(n14720), .ZN(n14722) );
  OAI21_X1 U16502 ( .B1(n14723), .B2(n14735), .A(n14722), .ZN(P1_U3261) );
  INV_X1 U16503 ( .A(n14740), .ZN(n14734) );
  NAND2_X1 U16504 ( .A1(n14726), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14730) );
  NAND2_X1 U16505 ( .A1(n14728), .A2(n14727), .ZN(n14729) );
  NAND2_X1 U16506 ( .A1(n14730), .A2(n14729), .ZN(n14732) );
  INV_X1 U16507 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14731) );
  XNOR2_X1 U16508 ( .A(n14732), .B(n14731), .ZN(n14736) );
  AOI22_X1 U16509 ( .A1(n14734), .A2(n14739), .B1(n14733), .B2(n14736), .ZN(
        n14742) );
  NOR2_X1 U16510 ( .A1(n14736), .A2(n14735), .ZN(n14738) );
  AOI211_X1 U16511 ( .C1(n14740), .C2(n14739), .A(n14738), .B(n14737), .ZN(
        n14741) );
  MUX2_X1 U16512 ( .A(n14742), .B(n14741), .S(n15296), .Z(n14744) );
  OAI211_X1 U16513 ( .C1(n7785), .C2(n14745), .A(n14744), .B(n14743), .ZN(
        P1_U3262) );
  NOR2_X1 U16514 ( .A1(n15305), .A2(n14746), .ZN(n14747) );
  NOR2_X1 U16515 ( .A1(n15307), .A2(n15027), .ZN(n14754) );
  AOI211_X1 U16516 ( .C1(n14748), .C2(n14980), .A(n14747), .B(n14754), .ZN(
        n14749) );
  OAI21_X1 U16517 ( .B1(n14750), .B2(n14984), .A(n14749), .ZN(P1_U3263) );
  OAI211_X1 U16518 ( .C1(n14752), .C2(n15124), .A(n6432), .B(n14751), .ZN(
        n15028) );
  NOR2_X1 U16519 ( .A1(n15305), .A2(n14753), .ZN(n14755) );
  AOI211_X1 U16520 ( .C1(n14756), .C2(n14980), .A(n14755), .B(n14754), .ZN(
        n14757) );
  OAI21_X1 U16521 ( .B1(n15028), .B2(n14984), .A(n14757), .ZN(P1_U3264) );
  INV_X1 U16522 ( .A(n14759), .ZN(n14760) );
  OAI211_X1 U16523 ( .C1(n14763), .C2(n14768), .A(n6432), .B(n14762), .ZN(
        n15043) );
  INV_X1 U16524 ( .A(n15043), .ZN(n14774) );
  NOR2_X1 U16525 ( .A1(n15305), .A2(n14764), .ZN(n14765) );
  AOI21_X1 U16526 ( .B1(n14766), .B2(n15301), .A(n14765), .ZN(n14767) );
  OAI21_X1 U16527 ( .B1(n14768), .B2(n15279), .A(n14767), .ZN(n14773) );
  NAND2_X1 U16528 ( .A1(n14771), .A2(n14770), .ZN(n15040) );
  AND3_X1 U16529 ( .A1(n14769), .A2(n15282), .A3(n15040), .ZN(n14772) );
  OAI21_X1 U16530 ( .B1(n15044), .B2(n15307), .A(n14775), .ZN(P1_U3265) );
  NAND2_X1 U16531 ( .A1(n14776), .A2(n15305), .ZN(n14782) );
  OAI22_X1 U16532 ( .A1(n14778), .A2(n14997), .B1(n14777), .B2(n15305), .ZN(
        n14779) );
  AOI21_X1 U16533 ( .B1(n14780), .B2(n14980), .A(n14779), .ZN(n14781) );
  OAI211_X1 U16534 ( .C1(n14984), .C2(n14783), .A(n14782), .B(n14781), .ZN(
        P1_U3266) );
  XNOR2_X1 U16535 ( .A(n14784), .B(n14787), .ZN(n14791) );
  OAI211_X1 U16536 ( .C1(n14787), .C2(n14786), .A(n14785), .B(n15078), .ZN(
        n14788) );
  INV_X1 U16537 ( .A(n14788), .ZN(n14789) );
  AOI211_X2 U16538 ( .C1(n14791), .C2(n14874), .A(n14790), .B(n14789), .ZN(
        n15047) );
  OAI21_X1 U16539 ( .B1(n14806), .B2(n15048), .A(n6432), .ZN(n14792) );
  INV_X1 U16540 ( .A(n15046), .ZN(n14797) );
  AOI22_X1 U16541 ( .A1(n14794), .A2(n15301), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15307), .ZN(n14795) );
  OAI21_X1 U16542 ( .B1(n15048), .B2(n15279), .A(n14795), .ZN(n14796) );
  AOI21_X1 U16543 ( .B1(n14797), .B2(n15273), .A(n14796), .ZN(n14798) );
  OAI21_X1 U16544 ( .B1(n15047), .B2(n15307), .A(n14798), .ZN(P1_U3267) );
  NAND2_X1 U16545 ( .A1(n14800), .A2(n14799), .ZN(n14818) );
  NOR2_X1 U16546 ( .A1(n14818), .A2(n14817), .ZN(n14821) );
  NOR2_X1 U16547 ( .A1(n14821), .A2(n14801), .ZN(n14803) );
  XNOR2_X1 U16548 ( .A(n14803), .B(n14802), .ZN(n14805) );
  AOI21_X1 U16549 ( .B1(n14805), .B2(n14874), .A(n14804), .ZN(n15052) );
  INV_X1 U16550 ( .A(n14828), .ZN(n14807) );
  AOI211_X1 U16551 ( .C1(n15050), .C2(n14807), .A(n15015), .B(n14806), .ZN(
        n15049) );
  AOI22_X1 U16552 ( .A1(n14808), .A2(n15301), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15307), .ZN(n14809) );
  OAI21_X1 U16553 ( .B1(n14810), .B2(n15279), .A(n14809), .ZN(n14815) );
  OAI21_X1 U16554 ( .B1(n14813), .B2(n14812), .A(n14811), .ZN(n15053) );
  NOR2_X1 U16555 ( .A1(n15053), .A2(n15023), .ZN(n14814) );
  AOI211_X1 U16556 ( .C1(n15049), .C2(n15273), .A(n14815), .B(n14814), .ZN(
        n14816) );
  OAI21_X1 U16557 ( .B1(n15052), .B2(n15307), .A(n14816), .ZN(P1_U3268) );
  NAND2_X1 U16558 ( .A1(n14818), .A2(n14817), .ZN(n14819) );
  NAND2_X1 U16559 ( .A1(n14819), .A2(n14874), .ZN(n14820) );
  OR2_X1 U16560 ( .A1(n14821), .A2(n14820), .ZN(n14823) );
  NAND2_X1 U16561 ( .A1(n14823), .A2(n14822), .ZN(n15059) );
  INV_X1 U16562 ( .A(n15059), .ZN(n14837) );
  NAND2_X1 U16563 ( .A1(n14825), .A2(n14824), .ZN(n14826) );
  NAND2_X1 U16564 ( .A1(n6570), .A2(n14826), .ZN(n15054) );
  NAND2_X1 U16565 ( .A1(n14844), .A2(n14833), .ZN(n14827) );
  NAND2_X1 U16566 ( .A1(n14827), .A2(n6432), .ZN(n14829) );
  OR2_X1 U16567 ( .A1(n14829), .A2(n14828), .ZN(n15055) );
  OAI22_X1 U16568 ( .A1(n14831), .A2(n14997), .B1(n14830), .B2(n15305), .ZN(
        n14832) );
  AOI21_X1 U16569 ( .B1(n14833), .B2(n14980), .A(n14832), .ZN(n14834) );
  OAI21_X1 U16570 ( .B1(n15055), .B2(n14984), .A(n14834), .ZN(n14835) );
  AOI21_X1 U16571 ( .B1(n15054), .B2(n15282), .A(n14835), .ZN(n14836) );
  OAI21_X1 U16572 ( .B1(n14837), .B2(n15307), .A(n14836), .ZN(P1_U3269) );
  XNOR2_X1 U16573 ( .A(n14838), .B(n14849), .ZN(n14839) );
  NAND2_X1 U16574 ( .A1(n14839), .A2(n14874), .ZN(n14841) );
  NAND2_X1 U16575 ( .A1(n14841), .A2(n14840), .ZN(n15066) );
  INV_X1 U16576 ( .A(n15066), .ZN(n14854) );
  OAI22_X1 U16577 ( .A1(n14843), .A2(n14997), .B1(n14842), .B2(n15305), .ZN(
        n14847) );
  AOI21_X1 U16578 ( .B1(n14862), .B2(n15061), .A(n15015), .ZN(n14845) );
  NAND2_X1 U16579 ( .A1(n14845), .A2(n14844), .ZN(n15062) );
  NOR2_X1 U16580 ( .A1(n15062), .A2(n14984), .ZN(n14846) );
  AOI211_X1 U16581 ( .C1(n14980), .C2(n15061), .A(n14847), .B(n14846), .ZN(
        n14853) );
  INV_X1 U16582 ( .A(n14848), .ZN(n14850) );
  NAND2_X1 U16583 ( .A1(n14850), .A2(n14849), .ZN(n15060) );
  NAND3_X1 U16584 ( .A1(n15060), .A2(n15282), .A3(n14851), .ZN(n14852) );
  OAI211_X1 U16585 ( .C1(n14854), .C2(n15307), .A(n14853), .B(n14852), .ZN(
        P1_U3270) );
  INV_X1 U16586 ( .A(n14897), .ZN(n14855) );
  NAND2_X1 U16587 ( .A1(n14855), .A2(n14911), .ZN(n14899) );
  INV_X1 U16588 ( .A(n14856), .ZN(n14892) );
  AOI21_X1 U16589 ( .B1(n14899), .B2(n14873), .A(n14892), .ZN(n14877) );
  INV_X1 U16590 ( .A(n14857), .ZN(n14858) );
  OAI21_X1 U16591 ( .B1(n14877), .B2(n14858), .A(n14869), .ZN(n14859) );
  AOI21_X1 U16592 ( .B1(n14861), .B2(n14874), .A(n14860), .ZN(n15070) );
  INV_X1 U16593 ( .A(n14885), .ZN(n14864) );
  INV_X1 U16594 ( .A(n14862), .ZN(n14863) );
  AOI211_X1 U16595 ( .C1(n15068), .C2(n14864), .A(n15015), .B(n14863), .ZN(
        n15067) );
  AOI22_X1 U16596 ( .A1(n14865), .A2(n15301), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15307), .ZN(n14866) );
  OAI21_X1 U16597 ( .B1(n14867), .B2(n15279), .A(n14866), .ZN(n14871) );
  XNOR2_X1 U16598 ( .A(n14869), .B(n14868), .ZN(n15071) );
  NOR2_X1 U16599 ( .A1(n15071), .A2(n15023), .ZN(n14870) );
  AOI211_X1 U16600 ( .C1(n15067), .C2(n15273), .A(n14871), .B(n14870), .ZN(
        n14872) );
  OAI21_X1 U16601 ( .B1(n15070), .B2(n15307), .A(n14872), .ZN(P1_U3271) );
  NAND3_X1 U16602 ( .A1(n14899), .A2(n14892), .A3(n14873), .ZN(n14875) );
  NAND2_X1 U16603 ( .A1(n14875), .A2(n14874), .ZN(n14876) );
  OR2_X1 U16604 ( .A1(n14877), .A2(n14876), .ZN(n14881) );
  AOI22_X1 U16605 ( .A1(n14879), .A2(n15008), .B1(n15010), .B2(n14878), .ZN(
        n14880) );
  OAI22_X1 U16606 ( .A1(n14883), .A2(n14997), .B1(n14882), .B2(n15305), .ZN(
        n14887) );
  OAI21_X1 U16607 ( .B1(n14907), .B2(n15135), .A(n6432), .ZN(n14884) );
  OR2_X1 U16608 ( .A1(n14885), .A2(n14884), .ZN(n15072) );
  NOR2_X1 U16609 ( .A1(n15072), .A2(n14984), .ZN(n14886) );
  AOI211_X1 U16610 ( .C1(n14980), .C2(n14888), .A(n14887), .B(n14886), .ZN(
        n14895) );
  INV_X1 U16611 ( .A(n14889), .ZN(n14890) );
  NAND2_X1 U16612 ( .A1(n14890), .A2(n14896), .ZN(n15079) );
  NAND2_X1 U16613 ( .A1(n15079), .A2(n14891), .ZN(n14893) );
  XNOR2_X1 U16614 ( .A(n14893), .B(n14892), .ZN(n15074) );
  OR2_X1 U16615 ( .A1(n15074), .A2(n15023), .ZN(n14894) );
  OAI211_X1 U16616 ( .C1(n15073), .C2(n15307), .A(n14895), .B(n14894), .ZN(
        P1_U3272) );
  AOI21_X1 U16617 ( .B1(n14897), .B2(n14896), .A(n14988), .ZN(n14898) );
  NAND2_X1 U16618 ( .A1(n14899), .A2(n14898), .ZN(n14903) );
  AOI22_X1 U16619 ( .A1(n15008), .A2(n14901), .B1(n14900), .B2(n15010), .ZN(
        n14902) );
  NAND2_X1 U16620 ( .A1(n14903), .A2(n14902), .ZN(n15084) );
  INV_X1 U16621 ( .A(n15084), .ZN(n14914) );
  OAI22_X1 U16622 ( .A1(n14905), .A2(n14997), .B1(n14904), .B2(n15305), .ZN(
        n14909) );
  OAI21_X1 U16623 ( .B1(n14918), .B2(n15082), .A(n6432), .ZN(n14906) );
  OR2_X1 U16624 ( .A1(n14907), .A2(n14906), .ZN(n15080) );
  NOR2_X1 U16625 ( .A1(n15080), .A2(n14984), .ZN(n14908) );
  AOI211_X1 U16626 ( .C1(n14980), .C2(n14910), .A(n14909), .B(n14908), .ZN(
        n14913) );
  NAND2_X1 U16627 ( .A1(n14889), .A2(n14911), .ZN(n15077) );
  NAND3_X1 U16628 ( .A1(n15079), .A2(n15282), .A3(n15077), .ZN(n14912) );
  OAI211_X1 U16629 ( .C1(n14914), .C2(n15307), .A(n14913), .B(n14912), .ZN(
        P1_U3273) );
  OAI21_X1 U16630 ( .B1(n6598), .B2(n14924), .A(n14915), .ZN(n14917) );
  AOI21_X1 U16631 ( .B1(n14917), .B2(n14874), .A(n14916), .ZN(n15090) );
  AOI211_X1 U16632 ( .C1(n15088), .C2(n14937), .A(n15015), .B(n14918), .ZN(
        n15087) );
  INV_X1 U16633 ( .A(n14919), .ZN(n14920) );
  AOI22_X1 U16634 ( .A1(n14920), .A2(n15301), .B1(P1_REG2_REG_19__SCAN_IN), 
        .B2(n15307), .ZN(n14921) );
  OAI21_X1 U16635 ( .B1(n14922), .B2(n15279), .A(n14921), .ZN(n14926) );
  XNOR2_X1 U16636 ( .A(n14923), .B(n14924), .ZN(n15091) );
  NOR2_X1 U16637 ( .A1(n15091), .A2(n15023), .ZN(n14925) );
  AOI211_X1 U16638 ( .C1(n15087), .C2(n15273), .A(n14926), .B(n14925), .ZN(
        n14927) );
  OAI21_X1 U16639 ( .B1(n15090), .B2(n15307), .A(n14927), .ZN(P1_U3274) );
  XNOR2_X1 U16640 ( .A(n14928), .B(n14929), .ZN(n14936) );
  OAI211_X1 U16641 ( .C1(n14931), .C2(n6905), .A(n14930), .B(n14874), .ZN(
        n14935) );
  OAI22_X1 U16642 ( .A1(n14932), .A2(n14993), .B1(n14967), .B2(n15032), .ZN(
        n14933) );
  INV_X1 U16643 ( .A(n14933), .ZN(n14934) );
  OAI211_X1 U16644 ( .C1(n14936), .C2(n15314), .A(n14935), .B(n14934), .ZN(
        n15093) );
  INV_X1 U16645 ( .A(n15093), .ZN(n14945) );
  INV_X1 U16646 ( .A(n14953), .ZN(n14939) );
  INV_X1 U16647 ( .A(n14937), .ZN(n14938) );
  AOI211_X1 U16648 ( .C1(n14940), .C2(n14939), .A(n15015), .B(n14938), .ZN(
        n15092) );
  AOI22_X1 U16649 ( .A1(n15307), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14941), 
        .B2(n15301), .ZN(n14942) );
  OAI21_X1 U16650 ( .B1(n15144), .B2(n15279), .A(n14942), .ZN(n14943) );
  AOI21_X1 U16651 ( .B1(n15092), .B2(n15273), .A(n14943), .ZN(n14944) );
  OAI21_X1 U16652 ( .B1(n14945), .B2(n15307), .A(n14944), .ZN(P1_U3275) );
  XNOR2_X1 U16653 ( .A(n14946), .B(n14948), .ZN(n15101) );
  OAI211_X1 U16654 ( .C1(n14949), .C2(n14948), .A(n14947), .B(n14874), .ZN(
        n14952) );
  AOI22_X1 U16655 ( .A1(n14950), .A2(n15008), .B1(n15010), .B2(n6981), .ZN(
        n14951) );
  NAND2_X1 U16656 ( .A1(n14952), .A2(n14951), .ZN(n15097) );
  NAND2_X1 U16657 ( .A1(n15097), .A2(n15305), .ZN(n14961) );
  INV_X1 U16658 ( .A(n14964), .ZN(n14954) );
  AOI211_X1 U16659 ( .C1(n15099), .C2(n14954), .A(n15015), .B(n14953), .ZN(
        n15098) );
  NOR2_X1 U16660 ( .A1(n14955), .A2(n15279), .ZN(n14959) );
  OAI22_X1 U16661 ( .A1(n15305), .A2(n14957), .B1(n14956), .B2(n14997), .ZN(
        n14958) );
  AOI211_X1 U16662 ( .C1(n15098), .C2(n15273), .A(n14959), .B(n14958), .ZN(
        n14960) );
  OAI211_X1 U16663 ( .C1(n15101), .C2(n15023), .A(n14961), .B(n14960), .ZN(
        P1_U3276) );
  NAND2_X1 U16664 ( .A1(n15000), .A2(n14981), .ZN(n14963) );
  NAND2_X1 U16665 ( .A1(n14963), .A2(n6432), .ZN(n14965) );
  OAI22_X1 U16666 ( .A1(n14967), .A2(n14993), .B1(n14966), .B2(n15032), .ZN(
        n14976) );
  INV_X1 U16667 ( .A(n14968), .ZN(n14970) );
  NOR2_X1 U16668 ( .A1(n14970), .A2(n14969), .ZN(n14971) );
  OAI22_X1 U16669 ( .A1(n6521), .A2(n14988), .B1(n14971), .B2(n15314), .ZN(
        n14974) );
  INV_X1 U16670 ( .A(n14971), .ZN(n14972) );
  NOR2_X1 U16671 ( .A1(n14972), .A2(n15314), .ZN(n14973) );
  MUX2_X1 U16672 ( .A(n14974), .B(n14973), .S(n8337), .Z(n14975) );
  AOI211_X1 U16673 ( .C1(n6536), .C2(n14874), .A(n14976), .B(n14975), .ZN(
        n15103) );
  OR2_X1 U16674 ( .A1(n15103), .A2(n15307), .ZN(n14983) );
  INV_X1 U16675 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14978) );
  OAI22_X1 U16676 ( .A1(n15305), .A2(n14978), .B1(n14977), .B2(n14997), .ZN(
        n14979) );
  AOI21_X1 U16677 ( .B1(n14981), .B2(n14980), .A(n14979), .ZN(n14982) );
  OAI211_X1 U16678 ( .C1(n15102), .C2(n14984), .A(n14983), .B(n14982), .ZN(
        P1_U3277) );
  NAND2_X1 U16679 ( .A1(n15022), .A2(n14986), .ZN(n14987) );
  XNOR2_X1 U16680 ( .A(n14987), .B(n14989), .ZN(n15110) );
  AOI21_X1 U16681 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14996) );
  OAI22_X1 U16682 ( .A1(n14994), .A2(n14993), .B1(n14992), .B2(n15032), .ZN(
        n14995) );
  AOI21_X1 U16683 ( .B1(n14996), .B2(n7428), .A(n14995), .ZN(n15109) );
  OAI21_X1 U16684 ( .B1(n14998), .B2(n14997), .A(n15109), .ZN(n14999) );
  NAND2_X1 U16685 ( .A1(n14999), .A2(n15305), .ZN(n15006) );
  AOI21_X1 U16686 ( .B1(n15013), .B2(n15107), .A(n15015), .ZN(n15001) );
  AND2_X1 U16687 ( .A1(n15001), .A2(n15000), .ZN(n15106) );
  OAI22_X1 U16688 ( .A1(n15003), .A2(n15279), .B1(n15002), .B2(n15305), .ZN(
        n15004) );
  AOI21_X1 U16689 ( .B1(n15106), .B2(n15273), .A(n15004), .ZN(n15005) );
  OAI211_X1 U16690 ( .C1(n15110), .C2(n15023), .A(n15006), .B(n15005), .ZN(
        P1_U3278) );
  XOR2_X1 U16691 ( .A(n15007), .B(n15020), .Z(n15012) );
  AOI222_X1 U16692 ( .A1(n14874), .A2(n15012), .B1(n15011), .B2(n15010), .C1(
        n15009), .C2(n15008), .ZN(n15114) );
  INV_X1 U16693 ( .A(n15013), .ZN(n15014) );
  AOI211_X1 U16694 ( .C1(n15112), .C2(n15016), .A(n15015), .B(n15014), .ZN(
        n15111) );
  AOI22_X1 U16695 ( .A1(n15307), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n15017), 
        .B2(n15301), .ZN(n15018) );
  OAI21_X1 U16696 ( .B1(n15019), .B2(n15279), .A(n15018), .ZN(n15025) );
  NAND2_X1 U16697 ( .A1(n14985), .A2(n15020), .ZN(n15021) );
  NAND2_X1 U16698 ( .A1(n15022), .A2(n15021), .ZN(n15115) );
  NOR2_X1 U16699 ( .A1(n15115), .A2(n15023), .ZN(n15024) );
  AOI211_X1 U16700 ( .C1(n15111), .C2(n15273), .A(n15025), .B(n15024), .ZN(
        n15026) );
  OAI21_X1 U16701 ( .B1(n15114), .B2(n15307), .A(n15026), .ZN(P1_U3279) );
  INV_X1 U16702 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n15029) );
  AND2_X1 U16703 ( .A1(n15028), .A2(n15027), .ZN(n15121) );
  MUX2_X1 U16704 ( .A(n15029), .B(n15121), .S(n15322), .Z(n15030) );
  OAI21_X1 U16705 ( .B1(n15124), .B2(n15096), .A(n15030), .ZN(P1_U3558) );
  OAI21_X1 U16706 ( .B1(n15033), .B2(n15032), .A(n15031), .ZN(n15035) );
  MUX2_X1 U16707 ( .A(n15125), .B(P1_REG1_REG_29__SCAN_IN), .S(n15320), .Z(
        P1_U3557) );
  NAND3_X1 U16708 ( .A1(n14769), .A2(n15078), .A3(n15040), .ZN(n15045) );
  NAND2_X1 U16709 ( .A1(n15041), .A2(n15311), .ZN(n15042) );
  MUX2_X1 U16710 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15126), .S(n15322), .Z(
        P1_U3556) );
  INV_X1 U16711 ( .A(n15311), .ZN(n15104) );
  OAI211_X1 U16712 ( .C1(n15048), .C2(n15104), .A(n15047), .B(n15046), .ZN(
        n15127) );
  MUX2_X1 U16713 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15127), .S(n15322), .Z(
        P1_U3554) );
  AOI21_X1 U16714 ( .B1(n15311), .B2(n15050), .A(n15049), .ZN(n15051) );
  OAI211_X1 U16715 ( .C1(n15314), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        n15128) );
  MUX2_X1 U16716 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15128), .S(n15322), .Z(
        P1_U3553) );
  NAND2_X1 U16717 ( .A1(n15054), .A2(n15078), .ZN(n15056) );
  OAI211_X1 U16718 ( .C1(n15057), .C2(n15104), .A(n15056), .B(n15055), .ZN(
        n15058) );
  MUX2_X1 U16719 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15129), .S(n15322), .Z(
        P1_U3552) );
  NAND3_X1 U16720 ( .A1(n15060), .A2(n15078), .A3(n14851), .ZN(n15064) );
  NAND2_X1 U16721 ( .A1(n15061), .A2(n15311), .ZN(n15063) );
  NAND3_X1 U16722 ( .A1(n15064), .A2(n15063), .A3(n15062), .ZN(n15065) );
  MUX2_X1 U16723 ( .A(n15130), .B(P1_REG1_REG_23__SCAN_IN), .S(n15320), .Z(
        P1_U3551) );
  AOI21_X1 U16724 ( .B1(n15311), .B2(n15068), .A(n15067), .ZN(n15069) );
  OAI211_X1 U16725 ( .C1(n15314), .C2(n15071), .A(n15070), .B(n15069), .ZN(
        n15131) );
  MUX2_X1 U16726 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15131), .S(n15322), .Z(
        P1_U3550) );
  OAI211_X1 U16727 ( .C1(n15074), .C2(n15314), .A(n15073), .B(n15072), .ZN(
        n15132) );
  MUX2_X1 U16728 ( .A(n15132), .B(P1_REG1_REG_21__SCAN_IN), .S(n15320), .Z(
        n15075) );
  INV_X1 U16729 ( .A(n15075), .ZN(n15076) );
  OAI21_X1 U16730 ( .B1(n15135), .B2(n15096), .A(n15076), .ZN(P1_U3549) );
  INV_X1 U16731 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15085) );
  NAND3_X1 U16732 ( .A1(n15079), .A2(n15078), .A3(n15077), .ZN(n15081) );
  OAI211_X1 U16733 ( .C1(n15082), .C2(n15104), .A(n15081), .B(n15080), .ZN(
        n15083) );
  NOR2_X1 U16734 ( .A1(n15084), .A2(n15083), .ZN(n15136) );
  MUX2_X1 U16735 ( .A(n15085), .B(n15136), .S(n15322), .Z(n15086) );
  INV_X1 U16736 ( .A(n15086), .ZN(P1_U3548) );
  AOI21_X1 U16737 ( .B1(n15311), .B2(n15088), .A(n15087), .ZN(n15089) );
  OAI211_X1 U16738 ( .C1(n15314), .C2(n15091), .A(n15090), .B(n15089), .ZN(
        n15139) );
  MUX2_X1 U16739 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15139), .S(n15322), .Z(
        P1_U3547) );
  NOR2_X1 U16740 ( .A1(n15093), .A2(n15092), .ZN(n15141) );
  MUX2_X1 U16741 ( .A(n15141), .B(n15094), .S(n15320), .Z(n15095) );
  OAI21_X1 U16742 ( .B1(n15144), .B2(n15096), .A(n15095), .ZN(P1_U3546) );
  AOI211_X1 U16743 ( .C1(n15311), .C2(n15099), .A(n15098), .B(n15097), .ZN(
        n15100) );
  OAI21_X1 U16744 ( .B1(n15314), .B2(n15101), .A(n15100), .ZN(n15145) );
  MUX2_X1 U16745 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15145), .S(n15322), .Z(
        P1_U3545) );
  OAI211_X1 U16746 ( .C1(n15105), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        n15146) );
  MUX2_X1 U16747 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15146), .S(n15322), .Z(
        P1_U3544) );
  AOI21_X1 U16748 ( .B1(n15311), .B2(n15107), .A(n15106), .ZN(n15108) );
  OAI211_X1 U16749 ( .C1(n15110), .C2(n15314), .A(n15109), .B(n15108), .ZN(
        n15147) );
  MUX2_X1 U16750 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15147), .S(n15322), .Z(
        P1_U3543) );
  AOI21_X1 U16751 ( .B1(n15311), .B2(n15112), .A(n15111), .ZN(n15113) );
  OAI211_X1 U16752 ( .C1(n15314), .C2(n15115), .A(n15114), .B(n15113), .ZN(
        n15148) );
  MUX2_X1 U16753 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15148), .S(n15322), .Z(
        P1_U3542) );
  AOI21_X1 U16754 ( .B1(n15311), .B2(n15117), .A(n15116), .ZN(n15118) );
  OAI211_X1 U16755 ( .C1(n15314), .C2(n15120), .A(n15119), .B(n15118), .ZN(
        n15149) );
  MUX2_X1 U16756 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15149), .S(n15322), .Z(
        P1_U3539) );
  INV_X1 U16757 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15122) );
  MUX2_X1 U16758 ( .A(n15122), .B(n15121), .S(n15319), .Z(n15123) );
  OAI21_X1 U16759 ( .B1(n15124), .B2(n15143), .A(n15123), .ZN(P1_U3526) );
  MUX2_X1 U16760 ( .A(n15125), .B(P1_REG0_REG_29__SCAN_IN), .S(n15317), .Z(
        P1_U3525) );
  MUX2_X1 U16761 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15126), .S(n15319), .Z(
        P1_U3524) );
  MUX2_X1 U16762 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15127), .S(n15319), .Z(
        P1_U3522) );
  MUX2_X1 U16763 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15128), .S(n15319), .Z(
        P1_U3521) );
  MUX2_X1 U16764 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15129), .S(n15319), .Z(
        P1_U3520) );
  MUX2_X1 U16765 ( .A(n15130), .B(P1_REG0_REG_23__SCAN_IN), .S(n15317), .Z(
        P1_U3519) );
  MUX2_X1 U16766 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15131), .S(n15319), .Z(
        P1_U3518) );
  MUX2_X1 U16767 ( .A(n15132), .B(P1_REG0_REG_21__SCAN_IN), .S(n15317), .Z(
        n15133) );
  INV_X1 U16768 ( .A(n15133), .ZN(n15134) );
  OAI21_X1 U16769 ( .B1(n15135), .B2(n15143), .A(n15134), .ZN(P1_U3517) );
  INV_X1 U16770 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15137) );
  MUX2_X1 U16771 ( .A(n15137), .B(n15136), .S(n15319), .Z(n15138) );
  INV_X1 U16772 ( .A(n15138), .ZN(P1_U3516) );
  MUX2_X1 U16773 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15139), .S(n15319), .Z(
        P1_U3515) );
  INV_X1 U16774 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n15140) );
  MUX2_X1 U16775 ( .A(n15141), .B(n15140), .S(n15317), .Z(n15142) );
  OAI21_X1 U16776 ( .B1(n15144), .B2(n15143), .A(n15142), .ZN(P1_U3513) );
  MUX2_X1 U16777 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15145), .S(n15319), .Z(
        P1_U3510) );
  MUX2_X1 U16778 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15146), .S(n15319), .Z(
        P1_U3507) );
  MUX2_X1 U16779 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15147), .S(n15319), .Z(
        P1_U3504) );
  MUX2_X1 U16780 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15148), .S(n15319), .Z(
        P1_U3501) );
  MUX2_X1 U16781 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15149), .S(n15319), .Z(
        P1_U3492) );
  NOR4_X1 U16782 ( .A1(n15152), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15151), .A4(
        P1_U3086), .ZN(n15153) );
  AOI21_X1 U16783 ( .B1(n15154), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15153), 
        .ZN(n15155) );
  OAI21_X1 U16784 ( .B1(n15156), .B2(n15159), .A(n15155), .ZN(P1_U3324) );
  OAI222_X1 U16785 ( .A1(P1_U3086), .A2(n15160), .B1(n15159), .B2(n15158), 
        .C1(n15157), .C2(n15165), .ZN(P1_U3326) );
  NAND2_X1 U16786 ( .A1(n15162), .A2(n15161), .ZN(n15164) );
  OAI211_X1 U16787 ( .C1(n15166), .C2(n15165), .A(n15164), .B(n15163), .ZN(
        P1_U3328) );
  MUX2_X1 U16788 ( .A(n15167), .B(n8371), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16789 ( .A(n15168), .ZN(n15169) );
  MUX2_X1 U16790 ( .A(n15169), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U16791 ( .A(n15171), .B(n15170), .Z(SUB_1596_U57) );
  XOR2_X1 U16792 ( .A(n15172), .B(n15173), .Z(SUB_1596_U56) );
  XOR2_X1 U16793 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n15174), .Z(SUB_1596_U54) );
  INV_X1 U16794 ( .A(n15176), .ZN(n15177) );
  NAND2_X1 U16795 ( .A1(n15178), .A2(n15177), .ZN(n15179) );
  INV_X1 U16796 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15183) );
  NAND2_X1 U16797 ( .A1(n15183), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n15195) );
  NAND2_X1 U16798 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15184), .ZN(n15193) );
  NAND2_X1 U16799 ( .A1(n15195), .A2(n15193), .ZN(n15185) );
  XNOR2_X1 U16800 ( .A(n15194), .B(n15185), .ZN(n15187) );
  INV_X1 U16801 ( .A(n15187), .ZN(n15186) );
  NAND2_X1 U16802 ( .A1(n15188), .A2(n15187), .ZN(n15191) );
  NAND2_X1 U16803 ( .A1(n15190), .A2(n15191), .ZN(n15189) );
  XNOR2_X1 U16804 ( .A(n15189), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  INV_X1 U16805 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15403) );
  NAND2_X1 U16806 ( .A1(n15190), .A2(n15403), .ZN(n15192) );
  NAND2_X1 U16807 ( .A1(n15194), .A2(n15193), .ZN(n15196) );
  NAND2_X1 U16808 ( .A1(n15196), .A2(n15195), .ZN(n15201) );
  INV_X1 U16809 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U16810 ( .A1(n15197), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n15209) );
  INV_X1 U16811 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15198) );
  NAND2_X1 U16812 ( .A1(n15198), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15199) );
  AND2_X1 U16813 ( .A1(n15209), .A2(n15199), .ZN(n15200) );
  NAND2_X1 U16814 ( .A1(n15201), .A2(n15200), .ZN(n15210) );
  OR2_X1 U16815 ( .A1(n15201), .A2(n15200), .ZN(n15202) );
  AND2_X1 U16816 ( .A1(n15210), .A2(n15202), .ZN(n15203) );
  INV_X1 U16817 ( .A(n15208), .ZN(n15205) );
  NAND2_X1 U16818 ( .A1(n15205), .A2(n15207), .ZN(n15206) );
  XNOR2_X1 U16819 ( .A(n15206), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  NAND2_X1 U16820 ( .A1(n15210), .A2(n15209), .ZN(n15218) );
  INV_X1 U16821 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15219) );
  XNOR2_X1 U16822 ( .A(n15219), .B(P3_ADDR_REG_15__SCAN_IN), .ZN(n15211) );
  XNOR2_X1 U16823 ( .A(n15218), .B(n15211), .ZN(n15215) );
  XNOR2_X1 U16824 ( .A(n15215), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(n15212) );
  XNOR2_X1 U16825 ( .A(n15213), .B(n15212), .ZN(SUB_1596_U65) );
  INV_X1 U16826 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15214) );
  INV_X1 U16827 ( .A(n15215), .ZN(n15216) );
  OR2_X1 U16828 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15219), .ZN(n15217) );
  NAND2_X1 U16829 ( .A1(n15218), .A2(n15217), .ZN(n15221) );
  NAND2_X1 U16830 ( .A1(n15219), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n15220) );
  NAND2_X1 U16831 ( .A1(n15221), .A2(n15220), .ZN(n15228) );
  XOR2_X1 U16832 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .Z(n15222) );
  XNOR2_X1 U16833 ( .A(n15228), .B(n15222), .ZN(n15223) );
  NAND2_X1 U16834 ( .A1(n6578), .A2(n15225), .ZN(n15224) );
  XNOR2_X1 U16835 ( .A(n15224), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  INV_X1 U16836 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15230) );
  INV_X1 U16837 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15226) );
  NOR2_X1 U16838 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15226), .ZN(n15227) );
  OAI21_X1 U16839 ( .B1(n15230), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n15229), 
        .ZN(n15236) );
  XNOR2_X1 U16840 ( .A(n15236), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n15235) );
  XNOR2_X1 U16841 ( .A(n15235), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15231) );
  NAND2_X1 U16842 ( .A1(n15232), .A2(n15231), .ZN(n15234) );
  NAND2_X1 U16843 ( .A1(n7303), .A2(n15234), .ZN(n15233) );
  XNOR2_X1 U16844 ( .A(n15233), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  INV_X1 U16845 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15247) );
  NAND2_X1 U16846 ( .A1(n15247), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n15248) );
  OAI21_X1 U16847 ( .B1(n15247), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n15248), 
        .ZN(n15239) );
  INV_X1 U16848 ( .A(n15235), .ZN(n15238) );
  NOR2_X1 U16849 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15236), .ZN(n15237) );
  AOI21_X1 U16850 ( .B1(n15238), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n15237), 
        .ZN(n15251) );
  XOR2_X1 U16851 ( .A(n15239), .B(n15251), .Z(n15240) );
  AOI21_X1 U16852 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15242), .A(n15246), 
        .ZN(n15243) );
  INV_X1 U16853 ( .A(n15243), .ZN(SUB_1596_U62) );
  INV_X1 U16854 ( .A(n15244), .ZN(n15245) );
  OR2_X1 U16855 ( .A1(n15247), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n15250) );
  INV_X1 U16856 ( .A(n15248), .ZN(n15249) );
  AOI21_X1 U16857 ( .B1(n15251), .B2(n15250), .A(n15249), .ZN(n15254) );
  XNOR2_X1 U16858 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15252) );
  XNOR2_X1 U16859 ( .A(n15252), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n15253) );
  AOI21_X1 U16860 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15255) );
  OAI21_X1 U16861 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15255), 
        .ZN(U28) );
  AOI21_X1 U16862 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15256) );
  OAI21_X1 U16863 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15256), 
        .ZN(U29) );
  AND2_X1 U16864 ( .A1(n15258), .A2(n15257), .ZN(n15260) );
  XNOR2_X1 U16865 ( .A(n15260), .B(n15259), .ZN(SUB_1596_U61) );
  NOR2_X1 U16866 ( .A1(n15261), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15263) );
  OR2_X1 U16867 ( .A1(n15262), .A2(n15263), .ZN(n15266) );
  INV_X1 U16868 ( .A(n15263), .ZN(n15265) );
  MUX2_X1 U16869 ( .A(n15266), .B(n15265), .S(n15264), .Z(n15268) );
  NAND2_X1 U16870 ( .A1(n15268), .A2(n15267), .ZN(n15271) );
  AOI22_X1 U16871 ( .A1(n15269), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15270) );
  OAI21_X1 U16872 ( .B1(n15272), .B2(n15271), .A(n15270), .ZN(P1_U3243) );
  NAND2_X1 U16873 ( .A1(n15274), .A2(n15273), .ZN(n15278) );
  INV_X1 U16874 ( .A(n15275), .ZN(n15276) );
  AOI22_X1 U16875 ( .A1(n15307), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n15276), 
        .B2(n15301), .ZN(n15277) );
  OAI211_X1 U16876 ( .C1(n15280), .C2(n15279), .A(n15278), .B(n15277), .ZN(
        n15281) );
  AOI21_X1 U16877 ( .B1(n15283), .B2(n15282), .A(n15281), .ZN(n15284) );
  OAI21_X1 U16878 ( .B1(n15307), .B2(n15285), .A(n15284), .ZN(P1_U3285) );
  AOI21_X1 U16879 ( .B1(n15301), .B2(P1_REG3_REG_1__SCAN_IN), .A(n15286), .ZN(
        n15295) );
  INV_X1 U16880 ( .A(n15287), .ZN(n15290) );
  NAND2_X1 U16881 ( .A1(n15288), .A2(n8398), .ZN(n15289) );
  OAI211_X1 U16882 ( .C1(n15292), .C2(n15291), .A(n15290), .B(n15289), .ZN(
        n15293) );
  NOR2_X1 U16883 ( .A1(n15307), .A2(n15293), .ZN(n15294) );
  AOI22_X1 U16884 ( .A1(n10342), .A2(n15307), .B1(n15295), .B2(n15294), .ZN(
        P1_U3292) );
  NAND2_X1 U16885 ( .A1(n15297), .A2(n15296), .ZN(n15299) );
  AOI21_X1 U16886 ( .B1(n15300), .B2(n15299), .A(n15298), .ZN(n15306) );
  INV_X1 U16887 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U16888 ( .A1(n15302), .A2(n15305), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n15301), .ZN(n15303) );
  OAI221_X1 U16889 ( .B1(n15307), .B2(n15306), .C1(n15305), .C2(n15304), .A(
        n15303), .ZN(P1_U3293) );
  AND2_X1 U16890 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15308), .ZN(P1_U3294) );
  AND2_X1 U16891 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15308), .ZN(P1_U3295) );
  AND2_X1 U16892 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15308), .ZN(P1_U3296) );
  AND2_X1 U16893 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15308), .ZN(P1_U3297) );
  AND2_X1 U16894 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15308), .ZN(P1_U3298) );
  AND2_X1 U16895 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15308), .ZN(P1_U3299) );
  AND2_X1 U16896 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15308), .ZN(P1_U3300) );
  AND2_X1 U16897 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15308), .ZN(P1_U3301) );
  AND2_X1 U16898 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15308), .ZN(P1_U3302) );
  AND2_X1 U16899 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15308), .ZN(P1_U3303) );
  AND2_X1 U16900 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15308), .ZN(P1_U3304) );
  AND2_X1 U16901 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15308), .ZN(P1_U3305) );
  AND2_X1 U16902 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15308), .ZN(P1_U3306) );
  AND2_X1 U16903 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15308), .ZN(P1_U3307) );
  AND2_X1 U16904 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15308), .ZN(P1_U3308) );
  AND2_X1 U16905 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15308), .ZN(P1_U3309) );
  AND2_X1 U16906 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15308), .ZN(P1_U3310) );
  AND2_X1 U16907 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15308), .ZN(P1_U3311) );
  AND2_X1 U16908 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15308), .ZN(P1_U3312) );
  AND2_X1 U16909 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15308), .ZN(P1_U3313) );
  AND2_X1 U16910 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15308), .ZN(P1_U3314) );
  AND2_X1 U16911 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15308), .ZN(P1_U3315) );
  AND2_X1 U16912 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15308), .ZN(P1_U3316) );
  AND2_X1 U16913 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15308), .ZN(P1_U3317) );
  AND2_X1 U16914 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15308), .ZN(P1_U3318) );
  AND2_X1 U16915 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15308), .ZN(P1_U3319) );
  AND2_X1 U16916 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15308), .ZN(P1_U3320) );
  AND2_X1 U16917 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15308), .ZN(P1_U3321) );
  AND2_X1 U16918 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15308), .ZN(P1_U3322) );
  AND2_X1 U16919 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15308), .ZN(P1_U3323) );
  AOI21_X1 U16920 ( .B1(n15311), .B2(n6430), .A(n15309), .ZN(n15312) );
  OAI211_X1 U16921 ( .C1(n15315), .C2(n15314), .A(n15313), .B(n15312), .ZN(
        n15316) );
  INV_X1 U16922 ( .A(n15316), .ZN(n15321) );
  INV_X1 U16923 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15318) );
  AOI22_X1 U16924 ( .A1(n15319), .A2(n15321), .B1(n15318), .B2(n15317), .ZN(
        P1_U3471) );
  AOI22_X1 U16925 ( .A1(n15322), .A2(n15321), .B1(n10318), .B2(n15320), .ZN(
        P1_U3532) );
  NOR2_X1 U16926 ( .A1(n15373), .A2(P2_U3947), .ZN(P2_U3087) );
  OR2_X1 U16927 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15323), .ZN(n15347) );
  OAI21_X1 U16928 ( .B1(n15325), .B2(n15324), .A(n15347), .ZN(n15331) );
  AOI211_X1 U16929 ( .C1(n15329), .C2(n15328), .A(n15327), .B(n15326), .ZN(
        n15330) );
  AOI211_X1 U16930 ( .C1(n15471), .C2(n15332), .A(n15331), .B(n15330), .ZN(
        n15333) );
  OAI21_X1 U16931 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n15334), .A(n15333), .ZN(
        P2_U3190) );
  OAI21_X1 U16932 ( .B1(n15361), .B2(n15335), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15336) );
  OAI21_X1 U16933 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15336), .ZN(n15346) );
  OAI211_X1 U16934 ( .C1(n15339), .C2(n15338), .A(n15423), .B(n15337), .ZN(
        n15345) );
  NAND2_X1 U16935 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15373), .ZN(n15344) );
  NOR2_X1 U16936 ( .A1(n6914), .A2(n10635), .ZN(n15342) );
  OAI211_X1 U16937 ( .C1(n15342), .C2(n15341), .A(n15419), .B(n15340), .ZN(
        n15343) );
  NAND4_X1 U16938 ( .A1(n15346), .A2(n15345), .A3(n15344), .A4(n15343), .ZN(
        P2_U3215) );
  OAI21_X1 U16939 ( .B1(n15408), .B2(n15348), .A(n15347), .ZN(n15349) );
  AOI21_X1 U16940 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15373), .A(n15349), .ZN(
        n15359) );
  OAI211_X1 U16941 ( .C1(n15352), .C2(n15351), .A(n15423), .B(n15350), .ZN(
        n15358) );
  NAND2_X1 U16942 ( .A1(n15354), .A2(n15353), .ZN(n15355) );
  NAND3_X1 U16943 ( .A1(n15419), .A2(n15356), .A3(n15355), .ZN(n15357) );
  NAND3_X1 U16944 ( .A1(n15359), .A2(n15358), .A3(n15357), .ZN(P2_U3217) );
  OAI21_X1 U16945 ( .B1(n15361), .B2(n15360), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15362) );
  OAI21_X1 U16946 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15362), .ZN(n15372) );
  OAI211_X1 U16947 ( .C1(n15365), .C2(n15364), .A(n15419), .B(n15363), .ZN(
        n15371) );
  OAI211_X1 U16948 ( .C1(n15368), .C2(n15367), .A(n15423), .B(n15366), .ZN(
        n15370) );
  NAND2_X1 U16949 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15373), .ZN(n15369) );
  NAND4_X1 U16950 ( .A1(n15372), .A2(n15371), .A3(n15370), .A4(n15369), .ZN(
        P2_U3218) );
  NAND2_X1 U16951 ( .A1(n15373), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n15376) );
  INV_X1 U16952 ( .A(n15374), .ZN(n15375) );
  OAI211_X1 U16953 ( .C1(n15408), .C2(n15377), .A(n15376), .B(n15375), .ZN(
        n15378) );
  INV_X1 U16954 ( .A(n15378), .ZN(n15388) );
  AOI211_X1 U16955 ( .C1(n15381), .C2(n15380), .A(n15392), .B(n15379), .ZN(
        n15382) );
  INV_X1 U16956 ( .A(n15382), .ZN(n15387) );
  OAI211_X1 U16957 ( .C1(n15385), .C2(n15384), .A(n15423), .B(n15383), .ZN(
        n15386) );
  NAND3_X1 U16958 ( .A1(n15388), .A2(n15387), .A3(n15386), .ZN(P2_U3221) );
  OR2_X1 U16959 ( .A1(n15390), .A2(n15389), .ZN(n15393) );
  AOI211_X1 U16960 ( .C1(n15394), .C2(n15393), .A(n15392), .B(n15391), .ZN(
        n15395) );
  AOI211_X1 U16961 ( .C1(n15421), .C2(n15397), .A(n15396), .B(n15395), .ZN(
        n15402) );
  OAI211_X1 U16962 ( .C1(n15400), .C2(n15399), .A(n15398), .B(n15423), .ZN(
        n15401) );
  OAI211_X1 U16963 ( .C1(n15427), .C2(n15403), .A(n15402), .B(n15401), .ZN(
        P2_U3227) );
  XOR2_X1 U16964 ( .A(n15405), .B(n15404), .Z(n15410) );
  OAI21_X1 U16965 ( .B1(n15408), .B2(n15407), .A(n15406), .ZN(n15409) );
  AOI21_X1 U16966 ( .B1(n15410), .B2(n15419), .A(n15409), .ZN(n15414) );
  XOR2_X1 U16967 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n15411), .Z(n15412) );
  NAND2_X1 U16968 ( .A1(n15412), .A2(n15423), .ZN(n15413) );
  OAI211_X1 U16969 ( .C1(n15427), .C2(n7308), .A(n15414), .B(n15413), .ZN(
        P2_U3228) );
  INV_X1 U16970 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15428) );
  NAND2_X1 U16971 ( .A1(n15415), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n15416) );
  NAND2_X1 U16972 ( .A1(n15417), .A2(n15416), .ZN(n15424) );
  XOR2_X1 U16973 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n15418), .Z(n15420) );
  AOI222_X1 U16974 ( .A1(n15424), .A2(n15423), .B1(n15422), .B2(n15421), .C1(
        n15420), .C2(n15419), .ZN(n15426) );
  OAI211_X1 U16975 ( .C1(n15428), .C2(n15427), .A(n15426), .B(n15425), .ZN(
        P2_U3232) );
  XNOR2_X1 U16976 ( .A(n15430), .B(n15429), .ZN(n15432) );
  AOI21_X1 U16977 ( .B1(n15432), .B2(n15479), .A(n15431), .ZN(n15483) );
  NOR2_X1 U16978 ( .A1(n15434), .A2(n15433), .ZN(n15435) );
  AOI21_X1 U16979 ( .B1(n6438), .B2(P2_REG2_REG_4__SCAN_IN), .A(n15435), .ZN(
        n15436) );
  OAI21_X1 U16980 ( .B1(n15437), .B2(n15482), .A(n15436), .ZN(n15438) );
  INV_X1 U16981 ( .A(n15438), .ZN(n15448) );
  XNOR2_X1 U16982 ( .A(n15440), .B(n15439), .ZN(n15486) );
  OR2_X1 U16983 ( .A1(n15441), .A2(n15482), .ZN(n15442) );
  AND3_X1 U16984 ( .A1(n15444), .A2(n15443), .A3(n15442), .ZN(n15480) );
  AOI22_X1 U16985 ( .A1(n15486), .A2(n15446), .B1(n15445), .B2(n15480), .ZN(
        n15447) );
  OAI211_X1 U16986 ( .C1(n6438), .C2(n15483), .A(n15448), .B(n15447), .ZN(
        P2_U3261) );
  AND2_X1 U16987 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15455), .ZN(P2_U3266) );
  AND2_X1 U16988 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15455), .ZN(P2_U3267) );
  AND2_X1 U16989 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15455), .ZN(P2_U3268) );
  AND2_X1 U16990 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15455), .ZN(P2_U3269) );
  AND2_X1 U16991 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15455), .ZN(P2_U3270) );
  AND2_X1 U16992 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15455), .ZN(P2_U3271) );
  AND2_X1 U16993 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15455), .ZN(P2_U3272) );
  AND2_X1 U16994 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15455), .ZN(P2_U3273) );
  AND2_X1 U16995 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15455), .ZN(P2_U3274) );
  AND2_X1 U16996 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15455), .ZN(P2_U3275) );
  AND2_X1 U16997 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15455), .ZN(P2_U3276) );
  AND2_X1 U16998 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15455), .ZN(P2_U3277) );
  INV_X1 U16999 ( .A(n15455), .ZN(n15454) );
  NOR2_X1 U17000 ( .A1(n15454), .A2(n15450), .ZN(P2_U3278) );
  AND2_X1 U17001 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15455), .ZN(P2_U3279) );
  AND2_X1 U17002 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15455), .ZN(P2_U3280) );
  AND2_X1 U17003 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15455), .ZN(P2_U3281) );
  NOR2_X1 U17004 ( .A1(n15454), .A2(n15451), .ZN(P2_U3282) );
  AND2_X1 U17005 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15455), .ZN(P2_U3283) );
  AND2_X1 U17006 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15455), .ZN(P2_U3284) );
  AND2_X1 U17007 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15455), .ZN(P2_U3285) );
  AND2_X1 U17008 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15455), .ZN(P2_U3286) );
  AND2_X1 U17009 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15455), .ZN(P2_U3287) );
  AND2_X1 U17010 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15455), .ZN(P2_U3288) );
  AND2_X1 U17011 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15455), .ZN(P2_U3289) );
  INV_X1 U17012 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15452) );
  NOR2_X1 U17013 ( .A1(n15454), .A2(n15452), .ZN(P2_U3290) );
  AND2_X1 U17014 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15455), .ZN(P2_U3291) );
  NOR2_X1 U17015 ( .A1(n15454), .A2(n15453), .ZN(P2_U3292) );
  AND2_X1 U17016 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15455), .ZN(P2_U3293) );
  AND2_X1 U17017 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15455), .ZN(P2_U3294) );
  AND2_X1 U17018 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15455), .ZN(P2_U3295) );
  INV_X1 U17019 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15457) );
  OAI21_X1 U17020 ( .B1(n15459), .B2(n15457), .A(n15456), .ZN(P2_U3416) );
  INV_X1 U17021 ( .A(n15458), .ZN(n15460) );
  OAI22_X1 U17022 ( .A1(n15461), .A2(n15460), .B1(P2_D_REG_1__SCAN_IN), .B2(
        n15459), .ZN(n15462) );
  INV_X1 U17023 ( .A(n15462), .ZN(P2_U3417) );
  AND2_X1 U17024 ( .A1(n8826), .A2(n15463), .ZN(n15468) );
  OAI211_X1 U17025 ( .C1(n15490), .C2(n15466), .A(n15465), .B(n15464), .ZN(
        n15467) );
  AOI211_X1 U17026 ( .C1(n15469), .C2(n15479), .A(n15468), .B(n15467), .ZN(
        n15497) );
  AOI22_X1 U17027 ( .A1(n15496), .A2(n15497), .B1(n8449), .B2(n6954), .ZN(
        P2_U3433) );
  AOI21_X1 U17028 ( .B1(n15472), .B2(n15471), .A(n15470), .ZN(n15474) );
  OAI211_X1 U17029 ( .C1(n15476), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        n15477) );
  AOI21_X1 U17030 ( .B1(n15479), .B2(n15478), .A(n15477), .ZN(n15498) );
  AOI22_X1 U17031 ( .A1(n15496), .A2(n15498), .B1(n8484), .B2(n6954), .ZN(
        P2_U3439) );
  INV_X1 U17032 ( .A(n15480), .ZN(n15481) );
  OAI21_X1 U17033 ( .B1(n15482), .B2(n15490), .A(n15481), .ZN(n15485) );
  INV_X1 U17034 ( .A(n15483), .ZN(n15484) );
  AOI211_X1 U17035 ( .C1(n15486), .C2(n8826), .A(n15485), .B(n15484), .ZN(
        n15499) );
  INV_X1 U17036 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15487) );
  AOI22_X1 U17037 ( .A1(n15496), .A2(n15499), .B1(n15487), .B2(n6954), .ZN(
        P2_U3442) );
  INV_X1 U17038 ( .A(n15488), .ZN(n15489) );
  OAI21_X1 U17039 ( .B1(n15491), .B2(n15490), .A(n15489), .ZN(n15492) );
  AOI211_X1 U17040 ( .C1(n15495), .C2(n15494), .A(n15493), .B(n15492), .ZN(
        n15501) );
  AOI22_X1 U17041 ( .A1(n15496), .A2(n15501), .B1(n8535), .B2(n6954), .ZN(
        P2_U3448) );
  AOI22_X1 U17042 ( .A1(n15502), .A2(n15497), .B1(n10423), .B2(n15500), .ZN(
        P2_U3500) );
  AOI22_X1 U17043 ( .A1(n15502), .A2(n15498), .B1(n10484), .B2(n15500), .ZN(
        P2_U3502) );
  AOI22_X1 U17044 ( .A1(n15502), .A2(n15499), .B1(n10485), .B2(n15500), .ZN(
        P2_U3503) );
  AOI22_X1 U17045 ( .A1(n15502), .A2(n15501), .B1(n8540), .B2(n15500), .ZN(
        P2_U3505) );
  NOR2_X1 U17046 ( .A1(P3_U3897), .A2(n15503), .ZN(P3_U3150) );
  XNOR2_X1 U17047 ( .A(n15505), .B(n15504), .ZN(n15515) );
  INV_X1 U17048 ( .A(n15515), .ZN(n15597) );
  XNOR2_X1 U17049 ( .A(n15507), .B(n15506), .ZN(n15513) );
  OAI22_X1 U17050 ( .A1(n15511), .A2(n15510), .B1(n15509), .B2(n15508), .ZN(
        n15512) );
  AOI21_X1 U17051 ( .B1(n15513), .B2(n10147), .A(n15512), .ZN(n15514) );
  OAI21_X1 U17052 ( .B1(n15551), .B2(n15515), .A(n15514), .ZN(n15594) );
  AOI21_X1 U17053 ( .B1(n15538), .B2(n15597), .A(n15594), .ZN(n15522) );
  NOR2_X1 U17054 ( .A1(n15516), .A2(n15541), .ZN(n15595) );
  AOI22_X1 U17055 ( .A1(n15519), .A2(n15595), .B1(n15518), .B2(n15517), .ZN(
        n15520) );
  OAI221_X1 U17056 ( .B1(n15561), .B2(n15522), .C1(n15559), .C2(n15521), .A(
        n15520), .ZN(P3_U3224) );
  XNOR2_X1 U17057 ( .A(n15523), .B(n15528), .ZN(n15536) );
  INV_X1 U17058 ( .A(n15536), .ZN(n15568) );
  NOR2_X1 U17059 ( .A1(n15541), .A2(n15524), .ZN(n15567) );
  INV_X1 U17060 ( .A(n15567), .ZN(n15525) );
  OAI22_X1 U17061 ( .A1(n15553), .A2(n15527), .B1(n15526), .B2(n15525), .ZN(
        n15537) );
  XNOR2_X1 U17062 ( .A(n15528), .B(n15529), .ZN(n15530) );
  NAND2_X1 U17063 ( .A1(n15530), .A2(n10147), .ZN(n15535) );
  AOI22_X1 U17064 ( .A1(n15546), .A2(n15533), .B1(n15532), .B2(n15531), .ZN(
        n15534) );
  OAI211_X1 U17065 ( .C1(n15536), .C2(n15551), .A(n15535), .B(n15534), .ZN(
        n15566) );
  AOI211_X1 U17066 ( .C1(n15538), .C2(n15568), .A(n15537), .B(n15566), .ZN(
        n15539) );
  AOI22_X1 U17067 ( .A1(n15561), .A2(n9573), .B1(n15539), .B2(n15559), .ZN(
        P3_U3231) );
  NOR2_X1 U17068 ( .A1(n15541), .A2(n15540), .ZN(n15564) );
  XNOR2_X1 U17069 ( .A(n12391), .B(n15542), .ZN(n15562) );
  AOI22_X1 U17070 ( .A1(n15546), .A2(n15545), .B1(n15544), .B2(n15543), .ZN(
        n15550) );
  XNOR2_X1 U17071 ( .A(n12391), .B(n15547), .ZN(n15548) );
  NAND2_X1 U17072 ( .A1(n15548), .A2(n10147), .ZN(n15549) );
  OAI211_X1 U17073 ( .C1(n15562), .C2(n15551), .A(n15550), .B(n15549), .ZN(
        n15563) );
  AOI21_X1 U17074 ( .B1(n15564), .B2(n15552), .A(n15563), .ZN(n15560) );
  OAI22_X1 U17075 ( .A1(n15555), .A2(n15562), .B1(n15554), .B2(n15553), .ZN(
        n15556) );
  INV_X1 U17076 ( .A(n15556), .ZN(n15557) );
  OAI221_X1 U17077 ( .B1(n15561), .B2(n15560), .C1(n15559), .C2(n15558), .A(
        n15557), .ZN(P3_U3232) );
  INV_X1 U17078 ( .A(n15562), .ZN(n15565) );
  AOI211_X1 U17079 ( .C1(n15596), .C2(n15565), .A(n15564), .B(n15563), .ZN(
        n15601) );
  AOI22_X1 U17080 ( .A1(n15600), .A2(n15601), .B1(n8930), .B2(n15598), .ZN(
        P3_U3393) );
  AOI211_X1 U17081 ( .C1(n15568), .C2(n15596), .A(n15567), .B(n15566), .ZN(
        n15602) );
  AOI22_X1 U17082 ( .A1(n15600), .A2(n15602), .B1(n8956), .B2(n15598), .ZN(
        P3_U3396) );
  INV_X1 U17083 ( .A(n15569), .ZN(n15570) );
  AOI211_X1 U17084 ( .C1(n15572), .C2(n15596), .A(n15571), .B(n15570), .ZN(
        n15603) );
  AOI22_X1 U17085 ( .A1(n15600), .A2(n15603), .B1(n11995), .B2(n15598), .ZN(
        P3_U3399) );
  INV_X1 U17086 ( .A(n15573), .ZN(n15575) );
  AOI211_X1 U17087 ( .C1(n15576), .C2(n15596), .A(n15575), .B(n15574), .ZN(
        n15604) );
  AOI22_X1 U17088 ( .A1(n15600), .A2(n15604), .B1(n8980), .B2(n15598), .ZN(
        P3_U3402) );
  INV_X1 U17089 ( .A(n15577), .ZN(n15581) );
  INV_X1 U17090 ( .A(n15578), .ZN(n15579) );
  AOI211_X1 U17091 ( .C1(n15581), .C2(n15596), .A(n15580), .B(n15579), .ZN(
        n15605) );
  AOI22_X1 U17092 ( .A1(n15600), .A2(n15605), .B1(n8998), .B2(n15598), .ZN(
        P3_U3405) );
  INV_X1 U17093 ( .A(n15582), .ZN(n15584) );
  AOI211_X1 U17094 ( .C1(n15596), .C2(n15585), .A(n15584), .B(n15583), .ZN(
        n15606) );
  AOI22_X1 U17095 ( .A1(n15600), .A2(n15606), .B1(n9016), .B2(n15598), .ZN(
        P3_U3408) );
  INV_X1 U17096 ( .A(n15586), .ZN(n15588) );
  AOI211_X1 U17097 ( .C1(n15589), .C2(n15596), .A(n15588), .B(n15587), .ZN(
        n15607) );
  AOI22_X1 U17098 ( .A1(n15600), .A2(n15607), .B1(n9033), .B2(n15598), .ZN(
        P3_U3411) );
  INV_X1 U17099 ( .A(n15590), .ZN(n15592) );
  AOI211_X1 U17100 ( .C1(n15596), .C2(n15593), .A(n15592), .B(n15591), .ZN(
        n15608) );
  AOI22_X1 U17101 ( .A1(n15600), .A2(n15608), .B1(n9062), .B2(n15598), .ZN(
        P3_U3414) );
  AOI211_X1 U17102 ( .C1(n15597), .C2(n15596), .A(n15595), .B(n15594), .ZN(
        n15611) );
  INV_X1 U17103 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15599) );
  AOI22_X1 U17104 ( .A1(n15600), .A2(n15611), .B1(n15599), .B2(n15598), .ZN(
        P3_U3417) );
  AOI22_X1 U17105 ( .A1(n15612), .A2(n15601), .B1(n10627), .B2(n15609), .ZN(
        P3_U3460) );
  AOI22_X1 U17106 ( .A1(n15612), .A2(n15602), .B1(n9572), .B2(n15609), .ZN(
        P3_U3461) );
  AOI22_X1 U17107 ( .A1(n15612), .A2(n15603), .B1(n10450), .B2(n15609), .ZN(
        P3_U3462) );
  AOI22_X1 U17108 ( .A1(n15612), .A2(n15604), .B1(n8978), .B2(n15609), .ZN(
        P3_U3463) );
  AOI22_X1 U17109 ( .A1(n15612), .A2(n15605), .B1(n9584), .B2(n15609), .ZN(
        P3_U3464) );
  AOI22_X1 U17110 ( .A1(n15612), .A2(n15606), .B1(n9012), .B2(n15609), .ZN(
        P3_U3465) );
  AOI22_X1 U17111 ( .A1(n15612), .A2(n15607), .B1(n9030), .B2(n15609), .ZN(
        P3_U3466) );
  AOI22_X1 U17112 ( .A1(n15612), .A2(n15608), .B1(n9059), .B2(n15609), .ZN(
        P3_U3467) );
  AOI22_X1 U17113 ( .A1(n15612), .A2(n15611), .B1(n15610), .B2(n15609), .ZN(
        P3_U3468) );
  XNOR2_X1 U17114 ( .A(n15614), .B(n15613), .ZN(n15615) );
  XNOR2_X1 U17115 ( .A(n15615), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U17116 ( .A(n15617), .B(n15616), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7177 ( .A(n14962), .Z(n6432) );
  BUF_X1 U7180 ( .A(n9075), .Z(n9814) );
  NAND2_X2 U7184 ( .A1(n7856), .A2(n10193), .ZN(n8262) );
  XNOR2_X1 U7236 ( .A(n9415), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12394) );
  NAND2_X2 U7459 ( .A1(n7809), .A2(n10433), .ZN(n7856) );
  CLKBUF_X2 U9683 ( .A(n9424), .Z(n13714) );
endmodule

