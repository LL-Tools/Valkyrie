

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150;

  NAND2_X1 U5152 ( .A1(n6197), .A2(n6196), .ZN(n6225) );
  CLKBUF_X2 U5153 ( .A(n6548), .Z(n6639) );
  CLKBUF_X2 U5154 ( .A(n6125), .Z(n5102) );
  CLKBUF_X2 U5155 ( .A(n5100), .Z(n6121) );
  INV_X2 U5156 ( .A(n8670), .ZN(n8679) );
  CLKBUF_X2 U5158 ( .A(n7223), .Z(n8540) );
  CLKBUF_X3 U5159 ( .A(n5126), .Z(n8643) );
  INV_X1 U5160 ( .A(n5845), .ZN(n5090) );
  NAND4_X1 U5161 ( .A1(n7005), .A2(n7004), .A3(n7003), .A4(n7002), .ZN(n9074)
         );
  NAND2_X1 U5162 ( .A1(n5805), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U5163 ( .A1(n5802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U5164 ( .A1(n5104), .A2(n5848), .ZN(n5913) );
  NAND2_X1 U5166 ( .A1(n7406), .A2(n10930), .ZN(n8462) );
  CLKBUF_X2 U5168 ( .A(n5954), .Z(n6519) );
  BUF_X1 U5169 ( .A(n5785), .Z(n5786) );
  NAND2_X1 U5170 ( .A1(n5793), .A2(n10735), .ZN(n5802) );
  INV_X1 U5171 ( .A(n5876), .ZN(n10334) );
  NAND2_X1 U5172 ( .A1(n5796), .A2(n5802), .ZN(n7908) );
  INV_X1 U5173 ( .A(n5867), .ZN(n5091) );
  INV_X1 U5174 ( .A(n7226), .ZN(n5106) );
  AND2_X2 U5175 ( .A1(n5768), .A2(n5831), .ZN(n5931) );
  AOI211_X2 U5176 ( .C1(n8565), .C2(n8343), .A(n8342), .B(n8341), .ZN(n8344)
         );
  OAI21_X2 U5177 ( .B1(n6324), .B2(n6323), .A(n6322), .ZN(n6349) );
  NAND2_X2 U5178 ( .A1(n9948), .A2(n9947), .ZN(n9961) );
  OAI211_X4 U5179 ( .C1(n9730), .C2(n7041), .A(n5874), .B(n5873), .ZN(n7523)
         );
  AND2_X1 U5180 ( .A1(n7301), .A2(n7302), .ZN(n5946) );
  AND4_X2 U5181 ( .A1(n6670), .A2(n6669), .A3(n6668), .A4(n6667), .ZN(n5127)
         );
  INV_X1 U5182 ( .A(n8451), .ZN(n8774) );
  NAND2_X2 U5183 ( .A1(n7346), .A2(n8449), .ZN(n8456) );
  NAND2_X2 U5184 ( .A1(n8448), .A2(n8741), .ZN(n7346) );
  NAND2_X1 U5185 ( .A1(n8198), .A2(n8760), .ZN(n8701) );
  OR2_X1 U5186 ( .A1(n5843), .A2(n5841), .ZN(n7637) );
  NAND3_X4 U5187 ( .A1(n5816), .A2(n5817), .A3(n5815), .ZN(n5857) );
  NAND4_X2 U5188 ( .A1(n5863), .A2(n5862), .A3(n5861), .A4(n5860), .ZN(n6953)
         );
  NAND2_X2 U5189 ( .A1(n6770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6772) );
  OAI211_X2 U5190 ( .C1(n6013), .C2(n6730), .A(n5989), .B(n5988), .ZN(n7783)
         );
  OAI21_X2 U5191 ( .B1(n6225), .B2(n6224), .A(n6223), .ZN(n6248) );
  OAI21_X2 U5192 ( .B1(n9199), .B2(n8725), .A(n8724), .ZN(n9184) );
  NAND2_X2 U5193 ( .A1(n9394), .A2(n8722), .ZN(n9199) );
  AND2_X1 U5194 ( .A1(n5876), .A2(n5877), .ZN(n6125) );
  NOR2_X2 U5195 ( .A1(n9966), .A2(n9965), .ZN(n9972) );
  NOR2_X2 U5196 ( .A1(n7166), .A2(n5211), .ZN(n7267) );
  AOI21_X4 U5197 ( .B1(n9271), .B2(n8711), .A(n8710), .ZN(n9275) );
  CLKBUF_X2 U5198 ( .A(n7562), .Z(n5088) );
  OAI21_X2 U5199 ( .B1(n6712), .B2(n6714), .A(n6713), .ZN(n6716) );
  NAND2_X1 U5200 ( .A1(n8820), .A2(n8819), .ZN(n8973) );
  NAND2_X1 U5201 ( .A1(n8001), .A2(n8509), .ZN(n8005) );
  INV_X2 U5202 ( .A(n8758), .ZN(n8518) );
  NAND2_X2 U5203 ( .A1(n8506), .A2(n8496), .ZN(n8751) );
  AND2_X1 U5204 ( .A1(n9851), .A2(n9660), .ZN(n9658) );
  INV_X1 U5206 ( .A(n9068), .ZN(n7737) );
  INV_X1 U5207 ( .A(n9067), .ZN(n7827) );
  NAND2_X1 U5208 ( .A1(n9844), .A2(n9650), .ZN(n10908) );
  INV_X1 U5209 ( .A(n10970), .ZN(n11011) );
  INV_X1 U5210 ( .A(n9069), .ZN(n7567) );
  INV_X1 U5211 ( .A(n9070), .ZN(n7405) );
  INV_X1 U5212 ( .A(n9071), .ZN(n7406) );
  INV_X2 U5213 ( .A(n5091), .ZN(n6638) );
  INV_X1 U5214 ( .A(n9909), .ZN(n7628) );
  NAND4_X1 U5215 ( .A1(n7230), .A2(n7229), .A3(n7228), .A4(n7227), .ZN(n9070)
         );
  INV_X1 U5216 ( .A(n7562), .ZN(n10937) );
  CLKBUF_X2 U5217 ( .A(n8110), .Z(n8689) );
  BUF_X1 U5218 ( .A(n5951), .Z(n5100) );
  NAND2_X1 U5219 ( .A1(n6787), .A2(n7036), .ZN(n9730) );
  CLKBUF_X1 U5220 ( .A(n5841), .Z(n10179) );
  INV_X2 U5221 ( .A(n7502), .ZN(n7561) );
  CLKBUF_X2 U5223 ( .A(n5827), .Z(n8684) );
  NOR2_X4 U5224 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6712) );
  NAND2_X1 U5225 ( .A1(n9619), .A2(n6532), .ZN(n9620) );
  NAND2_X1 U5226 ( .A1(n8777), .A2(n8776), .ZN(n8781) );
  NAND2_X1 U5227 ( .A1(n5646), .A2(n5170), .ZN(n9580) );
  OR2_X1 U5228 ( .A1(n9600), .A2(n9521), .ZN(n5651) );
  AND2_X1 U5229 ( .A1(n5653), .A2(n5652), .ZN(n9522) );
  INV_X1 U5230 ( .A(n9380), .ZN(n9381) );
  OR2_X1 U5231 ( .A1(n9379), .A2(n8883), .ZN(n5464) );
  AND2_X1 U5232 ( .A1(n10246), .A2(n5209), .ZN(n5671) );
  NOR2_X1 U5233 ( .A1(n10244), .A2(n5185), .ZN(n5209) );
  NAND3_X1 U5234 ( .A1(n5626), .A2(n5628), .A3(n5625), .ZN(n9564) );
  AND2_X1 U5235 ( .A1(n8983), .A2(n8837), .ZN(n8836) );
  NAND2_X1 U5236 ( .A1(n8215), .A2(n6192), .ZN(n6219) );
  NAND2_X1 U5237 ( .A1(n9732), .A2(n9731), .ZN(n10245) );
  XNOR2_X1 U5238 ( .A(n8688), .B(n8687), .ZN(n9645) );
  XNOR2_X1 U5239 ( .A(n8683), .B(n8682), .ZN(n9734) );
  NAND2_X1 U5240 ( .A1(n5700), .A2(n5703), .ZN(n10138) );
  NAND2_X1 U5241 ( .A1(n8973), .A2(n5745), .ZN(n9022) );
  OAI21_X1 U5242 ( .B1(n8250), .B2(n5298), .A(n5295), .ZN(n8967) );
  NAND2_X1 U5243 ( .A1(n8178), .A2(n8177), .ZN(n8183) );
  OR2_X1 U5244 ( .A1(n8176), .A2(n9061), .ZN(n8177) );
  AND2_X1 U5245 ( .A1(n8144), .A2(n9911), .ZN(n9922) );
  OAI21_X1 U5246 ( .B1(n11071), .B2(n11070), .A(n11069), .ZN(n11074) );
  OAI21_X1 U5247 ( .B1(n8041), .B2(n8040), .A(n8039), .ZN(n8042) );
  NOR2_X1 U5248 ( .A1(n8237), .A2(n8238), .ZN(n8240) );
  NOR2_X1 U5249 ( .A1(n8052), .A2(n11090), .ZN(n8237) );
  NAND2_X1 U5250 ( .A1(n7647), .A2(n7646), .ZN(n7763) );
  OAI21_X1 U5251 ( .B1(n5309), .B2(n5308), .A(n5306), .ZN(n7647) );
  NAND2_X1 U5252 ( .A1(n7729), .A2(n5445), .ZN(n7924) );
  OR2_X1 U5253 ( .A1(n7584), .A2(n5305), .ZN(n5306) );
  INV_X1 U5254 ( .A(n6083), .ZN(n5089) );
  NOR2_X1 U5255 ( .A1(n7854), .A2(n7853), .ZN(n7857) );
  OAI21_X1 U5256 ( .B1(n5750), .B2(n5752), .A(n5748), .ZN(n7584) );
  NAND2_X1 U5257 ( .A1(n8119), .A2(n8118), .ZN(n11107) );
  NAND2_X1 U5258 ( .A1(n5749), .A2(n5754), .ZN(n5748) );
  NAND2_X1 U5259 ( .A1(n6069), .A2(n6068), .ZN(n7712) );
  OAI21_X1 U5260 ( .B1(n7427), .B2(n7417), .A(n7416), .ZN(n7563) );
  AND2_X1 U5261 ( .A1(n8499), .A2(n8484), .ZN(n8746) );
  NOR2_X1 U5262 ( .A1(n5610), .A2(n7498), .ZN(n7669) );
  INV_X2 U5263 ( .A(n11111), .ZN(n9352) );
  NAND2_X1 U5264 ( .A1(n5501), .A2(n5500), .ZN(n5499) );
  AOI21_X1 U5265 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7561), .A(n7494), .ZN(
        n7495) );
  OAI21_X1 U5266 ( .B1(n7167), .B2(n5617), .A(n5616), .ZN(n7494) );
  INV_X1 U5267 ( .A(n6636), .ZN(n5992) );
  NAND4_X2 U5268 ( .A1(n7198), .A2(n7197), .A3(n7196), .A4(n7195), .ZN(n9071)
         );
  NOR2_X2 U5269 ( .A1(n9193), .A2(n8670), .ZN(n7120) );
  AND4_X1 U5270 ( .A1(n7149), .A2(n7148), .A3(n7147), .A4(n7146), .ZN(n7413)
         );
  NAND4_X1 U5271 ( .A1(n5900), .A2(n5899), .A3(n5898), .A4(n5897), .ZN(n9909)
         );
  OAI211_X1 U5272 ( .C1(n8399), .C2(n7234), .A(n7233), .B(n7232), .ZN(n7562)
         );
  INV_X1 U5273 ( .A(n7523), .ZN(n10880) );
  XNOR2_X1 U5274 ( .A(n7267), .B(n7377), .ZN(n7167) );
  BUF_X2 U5275 ( .A(n6143), .Z(n9644) );
  OR2_X1 U5276 ( .A1(n5954), .A2(n5778), .ZN(n5784) );
  NAND2_X1 U5277 ( .A1(n5359), .A2(n5358), .ZN(n6947) );
  NAND2_X1 U5278 ( .A1(n5614), .A2(n5613), .ZN(n7166) );
  INV_X2 U5279 ( .A(n7037), .ZN(n8578) );
  NAND2_X1 U5280 ( .A1(n7932), .A2(n8579), .ZN(n8785) );
  NAND2_X1 U5281 ( .A1(n7037), .A2(n8684), .ZN(n8399) );
  INV_X1 U5282 ( .A(n6773), .ZN(n9514) );
  AND2_X2 U5283 ( .A1(n6787), .A2(n8684), .ZN(n5979) );
  NAND2_X1 U5284 ( .A1(n5841), .A2(n7908), .ZN(n6948) );
  NAND2_X1 U5285 ( .A1(n9835), .A2(n7908), .ZN(n5843) );
  NAND2_X2 U5286 ( .A1(n5780), .A2(n10334), .ZN(n5954) );
  NAND2_X1 U5287 ( .A1(n5777), .A2(n5776), .ZN(n5780) );
  XNOR2_X1 U5288 ( .A(n5814), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6574) );
  XNOR2_X1 U5289 ( .A(n5792), .B(n5791), .ZN(n5841) );
  AND2_X1 U5290 ( .A1(n5813), .A2(n5811), .ZN(n5797) );
  MUX2_X1 U5291 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6704), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n6708) );
  XNOR2_X1 U5292 ( .A(n5813), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9835) );
  XNOR2_X1 U5293 ( .A(n6702), .B(n6705), .ZN(n6834) );
  OR2_X1 U5294 ( .A1(n6602), .A2(n10748), .ZN(n6797) );
  OR2_X1 U5295 ( .A1(n5790), .A2(n5789), .ZN(n5792) );
  NOR2_X1 U5296 ( .A1(n6899), .A2(n7235), .ZN(n7072) );
  MUX2_X1 U5297 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5775), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5777) );
  NOR2_X1 U5298 ( .A1(n6277), .A2(n5788), .ZN(n5790) );
  INV_X1 U5299 ( .A(n5802), .ZN(n5800) );
  OAI21_X1 U5300 ( .B1(n7491), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6992) );
  XNOR2_X1 U5301 ( .A(n5982), .B(n5965), .ZN(n5980) );
  NOR2_X1 U5302 ( .A1(n6731), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6739) );
  OR2_X1 U5303 ( .A1(n6721), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6731) );
  NAND2_X2 U5304 ( .A1(n8684), .A2(P2_U3151), .ZN(n9518) );
  AND2_X1 U5305 ( .A1(n5127), .A2(n5725), .ZN(n5210) );
  INV_X1 U5306 ( .A(n5725), .ZN(n6721) );
  AND2_X1 U5307 ( .A1(n5552), .A2(n6707), .ZN(n5551) );
  INV_X1 U5308 ( .A(n5827), .ZN(n5824) );
  OR2_X1 U5309 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(n5787), .ZN(n5788) );
  AND2_X1 U5310 ( .A1(n5759), .A2(n6684), .ZN(n5552) );
  AND2_X1 U5311 ( .A1(n5178), .A2(n6686), .ZN(n5759) );
  CLKBUF_X1 U5312 ( .A(n5931), .Z(n5934) );
  NAND3_X1 U5313 ( .A1(n6662), .A2(n5589), .A3(n5590), .ZN(n6724) );
  AND3_X1 U5314 ( .A1(n5624), .A2(n5623), .A3(n5622), .ZN(n6144) );
  AND2_X1 U5315 ( .A1(n10736), .A2(n5366), .ZN(n5808) );
  AND3_X1 U5316 ( .A1(n6738), .A2(n6666), .A3(n6665), .ZN(n6670) );
  INV_X1 U5317 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6662) );
  INV_X4 U5318 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5319 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10730) );
  INV_X1 U5320 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10729) );
  INV_X1 U5321 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5590) );
  INV_X1 U5322 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5791) );
  NOR2_X1 U5323 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5769) );
  INV_X1 U5324 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6684) );
  INV_X1 U5325 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6679) );
  INV_X1 U5326 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10743) );
  NOR2_X1 U5327 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5624) );
  NOR2_X1 U5328 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5623) );
  NOR2_X1 U5329 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5622) );
  INV_X1 U5330 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10737) );
  INV_X1 U5331 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7490) );
  NOR2_X2 U5332 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5831) );
  NOR2_X1 U5333 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5768) );
  INV_X1 U5334 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5933) );
  INV_X1 U5335 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5228) );
  INV_X4 U5336 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U5337 ( .A1(n5093), .A2(n5946), .ZN(n5092) );
  CLKBUF_X1 U5338 ( .A(n7211), .Z(n5093) );
  CLKBUF_X1 U5339 ( .A(n7793), .Z(n5094) );
  NAND2_X1 U5340 ( .A1(n9536), .A2(n5097), .ZN(n5095) );
  AND2_X1 U5341 ( .A1(n5095), .A2(n5096), .ZN(n6106) );
  OR2_X1 U5342 ( .A1(n5089), .A2(n5145), .ZN(n5096) );
  AND2_X1 U5343 ( .A1(n6054), .A2(n6083), .ZN(n5097) );
  NAND2_X1 U5344 ( .A1(n7210), .A2(n7209), .ZN(n7211) );
  XNOR2_X2 U5345 ( .A(n5801), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6573) );
  NAND2_X2 U5346 ( .A1(n9514), .A2(n9519), .ZN(n7044) );
  INV_X1 U5347 ( .A(n7239), .ZN(n5098) );
  INV_X4 U5348 ( .A(n5098), .ZN(n5099) );
  OAI21_X1 U5349 ( .B1(n7342), .B2(n7033), .A(n7034), .ZN(n7239) );
  AND2_X2 U5350 ( .A1(n5857), .A2(n5837), .ZN(n5867) );
  AND2_X1 U5351 ( .A1(n6410), .A2(n5183), .ZN(n9600) );
  NAND2_X2 U5352 ( .A1(n7568), .A2(n8746), .ZN(n7729) );
  AND3_X1 U5353 ( .A1(n5150), .A2(n5785), .A3(n5721), .ZN(n5818) );
  NAND4_X2 U5354 ( .A1(n5784), .A2(n5783), .A3(n5782), .A4(n5781), .ZN(n5839)
         );
  OR2_X2 U5355 ( .A1(n9325), .A2(n9324), .ZN(n9427) );
  OR4_X4 U5356 ( .A1(n6658), .A2(n6642), .A3(n6643), .A4(n9616), .ZN(n6660) );
  AOI22_X2 U5357 ( .A1(n8261), .A2(n8260), .B1(n9899), .B2(n8259), .ZN(n10015)
         );
  NAND2_X2 U5358 ( .A1(n8005), .A2(n8755), .ZN(n8134) );
  AOI21_X2 U5359 ( .B1(n10961), .B2(n10966), .A(n7635), .ZN(n7781) );
  NAND2_X2 U5360 ( .A1(n7633), .A2(n9846), .ZN(n10966) );
  NAND2_X1 U5361 ( .A1(n7632), .A2(n7631), .ZN(n10961) );
  NAND2_X2 U5362 ( .A1(n8134), .A2(n8512), .ZN(n8135) );
  OAI21_X2 U5363 ( .B1(n8135), .B2(n5136), .A(n5431), .ZN(n8198) );
  NAND2_X1 U5364 ( .A1(n8720), .A2(n8719), .ZN(n9229) );
  NAND2_X2 U5365 ( .A1(n9427), .A2(n5475), .ZN(n9271) );
  OR2_X1 U5366 ( .A1(n5954), .A2(n5859), .ZN(n5863) );
  INV_X4 U5367 ( .A(n7248), .ZN(n8597) );
  NAND2_X2 U5368 ( .A1(n9557), .A2(n9558), .ZN(n9619) );
  NAND2_X1 U5369 ( .A1(n7413), .A2(n7347), .ZN(n8461) );
  OR2_X1 U5370 ( .A1(n7044), .A2(n6775), .ZN(n6777) );
  AND2_X2 U5371 ( .A1(n6774), .A2(n9514), .ZN(n5126) );
  OAI222_X1 U5372 ( .A1(n10340), .A2(n8105), .B1(P1_U3086), .B2(n6573), .C1(
        n10687), .C2(n10337), .ZN(P1_U3330) );
  NAND2_X1 U5373 ( .A1(n6769), .A2(n6770), .ZN(n9519) );
  XNOR2_X1 U5374 ( .A(n5849), .B(n5992), .ZN(n5850) );
  NOR2_X1 U5375 ( .A1(n5876), .A2(n5780), .ZN(n5951) );
  OAI21_X1 U5376 ( .B1(n9379), .B2(n10954), .A(n9378), .ZN(n9380) );
  XNOR2_X1 U5377 ( .A(n6722), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7231) );
  OAI211_X1 U5378 ( .C1(n6948), .C2(n9893), .A(n7637), .B(n5857), .ZN(n5104)
         );
  OAI211_X1 U5379 ( .C1(n6948), .C2(n9893), .A(n7637), .B(n5857), .ZN(n5105)
         );
  OAI211_X1 U5380 ( .C1(n6948), .C2(n9893), .A(n7637), .B(n5857), .ZN(n5845)
         );
  INV_X1 U5381 ( .A(n5106), .ZN(n5107) );
  XNOR2_X2 U5382 ( .A(n6772), .B(n6771), .ZN(n6773) );
  NAND2_X1 U5383 ( .A1(n8187), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7228) );
  XNOR2_X2 U5384 ( .A(n5807), .B(n5806), .ZN(n6576) );
  AND2_X1 U5385 ( .A1(n6787), .A2(n8684), .ZN(n5108) );
  AND2_X1 U5386 ( .A1(n6787), .A2(n8684), .ZN(n5109) );
  INV_X1 U5387 ( .A(n5091), .ZN(n6528) );
  OAI222_X1 U5388 ( .A1(n9519), .A2(P2_U3151), .B1(n9518), .B2(n10336), .C1(
        n9517), .C2(n9516), .ZN(P2_U3266) );
  INV_X1 U5389 ( .A(n9513), .ZN(n9516) );
  NOR2_X1 U5390 ( .A1(n5268), .A2(n5267), .ZN(n5266) );
  NOR2_X1 U5391 ( .A1(n5258), .A2(n9782), .ZN(n5268) );
  NAND2_X1 U5392 ( .A1(n6250), .A2(n6249), .ZN(n6271) );
  INV_X1 U5393 ( .A(SI_16_), .ZN(n6249) );
  NAND2_X1 U5394 ( .A1(n6199), .A2(n6198), .ZN(n6223) );
  INV_X1 U5395 ( .A(SI_14_), .ZN(n6198) );
  NAND2_X1 U5396 ( .A1(n8401), .A2(n5437), .ZN(n8737) );
  AND2_X1 U5397 ( .A1(n5438), .A2(n8400), .ZN(n5437) );
  OR2_X1 U5398 ( .A1(n8934), .A2(n9290), .ZN(n8708) );
  NAND2_X1 U5399 ( .A1(n6484), .A2(n6483), .ZN(n6486) );
  NAND2_X1 U5400 ( .A1(n6457), .A2(n6456), .ZN(n6484) );
  NOR2_X1 U5401 ( .A1(n6140), .A2(n5462), .ZN(n5461) );
  INV_X1 U5402 ( .A(n6110), .ZN(n5462) );
  OR2_X1 U5403 ( .A1(n6061), .A2(n5247), .ZN(n5246) );
  NAND2_X1 U5404 ( .A1(n5765), .A2(n5248), .ZN(n5247) );
  INV_X1 U5405 ( .A(n6060), .ZN(n5248) );
  NAND2_X1 U5406 ( .A1(n10075), .A2(n9747), .ZN(n5276) );
  AOI21_X1 U5407 ( .B1(n5281), .B2(n5279), .A(n9742), .ZN(n5278) );
  INV_X1 U5408 ( .A(n5273), .ZN(n5272) );
  OR2_X1 U5409 ( .A1(n10245), .A2(n9733), .ZN(n9750) );
  OR2_X1 U5410 ( .A1(n6414), .A2(n6413), .ZN(n6417) );
  NAND2_X1 U5411 ( .A1(n5195), .A2(n6372), .ZN(n5450) );
  NAND2_X1 U5412 ( .A1(n6348), .A2(n6347), .ZN(n5452) );
  OAI21_X1 U5413 ( .B1(n5731), .B2(n5730), .A(n8072), .ZN(n5729) );
  NAND2_X1 U5414 ( .A1(n8945), .A2(n5757), .ZN(n5756) );
  INV_X1 U5415 ( .A(n8828), .ZN(n5757) );
  INV_X1 U5416 ( .A(n8801), .ZN(n5302) );
  INV_X1 U5417 ( .A(n9519), .ZN(n6774) );
  NAND2_X1 U5418 ( .A1(n5491), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5490) );
  OAI21_X1 U5419 ( .B1(n5549), .B2(n5547), .A(n5188), .ZN(n5546) );
  INV_X1 U5420 ( .A(n8878), .ZN(n5547) );
  OR2_X1 U5421 ( .A1(n8896), .A2(n9209), .ZN(n8723) );
  NAND2_X1 U5422 ( .A1(n8896), .A2(n9209), .ZN(n8724) );
  OR2_X1 U5423 ( .A1(n9232), .A2(n9248), .ZN(n8872) );
  AND2_X1 U5424 ( .A1(n9232), .A2(n9248), .ZN(n8870) );
  INV_X1 U5425 ( .A(n9293), .ZN(n5536) );
  NAND2_X1 U5426 ( .A1(n5522), .A2(n9061), .ZN(n5518) );
  INV_X1 U5427 ( .A(n8183), .ZN(n5531) );
  NAND4_X1 U5428 ( .A1(n5725), .A2(n5114), .A3(n5127), .A4(n6684), .ZN(n5321)
         );
  AOI21_X1 U5429 ( .B1(n5266), .B2(n5118), .A(n9884), .ZN(n5264) );
  NOR2_X1 U5430 ( .A1(n5256), .A2(n5255), .ZN(n5254) );
  INV_X1 U5431 ( .A(n9782), .ZN(n5257) );
  INV_X1 U5432 ( .A(n5263), .ZN(n5260) );
  OR2_X1 U5433 ( .A1(n10248), .A2(n10029), .ZN(n9749) );
  OR2_X1 U5434 ( .A1(n10254), .A2(n10080), .ZN(n10047) );
  OR2_X1 U5435 ( .A1(n10259), .A2(n10096), .ZN(n9751) );
  NOR2_X1 U5436 ( .A1(n10114), .A2(n9791), .ZN(n5678) );
  OR2_X1 U5437 ( .A1(n10277), .A2(n10162), .ZN(n10001) );
  NAND2_X1 U5438 ( .A1(n10001), .A2(n9717), .ZN(n10021) );
  OR2_X1 U5439 ( .A1(n10299), .A2(n9709), .ZN(n9794) );
  OR2_X1 U5440 ( .A1(n10100), .A2(n10259), .ZN(n10065) );
  NAND2_X1 U5441 ( .A1(n8398), .A2(n8391), .ZN(n8683) );
  OR2_X1 U5442 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  NAND2_X1 U5443 ( .A1(n5467), .A2(n5465), .ZN(n6627) );
  AOI21_X1 U5444 ( .B1(n5469), .B2(n5471), .A(n5466), .ZN(n5465) );
  INV_X1 U5445 ( .A(n6543), .ZN(n5466) );
  AOI21_X1 U5446 ( .B1(n6248), .B2(n5425), .A(n5422), .ZN(n5421) );
  NAND2_X1 U5447 ( .A1(n5423), .A2(n6299), .ZN(n5422) );
  NAND2_X1 U5448 ( .A1(n5425), .A2(n5427), .ZN(n5423) );
  AND2_X1 U5449 ( .A1(n6299), .A2(n6276), .ZN(n6297) );
  NAND2_X1 U5450 ( .A1(n6271), .A2(n6252), .ZN(n6272) );
  AOI21_X1 U5451 ( .B1(n5455), .B2(n5457), .A(n6193), .ZN(n5454) );
  NAND2_X1 U5452 ( .A1(n6139), .A2(n6116), .ZN(n6140) );
  AOI21_X1 U5453 ( .B1(n5765), .B2(n5251), .A(n5250), .ZN(n5249) );
  INV_X1 U5454 ( .A(n6085), .ZN(n5250) );
  INV_X1 U5455 ( .A(n6059), .ZN(n5251) );
  NAND2_X1 U5456 ( .A1(n6041), .A2(n6040), .ZN(n6061) );
  INV_X1 U5457 ( .A(n6036), .ZN(n6037) );
  INV_X1 U5458 ( .A(n5312), .ZN(n5308) );
  AOI21_X1 U5459 ( .B1(n8674), .B2(n8673), .A(n8672), .ZN(n8675) );
  OAI21_X1 U5460 ( .B1(n8781), .B2(n5215), .A(n5214), .ZN(n5213) );
  AOI21_X1 U5461 ( .B1(n8786), .B2(n8779), .A(n8792), .ZN(n5214) );
  NAND2_X1 U5462 ( .A1(n5217), .A2(n5216), .ZN(n5215) );
  INV_X1 U5463 ( .A(n8778), .ZN(n5216) );
  INV_X1 U5464 ( .A(n7281), .ZN(n5500) );
  AOI21_X1 U5465 ( .B1(n8293), .B2(n8305), .A(n9095), .ZN(n5502) );
  NAND2_X1 U5466 ( .A1(n5497), .A2(n5496), .ZN(n5495) );
  INV_X1 U5467 ( .A(n9140), .ZN(n5496) );
  NAND2_X1 U5468 ( .A1(n5486), .A2(n8300), .ZN(n5484) );
  NOR2_X1 U5469 ( .A1(n9434), .A2(n9160), .ZN(n9159) );
  AND2_X1 U5470 ( .A1(n8708), .A2(n8707), .ZN(n5475) );
  OR2_X1 U5471 ( .A1(n9428), .A2(n8940), .ZN(n8707) );
  NAND2_X1 U5472 ( .A1(n8401), .A2(n8400), .ZN(n5442) );
  AND2_X2 U5473 ( .A1(n5210), .A2(n5114), .ZN(n6685) );
  NOR2_X1 U5474 ( .A1(n6319), .A2(n9611), .ZN(n5641) );
  AND2_X1 U5475 ( .A1(n9749), .A2(n10007), .ZN(n10049) );
  NOR2_X1 U5476 ( .A1(n9764), .A2(n5335), .ZN(n5334) );
  INV_X1 U5477 ( .A(n9793), .ZN(n5335) );
  INV_X1 U5478 ( .A(n9999), .ZN(n5332) );
  NOR2_X1 U5479 ( .A1(n10176), .A2(n5709), .ZN(n5708) );
  NOR2_X1 U5480 ( .A1(n5111), .A2(n10018), .ZN(n5709) );
  NAND2_X1 U5481 ( .A1(n5662), .A2(n10191), .ZN(n10194) );
  NAND2_X1 U5482 ( .A1(n5327), .A2(n5663), .ZN(n5662) );
  AOI21_X1 U5483 ( .B1(n5666), .B2(n5664), .A(n9762), .ZN(n5663) );
  OR2_X1 U5484 ( .A1(n10299), .A2(n10223), .ZN(n5212) );
  AND2_X1 U5485 ( .A1(n7898), .A2(n9903), .ZN(n5207) );
  INV_X1 U5486 ( .A(n7897), .ZN(n5208) );
  OR2_X1 U5487 ( .A1(n9543), .A2(n9906), .ZN(n5694) );
  INV_X2 U5488 ( .A(n6787), .ZN(n6329) );
  XNOR2_X1 U5489 ( .A(n6538), .B(n6537), .ZN(n8426) );
  NAND2_X1 U5490 ( .A1(n5468), .A2(n6504), .ZN(n6538) );
  XNOR2_X1 U5491 ( .A(n6484), .B(n6483), .ZN(n8636) );
  XNOR2_X1 U5493 ( .A(n8833), .B(n8834), .ZN(n8919) );
  NAND2_X1 U5494 ( .A1(n10391), .A2(SI_26_), .ZN(n10393) );
  NAND2_X1 U5495 ( .A1(n10597), .A2(keyinput_6), .ZN(n10392) );
  NAND2_X1 U5496 ( .A1(n5388), .A2(n5387), .ZN(n5386) );
  INV_X1 U5497 ( .A(n10624), .ZN(n5387) );
  NAND2_X1 U5498 ( .A1(n10615), .A2(n5389), .ZN(n5388) );
  AND2_X1 U5499 ( .A1(n10622), .A2(n10623), .ZN(n5385) );
  AOI21_X1 U5500 ( .B1(n5582), .B2(n5581), .A(n5578), .ZN(n10463) );
  NAND2_X1 U5501 ( .A1(n5580), .A2(n5579), .ZN(n5578) );
  AOI22_X1 U5502 ( .A1(n7023), .A2(n10452), .B1(keyinput_50), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n5581) );
  OAI21_X1 U5503 ( .B1(n10449), .B2(n5586), .A(n5583), .ZN(n5582) );
  OAI21_X1 U5504 ( .B1(n5113), .B2(n5242), .A(n5119), .ZN(n5239) );
  INV_X1 U5505 ( .A(n9668), .ZN(n5242) );
  OR2_X1 U5506 ( .A1(n9682), .A2(n9747), .ZN(n5238) );
  OAI21_X1 U5507 ( .B1(n9856), .B2(n5237), .A(n9747), .ZN(n5236) );
  AND2_X1 U5508 ( .A1(n9681), .A2(n9853), .ZN(n5237) );
  NAND2_X1 U5509 ( .A1(n9857), .A2(n9747), .ZN(n5244) );
  OAI21_X1 U5510 ( .B1(n10479), .B2(n5577), .A(n5576), .ZN(n5575) );
  AND2_X1 U5511 ( .A1(n10685), .A2(keyinput_70), .ZN(n5577) );
  AOI22_X1 U5512 ( .A1(n10687), .A2(n10480), .B1(keyinput_71), .B2(
        P2_DATAO_REG_25__SCAN_IN), .ZN(n5576) );
  AOI21_X1 U5513 ( .B1(n10684), .B2(n5381), .A(n5380), .ZN(n5379) );
  NAND2_X1 U5514 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n5382), .ZN(n5381) );
  OAI22_X1 U5515 ( .A1(n10687), .A2(n10686), .B1(P2_DATAO_REG_25__SCAN_IN), 
        .B2(keyinput_199), .ZN(n5380) );
  NAND2_X1 U5516 ( .A1(n5404), .A2(n5401), .ZN(n5400) );
  AND2_X1 U5517 ( .A1(n5403), .A2(n5402), .ZN(n5401) );
  OR2_X1 U5518 ( .A1(n10693), .A2(n5405), .ZN(n5404) );
  NAND2_X1 U5519 ( .A1(n10696), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n5402) );
  NOR2_X1 U5520 ( .A1(n5117), .A2(n5160), .ZN(n5289) );
  INV_X1 U5521 ( .A(n5287), .ZN(n5286) );
  OAI21_X1 U5522 ( .B1(n5293), .B2(n9742), .A(n5288), .ZN(n5287) );
  AND2_X1 U5523 ( .A1(n9761), .A2(n9794), .ZN(n5293) );
  NOR2_X1 U5524 ( .A1(n9877), .A2(n5189), .ZN(n5288) );
  AOI21_X1 U5525 ( .B1(n5559), .B2(n10512), .A(n5203), .ZN(n10515) );
  OAI21_X1 U5526 ( .B1(n10504), .B2(n5562), .A(n5560), .ZN(n5559) );
  OAI21_X1 U5527 ( .B1(n5554), .B2(n5202), .A(n5553), .ZN(n10536) );
  NOR2_X1 U5528 ( .A1(n10531), .A2(n10532), .ZN(n5553) );
  AOI21_X1 U5529 ( .B1(n5558), .B2(n5556), .A(n5555), .ZN(n5554) );
  NAND2_X1 U5530 ( .A1(n10718), .A2(n10717), .ZN(n5375) );
  INV_X1 U5531 ( .A(n5276), .ZN(n5275) );
  INV_X1 U5532 ( .A(n5278), .ZN(n5274) );
  AOI21_X1 U5533 ( .B1(n5277), .B2(n5276), .A(n5154), .ZN(n5273) );
  NAND2_X1 U5534 ( .A1(n5162), .A2(n10075), .ZN(n5277) );
  INV_X1 U5535 ( .A(n5281), .ZN(n5280) );
  INV_X1 U5536 ( .A(n9725), .ZN(n5283) );
  NOR2_X1 U5537 ( .A1(n8599), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8598) );
  INV_X1 U5538 ( .A(n5980), .ZN(n5231) );
  INV_X1 U5539 ( .A(n5983), .ZN(n5233) );
  INV_X1 U5540 ( .A(n8995), .ZN(n5758) );
  INV_X1 U5541 ( .A(n8823), .ZN(n5320) );
  OAI21_X1 U5542 ( .B1(n8677), .B2(n9385), .A(n8415), .ZN(n8674) );
  NOR2_X1 U5543 ( .A1(n7669), .A2(n5612), .ZN(n7851) );
  AND2_X1 U5544 ( .A1(n7670), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5612) );
  AOI21_X1 U5545 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n8054), .A(n8053), .ZN(
        n8222) );
  AND2_X1 U5546 ( .A1(n5495), .A2(n5494), .ZN(n8298) );
  NAND2_X1 U5547 ( .A1(n8335), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U5548 ( .A1(n5168), .A2(n5125), .ZN(n5549) );
  NAND2_X1 U5549 ( .A1(n5138), .A2(n8875), .ZN(n5550) );
  OR2_X1 U5550 ( .A1(n9392), .A2(n9059), .ZN(n8875) );
  OR2_X1 U5551 ( .A1(n9392), .A2(n9224), .ZN(n8722) );
  OR2_X1 U5552 ( .A1(n9220), .A2(n9237), .ZN(n8655) );
  OR2_X1 U5553 ( .A1(n9253), .A2(n9238), .ZN(n8717) );
  INV_X1 U5554 ( .A(n8136), .ZN(n5434) );
  AOI21_X1 U5555 ( .B1(n8758), .B2(n5520), .A(n5152), .ZN(n5519) );
  INV_X1 U5556 ( .A(n8114), .ZN(n5520) );
  INV_X1 U5557 ( .A(n5513), .ZN(n5512) );
  OAI21_X1 U5558 ( .B1(n8749), .B2(n5514), .A(n8751), .ZN(n5513) );
  INV_X1 U5559 ( .A(n7920), .ZN(n5514) );
  AND2_X1 U5560 ( .A1(n5142), .A2(n5544), .ZN(n5542) );
  OR2_X1 U5561 ( .A1(n9070), .A2(n5088), .ZN(n5544) );
  NAND2_X1 U5562 ( .A1(n8462), .A2(n8471), .ZN(n5222) );
  INV_X1 U5563 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U5564 ( .A1(n6058), .A2(n5145), .ZN(n5655) );
  INV_X1 U5565 ( .A(n6057), .ZN(n5656) );
  NAND2_X1 U5566 ( .A1(n5913), .A2(n6947), .ZN(n5870) );
  AOI21_X1 U5567 ( .B1(n5264), .B2(n5265), .A(n9748), .ZN(n5263) );
  INV_X1 U5568 ( .A(n5266), .ZN(n5265) );
  OR3_X1 U5569 ( .A1(n9780), .A2(n9757), .A3(n9772), .ZN(n9879) );
  NOR2_X1 U5570 ( .A1(n10245), .A2(n5364), .ZN(n5363) );
  INV_X1 U5571 ( .A(n5365), .ZN(n5364) );
  NOR2_X1 U5572 ( .A1(n10248), .A2(n10254), .ZN(n5365) );
  NOR2_X1 U5573 ( .A1(n5705), .A2(n5702), .ZN(n5701) );
  INV_X1 U5574 ( .A(n5708), .ZN(n5702) );
  NOR2_X1 U5575 ( .A1(n9760), .A2(n5670), .ZN(n5669) );
  INV_X1 U5576 ( .A(n9864), .ZN(n5670) );
  NOR2_X1 U5577 ( .A1(n8259), .A2(n10307), .ZN(n5346) );
  NOR2_X1 U5578 ( .A1(n9808), .A2(n5715), .ZN(n5713) );
  INV_X1 U5579 ( .A(n9676), .ZN(n9683) );
  NAND2_X1 U5580 ( .A1(n5324), .A2(n5323), .ZN(n5661) );
  INV_X1 U5581 ( .A(n9854), .ZN(n5324) );
  NAND2_X1 U5582 ( .A1(n9849), .A2(n11012), .ZN(n5323) );
  NAND2_X1 U5583 ( .A1(n11050), .A2(n7722), .ZN(n5693) );
  NAND2_X1 U5584 ( .A1(n9668), .A2(n5694), .ZN(n5692) );
  NAND2_X1 U5585 ( .A1(n10978), .A2(n10946), .ZN(n5349) );
  NAND2_X1 U5586 ( .A1(n6627), .A2(n6626), .ZN(n8385) );
  NAND2_X1 U5587 ( .A1(n5472), .A2(n6504), .ZN(n5471) );
  INV_X1 U5588 ( .A(n6537), .ZN(n5472) );
  INV_X1 U5589 ( .A(n5470), .ZN(n5469) );
  OAI21_X1 U5590 ( .B1(n5473), .B2(n5471), .A(n6536), .ZN(n5470) );
  AOI21_X1 U5591 ( .B1(n5450), .B2(n5448), .A(n5194), .ZN(n5447) );
  INV_X1 U5592 ( .A(n5451), .ZN(n5448) );
  INV_X1 U5593 ( .A(n5450), .ZN(n5449) );
  AND4_X1 U5594 ( .A1(n5791), .A2(n10721), .A3(n10729), .A4(n10730), .ZN(n5771) );
  AND2_X1 U5595 ( .A1(n6372), .A2(n6353), .ZN(n6370) );
  INV_X1 U5596 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5770) );
  AOI21_X1 U5597 ( .B1(n5461), .B2(n6111), .A(n5460), .ZN(n5459) );
  INV_X1 U5598 ( .A(n6139), .ZN(n5460) );
  NAND2_X1 U5599 ( .A1(n6042), .A2(n10618), .ZN(n6059) );
  NAND2_X1 U5600 ( .A1(n5907), .A2(n5906), .ZN(n5928) );
  OR2_X1 U5601 ( .A1(n7036), .A2(n5905), .ZN(n5907) );
  AND2_X1 U5602 ( .A1(n5227), .A2(n5223), .ZN(n5827) );
  OR2_X1 U5603 ( .A1(n5730), .A2(n5141), .ZN(n5726) );
  INV_X1 U5604 ( .A(n5729), .ZN(n5728) );
  NAND2_X1 U5605 ( .A1(n7762), .A2(n7827), .ZN(n5733) );
  XNOR2_X1 U5606 ( .A(n8628), .B(n5099), .ZN(n8829) );
  NAND2_X1 U5607 ( .A1(n5751), .A2(n5755), .ZN(n5749) );
  OR2_X1 U5608 ( .A1(n7406), .A2(n7243), .ZN(n5755) );
  NAND2_X1 U5609 ( .A1(n8927), .A2(n8926), .ZN(n8925) );
  NAND2_X1 U5610 ( .A1(n8818), .A2(n8562), .ZN(n5747) );
  AND2_X1 U5611 ( .A1(n5552), .A2(n6705), .ZN(n5443) );
  OR4_X1 U5612 ( .A1(n8773), .A2(n8772), .A3(n8881), .A4(n8771), .ZN(n8775) );
  NAND2_X1 U5613 ( .A1(n7186), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6860) );
  OR2_X1 U5614 ( .A1(n7186), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6861) );
  OR2_X1 U5615 ( .A1(n7186), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6870) );
  NAND2_X1 U5616 ( .A1(n6662), .A2(n9510), .ZN(n6713) );
  NAND2_X1 U5617 ( .A1(n5492), .A2(n7235), .ZN(n5491) );
  NAND2_X1 U5618 ( .A1(n6894), .A2(n6893), .ZN(n5493) );
  NOR2_X1 U5619 ( .A1(n5103), .A2(n7073), .ZN(n5211) );
  OR2_X1 U5620 ( .A1(n7279), .A2(n7280), .ZN(n5501) );
  XNOR2_X1 U5621 ( .A(n7513), .B(n7512), .ZN(n10345) );
  NOR2_X1 U5622 ( .A1(n7516), .A2(n7515), .ZN(n7660) );
  AOI21_X1 U5623 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7670), .A(n7660), .ZN(
        n7845) );
  NOR2_X1 U5624 ( .A1(n7857), .A2(n7856), .ZN(n8051) );
  OR2_X1 U5625 ( .A1(n8051), .A2(n5593), .ZN(n5592) );
  NOR2_X1 U5626 ( .A1(n7937), .A2(n5594), .ZN(n5593) );
  NAND2_X1 U5627 ( .A1(n5595), .A2(n5596), .ZN(n5598) );
  INV_X1 U5628 ( .A(n8239), .ZN(n5596) );
  NAND2_X1 U5629 ( .A1(n5600), .A2(n5599), .ZN(n8327) );
  AOI21_X1 U5630 ( .B1(n8239), .B2(n5601), .A(n9087), .ZN(n5599) );
  NAND2_X1 U5631 ( .A1(n8240), .A2(n5601), .ZN(n5600) );
  INV_X1 U5632 ( .A(n8324), .ZN(n5601) );
  NAND2_X1 U5633 ( .A1(n9078), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9077) );
  NOR2_X1 U5634 ( .A1(n9091), .A2(n8331), .ZN(n8332) );
  OR2_X1 U5635 ( .A1(n9119), .A2(n8297), .ZN(n5497) );
  NOR2_X1 U5636 ( .A1(n8357), .A2(n8356), .ZN(n8364) );
  NAND2_X1 U5637 ( .A1(n8737), .A2(n8736), .ZN(n8881) );
  XNOR2_X1 U5638 ( .A(n8877), .B(n9058), .ZN(n9183) );
  NAND2_X1 U5639 ( .A1(n8723), .A2(n8724), .ZN(n9198) );
  XNOR2_X1 U5640 ( .A(n9392), .B(n9224), .ZN(n9216) );
  OAI21_X1 U5641 ( .B1(n8869), .B2(n5133), .A(n5524), .ZN(n9222) );
  INV_X1 U5642 ( .A(n5525), .ZN(n5524) );
  OAI21_X1 U5643 ( .B1(n5526), .B2(n5133), .A(n8872), .ZN(n5525) );
  AOI21_X1 U5644 ( .B1(n5534), .B2(n5533), .A(n5156), .ZN(n5532) );
  OR2_X1 U5645 ( .A1(n9295), .A2(n8826), .ZN(n9273) );
  AND2_X1 U5646 ( .A1(n9273), .A2(n8738), .ZN(n9293) );
  NAND2_X1 U5647 ( .A1(n9302), .A2(n9307), .ZN(n9301) );
  NAND2_X1 U5648 ( .A1(n8707), .A2(n8574), .ZN(n9324) );
  AOI21_X1 U5649 ( .B1(n5531), .B2(n5530), .A(n5527), .ZN(n9346) );
  AND2_X1 U5650 ( .A1(n8858), .A2(n8182), .ZN(n5530) );
  NAND2_X1 U5651 ( .A1(n5164), .A2(n5528), .ZN(n5527) );
  NAND2_X1 U5652 ( .A1(n5516), .A2(n5519), .ZN(n8176) );
  NAND2_X1 U5653 ( .A1(n5523), .A2(n5517), .ZN(n5516) );
  NOR2_X1 U5654 ( .A1(n8518), .A2(n8115), .ZN(n5517) );
  NAND2_X1 U5655 ( .A1(n8135), .A2(n8518), .ZN(n8166) );
  NAND2_X1 U5656 ( .A1(n8008), .A2(n8007), .ZN(n8116) );
  AND2_X1 U5657 ( .A1(n7730), .A2(n8499), .ZN(n5445) );
  INV_X1 U5658 ( .A(n9363), .ZN(n9291) );
  INV_X1 U5659 ( .A(n7120), .ZN(n9289) );
  NAND2_X1 U5660 ( .A1(n8418), .A2(n8417), .ZN(n8896) );
  NAND2_X1 U5661 ( .A1(n8581), .A2(n8580), .ZN(n8934) );
  NAND2_X1 U5662 ( .A1(n8539), .A2(n8538), .ZN(n8964) );
  NAND2_X1 U5663 ( .A1(n5321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6700) );
  AOI22_X1 U5664 ( .A1(n6319), .A2(n5640), .B1(n5642), .B2(n9611), .ZN(n5639)
         );
  INV_X1 U5665 ( .A(n6295), .ZN(n5640) );
  NAND2_X1 U5666 ( .A1(n6295), .A2(n5643), .ZN(n5642) );
  AND2_X1 U5667 ( .A1(n5632), .A2(n6221), .ZN(n5627) );
  NAND2_X1 U5668 ( .A1(n6219), .A2(n6220), .ZN(n8202) );
  AND2_X1 U5669 ( .A1(n5632), .A2(n8204), .ZN(n5630) );
  NAND2_X1 U5670 ( .A1(n5633), .A2(n9631), .ZN(n5632) );
  NOR2_X1 U5671 ( .A1(n5633), .A2(n9631), .ZN(n5629) );
  NAND2_X1 U5672 ( .A1(n5135), .A2(n5183), .ZN(n5644) );
  XNOR2_X1 U5673 ( .A(n5941), .B(n6636), .ZN(n5949) );
  XNOR2_X1 U5674 ( .A(n5916), .B(n6636), .ZN(n5943) );
  NAND2_X1 U5675 ( .A1(n9574), .A2(n6294), .ZN(n6296) );
  NAND2_X1 U5676 ( .A1(n5634), .A2(n8203), .ZN(n5631) );
  NAND2_X1 U5677 ( .A1(n6222), .A2(n6221), .ZN(n8203) );
  INV_X1 U5678 ( .A(n5780), .ZN(n5877) );
  INV_X1 U5679 ( .A(n5363), .ZN(n5362) );
  INV_X1 U5680 ( .A(n10065), .ZN(n10081) );
  NAND2_X1 U5681 ( .A1(n9736), .A2(n9735), .ZN(n9789) );
  AND2_X1 U5682 ( .A1(n10056), .A2(n10047), .ZN(n10050) );
  NAND2_X1 U5683 ( .A1(n10130), .A2(n5678), .ZN(n5679) );
  OR2_X1 U5684 ( .A1(n10094), .A2(n10004), .ZN(n5674) );
  NOR2_X1 U5685 ( .A1(n10094), .A2(n5677), .ZN(n5676) );
  INV_X1 U5686 ( .A(n9898), .ZN(n10115) );
  NAND2_X1 U5687 ( .A1(n5333), .A2(n5149), .ZN(n10144) );
  AOI21_X1 U5688 ( .B1(n5708), .B2(n5111), .A(n5120), .ZN(n5706) );
  AND2_X1 U5689 ( .A1(n9793), .A2(n10156), .ZN(n10176) );
  INV_X1 U5690 ( .A(n9869), .ZN(n5667) );
  NAND2_X1 U5691 ( .A1(n9758), .A2(n5669), .ZN(n5668) );
  NAND2_X1 U5692 ( .A1(n5329), .A2(n5326), .ZN(n8265) );
  NAND2_X1 U5693 ( .A1(n5167), .A2(n9700), .ZN(n5329) );
  NAND2_X1 U5694 ( .A1(n8265), .A2(n10014), .ZN(n9758) );
  NAND2_X1 U5695 ( .A1(n8041), .A2(n8040), .ZN(n5717) );
  AND2_X1 U5696 ( .A1(n9860), .A2(n9694), .ZN(n9810) );
  NAND2_X1 U5697 ( .A1(n5681), .A2(n7966), .ZN(n5680) );
  INV_X1 U5698 ( .A(n5685), .ZN(n5684) );
  INV_X1 U5699 ( .A(n9905), .ZN(n7722) );
  NOR2_X1 U5700 ( .A1(n7704), .A2(n7712), .ZN(n7723) );
  OR2_X1 U5701 ( .A1(n10338), .A2(n7528), .ZN(n11010) );
  NOR2_X1 U5702 ( .A1(n7523), .A2(n6947), .ZN(n7749) );
  AND2_X1 U5703 ( .A1(n10338), .A2(n9787), .ZN(n10969) );
  NAND2_X1 U5704 ( .A1(n6797), .A2(n5820), .ZN(n5357) );
  AND2_X1 U5705 ( .A1(n6598), .A2(n7908), .ZN(n11006) );
  NAND2_X1 U5706 ( .A1(n5771), .A2(n10735), .ZN(n5723) );
  NAND2_X1 U5707 ( .A1(n5776), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5773) );
  XNOR2_X1 U5708 ( .A(n8385), .B(n8384), .ZN(n8406) );
  XNOR2_X1 U5709 ( .A(n6506), .B(n6501), .ZN(n8436) );
  XNOR2_X1 U5710 ( .A(n6397), .B(n6412), .ZN(n8618) );
  NAND2_X1 U5711 ( .A1(n6396), .A2(n6419), .ZN(n6397) );
  XNOR2_X1 U5712 ( .A(n6374), .B(n6415), .ZN(n8614) );
  INV_X1 U5713 ( .A(n6416), .ZN(n6374) );
  INV_X1 U5714 ( .A(n5424), .ZN(n6298) );
  AOI21_X1 U5715 ( .B1(n6248), .B2(n5429), .A(n5427), .ZN(n5424) );
  NAND2_X1 U5716 ( .A1(n5699), .A2(n5695), .ZN(n5696) );
  OAI21_X1 U5717 ( .B1(n6112), .B2(n5457), .A(n5455), .ZN(n6194) );
  NAND2_X1 U5718 ( .A1(n5252), .A2(n6110), .ZN(n6141) );
  XNOR2_X1 U5719 ( .A(n6084), .B(n5765), .ZN(n7807) );
  NAND2_X1 U5720 ( .A1(n5253), .A2(n6059), .ZN(n6084) );
  OR2_X1 U5721 ( .A1(n6061), .A2(n6060), .ZN(n5253) );
  NAND2_X1 U5722 ( .A1(n5964), .A2(n5963), .ZN(n5981) );
  NAND2_X1 U5723 ( .A1(n5414), .A2(n5904), .ZN(n5927) );
  NAND2_X1 U5724 ( .A1(n9022), .A2(n8823), .ZN(n8937) );
  INV_X1 U5725 ( .A(n9059), .ZN(n9224) );
  AOI21_X1 U5726 ( .B1(n5297), .B2(n5296), .A(n5190), .ZN(n5295) );
  INV_X1 U5727 ( .A(n5299), .ZN(n5296) );
  INV_X1 U5728 ( .A(n9062), .ZN(n9007) );
  NAND2_X1 U5729 ( .A1(n5316), .A2(n5314), .ZN(n9012) );
  AOI21_X1 U5730 ( .B1(n5317), .B2(n5318), .A(n5315), .ZN(n5314) );
  INV_X1 U5731 ( .A(n9013), .ZN(n5315) );
  OAI21_X1 U5732 ( .B1(n9022), .B2(n5318), .A(n5317), .ZN(n9014) );
  AND2_X1 U5733 ( .A1(n5418), .A2(n5417), .ZN(n8787) );
  INV_X1 U5734 ( .A(n6834), .ZN(n8788) );
  XNOR2_X1 U5735 ( .A(n7496), .B(n7512), .ZN(n10344) );
  NAND2_X1 U5736 ( .A1(n5408), .A2(n5407), .ZN(n5406) );
  NOR2_X1 U5737 ( .A1(n10763), .A2(n10762), .ZN(n5407) );
  INV_X1 U5738 ( .A(n10764), .ZN(n5408) );
  NAND2_X1 U5739 ( .A1(n5412), .A2(n5411), .ZN(n5410) );
  NOR2_X1 U5740 ( .A1(n10753), .A2(n10752), .ZN(n5411) );
  NAND2_X1 U5741 ( .A1(n5413), .A2(n10754), .ZN(n5412) );
  AND3_X1 U5742 ( .A1(n8327), .A2(n5597), .A3(P2_REG2_REG_13__SCAN_IN), .ZN(
        n9075) );
  OR2_X1 U5743 ( .A1(n5607), .A2(n8364), .ZN(n5606) );
  OR2_X1 U5744 ( .A1(n8363), .A2(n8361), .ZN(n5607) );
  NAND2_X1 U5745 ( .A1(n9159), .A2(n5200), .ZN(n5481) );
  INV_X1 U5746 ( .A(n5604), .ZN(n5603) );
  AOI21_X1 U5747 ( .B1(n8367), .B2(n10352), .A(n8366), .ZN(n5604) );
  INV_X1 U5748 ( .A(n8894), .ZN(n5440) );
  NAND2_X1 U5749 ( .A1(n7446), .A2(n11102), .ZN(n11111) );
  INV_X1 U5750 ( .A(n6765), .ZN(n6768) );
  NAND2_X1 U5751 ( .A1(n6331), .A2(n6330), .ZN(n10293) );
  NAND2_X1 U5752 ( .A1(n6048), .A2(n6047), .ZN(n9543) );
  NAND2_X1 U5753 ( .A1(n6462), .A2(n6461), .ZN(n10268) );
  NAND2_X1 U5754 ( .A1(n6309), .A2(n6308), .ZN(n10299) );
  NAND2_X1 U5755 ( .A1(n6512), .A2(n6511), .ZN(n10259) );
  NAND2_X1 U5756 ( .A1(n8426), .A2(n9644), .ZN(n6512) );
  AND2_X1 U5757 ( .A1(n6600), .A2(n6595), .ZN(n9633) );
  AOI21_X1 U5758 ( .B1(n9829), .B2(n9828), .A(n7908), .ZN(n9830) );
  AND2_X1 U5759 ( .A1(n9647), .A2(n9646), .ZN(n10239) );
  AND2_X1 U5760 ( .A1(n6607), .A2(n6552), .ZN(n10066) );
  OR2_X1 U5761 ( .A1(n6943), .A2(n6939), .ZN(n10227) );
  OAI21_X1 U5762 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(n10404) );
  AOI22_X1 U5763 ( .A1(n10589), .A2(keyinput_131), .B1(SI_30_), .B2(
        keyinput_130), .ZN(n10588) );
  AND2_X1 U5764 ( .A1(n5568), .A2(n5567), .ZN(n5566) );
  NAND2_X1 U5765 ( .A1(n10412), .A2(SI_13_), .ZN(n5567) );
  NAND2_X1 U5766 ( .A1(n10613), .A2(keyinput_19), .ZN(n5568) );
  NAND2_X1 U5767 ( .A1(n5565), .A2(n5563), .ZN(n10419) );
  NOR2_X1 U5768 ( .A1(n10415), .A2(n5564), .ZN(n5563) );
  OAI21_X1 U5769 ( .B1(n10411), .B2(n5193), .A(n5566), .ZN(n5565) );
  XNOR2_X1 U5770 ( .A(SI_11_), .B(keyinput_21), .ZN(n5564) );
  AND2_X1 U5771 ( .A1(n10616), .A2(n5390), .ZN(n5389) );
  XNOR2_X1 U5772 ( .A(n5391), .B(SI_12_), .ZN(n5390) );
  INV_X1 U5773 ( .A(keyinput_148), .ZN(n5391) );
  AOI21_X1 U5774 ( .B1(n5384), .B2(n10639), .A(n5383), .ZN(n10646) );
  OR2_X1 U5775 ( .A1(n10638), .A2(n10637), .ZN(n5383) );
  NAND2_X1 U5776 ( .A1(n5386), .A2(n5385), .ZN(n5384) );
  NAND2_X1 U5777 ( .A1(n5588), .A2(n5587), .ZN(n5586) );
  NAND2_X1 U5778 ( .A1(n10450), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U5779 ( .A1(n10655), .A2(keyinput_48), .ZN(n5588) );
  AND2_X1 U5780 ( .A1(n5585), .A2(n5584), .ZN(n5583) );
  NAND2_X1 U5781 ( .A1(n10451), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U5782 ( .A1(n10658), .A2(keyinput_49), .ZN(n5585) );
  NAND2_X1 U5783 ( .A1(n10660), .A2(keyinput_51), .ZN(n5580) );
  NAND2_X1 U5784 ( .A1(n10453), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5579) );
  INV_X1 U5785 ( .A(n5398), .ZN(n5397) );
  OAI22_X1 U5786 ( .A1(n10657), .A2(n10658), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        keyinput_177), .ZN(n5398) );
  OAI22_X1 U5787 ( .A1(n7023), .A2(keyinput_178), .B1(n10659), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n5396) );
  AND2_X1 U5788 ( .A1(n10663), .A2(n10664), .ZN(n5393) );
  NOR4_X1 U5789 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10469) );
  OAI21_X1 U5790 ( .B1(n5395), .B2(n5394), .A(n5392), .ZN(n10669) );
  OAI22_X1 U5791 ( .A1(n10660), .A2(keyinput_179), .B1(n10661), .B2(
        P2_REG3_REG_24__SCAN_IN), .ZN(n5394) );
  AND2_X1 U5792 ( .A1(n10662), .A2(n5393), .ZN(n5392) );
  AOI21_X1 U5793 ( .B1(n10656), .B2(n5397), .A(n5396), .ZN(n5395) );
  NAND2_X1 U5794 ( .A1(n9667), .A2(n9747), .ZN(n5241) );
  NAND2_X1 U5795 ( .A1(n9666), .A2(n9742), .ZN(n5240) );
  INV_X1 U5796 ( .A(keyinput_198), .ZN(n5382) );
  AND2_X1 U5797 ( .A1(n5243), .A2(n5235), .ZN(n9696) );
  AND2_X1 U5798 ( .A1(n5245), .A2(n5244), .ZN(n5243) );
  NAND2_X1 U5799 ( .A1(n9686), .A2(n9742), .ZN(n5245) );
  NAND2_X1 U5800 ( .A1(n5571), .A2(n5570), .ZN(n5569) );
  NAND2_X1 U5801 ( .A1(n10482), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U5802 ( .A1(n6424), .A2(keyinput_73), .ZN(n5571) );
  AND2_X1 U5803 ( .A1(n5574), .A2(n5573), .ZN(n5572) );
  NAND2_X1 U5804 ( .A1(n10481), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U5805 ( .A1(n10688), .A2(keyinput_72), .ZN(n5574) );
  INV_X1 U5806 ( .A(n5377), .ZN(n5376) );
  OAI22_X1 U5807 ( .A1(n6424), .A2(n10690), .B1(P2_DATAO_REG_23__SCAN_IN), 
        .B2(keyinput_201), .ZN(n5377) );
  OAI22_X1 U5808 ( .A1(n10688), .A2(keyinput_200), .B1(n10689), .B2(
        P2_DATAO_REG_24__SCAN_IN), .ZN(n5378) );
  AOI21_X1 U5809 ( .B1(n5575), .B2(n5572), .A(n5569), .ZN(n10489) );
  OAI21_X1 U5810 ( .B1(n5379), .B2(n5378), .A(n5376), .ZN(n10691) );
  AND2_X1 U5811 ( .A1(n10694), .A2(keyinput_204), .ZN(n5405) );
  NAND2_X1 U5812 ( .A1(n10695), .A2(keyinput_205), .ZN(n5403) );
  INV_X1 U5813 ( .A(n10505), .ZN(n5562) );
  XNOR2_X1 U5814 ( .A(n10506), .B(n5561), .ZN(n5560) );
  INV_X1 U5815 ( .A(keyinput_89), .ZN(n5561) );
  XNOR2_X1 U5816 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n5399)
         );
  AOI21_X1 U5817 ( .B1(n5400), .B2(n5198), .A(n5399), .ZN(n10697) );
  NAND2_X1 U5818 ( .A1(n5292), .A2(n5291), .ZN(n5290) );
  INV_X1 U5819 ( .A(n9714), .ZN(n5291) );
  OAI21_X1 U5820 ( .B1(n10521), .B2(n10520), .A(n10519), .ZN(n5558) );
  INV_X1 U5821 ( .A(n10526), .ZN(n5555) );
  INV_X1 U5822 ( .A(n5557), .ZN(n5556) );
  OAI22_X1 U5823 ( .A1(n10719), .A2(n10522), .B1(P1_IR_REG_11__SCAN_IN), .B2(
        keyinput_101), .ZN(n5557) );
  AOI21_X1 U5824 ( .B1(n10076), .B2(n9769), .A(n5282), .ZN(n5281) );
  INV_X1 U5825 ( .A(n9723), .ZN(n5282) );
  INV_X1 U5826 ( .A(n10716), .ZN(n5374) );
  OR2_X1 U5827 ( .A1(n9684), .A2(n9680), .ZN(n9856) );
  NAND2_X1 U5828 ( .A1(n9683), .A2(n9693), .ZN(n9857) );
  INV_X1 U5829 ( .A(SI_26_), .ZN(n10597) );
  INV_X1 U5830 ( .A(SI_17_), .ZN(n10606) );
  NOR3_X1 U5831 ( .A1(n10539), .A2(n10538), .A3(n10537), .ZN(n10543) );
  NAND2_X1 U5832 ( .A1(n5373), .A2(n5372), .ZN(n5371) );
  AOI21_X1 U5833 ( .B1(n10719), .B2(keyinput_229), .A(n5205), .ZN(n5372) );
  NAND2_X1 U5834 ( .A1(n5375), .A2(n5374), .ZN(n5373) );
  INV_X1 U5835 ( .A(n10733), .ZN(n5370) );
  INV_X1 U5836 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5760) );
  INV_X1 U5837 ( .A(n9740), .ZN(n5256) );
  AOI21_X1 U5838 ( .B1(n5121), .B2(n5273), .A(n5166), .ZN(n5271) );
  NOR2_X1 U5839 ( .A1(n9679), .A2(n7716), .ZN(n9849) );
  AND2_X1 U5840 ( .A1(n9802), .A2(n7719), .ZN(n9854) );
  INV_X1 U5841 ( .A(SI_23_), .ZN(n10599) );
  AND2_X1 U5842 ( .A1(n6372), .A2(n6347), .ZN(n5451) );
  INV_X1 U5843 ( .A(SI_19_), .ZN(n10582) );
  INV_X1 U5844 ( .A(SI_18_), .ZN(n10583) );
  INV_X1 U5845 ( .A(n5426), .ZN(n5425) );
  OAI21_X1 U5846 ( .B1(n5427), .B2(n5429), .A(n6297), .ZN(n5426) );
  INV_X1 U5847 ( .A(SI_15_), .ZN(n10379) );
  INV_X1 U5848 ( .A(SI_10_), .ZN(n10414) );
  NAND2_X1 U5849 ( .A1(n6063), .A2(n10619), .ZN(n6085) );
  INV_X1 U5850 ( .A(n7583), .ZN(n5307) );
  NAND2_X1 U5851 ( .A1(n7645), .A2(n9068), .ZN(n5312) );
  INV_X1 U5852 ( .A(n5131), .ZN(n5730) );
  NOR2_X1 U5853 ( .A1(n8542), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8541) );
  AND2_X1 U5854 ( .A1(n8598), .A2(n7024), .ZN(n8608) );
  AND2_X1 U5855 ( .A1(n8541), .A2(n7023), .ZN(n8555) );
  NAND2_X1 U5856 ( .A1(n8405), .A2(n8732), .ZN(n8677) );
  INV_X1 U5857 ( .A(n8786), .ZN(n5217) );
  AOI21_X1 U5858 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n6898), .A(n6897), .ZN(
        n6899) );
  INV_X1 U5859 ( .A(n7072), .ZN(n6901) );
  NOR2_X1 U5860 ( .A1(n7177), .A2(n7176), .ZN(n7278) );
  NOR2_X1 U5861 ( .A1(n5103), .A2(n10942), .ZN(n7176) );
  AOI21_X1 U5862 ( .B1(n5369), .B2(n5368), .A(n5367), .ZN(n10747) );
  AND2_X1 U5863 ( .A1(n10732), .A2(n10731), .ZN(n5368) );
  NAND2_X1 U5864 ( .A1(n10742), .A2(n10741), .ZN(n5367) );
  NAND2_X1 U5865 ( .A1(n5371), .A2(n5370), .ZN(n5369) );
  NAND2_X1 U5866 ( .A1(n5499), .A2(n5498), .ZN(n7513) );
  NAND2_X1 U5867 ( .A1(n7561), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5498) );
  AND2_X1 U5868 ( .A1(n5505), .A2(n5504), .ZN(n8296) );
  NAND2_X1 U5869 ( .A1(n8330), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5504) );
  AND2_X1 U5870 ( .A1(n6672), .A2(n6671), .ZN(n6681) );
  OR2_X1 U5871 ( .A1(n8336), .A2(n9165), .ZN(n8359) );
  AND2_X1 U5872 ( .A1(n9246), .A2(n8868), .ZN(n5526) );
  OR2_X1 U5873 ( .A1(n8628), .A2(n9261), .ZN(n8865) );
  OR2_X1 U5874 ( .A1(n8964), .A2(n9051), .ZN(n8740) );
  NAND2_X1 U5875 ( .A1(n8858), .A2(n5529), .ZN(n5528) );
  INV_X1 U5876 ( .A(n8855), .ZN(n5529) );
  NOR2_X1 U5877 ( .A1(n8108), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8107) );
  AND2_X1 U5878 ( .A1(n7551), .A2(n7021), .ZN(n7649) );
  INV_X1 U5879 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10658) );
  OR2_X1 U5880 ( .A1(n10336), .A2(n8399), .ZN(n8401) );
  AND2_X1 U5881 ( .A1(n6739), .A2(n6738), .ZN(n6761) );
  INV_X1 U5882 ( .A(n9602), .ZN(n5652) );
  NAND2_X1 U5883 ( .A1(n5844), .A2(n5857), .ZN(n5848) );
  AND2_X1 U5884 ( .A1(n6949), .A2(n5843), .ZN(n5844) );
  NAND2_X1 U5885 ( .A1(n5650), .A2(n5648), .ZN(n5647) );
  INV_X1 U5886 ( .A(n5135), .ZN(n5648) );
  NAND2_X1 U5887 ( .A1(n5649), .A2(n9521), .ZN(n5645) );
  INV_X1 U5888 ( .A(n5843), .ZN(n5837) );
  INV_X1 U5889 ( .A(n5678), .ZN(n5677) );
  NAND2_X1 U5890 ( .A1(n10168), .A2(n5355), .ZN(n5354) );
  NAND2_X1 U5891 ( .A1(n5353), .A2(n10143), .ZN(n5352) );
  INV_X1 U5892 ( .A(n5354), .ZN(n5353) );
  NOR2_X1 U5893 ( .A1(n5665), .A2(n5328), .ZN(n5325) );
  INV_X1 U5894 ( .A(n5666), .ZN(n5665) );
  INV_X1 U5895 ( .A(n5669), .ZN(n5664) );
  AND2_X1 U5896 ( .A1(n8159), .A2(n5343), .ZN(n10210) );
  NOR2_X1 U5897 ( .A1(n5345), .A2(n10234), .ZN(n5343) );
  INV_X1 U5898 ( .A(n6311), .ZN(n6310) );
  NAND2_X1 U5899 ( .A1(n8157), .A2(n9689), .ZN(n5331) );
  INV_X1 U5900 ( .A(n6256), .ZN(n6257) );
  NAND2_X1 U5901 ( .A1(n6257), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6283) );
  AND2_X1 U5902 ( .A1(n8046), .A2(n11114), .ZN(n8159) );
  AND2_X1 U5903 ( .A1(n6176), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6207) );
  NOR2_X1 U5904 ( .A1(n6123), .A2(n6122), .ZN(n6151) );
  OR2_X1 U5905 ( .A1(n6093), .A2(n6092), .ZN(n6123) );
  OR2_X1 U5906 ( .A1(n6071), .A2(n6070), .ZN(n6093) );
  NAND2_X1 U5907 ( .A1(n5973), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6005) );
  OR2_X1 U5908 ( .A1(n10123), .A2(n10268), .ZN(n10102) );
  NOR2_X1 U5909 ( .A1(n10186), .A2(n10289), .ZN(n10174) );
  NAND2_X1 U5910 ( .A1(n8387), .A2(n8386), .ZN(n8390) );
  NAND2_X1 U5911 ( .A1(n8385), .A2(n8384), .ZN(n8387) );
  NOR2_X1 U5912 ( .A1(n6505), .A2(n5474), .ZN(n5473) );
  INV_X1 U5913 ( .A(n6485), .ZN(n5474) );
  NAND2_X1 U5914 ( .A1(n5446), .A2(n5450), .ZN(n6416) );
  NAND2_X1 U5915 ( .A1(n6349), .A2(n5451), .ZN(n5446) );
  NOR2_X1 U5916 ( .A1(n6272), .A2(n5430), .ZN(n5429) );
  INV_X1 U5917 ( .A(n6246), .ZN(n5430) );
  NAND2_X1 U5918 ( .A1(n5428), .A2(n6271), .ZN(n5427) );
  NAND2_X1 U5919 ( .A1(n5429), .A2(n6247), .ZN(n5428) );
  AND2_X1 U5920 ( .A1(n5769), .A2(n5933), .ZN(n5699) );
  AOI21_X1 U5921 ( .B1(n5115), .B2(n5456), .A(n5159), .ZN(n5455) );
  INV_X1 U5922 ( .A(n5461), .ZN(n5456) );
  INV_X1 U5923 ( .A(n5115), .ZN(n5457) );
  CLKBUF_X1 U5924 ( .A(n6144), .Z(n6145) );
  NAND2_X1 U5925 ( .A1(n6059), .A2(n6044), .ZN(n6060) );
  XNOR2_X1 U5926 ( .A(n6039), .B(SI_7_), .ZN(n6036) );
  NAND2_X1 U5927 ( .A1(n5230), .A2(n5232), .ZN(n6038) );
  AOI21_X1 U5928 ( .B1(n6016), .B2(n5233), .A(n5158), .ZN(n5232) );
  NOR2_X1 U5929 ( .A1(n6015), .A2(n5231), .ZN(n5229) );
  OR2_X1 U5930 ( .A1(n7383), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7552) );
  NAND2_X1 U5931 ( .A1(n8075), .A2(n8074), .ZN(n8246) );
  INV_X1 U5932 ( .A(n5742), .ZN(n5741) );
  OAI21_X1 U5933 ( .B1(n5137), .B2(n5743), .A(n8848), .ZN(n5742) );
  AND2_X1 U5934 ( .A1(n9074), .A2(n7449), .ZN(n7144) );
  NOR2_X1 U5935 ( .A1(n5151), .A2(n5301), .ZN(n5300) );
  NOR2_X1 U5936 ( .A1(n5303), .A2(n5302), .ZN(n5301) );
  NOR2_X1 U5937 ( .A1(n7805), .A2(n5732), .ZN(n5731) );
  INV_X1 U5938 ( .A(n5733), .ZN(n5732) );
  NAND2_X1 U5939 ( .A1(n8935), .A2(n5134), .ZN(n8992) );
  NAND2_X1 U5940 ( .A1(n5122), .A2(n5110), .ZN(n5317) );
  NAND2_X1 U5941 ( .A1(n8936), .A2(n5320), .ZN(n5319) );
  NAND2_X1 U5942 ( .A1(n5110), .A2(n8936), .ZN(n5318) );
  XNOR2_X1 U5943 ( .A(n5099), .B(n8454), .ZN(n7190) );
  NAND2_X1 U5944 ( .A1(n8555), .A2(n10666), .ZN(n8582) );
  INV_X1 U5945 ( .A(n5313), .ZN(n5310) );
  NAND2_X1 U5946 ( .A1(n7582), .A2(n7567), .ZN(n5313) );
  OR2_X1 U5947 ( .A1(n7584), .A2(n7583), .ZN(n5311) );
  OR2_X1 U5948 ( .A1(n8812), .A2(n8811), .ZN(n9042) );
  NOR2_X1 U5949 ( .A1(n5130), .A2(n5302), .ZN(n5299) );
  OR2_X1 U5950 ( .A1(n6841), .A2(n6775), .ZN(n6868) );
  OR2_X1 U5951 ( .A1(n6837), .A2(n6836), .ZN(n6863) );
  NAND2_X1 U5952 ( .A1(n6868), .A2(n6867), .ZN(n6871) );
  AND2_X1 U5953 ( .A1(n6871), .A2(n6872), .ZN(n6897) );
  INV_X1 U5954 ( .A(n5490), .ZN(n5489) );
  AND2_X1 U5955 ( .A1(n5490), .A2(n5493), .ZN(n7076) );
  NOR2_X1 U5956 ( .A1(n7076), .A2(n7075), .ZN(n7177) );
  AOI22_X1 U5957 ( .A1(n5103), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n7073), .B2(
        n7175), .ZN(n7074) );
  NOR2_X1 U5958 ( .A1(n6903), .A2(n6902), .ZN(n7071) );
  AOI22_X1 U5959 ( .A1(n10345), .A2(P2_REG1_REG_7__SCAN_IN), .B1(n7513), .B2(
        n10356), .ZN(n7516) );
  NOR2_X1 U5960 ( .A1(n7847), .A2(n7846), .ZN(n7850) );
  NOR2_X1 U5961 ( .A1(n7850), .A2(n7849), .ZN(n8053) );
  INV_X1 U5962 ( .A(n5592), .ZN(n8235) );
  NAND2_X1 U5963 ( .A1(n5725), .A2(n5127), .ZN(n7126) );
  AOI21_X1 U5964 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8335), .A(n9130), .ZN(
        n8336) );
  XNOR2_X1 U5965 ( .A(n8298), .B(n9165), .ZN(n9160) );
  INV_X1 U5966 ( .A(n8359), .ZN(n8358) );
  AOI21_X1 U5967 ( .B1(n8299), .B2(n5488), .A(n8347), .ZN(n5487) );
  AND2_X1 U5968 ( .A1(n5143), .A2(n8878), .ZN(n5548) );
  NAND2_X1 U5969 ( .A1(n5545), .A2(n5549), .ZN(n9178) );
  INV_X1 U5970 ( .A(n9180), .ZN(n9209) );
  AND2_X1 U5971 ( .A1(n8655), .A2(n8721), .ZN(n9221) );
  OR2_X1 U5972 ( .A1(n8650), .A2(n8870), .ZN(n9242) );
  AND2_X1 U5973 ( .A1(n7031), .A2(n7030), .ZN(n9238) );
  OR2_X1 U5974 ( .A1(n8623), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8640) );
  NOR2_X1 U5975 ( .A1(n8640), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8639) );
  INV_X1 U5976 ( .A(n9251), .ZN(n9246) );
  NAND2_X1 U5977 ( .A1(n8869), .A2(n5526), .ZN(n9245) );
  AND2_X1 U5978 ( .A1(n8717), .A2(n8656), .ZN(n9251) );
  INV_X1 U5979 ( .A(n8859), .ZN(n9334) );
  NAND2_X1 U5980 ( .A1(n8856), .A2(n8855), .ZN(n9360) );
  INV_X1 U5981 ( .A(n5515), .ZN(n8175) );
  NAND2_X1 U5982 ( .A1(n5531), .A2(n8182), .ZN(n8856) );
  NOR2_X1 U5983 ( .A1(n5433), .A2(n5432), .ZN(n5431) );
  NOR2_X1 U5984 ( .A1(n8518), .A2(n5136), .ZN(n5433) );
  OR2_X1 U5985 ( .A1(n7942), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8009) );
  OR2_X1 U5986 ( .A1(n8009), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8108) );
  AND2_X1 U5987 ( .A1(n8514), .A2(n8512), .ZN(n8755) );
  NAND2_X1 U5988 ( .A1(n5510), .A2(n5509), .ZN(n8006) );
  AOI21_X1 U5989 ( .B1(n5512), .B2(n5514), .A(n5155), .ZN(n5509) );
  OR2_X1 U5990 ( .A1(n7733), .A2(n9068), .ZN(n5543) );
  NOR2_X1 U5991 ( .A1(n5541), .A2(n7734), .ZN(n5539) );
  NAND2_X1 U5992 ( .A1(n5542), .A2(n5132), .ZN(n5538) );
  OAI21_X1 U5993 ( .B1(n7563), .B2(n5132), .A(n5544), .ZN(n7594) );
  NAND2_X1 U5994 ( .A1(n8462), .A2(n5222), .ZN(n5435) );
  NAND2_X1 U5995 ( .A1(n7407), .A2(n8461), .ZN(n7426) );
  INV_X1 U5996 ( .A(n5222), .ZN(n8742) );
  INV_X1 U5997 ( .A(n8741), .ZN(n7350) );
  NAND2_X1 U5998 ( .A1(n6976), .A2(n6975), .ZN(n7342) );
  INV_X1 U5999 ( .A(n9074), .ZN(n5420) );
  NAND2_X1 U6000 ( .A1(n8394), .A2(n8393), .ZN(n9175) );
  NAND2_X1 U6001 ( .A1(n5521), .A2(n8114), .ZN(n8167) );
  NAND2_X1 U6002 ( .A1(n5523), .A2(n5522), .ZN(n5521) );
  INV_X1 U6003 ( .A(n5321), .ZN(n6690) );
  NOR2_X1 U6004 ( .A1(n6105), .A2(n5089), .ZN(n5654) );
  NAND2_X1 U6005 ( .A1(n6106), .A2(n6105), .ZN(n7794) );
  NOR2_X1 U6006 ( .A1(n6005), .A2(n6004), .ZN(n6028) );
  OR2_X1 U6007 ( .A1(n9550), .A2(n9549), .ZN(n5206) );
  AND3_X1 U6008 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5973) );
  AND2_X1 U6009 ( .A1(n6482), .A2(n6481), .ZN(n9581) );
  CLKBUF_X1 U6010 ( .A(n8025), .Z(n8026) );
  AOI21_X1 U6011 ( .B1(n5839), .B2(n5090), .A(n5838), .ZN(n5851) );
  NAND2_X1 U6012 ( .A1(n5998), .A2(n5997), .ZN(n5657) );
  INV_X1 U6013 ( .A(n5996), .ZN(n5997) );
  INV_X1 U6014 ( .A(n6231), .ZN(n6232) );
  NAND2_X1 U6015 ( .A1(n6232), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6256) );
  INV_X1 U6016 ( .A(n5333), .ZN(n10000) );
  AOI21_X1 U6017 ( .B1(n5263), .B2(n5262), .A(n9822), .ZN(n5261) );
  OR2_X1 U6018 ( .A1(n9741), .A2(n5260), .ZN(n5259) );
  INV_X1 U6019 ( .A(n5264), .ZN(n5262) );
  OR2_X1 U6020 ( .A1(n5954), .A2(n5875), .ZN(n5881) );
  AOI21_X1 U6021 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6800), .A(n6817), .ZN(
        n10865) );
  AOI21_X1 U6022 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6932), .A(n6931), .ZN(
        n6935) );
  AOI21_X1 U6023 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7317), .A(n7316), .ZN(
        n7319) );
  AOI21_X1 U6024 ( .B1(n7881), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7880), .ZN(
        n10844) );
  OR2_X1 U6025 ( .A1(n7883), .A2(n7882), .ZN(n5219) );
  AND2_X1 U6026 ( .A1(n5219), .A2(n5218), .ZN(n8098) );
  NAND2_X1 U6027 ( .A1(n8093), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5218) );
  OR2_X1 U6028 ( .A1(n8098), .A2(n8097), .ZN(n8142) );
  INV_X1 U6029 ( .A(n9925), .ZN(n5220) );
  AND2_X1 U6030 ( .A1(n9945), .A2(n9944), .ZN(n9948) );
  AND2_X1 U6031 ( .A1(n10081), .A2(n5363), .ZN(n10033) );
  OR2_X1 U6032 ( .A1(n10336), .A2(n9730), .ZN(n9732) );
  AOI21_X1 U6033 ( .B1(n5719), .B2(n10075), .A(n5192), .ZN(n5718) );
  NOR2_X1 U6034 ( .A1(n10078), .A2(n10006), .ZN(n10058) );
  NAND2_X1 U6035 ( .A1(n10058), .A2(n10057), .ZN(n10056) );
  INV_X1 U6036 ( .A(n10051), .ZN(n10080) );
  AND2_X1 U6037 ( .A1(n5337), .A2(n5336), .ZN(n10078) );
  NOR2_X1 U6038 ( .A1(n10073), .A2(n5279), .ZN(n5336) );
  INV_X1 U6039 ( .A(n10102), .ZN(n10108) );
  NOR2_X1 U6040 ( .A1(n10186), .A2(n5354), .ZN(n10163) );
  INV_X1 U6041 ( .A(n5704), .ZN(n5703) );
  NAND2_X1 U6042 ( .A1(n10185), .A2(n5701), .ZN(n5700) );
  OAI21_X1 U6043 ( .B1(n5706), .B2(n5705), .A(n10019), .ZN(n5704) );
  OR2_X1 U6044 ( .A1(n10211), .A2(n10293), .ZN(n10186) );
  NAND2_X1 U6045 ( .A1(n6281), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6311) );
  INV_X1 U6046 ( .A(n6283), .ZN(n6281) );
  INV_X1 U6047 ( .A(n6332), .ZN(n6356) );
  NAND2_X1 U6048 ( .A1(n8159), .A2(n5346), .ZN(n8262) );
  INV_X1 U6049 ( .A(n5711), .ZN(n5710) );
  OAI22_X1 U6050 ( .A1(n9808), .A2(n5716), .B1(n9688), .B2(n8280), .ZN(n5711)
         );
  OR2_X1 U6051 ( .A1(n8043), .A2(n8040), .ZN(n9693) );
  NAND2_X1 U6052 ( .A1(n5660), .A2(n9683), .ZN(n8035) );
  NAND2_X1 U6053 ( .A1(n5659), .A2(n5129), .ZN(n5660) );
  NAND2_X1 U6054 ( .A1(n5661), .A2(n7865), .ZN(n5659) );
  NOR2_X1 U6055 ( .A1(n7903), .A2(n8043), .ZN(n8046) );
  OR2_X1 U6056 ( .A1(n7873), .A2(n7898), .ZN(n7903) );
  INV_X1 U6057 ( .A(n5661), .ZN(n7720) );
  NOR2_X1 U6058 ( .A1(n7720), .A2(n5683), .ZN(n7900) );
  AND2_X1 U6059 ( .A1(n5693), .A2(n5694), .ZN(n5690) );
  NOR2_X1 U6060 ( .A1(n5692), .A2(n5691), .ZN(n5687) );
  INV_X1 U6061 ( .A(n5693), .ZN(n5691) );
  INV_X1 U6062 ( .A(n5349), .ZN(n5347) );
  NOR2_X1 U6063 ( .A1(n7783), .A2(n10903), .ZN(n5348) );
  OR2_X1 U6064 ( .A1(n11005), .A2(n9543), .ZN(n7704) );
  NOR2_X1 U6065 ( .A1(n5349), .A2(n10903), .ZN(n10962) );
  NAND2_X1 U6066 ( .A1(n10962), .A2(n10997), .ZN(n11004) );
  NOR2_X1 U6067 ( .A1(n10903), .A2(n7692), .ZN(n10964) );
  NAND2_X1 U6068 ( .A1(n7334), .A2(n10907), .ZN(n10909) );
  NAND2_X1 U6069 ( .A1(n6633), .A2(n6632), .ZN(n10248) );
  NAND2_X1 U6070 ( .A1(n6435), .A2(n6434), .ZN(n10273) );
  OAI22_X1 U6071 ( .A1(n8683), .A2(n8682), .B1(SI_30_), .B2(n8681), .ZN(n8688)
         );
  INV_X1 U6072 ( .A(SI_29_), .ZN(n10589) );
  XNOR2_X1 U6073 ( .A(n8390), .B(n8388), .ZN(n8395) );
  NAND2_X1 U6074 ( .A1(n8395), .A2(SI_29_), .ZN(n8398) );
  INV_X1 U6075 ( .A(n5723), .ZN(n5721) );
  OAI21_X1 U6076 ( .B1(n6486), .B2(n5471), .A(n5469), .ZN(n6544) );
  OR2_X1 U6077 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  OR2_X1 U6078 ( .A1(n5797), .A2(n10736), .ZN(n5840) );
  OAI21_X1 U6079 ( .B1(n6248), .B2(n6247), .A(n6246), .ZN(n6273) );
  NAND2_X1 U6080 ( .A1(n5458), .A2(n5459), .ZN(n6170) );
  OR2_X1 U6081 ( .A1(n5984), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U6082 ( .A1(n5234), .A2(n5983), .ZN(n6017) );
  NAND2_X1 U6083 ( .A1(n5981), .A2(n5980), .ZN(n5234) );
  NAND2_X1 U6084 ( .A1(n5658), .A2(n5929), .ZN(n5961) );
  NAND2_X1 U6085 ( .A1(n5415), .A2(n5830), .ZN(n5902) );
  NAND2_X1 U6086 ( .A1(n8181), .A2(n8180), .ZN(n8916) );
  NAND2_X1 U6087 ( .A1(n8635), .A2(n8634), .ZN(n9253) );
  NAND2_X1 U6088 ( .A1(n8937), .A2(n8936), .ZN(n8935) );
  OAI21_X1 U6089 ( .B1(n5741), .B2(n8849), .A(n5736), .ZN(n5735) );
  NAND2_X1 U6090 ( .A1(n5741), .A2(n5737), .ZN(n5736) );
  NAND2_X1 U6091 ( .A1(n5743), .A2(n5738), .ZN(n5737) );
  NAND2_X1 U6092 ( .A1(n5744), .A2(n8849), .ZN(n5739) );
  NAND2_X1 U6093 ( .A1(n8408), .A2(n8407), .ZN(n8877) );
  NAND2_X1 U6094 ( .A1(n7763), .A2(n5733), .ZN(n7806) );
  XNOR2_X1 U6095 ( .A(n7190), .B(n7354), .ZN(n5724) );
  AOI21_X1 U6096 ( .B1(n7035), .B2(n7140), .A(n7144), .ZN(n7042) );
  NAND2_X1 U6097 ( .A1(n8992), .A2(n8828), .ZN(n8944) );
  NAND2_X1 U6098 ( .A1(n5304), .A2(n5303), .ZN(n8802) );
  INV_X1 U6099 ( .A(n8250), .ZN(n5304) );
  AND2_X1 U6100 ( .A1(n8956), .A2(n8955), .ZN(n8957) );
  NAND2_X1 U6101 ( .A1(n8438), .A2(n8437), .ZN(n9220) );
  NAND2_X1 U6102 ( .A1(n8554), .A2(n8553), .ZN(n9336) );
  NAND2_X1 U6103 ( .A1(n8638), .A2(n8637), .ZN(n9232) );
  INV_X1 U6104 ( .A(n5749), .ZN(n5753) );
  NAND2_X1 U6105 ( .A1(n8925), .A2(n5755), .ZN(n7244) );
  NAND2_X1 U6106 ( .A1(n5727), .A2(n5131), .ZN(n8073) );
  NAND2_X1 U6107 ( .A1(n7763), .A2(n5731), .ZN(n5727) );
  NAND2_X1 U6108 ( .A1(n8935), .A2(n8825), .ZN(n8994) );
  NAND2_X1 U6109 ( .A1(n8596), .A2(n8595), .ZN(n9295) );
  NOR2_X1 U6110 ( .A1(n9020), .A2(n5746), .ZN(n5745) );
  INV_X1 U6111 ( .A(n5747), .ZN(n5746) );
  NAND2_X1 U6112 ( .A1(n8973), .A2(n5747), .ZN(n9021) );
  INV_X1 U6113 ( .A(n9207), .ZN(n9237) );
  NAND2_X1 U6114 ( .A1(n5294), .A2(n5297), .ZN(n9046) );
  NAND2_X1 U6115 ( .A1(n8250), .A2(n5299), .ZN(n5294) );
  NOR2_X1 U6116 ( .A1(n9455), .A2(n9172), .ZN(n8786) );
  NAND2_X1 U6117 ( .A1(n5444), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6704) );
  NAND2_X1 U6118 ( .A1(n8787), .A2(n6999), .ZN(n5416) );
  INV_X1 U6119 ( .A(n5213), .ZN(n8783) );
  NAND2_X1 U6120 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6714) );
  NAND2_X1 U6121 ( .A1(n5491), .A2(n5493), .ZN(n6895) );
  NOR2_X1 U6122 ( .A1(n7167), .A2(n7168), .ZN(n7269) );
  INV_X1 U6123 ( .A(n5501), .ZN(n7282) );
  INV_X1 U6124 ( .A(n5499), .ZN(n7511) );
  NAND2_X1 U6125 ( .A1(n5618), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5617) );
  INV_X1 U6126 ( .A(n7270), .ZN(n5618) );
  INV_X1 U6127 ( .A(n10756), .ZN(n5409) );
  NAND2_X1 U6128 ( .A1(n7496), .A2(n5611), .ZN(n5609) );
  NOR2_X1 U6129 ( .A1(n5139), .A2(n10356), .ZN(n5611) );
  INV_X1 U6130 ( .A(n5479), .ZN(n8224) );
  OR2_X1 U6131 ( .A1(n8056), .A2(n8055), .ZN(n5479) );
  INV_X1 U6132 ( .A(n8223), .ZN(n5478) );
  OAI21_X1 U6133 ( .B1(n8056), .B2(n5477), .A(n5476), .ZN(n8289) );
  NAND2_X1 U6134 ( .A1(n5480), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5477) );
  INV_X1 U6135 ( .A(n8225), .ZN(n5480) );
  NAND2_X1 U6136 ( .A1(n8327), .A2(n5597), .ZN(n9076) );
  NOR2_X1 U6137 ( .A1(n9075), .A2(n8328), .ZN(n9093) );
  AND2_X1 U6138 ( .A1(n9077), .A2(n8293), .ZN(n9096) );
  NOR2_X1 U6139 ( .A1(n9112), .A2(n9368), .ZN(n9111) );
  INV_X1 U6140 ( .A(n5497), .ZN(n9141) );
  INV_X1 U6141 ( .A(n5495), .ZN(n9139) );
  OAI21_X1 U6142 ( .B1(n9112), .B2(n5620), .A(n5619), .ZN(n9130) );
  NAND2_X1 U6143 ( .A1(n5621), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U6144 ( .A1(n8333), .A2(n5621), .ZN(n5619) );
  INV_X1 U6145 ( .A(n9131), .ZN(n5621) );
  INV_X1 U6146 ( .A(n10357), .ZN(n9166) );
  OR2_X1 U6147 ( .A1(P2_U3150), .A2(n6832), .ZN(n9158) );
  OAI21_X1 U6148 ( .B1(n9197), .B2(n9287), .A(n9196), .ZN(n9388) );
  INV_X1 U6149 ( .A(n9195), .ZN(n9196) );
  OAI22_X1 U6150 ( .A1(n9194), .A2(n9193), .B1(n9291), .B2(n9224), .ZN(n9195)
         );
  NAND2_X1 U6151 ( .A1(n8428), .A2(n8427), .ZN(n9392) );
  NAND2_X1 U6152 ( .A1(n8426), .A2(n8689), .ZN(n8428) );
  NAND2_X1 U6153 ( .A1(n8620), .A2(n8619), .ZN(n9411) );
  NAND2_X1 U6154 ( .A1(n9301), .A2(n8863), .ZN(n9285) );
  NAND2_X1 U6155 ( .A1(n9427), .A2(n8707), .ZN(n9308) );
  NAND2_X1 U6156 ( .A1(n8567), .A2(n8566), .ZN(n9428) );
  NAND2_X1 U6157 ( .A1(n8536), .A2(n8535), .ZN(n9370) );
  NAND2_X1 U6158 ( .A1(n8166), .A2(n8136), .ZN(n8197) );
  NAND2_X1 U6159 ( .A1(n5511), .A2(n7920), .ZN(n7935) );
  NAND2_X1 U6160 ( .A1(n7918), .A2(n8749), .ZN(n5511) );
  NAND2_X1 U6161 ( .A1(n7729), .A2(n8499), .ZN(n7731) );
  OR2_X1 U6162 ( .A1(n7446), .A2(n9233), .ZN(n9354) );
  OAI21_X1 U6163 ( .B1(n8884), .B2(n5589), .A(n5419), .ZN(n7449) );
  NAND2_X1 U6164 ( .A1(n8884), .A2(n9520), .ZN(n5419) );
  INV_X1 U6165 ( .A(n11102), .ZN(n11086) );
  INV_X1 U6166 ( .A(n11127), .ZN(n11126) );
  INV_X1 U6167 ( .A(n9175), .ZN(n9458) );
  AND2_X1 U6168 ( .A1(n9396), .A2(n9395), .ZN(n9465) );
  AND2_X1 U6169 ( .A1(n9442), .A2(n9441), .ZN(n9500) );
  NAND2_X1 U6170 ( .A1(n8004), .A2(n8003), .ZN(n11085) );
  INV_X1 U6171 ( .A(n8454), .ZN(n7440) );
  INV_X1 U6172 ( .A(n11131), .ZN(n11128) );
  INV_X1 U6173 ( .A(n7449), .ZN(n7140) );
  NAND2_X1 U6174 ( .A1(n6765), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U6175 ( .A1(n5508), .A2(n5506), .ZN(n6851) );
  NAND2_X1 U6176 ( .A1(n5590), .A2(n5507), .ZN(n5506) );
  NAND2_X1 U6178 ( .A1(n5637), .A2(n5639), .ZN(n5636) );
  INV_X1 U6179 ( .A(n9531), .ZN(n5637) );
  INV_X1 U6180 ( .A(n5638), .ZN(n5635) );
  AND2_X1 U6181 ( .A1(n6565), .A2(n6564), .ZN(n6642) );
  NAND2_X1 U6182 ( .A1(n6376), .A2(n6375), .ZN(n10284) );
  NAND2_X1 U6183 ( .A1(n5632), .A2(n5629), .ZN(n5628) );
  NAND2_X1 U6184 ( .A1(n6222), .A2(n5627), .ZN(n5625) );
  NAND2_X1 U6185 ( .A1(n6058), .A2(n6057), .ZN(n7544) );
  NAND2_X1 U6186 ( .A1(n6399), .A2(n6398), .ZN(n10277) );
  CLKBUF_X1 U6187 ( .A(n7331), .Z(n7332) );
  AND2_X1 U6188 ( .A1(n7161), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9624) );
  AND2_X1 U6189 ( .A1(n6620), .A2(n7053), .ZN(n9623) );
  AND2_X1 U6190 ( .A1(n6620), .A2(n10338), .ZN(n9640) );
  NAND2_X1 U6191 ( .A1(n5631), .A2(n6243), .ZN(n9630) );
  OR2_X1 U6192 ( .A1(n6645), .A2(n5922), .ZN(n5923) );
  NAND2_X1 U6193 ( .A1(n5100), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5899) );
  OR2_X1 U6194 ( .A1(n6645), .A2(n5896), .ZN(n5897) );
  NOR2_X1 U6195 ( .A1(n10831), .A2(n5140), .ZN(n7057) );
  AOI21_X1 U6196 ( .B1(n7093), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7090), .ZN(
        n7092) );
  OAI21_X1 U6197 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7363), .A(n7362), .ZN(
        n7365) );
  AOI21_X1 U6198 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7478), .A(n7477), .ZN(
        n7480) );
  OAI21_X1 U6199 ( .B1(n7886), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10843), .ZN(
        n7883) );
  INV_X1 U6200 ( .A(n5219), .ZN(n8092) );
  INV_X1 U6201 ( .A(n10855), .ZN(n10862) );
  AND2_X1 U6202 ( .A1(n6789), .A2(n6795), .ZN(n10861) );
  NOR2_X1 U6203 ( .A1(n9789), .A2(n5362), .ZN(n5361) );
  NAND2_X1 U6204 ( .A1(n5673), .A2(n10972), .ZN(n5672) );
  XNOR2_X1 U6205 ( .A(n10008), .B(n5269), .ZN(n5673) );
  AND2_X1 U6206 ( .A1(n5342), .A2(n5341), .ZN(n10250) );
  AOI21_X1 U6207 ( .B1(n10052), .B2(n10969), .A(n5184), .ZN(n5341) );
  NAND2_X1 U6208 ( .A1(n10053), .A2(n10972), .ZN(n5342) );
  NAND2_X1 U6209 ( .A1(n10072), .A2(n10028), .ZN(n10055) );
  AND2_X1 U6210 ( .A1(n5679), .A2(n10004), .ZN(n10095) );
  NAND2_X1 U6211 ( .A1(n6488), .A2(n6487), .ZN(n10263) );
  NAND2_X1 U6212 ( .A1(n10130), .A2(n10003), .ZN(n10113) );
  INV_X1 U6213 ( .A(n10268), .ZN(n10111) );
  AND2_X1 U6214 ( .A1(n5333), .A2(n5332), .ZN(n10146) );
  NAND2_X1 U6215 ( .A1(n10175), .A2(n9793), .ZN(n10157) );
  NAND2_X1 U6216 ( .A1(n5707), .A2(n5706), .ZN(n10155) );
  NAND2_X1 U6217 ( .A1(n10185), .A2(n5708), .ZN(n5707) );
  AOI21_X1 U6218 ( .B1(n10185), .B2(n10018), .A(n5111), .ZN(n10171) );
  AND2_X1 U6219 ( .A1(n5668), .A2(n5666), .ZN(n10196) );
  NAND2_X1 U6220 ( .A1(n5668), .A2(n9869), .ZN(n10205) );
  NAND2_X1 U6221 ( .A1(n9758), .A2(n9864), .ZN(n10221) );
  NAND2_X1 U6222 ( .A1(n6230), .A2(n6229), .ZN(n8259) );
  AOI21_X1 U6223 ( .B1(n8042), .B2(n5714), .A(n5766), .ZN(n8273) );
  NAND2_X1 U6224 ( .A1(n6175), .A2(n6174), .ZN(n8220) );
  NAND2_X1 U6225 ( .A1(n8042), .A2(n5717), .ZN(n8155) );
  NAND2_X1 U6226 ( .A1(n7807), .A2(n9644), .ZN(n6069) );
  OAI21_X1 U6227 ( .B1(n7699), .B2(n9668), .A(n5694), .ZN(n7714) );
  NOR2_X1 U6228 ( .A1(n10180), .A2(n7638), .ZN(n10982) );
  OR2_X1 U6229 ( .A1(n11028), .A2(n7534), .ZN(n11031) );
  INV_X1 U6230 ( .A(n10982), .ZN(n10220) );
  OR2_X1 U6231 ( .A1(n6787), .A2(n6790), .ZN(n5873) );
  NAND2_X1 U6232 ( .A1(n5108), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5874) );
  AND2_X1 U6233 ( .A1(n5822), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n5356) );
  INV_X1 U6234 ( .A(n11031), .ZN(n10235) );
  NOR2_X1 U6235 ( .A1(n5723), .A2(n5157), .ZN(n5722) );
  CLKBUF_X1 U6236 ( .A(n6574), .Z(n8140) );
  INV_X1 U6237 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6747) );
  AOI21_X1 U6238 ( .B1(n5410), .B2(n5409), .A(n5406), .ZN(n10765) );
  AOI21_X1 U6239 ( .B1(n5605), .B2(n6873), .A(n5603), .ZN(n5602) );
  OR2_X1 U6240 ( .A1(n8368), .A2(n10346), .ZN(n5608) );
  NAND2_X1 U6241 ( .A1(n8365), .A2(n5606), .ZN(n5605) );
  NOR2_X1 U6242 ( .A1(n8893), .A2(n5439), .ZN(n8895) );
  NAND2_X1 U6243 ( .A1(n5441), .A2(n5440), .ZN(n5439) );
  OAI21_X1 U6244 ( .B1(n6658), .B2(n6596), .A(n9633), .ZN(n6625) );
  OAI21_X1 U6245 ( .B1(n10250), .B2(n10180), .A(n5338), .ZN(P1_U3265) );
  INV_X1 U6246 ( .A(n5339), .ZN(n5338) );
  OAI21_X1 U6247 ( .B1(n10251), .B2(n10220), .A(n5340), .ZN(n5339) );
  AOI21_X1 U6248 ( .B1(n10247), .B2(n11035), .A(n10054), .ZN(n5340) );
  AND2_X1 U6249 ( .A1(n5756), .A2(n5148), .ZN(n5110) );
  AND2_X1 U6250 ( .A1(n10190), .A2(n10209), .ZN(n5111) );
  OR2_X1 U6251 ( .A1(n7898), .A2(n9903), .ZN(n5112) );
  AND3_X1 U6252 ( .A1(n9663), .A2(n9662), .A3(n9661), .ZN(n5113) );
  AND4_X1 U6253 ( .A1(n6681), .A2(n6680), .A3(n7490), .A4(n6679), .ZN(n5114)
         );
  NAND4_X2 U6254 ( .A1(n7252), .A2(n7251), .A3(n7250), .A4(n7249), .ZN(n9069)
         );
  INV_X1 U6255 ( .A(n6243), .ZN(n5633) );
  AND2_X1 U6256 ( .A1(n5459), .A2(n6168), .ZN(n5115) );
  OR2_X1 U6257 ( .A1(n8900), .A2(n8897), .ZN(n5116) );
  INV_X1 U6258 ( .A(n9307), .ZN(n5533) );
  OR2_X1 U6259 ( .A1(n8259), .A2(n8271), .ZN(n9700) );
  NAND2_X1 U6260 ( .A1(n6355), .A2(n6354), .ZN(n10289) );
  INV_X1 U6261 ( .A(n10289), .ZN(n5355) );
  NAND2_X1 U6262 ( .A1(n6091), .A2(n6090), .ZN(n7864) );
  INV_X1 U6263 ( .A(n7864), .ZN(n5681) );
  OR2_X1 U6264 ( .A1(n10263), .A2(n10115), .ZN(n10076) );
  INV_X1 U6265 ( .A(n10076), .ZN(n5279) );
  OR2_X1 U6266 ( .A1(n9175), .A2(n8886), .ZN(n8732) );
  NAND2_X1 U6267 ( .A1(n6120), .A2(n6119), .ZN(n7898) );
  NOR2_X1 U6268 ( .A1(n9832), .A2(n9742), .ZN(n5117) );
  NAND2_X1 U6269 ( .A1(n6280), .A2(n6279), .ZN(n10234) );
  NAND2_X1 U6270 ( .A1(n5257), .A2(n5254), .ZN(n5118) );
  AND2_X1 U6271 ( .A1(n5241), .A2(n5240), .ZN(n5119) );
  AND2_X1 U6272 ( .A1(n5355), .A2(n10161), .ZN(n5120) );
  AND2_X1 U6273 ( .A1(n5275), .A2(n5274), .ZN(n5121) );
  NAND2_X1 U6274 ( .A1(n5169), .A2(n5319), .ZN(n5122) );
  INV_X1 U6275 ( .A(n6455), .ZN(n9582) );
  OR2_X1 U6276 ( .A1(n5519), .A2(n8803), .ZN(n5123) );
  AND2_X1 U6277 ( .A1(n6187), .A2(n6167), .ZN(n5124) );
  INV_X1 U6278 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5360) );
  INV_X1 U6279 ( .A(n6319), .ZN(n5643) );
  OR2_X1 U6280 ( .A1(n8896), .A2(n9180), .ZN(n5125) );
  NAND2_X1 U6281 ( .A1(n8026), .A2(n6167), .ZN(n8214) );
  INV_X1 U6282 ( .A(n5979), .ZN(n6013) );
  XNOR2_X1 U6283 ( .A(n6727), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7377) );
  NAND2_X1 U6284 ( .A1(n10202), .A2(n5212), .ZN(n10185) );
  NAND2_X1 U6285 ( .A1(n8616), .A2(n8615), .ZN(n8628) );
  OAI211_X1 U6286 ( .C1(n9730), .C2(n7234), .A(n5938), .B(n5937), .ZN(n7692)
         );
  OR2_X1 U6287 ( .A1(n10268), .A2(n10097), .ZN(n10004) );
  INV_X1 U6288 ( .A(n7231), .ZN(n7175) );
  AND2_X1 U6289 ( .A1(n9700), .A2(n9689), .ZN(n5330) );
  INV_X1 U6290 ( .A(n10158), .ZN(n5705) );
  OR2_X1 U6291 ( .A1(n6694), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n5128) );
  AND2_X1 U6292 ( .A1(n7899), .A2(n9672), .ZN(n5129) );
  NAND2_X1 U6293 ( .A1(n6150), .A2(n6149), .ZN(n8043) );
  NOR2_X1 U6294 ( .A1(n9044), .A2(n9042), .ZN(n5130) );
  OR2_X1 U6295 ( .A1(n7804), .A2(n7922), .ZN(n5131) );
  AND2_X1 U6296 ( .A1(n9070), .A2(n5088), .ZN(n5132) );
  NAND2_X1 U6297 ( .A1(n9234), .A2(n8871), .ZN(n5133) );
  AND2_X1 U6298 ( .A1(n8825), .A2(n5758), .ZN(n5134) );
  AND2_X1 U6299 ( .A1(n6455), .A2(n5652), .ZN(n5135) );
  XNOR2_X1 U6300 ( .A(n8332), .B(n8534), .ZN(n9112) );
  INV_X1 U6301 ( .A(n9784), .ZN(n5255) );
  INV_X1 U6302 ( .A(n7194), .ZN(n7248) );
  OAI211_X1 U6303 ( .C1(n9730), .C2(n7189), .A(n5836), .B(n5835), .ZN(n7334)
         );
  AND2_X1 U6304 ( .A1(n9751), .A2(n10005), .ZN(n10075) );
  INV_X1 U6305 ( .A(n10075), .ZN(n10073) );
  OR2_X1 U6306 ( .A1(n8525), .A2(n5434), .ZN(n5136) );
  AND2_X1 U6307 ( .A1(n5116), .A2(n8840), .ZN(n5137) );
  AND2_X1 U6308 ( .A1(n9392), .A2(n9059), .ZN(n5138) );
  INV_X1 U6309 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9510) );
  NAND2_X1 U6310 ( .A1(n6255), .A2(n6254), .ZN(n10303) );
  AND2_X1 U6311 ( .A1(n7512), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5139) );
  AND2_X1 U6312 ( .A1(n10835), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6313 ( .A1(n6206), .A2(n6205), .ZN(n10307) );
  AND2_X1 U6314 ( .A1(n8071), .A2(n9065), .ZN(n5141) );
  OR2_X1 U6315 ( .A1(n9069), .A2(n7602), .ZN(n5142) );
  NAND2_X1 U6316 ( .A1(n6685), .A2(n5552), .ZN(n6703) );
  NAND2_X1 U6317 ( .A1(n5740), .A2(n5744), .ZN(n8902) );
  XNOR2_X1 U6318 ( .A(n9307), .B(n8842), .ZN(n8936) );
  AND2_X1 U6319 ( .A1(n5125), .A2(n8875), .ZN(n5143) );
  NOR2_X1 U6320 ( .A1(n9111), .A2(n8333), .ZN(n5144) );
  NOR2_X1 U6321 ( .A1(n7543), .A2(n5656), .ZN(n5145) );
  INV_X1 U6322 ( .A(n7235), .ZN(n6893) );
  AND2_X1 U6323 ( .A1(n6726), .A2(n6721), .ZN(n7235) );
  INV_X1 U6324 ( .A(n6108), .ZN(n6111) );
  XNOR2_X1 U6325 ( .A(n6109), .B(n10414), .ZN(n6108) );
  INV_X1 U6326 ( .A(n6015), .ZN(n6016) );
  XNOR2_X1 U6327 ( .A(n6018), .B(SI_6_), .ZN(n6015) );
  AND2_X1 U6328 ( .A1(n10072), .A2(n5719), .ZN(n5146) );
  XNOR2_X1 U6329 ( .A(n6169), .B(n6142), .ZN(n6168) );
  AND2_X1 U6330 ( .A1(n9868), .A2(n9864), .ZN(n10014) );
  INV_X1 U6331 ( .A(n10014), .ZN(n5328) );
  AND2_X1 U6332 ( .A1(n9182), .A2(n9181), .ZN(n5147) );
  INV_X1 U6333 ( .A(n10254), .ZN(n10069) );
  NAND2_X1 U6334 ( .A1(n6547), .A2(n6546), .ZN(n10254) );
  NAND2_X1 U6335 ( .A1(n8829), .A2(n9288), .ZN(n5148) );
  AND2_X1 U6336 ( .A1(n5332), .A2(n10145), .ZN(n5149) );
  NOR2_X1 U6337 ( .A1(n5803), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6338 ( .A1(n9041), .A2(n8805), .ZN(n5151) );
  INV_X1 U6339 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10735) );
  AND2_X1 U6340 ( .A1(n11107), .A2(n9062), .ZN(n5152) );
  AND2_X1 U6341 ( .A1(n9301), .A2(n5534), .ZN(n5153) );
  INV_X1 U6342 ( .A(n9789), .ZN(n10242) );
  AND2_X1 U6343 ( .A1(n5278), .A2(n5280), .ZN(n5154) );
  NAND2_X1 U6344 ( .A1(n7405), .A2(n7381), .ZN(n5754) );
  NOR2_X1 U6345 ( .A1(n7976), .A2(n9065), .ZN(n5155) );
  NOR2_X1 U6346 ( .A1(n9295), .A2(n9304), .ZN(n5156) );
  NAND2_X1 U6347 ( .A1(n5819), .A2(n5772), .ZN(n5157) );
  INV_X1 U6348 ( .A(n5345), .ZN(n5344) );
  NAND2_X1 U6349 ( .A1(n5346), .A2(n10012), .ZN(n5345) );
  INV_X1 U6350 ( .A(n6645), .ZN(n5779) );
  AND2_X1 U6351 ( .A1(n6018), .A2(SI_6_), .ZN(n5158) );
  AND2_X1 U6352 ( .A1(n6169), .A2(SI_12_), .ZN(n5159) );
  NOR2_X1 U6353 ( .A1(n9710), .A2(n9747), .ZN(n5160) );
  INV_X1 U6354 ( .A(n5298), .ZN(n5297) );
  NOR2_X1 U6355 ( .A1(n5300), .A2(n5130), .ZN(n5298) );
  INV_X1 U6356 ( .A(n5766), .ZN(n5716) );
  INV_X1 U6357 ( .A(n5715), .ZN(n5714) );
  NAND2_X1 U6358 ( .A1(n5163), .A2(n5717), .ZN(n5715) );
  AND2_X1 U6359 ( .A1(n10047), .A2(n9774), .ZN(n10057) );
  INV_X1 U6360 ( .A(n10057), .ZN(n5284) );
  XNOR2_X1 U6361 ( .A(n6195), .B(SI_13_), .ZN(n6193) );
  AND2_X1 U6362 ( .A1(n10356), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5161) );
  INV_X1 U6363 ( .A(n5720), .ZN(n5719) );
  NAND2_X1 U6364 ( .A1(n5284), .A2(n10028), .ZN(n5720) );
  AND2_X1 U6365 ( .A1(n9746), .A2(n9745), .ZN(n9884) );
  AND2_X1 U6366 ( .A1(n10088), .A2(n10004), .ZN(n5162) );
  OR2_X1 U6367 ( .A1(n8220), .A2(n9901), .ZN(n5163) );
  INV_X1 U6368 ( .A(n5650), .ZN(n5649) );
  OAI21_X1 U6369 ( .B1(n9521), .B2(n5183), .A(n6455), .ZN(n5650) );
  OR2_X1 U6370 ( .A1(n8857), .A2(n9345), .ZN(n5164) );
  NAND2_X1 U6371 ( .A1(n8899), .A2(n8844), .ZN(n5165) );
  INV_X1 U6372 ( .A(n5744), .ZN(n5743) );
  NAND2_X1 U6373 ( .A1(n5165), .A2(n5116), .ZN(n5744) );
  OR2_X1 U6374 ( .A1(n5284), .A2(n5283), .ZN(n5166) );
  NAND2_X1 U6375 ( .A1(n9811), .A2(n5331), .ZN(n5167) );
  NAND2_X1 U6376 ( .A1(n9198), .A2(n5550), .ZN(n5168) );
  INV_X1 U6377 ( .A(n8527), .ZN(n5432) );
  AND2_X1 U6378 ( .A1(n5134), .A2(n8945), .ZN(n5169) );
  AND3_X1 U6379 ( .A1(n5645), .A2(n9581), .A3(n5644), .ZN(n5170) );
  AND2_X1 U6380 ( .A1(n5249), .A2(n6108), .ZN(n5171) );
  AND2_X1 U6381 ( .A1(n8869), .A2(n8868), .ZN(n5172) );
  AND2_X1 U6382 ( .A1(n5672), .A2(n10011), .ZN(n5173) );
  AND2_X1 U6383 ( .A1(n8889), .A2(n5463), .ZN(n5174) );
  AND2_X1 U6384 ( .A1(n9853), .A2(n9672), .ZN(n7865) );
  INV_X1 U6385 ( .A(n7865), .ZN(n5683) );
  NOR2_X1 U6386 ( .A1(n8301), .A2(n8300), .ZN(n5175) );
  NAND2_X1 U6387 ( .A1(n5675), .A2(n5674), .ZN(n10093) );
  INV_X1 U6388 ( .A(n10093), .ZN(n5337) );
  AND2_X1 U6389 ( .A1(n5741), .A2(n5738), .ZN(n5176) );
  AND2_X1 U6390 ( .A1(n9713), .A2(n5705), .ZN(n5177) );
  AND2_X1 U6391 ( .A1(n6688), .A2(n5760), .ZN(n5178) );
  NAND2_X1 U6392 ( .A1(n9750), .A2(n9779), .ZN(n10031) );
  INV_X1 U6393 ( .A(n10031), .ZN(n5269) );
  INV_X1 U6394 ( .A(n8728), .ZN(n9455) );
  NAND2_X1 U6395 ( .A1(n8691), .A2(n8690), .ZN(n8728) );
  INV_X1 U6396 ( .A(n5535), .ZN(n5534) );
  NAND2_X1 U6397 ( .A1(n5536), .A2(n8863), .ZN(n5535) );
  OR2_X1 U6398 ( .A1(n8518), .A2(n5518), .ZN(n5179) );
  INV_X1 U6399 ( .A(n7035), .ZN(n8842) );
  NAND2_X1 U6400 ( .A1(n8802), .A2(n8801), .ZN(n8908) );
  NAND2_X1 U6401 ( .A1(n8202), .A2(n8204), .ZN(n5634) );
  AND2_X1 U6402 ( .A1(n8159), .A2(n8280), .ZN(n5180) );
  AND2_X1 U6403 ( .A1(n8159), .A2(n5344), .ZN(n5181) );
  OR2_X1 U6404 ( .A1(n5698), .A2(n5696), .ZN(n5182) );
  XOR2_X1 U6405 ( .A(n6409), .B(n6636), .Z(n5183) );
  NAND2_X1 U6406 ( .A1(n6296), .A2(n6295), .ZN(n9610) );
  NOR2_X1 U6407 ( .A1(n9870), .A2(n5667), .ZN(n5666) );
  AND2_X1 U6408 ( .A1(n10051), .A2(n10967), .ZN(n5184) );
  AND2_X1 U6409 ( .A1(n10245), .A2(n10308), .ZN(n5185) );
  NAND2_X1 U6410 ( .A1(n5635), .A2(n5639), .ZN(n9529) );
  NOR3_X1 U6411 ( .A1(n10186), .A2(n10273), .A3(n5352), .ZN(n5350) );
  NOR2_X1 U6412 ( .A1(n8324), .A2(n8326), .ZN(n5186) );
  AND2_X1 U6413 ( .A1(n5479), .A2(n5478), .ZN(n5187) );
  INV_X1 U6414 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5695) );
  INV_X1 U6415 ( .A(n5351), .ZN(n10139) );
  NOR2_X1 U6416 ( .A1(n10186), .A2(n5352), .ZN(n5351) );
  NAND2_X1 U6417 ( .A1(n8877), .A2(n9058), .ZN(n5188) );
  NOR2_X1 U6418 ( .A1(n10192), .A2(n9747), .ZN(n5189) );
  NOR2_X1 U6419 ( .A1(n8814), .A2(n8813), .ZN(n5190) );
  NAND3_X1 U6420 ( .A1(n5634), .A2(n8203), .A3(n5633), .ZN(n5191) );
  AND2_X1 U6421 ( .A1(n10069), .A2(n10080), .ZN(n5192) );
  AND2_X1 U6422 ( .A1(SI_14_), .A2(keyinput_18), .ZN(n5193) );
  NAND2_X1 U6423 ( .A1(n6415), .A2(n6417), .ZN(n5194) );
  NAND2_X1 U6424 ( .A1(n5452), .A2(n6370), .ZN(n5195) );
  AND4_X1 U6425 ( .A1(n8695), .A2(n8404), .A3(n8403), .A4(n8402), .ZN(n9057)
         );
  INV_X1 U6426 ( .A(n9057), .ZN(n5438) );
  CLKBUF_X3 U6427 ( .A(n7376), .Z(n8392) );
  INV_X1 U6428 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5366) );
  INV_X1 U6429 ( .A(n8236), .ZN(n5591) );
  AND2_X1 U6430 ( .A1(n5311), .A2(n5309), .ZN(n5196) );
  INV_X1 U6431 ( .A(n7564), .ZN(n5541) );
  AND2_X1 U6432 ( .A1(n5753), .A2(n8925), .ZN(n5197) );
  INV_X1 U6433 ( .A(n11016), .ZN(n10972) );
  AND4_X1 U6434 ( .A1(n10566), .A2(n10565), .A3(n10564), .A4(n10563), .ZN(
        n5198) );
  INV_X1 U6435 ( .A(n8300), .ZN(n5488) );
  NOR2_X1 U6436 ( .A1(n7269), .A2(n7268), .ZN(n5199) );
  OAI21_X1 U6437 ( .B1(n7496), .B2(n5161), .A(n5609), .ZN(n5610) );
  AND2_X1 U6438 ( .A1(n8349), .A2(n5488), .ZN(n5200) );
  INV_X1 U6439 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5594) );
  XNOR2_X1 U6440 ( .A(n6678), .B(n6677), .ZN(n8451) );
  NOR2_X1 U6441 ( .A1(n7071), .A2(n7072), .ZN(n5201) );
  OR2_X1 U6442 ( .A1(n10524), .A2(n10525), .ZN(n5202) );
  OR2_X1 U6443 ( .A1(n10510), .A2(n10511), .ZN(n5203) );
  AND2_X1 U6444 ( .A1(n5489), .A2(n5493), .ZN(n5204) );
  AND2_X1 U6445 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(n10720), .ZN(n5205) );
  NAND2_X2 U6446 ( .A1(n8883), .A2(n10954), .ZN(n11119) );
  NOR2_X2 U6447 ( .A1(n9590), .A2(n5206), .ZN(n9548) );
  NAND2_X1 U6448 ( .A1(n8025), .A2(n5124), .ZN(n8215) );
  OAI21_X1 U6449 ( .B1(n7395), .B2(n7396), .A(n7397), .ZN(n6027) );
  AND2_X1 U6450 ( .A1(n5870), .A2(n5858), .ZN(n5865) );
  NAND2_X1 U6451 ( .A1(n6164), .A2(n6163), .ZN(n8025) );
  OAI21_X2 U6452 ( .B1(n9229), .B2(n9228), .A(n8721), .ZN(n9217) );
  NAND2_X1 U6453 ( .A1(n5800), .A2(n5804), .ZN(n5805) );
  XNOR2_X2 U6454 ( .A(n8882), .B(n8881), .ZN(n9379) );
  AOI21_X2 U6455 ( .B1(n5208), .B2(n5112), .A(n5207), .ZN(n8039) );
  OAI21_X2 U6456 ( .B1(n10074), .B2(n5720), .A(n5718), .ZN(n10041) );
  OAI22_X1 U6457 ( .A1(n10015), .A2(n10014), .B1(n10013), .B2(n10012), .ZN(
        n10225) );
  NAND2_X1 U6458 ( .A1(n6768), .A2(n6767), .ZN(n6770) );
  NAND2_X1 U6459 ( .A1(n7924), .A2(n8507), .ZN(n7952) );
  NAND2_X1 U6460 ( .A1(n7590), .A2(n8745), .ZN(n7569) );
  NOR2_X2 U6461 ( .A1(n9148), .A2(n8358), .ZN(n8337) );
  NAND2_X1 U6462 ( .A1(n8456), .A2(n8743), .ZN(n7407) );
  NAND2_X2 U6463 ( .A1(n5126), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6778) );
  NAND3_X1 U6464 ( .A1(n5150), .A2(n5722), .A3(n5786), .ZN(n5776) );
  NOR2_X1 U6465 ( .A1(n5687), .A2(n5686), .ZN(n5685) );
  INV_X1 U6466 ( .A(n8743), .ZN(n8468) );
  AND2_X1 U6467 ( .A1(n8463), .A2(n8461), .ZN(n8743) );
  NAND3_X1 U6468 ( .A1(n5436), .A2(n5435), .A3(n8747), .ZN(n7566) );
  XNOR2_X2 U6469 ( .A(n7354), .B(n8454), .ZN(n8741) );
  OAI21_X2 U6470 ( .B1(n7959), .B2(n7961), .A(n7960), .ZN(n8028) );
  NOR2_X1 U6471 ( .A1(n9592), .A2(n9591), .ZN(n9590) );
  NOR2_X1 U6472 ( .A1(n5638), .A2(n5636), .ZN(n9530) );
  INV_X1 U6473 ( .A(n5221), .ZN(n9926) );
  NAND2_X1 U6474 ( .A1(n5221), .A2(n5220), .ZN(n9945) );
  OR2_X1 U6475 ( .A1(n9921), .A2(n9922), .ZN(n5221) );
  NOR2_X1 U6476 ( .A1(n7057), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U6477 ( .A1(n5712), .A2(n5710), .ZN(n8261) );
  NOR2_X1 U6478 ( .A1(n7480), .A2(n7479), .ZN(n7880) );
  NAND2_X1 U6479 ( .A1(n5173), .A2(n5671), .ZN(n10316) );
  NAND2_X2 U6480 ( .A1(n6685), .A2(n5551), .ZN(n6765) );
  INV_X1 U6481 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5226) );
  INV_X1 U6482 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5224) );
  INV_X1 U6483 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5225) );
  NAND3_X1 U6484 ( .A1(n5226), .A2(n5225), .A3(n5224), .ZN(n5223) );
  NAND3_X1 U6485 ( .A1(n5228), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6486 ( .A1(n5981), .A2(n5229), .ZN(n5230) );
  NAND3_X1 U6487 ( .A1(n5239), .A2(n5238), .A3(n5236), .ZN(n5235) );
  NAND2_X1 U6488 ( .A1(n5246), .A2(n5249), .ZN(n6112) );
  NAND2_X1 U6489 ( .A1(n5246), .A2(n5171), .ZN(n5252) );
  INV_X1 U6490 ( .A(n9744), .ZN(n5267) );
  NAND3_X1 U6491 ( .A1(n9740), .A2(n9784), .A3(n10031), .ZN(n5258) );
  NAND2_X1 U6492 ( .A1(n5259), .A2(n5261), .ZN(n9829) );
  NAND2_X1 U6493 ( .A1(n5270), .A2(n5271), .ZN(n9727) );
  OR2_X1 U6494 ( .A1(n9722), .A2(n5272), .ZN(n5270) );
  OR2_X1 U6495 ( .A1(n9711), .A2(n5289), .ZN(n5285) );
  NAND2_X1 U6496 ( .A1(n5285), .A2(n5286), .ZN(n5292) );
  NAND2_X1 U6497 ( .A1(n5290), .A2(n5177), .ZN(n9716) );
  INV_X1 U6498 ( .A(n8249), .ZN(n5303) );
  NAND2_X1 U6499 ( .A1(n5307), .A2(n5312), .ZN(n5305) );
  NAND2_X1 U6500 ( .A1(n5311), .A2(n5313), .ZN(n7585) );
  NOR2_X1 U6501 ( .A1(n7586), .A2(n5310), .ZN(n5309) );
  NAND2_X1 U6502 ( .A1(n9022), .A2(n5317), .ZN(n5316) );
  NAND2_X1 U6503 ( .A1(n7008), .A2(n5855), .ZN(n5322) );
  NAND2_X1 U6504 ( .A1(n5322), .A2(n5871), .ZN(n5415) );
  XNOR2_X1 U6505 ( .A(n5322), .B(n5871), .ZN(n7041) );
  NAND2_X1 U6506 ( .A1(n8265), .A2(n5325), .ZN(n5327) );
  NAND2_X1 U6507 ( .A1(n8270), .A2(n5330), .ZN(n5326) );
  OAI21_X1 U6508 ( .B1(n8270), .B2(n8157), .A(n9689), .ZN(n8264) );
  NAND2_X1 U6509 ( .A1(n10175), .A2(n5334), .ZN(n5333) );
  NAND3_X1 U6510 ( .A1(n5348), .A2(n5347), .A3(n11030), .ZN(n11005) );
  INV_X1 U6511 ( .A(n5350), .ZN(n10123) );
  NAND2_X2 U6512 ( .A1(n5357), .A2(n5822), .ZN(n6787) );
  NAND2_X1 U6513 ( .A1(n5357), .A2(n5356), .ZN(n5359) );
  NAND2_X1 U6514 ( .A1(n6787), .A2(n10341), .ZN(n5358) );
  NAND2_X1 U6515 ( .A1(n10081), .A2(n5361), .ZN(n9987) );
  NAND2_X1 U6516 ( .A1(n10081), .A2(n5365), .ZN(n10042) );
  NAND2_X1 U6517 ( .A1(n10081), .A2(n10069), .ZN(n10063) );
  NAND4_X1 U6518 ( .A1(n5808), .A2(n10743), .A3(n10737), .A4(n5798), .ZN(n5803) );
  NAND3_X1 U6519 ( .A1(n10751), .A2(n10749), .A3(n10750), .ZN(n5413) );
  NAND2_X1 U6520 ( .A1(n5902), .A2(n5901), .ZN(n5414) );
  NAND3_X1 U6521 ( .A1(n8783), .A2(n8782), .A3(n5416), .ZN(n8796) );
  INV_X1 U6522 ( .A(n8699), .ZN(n5417) );
  NOR2_X1 U6523 ( .A1(n8698), .A2(n8773), .ZN(n5418) );
  AND2_X1 U6524 ( .A1(n5420), .A2(n7449), .ZN(n8448) );
  INV_X1 U6525 ( .A(n5421), .ZN(n6324) );
  NAND3_X1 U6526 ( .A1(n7407), .A2(n8462), .A3(n8461), .ZN(n5436) );
  NAND2_X1 U6527 ( .A1(n7426), .A2(n8742), .ZN(n7425) );
  NAND2_X1 U6528 ( .A1(n5442), .A2(n9057), .ZN(n8736) );
  NAND2_X1 U6529 ( .A1(n5442), .A2(n11121), .ZN(n9378) );
  NAND2_X1 U6530 ( .A1(n5442), .A2(n11106), .ZN(n5441) );
  NAND2_X1 U6531 ( .A1(n6685), .A2(n5443), .ZN(n5444) );
  OAI21_X1 U6532 ( .B1(n6349), .B2(n5449), .A(n5447), .ZN(n6423) );
  OAI21_X1 U6533 ( .B1(n6349), .B2(n6348), .A(n6347), .ZN(n6371) );
  NAND2_X1 U6534 ( .A1(n6112), .A2(n5455), .ZN(n5453) );
  NAND2_X1 U6535 ( .A1(n5453), .A2(n5454), .ZN(n6197) );
  NAND2_X1 U6536 ( .A1(n6112), .A2(n5461), .ZN(n5458) );
  AND2_X2 U6537 ( .A1(n5464), .A2(n5174), .ZN(n9382) );
  INV_X1 U6538 ( .A(n8888), .ZN(n5463) );
  OR2_X2 U6539 ( .A1(n9217), .A2(n9216), .ZN(n9394) );
  NAND2_X1 U6540 ( .A1(n6486), .A2(n5469), .ZN(n5467) );
  NAND2_X1 U6541 ( .A1(n6486), .A2(n5473), .ZN(n5468) );
  NAND2_X1 U6542 ( .A1(n6486), .A2(n6485), .ZN(n6506) );
  NAND2_X1 U6543 ( .A1(n8223), .A2(n5480), .ZN(n5476) );
  XNOR2_X1 U6544 ( .A(n8222), .B(n8236), .ZN(n8056) );
  NOR2_X1 U6545 ( .A1(n9159), .A2(n8299), .ZN(n8301) );
  OAI211_X1 U6546 ( .C1(n9159), .C2(n5485), .A(n5482), .B(n5481), .ZN(n8368)
         );
  OAI21_X1 U6547 ( .B1(n5487), .B2(n8349), .A(n5483), .ZN(n5482) );
  NAND2_X1 U6548 ( .A1(n5487), .A2(n5484), .ZN(n5483) );
  NAND2_X1 U6549 ( .A1(n5487), .A2(n5486), .ZN(n5485) );
  INV_X1 U6550 ( .A(n8349), .ZN(n5486) );
  INV_X1 U6551 ( .A(n6894), .ZN(n5492) );
  INV_X1 U6552 ( .A(n8293), .ZN(n5503) );
  OAI21_X1 U6553 ( .B1(n9078), .B2(n5503), .A(n5502), .ZN(n5505) );
  INV_X1 U6554 ( .A(n5505), .ZN(n9094) );
  NAND2_X1 U6555 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5507) );
  NAND3_X1 U6556 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U6557 ( .A1(n6861), .A2(n6860), .ZN(n6865) );
  NAND2_X1 U6558 ( .A1(n5608), .A2(n5602), .ZN(P2_U3201) );
  NAND2_X1 U6559 ( .A1(n6865), .A2(n6864), .ZN(n6892) );
  NAND2_X1 U6560 ( .A1(n7918), .A2(n5512), .ZN(n5510) );
  INV_X1 U6561 ( .A(n8116), .ZN(n5523) );
  OAI21_X1 U6562 ( .B1(n8116), .B2(n5179), .A(n5123), .ZN(n5515) );
  INV_X1 U6563 ( .A(n8115), .ZN(n5522) );
  OAI21_X1 U6564 ( .B1(n9302), .B2(n5535), .A(n5532), .ZN(n9278) );
  NAND2_X1 U6565 ( .A1(n7563), .A2(n5542), .ZN(n5540) );
  NAND2_X1 U6566 ( .A1(n5537), .A2(n5543), .ZN(n7822) );
  NAND3_X1 U6567 ( .A1(n5540), .A2(n5538), .A3(n5539), .ZN(n5537) );
  NAND3_X1 U6568 ( .A1(n5540), .A2(n5538), .A3(n7564), .ZN(n7735) );
  NAND2_X1 U6569 ( .A1(n9206), .A2(n5143), .ZN(n5545) );
  AOI21_X1 U6570 ( .B1(n9206), .B2(n5548), .A(n5546), .ZN(n8879) );
  OAI21_X1 U6571 ( .B1(n9206), .B2(n5138), .A(n8875), .ZN(n9192) );
  INV_X2 U6572 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5589) );
  XNOR2_X2 U6573 ( .A(n5592), .B(n5591), .ZN(n8052) );
  INV_X1 U6574 ( .A(n8240), .ZN(n5595) );
  NAND2_X1 U6575 ( .A1(n5598), .A2(n5186), .ZN(n5597) );
  INV_X1 U6576 ( .A(n5598), .ZN(n8325) );
  NAND2_X1 U6577 ( .A1(n6901), .A2(n6900), .ZN(n6903) );
  NAND2_X1 U6578 ( .A1(n5615), .A2(n7072), .ZN(n5613) );
  NAND4_X1 U6579 ( .A1(n5615), .A2(n6901), .A3(P2_REG2_REG_3__SCAN_IN), .A4(
        n6900), .ZN(n5614) );
  INV_X1 U6580 ( .A(n7074), .ZN(n5615) );
  NAND2_X1 U6581 ( .A1(n7268), .A2(n5618), .ZN(n5616) );
  NAND2_X1 U6582 ( .A1(n8202), .A2(n5630), .ZN(n5626) );
  NOR2_X2 U6583 ( .A1(n6296), .A2(n5641), .ZN(n5638) );
  NAND2_X1 U6584 ( .A1(n6410), .A2(n5647), .ZN(n5646) );
  OR2_X2 U6585 ( .A1(n6410), .A2(n5183), .ZN(n5653) );
  NOR2_X2 U6586 ( .A1(n5651), .A2(n9522), .ZN(n9583) );
  INV_X1 U6587 ( .A(n5653), .ZN(n9599) );
  NAND2_X1 U6588 ( .A1(n5655), .A2(n5654), .ZN(n7793) );
  NAND3_X1 U6589 ( .A1(n7289), .A2(n7291), .A3(n5657), .ZN(n6003) );
  NAND2_X1 U6590 ( .A1(n7308), .A2(n5657), .ZN(n7310) );
  NAND2_X1 U6591 ( .A1(n7289), .A2(n5657), .ZN(n7293) );
  AND2_X2 U6592 ( .A1(n5785), .A2(n5771), .ZN(n5793) );
  AND2_X2 U6593 ( .A1(n6203), .A2(n10365), .ZN(n5785) );
  NOR2_X2 U6594 ( .A1(n5698), .A2(n5697), .ZN(n6203) );
  NAND2_X1 U6595 ( .A1(n5927), .A2(n5926), .ZN(n5658) );
  NAND2_X1 U6596 ( .A1(n8035), .A2(n9795), .ZN(n8036) );
  NAND2_X1 U6597 ( .A1(n10130), .A2(n5676), .ZN(n5675) );
  INV_X1 U6598 ( .A(n5679), .ZN(n10112) );
  MUX2_X1 U6599 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5827), .Z(n5829) );
  NAND2_X1 U6600 ( .A1(n5685), .A2(n5689), .ZN(n7866) );
  OAI21_X2 U6601 ( .B1(n5684), .B2(n5682), .A(n5680), .ZN(n7897) );
  NAND2_X1 U6602 ( .A1(n5689), .A2(n5683), .ZN(n5682) );
  INV_X1 U6603 ( .A(n7713), .ZN(n5688) );
  AND2_X1 U6604 ( .A1(n5688), .A2(n5693), .ZN(n5686) );
  NAND2_X1 U6605 ( .A1(n7699), .A2(n5690), .ZN(n5689) );
  NAND4_X1 U6606 ( .A1(n5769), .A2(n5933), .A3(n5770), .A4(n5695), .ZN(n5697)
         );
  NAND2_X1 U6607 ( .A1(n6144), .A2(n5931), .ZN(n5698) );
  NAND3_X1 U6608 ( .A1(n6145), .A2(n5934), .A3(n5699), .ZN(n6171) );
  NAND2_X1 U6609 ( .A1(n8042), .A2(n5713), .ZN(n5712) );
  NAND2_X1 U6610 ( .A1(n10074), .A2(n10073), .ZN(n10072) );
  NAND2_X1 U6611 ( .A1(n5724), .A2(n7042), .ZN(n7191) );
  OAI21_X1 U6612 ( .B1(n7042), .B2(n5724), .A(n7191), .ZN(n7043) );
  NAND2_X2 U6613 ( .A1(n8789), .A2(n6834), .ZN(n7037) );
  NAND3_X1 U6614 ( .A1(n8789), .A2(n6834), .A3(n7038), .ZN(n7039) );
  NAND2_X2 U6615 ( .A1(n6765), .A2(n6708), .ZN(n8789) );
  AND2_X2 U6616 ( .A1(n6664), .A2(n6663), .ZN(n5725) );
  OAI22_X1 U6617 ( .A1(n7763), .A2(n5726), .B1(n5141), .B2(n5728), .ZN(n8075)
         );
  NAND2_X1 U6618 ( .A1(n8956), .A2(n5137), .ZN(n5740) );
  NAND2_X1 U6619 ( .A1(n8956), .A2(n8840), .ZN(n9031) );
  OAI211_X1 U6620 ( .C1(n8956), .C2(n5739), .A(n5735), .B(n5734), .ZN(n8854)
         );
  NAND2_X1 U6621 ( .A1(n8956), .A2(n5176), .ZN(n5734) );
  INV_X1 U6622 ( .A(n8849), .ZN(n5738) );
  INV_X1 U6623 ( .A(n8927), .ZN(n5750) );
  INV_X1 U6624 ( .A(n7245), .ZN(n5751) );
  NAND2_X1 U6625 ( .A1(n8926), .A2(n5754), .ZN(n5752) );
  NAND2_X1 U6626 ( .A1(n6690), .A2(n6686), .ZN(n6694) );
  NAND2_X1 U6627 ( .A1(n5779), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5860) );
  NAND4_X2 U6628 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5767), .ZN(n5886)
         );
  NAND2_X1 U6629 ( .A1(n8734), .A2(n8733), .ZN(n8735) );
  INV_X1 U6630 ( .A(n5995), .ZN(n5998) );
  AOI21_X1 U6631 ( .B1(n10057), .B2(n10055), .A(n5146), .ZN(n10256) );
  OR2_X2 U6632 ( .A1(n9548), .A2(n5764), .ZN(n6410) );
  NAND2_X1 U6633 ( .A1(n5147), .A2(n9387), .ZN(n9460) );
  OR2_X1 U6634 ( .A1(n9222), .A2(n9221), .ZN(n8874) );
  NAND4_X1 U6635 ( .A1(n7149), .A2(n7148), .A3(n7147), .A4(n7146), .ZN(n9072)
         );
  NAND2_X1 U6636 ( .A1(n7226), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7147) );
  AOI21_X2 U6637 ( .B1(n9564), .B2(n9565), .A(n5763), .ZN(n9574) );
  INV_X1 U6638 ( .A(n6724), .ZN(n6664) );
  AND2_X1 U6639 ( .A1(n5808), .A2(n10737), .ZN(n5761) );
  INV_X1 U6640 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5905) );
  AND2_X1 U6641 ( .A1(n10027), .A2(n10115), .ZN(n5762) );
  AND2_X1 U6642 ( .A1(n6270), .A2(n6269), .ZN(n5763) );
  AND2_X1 U6643 ( .A1(n6394), .A2(n6393), .ZN(n5764) );
  AND2_X1 U6644 ( .A1(n6085), .A2(n6065), .ZN(n5765) );
  AND2_X1 U6645 ( .A1(n11111), .A2(n11083), .ZN(n11104) );
  INV_X1 U6646 ( .A(n10835), .ZN(n6790) );
  INV_X1 U6647 ( .A(n7044), .ZN(n7226) );
  INV_X1 U6648 ( .A(n8220), .ZN(n11114) );
  AND2_X1 U6649 ( .A1(n8220), .A2(n9901), .ZN(n5766) );
  CLKBUF_X2 U6650 ( .A(P1_U3973), .Z(n9910) );
  INV_X1 U6651 ( .A(n10218), .ZN(n10180) );
  INV_X1 U6652 ( .A(n11028), .ZN(n10218) );
  OR2_X1 U6653 ( .A1(n5878), .A2(n5877), .ZN(n5767) );
  OAI221_X1 U6654 ( .B1(SI_30_), .B2(n10384), .C1(n10589), .C2(n10383), .A(
        n10382), .ZN(n10385) );
  INV_X1 U6655 ( .A(n10395), .ZN(n10396) );
  AND2_X1 U6656 ( .A1(n10402), .A2(n10401), .ZN(n10403) );
  NAND2_X1 U6657 ( .A1(n10404), .A2(n10403), .ZN(n10408) );
  INV_X1 U6658 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10485) );
  XNOR2_X1 U6659 ( .A(n10485), .B(keyinput_75), .ZN(n10486) );
  NAND2_X1 U6660 ( .A1(n10487), .A2(n10486), .ZN(n10488) );
  OR2_X1 U6661 ( .A1(n10489), .A2(n10488), .ZN(n10490) );
  XNOR2_X1 U6662 ( .A(n10500), .B(keyinput_86), .ZN(n10501) );
  AOI21_X1 U6663 ( .B1(n10503), .B2(n10502), .A(n10501), .ZN(n10504) );
  INV_X1 U6664 ( .A(n9785), .ZN(n9743) );
  NAND2_X1 U6665 ( .A1(n8451), .A2(n8785), .ZN(n7033) );
  NAND2_X1 U6666 ( .A1(n7186), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6869) );
  OR2_X1 U6667 ( .A1(n9572), .A2(n9571), .ZN(n6294) );
  INV_X1 U6668 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5798) );
  OR2_X1 U6669 ( .A1(n8847), .A2(n9033), .ZN(n8897) );
  INV_X1 U6670 ( .A(n10356), .ZN(n7512) );
  INV_X1 U6671 ( .A(n8399), .ZN(n8110) );
  AND2_X1 U6672 ( .A1(n6706), .A2(n6705), .ZN(n6707) );
  NAND2_X1 U6673 ( .A1(n9572), .A2(n9571), .ZN(n6295) );
  INV_X1 U6674 ( .A(n9884), .ZN(n9818) );
  INV_X1 U6675 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U6676 ( .A1(n5109), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5938) );
  INV_X1 U6677 ( .A(n10263), .ZN(n10027) );
  NAND2_X1 U6678 ( .A1(n5842), .A2(n5841), .ZN(n6949) );
  AND2_X1 U6679 ( .A1(n5761), .A2(n5798), .ZN(n5799) );
  INV_X1 U6680 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10365) );
  INV_X1 U6681 ( .A(SI_8_), .ZN(n10618) );
  NOR2_X1 U6682 ( .A1(n7552), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7551) );
  OR2_X1 U6683 ( .A1(n8800), .A2(n9007), .ZN(n8801) );
  AND2_X1 U6684 ( .A1(n8955), .A2(n8958), .ZN(n8840) );
  NAND2_X1 U6685 ( .A1(n8775), .A2(n8451), .ZN(n8776) );
  AND2_X1 U6686 ( .A1(n8330), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8331) );
  NOR2_X1 U6687 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7224) );
  AND2_X1 U6688 ( .A1(n9621), .A2(n9618), .ZN(n6532) );
  NAND2_X1 U6689 ( .A1(n6310), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6332) );
  AND2_X1 U6690 ( .A1(n6151), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6176) );
  OR2_X1 U6691 ( .A1(n6787), .A2(n7063), .ZN(n5835) );
  NAND2_X1 U6692 ( .A1(n10027), .A2(n10108), .ZN(n10100) );
  INV_X1 U6693 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10748) );
  INV_X1 U6694 ( .A(n6431), .ZN(n6429) );
  NAND2_X1 U6695 ( .A1(n6114), .A2(n6113), .ZN(n6139) );
  NAND2_X1 U6696 ( .A1(n7036), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5906) );
  AOI21_X1 U6697 ( .B1(n9031), .B2(n8899), .A(n8898), .ZN(n8901) );
  OR2_X1 U6698 ( .A1(n8582), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8599) );
  OR2_X1 U6699 ( .A1(n8839), .A2(n8986), .ZN(n8955) );
  NAND2_X1 U6700 ( .A1(n7649), .A2(n7022), .ZN(n7942) );
  OR2_X1 U6701 ( .A1(n8185), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8542) );
  INV_X1 U6702 ( .A(n9221), .ZN(n9228) );
  NAND2_X1 U6703 ( .A1(n8708), .A2(n9292), .ZN(n9307) );
  INV_X1 U6704 ( .A(n8785), .ZN(n7348) );
  INV_X1 U6705 ( .A(n9065), .ZN(n8081) );
  INV_X1 U6706 ( .A(n9066), .ZN(n7922) );
  AOI21_X1 U6707 ( .B1(n6735), .B2(n8104), .A(n8285), .ZN(n6974) );
  NOR2_X1 U6708 ( .A1(n6369), .A2(n6368), .ZN(n9550) );
  NAND2_X1 U6709 ( .A1(n9580), .A2(n6482), .ZN(n9557) );
  AND2_X1 U6710 ( .A1(n10035), .A2(n6608), .ZN(n10044) );
  NAND2_X1 U6711 ( .A1(n5100), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5880) );
  INV_X1 U6712 ( .A(n7063), .ZN(n6801) );
  NAND2_X1 U6713 ( .A1(n10076), .A2(n9723), .ZN(n10094) );
  AOI22_X1 U6714 ( .A1(n10225), .A2(n10226), .B1(n10234), .B2(n10016), .ZN(
        n10203) );
  AND2_X1 U6715 ( .A1(n6580), .A2(n6754), .ZN(n7524) );
  AND2_X1 U6716 ( .A1(n9826), .A2(n6952), .ZN(n11016) );
  AND2_X1 U6717 ( .A1(n7717), .A2(n7715), .ZN(n9668) );
  NAND2_X1 U6718 ( .A1(n6223), .A2(n6201), .ZN(n6224) );
  BUF_X8 U6719 ( .A(n5824), .Z(n7036) );
  AOI22_X1 U6720 ( .A1(n7242), .A2(n7241), .B1(n7413), .B2(n7240), .ZN(n8927)
         );
  INV_X1 U6721 ( .A(n11079), .ZN(n9053) );
  AND4_X1 U6722 ( .A1(n8587), .A2(n8586), .A3(n8585), .A4(n8584), .ZN(n9290)
         );
  AND4_X1 U6723 ( .A1(n8123), .A2(n8122), .A3(n8121), .A4(n8120), .ZN(n8803)
         );
  OR2_X1 U6724 ( .A1(n7044), .A2(n6847), .ZN(n7005) );
  AOI21_X1 U6725 ( .B1(n9162), .B2(n9161), .A(n10346), .ZN(n9163) );
  AND2_X1 U6726 ( .A1(n9193), .A2(n8679), .ZN(n9363) );
  INV_X1 U6727 ( .A(n9354), .ZN(n11106) );
  AND2_X1 U6728 ( .A1(n6643), .A2(n9633), .ZN(n6657) );
  AND2_X1 U6729 ( .A1(n6592), .A2(n5840), .ZN(n9893) );
  NOR2_X1 U6730 ( .A1(n7365), .A2(n7364), .ZN(n7477) );
  INV_X1 U6731 ( .A(n10021), .ZN(n10145) );
  AND2_X1 U6732 ( .A1(n9761), .A2(n9763), .ZN(n10191) );
  AND2_X1 U6733 ( .A1(n9693), .A2(n9687), .ZN(n9795) );
  INV_X1 U6734 ( .A(n11010), .ZN(n10967) );
  AND2_X1 U6735 ( .A1(n6578), .A2(n6756), .ZN(n7981) );
  INV_X1 U6736 ( .A(n11144), .ZN(n10885) );
  OR2_X1 U6737 ( .A1(n6788), .A2(n6661), .ZN(n6943) );
  AND2_X1 U6738 ( .A1(n6089), .A2(n6117), .ZN(n7478) );
  XNOR2_X1 U6739 ( .A(n5962), .B(n5930), .ZN(n5960) );
  INV_X1 U6740 ( .A(n7759), .ZN(n7823) );
  AND2_X1 U6741 ( .A1(n7001), .A2(n7000), .ZN(n11079) );
  OR2_X1 U6742 ( .A1(n7011), .A2(n7010), .ZN(n11072) );
  AOI21_X1 U6743 ( .B1(n9211), .B2(n9358), .A(n9210), .ZN(n9396) );
  AND2_X1 U6744 ( .A1(n9365), .A2(n9364), .ZN(n9442) );
  OR3_X1 U6745 ( .A1(n9431), .A2(n9430), .A3(n9429), .ZN(n9491) );
  AOI21_X1 U6746 ( .B1(n6658), .B2(n6657), .A(n6656), .ZN(n6659) );
  INV_X1 U6747 ( .A(n9633), .ZN(n9616) );
  OAI21_X1 U6748 ( .B1(n9891), .B2(n9890), .A(n9889), .ZN(n9897) );
  AND2_X1 U6749 ( .A1(n7535), .A2(n10227), .ZN(n11028) );
  INV_X1 U6750 ( .A(n11147), .ZN(n11146) );
  INV_X1 U6751 ( .A(n11150), .ZN(n11148) );
  INV_X1 U6752 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10552) );
  INV_X1 U6753 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10721) );
  INV_X1 U6754 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5806) );
  NOR2_X1 U6755 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5819) );
  INV_X1 U6756 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5772) );
  XNOR2_X2 U6757 ( .A(n5773), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U6758 ( .A1(n5818), .A2(n5819), .ZN(n5774) );
  NAND2_X1 U6759 ( .A1(n5774), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5775) );
  INV_X1 U6760 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5778) );
  NAND2_X4 U6761 ( .A1(n5780), .A2(n5876), .ZN(n6645) );
  NAND2_X1 U6762 ( .A1(n5779), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6763 ( .A1(n5100), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U6764 ( .A1(n6125), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5781) );
  INV_X1 U6765 ( .A(n5786), .ZN(n6277) );
  AND2_X1 U6766 ( .A1(n10729), .A2(n10730), .ZN(n6302) );
  INV_X1 U6767 ( .A(n6302), .ZN(n5787) );
  INV_X1 U6768 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5789) );
  INV_X1 U6769 ( .A(n5793), .ZN(n5794) );
  NAND2_X1 U6770 ( .A1(n5794), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5795) );
  MUX2_X1 U6771 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5795), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5796) );
  OR2_X1 U6772 ( .A1(n5789), .A2(n10737), .ZN(n5811) );
  INV_X1 U6773 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10736) );
  NAND2_X1 U6774 ( .A1(n5797), .A2(n10736), .ZN(n6592) );
  AOI21_X1 U6775 ( .B1(n5800), .B2(n5799), .A(n5789), .ZN(n5801) );
  INV_X1 U6776 ( .A(n6573), .ZN(n5817) );
  INV_X1 U6777 ( .A(n5803), .ZN(n5804) );
  INV_X1 U6778 ( .A(n6576), .ZN(n5816) );
  INV_X1 U6779 ( .A(n5808), .ZN(n5809) );
  NAND2_X1 U6780 ( .A1(n5809), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5810) );
  AND2_X1 U6781 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  NAND2_X1 U6782 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  INV_X1 U6783 ( .A(n6574), .ZN(n5815) );
  INV_X1 U6784 ( .A(n5818), .ZN(n5821) );
  NAND2_X1 U6785 ( .A1(n5821), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6602) );
  INV_X1 U6786 ( .A(n5819), .ZN(n5820) );
  INV_X1 U6787 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6603) );
  NAND3_X1 U6788 ( .A1(n5821), .A2(P1_IR_REG_31__SCAN_IN), .A3(n6603), .ZN(
        n5822) );
  MUX2_X1 U6789 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5824), .Z(n5903) );
  INV_X1 U6790 ( .A(SI_2_), .ZN(n5823) );
  XNOR2_X1 U6791 ( .A(n5903), .B(n5823), .ZN(n5901) );
  INV_X1 U6792 ( .A(SI_1_), .ZN(n5825) );
  XNOR2_X1 U6793 ( .A(n5829), .B(n5825), .ZN(n5871) );
  AND2_X1 U6794 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U6795 ( .A1(n5824), .A2(n5826), .ZN(n5855) );
  AND2_X1 U6796 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U6797 ( .A1(n8684), .A2(n5828), .ZN(n7008) );
  NAND2_X1 U6798 ( .A1(n5829), .A2(SI_1_), .ZN(n5830) );
  XNOR2_X1 U6799 ( .A(n5902), .B(n5901), .ZN(n7189) );
  NAND2_X1 U6800 ( .A1(n5109), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5836) );
  INV_X1 U6801 ( .A(n5831), .ZN(n5832) );
  NAND2_X1 U6802 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5832), .ZN(n5833) );
  MUX2_X1 U6803 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5833), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n5834) );
  INV_X1 U6804 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U6805 ( .A1(n10508), .A2(n5831), .ZN(n5909) );
  NAND2_X1 U6806 ( .A1(n5834), .A2(n5909), .ZN(n7063) );
  AND2_X1 U6807 ( .A1(n7334), .A2(n5867), .ZN(n5838) );
  NAND2_X1 U6808 ( .A1(n5839), .A2(n5867), .ZN(n5847) );
  NAND2_X1 U6809 ( .A1(n5840), .A2(n6592), .ZN(n6594) );
  INV_X1 U6810 ( .A(n6594), .ZN(n5842) );
  INV_X1 U6811 ( .A(n5841), .ZN(n6328) );
  NAND2_X1 U6812 ( .A1(n5913), .A2(n7334), .ZN(n5846) );
  NAND2_X1 U6813 ( .A1(n5847), .A2(n5846), .ZN(n5849) );
  BUF_X4 U6814 ( .A(n5848), .Z(n6636) );
  NAND2_X1 U6815 ( .A1(n5850), .A2(n5851), .ZN(n5894) );
  OAI21_X1 U6816 ( .B1(n5851), .B2(n5850), .A(n5894), .ZN(n5852) );
  INV_X1 U6817 ( .A(n5852), .ZN(n7333) );
  INV_X1 U6818 ( .A(SI_0_), .ZN(n5854) );
  INV_X1 U6819 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5853) );
  OAI21_X1 U6820 ( .B1(n8684), .B2(n5854), .A(n5853), .ZN(n5856) );
  AND2_X1 U6821 ( .A1(n5856), .A2(n5855), .ZN(n10341) );
  INV_X1 U6822 ( .A(n5857), .ZN(n6788) );
  NAND2_X1 U6823 ( .A1(n6788), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5858) );
  INV_X1 U6824 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U6825 ( .A1(n5100), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U6826 ( .A1(n6125), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5861) );
  INV_X1 U6827 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10825) );
  NAND2_X1 U6828 ( .A1(n6953), .A2(n5867), .ZN(n5864) );
  NAND2_X1 U6829 ( .A1(n5865), .A2(n5864), .ZN(n7048) );
  NAND2_X1 U6830 ( .A1(n6953), .A2(n5090), .ZN(n5869) );
  NOR2_X1 U6831 ( .A1(n5857), .A2(n5360), .ZN(n5866) );
  AOI21_X1 U6832 ( .B1(n6947), .B2(n5867), .A(n5866), .ZN(n5868) );
  NAND2_X1 U6833 ( .A1(n5869), .A2(n5868), .ZN(n7049) );
  NAND2_X1 U6834 ( .A1(n7048), .A2(n7049), .ZN(n5889) );
  NAND2_X1 U6835 ( .A1(n5870), .A2(n5992), .ZN(n5888) );
  NAND2_X1 U6836 ( .A1(n5889), .A2(n5888), .ZN(n5885) );
  NAND2_X1 U6837 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5872) );
  XNOR2_X2 U6838 ( .A(n5872), .B(P1_IR_REG_1__SCAN_IN), .ZN(n10835) );
  NAND2_X1 U6839 ( .A1(n7523), .A2(n5913), .ZN(n5883) );
  INV_X1 U6840 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U6841 ( .A1(n6125), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U6842 ( .A1(n5876), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U6843 ( .A1(n5886), .A2(n5867), .ZN(n5882) );
  NAND2_X1 U6844 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  XNOR2_X1 U6845 ( .A(n5884), .B(n6636), .ZN(n5890) );
  NAND2_X1 U6846 ( .A1(n5885), .A2(n5890), .ZN(n7157) );
  AND2_X1 U6847 ( .A1(n7523), .A2(n5867), .ZN(n5887) );
  AOI21_X1 U6848 ( .B1(n5886), .B2(n5101), .A(n5887), .ZN(n7159) );
  NAND2_X1 U6849 ( .A1(n7157), .A2(n7159), .ZN(n5893) );
  AND2_X1 U6850 ( .A1(n5889), .A2(n5888), .ZN(n5892) );
  INV_X1 U6851 ( .A(n5890), .ZN(n5891) );
  NAND2_X1 U6852 ( .A1(n5892), .A2(n5891), .ZN(n7158) );
  NAND2_X1 U6853 ( .A1(n5893), .A2(n7158), .ZN(n7330) );
  NAND2_X1 U6854 ( .A1(n7333), .A2(n7330), .ZN(n7331) );
  NAND2_X1 U6855 ( .A1(n7331), .A2(n5894), .ZN(n7210) );
  INV_X1 U6856 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10919) );
  NAND2_X1 U6857 ( .A1(n6125), .A2(n10919), .ZN(n5900) );
  INV_X1 U6858 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5895) );
  OR2_X1 U6859 ( .A1(n5954), .A2(n5895), .ZN(n5898) );
  INV_X1 U6860 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U6861 ( .A1(n9909), .A2(n5867), .ZN(n5915) );
  NAND2_X1 U6862 ( .A1(n5903), .A2(SI_2_), .ZN(n5904) );
  INV_X1 U6863 ( .A(SI_3_), .ZN(n5908) );
  XNOR2_X1 U6864 ( .A(n5928), .B(n5908), .ZN(n5926) );
  XNOR2_X1 U6865 ( .A(n5927), .B(n5926), .ZN(n7238) );
  NAND2_X1 U6866 ( .A1(n5109), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U6867 ( .A1(n5909), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5910) );
  XNOR2_X1 U6868 ( .A(n5910), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U6869 ( .A1(n6329), .A2(n6800), .ZN(n5911) );
  OAI211_X1 U6870 ( .C1(n9730), .C2(n7238), .A(n5912), .B(n5911), .ZN(n7617)
         );
  NAND2_X1 U6871 ( .A1(n7617), .A2(n6548), .ZN(n5914) );
  NAND2_X1 U6872 ( .A1(n5915), .A2(n5914), .ZN(n5916) );
  AND2_X1 U6873 ( .A1(n7617), .A2(n6528), .ZN(n5917) );
  AOI21_X1 U6874 ( .B1(n9909), .B2(n5101), .A(n5917), .ZN(n5944) );
  XNOR2_X1 U6875 ( .A(n5943), .B(n5944), .ZN(n7209) );
  NAND2_X1 U6876 ( .A1(n5100), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5920) );
  INV_X1 U6877 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5918) );
  XNOR2_X1 U6878 ( .A(n5918), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U6879 ( .A1(n6125), .A2(n7691), .ZN(n5919) );
  AND2_X1 U6880 ( .A1(n5920), .A2(n5919), .ZN(n5925) );
  INV_X1 U6881 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5921) );
  OR2_X1 U6882 ( .A1(n5954), .A2(n5921), .ZN(n5924) );
  INV_X1 U6883 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U6885 ( .A1(n10968), .A2(n5867), .ZN(n5940) );
  NAND2_X1 U6886 ( .A1(n5928), .A2(SI_3_), .ZN(n5929) );
  MUX2_X1 U6887 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7036), .Z(n5962) );
  INV_X1 U6888 ( .A(SI_4_), .ZN(n5930) );
  XNOR2_X1 U6889 ( .A(n5961), .B(n5960), .ZN(n7234) );
  NOR2_X1 U6890 ( .A1(n5934), .A2(n5789), .ZN(n5932) );
  MUX2_X1 U6891 ( .A(n5789), .B(n5932), .S(P1_IR_REG_4__SCAN_IN), .Z(n5936) );
  NAND2_X1 U6892 ( .A1(n5934), .A2(n5933), .ZN(n5984) );
  INV_X1 U6893 ( .A(n5984), .ZN(n5935) );
  NOR2_X1 U6894 ( .A1(n5936), .A2(n5935), .ZN(n10868) );
  NAND2_X1 U6895 ( .A1(n6329), .A2(n10868), .ZN(n5937) );
  NAND2_X1 U6896 ( .A1(n7692), .A2(n6548), .ZN(n5939) );
  NAND2_X1 U6897 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  AND2_X1 U6898 ( .A1(n7692), .A2(n6528), .ZN(n5942) );
  AOI21_X1 U6899 ( .B1(n10968), .B2(n5101), .A(n5942), .ZN(n5947) );
  XNOR2_X1 U6900 ( .A(n5949), .B(n5947), .ZN(n7301) );
  INV_X1 U6901 ( .A(n5943), .ZN(n5945) );
  NAND2_X1 U6902 ( .A1(n5945), .A2(n5944), .ZN(n7302) );
  NAND2_X1 U6903 ( .A1(n7211), .A2(n5946), .ZN(n7300) );
  INV_X1 U6904 ( .A(n5947), .ZN(n5948) );
  NAND2_X1 U6905 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  NAND2_X1 U6906 ( .A1(n7300), .A2(n5950), .ZN(n5995) );
  NAND2_X1 U6907 ( .A1(n6121), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5959) );
  AOI21_X1 U6908 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5952) );
  NOR2_X1 U6909 ( .A1(n5952), .A2(n5973), .ZN(n10976) );
  NAND2_X1 U6910 ( .A1(n5102), .A2(n10976), .ZN(n5958) );
  INV_X1 U6911 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5953) );
  OR2_X1 U6912 ( .A1(n6645), .A2(n5953), .ZN(n5957) );
  INV_X1 U6913 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5955) );
  OR2_X1 U6914 ( .A1(n6519), .A2(n5955), .ZN(n5956) );
  NAND4_X1 U6915 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n9908)
         );
  NAND2_X1 U6916 ( .A1(n9908), .A2(n6638), .ZN(n5970) );
  NAND2_X1 U6917 ( .A1(n5961), .A2(n5960), .ZN(n5964) );
  NAND2_X1 U6918 ( .A1(n5962), .A2(SI_4_), .ZN(n5963) );
  MUX2_X1 U6919 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n7036), .Z(n5982) );
  INV_X1 U6920 ( .A(SI_5_), .ZN(n5965) );
  XNOR2_X1 U6921 ( .A(n5981), .B(n5980), .ZN(n7380) );
  NAND2_X1 U6922 ( .A1(n5108), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U6923 ( .A1(n5984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5966) );
  XNOR2_X1 U6924 ( .A(n5966), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6932) );
  NAND2_X1 U6925 ( .A1(n6329), .A2(n6932), .ZN(n5967) );
  OAI211_X1 U6926 ( .C1(n9730), .C2(n7380), .A(n5968), .B(n5967), .ZN(n7634)
         );
  NAND2_X1 U6927 ( .A1(n7634), .A2(n6639), .ZN(n5969) );
  NAND2_X1 U6928 ( .A1(n5970), .A2(n5969), .ZN(n5971) );
  XNOR2_X1 U6929 ( .A(n5971), .B(n6636), .ZN(n5996) );
  NAND2_X1 U6930 ( .A1(n5995), .A2(n5996), .ZN(n7308) );
  AND2_X1 U6931 ( .A1(n7634), .A2(n6638), .ZN(n5972) );
  AOI21_X1 U6932 ( .B1(n9908), .B2(n5101), .A(n5972), .ZN(n7309) );
  NAND2_X1 U6933 ( .A1(n7308), .A2(n7309), .ZN(n7289) );
  NAND2_X1 U6934 ( .A1(n6121), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5978) );
  OAI21_X1 U6935 ( .B1(n5973), .B2(P1_REG3_REG_6__SCAN_IN), .A(n6005), .ZN(
        n7294) );
  INV_X1 U6936 ( .A(n7294), .ZN(n7782) );
  NAND2_X1 U6937 ( .A1(n5102), .A2(n7782), .ZN(n5977) );
  INV_X1 U6938 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6933) );
  OR2_X1 U6939 ( .A1(n6645), .A2(n6933), .ZN(n5976) );
  INV_X1 U6940 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5974) );
  OR2_X1 U6941 ( .A1(n6519), .A2(n5974), .ZN(n5975) );
  NAND4_X1 U6942 ( .A1(n5978), .A2(n5977), .A3(n5976), .A4(n5975), .ZN(n10970)
         );
  NAND2_X1 U6943 ( .A1(n10970), .A2(n6638), .ZN(n5991) );
  INV_X1 U6944 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6730) );
  INV_X1 U6945 ( .A(n9730), .ZN(n6143) );
  NAND2_X1 U6946 ( .A1(n5982), .A2(SI_5_), .ZN(n5983) );
  MUX2_X1 U6947 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7036), .Z(n6018) );
  XNOR2_X1 U6948 ( .A(n6017), .B(n6015), .ZN(n7558) );
  NAND2_X1 U6949 ( .A1(n6143), .A2(n7558), .ZN(n5989) );
  NAND2_X1 U6950 ( .A1(n6147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5985) );
  MUX2_X1 U6951 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5985), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5987) );
  NOR2_X1 U6952 ( .A1(n6147), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6045) );
  INV_X1 U6953 ( .A(n6045), .ZN(n5986) );
  NAND2_X1 U6954 ( .A1(n5987), .A2(n5986), .ZN(n6962) );
  INV_X1 U6955 ( .A(n6962), .ZN(n6966) );
  NAND2_X1 U6956 ( .A1(n6329), .A2(n6966), .ZN(n5988) );
  NAND2_X1 U6957 ( .A1(n7783), .A2(n6639), .ZN(n5990) );
  NAND2_X1 U6958 ( .A1(n5991), .A2(n5990), .ZN(n5993) );
  XNOR2_X1 U6959 ( .A(n5993), .B(n6561), .ZN(n5999) );
  AND2_X1 U6960 ( .A1(n7783), .A2(n6638), .ZN(n5994) );
  AOI21_X1 U6961 ( .B1(n10970), .B2(n5101), .A(n5994), .ZN(n6000) );
  NAND2_X1 U6962 ( .A1(n5999), .A2(n6000), .ZN(n7291) );
  INV_X1 U6963 ( .A(n5999), .ZN(n6002) );
  INV_X1 U6964 ( .A(n6000), .ZN(n6001) );
  NAND2_X1 U6965 ( .A1(n6002), .A2(n6001), .ZN(n7290) );
  NAND2_X1 U6966 ( .A1(n6003), .A2(n7290), .ZN(n7395) );
  NAND2_X1 U6967 ( .A1(n6121), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6012) );
  AND2_X1 U6968 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  NOR2_X1 U6969 ( .A1(n6028), .A2(n6006), .ZN(n11027) );
  NAND2_X1 U6970 ( .A1(n5102), .A2(n11027), .ZN(n6011) );
  INV_X1 U6971 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6007) );
  OR2_X1 U6972 ( .A1(n6645), .A2(n6007), .ZN(n6010) );
  INV_X1 U6973 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6008) );
  OR2_X1 U6974 ( .A1(n6519), .A2(n6008), .ZN(n6009) );
  NAND4_X1 U6975 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n9907)
         );
  NAND2_X1 U6976 ( .A1(n9907), .A2(n5101), .ZN(n6022) );
  OR2_X1 U6977 ( .A1(n6045), .A2(n5789), .ZN(n6014) );
  XNOR2_X1 U6978 ( .A(n6014), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7093) );
  AOI22_X1 U6979 ( .A1(n5979), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6329), .B2(
        n7093), .ZN(n6020) );
  MUX2_X1 U6980 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7036), .Z(n6039) );
  XNOR2_X1 U6981 ( .A(n6038), .B(n6036), .ZN(n7641) );
  NAND2_X1 U6982 ( .A1(n7641), .A2(n9644), .ZN(n6019) );
  NAND2_X1 U6983 ( .A1(n6020), .A2(n6019), .ZN(n7618) );
  NAND2_X1 U6984 ( .A1(n7618), .A2(n6528), .ZN(n6021) );
  NAND2_X1 U6985 ( .A1(n6022), .A2(n6021), .ZN(n7396) );
  NAND2_X1 U6986 ( .A1(n9907), .A2(n6638), .ZN(n6024) );
  NAND2_X1 U6987 ( .A1(n7618), .A2(n6639), .ZN(n6023) );
  NAND2_X1 U6988 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  XNOR2_X1 U6989 ( .A(n6025), .B(n6636), .ZN(n7397) );
  NAND2_X1 U6990 ( .A1(n7395), .A2(n7396), .ZN(n6026) );
  NAND2_X1 U6991 ( .A1(n6027), .A2(n6026), .ZN(n9536) );
  NAND2_X1 U6992 ( .A1(n6121), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U6993 ( .A1(n6028), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6071) );
  OR2_X1 U6994 ( .A1(n6028), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6029) );
  AND2_X1 U6995 ( .A1(n6071), .A2(n6029), .ZN(n9542) );
  NAND2_X1 U6996 ( .A1(n5102), .A2(n9542), .ZN(n6034) );
  INV_X1 U6997 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6030) );
  OR2_X1 U6998 ( .A1(n6645), .A2(n6030), .ZN(n6033) );
  INV_X1 U6999 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6031) );
  OR2_X1 U7000 ( .A1(n6519), .A2(n6031), .ZN(n6032) );
  NAND4_X1 U7001 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n9906)
         );
  NAND2_X1 U7002 ( .A1(n9906), .A2(n6638), .ZN(n6050) );
  NAND2_X1 U7003 ( .A1(n6038), .A2(n6037), .ZN(n6041) );
  NAND2_X1 U7004 ( .A1(n6039), .A2(SI_7_), .ZN(n6040) );
  INV_X1 U7005 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6752) );
  MUX2_X1 U7006 ( .A(n6752), .B(n6747), .S(n7036), .Z(n6042) );
  INV_X1 U7007 ( .A(n6042), .ZN(n6043) );
  NAND2_X1 U7008 ( .A1(n6043), .A2(SI_8_), .ZN(n6044) );
  XNOR2_X1 U7009 ( .A(n6061), .B(n6060), .ZN(n7764) );
  NAND2_X1 U7010 ( .A1(n7764), .A2(n9644), .ZN(n6048) );
  INV_X1 U7011 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10517) );
  NAND2_X1 U7012 ( .A1(n6045), .A2(n10517), .ZN(n6066) );
  NAND2_X1 U7013 ( .A1(n6066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6046) );
  XNOR2_X1 U7014 ( .A(n6046), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7317) );
  AOI22_X1 U7015 ( .A1(n5979), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6329), .B2(
        n7317), .ZN(n6047) );
  NAND2_X1 U7016 ( .A1(n9543), .A2(n6639), .ZN(n6049) );
  NAND2_X1 U7017 ( .A1(n6050), .A2(n6049), .ZN(n6051) );
  XNOR2_X1 U7018 ( .A(n6051), .B(n6561), .ZN(n9538) );
  NAND2_X1 U7019 ( .A1(n9906), .A2(n5101), .ZN(n6053) );
  NAND2_X1 U7020 ( .A1(n9543), .A2(n6638), .ZN(n6052) );
  AND2_X1 U7021 ( .A1(n6053), .A2(n6052), .ZN(n9537) );
  NAND2_X1 U7022 ( .A1(n9538), .A2(n9537), .ZN(n6054) );
  NAND2_X1 U7023 ( .A1(n9536), .A2(n6054), .ZN(n6058) );
  INV_X1 U7024 ( .A(n9538), .ZN(n6056) );
  INV_X1 U7025 ( .A(n9537), .ZN(n6055) );
  NAND2_X1 U7026 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  INV_X1 U7027 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6062) );
  MUX2_X1 U7028 ( .A(n6062), .B(n10552), .S(n7036), .Z(n6063) );
  INV_X1 U7029 ( .A(SI_9_), .ZN(n10619) );
  INV_X1 U7030 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7031 ( .A1(n6064), .A2(SI_9_), .ZN(n6065) );
  OR2_X1 U7032 ( .A1(n6066), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7033 ( .A1(n6067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6086) );
  XNOR2_X1 U7034 ( .A(n6086), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7363) );
  AOI22_X1 U7035 ( .A1(n5979), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6329), .B2(
        n7363), .ZN(n6068) );
  NAND2_X1 U7036 ( .A1(n7712), .A2(n6639), .ZN(n6079) );
  NAND2_X1 U7037 ( .A1(n6121), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6077) );
  INV_X1 U7038 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7039 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  AND2_X1 U7040 ( .A1(n6093), .A2(n6072), .ZN(n7614) );
  NAND2_X1 U7041 ( .A1(n5102), .A2(n7614), .ZN(n6076) );
  INV_X1 U7042 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7616) );
  OR2_X1 U7043 ( .A1(n6645), .A2(n7616), .ZN(n6075) );
  INV_X1 U7044 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6073) );
  OR2_X1 U7045 ( .A1(n6519), .A2(n6073), .ZN(n6074) );
  NAND4_X1 U7046 ( .A1(n6077), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n9905)
         );
  NAND2_X1 U7047 ( .A1(n9905), .A2(n6638), .ZN(n6078) );
  NAND2_X1 U7048 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  XNOR2_X1 U7049 ( .A(n6080), .B(n6561), .ZN(n6082) );
  AOI22_X1 U7050 ( .A1(n7712), .A2(n6638), .B1(n5101), .B2(n9905), .ZN(n6081)
         );
  XNOR2_X1 U7051 ( .A(n6082), .B(n6081), .ZN(n7543) );
  NAND2_X1 U7052 ( .A1(n6082), .A2(n6081), .ZN(n6083) );
  MUX2_X1 U7053 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7036), .Z(n6109) );
  XNOR2_X1 U7054 ( .A(n6112), .B(n6108), .ZN(n7936) );
  NAND2_X1 U7055 ( .A1(n7936), .A2(n9644), .ZN(n6091) );
  INV_X1 U7056 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10715) );
  NAND2_X1 U7057 ( .A1(n6086), .A2(n10715), .ZN(n6087) );
  NAND2_X1 U7058 ( .A1(n6087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6088) );
  INV_X1 U7059 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10714) );
  OR2_X1 U7060 ( .A1(n6088), .A2(n10714), .ZN(n6089) );
  NAND2_X1 U7061 ( .A1(n6088), .A2(n10714), .ZN(n6117) );
  AOI22_X1 U7062 ( .A1(n5979), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6329), .B2(
        n7478), .ZN(n6090) );
  NAND2_X1 U7063 ( .A1(n7864), .A2(n6639), .ZN(n6102) );
  NAND2_X1 U7064 ( .A1(n6121), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6100) );
  INV_X1 U7065 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7066 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  AND2_X1 U7067 ( .A1(n6123), .A2(n6094), .ZN(n7797) );
  NAND2_X1 U7068 ( .A1(n5102), .A2(n7797), .ZN(n6099) );
  INV_X1 U7069 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6095) );
  OR2_X1 U7070 ( .A1(n6645), .A2(n6095), .ZN(n6098) );
  INV_X1 U7071 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6096) );
  OR2_X1 U7072 ( .A1(n6519), .A2(n6096), .ZN(n6097) );
  NAND4_X1 U7073 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(n9904)
         );
  NAND2_X1 U7074 ( .A1(n9904), .A2(n6638), .ZN(n6101) );
  NAND2_X1 U7075 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  XNOR2_X1 U7076 ( .A(n6103), .B(n6561), .ZN(n6105) );
  AND2_X1 U7077 ( .A1(n9904), .A2(n5101), .ZN(n6104) );
  AOI21_X1 U7078 ( .B1(n7864), .B2(n6638), .A(n6104), .ZN(n7795) );
  NAND2_X1 U7079 ( .A1(n7793), .A2(n7795), .ZN(n6107) );
  NAND2_X1 U7080 ( .A1(n6107), .A2(n7794), .ZN(n7959) );
  NAND2_X1 U7081 ( .A1(n6109), .A2(SI_10_), .ZN(n6110) );
  INV_X1 U7082 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6916) );
  INV_X1 U7083 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6918) );
  MUX2_X1 U7084 ( .A(n6916), .B(n6918), .S(n7036), .Z(n6114) );
  INV_X1 U7085 ( .A(SI_11_), .ZN(n6113) );
  INV_X1 U7086 ( .A(n6114), .ZN(n6115) );
  NAND2_X1 U7087 ( .A1(n6115), .A2(SI_11_), .ZN(n6116) );
  XNOR2_X1 U7088 ( .A(n6141), .B(n6140), .ZN(n8002) );
  NAND2_X1 U7089 ( .A1(n8002), .A2(n9644), .ZN(n6120) );
  NAND2_X1 U7090 ( .A1(n6117), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6118) );
  XNOR2_X1 U7091 ( .A(n6118), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7881) );
  AOI22_X1 U7092 ( .A1(n5979), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6329), .B2(
        n7881), .ZN(n6119) );
  NAND2_X1 U7093 ( .A1(n7898), .A2(n6639), .ZN(n6132) );
  NAND2_X1 U7094 ( .A1(n6121), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6130) );
  INV_X1 U7095 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6122) );
  AND2_X1 U7096 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  NOR2_X1 U7097 ( .A1(n6151), .A2(n6124), .ZN(n7871) );
  NAND2_X1 U7098 ( .A1(n5102), .A2(n7871), .ZN(n6129) );
  INV_X1 U7099 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7872) );
  OR2_X1 U7100 ( .A1(n6645), .A2(n7872), .ZN(n6128) );
  INV_X1 U7101 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6126) );
  OR2_X1 U7102 ( .A1(n6519), .A2(n6126), .ZN(n6127) );
  NAND4_X1 U7103 ( .A1(n6130), .A2(n6129), .A3(n6128), .A4(n6127), .ZN(n9903)
         );
  NAND2_X1 U7104 ( .A1(n9903), .A2(n6528), .ZN(n6131) );
  NAND2_X1 U7105 ( .A1(n6132), .A2(n6131), .ZN(n6133) );
  XNOR2_X1 U7106 ( .A(n6133), .B(n6561), .ZN(n6135) );
  AND2_X1 U7107 ( .A1(n9903), .A2(n5101), .ZN(n6134) );
  AOI21_X1 U7108 ( .B1(n7898), .B2(n6638), .A(n6134), .ZN(n6136) );
  AND2_X1 U7109 ( .A1(n6135), .A2(n6136), .ZN(n7961) );
  INV_X1 U7110 ( .A(n6135), .ZN(n6138) );
  INV_X1 U7111 ( .A(n6136), .ZN(n6137) );
  NAND2_X1 U7112 ( .A1(n6138), .A2(n6137), .ZN(n7960) );
  INV_X1 U7113 ( .A(n8028), .ZN(n6164) );
  MUX2_X1 U7114 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7036), .Z(n6169) );
  INV_X1 U7115 ( .A(SI_12_), .ZN(n6142) );
  XNOR2_X1 U7116 ( .A(n6170), .B(n6168), .ZN(n8117) );
  NAND2_X1 U7117 ( .A1(n8117), .A2(n9644), .ZN(n6150) );
  INV_X1 U7118 ( .A(n6145), .ZN(n6146) );
  OAI21_X1 U7119 ( .B1(n6147), .B2(n6146), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6148) );
  XNOR2_X1 U7120 ( .A(n6148), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7886) );
  AOI22_X1 U7121 ( .A1(n5979), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6329), .B2(
        n7886), .ZN(n6149) );
  NAND2_X1 U7122 ( .A1(n8043), .A2(n6639), .ZN(n6160) );
  NAND2_X1 U7123 ( .A1(n6121), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6158) );
  NOR2_X1 U7124 ( .A1(n6151), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6152) );
  NOR2_X1 U7125 ( .A1(n6176), .A2(n6152), .ZN(n8030) );
  NAND2_X1 U7126 ( .A1(n5102), .A2(n8030), .ZN(n6157) );
  INV_X1 U7127 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6153) );
  OR2_X1 U7128 ( .A1(n6645), .A2(n6153), .ZN(n6156) );
  INV_X1 U7129 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6154) );
  OR2_X1 U7130 ( .A1(n6519), .A2(n6154), .ZN(n6155) );
  NAND4_X1 U7131 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n9902)
         );
  NAND2_X1 U7132 ( .A1(n9902), .A2(n6638), .ZN(n6159) );
  NAND2_X1 U7133 ( .A1(n6160), .A2(n6159), .ZN(n6161) );
  XNOR2_X1 U7134 ( .A(n6161), .B(n6561), .ZN(n6166) );
  AND2_X1 U7135 ( .A1(n9902), .A2(n5101), .ZN(n6162) );
  AOI21_X1 U7136 ( .B1(n8043), .B2(n6528), .A(n6162), .ZN(n6165) );
  XNOR2_X1 U7137 ( .A(n6166), .B(n6165), .ZN(n8029) );
  INV_X1 U7138 ( .A(n8029), .ZN(n6163) );
  NAND2_X1 U7139 ( .A1(n6166), .A2(n6165), .ZN(n6167) );
  MUX2_X1 U7140 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7036), .Z(n6195) );
  XNOR2_X1 U7141 ( .A(n6194), .B(n6193), .ZN(n8111) );
  NAND2_X1 U7142 ( .A1(n8111), .A2(n9644), .ZN(n6175) );
  NAND2_X1 U7143 ( .A1(n6171), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6172) );
  MUX2_X1 U7144 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6172), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6173) );
  AND2_X1 U7145 ( .A1(n6173), .A2(n5182), .ZN(n8093) );
  AOI22_X1 U7146 ( .A1(n5979), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6329), .B2(
        n8093), .ZN(n6174) );
  NAND2_X1 U7147 ( .A1(n8220), .A2(n6639), .ZN(n6184) );
  NAND2_X1 U7148 ( .A1(n6121), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6182) );
  NOR2_X1 U7149 ( .A1(n6176), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6177) );
  NOR2_X1 U7150 ( .A1(n6207), .A2(n6177), .ZN(n8211) );
  NAND2_X1 U7151 ( .A1(n5102), .A2(n8211), .ZN(n6181) );
  INV_X1 U7152 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n8045) );
  OR2_X1 U7153 ( .A1(n6645), .A2(n8045), .ZN(n6180) );
  INV_X1 U7154 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6178) );
  OR2_X1 U7155 ( .A1(n6519), .A2(n6178), .ZN(n6179) );
  NAND4_X1 U7156 ( .A1(n6182), .A2(n6181), .A3(n6180), .A4(n6179), .ZN(n9901)
         );
  NAND2_X1 U7157 ( .A1(n9901), .A2(n6528), .ZN(n6183) );
  NAND2_X1 U7158 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  XNOR2_X1 U7159 ( .A(n6185), .B(n6561), .ZN(n6188) );
  AND2_X1 U7160 ( .A1(n9901), .A2(n5101), .ZN(n6186) );
  AOI21_X1 U7161 ( .B1(n8220), .B2(n6638), .A(n6186), .ZN(n6189) );
  XNOR2_X1 U7162 ( .A(n6188), .B(n6189), .ZN(n8217) );
  INV_X1 U7163 ( .A(n8217), .ZN(n6187) );
  INV_X1 U7164 ( .A(n6188), .ZN(n6191) );
  INV_X1 U7165 ( .A(n6189), .ZN(n6190) );
  NAND2_X1 U7166 ( .A1(n6191), .A2(n6190), .ZN(n6192) );
  NAND2_X1 U7167 ( .A1(n6195), .A2(SI_13_), .ZN(n6196) );
  INV_X1 U7168 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7207) );
  INV_X1 U7169 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10557) );
  MUX2_X1 U7170 ( .A(n7207), .B(n10557), .S(n7036), .Z(n6199) );
  INV_X1 U7171 ( .A(n6199), .ZN(n6200) );
  NAND2_X1 U7172 ( .A1(n6200), .A2(SI_14_), .ZN(n6201) );
  XNOR2_X1 U7173 ( .A(n6225), .B(n6224), .ZN(n8179) );
  NAND2_X1 U7174 ( .A1(n8179), .A2(n9644), .ZN(n6206) );
  NAND2_X1 U7175 ( .A1(n5182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6202) );
  MUX2_X1 U7176 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6202), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6204) );
  INV_X1 U7177 ( .A(n6203), .ZN(n6226) );
  NAND2_X1 U7178 ( .A1(n6204), .A2(n6226), .ZN(n8103) );
  INV_X1 U7179 ( .A(n8103), .ZN(n8147) );
  AOI22_X1 U7180 ( .A1(n5979), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6329), .B2(
        n8147), .ZN(n6205) );
  NAND2_X1 U7181 ( .A1(n10307), .A2(n6639), .ZN(n6216) );
  NAND2_X1 U7182 ( .A1(n6121), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6214) );
  OR2_X1 U7183 ( .A1(n6207), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7184 ( .A1(n6207), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6231) );
  AND2_X1 U7185 ( .A1(n6208), .A2(n6231), .ZN(n8278) );
  NAND2_X1 U7186 ( .A1(n5102), .A2(n8278), .ZN(n6213) );
  INV_X1 U7187 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6209) );
  OR2_X1 U7188 ( .A1(n6645), .A2(n6209), .ZN(n6212) );
  INV_X1 U7189 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6210) );
  OR2_X1 U7190 ( .A1(n6519), .A2(n6210), .ZN(n6211) );
  NAND4_X1 U7191 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n9900)
         );
  NAND2_X1 U7192 ( .A1(n9900), .A2(n6638), .ZN(n6215) );
  NAND2_X1 U7193 ( .A1(n6216), .A2(n6215), .ZN(n6217) );
  XNOR2_X1 U7194 ( .A(n6217), .B(n6636), .ZN(n6220) );
  AND2_X1 U7195 ( .A1(n9900), .A2(n5101), .ZN(n6218) );
  AOI21_X1 U7196 ( .B1(n10307), .B2(n6638), .A(n6218), .ZN(n8204) );
  INV_X1 U7197 ( .A(n6219), .ZN(n6222) );
  INV_X1 U7198 ( .A(n6220), .ZN(n6221) );
  MUX2_X1 U7199 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7036), .Z(n6245) );
  XNOR2_X1 U7200 ( .A(n6245), .B(n10379), .ZN(n6244) );
  XNOR2_X1 U7201 ( .A(n6248), .B(n6244), .ZN(n8533) );
  NAND2_X1 U7202 ( .A1(n8533), .A2(n9644), .ZN(n6230) );
  NAND2_X1 U7203 ( .A1(n6226), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6227) );
  MUX2_X1 U7204 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6227), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6228) );
  NAND2_X1 U7205 ( .A1(n6228), .A2(n6277), .ZN(n8154) );
  INV_X1 U7206 ( .A(n8154), .ZN(n9911) );
  AOI22_X1 U7207 ( .A1(n5979), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6329), .B2(
        n9911), .ZN(n6229) );
  NAND2_X1 U7208 ( .A1(n8259), .A2(n6639), .ZN(n6241) );
  OAI21_X1 U7209 ( .B1(n6232), .B2(P1_REG3_REG_15__SCAN_IN), .A(n6256), .ZN(
        n9635) );
  INV_X1 U7210 ( .A(n9635), .ZN(n6233) );
  NAND2_X1 U7211 ( .A1(n5102), .A2(n6233), .ZN(n6239) );
  NAND2_X1 U7212 ( .A1(n6121), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6238) );
  INV_X1 U7213 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n6234) );
  OR2_X1 U7214 ( .A1(n6519), .A2(n6234), .ZN(n6237) );
  INV_X1 U7215 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6235) );
  OR2_X1 U7216 ( .A1(n6645), .A2(n6235), .ZN(n6236) );
  NAND4_X1 U7217 ( .A1(n6239), .A2(n6238), .A3(n6237), .A4(n6236), .ZN(n9899)
         );
  NAND2_X1 U7218 ( .A1(n9899), .A2(n6638), .ZN(n6240) );
  NAND2_X1 U7219 ( .A1(n6241), .A2(n6240), .ZN(n6242) );
  XNOR2_X1 U7220 ( .A(n6242), .B(n6561), .ZN(n6243) );
  INV_X1 U7221 ( .A(n8259), .ZN(n11134) );
  INV_X1 U7222 ( .A(n9899), .ZN(n8271) );
  OAI22_X1 U7223 ( .A1(n11134), .A2(n5091), .B1(n8271), .B2(n5105), .ZN(n9631)
         );
  INV_X1 U7224 ( .A(n6244), .ZN(n6247) );
  NAND2_X1 U7225 ( .A1(n6245), .A2(SI_15_), .ZN(n6246) );
  INV_X1 U7226 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7438) );
  INV_X1 U7227 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10558) );
  MUX2_X1 U7228 ( .A(n7438), .B(n10558), .S(n7036), .Z(n6250) );
  INV_X1 U7229 ( .A(n6250), .ZN(n6251) );
  NAND2_X1 U7230 ( .A1(n6251), .A2(SI_16_), .ZN(n6252) );
  XNOR2_X1 U7231 ( .A(n6273), .B(n6272), .ZN(n8537) );
  NAND2_X1 U7232 ( .A1(n8537), .A2(n9644), .ZN(n6255) );
  NAND2_X1 U7233 ( .A1(n6277), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6253) );
  XNOR2_X1 U7234 ( .A(n6253), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9932) );
  AOI22_X1 U7235 ( .A1(n5979), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6329), .B2(
        n9932), .ZN(n6254) );
  NAND2_X1 U7236 ( .A1(n10303), .A2(n6639), .ZN(n6266) );
  OAI21_X1 U7237 ( .B1(n6257), .B2(P1_REG3_REG_16__SCAN_IN), .A(n6283), .ZN(
        n6258) );
  INV_X1 U7238 ( .A(n6258), .ZN(n9566) );
  NAND2_X1 U7239 ( .A1(n5102), .A2(n9566), .ZN(n6264) );
  NAND2_X1 U7240 ( .A1(n6121), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6263) );
  INV_X1 U7241 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6259) );
  OR2_X1 U7242 ( .A1(n6645), .A2(n6259), .ZN(n6262) );
  INV_X1 U7243 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6260) );
  OR2_X1 U7244 ( .A1(n6519), .A2(n6260), .ZN(n6261) );
  NAND4_X1 U7245 ( .A1(n6264), .A2(n6263), .A3(n6262), .A4(n6261), .ZN(n10222)
         );
  NAND2_X1 U7246 ( .A1(n10222), .A2(n6638), .ZN(n6265) );
  NAND2_X1 U7247 ( .A1(n6266), .A2(n6265), .ZN(n6267) );
  XNOR2_X1 U7248 ( .A(n6267), .B(n6636), .ZN(n6268) );
  AOI22_X1 U7249 ( .A1(n10303), .A2(n6638), .B1(n5101), .B2(n10222), .ZN(n6269) );
  XNOR2_X1 U7250 ( .A(n6268), .B(n6269), .ZN(n9565) );
  INV_X1 U7251 ( .A(n6268), .ZN(n6270) );
  INV_X1 U7252 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7456) );
  INV_X1 U7253 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10555) );
  MUX2_X1 U7254 ( .A(n7456), .B(n10555), .S(n7036), .Z(n6274) );
  NAND2_X1 U7255 ( .A1(n6274), .A2(n10606), .ZN(n6299) );
  INV_X1 U7256 ( .A(n6274), .ZN(n6275) );
  NAND2_X1 U7257 ( .A1(n6275), .A2(SI_17_), .ZN(n6276) );
  XNOR2_X1 U7258 ( .A(n6298), .B(n6297), .ZN(n8552) );
  NAND2_X1 U7259 ( .A1(n8552), .A2(n9644), .ZN(n6280) );
  OR2_X1 U7260 ( .A1(n6277), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7261 ( .A1(n6278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6303) );
  XNOR2_X1 U7262 ( .A(n6303), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U7263 ( .A1(n5979), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6329), .B2(
        n9962), .ZN(n6279) );
  NAND2_X1 U7264 ( .A1(n10234), .A2(n6639), .ZN(n6290) );
  NAND2_X1 U7265 ( .A1(n6121), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6288) );
  INV_X1 U7266 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6282) );
  AOI21_X1 U7267 ( .B1(n6283), .B2(n6282), .A(n6310), .ZN(n9576) );
  NAND2_X1 U7268 ( .A1(n5102), .A2(n9576), .ZN(n6287) );
  INV_X1 U7269 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10229) );
  OR2_X1 U7270 ( .A1(n6645), .A2(n10229), .ZN(n6286) );
  INV_X1 U7271 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n6284) );
  OR2_X1 U7272 ( .A1(n6519), .A2(n6284), .ZN(n6285) );
  NAND4_X1 U7273 ( .A1(n6288), .A2(n6287), .A3(n6286), .A4(n6285), .ZN(n10016)
         );
  NAND2_X1 U7274 ( .A1(n10016), .A2(n6638), .ZN(n6289) );
  NAND2_X1 U7275 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  XNOR2_X1 U7276 ( .A(n6291), .B(n6636), .ZN(n9572) );
  NAND2_X1 U7277 ( .A1(n10234), .A2(n6638), .ZN(n6293) );
  NAND2_X1 U7278 ( .A1(n10016), .A2(n5101), .ZN(n6292) );
  NAND2_X1 U7279 ( .A1(n6293), .A2(n6292), .ZN(n9571) );
  MUX2_X1 U7280 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7036), .Z(n6321) );
  XNOR2_X1 U7281 ( .A(n6321), .B(n10583), .ZN(n6320) );
  XNOR2_X1 U7282 ( .A(n6324), .B(n6320), .ZN(n8564) );
  NAND2_X1 U7283 ( .A1(n8564), .A2(n9644), .ZN(n6309) );
  NAND2_X1 U7284 ( .A1(n6303), .A2(n10729), .ZN(n6300) );
  NAND2_X1 U7285 ( .A1(n6300), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6301) );
  OR2_X1 U7286 ( .A1(n6301), .A2(n10730), .ZN(n6307) );
  NAND2_X1 U7287 ( .A1(n6303), .A2(n6302), .ZN(n6305) );
  OR2_X1 U7288 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6304) );
  AND2_X1 U7289 ( .A1(n6305), .A2(n6304), .ZN(n6306) );
  AND2_X1 U7290 ( .A1(n6307), .A2(n6306), .ZN(n9975) );
  AOI22_X1 U7291 ( .A1(n5979), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6329), .B2(
        n9975), .ZN(n6308) );
  INV_X1 U7292 ( .A(n10299), .ZN(n10216) );
  NAND2_X1 U7293 ( .A1(n6121), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6317) );
  INV_X1 U7294 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6312) );
  AOI21_X1 U7295 ( .B1(n6312), .B2(n6311), .A(n6356), .ZN(n10213) );
  NAND2_X1 U7296 ( .A1(n5102), .A2(n10213), .ZN(n6316) );
  INV_X1 U7297 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9963) );
  OR2_X1 U7298 ( .A1(n6645), .A2(n9963), .ZN(n6315) );
  INV_X1 U7299 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n6313) );
  OR2_X1 U7300 ( .A1(n6519), .A2(n6313), .ZN(n6314) );
  NAND4_X1 U7301 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n10223)
         );
  INV_X1 U7302 ( .A(n10223), .ZN(n9709) );
  OAI22_X1 U7303 ( .A1(n10216), .A2(n5091), .B1(n9709), .B2(n5845), .ZN(n6319)
         );
  AOI22_X1 U7304 ( .A1(n10299), .A2(n6639), .B1(n6638), .B2(n10223), .ZN(n6318) );
  XOR2_X1 U7305 ( .A(n6636), .B(n6318), .Z(n9611) );
  INV_X1 U7306 ( .A(n6320), .ZN(n6323) );
  NAND2_X1 U7307 ( .A1(n6321), .A2(SI_18_), .ZN(n6322) );
  INV_X1 U7308 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7698) );
  INV_X1 U7309 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10695) );
  MUX2_X1 U7310 ( .A(n7698), .B(n10695), .S(n7036), .Z(n6325) );
  NAND2_X1 U7311 ( .A1(n6325), .A2(n10582), .ZN(n6347) );
  INV_X1 U7312 ( .A(n6325), .ZN(n6326) );
  NAND2_X1 U7313 ( .A1(n6326), .A2(SI_19_), .ZN(n6327) );
  NAND2_X1 U7314 ( .A1(n6347), .A2(n6327), .ZN(n6348) );
  XNOR2_X1 U7315 ( .A(n6349), .B(n6348), .ZN(n8577) );
  NAND2_X1 U7316 ( .A1(n8577), .A2(n9644), .ZN(n6331) );
  AOI22_X1 U7317 ( .A1(n5979), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6328), .B2(
        n6329), .ZN(n6330) );
  NAND2_X1 U7318 ( .A1(n10293), .A2(n6639), .ZN(n6340) );
  NAND2_X1 U7319 ( .A1(n6121), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6338) );
  XNOR2_X1 U7320 ( .A(P1_REG3_REG_19__SCAN_IN), .B(n6332), .ZN(n10188) );
  NAND2_X1 U7321 ( .A1(n5102), .A2(n10188), .ZN(n6337) );
  INV_X1 U7322 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6333) );
  OR2_X1 U7323 ( .A1(n6645), .A2(n6333), .ZN(n6336) );
  INV_X1 U7324 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n6334) );
  OR2_X1 U7325 ( .A1(n6519), .A2(n6334), .ZN(n6335) );
  NAND4_X1 U7326 ( .A1(n6338), .A2(n6337), .A3(n6336), .A4(n6335), .ZN(n10017)
         );
  NAND2_X1 U7327 ( .A1(n10017), .A2(n6638), .ZN(n6339) );
  NAND2_X1 U7328 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  XNOR2_X1 U7329 ( .A(n6341), .B(n6561), .ZN(n6344) );
  AND2_X1 U7330 ( .A1(n10017), .A2(n5101), .ZN(n6342) );
  AOI21_X1 U7331 ( .B1(n10293), .B2(n6638), .A(n6342), .ZN(n6343) );
  NAND2_X1 U7332 ( .A1(n6344), .A2(n6343), .ZN(n6345) );
  OAI21_X1 U7333 ( .B1(n6344), .B2(n6343), .A(n6345), .ZN(n9531) );
  INV_X1 U7334 ( .A(n6345), .ZN(n6346) );
  NOR2_X2 U7335 ( .A1(n9530), .A2(n6346), .ZN(n9592) );
  INV_X1 U7336 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7934) );
  INV_X1 U7337 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10694) );
  MUX2_X1 U7338 ( .A(n7934), .B(n10694), .S(n7036), .Z(n6351) );
  INV_X1 U7339 ( .A(SI_20_), .ZN(n6350) );
  NAND2_X1 U7340 ( .A1(n6351), .A2(n6350), .ZN(n6372) );
  INV_X1 U7341 ( .A(n6351), .ZN(n6352) );
  NAND2_X1 U7342 ( .A1(n6352), .A2(SI_20_), .ZN(n6353) );
  XNOR2_X1 U7343 ( .A(n6371), .B(n6370), .ZN(n8594) );
  NAND2_X1 U7344 ( .A1(n8594), .A2(n9644), .ZN(n6355) );
  NAND2_X1 U7345 ( .A1(n5979), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U7346 ( .A1(n6121), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6363) );
  NAND3_X1 U7347 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_REG3_REG_20__SCAN_IN), 
        .A3(n6356), .ZN(n6379) );
  INV_X1 U7348 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U7349 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(n6356), .ZN(n6357) );
  NAND2_X1 U7350 ( .A1(n9593), .A2(n6357), .ZN(n6358) );
  AND2_X1 U7351 ( .A1(n6379), .A2(n6358), .ZN(n9594) );
  NAND2_X1 U7352 ( .A1(n5102), .A2(n9594), .ZN(n6362) );
  INV_X1 U7353 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10173) );
  OR2_X1 U7354 ( .A1(n6645), .A2(n10173), .ZN(n6361) );
  INV_X1 U7355 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6359) );
  OR2_X1 U7356 ( .A1(n6519), .A2(n6359), .ZN(n6360) );
  NAND4_X1 U7357 ( .A1(n6363), .A2(n6362), .A3(n6361), .A4(n6360), .ZN(n10197)
         );
  AOI22_X1 U7358 ( .A1(n10289), .A2(n6639), .B1(n6638), .B2(n10197), .ZN(n6364) );
  XNOR2_X1 U7359 ( .A(n6364), .B(n6636), .ZN(n6366) );
  AND2_X1 U7360 ( .A1(n10197), .A2(n5101), .ZN(n6365) );
  AOI21_X1 U7361 ( .B1(n10289), .B2(n6638), .A(n6365), .ZN(n6367) );
  XNOR2_X1 U7362 ( .A(n6366), .B(n6367), .ZN(n9591) );
  INV_X1 U7363 ( .A(n6366), .ZN(n6369) );
  INV_X1 U7364 ( .A(n6367), .ZN(n6368) );
  MUX2_X1 U7365 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7036), .Z(n6395) );
  INV_X1 U7366 ( .A(SI_21_), .ZN(n6373) );
  XNOR2_X1 U7367 ( .A(n6395), .B(n6373), .ZN(n6415) );
  NAND2_X1 U7368 ( .A1(n8614), .A2(n9644), .ZN(n6376) );
  NAND2_X1 U7369 ( .A1(n5979), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U7370 ( .A1(n10284), .A2(n6639), .ZN(n6388) );
  INV_X1 U7371 ( .A(n6379), .ZN(n6377) );
  NAND2_X1 U7372 ( .A1(n6377), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6401) );
  INV_X1 U7373 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U7374 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  AND2_X1 U7375 ( .A1(n6401), .A2(n6380), .ZN(n10165) );
  NAND2_X1 U7376 ( .A1(n5102), .A2(n10165), .ZN(n6386) );
  NAND2_X1 U7377 ( .A1(n6121), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6385) );
  INV_X1 U7378 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6381) );
  OR2_X1 U7379 ( .A1(n6645), .A2(n6381), .ZN(n6384) );
  INV_X1 U7380 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n6382) );
  OR2_X1 U7381 ( .A1(n6519), .A2(n6382), .ZN(n6383) );
  NAND4_X1 U7382 ( .A1(n6386), .A2(n6385), .A3(n6384), .A4(n6383), .ZN(n10148)
         );
  NAND2_X1 U7383 ( .A1(n10148), .A2(n6638), .ZN(n6387) );
  NAND2_X1 U7384 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  XNOR2_X1 U7385 ( .A(n6389), .B(n6561), .ZN(n6391) );
  AND2_X1 U7386 ( .A1(n10148), .A2(n5101), .ZN(n6390) );
  AOI21_X1 U7387 ( .B1(n10284), .B2(n6638), .A(n6390), .ZN(n6392) );
  XNOR2_X1 U7388 ( .A(n6391), .B(n6392), .ZN(n9549) );
  INV_X1 U7389 ( .A(n6391), .ZN(n6394) );
  INV_X1 U7390 ( .A(n6392), .ZN(n6393) );
  NAND2_X1 U7391 ( .A1(n6416), .A2(n6415), .ZN(n6396) );
  NAND2_X1 U7392 ( .A1(n6395), .A2(SI_21_), .ZN(n6419) );
  MUX2_X1 U7393 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n7036), .Z(n6411) );
  XNOR2_X1 U7394 ( .A(n6411), .B(SI_22_), .ZN(n6412) );
  NAND2_X1 U7395 ( .A1(n8618), .A2(n9644), .ZN(n6399) );
  NAND2_X1 U7396 ( .A1(n5979), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6398) );
  INV_X1 U7397 ( .A(n6401), .ZN(n6400) );
  NAND2_X1 U7398 ( .A1(n6400), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6438) );
  INV_X1 U7399 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U7400 ( .A1(n6401), .A2(n9603), .ZN(n6402) );
  AND2_X1 U7401 ( .A1(n6438), .A2(n6402), .ZN(n10141) );
  NAND2_X1 U7402 ( .A1(n5102), .A2(n10141), .ZN(n6408) );
  NAND2_X1 U7403 ( .A1(n6121), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6407) );
  INV_X1 U7404 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6403) );
  OR2_X1 U7405 ( .A1(n6645), .A2(n6403), .ZN(n6406) );
  INV_X1 U7406 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6404) );
  OR2_X1 U7407 ( .A1(n5954), .A2(n6404), .ZN(n6405) );
  NAND4_X1 U7408 ( .A1(n6408), .A2(n6407), .A3(n6406), .A4(n6405), .ZN(n10132)
         );
  AOI22_X1 U7409 ( .A1(n10277), .A2(n6639), .B1(n6638), .B2(n10132), .ZN(n6409) );
  AOI22_X1 U7410 ( .A1(n10277), .A2(n6638), .B1(n5101), .B2(n10132), .ZN(n9602) );
  NAND2_X1 U7411 ( .A1(n6411), .A2(SI_22_), .ZN(n6418) );
  INV_X1 U7412 ( .A(n6418), .ZN(n6414) );
  INV_X1 U7413 ( .A(n6412), .ZN(n6413) );
  INV_X1 U7414 ( .A(n6417), .ZN(n6421) );
  AND2_X1 U7415 ( .A1(n6419), .A2(n6418), .ZN(n6420) );
  NAND2_X1 U7416 ( .A1(n6423), .A2(n6422), .ZN(n6432) );
  INV_X1 U7417 ( .A(n6432), .ZN(n6430) );
  INV_X1 U7418 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n6425) );
  INV_X1 U7419 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6424) );
  MUX2_X1 U7420 ( .A(n6425), .B(n6424), .S(n7036), .Z(n6426) );
  NAND2_X1 U7421 ( .A1(n6426), .A2(n10599), .ZN(n6456) );
  INV_X1 U7422 ( .A(n6426), .ZN(n6427) );
  NAND2_X1 U7423 ( .A1(n6427), .A2(SI_23_), .ZN(n6428) );
  NAND2_X1 U7424 ( .A1(n6456), .A2(n6428), .ZN(n6431) );
  NAND2_X1 U7425 ( .A1(n6430), .A2(n6429), .ZN(n6457) );
  NAND2_X1 U7426 ( .A1(n6432), .A2(n6431), .ZN(n6433) );
  NAND2_X1 U7427 ( .A1(n6457), .A2(n6433), .ZN(n8633) );
  NAND2_X1 U7428 ( .A1(n8633), .A2(n9644), .ZN(n6435) );
  NAND2_X1 U7429 ( .A1(n5979), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U7430 ( .A1(n10273), .A2(n6639), .ZN(n6447) );
  INV_X1 U7431 ( .A(n6438), .ZN(n6436) );
  NAND2_X1 U7432 ( .A1(n6436), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6465) );
  INV_X1 U7433 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U7434 ( .A1(n6438), .A2(n6437), .ZN(n6439) );
  AND2_X1 U7435 ( .A1(n6465), .A2(n6439), .ZN(n10124) );
  NAND2_X1 U7436 ( .A1(n5102), .A2(n10124), .ZN(n6445) );
  NAND2_X1 U7437 ( .A1(n6121), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6444) );
  INV_X1 U7438 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6440) );
  OR2_X1 U7439 ( .A1(n6645), .A2(n6440), .ZN(n6443) );
  INV_X1 U7440 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6441) );
  OR2_X1 U7441 ( .A1(n6519), .A2(n6441), .ZN(n6442) );
  NAND4_X1 U7442 ( .A1(n6445), .A2(n6444), .A3(n6443), .A4(n6442), .ZN(n10147)
         );
  NAND2_X1 U7443 ( .A1(n10147), .A2(n6638), .ZN(n6446) );
  NAND2_X1 U7444 ( .A1(n6447), .A2(n6446), .ZN(n6448) );
  XNOR2_X1 U7445 ( .A(n6448), .B(n6561), .ZN(n6450) );
  AND2_X1 U7446 ( .A1(n10147), .A2(n5101), .ZN(n6449) );
  AOI21_X1 U7447 ( .B1(n10273), .B2(n6638), .A(n6449), .ZN(n6451) );
  NAND2_X1 U7448 ( .A1(n6450), .A2(n6451), .ZN(n6455) );
  INV_X1 U7449 ( .A(n6450), .ZN(n6453) );
  INV_X1 U7450 ( .A(n6451), .ZN(n6452) );
  NAND2_X1 U7451 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  NAND2_X1 U7452 ( .A1(n6455), .A2(n6454), .ZN(n9521) );
  INV_X1 U7453 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8799) );
  INV_X1 U7454 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10688) );
  MUX2_X1 U7455 ( .A(n8799), .B(n10688), .S(n7036), .Z(n6458) );
  INV_X1 U7456 ( .A(SI_24_), .ZN(n10585) );
  NAND2_X1 U7457 ( .A1(n6458), .A2(n10585), .ZN(n6485) );
  INV_X1 U7458 ( .A(n6458), .ZN(n6459) );
  NAND2_X1 U7459 ( .A1(n6459), .A2(SI_24_), .ZN(n6460) );
  AND2_X1 U7460 ( .A1(n6485), .A2(n6460), .ZN(n6483) );
  NAND2_X1 U7461 ( .A1(n8636), .A2(n9644), .ZN(n6462) );
  NAND2_X1 U7462 ( .A1(n5979), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U7463 ( .A1(n10268), .A2(n6639), .ZN(n6474) );
  NAND2_X1 U7464 ( .A1(n6121), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6472) );
  INV_X1 U7465 ( .A(n6465), .ZN(n6463) );
  NAND2_X1 U7466 ( .A1(n6463), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6491) );
  INV_X1 U7467 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U7468 ( .A1(n6465), .A2(n6464), .ZN(n6466) );
  AND2_X1 U7469 ( .A1(n6491), .A2(n6466), .ZN(n10109) );
  NAND2_X1 U7470 ( .A1(n5102), .A2(n10109), .ZN(n6471) );
  INV_X1 U7471 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6467) );
  OR2_X1 U7472 ( .A1(n6645), .A2(n6467), .ZN(n6470) );
  INV_X1 U7473 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6468) );
  OR2_X1 U7474 ( .A1(n6519), .A2(n6468), .ZN(n6469) );
  NAND4_X1 U7475 ( .A1(n6472), .A2(n6471), .A3(n6470), .A4(n6469), .ZN(n10133)
         );
  NAND2_X1 U7476 ( .A1(n10133), .A2(n6638), .ZN(n6473) );
  NAND2_X1 U7477 ( .A1(n6474), .A2(n6473), .ZN(n6475) );
  XNOR2_X1 U7478 ( .A(n6475), .B(n6561), .ZN(n6477) );
  AND2_X1 U7479 ( .A1(n10133), .A2(n5101), .ZN(n6476) );
  AOI21_X1 U7480 ( .B1(n10268), .B2(n6638), .A(n6476), .ZN(n6478) );
  NAND2_X1 U7481 ( .A1(n6477), .A2(n6478), .ZN(n6482) );
  INV_X1 U7482 ( .A(n6477), .ZN(n6480) );
  INV_X1 U7483 ( .A(n6478), .ZN(n6479) );
  NAND2_X1 U7484 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  INV_X1 U7485 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8106) );
  INV_X1 U7486 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10687) );
  MUX2_X1 U7487 ( .A(n8106), .B(n10687), .S(n7036), .Z(n6502) );
  XNOR2_X1 U7488 ( .A(n6502), .B(SI_25_), .ZN(n6501) );
  NAND2_X1 U7489 ( .A1(n8436), .A2(n9644), .ZN(n6488) );
  NAND2_X1 U7490 ( .A1(n5979), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7491 ( .A1(n10263), .A2(n6639), .ZN(n6499) );
  NAND2_X1 U7492 ( .A1(n6121), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6497) );
  INV_X1 U7493 ( .A(n6491), .ZN(n6489) );
  NAND2_X1 U7494 ( .A1(n6489), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6515) );
  INV_X1 U7495 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U7496 ( .A1(n6491), .A2(n6490), .ZN(n6492) );
  AND2_X1 U7497 ( .A1(n6515), .A2(n6492), .ZN(n10090) );
  NAND2_X1 U7498 ( .A1(n5102), .A2(n10090), .ZN(n6496) );
  INV_X1 U7499 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10092) );
  OR2_X1 U7500 ( .A1(n6645), .A2(n10092), .ZN(n6495) );
  INV_X1 U7501 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6493) );
  OR2_X1 U7502 ( .A1(n5954), .A2(n6493), .ZN(n6494) );
  NAND4_X1 U7503 ( .A1(n6497), .A2(n6496), .A3(n6495), .A4(n6494), .ZN(n9898)
         );
  NAND2_X1 U7504 ( .A1(n9898), .A2(n6638), .ZN(n6498) );
  NAND2_X1 U7505 ( .A1(n6499), .A2(n6498), .ZN(n6500) );
  XNOR2_X1 U7506 ( .A(n6500), .B(n6636), .ZN(n6529) );
  AOI22_X1 U7507 ( .A1(n10263), .A2(n6638), .B1(n5101), .B2(n9898), .ZN(n6530)
         );
  XNOR2_X1 U7508 ( .A(n6529), .B(n6530), .ZN(n9558) );
  INV_X1 U7509 ( .A(n6501), .ZN(n6505) );
  INV_X1 U7510 ( .A(n6502), .ZN(n6503) );
  NAND2_X1 U7511 ( .A1(n6503), .A2(SI_25_), .ZN(n6504) );
  INV_X1 U7512 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6507) );
  INV_X1 U7513 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10685) );
  MUX2_X1 U7514 ( .A(n6507), .B(n10685), .S(n7036), .Z(n6508) );
  NAND2_X1 U7515 ( .A1(n6508), .A2(n10597), .ZN(n6536) );
  INV_X1 U7516 ( .A(n6508), .ZN(n6509) );
  NAND2_X1 U7517 ( .A1(n6509), .A2(SI_26_), .ZN(n6510) );
  NAND2_X1 U7518 ( .A1(n6536), .A2(n6510), .ZN(n6537) );
  NAND2_X1 U7519 ( .A1(n5979), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U7520 ( .A1(n10259), .A2(n6639), .ZN(n6525) );
  NAND2_X1 U7521 ( .A1(n6121), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6523) );
  INV_X1 U7522 ( .A(n6515), .ZN(n6513) );
  NAND2_X1 U7523 ( .A1(n6513), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6551) );
  INV_X1 U7524 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U7525 ( .A1(n6515), .A2(n6514), .ZN(n6516) );
  AND2_X1 U7526 ( .A1(n6551), .A2(n6516), .ZN(n10082) );
  NAND2_X1 U7527 ( .A1(n5102), .A2(n10082), .ZN(n6522) );
  INV_X1 U7528 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6517) );
  OR2_X1 U7529 ( .A1(n6645), .A2(n6517), .ZN(n6521) );
  INV_X1 U7530 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6518) );
  OR2_X1 U7531 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  NAND4_X1 U7532 ( .A1(n6523), .A2(n6522), .A3(n6521), .A4(n6520), .ZN(n10060)
         );
  NAND2_X1 U7533 ( .A1(n10060), .A2(n6638), .ZN(n6524) );
  NAND2_X1 U7534 ( .A1(n6525), .A2(n6524), .ZN(n6526) );
  XNOR2_X1 U7535 ( .A(n6526), .B(n6636), .ZN(n6535) );
  AND2_X1 U7536 ( .A1(n10060), .A2(n5101), .ZN(n6527) );
  AOI21_X1 U7537 ( .B1(n10259), .B2(n6638), .A(n6527), .ZN(n6533) );
  XNOR2_X1 U7538 ( .A(n6535), .B(n6533), .ZN(n9621) );
  INV_X1 U7539 ( .A(n6529), .ZN(n6531) );
  NAND2_X1 U7540 ( .A1(n6531), .A2(n6530), .ZN(n9618) );
  INV_X1 U7541 ( .A(n6533), .ZN(n6534) );
  NAND2_X1 U7542 ( .A1(n6535), .A2(n6534), .ZN(n6569) );
  INV_X1 U7543 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8383) );
  INV_X1 U7544 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10570) );
  MUX2_X1 U7545 ( .A(n8383), .B(n10570), .S(n7036), .Z(n6540) );
  INV_X1 U7546 ( .A(SI_27_), .ZN(n6539) );
  NAND2_X1 U7547 ( .A1(n6540), .A2(n6539), .ZN(n6626) );
  INV_X1 U7548 ( .A(n6540), .ZN(n6541) );
  NAND2_X1 U7549 ( .A1(n6541), .A2(SI_27_), .ZN(n6542) );
  AND2_X1 U7550 ( .A1(n6626), .A2(n6542), .ZN(n6543) );
  OR2_X1 U7551 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  NAND2_X1 U7552 ( .A1(n6627), .A2(n6545), .ZN(n8416) );
  NAND2_X1 U7553 ( .A1(n8416), .A2(n9644), .ZN(n6547) );
  NAND2_X1 U7554 ( .A1(n5979), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U7555 ( .A1(n10254), .A2(n6639), .ZN(n6560) );
  INV_X1 U7556 ( .A(n6551), .ZN(n6549) );
  NAND2_X1 U7557 ( .A1(n6549), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6607) );
  INV_X1 U7558 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U7559 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  NAND2_X1 U7560 ( .A1(n5102), .A2(n10066), .ZN(n6558) );
  NAND2_X1 U7561 ( .A1(n6121), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6557) );
  INV_X1 U7562 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6553) );
  OR2_X1 U7563 ( .A1(n6645), .A2(n6553), .ZN(n6556) );
  INV_X1 U7564 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6554) );
  OR2_X1 U7565 ( .A1(n6519), .A2(n6554), .ZN(n6555) );
  NAND4_X1 U7566 ( .A1(n6558), .A2(n6557), .A3(n6556), .A4(n6555), .ZN(n10051)
         );
  NAND2_X1 U7567 ( .A1(n10051), .A2(n6638), .ZN(n6559) );
  NAND2_X1 U7568 ( .A1(n6560), .A2(n6559), .ZN(n6562) );
  XNOR2_X1 U7569 ( .A(n6562), .B(n6561), .ZN(n6565) );
  INV_X1 U7570 ( .A(n6565), .ZN(n6567) );
  AND2_X1 U7571 ( .A1(n10051), .A2(n5101), .ZN(n6563) );
  AOI21_X1 U7572 ( .B1(n10254), .B2(n6638), .A(n6563), .ZN(n6564) );
  INV_X1 U7573 ( .A(n6564), .ZN(n6566) );
  AOI21_X1 U7574 ( .B1(n6567), .B2(n6566), .A(n6642), .ZN(n6568) );
  AOI21_X1 U7575 ( .B1(n9620), .B2(n6569), .A(n6568), .ZN(n6596) );
  INV_X1 U7576 ( .A(n6568), .ZN(n6571) );
  INV_X1 U7577 ( .A(n6569), .ZN(n6570) );
  NOR2_X1 U7578 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  AND2_X2 U7579 ( .A1(n9620), .A2(n6572), .ZN(n6658) );
  NAND2_X1 U7580 ( .A1(n6573), .A2(P1_B_REG_SCAN_IN), .ZN(n6575) );
  MUX2_X1 U7581 ( .A(P1_B_REG_SCAN_IN), .B(n6575), .S(n8140), .Z(n6577) );
  INV_X1 U7582 ( .A(n6576), .ZN(n6579) );
  NAND2_X1 U7583 ( .A1(n6577), .A2(n6579), .ZN(n6753) );
  OR2_X1 U7584 ( .A1(n6753), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6578) );
  OR2_X1 U7585 ( .A1(n6579), .A2(n5815), .ZN(n6756) );
  OR2_X1 U7586 ( .A1(n6753), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U7587 ( .A1(n6576), .A2(n6573), .ZN(n6754) );
  NOR4_X1 U7588 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6584) );
  NOR4_X1 U7589 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6583) );
  NOR4_X1 U7590 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6582) );
  NOR4_X1 U7591 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6581) );
  NAND4_X1 U7592 ( .A1(n6584), .A2(n6583), .A3(n6582), .A4(n6581), .ZN(n6590)
         );
  NOR2_X1 U7593 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n6588) );
  NOR4_X1 U7594 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6587) );
  NOR4_X1 U7595 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6586) );
  NOR4_X1 U7596 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6585) );
  NAND4_X1 U7597 ( .A1(n6588), .A2(n6587), .A3(n6586), .A4(n6585), .ZN(n6589)
         );
  NOR2_X1 U7598 ( .A1(n6590), .A2(n6589), .ZN(n6591) );
  OR2_X1 U7599 ( .A1(n6753), .A2(n6591), .ZN(n6945) );
  AND3_X1 U7600 ( .A1(n7981), .A2(n7524), .A3(n6945), .ZN(n6600) );
  NAND2_X1 U7601 ( .A1(n6592), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6593) );
  XNOR2_X1 U7602 ( .A(n6593), .B(n5366), .ZN(n7995) );
  NAND2_X1 U7603 ( .A1(n7995), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6661) );
  INV_X1 U7604 ( .A(n9835), .ZN(n9822) );
  AND2_X1 U7605 ( .A1(n6594), .A2(n9822), .ZN(n6598) );
  NAND2_X1 U7606 ( .A1(n6598), .A2(n6948), .ZN(n11141) );
  OR2_X1 U7607 ( .A1(n6594), .A2(n9822), .ZN(n7528) );
  NAND2_X1 U7608 ( .A1(n11141), .A2(n7528), .ZN(n6615) );
  NOR2_X1 U7609 ( .A1(n6943), .A2(n6615), .ZN(n6595) );
  INV_X1 U7610 ( .A(n6598), .ZN(n6958) );
  OR2_X1 U7611 ( .A1(n6958), .A2(n7908), .ZN(n7534) );
  NOR2_X1 U7612 ( .A1(n6943), .A2(n7534), .ZN(n6597) );
  NAND2_X1 U7613 ( .A1(n6600), .A2(n6597), .ZN(n6599) );
  NAND2_X1 U7614 ( .A1(n11006), .A2(n6328), .ZN(n6939) );
  NAND2_X1 U7615 ( .A1(n6599), .A2(n10227), .ZN(n9625) );
  NAND2_X1 U7616 ( .A1(n10254), .A2(n9625), .ZN(n6624) );
  INV_X1 U7617 ( .A(n6600), .ZN(n6617) );
  INV_X1 U7618 ( .A(n7528), .ZN(n9787) );
  INV_X1 U7619 ( .A(n6948), .ZN(n6601) );
  NAND2_X1 U7620 ( .A1(n9787), .A2(n6601), .ZN(n6950) );
  OR2_X1 U7621 ( .A1(n6943), .A2(n6950), .ZN(n9892) );
  NOR2_X1 U7622 ( .A1(n6617), .A2(n9892), .ZN(n6620) );
  NAND2_X1 U7623 ( .A1(n6602), .A2(n10748), .ZN(n6796) );
  NAND2_X1 U7624 ( .A1(n6796), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6604) );
  XNOR2_X1 U7625 ( .A(n6604), .B(n6603), .ZN(n10338) );
  NAND2_X1 U7626 ( .A1(n6121), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6614) );
  INV_X1 U7627 ( .A(n6607), .ZN(n6605) );
  NAND2_X1 U7628 ( .A1(n6605), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n10035) );
  INV_X1 U7629 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U7630 ( .A1(n6607), .A2(n6606), .ZN(n6608) );
  NAND2_X1 U7631 ( .A1(n5102), .A2(n10044), .ZN(n6613) );
  INV_X1 U7632 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6609) );
  OR2_X1 U7633 ( .A1(n6645), .A2(n6609), .ZN(n6612) );
  INV_X1 U7634 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6610) );
  OR2_X1 U7635 ( .A1(n5954), .A2(n6610), .ZN(n6611) );
  NAND4_X1 U7636 ( .A1(n6614), .A2(n6613), .A3(n6612), .A4(n6611), .ZN(n10059)
         );
  NAND3_X1 U7637 ( .A1(n9892), .A2(n6615), .A3(n7534), .ZN(n6616) );
  NAND2_X1 U7638 ( .A1(n6617), .A2(n6616), .ZN(n6619) );
  NAND2_X1 U7639 ( .A1(n9787), .A2(n6948), .ZN(n6941) );
  AND3_X1 U7640 ( .A1(n6941), .A2(n5857), .A3(n7995), .ZN(n6618) );
  NAND2_X1 U7641 ( .A1(n6619), .A2(n6618), .ZN(n7161) );
  AOI22_X1 U7642 ( .A1(n9640), .A2(n10059), .B1(n9624), .B2(n10066), .ZN(n6622) );
  INV_X1 U7643 ( .A(n10338), .ZN(n7053) );
  AOI22_X1 U7644 ( .A1(n9623), .A2(n10060), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6621) );
  AND2_X1 U7645 ( .A1(n6622), .A2(n6621), .ZN(n6623) );
  NAND3_X1 U7646 ( .A1(n6625), .A2(n6624), .A3(n6623), .ZN(P1_U3214) );
  INV_X1 U7647 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6628) );
  INV_X1 U7648 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10373) );
  MUX2_X1 U7649 ( .A(n6628), .B(n10373), .S(n7036), .Z(n6629) );
  NAND2_X1 U7650 ( .A1(n6629), .A2(n10591), .ZN(n8386) );
  INV_X1 U7651 ( .A(n6629), .ZN(n6630) );
  NAND2_X1 U7652 ( .A1(n6630), .A2(SI_28_), .ZN(n6631) );
  AND2_X1 U7653 ( .A1(n8386), .A2(n6631), .ZN(n8384) );
  NAND2_X1 U7654 ( .A1(n8406), .A2(n9644), .ZN(n6633) );
  NAND2_X1 U7655 ( .A1(n5979), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6632) );
  NAND2_X1 U7656 ( .A1(n10248), .A2(n6638), .ZN(n6635) );
  NAND2_X1 U7657 ( .A1(n10059), .A2(n5101), .ZN(n6634) );
  NAND2_X1 U7658 ( .A1(n6635), .A2(n6634), .ZN(n6637) );
  XNOR2_X1 U7659 ( .A(n6637), .B(n6636), .ZN(n6641) );
  AOI22_X1 U7660 ( .A1(n10248), .A2(n6639), .B1(n6638), .B2(n10059), .ZN(n6640) );
  XNOR2_X1 U7661 ( .A(n6641), .B(n6640), .ZN(n6643) );
  NAND3_X1 U7662 ( .A1(n6643), .A2(n9633), .A3(n6642), .ZN(n6655) );
  AOI22_X1 U7663 ( .A1(n9623), .A2(n10051), .B1(n9624), .B2(n10044), .ZN(n6652) );
  NAND2_X1 U7664 ( .A1(n6121), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6650) );
  INV_X1 U7665 ( .A(n10035), .ZN(n6644) );
  NAND2_X1 U7666 ( .A1(n5102), .A2(n6644), .ZN(n6649) );
  INV_X1 U7667 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n10036) );
  OR2_X1 U7668 ( .A1(n6645), .A2(n10036), .ZN(n6648) );
  INV_X1 U7669 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6646) );
  OR2_X1 U7670 ( .A1(n5954), .A2(n6646), .ZN(n6647) );
  NAND4_X1 U7671 ( .A1(n6650), .A2(n6649), .A3(n6648), .A4(n6647), .ZN(n10052)
         );
  AOI22_X1 U7672 ( .A1(n9640), .A2(n10052), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6651) );
  NAND2_X1 U7673 ( .A1(n6652), .A2(n6651), .ZN(n6653) );
  AOI21_X1 U7674 ( .B1(n10248), .B2(n9625), .A(n6653), .ZN(n6654) );
  NAND2_X1 U7675 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  NAND2_X1 U7676 ( .A1(n6660), .A2(n6659), .ZN(P1_U3220) );
  NOR2_X1 U7677 ( .A1(n6661), .A2(n5857), .ZN(P1_U3973) );
  INV_X1 U7678 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6666) );
  INV_X1 U7679 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6665) );
  NOR2_X1 U7680 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6669) );
  NOR2_X1 U7681 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6668) );
  NOR2_X1 U7682 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6667) );
  OAI21_X1 U7683 ( .B1(n7126), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7205) );
  NOR2_X1 U7684 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6672) );
  NOR2_X1 U7685 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6671) );
  INV_X1 U7686 ( .A(n6681), .ZN(n6673) );
  NAND2_X1 U7687 ( .A1(n6673), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6674) );
  NAND2_X1 U7688 ( .A1(n7205), .A2(n6674), .ZN(n7491) );
  NAND2_X1 U7689 ( .A1(n6992), .A2(n6679), .ZN(n6675) );
  NAND2_X1 U7690 ( .A1(n6675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6991) );
  INV_X1 U7691 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U7692 ( .A1(n6991), .A2(n6990), .ZN(n6676) );
  NAND2_X1 U7693 ( .A1(n6676), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6678) );
  INV_X1 U7694 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6677) );
  NOR3_X1 U7695 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n6680) );
  INV_X1 U7696 ( .A(n6685), .ZN(n6682) );
  NAND2_X1 U7697 ( .A1(n6682), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6683) );
  XNOR2_X1 U7698 ( .A(n6683), .B(n6684), .ZN(n7997) );
  INV_X1 U7699 ( .A(n7997), .ZN(n8791) );
  NAND2_X2 U7700 ( .A1(n8774), .A2(n8791), .ZN(n8670) );
  NOR2_X1 U7701 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n6686) );
  NAND2_X1 U7702 ( .A1(n5128), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6687) );
  MUX2_X1 U7703 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6687), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6689) );
  INV_X1 U7704 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6688) );
  NAND2_X1 U7705 ( .A1(n6689), .A2(n6703), .ZN(n8285) );
  INV_X1 U7706 ( .A(n8285), .ZN(n6698) );
  INV_X1 U7707 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U7708 ( .A1(n6700), .A2(n6699), .ZN(n6691) );
  NAND2_X1 U7709 ( .A1(n6691), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6693) );
  INV_X1 U7710 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6692) );
  XNOR2_X1 U7711 ( .A(n6693), .B(n6692), .ZN(n8797) );
  NAND2_X1 U7712 ( .A1(n6694), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6695) );
  MUX2_X1 U7713 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6695), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6696) );
  NAND2_X1 U7714 ( .A1(n6696), .A2(n5128), .ZN(n8104) );
  NOR2_X1 U7715 ( .A1(n8797), .A2(n8104), .ZN(n6697) );
  NAND2_X1 U7716 ( .A1(n6698), .A2(n6697), .ZN(n6997) );
  NAND2_X1 U7717 ( .A1(n8670), .A2(n6997), .ZN(n6701) );
  XNOR2_X1 U7718 ( .A(n6700), .B(n6699), .ZN(n7991) );
  NAND2_X1 U7719 ( .A1(n6701), .A2(n7991), .ZN(n6833) );
  NAND2_X1 U7720 ( .A1(n6703), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6702) );
  INV_X1 U7721 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6705) );
  INV_X1 U7722 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6706) );
  NAND2_X1 U7723 ( .A1(n6833), .A2(n8884), .ZN(n6709) );
  NAND2_X1 U7724 ( .A1(n6709), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X1 U7725 ( .A1(n7991), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6736) );
  INV_X1 U7726 ( .A(n6736), .ZN(n6710) );
  NOR2_X1 U7727 ( .A1(n6997), .A2(n6710), .ZN(P2_U3893) );
  AND2_X1 U7728 ( .A1(n7036), .A2(P1_U3086), .ZN(n7994) );
  INV_X2 U7729 ( .A(n7994), .ZN(n10340) );
  AND2_X1 U7730 ( .A1(n8684), .A2(P1_U3086), .ZN(n10331) );
  INV_X2 U7731 ( .A(n10331), .ZN(n10337) );
  INV_X1 U7732 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6781) );
  OAI222_X1 U7733 ( .A1(n6790), .A2(P1_U3086), .B1(n10340), .B2(n7041), .C1(
        n10337), .C2(n6781), .ZN(P1_U3354) );
  INV_X1 U7734 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6711) );
  OAI222_X1 U7735 ( .A1(n10337), .A2(n6711), .B1(n10340), .B2(n7189), .C1(
        P1_U3086), .C2(n7063), .ZN(P1_U3353) );
  NOR2_X1 U7736 ( .A1(n8684), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9513) );
  INV_X1 U7737 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6717) );
  INV_X1 U7738 ( .A(n6724), .ZN(n6715) );
  NOR2_X4 U7739 ( .A1(n6716), .A2(n6715), .ZN(n7186) );
  INV_X1 U7740 ( .A(n7186), .ZN(n6898) );
  OAI222_X1 U7741 ( .A1(n9516), .A2(n6717), .B1(n9518), .B2(n7189), .C1(
        P2_U3151), .C2(n6898), .ZN(P2_U3293) );
  INV_X1 U7742 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6718) );
  INV_X1 U7743 ( .A(n6800), .ZN(n6825) );
  OAI222_X1 U7744 ( .A1(n10337), .A2(n6718), .B1(n10340), .B2(n7238), .C1(
        P1_U3086), .C2(n6825), .ZN(P1_U3352) );
  INV_X1 U7745 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6719) );
  INV_X1 U7746 ( .A(n10868), .ZN(n6807) );
  OAI222_X1 U7747 ( .A1(n10337), .A2(n6719), .B1(n10340), .B2(n7234), .C1(
        P1_U3086), .C2(n6807), .ZN(P1_U3351) );
  INV_X1 U7748 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6720) );
  OAI222_X1 U7749 ( .A1(n9516), .A2(n6720), .B1(n9518), .B2(n7041), .C1(
        P2_U3151), .C2(n6851), .ZN(P2_U3294) );
  INV_X1 U7750 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U7751 ( .A1(n6721), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6722) );
  OAI222_X1 U7752 ( .A1(n9516), .A2(n6723), .B1(n9518), .B2(n7234), .C1(
        P2_U3151), .C2(n7175), .ZN(P2_U3291) );
  NAND2_X1 U7753 ( .A1(n6724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6725) );
  MUX2_X1 U7754 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6725), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6726) );
  OAI222_X1 U7755 ( .A1(n9516), .A2(n5905), .B1(n9518), .B2(n7238), .C1(
        P2_U3151), .C2(n6893), .ZN(P2_U3292) );
  INV_X1 U7756 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6728) );
  NAND2_X1 U7757 ( .A1(n6731), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6727) );
  INV_X1 U7758 ( .A(n7377), .ZN(n7178) );
  OAI222_X1 U7759 ( .A1(n9516), .A2(n6728), .B1(n9518), .B2(n7380), .C1(
        P2_U3151), .C2(n7178), .ZN(P2_U3290) );
  INV_X1 U7760 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6729) );
  INV_X1 U7761 ( .A(n6932), .ZN(n6814) );
  OAI222_X1 U7762 ( .A1(n10337), .A2(n6729), .B1(n10340), .B2(n7380), .C1(
        P1_U3086), .C2(n6814), .ZN(P1_U3350) );
  INV_X1 U7763 ( .A(n7558), .ZN(n6733) );
  OAI222_X1 U7764 ( .A1(n10337), .A2(n6730), .B1(n10340), .B2(n6733), .C1(
        P1_U3086), .C2(n6962), .ZN(P1_U3349) );
  INV_X1 U7765 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6734) );
  OR2_X1 U7766 ( .A1(n6739), .A2(n9510), .ZN(n6732) );
  XNOR2_X1 U7767 ( .A(n6732), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7502) );
  OAI222_X1 U7768 ( .A1(n9516), .A2(n6734), .B1(n9518), .B2(n6733), .C1(
        P2_U3151), .C2(n7561), .ZN(P2_U3289) );
  NAND2_X1 U7769 ( .A1(n6997), .A2(n6736), .ZN(n9508) );
  XNOR2_X1 U7770 ( .A(n8797), .B(P2_B_REG_SCAN_IN), .ZN(n6735) );
  OR2_X1 U7771 ( .A1(n9508), .A2(n6974), .ZN(n8288) );
  INV_X1 U7772 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U7773 ( .A1(n8285), .A2(n8797), .ZN(n6975) );
  INV_X1 U7774 ( .A(n6975), .ZN(n6737) );
  AOI22_X1 U7775 ( .A1(n8288), .A2(n6973), .B1(n6737), .B2(n6736), .ZN(
        P2_U3376) );
  INV_X1 U7776 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6744) );
  INV_X1 U7777 ( .A(n7641), .ZN(n6746) );
  INV_X1 U7778 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6738) );
  INV_X1 U7779 ( .A(n6761), .ZN(n6740) );
  NAND2_X1 U7780 ( .A1(n6740), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6742) );
  INV_X1 U7781 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6741) );
  NAND2_X1 U7782 ( .A1(n6742), .A2(n6741), .ZN(n6748) );
  OR2_X1 U7783 ( .A1(n6742), .A2(n6741), .ZN(n6743) );
  NAND2_X1 U7784 ( .A1(n6748), .A2(n6743), .ZN(n10356) );
  OAI222_X1 U7785 ( .A1(n9516), .A2(n6744), .B1(n9518), .B2(n6746), .C1(
        P2_U3151), .C2(n10356), .ZN(P2_U3288) );
  INV_X1 U7786 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10506) );
  INV_X1 U7787 ( .A(n7093), .ZN(n6745) );
  OAI222_X1 U7788 ( .A1(n10337), .A2(n10506), .B1(n10340), .B2(n6746), .C1(
        P1_U3086), .C2(n6745), .ZN(P1_U3348) );
  INV_X1 U7789 ( .A(n7764), .ZN(n6751) );
  INV_X1 U7790 ( .A(n7317), .ZN(n7323) );
  OAI222_X1 U7791 ( .A1(n10337), .A2(n6747), .B1(n10340), .B2(n6751), .C1(
        P1_U3086), .C2(n7323), .ZN(P1_U3347) );
  NAND2_X1 U7792 ( .A1(n6748), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6750) );
  INV_X1 U7793 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6749) );
  XNOR2_X1 U7794 ( .A(n6750), .B(n6749), .ZN(n7670) );
  OAI222_X1 U7795 ( .A1(n9516), .A2(n6752), .B1(n9518), .B2(n6751), .C1(
        P2_U3151), .C2(n7670), .ZN(P2_U3287) );
  INV_X1 U7796 ( .A(n6943), .ZN(n6758) );
  NAND2_X1 U7797 ( .A1(n6758), .A2(n6753), .ZN(n10343) );
  INV_X1 U7798 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10362) );
  INV_X1 U7799 ( .A(n6754), .ZN(n6755) );
  AOI22_X1 U7800 ( .A1(n10343), .A2(n10362), .B1(n6758), .B2(n6755), .ZN(
        P1_U3440) );
  INV_X1 U7801 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6759) );
  INV_X1 U7802 ( .A(n6756), .ZN(n6757) );
  AOI22_X1 U7803 ( .A1(n10343), .A2(n6759), .B1(n6758), .B2(n6757), .ZN(
        P1_U3439) );
  INV_X1 U7804 ( .A(n7807), .ZN(n6764) );
  NOR2_X1 U7805 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6760) );
  NAND2_X1 U7806 ( .A1(n6761), .A2(n6760), .ZN(n6782) );
  NAND2_X1 U7807 ( .A1(n6782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6762) );
  XNOR2_X1 U7808 ( .A(n6762), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7852) );
  AOI22_X1 U7809 ( .A1(n7852), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9513), .ZN(n6763) );
  OAI21_X1 U7810 ( .B1(n6764), .B2(n9518), .A(n6763), .ZN(P2_U3286) );
  INV_X1 U7811 ( .A(n7363), .ZN(n7367) );
  OAI222_X1 U7812 ( .A1(n10340), .A2(n6764), .B1(n7367), .B2(P1_U3086), .C1(
        n10552), .C2(n10337), .ZN(P1_U3346) );
  MUX2_X1 U7813 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6766), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6769) );
  INV_X1 U7814 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6767) );
  INV_X1 U7815 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6771) );
  AND2_X2 U7816 ( .A1(n6774), .A2(n6773), .ZN(n7223) );
  NAND2_X1 U7817 ( .A1(n7223), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6779) );
  INV_X1 U7818 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6775) );
  AND2_X2 U7819 ( .A1(n6773), .A2(n9519), .ZN(n7194) );
  NAND2_X1 U7820 ( .A1(n7194), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6776) );
  NAND4_X4 U7821 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n7354)
         );
  NAND2_X1 U7822 ( .A1(n7354), .A2(P2_U3893), .ZN(n6780) );
  OAI21_X1 U7823 ( .B1(P2_U3893), .B2(n6781), .A(n6780), .ZN(P2_U3492) );
  INV_X1 U7824 ( .A(n7936), .ZN(n6784) );
  INV_X1 U7825 ( .A(n7478), .ZN(n7483) );
  INV_X1 U7826 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10500) );
  OAI222_X1 U7827 ( .A1(n10340), .A2(n6784), .B1(n7483), .B2(P1_U3086), .C1(
        n10500), .C2(n10337), .ZN(P1_U3345) );
  INV_X1 U7828 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6785) );
  NOR2_X1 U7829 ( .A1(n6782), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6912) );
  OR2_X1 U7830 ( .A1(n6912), .A2(n9510), .ZN(n6783) );
  INV_X1 U7831 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6911) );
  XNOR2_X1 U7832 ( .A(n6783), .B(n6911), .ZN(n8054) );
  OAI222_X1 U7833 ( .A1(n9516), .A2(n6785), .B1(n9518), .B2(n6784), .C1(n8054), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  NAND2_X1 U7834 ( .A1(n7995), .A2(n9787), .ZN(n6786) );
  AND2_X1 U7835 ( .A1(n6787), .A2(n6786), .ZN(n6794) );
  INV_X1 U7836 ( .A(n6794), .ZN(n6789) );
  AOI21_X1 U7837 ( .B1(n6788), .B2(n7995), .A(P1_U3086), .ZN(n6795) );
  NOR2_X1 U7838 ( .A1(n10861), .A2(n9910), .ZN(P1_U3085) );
  INV_X1 U7839 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6791) );
  AOI22_X1 U7840 ( .A1(n10835), .A2(n6791), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n6790), .ZN(n10832) );
  NAND2_X1 U7841 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10833) );
  NOR2_X1 U7842 ( .A1(n10832), .A2(n10833), .ZN(n10831) );
  NAND2_X1 U7843 ( .A1(n6801), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6792) );
  OAI21_X1 U7844 ( .B1(n6801), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6792), .ZN(
        n7056) );
  AOI21_X1 U7845 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6801), .A(n7055), .ZN(
        n6819) );
  NAND2_X1 U7846 ( .A1(n6800), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6793) );
  OAI21_X1 U7847 ( .B1(n6800), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6793), .ZN(
        n6818) );
  NOR2_X1 U7848 ( .A1(n6819), .A2(n6818), .ZN(n6817) );
  XNOR2_X1 U7849 ( .A(n10868), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n10864) );
  NOR2_X1 U7850 ( .A1(n10865), .A2(n10864), .ZN(n10863) );
  AOI21_X1 U7851 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n10868), .A(n10863), .ZN(
        n6799) );
  AOI22_X1 U7852 ( .A1(n6932), .A2(n5953), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n6814), .ZN(n6798) );
  NOR2_X1 U7853 ( .A1(n6799), .A2(n6798), .ZN(n6931) );
  NAND2_X1 U7854 ( .A1(n6795), .A2(n6794), .ZN(n10830) );
  AND2_X1 U7855 ( .A1(n6797), .A2(n6796), .ZN(n9989) );
  INV_X1 U7856 ( .A(n9989), .ZN(n10823) );
  OR2_X1 U7857 ( .A1(n10823), .A2(n10338), .ZN(n10826) );
  NOR2_X1 U7858 ( .A1(n10830), .A2(n10826), .ZN(n10855) );
  AOI211_X1 U7859 ( .C1(n6799), .C2(n6798), .A(n6931), .B(n10862), .ZN(n6816)
         );
  OR2_X1 U7860 ( .A1(n10830), .A2(n7053), .ZN(n10849) );
  INV_X1 U7861 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U7862 ( .A1(n6800), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6806) );
  MUX2_X1 U7863 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10917), .S(n6800), .Z(n6821)
         );
  NAND2_X1 U7864 ( .A1(n6801), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6805) );
  INV_X1 U7865 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6802) );
  MUX2_X1 U7866 ( .A(n6802), .B(P1_REG1_REG_2__SCAN_IN), .S(n7063), .Z(n7060)
         );
  NAND2_X1 U7867 ( .A1(n10835), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6804) );
  INV_X1 U7868 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6803) );
  MUX2_X1 U7869 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6803), .S(n10835), .Z(n10838) );
  NAND3_X1 U7870 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(n10838), .ZN(n10837) );
  NAND2_X1 U7871 ( .A1(n6804), .A2(n10837), .ZN(n7059) );
  NAND2_X1 U7872 ( .A1(n7060), .A2(n7059), .ZN(n7058) );
  NAND2_X1 U7873 ( .A1(n6805), .A2(n7058), .ZN(n6822) );
  NAND2_X1 U7874 ( .A1(n6821), .A2(n6822), .ZN(n6820) );
  NAND2_X1 U7875 ( .A1(n6806), .A2(n6820), .ZN(n10873) );
  MUX2_X1 U7876 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6808), .S(n10868), .Z(n10872) );
  NAND2_X1 U7877 ( .A1(n10873), .A2(n10872), .ZN(n10870) );
  OAI21_X1 U7878 ( .B1(n6808), .B2(n6807), .A(n10870), .ZN(n6811) );
  INV_X1 U7879 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6809) );
  MUX2_X1 U7880 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6809), .S(n6932), .Z(n6810)
         );
  OR2_X1 U7881 ( .A1(n10830), .A2(n9989), .ZN(n10851) );
  INV_X1 U7882 ( .A(n10851), .ZN(n10871) );
  NAND2_X1 U7883 ( .A1(n6810), .A2(n6811), .ZN(n6925) );
  OAI211_X1 U7884 ( .C1(n6811), .C2(n6810), .A(n10871), .B(n6925), .ZN(n6813)
         );
  AND2_X1 U7885 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7312) );
  AOI21_X1 U7886 ( .B1(n10861), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n7312), .ZN(
        n6812) );
  OAI211_X1 U7887 ( .C1(n10849), .C2(n6814), .A(n6813), .B(n6812), .ZN(n6815)
         );
  OR2_X1 U7888 ( .A1(n6816), .A2(n6815), .ZN(P1_U3248) );
  AOI211_X1 U7889 ( .C1(n6819), .C2(n6818), .A(n6817), .B(n10862), .ZN(n6827)
         );
  OAI211_X1 U7890 ( .C1(n6822), .C2(n6821), .A(n10871), .B(n6820), .ZN(n6824)
         );
  AND2_X1 U7891 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7213) );
  AOI21_X1 U7892 ( .B1(n10861), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n7213), .ZN(
        n6823) );
  OAI211_X1 U7893 ( .C1(n10849), .C2(n6825), .A(n6824), .B(n6823), .ZN(n6826)
         );
  OR2_X1 U7894 ( .A1(n6827), .A2(n6826), .ZN(P1_U3246) );
  NAND2_X1 U7895 ( .A1(n6833), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6828) );
  INV_X2 U7896 ( .A(P2_U3893), .ZN(n9073) );
  INV_X1 U7897 ( .A(n8789), .ZN(n7014) );
  MUX2_X1 U7898 ( .A(n6828), .B(n9073), .S(n7014), .Z(n6829) );
  INV_X1 U7899 ( .A(n6829), .ZN(n6830) );
  NAND2_X1 U7900 ( .A1(n6830), .A2(n8884), .ZN(n10357) );
  INV_X1 U7901 ( .A(n7991), .ZN(n6831) );
  NOR2_X1 U7902 ( .A1(n6997), .A2(n6831), .ZN(n6832) );
  INV_X1 U7903 ( .A(n9158), .ZN(n10360) );
  INV_X1 U7904 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10649) );
  NOR2_X1 U7905 ( .A1(n8789), .A2(P2_U3151), .ZN(n8286) );
  NAND2_X1 U7906 ( .A1(n8286), .A2(n6833), .ZN(n6852) );
  OR2_X1 U7907 ( .A1(n6852), .A2(n8788), .ZN(n10346) );
  INV_X1 U7908 ( .A(n10346), .ZN(n9117) );
  AND2_X1 U7909 ( .A1(n5589), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U7910 ( .A1(n6712), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6862) );
  OAI21_X1 U7911 ( .B1(n6851), .B2(n6835), .A(n6862), .ZN(n6837) );
  INV_X1 U7912 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U7913 ( .A1(n6837), .A2(n6836), .ZN(n6838) );
  NAND2_X1 U7914 ( .A1(n6863), .A2(n6838), .ZN(n6839) );
  NAND2_X1 U7915 ( .A1(n9117), .A2(n6839), .ZN(n6845) );
  OR2_X1 U7916 ( .A1(n6852), .A2(n8381), .ZN(n10348) );
  INV_X1 U7917 ( .A(n10348), .ZN(n6873) );
  AND2_X1 U7918 ( .A1(n5589), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U7919 ( .A1(n6712), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6867) );
  OAI21_X1 U7920 ( .B1(n6851), .B2(n6840), .A(n6867), .ZN(n6841) );
  NAND2_X1 U7921 ( .A1(n6841), .A2(n6775), .ZN(n6842) );
  NAND2_X1 U7922 ( .A1(n6868), .A2(n6842), .ZN(n6843) );
  NAND2_X1 U7923 ( .A1(n6873), .A2(n6843), .ZN(n6844) );
  OAI211_X1 U7924 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10649), .A(n6845), .B(
        n6844), .ZN(n6846) );
  AOI21_X1 U7925 ( .B1(n10360), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n6846), .ZN(
        n6850) );
  MUX2_X1 U7926 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8381), .Z(n6879) );
  INV_X1 U7927 ( .A(n6851), .ZN(n7038) );
  XNOR2_X1 U7928 ( .A(n6879), .B(n7038), .ZN(n6848) );
  INV_X1 U7929 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6847) );
  INV_X1 U7930 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7139) );
  INV_X4 U7931 ( .A(n8788), .ZN(n8381) );
  MUX2_X1 U7932 ( .A(n6847), .B(n7139), .S(n8381), .Z(n6854) );
  NAND2_X1 U7933 ( .A1(n6854), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U7934 ( .A1(n6848), .A2(n6853), .ZN(n6880) );
  AND2_X1 U7935 ( .A1(P2_U3893), .A2(n8789), .ZN(n10352) );
  OAI211_X1 U7936 ( .C1(n6848), .C2(n6853), .A(n6880), .B(n10352), .ZN(n6849)
         );
  OAI211_X1 U7937 ( .C1(n10357), .C2(n6851), .A(n6850), .B(n6849), .ZN(
        P2_U3183) );
  INV_X1 U7938 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U7939 ( .A1(n9166), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6858) );
  INV_X1 U7940 ( .A(n10352), .ZN(n6909) );
  NAND2_X1 U7941 ( .A1(n6909), .A2(n6852), .ZN(n6856) );
  OAI21_X1 U7942 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6854), .A(n6853), .ZN(n6855) );
  AOI22_X1 U7943 ( .A1(n6856), .A2(n6855), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6857) );
  OAI211_X1 U7944 ( .C1(n9158), .C2(n6859), .A(n6858), .B(n6857), .ZN(P2_U3182) );
  INV_X1 U7945 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6877) );
  INV_X1 U7946 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U7947 ( .A1(n6863), .A2(n6862), .ZN(n6864) );
  OAI21_X1 U7948 ( .B1(n6865), .B2(n6864), .A(n6892), .ZN(n6866) );
  AOI22_X1 U7949 ( .A1(n9117), .A2(n6866), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n6876) );
  NAND2_X1 U7950 ( .A1(n6870), .A2(n6869), .ZN(n6872) );
  NOR2_X1 U7951 ( .A1(n6872), .A2(n6871), .ZN(n6874) );
  OAI21_X1 U7952 ( .B1(n6897), .B2(n6874), .A(n6873), .ZN(n6875) );
  OAI211_X1 U7953 ( .C1(n6877), .C2(n9158), .A(n6876), .B(n6875), .ZN(n6878)
         );
  AOI21_X1 U7954 ( .B1(n7186), .B2(n9166), .A(n6878), .ZN(n6885) );
  INV_X1 U7955 ( .A(n6879), .ZN(n6881) );
  OAI21_X1 U7956 ( .B1(n7038), .B2(n6881), .A(n6880), .ZN(n6883) );
  MUX2_X1 U7957 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8381), .Z(n6886) );
  XNOR2_X1 U7958 ( .A(n6886), .B(n7186), .ZN(n6882) );
  NAND2_X1 U7959 ( .A1(n6883), .A2(n6882), .ZN(n6887) );
  OAI211_X1 U7960 ( .C1(n6883), .C2(n6882), .A(n6887), .B(n10352), .ZN(n6884)
         );
  NAND2_X1 U7961 ( .A1(n6885), .A2(n6884), .ZN(P2_U3184) );
  MUX2_X1 U7962 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8381), .Z(n7066) );
  XOR2_X1 U7963 ( .A(n7235), .B(n7066), .Z(n6890) );
  INV_X1 U7964 ( .A(n6886), .ZN(n6888) );
  OAI21_X1 U7965 ( .B1(n7186), .B2(n6888), .A(n6887), .ZN(n6889) );
  NOR2_X1 U7966 ( .A1(n6889), .A2(n6890), .ZN(n7067) );
  AOI21_X1 U7967 ( .B1(n6890), .B2(n6889), .A(n7067), .ZN(n6910) );
  OR2_X1 U7968 ( .A1(n7186), .A2(n10898), .ZN(n6891) );
  NAND2_X1 U7969 ( .A1(n6892), .A2(n6891), .ZN(n6894) );
  INV_X1 U7970 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10934) );
  AOI21_X1 U7971 ( .B1(n6895), .B2(n10934), .A(n5204), .ZN(n6896) );
  NAND2_X1 U7972 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8928) );
  OAI21_X1 U7973 ( .B1(n10346), .B2(n6896), .A(n8928), .ZN(n6906) );
  NAND2_X1 U7974 ( .A1(n6899), .A2(n7235), .ZN(n6900) );
  INV_X1 U7975 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6902) );
  AOI21_X1 U7976 ( .B1(n6903), .B2(n6902), .A(n7071), .ZN(n6904) );
  NOR2_X1 U7977 ( .A1(n6904), .A2(n10348), .ZN(n6905) );
  AOI211_X1 U7978 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n10360), .A(n6906), .B(
        n6905), .ZN(n6908) );
  NAND2_X1 U7979 ( .A1(n9166), .A2(n7235), .ZN(n6907) );
  OAI211_X1 U7980 ( .C1(n6910), .C2(n6909), .A(n6908), .B(n6907), .ZN(P2_U3185) );
  INV_X1 U7981 ( .A(n8002), .ZN(n6917) );
  NAND2_X1 U7982 ( .A1(n6912), .A2(n6911), .ZN(n6913) );
  NAND2_X1 U7983 ( .A1(n6913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6914) );
  NAND2_X1 U7984 ( .A1(n6914), .A2(n6666), .ZN(n7086) );
  OR2_X1 U7985 ( .A1(n6914), .A2(n6666), .ZN(n6915) );
  AND2_X1 U7986 ( .A1(n7086), .A2(n6915), .ZN(n8236) );
  OAI222_X1 U7987 ( .A1(n9516), .A2(n6916), .B1(n9518), .B2(n6917), .C1(
        P2_U3151), .C2(n5591), .ZN(P2_U3284) );
  INV_X1 U7988 ( .A(n7881), .ZN(n7885) );
  OAI222_X1 U7989 ( .A1(n10337), .A2(n6918), .B1(n10340), .B2(n6917), .C1(
        P1_U3086), .C2(n7885), .ZN(P1_U3344) );
  INV_X1 U7990 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6924) );
  INV_X1 U7991 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6922) );
  NAND2_X1 U7992 ( .A1(n6121), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6921) );
  INV_X1 U7993 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6919) );
  OR2_X1 U7994 ( .A1(n5954), .A2(n6919), .ZN(n6920) );
  OAI211_X1 U7995 ( .C1(n6645), .C2(n6922), .A(n6921), .B(n6920), .ZN(n9991)
         );
  NAND2_X1 U7996 ( .A1(n9991), .A2(n9910), .ZN(n6923) );
  OAI21_X1 U7997 ( .B1(n9910), .B2(n6924), .A(n6923), .ZN(P1_U3585) );
  INV_X1 U7998 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11001) );
  MUX2_X1 U7999 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n11001), .S(n6962), .Z(n6928)
         );
  INV_X1 U8000 ( .A(n6925), .ZN(n6926) );
  AOI21_X1 U8001 ( .B1(n6932), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6926), .ZN(
        n6927) );
  OR2_X1 U8002 ( .A1(n6928), .A2(n6927), .ZN(n6961) );
  NAND2_X1 U8003 ( .A1(n6928), .A2(n6927), .ZN(n6929) );
  NAND3_X1 U8004 ( .A1(n10871), .A2(n6961), .A3(n6929), .ZN(n6938) );
  INV_X1 U8005 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6930) );
  NOR2_X1 U8006 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6930), .ZN(n7296) );
  MUX2_X1 U8007 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6933), .S(n6962), .Z(n6934)
         );
  NOR2_X1 U8008 ( .A1(n6935), .A2(n6934), .ZN(n6965) );
  AOI211_X1 U8009 ( .C1(n6935), .C2(n6934), .A(n6965), .B(n10862), .ZN(n6936)
         );
  AOI211_X1 U8010 ( .C1(n10861), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n7296), .B(
        n6936), .ZN(n6937) );
  OAI211_X1 U8011 ( .C1(n10849), .C2(n6962), .A(n6938), .B(n6937), .ZN(
        P1_U3249) );
  INV_X1 U8012 ( .A(n6939), .ZN(n6940) );
  NOR2_X1 U8013 ( .A1(n7524), .A2(n6940), .ZN(n6946) );
  INV_X1 U8014 ( .A(n6941), .ZN(n6942) );
  NOR2_X1 U8015 ( .A1(n6943), .A2(n6942), .ZN(n6944) );
  AND2_X1 U8016 ( .A1(n6945), .A2(n6944), .ZN(n7525) );
  AND2_X1 U8017 ( .A1(n6946), .A2(n7525), .ZN(n7982) );
  INV_X1 U8018 ( .A(n7981), .ZN(n7526) );
  AND2_X2 U8019 ( .A1(n7982), .A2(n7526), .ZN(n11150) );
  INV_X1 U8020 ( .A(n6947), .ZN(n6957) );
  AND2_X1 U8021 ( .A1(n6949), .A2(n6948), .ZN(n6951) );
  NAND2_X1 U8022 ( .A1(n6950), .A2(n6958), .ZN(n8374) );
  OR2_X1 U8023 ( .A1(n6951), .A2(n8374), .ZN(n10905) );
  OR2_X1 U8024 ( .A1(n10179), .A2(n9893), .ZN(n9747) );
  INV_X1 U8025 ( .A(n9747), .ZN(n9742) );
  NAND2_X1 U8026 ( .A1(n9742), .A2(n7908), .ZN(n10877) );
  NAND2_X1 U8027 ( .A1(n10905), .A2(n10877), .ZN(n11144) );
  NAND2_X1 U8028 ( .A1(n9893), .A2(n6328), .ZN(n9826) );
  INV_X1 U8029 ( .A(n7908), .ZN(n9827) );
  NAND2_X1 U8030 ( .A1(n9835), .A2(n9827), .ZN(n6952) );
  NOR2_X1 U8031 ( .A1(n6953), .A2(n6957), .ZN(n7529) );
  AND2_X1 U8032 ( .A1(n6953), .A2(n6957), .ZN(n9833) );
  NOR2_X1 U8033 ( .A1(n7529), .A2(n9833), .ZN(n9797) );
  INV_X1 U8034 ( .A(n9797), .ZN(n6954) );
  OAI21_X1 U8035 ( .B1(n11144), .B2(n10972), .A(n6954), .ZN(n6956) );
  INV_X1 U8036 ( .A(n5886), .ZN(n7623) );
  INV_X1 U8037 ( .A(n10969), .ZN(n11008) );
  NOR2_X1 U8038 ( .A1(n7623), .A2(n11008), .ZN(n8376) );
  INV_X1 U8039 ( .A(n8376), .ZN(n6955) );
  OAI211_X1 U8040 ( .C1(n6958), .C2(n6957), .A(n6956), .B(n6955), .ZN(n10313)
         );
  NAND2_X1 U8041 ( .A1(n10313), .A2(n11150), .ZN(n6959) );
  OAI21_X1 U8042 ( .B1(n11150), .B2(n5859), .A(n6959), .ZN(P1_U3453) );
  NAND2_X1 U8043 ( .A1(n10147), .A2(n9910), .ZN(n6960) );
  OAI21_X1 U8044 ( .B1(n9910), .B2(n6425), .A(n6960), .ZN(P1_U3577) );
  INV_X1 U8045 ( .A(n10849), .ZN(n10869) );
  OAI21_X1 U8046 ( .B1(n11001), .B2(n6962), .A(n6961), .ZN(n7096) );
  INV_X1 U8047 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n11024) );
  MUX2_X1 U8048 ( .A(n11024), .B(P1_REG1_REG_7__SCAN_IN), .S(n7093), .Z(n7094)
         );
  XOR2_X1 U8049 ( .A(n7096), .B(n7094), .Z(n6964) );
  AND2_X1 U8050 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7402) );
  AOI21_X1 U8051 ( .B1(n10861), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7402), .ZN(
        n6963) );
  OAI21_X1 U8052 ( .B1(n10851), .B2(n6964), .A(n6963), .ZN(n6971) );
  AOI21_X1 U8053 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6966), .A(n6965), .ZN(
        n6969) );
  NAND2_X1 U8054 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n7093), .ZN(n6967) );
  OAI21_X1 U8055 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7093), .A(n6967), .ZN(
        n6968) );
  NOR2_X1 U8056 ( .A1(n6969), .A2(n6968), .ZN(n7090) );
  AOI211_X1 U8057 ( .C1(n6969), .C2(n6968), .A(n7090), .B(n10862), .ZN(n6970)
         );
  AOI211_X1 U8058 ( .C1(n10869), .C2(n7093), .A(n6971), .B(n6970), .ZN(n6972)
         );
  INV_X1 U8059 ( .A(n6972), .ZN(P1_U3250) );
  NAND2_X1 U8060 ( .A1(n6974), .A2(n6973), .ZN(n6976) );
  INV_X1 U8061 ( .A(n7342), .ZN(n7134) );
  INV_X1 U8062 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U8063 ( .A1(n6974), .A2(n6977), .ZN(n6979) );
  NAND2_X1 U8064 ( .A1(n8285), .A2(n8104), .ZN(n6978) );
  AND2_X1 U8065 ( .A1(n6979), .A2(n6978), .ZN(n9509) );
  AND2_X1 U8066 ( .A1(n7134), .A2(n9509), .ZN(n7133) );
  NOR2_X1 U8067 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6983) );
  NOR4_X1 U8068 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6982) );
  NOR4_X1 U8069 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6981) );
  NOR4_X1 U8070 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6980) );
  NAND4_X1 U8071 ( .A1(n6983), .A2(n6982), .A3(n6981), .A4(n6980), .ZN(n6989)
         );
  NOR4_X1 U8072 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6987) );
  NOR4_X1 U8073 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6986) );
  NOR4_X1 U8074 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6985) );
  NOR4_X1 U8075 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6984) );
  NAND4_X1 U8076 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n6988)
         );
  OAI21_X1 U8077 ( .B1(n6989), .B2(n6988), .A(n6974), .ZN(n7130) );
  NAND2_X1 U8078 ( .A1(n7133), .A2(n7130), .ZN(n7109) );
  NAND2_X1 U8079 ( .A1(n8451), .A2(n7997), .ZN(n10987) );
  XNOR2_X1 U8080 ( .A(n6991), .B(n6990), .ZN(n7932) );
  XNOR2_X1 U8081 ( .A(n6992), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8579) );
  OR2_X1 U8082 ( .A1(n10987), .A2(n7348), .ZN(n9233) );
  INV_X1 U8083 ( .A(n7932), .ZN(n8780) );
  NAND2_X1 U8084 ( .A1(n8780), .A2(n8579), .ZN(n8778) );
  OR3_X1 U8085 ( .A1(n8774), .A2(n7997), .A3(n8778), .ZN(n7107) );
  NAND3_X1 U8086 ( .A1(n7107), .A2(n8670), .A3(n10987), .ZN(n6993) );
  NAND2_X1 U8087 ( .A1(n9233), .A2(n6993), .ZN(n7110) );
  NAND2_X1 U8088 ( .A1(n7109), .A2(n7110), .ZN(n6996) );
  INV_X1 U8089 ( .A(n9509), .ZN(n7340) );
  NAND3_X1 U8090 ( .A1(n7342), .A2(n7340), .A3(n7130), .ZN(n7112) );
  INV_X1 U8091 ( .A(n7107), .ZN(n6994) );
  NAND2_X1 U8092 ( .A1(n7112), .A2(n6994), .ZN(n6995) );
  NAND2_X1 U8093 ( .A1(n6996), .A2(n6995), .ZN(n7011) );
  INV_X1 U8094 ( .A(n8579), .ZN(n8779) );
  AND2_X1 U8095 ( .A1(n7932), .A2(n8779), .ZN(n6999) );
  OR2_X1 U8096 ( .A1(n8670), .A2(n6999), .ZN(n7136) );
  NAND3_X1 U8097 ( .A1(n7136), .A2(n6997), .A3(n7991), .ZN(n6998) );
  OAI21_X1 U8098 ( .B1(n7011), .B2(n6998), .A(P2_STATE_REG_SCAN_IN), .ZN(n7001) );
  INV_X1 U8099 ( .A(n6999), .ZN(n8784) );
  OR2_X1 U8100 ( .A1(n8670), .A2(n8784), .ZN(n8790) );
  NOR2_X1 U8101 ( .A1(n8790), .A2(n9508), .ZN(n7012) );
  NAND2_X1 U8102 ( .A1(n7112), .A2(n7012), .ZN(n7000) );
  NOR2_X1 U8103 ( .A1(n9053), .A2(P2_U3151), .ZN(n7200) );
  INV_X1 U8104 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10456) );
  NAND2_X1 U8105 ( .A1(n5126), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U8106 ( .A1(n7223), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U8107 ( .A1(n7194), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7002) );
  NAND2_X1 U8108 ( .A1(n8684), .A2(SI_0_), .ZN(n7007) );
  INV_X1 U8109 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7006) );
  NAND2_X1 U8110 ( .A1(n7007), .A2(n7006), .ZN(n7009) );
  AND2_X1 U8111 ( .A1(n7009), .A2(n7008), .ZN(n9520) );
  AND2_X1 U8112 ( .A1(n9074), .A2(n7140), .ZN(n8452) );
  NOR2_X1 U8113 ( .A1(n8448), .A2(n8452), .ZN(n8744) );
  INV_X1 U8114 ( .A(n8744), .ZN(n7019) );
  INV_X1 U8115 ( .A(n9508), .ZN(n7131) );
  NAND3_X1 U8116 ( .A1(n7131), .A2(n8670), .A3(n10987), .ZN(n7010) );
  INV_X1 U8117 ( .A(n11072), .ZN(n9011) );
  INV_X1 U8118 ( .A(n7354), .ZN(n8455) );
  INV_X1 U8119 ( .A(n7112), .ZN(n7013) );
  AND2_X1 U8120 ( .A1(n7013), .A2(n7012), .ZN(n8950) );
  INV_X1 U8121 ( .A(n8950), .ZN(n11067) );
  NAND2_X1 U8122 ( .A1(n7014), .A2(n8788), .ZN(n7015) );
  AND2_X1 U8123 ( .A1(n7015), .A2(n8884), .ZN(n9193) );
  OR2_X1 U8124 ( .A1(n11067), .A2(n9193), .ZN(n9050) );
  INV_X1 U8125 ( .A(n7109), .ZN(n7016) );
  NOR2_X1 U8126 ( .A1(n9508), .A2(n10987), .ZN(n7115) );
  NAND2_X1 U8127 ( .A1(n7016), .A2(n7115), .ZN(n7017) );
  NAND2_X1 U8128 ( .A1(n7115), .A2(n7348), .ZN(n11102) );
  NAND2_X1 U8129 ( .A1(n7017), .A2(n11102), .ZN(n11077) );
  INV_X1 U8130 ( .A(n11077), .ZN(n9056) );
  OAI22_X1 U8131 ( .A1(n8455), .A2(n9050), .B1(n9056), .B2(n7140), .ZN(n7018)
         );
  AOI21_X1 U8132 ( .B1(n7019), .B2(n9011), .A(n7018), .ZN(n7020) );
  OAI21_X1 U8133 ( .B1(n7200), .B2(n10456), .A(n7020), .ZN(P2_U3172) );
  NAND2_X1 U8134 ( .A1(n7224), .A2(n10658), .ZN(n7383) );
  INV_X1 U8135 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7021) );
  NOR2_X1 U8136 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n7022) );
  INV_X1 U8137 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10626) );
  NAND2_X1 U8138 ( .A1(n8107), .A2(n10626), .ZN(n8185) );
  INV_X1 U8139 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7023) );
  INV_X1 U8140 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10666) );
  INV_X1 U8141 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7024) );
  INV_X1 U8142 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10577) );
  NAND2_X1 U8143 ( .A1(n8608), .A2(n10577), .ZN(n8623) );
  NAND2_X1 U8144 ( .A1(n8623), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7025) );
  NAND2_X1 U8145 ( .A1(n8640), .A2(n7025), .ZN(n9254) );
  NAND2_X1 U8146 ( .A1(n9254), .A2(n8643), .ZN(n7031) );
  INV_X1 U8147 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n7028) );
  NAND2_X1 U8148 ( .A1(n8540), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U8149 ( .A1(n8597), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7026) );
  OAI211_X1 U8150 ( .C1(n5106), .C2(n7028), .A(n7027), .B(n7026), .ZN(n7029)
         );
  INV_X1 U8151 ( .A(n7029), .ZN(n7030) );
  INV_X1 U8152 ( .A(n9238), .ZN(n9260) );
  NAND2_X1 U8153 ( .A1(n9260), .A2(P2_U3893), .ZN(n7032) );
  OAI21_X1 U8154 ( .B1(P2_U3893), .B2(n6424), .A(n7032), .ZN(P2_U3514) );
  NAND2_X1 U8155 ( .A1(n8774), .A2(n7932), .ZN(n7034) );
  AND2_X2 U8156 ( .A1(n7037), .A2(n7036), .ZN(n7376) );
  NAND2_X1 U8157 ( .A1(n7376), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7040) );
  OAI211_X2 U8158 ( .C1(n8399), .C2(n7041), .A(n7040), .B(n7039), .ZN(n8454)
         );
  NAND2_X1 U8159 ( .A1(n7043), .A2(n9011), .ZN(n7047) );
  AND2_X1 U8160 ( .A1(n8950), .A2(n9193), .ZN(n9048) );
  NAND2_X1 U8161 ( .A1(n7223), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U8162 ( .A1(n5126), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7148) );
  NAND2_X1 U8163 ( .A1(n7194), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7146) );
  OAI22_X1 U8164 ( .A1(n7413), .A2(n9050), .B1(n9056), .B2(n7440), .ZN(n7045)
         );
  AOI21_X1 U8165 ( .B1(n9048), .B2(n9074), .A(n7045), .ZN(n7046) );
  OAI211_X1 U8166 ( .C1(n7200), .C2(n10649), .A(n7047), .B(n7046), .ZN(
        P2_U3162) );
  XOR2_X1 U8167 ( .A(n7049), .B(n7048), .Z(n8369) );
  NAND3_X1 U8168 ( .A1(n8369), .A2(n7053), .A3(n10823), .ZN(n7052) );
  NOR2_X1 U8169 ( .A1(n10338), .A2(n10825), .ZN(n7050) );
  OAI211_X1 U8170 ( .C1(n7050), .C2(P1_IR_REG_0__SCAN_IN), .A(n9989), .B(
        n10833), .ZN(n7051) );
  OAI211_X1 U8171 ( .C1(n7053), .C2(n5360), .A(n7052), .B(n7051), .ZN(n7054)
         );
  AND2_X1 U8172 ( .A1(n7054), .A2(P1_U3973), .ZN(n10866) );
  AOI211_X1 U8173 ( .C1(n7057), .C2(n7056), .A(n7055), .B(n10862), .ZN(n7065)
         );
  AOI22_X1 U8174 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .B1(
        P1_ADDR_REG_2__SCAN_IN), .B2(n10861), .ZN(n7062) );
  OAI211_X1 U8175 ( .C1(n7060), .C2(n7059), .A(n10871), .B(n7058), .ZN(n7061)
         );
  OAI211_X1 U8176 ( .C1(n10849), .C2(n7063), .A(n7062), .B(n7061), .ZN(n7064)
         );
  OR3_X1 U8177 ( .A1(n10866), .A2(n7065), .A3(n7064), .ZN(P1_U3245) );
  INV_X1 U8178 ( .A(n7066), .ZN(n7068) );
  AOI21_X1 U8179 ( .B1(n7235), .B2(n7068), .A(n7067), .ZN(n7070) );
  MUX2_X1 U8180 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8381), .Z(n7169) );
  XNOR2_X1 U8181 ( .A(n7169), .B(n5103), .ZN(n7069) );
  NAND2_X1 U8182 ( .A1(n7070), .A2(n7069), .ZN(n7170) );
  OAI211_X1 U8183 ( .C1(n7070), .C2(n7069), .A(n7170), .B(n10352), .ZN(n7084)
         );
  INV_X1 U8184 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7073) );
  AOI21_X1 U8185 ( .B1(n5201), .B2(n7074), .A(n7166), .ZN(n7081) );
  INV_X1 U8186 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U8187 ( .A1(n5103), .A2(P2_REG1_REG_4__SCAN_IN), .B1(n10942), .B2(
        n7175), .ZN(n7075) );
  AOI21_X1 U8188 ( .B1(n7076), .B2(n7075), .A(n7177), .ZN(n7077) );
  NAND2_X1 U8189 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7253) );
  OAI21_X1 U8190 ( .B1(n7077), .B2(n10346), .A(n7253), .ZN(n7078) );
  INV_X1 U8191 ( .A(n7078), .ZN(n7080) );
  NAND2_X1 U8192 ( .A1(n10360), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7079) );
  OAI211_X1 U8193 ( .C1(n7081), .C2(n10348), .A(n7080), .B(n7079), .ZN(n7082)
         );
  AOI21_X1 U8194 ( .B1(n5103), .B2(n9166), .A(n7082), .ZN(n7083) );
  NAND2_X1 U8195 ( .A1(n7084), .A2(n7083), .ZN(P2_U3186) );
  INV_X1 U8196 ( .A(n8117), .ZN(n7088) );
  INV_X1 U8197 ( .A(n7886), .ZN(n10850) );
  INV_X1 U8198 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7085) );
  OAI222_X1 U8199 ( .A1(n10340), .A2(n7088), .B1(n10850), .B2(P1_U3086), .C1(
        n7085), .C2(n10337), .ZN(P1_U3343) );
  INV_X1 U8200 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U8201 ( .A1(n7086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7087) );
  XNOR2_X1 U8202 ( .A(n7087), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8323) );
  INV_X1 U8203 ( .A(n8323), .ZN(n8308) );
  OAI222_X1 U8204 ( .A1(n9516), .A2(n7089), .B1(n9518), .B2(n7088), .C1(n8308), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  AOI22_X1 U8205 ( .A1(n7317), .A2(n6030), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n7323), .ZN(n7091) );
  NOR2_X1 U8206 ( .A1(n7092), .A2(n7091), .ZN(n7316) );
  AOI211_X1 U8207 ( .C1(n7092), .C2(n7091), .A(n7316), .B(n10862), .ZN(n7106)
         );
  NAND2_X1 U8208 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n7093), .ZN(n7098) );
  INV_X1 U8209 ( .A(n7094), .ZN(n7095) );
  NAND2_X1 U8210 ( .A1(n7096), .A2(n7095), .ZN(n7097) );
  NAND2_X1 U8211 ( .A1(n7098), .A2(n7097), .ZN(n7101) );
  INV_X1 U8212 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7099) );
  MUX2_X1 U8213 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7099), .S(n7317), .Z(n7100)
         );
  NAND2_X1 U8214 ( .A1(n7100), .A2(n7101), .ZN(n7322) );
  OAI211_X1 U8215 ( .C1(n7101), .C2(n7100), .A(n10871), .B(n7322), .ZN(n7104)
         );
  INV_X1 U8216 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7102) );
  NOR2_X1 U8217 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7102), .ZN(n9541) );
  AOI21_X1 U8218 ( .B1(n10861), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9541), .ZN(
        n7103) );
  OAI211_X1 U8219 ( .C1(n10849), .C2(n7323), .A(n7104), .B(n7103), .ZN(n7105)
         );
  OR2_X1 U8220 ( .A1(n7106), .A2(n7105), .ZN(P1_U3251) );
  AND2_X1 U8221 ( .A1(n8790), .A2(n7107), .ZN(n7108) );
  OR2_X1 U8222 ( .A1(n7109), .A2(n7108), .ZN(n7114) );
  INV_X1 U8223 ( .A(n7110), .ZN(n7111) );
  OR2_X1 U8224 ( .A1(n7112), .A2(n7111), .ZN(n7113) );
  NAND2_X1 U8225 ( .A1(n7114), .A2(n7113), .ZN(n7122) );
  NAND2_X1 U8226 ( .A1(n7122), .A2(n7115), .ZN(n9503) );
  AOI21_X1 U8227 ( .B1(n8780), .B2(n7997), .A(n8579), .ZN(n7116) );
  AND2_X1 U8228 ( .A1(n10987), .A2(n7116), .ZN(n7117) );
  NAND2_X1 U8229 ( .A1(n7117), .A2(n8790), .ZN(n8883) );
  NAND2_X1 U8230 ( .A1(n7348), .A2(n7997), .ZN(n10954) );
  OR2_X1 U8231 ( .A1(n8451), .A2(n7932), .ZN(n7119) );
  NAND2_X1 U8232 ( .A1(n8579), .A2(n8791), .ZN(n7118) );
  NAND2_X1 U8233 ( .A1(n7119), .A2(n7118), .ZN(n9358) );
  NOR2_X1 U8234 ( .A1(n11119), .A2(n9358), .ZN(n7121) );
  NAND2_X1 U8235 ( .A1(n7354), .A2(n7120), .ZN(n7452) );
  OAI21_X1 U8236 ( .B1(n8744), .B2(n7121), .A(n7452), .ZN(n7142) );
  AND2_X2 U8237 ( .A1(n7122), .A2(n7131), .ZN(n11131) );
  INV_X1 U8238 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7123) );
  NOR2_X1 U8239 ( .A1(n11131), .A2(n7123), .ZN(n7124) );
  AOI21_X1 U8240 ( .B1(n7142), .B2(n11131), .A(n7124), .ZN(n7125) );
  OAI21_X1 U8241 ( .B1(n7140), .B2(n9503), .A(n7125), .ZN(P2_U3390) );
  INV_X1 U8242 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7128) );
  INV_X1 U8243 ( .A(n8111), .ZN(n7129) );
  NAND2_X1 U8244 ( .A1(n7126), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7127) );
  XNOR2_X1 U8245 ( .A(n7127), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9087) );
  INV_X1 U8246 ( .A(n9087), .ZN(n8326) );
  OAI222_X1 U8247 ( .A1(n9516), .A2(n7128), .B1(n9518), .B2(n7129), .C1(
        P2_U3151), .C2(n8326), .ZN(P2_U3282) );
  INV_X1 U8248 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10561) );
  INV_X1 U8249 ( .A(n8093), .ZN(n7894) );
  OAI222_X1 U8250 ( .A1(n10337), .A2(n10561), .B1(n10340), .B2(n7129), .C1(
        P1_U3086), .C2(n7894), .ZN(P1_U3342) );
  NAND2_X1 U8251 ( .A1(n7131), .A2(n7130), .ZN(n7132) );
  NOR2_X1 U8252 ( .A1(n7133), .A2(n7132), .ZN(n7344) );
  OAI21_X1 U8253 ( .B1(n8785), .B2(n10987), .A(n7134), .ZN(n7137) );
  OR3_X1 U8254 ( .A1(n7932), .A2(n8579), .A3(n7997), .ZN(n7135) );
  NAND2_X1 U8255 ( .A1(n8670), .A2(n7135), .ZN(n7341) );
  NAND2_X1 U8256 ( .A1(n7136), .A2(n7341), .ZN(n7339) );
  AOI22_X1 U8257 ( .A1(n7137), .A2(n7339), .B1(n7340), .B2(n7341), .ZN(n7138)
         );
  AND2_X2 U8258 ( .A1(n7344), .A2(n7138), .ZN(n11127) );
  INV_X1 U8259 ( .A(n10987), .ZN(n11121) );
  NAND2_X1 U8260 ( .A1(n11127), .A2(n11121), .ZN(n9445) );
  OAI22_X1 U8261 ( .A1(n9445), .A2(n7140), .B1(n11127), .B2(n7139), .ZN(n7141)
         );
  AOI21_X1 U8262 ( .B1(n7142), .B2(n11127), .A(n7141), .ZN(n7143) );
  INV_X1 U8263 ( .A(n7143), .ZN(P2_U3459) );
  OAI21_X1 U8264 ( .B1(n8741), .B2(n8448), .A(n7346), .ZN(n7444) );
  INV_X1 U8265 ( .A(n7144), .ZN(n7349) );
  XNOR2_X1 U8266 ( .A(n7350), .B(n7349), .ZN(n7145) );
  NAND2_X1 U8267 ( .A1(n7145), .A2(n9358), .ZN(n7151) );
  AOI22_X1 U8268 ( .A1(n7120), .A2(n9072), .B1(n9074), .B2(n9363), .ZN(n7150)
         );
  NAND2_X1 U8269 ( .A1(n7151), .A2(n7150), .ZN(n7441) );
  AOI21_X1 U8270 ( .B1(n11119), .B2(n7444), .A(n7441), .ZN(n7156) );
  INV_X1 U8271 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7152) );
  OAI22_X1 U8272 ( .A1(n9503), .A2(n7440), .B1(n11131), .B2(n7152), .ZN(n7153)
         );
  INV_X1 U8273 ( .A(n7153), .ZN(n7154) );
  OAI21_X1 U8274 ( .B1(n7156), .B2(n11128), .A(n7154), .ZN(P2_U3393) );
  INV_X1 U8275 ( .A(n9445), .ZN(n8018) );
  AOI22_X1 U8276 ( .A1(n8018), .A2(n8454), .B1(n11126), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7155) );
  OAI21_X1 U8277 ( .B1(n7156), .B2(n11126), .A(n7155), .ZN(P2_U3460) );
  NAND2_X1 U8278 ( .A1(n7158), .A2(n7157), .ZN(n7160) );
  XNOR2_X1 U8279 ( .A(n7160), .B(n7159), .ZN(n7165) );
  AOI22_X1 U8280 ( .A1(n9640), .A2(n5839), .B1(n7523), .B2(n9625), .ZN(n7164)
         );
  NOR2_X1 U8281 ( .A1(n7161), .A2(P1_U3086), .ZN(n8373) );
  INV_X1 U8282 ( .A(n8373), .ZN(n7162) );
  AOI22_X1 U8283 ( .A1(n7162), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9623), .B2(
        n6953), .ZN(n7163) );
  OAI211_X1 U8284 ( .C1(n7165), .C2(n9616), .A(n7164), .B(n7163), .ZN(P1_U3222) );
  INV_X1 U8285 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7168) );
  AOI21_X1 U8286 ( .B1(n7168), .B2(n7167), .A(n7269), .ZN(n7185) );
  INV_X1 U8287 ( .A(n7169), .ZN(n7171) );
  OAI21_X1 U8288 ( .B1(n5103), .B2(n7171), .A(n7170), .ZN(n7173) );
  MUX2_X1 U8289 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8381), .Z(n7271) );
  XNOR2_X1 U8290 ( .A(n7271), .B(n7377), .ZN(n7172) );
  NAND2_X1 U8291 ( .A1(n7173), .A2(n7172), .ZN(n7272) );
  OAI211_X1 U8292 ( .C1(n7173), .C2(n7172), .A(n7272), .B(n10352), .ZN(n7184)
         );
  INV_X1 U8293 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7174) );
  NAND2_X1 U8294 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7382) );
  OAI21_X1 U8295 ( .B1(n9158), .B2(n7174), .A(n7382), .ZN(n7182) );
  INV_X1 U8296 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10958) );
  XOR2_X1 U8297 ( .A(n7178), .B(n7278), .Z(n7179) );
  NOR2_X1 U8298 ( .A1(n10958), .A2(n7179), .ZN(n7279) );
  AOI21_X1 U8299 ( .B1(n10958), .B2(n7179), .A(n7279), .ZN(n7180) );
  NOR2_X1 U8300 ( .A1(n7180), .A2(n10346), .ZN(n7181) );
  AOI211_X1 U8301 ( .C1(n9166), .C2(n7377), .A(n7182), .B(n7181), .ZN(n7183)
         );
  OAI211_X1 U8302 ( .C1(n7185), .C2(n10348), .A(n7184), .B(n7183), .ZN(
        P2_U3187) );
  NAND2_X1 U8303 ( .A1(n7376), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7188) );
  NAND2_X1 U8304 ( .A1(n8578), .A2(n7186), .ZN(n7187) );
  OAI211_X1 U8305 ( .C1(n8399), .C2(n7189), .A(n7188), .B(n7187), .ZN(n7347)
         );
  XNOR2_X1 U8306 ( .A(n7347), .B(n5099), .ZN(n7240) );
  XNOR2_X1 U8307 ( .A(n7240), .B(n9072), .ZN(n7241) );
  INV_X1 U8308 ( .A(n7190), .ZN(n7192) );
  OAI21_X1 U8309 ( .B1(n7192), .B2(n7354), .A(n7191), .ZN(n7242) );
  XOR2_X1 U8310 ( .A(n7241), .B(n7242), .Z(n7204) );
  NAND2_X1 U8311 ( .A1(n7223), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7198) );
  INV_X1 U8312 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7193) );
  NAND2_X1 U8313 ( .A1(n5126), .A2(n7193), .ZN(n7197) );
  NAND2_X1 U8314 ( .A1(n8187), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U8315 ( .A1(n7194), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7195) );
  INV_X1 U8316 ( .A(n7347), .ZN(n7412) );
  OAI22_X1 U8317 ( .A1(n7406), .A2(n9050), .B1(n9056), .B2(n7412), .ZN(n7202)
         );
  INV_X1 U8318 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7199) );
  NOR2_X1 U8319 ( .A1(n7200), .A2(n7199), .ZN(n7201) );
  AOI211_X1 U8320 ( .C1(n9048), .C2(n7354), .A(n7202), .B(n7201), .ZN(n7203)
         );
  OAI21_X1 U8321 ( .B1(n7204), .B2(n11072), .A(n7203), .ZN(P2_U3177) );
  INV_X1 U8322 ( .A(n8179), .ZN(n7206) );
  OAI222_X1 U8323 ( .A1(n10337), .A2(n10557), .B1(n10340), .B2(n7206), .C1(
        P1_U3086), .C2(n8103), .ZN(P1_U3341) );
  INV_X1 U8324 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7219) );
  XNOR2_X1 U8325 ( .A(n7205), .B(n7219), .ZN(n8330) );
  OAI222_X1 U8326 ( .A1(n9516), .A2(n7207), .B1(n9518), .B2(n7206), .C1(
        P2_U3151), .C2(n8330), .ZN(P2_U3281) );
  NAND2_X1 U8327 ( .A1(n10060), .A2(n9910), .ZN(n7208) );
  OAI21_X1 U8328 ( .B1(n6507), .B2(n9910), .A(n7208), .ZN(P1_U3580) );
  OAI21_X1 U8329 ( .B1(n7209), .B2(n7210), .A(n5093), .ZN(n7217) );
  INV_X1 U8330 ( .A(n9624), .ZN(n9636) );
  AOI22_X1 U8331 ( .A1(n9623), .A2(n5839), .B1(n9640), .B2(n10968), .ZN(n7215)
         );
  AOI21_X1 U8332 ( .B1(n9625), .B2(n7617), .A(n7213), .ZN(n7214) );
  OAI211_X1 U8333 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9636), .A(n7215), .B(
        n7214), .ZN(n7216) );
  AOI21_X1 U8334 ( .B1(n7217), .B2(n9633), .A(n7216), .ZN(n7218) );
  INV_X1 U8335 ( .A(n7218), .ZN(P1_U3218) );
  INV_X1 U8336 ( .A(n8533), .ZN(n7221) );
  INV_X1 U8337 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10554) );
  OAI222_X1 U8338 ( .A1(n10340), .A2(n7221), .B1(n8154), .B2(P1_U3086), .C1(
        n10554), .C2(n10337), .ZN(P1_U3340) );
  INV_X1 U8339 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7222) );
  NAND2_X1 U8340 ( .A1(n7205), .A2(n7219), .ZN(n7220) );
  NAND2_X1 U8341 ( .A1(n7220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7433) );
  XNOR2_X1 U8342 ( .A(n7433), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8534) );
  INV_X1 U8343 ( .A(n8534), .ZN(n9124) );
  OAI222_X1 U8344 ( .A1(n9516), .A2(n7222), .B1(n9518), .B2(n7221), .C1(n9124), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  NAND2_X1 U8345 ( .A1(n7223), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7230) );
  INV_X1 U8346 ( .A(n7224), .ZN(n7246) );
  NAND2_X1 U8347 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7225) );
  NAND2_X1 U8348 ( .A1(n7246), .A2(n7225), .ZN(n7422) );
  NAND2_X1 U8349 ( .A1(n5126), .A2(n7422), .ZN(n7229) );
  NAND2_X1 U8350 ( .A1(n7194), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8351 ( .A1(n8392), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7233) );
  NAND2_X1 U8352 ( .A1(n8578), .A2(n5103), .ZN(n7232) );
  XNOR2_X1 U8353 ( .A(n5088), .B(n7035), .ZN(n7381) );
  XOR2_X1 U8354 ( .A(n9070), .B(n7381), .Z(n7245) );
  NAND2_X1 U8355 ( .A1(n7376), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U8356 ( .A1(n8578), .A2(n7235), .ZN(n7236) );
  OAI211_X1 U8357 ( .C1(n8399), .C2(n7238), .A(n7237), .B(n7236), .ZN(n10930)
         );
  XNOR2_X1 U8358 ( .A(n10930), .B(n5099), .ZN(n7243) );
  XNOR2_X1 U8359 ( .A(n7243), .B(n9071), .ZN(n8926) );
  AOI21_X1 U8360 ( .B1(n7245), .B2(n7244), .A(n5197), .ZN(n7260) );
  INV_X1 U8361 ( .A(n7422), .ZN(n7257) );
  INV_X1 U8362 ( .A(n9050), .ZN(n9034) );
  NAND2_X1 U8363 ( .A1(n7223), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7252) );
  NAND2_X1 U8364 ( .A1(n7246), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7247) );
  NAND2_X1 U8365 ( .A1(n7383), .A2(n7247), .ZN(n7601) );
  NAND2_X1 U8366 ( .A1(n8643), .A2(n7601), .ZN(n7251) );
  NAND2_X1 U8367 ( .A1(n7226), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7250) );
  NAND2_X1 U8368 ( .A1(n8597), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7249) );
  INV_X1 U8369 ( .A(n7253), .ZN(n7254) );
  AOI21_X1 U8370 ( .B1(n9034), .B2(n9069), .A(n7254), .ZN(n7256) );
  AOI22_X1 U8371 ( .A1(n9048), .A2(n9071), .B1(n11077), .B2(n5088), .ZN(n7255)
         );
  OAI211_X1 U8372 ( .C1(n11079), .C2(n7257), .A(n7256), .B(n7255), .ZN(n7258)
         );
  INV_X1 U8373 ( .A(n7258), .ZN(n7259) );
  OAI21_X1 U8374 ( .B1(n7260), .B2(n11072), .A(n7259), .ZN(P2_U3170) );
  INV_X1 U8375 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7262) );
  INV_X1 U8376 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U8377 ( .A1(n8639), .A2(n8439), .ZN(n8441) );
  NOR2_X1 U8378 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n8441), .ZN(n8419) );
  INV_X1 U8379 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10425) );
  NAND2_X1 U8380 ( .A1(n8419), .A2(n10425), .ZN(n8420) );
  INV_X1 U8381 ( .A(n8420), .ZN(n7261) );
  NAND2_X1 U8382 ( .A1(n7262), .A2(n7261), .ZN(n8410) );
  INV_X1 U8383 ( .A(n8410), .ZN(n8890) );
  NAND2_X1 U8384 ( .A1(n8643), .A2(n8890), .ZN(n8695) );
  NAND2_X1 U8385 ( .A1(n5107), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7265) );
  NAND2_X1 U8386 ( .A1(n8540), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U8387 ( .A1(n8597), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7263) );
  AND4_X1 U8388 ( .A1(n8695), .A2(n7265), .A3(n7264), .A4(n7263), .ZN(n8886)
         );
  NAND2_X1 U8389 ( .A1(n9073), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7266) );
  OAI21_X1 U8390 ( .B1(n8886), .B2(n9073), .A(n7266), .ZN(P2_U3521) );
  NOR2_X1 U8391 ( .A1(n7377), .A2(n7267), .ZN(n7268) );
  INV_X1 U8392 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7573) );
  AOI22_X1 U8393 ( .A1(n7502), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7573), .B2(
        n7561), .ZN(n7270) );
  AOI21_X1 U8394 ( .B1(n5199), .B2(n7270), .A(n7494), .ZN(n7288) );
  INV_X1 U8395 ( .A(n7271), .ZN(n7273) );
  OAI21_X1 U8396 ( .B1(n7377), .B2(n7273), .A(n7272), .ZN(n7275) );
  MUX2_X1 U8397 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8381), .Z(n7499) );
  XNOR2_X1 U8398 ( .A(n7499), .B(n7561), .ZN(n7274) );
  NOR2_X1 U8399 ( .A1(n7275), .A2(n7274), .ZN(n7500) );
  AND2_X1 U8400 ( .A1(n7275), .A2(n7274), .ZN(n7276) );
  OAI21_X1 U8401 ( .B1(n7500), .B2(n7276), .A(n10352), .ZN(n7287) );
  INV_X1 U8402 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7277) );
  NAND2_X1 U8403 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n7578) );
  OAI21_X1 U8404 ( .B1(n9158), .B2(n7277), .A(n7578), .ZN(n7285) );
  NOR2_X1 U8405 ( .A1(n7377), .A2(n7278), .ZN(n7280) );
  INV_X1 U8406 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U8407 ( .A1(n7502), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n10992), .B2(
        n7561), .ZN(n7281) );
  AOI21_X1 U8408 ( .B1(n7282), .B2(n7281), .A(n7511), .ZN(n7283) );
  NOR2_X1 U8409 ( .A1(n7283), .A2(n10346), .ZN(n7284) );
  AOI211_X1 U8410 ( .C1(n9166), .C2(n7502), .A(n7285), .B(n7284), .ZN(n7286)
         );
  OAI211_X1 U8411 ( .C1(n7288), .C2(n10348), .A(n7287), .B(n7286), .ZN(
        P2_U3188) );
  NAND2_X1 U8412 ( .A1(n7291), .A2(n7290), .ZN(n7292) );
  XNOR2_X1 U8413 ( .A(n7293), .B(n7292), .ZN(n7299) );
  AOI22_X1 U8414 ( .A1(n9623), .A2(n9908), .B1(n7783), .B2(n9625), .ZN(n7298)
         );
  NOR2_X1 U8415 ( .A1(n9636), .A2(n7294), .ZN(n7295) );
  AOI211_X1 U8416 ( .C1(n9640), .C2(n9907), .A(n7296), .B(n7295), .ZN(n7297)
         );
  OAI211_X1 U8417 ( .C1(n7299), .C2(n9616), .A(n7298), .B(n7297), .ZN(P1_U3239) );
  NAND2_X1 U8418 ( .A1(n5092), .A2(n9633), .ZN(n7307) );
  AOI21_X1 U8419 ( .B1(n5093), .B2(n7302), .A(n7301), .ZN(n7306) );
  AOI22_X1 U8420 ( .A1(n9623), .A2(n9909), .B1(n9640), .B2(n9908), .ZN(n7305)
         );
  AND2_X1 U8421 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10860) );
  INV_X1 U8422 ( .A(n9625), .ZN(n9643) );
  INV_X1 U8423 ( .A(n7692), .ZN(n10946) );
  NOR2_X1 U8424 ( .A1(n9643), .A2(n10946), .ZN(n7303) );
  AOI211_X1 U8425 ( .C1(n9624), .C2(n7691), .A(n10860), .B(n7303), .ZN(n7304)
         );
  OAI211_X1 U8426 ( .C1(n7307), .C2(n7306), .A(n7305), .B(n7304), .ZN(P1_U3230) );
  XNOR2_X1 U8427 ( .A(n7310), .B(n7309), .ZN(n7315) );
  AOI22_X1 U8428 ( .A1(n9623), .A2(n10968), .B1(n9640), .B2(n10970), .ZN(n7314) );
  INV_X1 U8429 ( .A(n7634), .ZN(n10978) );
  NOR2_X1 U8430 ( .A1(n9643), .A2(n10978), .ZN(n7311) );
  AOI211_X1 U8431 ( .C1(n9624), .C2(n10976), .A(n7312), .B(n7311), .ZN(n7313)
         );
  OAI211_X1 U8432 ( .C1(n7315), .C2(n9616), .A(n7314), .B(n7313), .ZN(P1_U3227) );
  AOI22_X1 U8433 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n7363), .B1(n7367), .B2(
        n7616), .ZN(n7318) );
  NAND2_X1 U8434 ( .A1(n7318), .A2(n7319), .ZN(n7362) );
  AOI221_X1 U8435 ( .B1(n7319), .B2(n7362), .C1(n7318), .C2(n7362), .A(n10862), 
        .ZN(n7320) );
  INV_X1 U8436 ( .A(n7320), .ZN(n7329) );
  AND2_X1 U8437 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7545) );
  INV_X1 U8438 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7321) );
  MUX2_X1 U8439 ( .A(n7321), .B(P1_REG1_REG_9__SCAN_IN), .S(n7363), .Z(n7325)
         );
  OAI21_X1 U8440 ( .B1(n7323), .B2(n7099), .A(n7322), .ZN(n7324) );
  NOR2_X1 U8441 ( .A1(n7325), .A2(n7324), .ZN(n7366) );
  AOI21_X1 U8442 ( .B1(n7325), .B2(n7324), .A(n7366), .ZN(n7326) );
  NOR2_X1 U8443 ( .A1(n10851), .A2(n7326), .ZN(n7327) );
  AOI211_X1 U8444 ( .C1(n10861), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7545), .B(
        n7327), .ZN(n7328) );
  OAI211_X1 U8445 ( .C1(n10849), .C2(n7367), .A(n7329), .B(n7328), .ZN(
        P1_U3252) );
  OAI21_X1 U8446 ( .B1(n7333), .B2(n7330), .A(n7332), .ZN(n7337) );
  INV_X1 U8447 ( .A(n9640), .ZN(n9605) );
  INV_X1 U8448 ( .A(n7334), .ZN(n10888) );
  OAI22_X1 U8449 ( .A1(n9605), .A2(n7628), .B1(n10888), .B2(n9643), .ZN(n7336)
         );
  INV_X1 U8450 ( .A(n9623), .ZN(n9637) );
  INV_X1 U8451 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7750) );
  OAI22_X1 U8452 ( .A1(n9637), .A2(n7623), .B1(n8373), .B2(n7750), .ZN(n7335)
         );
  AOI211_X1 U8453 ( .C1(n7337), .C2(n9633), .A(n7336), .B(n7335), .ZN(n7338)
         );
  INV_X1 U8454 ( .A(n7338), .ZN(P1_U3237) );
  AOI22_X1 U8455 ( .A1(n7342), .A2(n7341), .B1(n7340), .B2(n7339), .ZN(n7343)
         );
  NAND2_X1 U8456 ( .A1(n7344), .A2(n7343), .ZN(n7446) );
  AND2_X1 U8457 ( .A1(n8774), .A2(n7348), .ZN(n7592) );
  INV_X1 U8458 ( .A(n7592), .ZN(n7345) );
  NAND2_X1 U8459 ( .A1(n8883), .A2(n7345), .ZN(n11083) );
  INV_X1 U8460 ( .A(n11104), .ZN(n7361) );
  NAND2_X1 U8461 ( .A1(n8455), .A2(n8454), .ZN(n8449) );
  NAND2_X1 U8462 ( .A1(n9072), .A2(n7412), .ZN(n8463) );
  XNOR2_X1 U8463 ( .A(n8456), .B(n8468), .ZN(n10894) );
  INV_X1 U8464 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7359) );
  NAND2_X1 U8465 ( .A1(n7347), .A2(n11121), .ZN(n10896) );
  NOR2_X1 U8466 ( .A1(n10896), .A2(n7348), .ZN(n7357) );
  NAND2_X1 U8467 ( .A1(n7350), .A2(n7349), .ZN(n7352) );
  NAND2_X1 U8468 ( .A1(n8455), .A2(n7440), .ZN(n7351) );
  NAND2_X1 U8469 ( .A1(n7352), .A2(n7351), .ZN(n7411) );
  XNOR2_X1 U8470 ( .A(n7411), .B(n8468), .ZN(n7353) );
  NAND2_X1 U8471 ( .A1(n7353), .A2(n9358), .ZN(n7356) );
  AOI22_X1 U8472 ( .A1(n9363), .A2(n7354), .B1(n9071), .B2(n7120), .ZN(n7355)
         );
  NAND2_X1 U8473 ( .A1(n7356), .A2(n7355), .ZN(n10893) );
  AOI211_X1 U8474 ( .C1(n11086), .C2(P2_REG3_REG_2__SCAN_IN), .A(n7357), .B(
        n10893), .ZN(n7358) );
  MUX2_X1 U8475 ( .A(n7359), .B(n7358), .S(n11111), .Z(n7360) );
  OAI21_X1 U8476 ( .B1(n7361), .B2(n10894), .A(n7360), .ZN(P2_U3231) );
  AOI22_X1 U8477 ( .A1(n7478), .A2(n6095), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n7483), .ZN(n7364) );
  AOI211_X1 U8478 ( .C1(n7365), .C2(n7364), .A(n7477), .B(n10862), .ZN(n7375)
         );
  AOI21_X1 U8479 ( .B1(n7367), .B2(n7321), .A(n7366), .ZN(n7370) );
  INV_X1 U8480 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7368) );
  MUX2_X1 U8481 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7368), .S(n7478), .Z(n7369)
         );
  NAND2_X1 U8482 ( .A1(n7370), .A2(n7369), .ZN(n7482) );
  OAI211_X1 U8483 ( .C1(n7370), .C2(n7369), .A(n10871), .B(n7482), .ZN(n7373)
         );
  NAND2_X1 U8484 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n7798) );
  INV_X1 U8485 ( .A(n7798), .ZN(n7371) );
  AOI21_X1 U8486 ( .B1(n10861), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7371), .ZN(
        n7372) );
  OAI211_X1 U8487 ( .C1(n10849), .C2(n7483), .A(n7373), .B(n7372), .ZN(n7374)
         );
  OR2_X1 U8488 ( .A1(n7375), .A2(n7374), .ZN(P1_U3253) );
  NAND2_X1 U8489 ( .A1(n8392), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7379) );
  NAND2_X1 U8490 ( .A1(n8578), .A2(n7377), .ZN(n7378) );
  OAI211_X1 U8491 ( .C1(n8399), .C2(n7380), .A(n7379), .B(n7378), .ZN(n7602)
         );
  XNOR2_X1 U8492 ( .A(n7602), .B(n7035), .ZN(n7582) );
  XOR2_X1 U8493 ( .A(n9069), .B(n7582), .Z(n7583) );
  XOR2_X1 U8494 ( .A(n7583), .B(n7584), .Z(n7394) );
  INV_X1 U8495 ( .A(n7602), .ZN(n10953) );
  INV_X1 U8496 ( .A(n7382), .ZN(n7390) );
  NAND2_X1 U8497 ( .A1(n7223), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7388) );
  NAND2_X1 U8498 ( .A1(n7383), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7384) );
  NAND2_X1 U8499 ( .A1(n7552), .A2(n7384), .ZN(n7572) );
  NAND2_X1 U8500 ( .A1(n8643), .A2(n7572), .ZN(n7387) );
  NAND2_X1 U8501 ( .A1(n8187), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U8502 ( .A1(n8597), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7385) );
  NAND4_X1 U8503 ( .A1(n7388), .A2(n7387), .A3(n7386), .A4(n7385), .ZN(n9068)
         );
  NOR2_X1 U8504 ( .A1(n7737), .A2(n9050), .ZN(n7389) );
  AOI211_X1 U8505 ( .C1(n9048), .C2(n9070), .A(n7390), .B(n7389), .ZN(n7391)
         );
  OAI21_X1 U8506 ( .B1(n10953), .B2(n9056), .A(n7391), .ZN(n7392) );
  AOI21_X1 U8507 ( .B1(n7601), .B2(n9053), .A(n7392), .ZN(n7393) );
  OAI21_X1 U8508 ( .B1(n7394), .B2(n11072), .A(n7393), .ZN(P2_U3167) );
  INV_X1 U8509 ( .A(n7618), .ZN(n11030) );
  XNOR2_X1 U8510 ( .A(n7397), .B(n7396), .ZN(n7398) );
  XNOR2_X1 U8511 ( .A(n7395), .B(n7398), .ZN(n7399) );
  NAND2_X1 U8512 ( .A1(n7399), .A2(n9633), .ZN(n7404) );
  INV_X1 U8513 ( .A(n11027), .ZN(n7400) );
  OAI22_X1 U8514 ( .A1(n11011), .A2(n9637), .B1(n9636), .B2(n7400), .ZN(n7401)
         );
  AOI211_X1 U8515 ( .C1(n9640), .C2(n9906), .A(n7402), .B(n7401), .ZN(n7403)
         );
  OAI211_X1 U8516 ( .C1(n11030), .C2(n9643), .A(n7404), .B(n7403), .ZN(
        P1_U3213) );
  NAND2_X1 U8517 ( .A1(n7405), .A2(n5088), .ZN(n8473) );
  NAND2_X1 U8518 ( .A1(n9070), .A2(n10937), .ZN(n8477) );
  AND2_X2 U8519 ( .A1(n8473), .A2(n8477), .ZN(n8747) );
  INV_X1 U8520 ( .A(n8462), .ZN(n8479) );
  NOR2_X1 U8521 ( .A1(n8747), .A2(n8479), .ZN(n7410) );
  INV_X1 U8522 ( .A(n10930), .ZN(n7408) );
  NAND2_X1 U8523 ( .A1(n9071), .A2(n7408), .ZN(n8471) );
  INV_X1 U8524 ( .A(n7566), .ZN(n7409) );
  AOI21_X1 U8525 ( .B1(n7410), .B2(n7425), .A(n7409), .ZN(n10939) );
  NAND2_X1 U8526 ( .A1(n7411), .A2(n8468), .ZN(n7415) );
  NAND2_X1 U8527 ( .A1(n7413), .A2(n7412), .ZN(n7414) );
  NAND2_X1 U8528 ( .A1(n7415), .A2(n7414), .ZN(n7427) );
  NOR2_X1 U8529 ( .A1(n9071), .A2(n10930), .ZN(n7417) );
  NAND2_X1 U8530 ( .A1(n9071), .A2(n10930), .ZN(n7416) );
  XNOR2_X1 U8531 ( .A(n7563), .B(n8747), .ZN(n7418) );
  NAND2_X1 U8532 ( .A1(n7418), .A2(n9358), .ZN(n7420) );
  AOI22_X1 U8533 ( .A1(n7120), .A2(n9069), .B1(n9071), .B2(n9363), .ZN(n7419)
         );
  NAND2_X1 U8534 ( .A1(n7420), .A2(n7419), .ZN(n10940) );
  MUX2_X1 U8535 ( .A(n10940), .B(P2_REG2_REG_4__SCAN_IN), .S(n9352), .Z(n7421)
         );
  INV_X1 U8536 ( .A(n7421), .ZN(n7424) );
  AOI22_X1 U8537 ( .A1(n11106), .A2(n5088), .B1(n11086), .B2(n7422), .ZN(n7423) );
  OAI211_X1 U8538 ( .C1(n10939), .C2(n7361), .A(n7424), .B(n7423), .ZN(
        P2_U3229) );
  OAI21_X1 U8539 ( .B1(n7426), .B2(n8742), .A(n7425), .ZN(n10931) );
  INV_X1 U8540 ( .A(n10931), .ZN(n7431) );
  XOR2_X1 U8541 ( .A(n8742), .B(n7427), .Z(n7428) );
  AOI222_X1 U8542 ( .A1(n9358), .A2(n7428), .B1(n9070), .B2(n7120), .C1(n9072), 
        .C2(n9363), .ZN(n10933) );
  MUX2_X1 U8543 ( .A(n6902), .B(n10933), .S(n11111), .Z(n7430) );
  AOI22_X1 U8544 ( .A1(n11106), .A2(n10930), .B1(n7193), .B2(n11086), .ZN(
        n7429) );
  OAI211_X1 U8545 ( .C1(n7431), .C2(n7361), .A(n7430), .B(n7429), .ZN(P2_U3230) );
  INV_X1 U8546 ( .A(n8537), .ZN(n7439) );
  INV_X1 U8547 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7432) );
  NAND2_X1 U8548 ( .A1(n7433), .A2(n7432), .ZN(n7434) );
  NAND2_X1 U8549 ( .A1(n7434), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7436) );
  INV_X1 U8550 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U8551 ( .A1(n7436), .A2(n7435), .ZN(n7453) );
  OR2_X1 U8552 ( .A1(n7436), .A2(n7435), .ZN(n7437) );
  AND2_X1 U8553 ( .A1(n7453), .A2(n7437), .ZN(n9145) );
  INV_X1 U8554 ( .A(n9145), .ZN(n8335) );
  OAI222_X1 U8555 ( .A1(n9516), .A2(n7438), .B1(n9518), .B2(n7439), .C1(
        P2_U3151), .C2(n8335), .ZN(P2_U3279) );
  INV_X1 U8556 ( .A(n9932), .ZN(n9931) );
  OAI222_X1 U8557 ( .A1(n10337), .A2(n10558), .B1(n10340), .B2(n7439), .C1(
        P1_U3086), .C2(n9931), .ZN(P1_U3339) );
  INV_X1 U8558 ( .A(n8552), .ZN(n7455) );
  INV_X1 U8559 ( .A(n9962), .ZN(n9953) );
  OAI222_X1 U8560 ( .A1(n10340), .A2(n7455), .B1(n9953), .B2(P1_U3086), .C1(
        n10555), .C2(n10337), .ZN(P1_U3338) );
  OAI22_X1 U8561 ( .A1(n9354), .A2(n7440), .B1(n10649), .B2(n11102), .ZN(n7443) );
  MUX2_X1 U8562 ( .A(n7441), .B(P2_REG2_REG_1__SCAN_IN), .S(n9352), .Z(n7442)
         );
  AOI211_X1 U8563 ( .C1(n11104), .C2(n7444), .A(n7443), .B(n7442), .ZN(n7445)
         );
  INV_X1 U8564 ( .A(n7445), .ZN(P2_U3232) );
  INV_X1 U8565 ( .A(n8790), .ZN(n7447) );
  NOR4_X1 U8566 ( .A1(n8744), .A2(n11121), .A3(n7447), .A4(n7446), .ZN(n7448)
         );
  AOI21_X1 U8567 ( .B1(n11086), .B2(P2_REG3_REG_0__SCAN_IN), .A(n7448), .ZN(
        n7451) );
  AOI22_X1 U8568 ( .A1(n9352), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n11106), .B2(
        n7449), .ZN(n7450) );
  OAI211_X1 U8569 ( .C1(n9352), .C2(n7452), .A(n7451), .B(n7450), .ZN(P2_U3233) );
  NAND2_X1 U8570 ( .A1(n7453), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7454) );
  XNOR2_X1 U8571 ( .A(n7454), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9165) );
  INV_X1 U8572 ( .A(n9165), .ZN(n8316) );
  OAI222_X1 U8573 ( .A1(n9516), .A2(n7456), .B1(n9518), .B2(n7455), .C1(n8316), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  NOR2_X1 U8574 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7457) );
  AOI21_X1 U8575 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7457), .ZN(n10822) );
  NOR2_X1 U8576 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7458) );
  AOI21_X1 U8577 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7458), .ZN(n10819) );
  NOR2_X1 U8578 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7459) );
  AOI21_X1 U8579 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7459), .ZN(n10816) );
  NOR2_X1 U8580 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7460) );
  AOI21_X1 U8581 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7460), .ZN(n10813) );
  NOR2_X1 U8582 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7461) );
  AOI21_X1 U8583 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7461), .ZN(n10810) );
  NOR2_X1 U8584 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7462) );
  AOI21_X1 U8585 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7462), .ZN(n10807) );
  NOR2_X1 U8586 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7463) );
  AOI21_X1 U8587 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7463), .ZN(n10804) );
  NOR2_X1 U8588 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7464) );
  AOI21_X1 U8589 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7464), .ZN(n10801) );
  NOR2_X1 U8590 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7465) );
  AOI21_X1 U8591 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7465), .ZN(n10798) );
  NOR2_X1 U8592 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7466) );
  AOI21_X1 U8593 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7466), .ZN(n10795) );
  NOR2_X1 U8594 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7467) );
  AOI21_X1 U8595 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7467), .ZN(n10792) );
  NOR2_X1 U8596 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7468) );
  AOI21_X1 U8597 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7468), .ZN(n10789) );
  NOR2_X1 U8598 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7469) );
  AOI21_X1 U8599 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7469), .ZN(n10786) );
  NOR2_X1 U8600 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7470) );
  AOI21_X1 U8601 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7470), .ZN(n10783) );
  AND2_X1 U8602 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n7471) );
  NOR2_X1 U8603 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7471), .ZN(n10768) );
  INV_X1 U8604 ( .A(n10768), .ZN(n10769) );
  INV_X1 U8605 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10771) );
  NAND3_X1 U8606 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10770) );
  NAND2_X1 U8607 ( .A1(n10771), .A2(n10770), .ZN(n10767) );
  NAND2_X1 U8608 ( .A1(n10769), .A2(n10767), .ZN(n10774) );
  NAND2_X1 U8609 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7472) );
  OAI21_X1 U8610 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7472), .ZN(n10773) );
  NOR2_X1 U8611 ( .A1(n10774), .A2(n10773), .ZN(n10772) );
  AOI21_X1 U8612 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10772), .ZN(n10777) );
  NAND2_X1 U8613 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7473) );
  OAI21_X1 U8614 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7473), .ZN(n10776) );
  NOR2_X1 U8615 ( .A1(n10777), .A2(n10776), .ZN(n10775) );
  AOI21_X1 U8616 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10775), .ZN(n10780) );
  NOR2_X1 U8617 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7474) );
  AOI21_X1 U8618 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7474), .ZN(n10779) );
  NAND2_X1 U8619 ( .A1(n10780), .A2(n10779), .ZN(n10778) );
  OAI21_X1 U8620 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10778), .ZN(n10782) );
  NAND2_X1 U8621 ( .A1(n10783), .A2(n10782), .ZN(n10781) );
  OAI21_X1 U8622 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10781), .ZN(n10785) );
  NAND2_X1 U8623 ( .A1(n10786), .A2(n10785), .ZN(n10784) );
  OAI21_X1 U8624 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10784), .ZN(n10788) );
  NAND2_X1 U8625 ( .A1(n10789), .A2(n10788), .ZN(n10787) );
  OAI21_X1 U8626 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10787), .ZN(n10791) );
  NAND2_X1 U8627 ( .A1(n10792), .A2(n10791), .ZN(n10790) );
  OAI21_X1 U8628 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10790), .ZN(n10794) );
  NAND2_X1 U8629 ( .A1(n10795), .A2(n10794), .ZN(n10793) );
  OAI21_X1 U8630 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10793), .ZN(n10797) );
  NAND2_X1 U8631 ( .A1(n10798), .A2(n10797), .ZN(n10796) );
  OAI21_X1 U8632 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10796), .ZN(n10800) );
  NAND2_X1 U8633 ( .A1(n10801), .A2(n10800), .ZN(n10799) );
  OAI21_X1 U8634 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10799), .ZN(n10803) );
  NAND2_X1 U8635 ( .A1(n10804), .A2(n10803), .ZN(n10802) );
  OAI21_X1 U8636 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10802), .ZN(n10806) );
  NAND2_X1 U8637 ( .A1(n10807), .A2(n10806), .ZN(n10805) );
  OAI21_X1 U8638 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10805), .ZN(n10809) );
  NAND2_X1 U8639 ( .A1(n10810), .A2(n10809), .ZN(n10808) );
  OAI21_X1 U8640 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10808), .ZN(n10812) );
  NAND2_X1 U8641 ( .A1(n10813), .A2(n10812), .ZN(n10811) );
  OAI21_X1 U8642 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10811), .ZN(n10815) );
  NAND2_X1 U8643 ( .A1(n10816), .A2(n10815), .ZN(n10814) );
  OAI21_X1 U8644 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10814), .ZN(n10818) );
  NAND2_X1 U8645 ( .A1(n10819), .A2(n10818), .ZN(n10817) );
  OAI21_X1 U8646 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10817), .ZN(n10821) );
  NAND2_X1 U8647 ( .A1(n10822), .A2(n10821), .ZN(n10820) );
  OAI21_X1 U8648 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10820), .ZN(n7476) );
  XNOR2_X1 U8649 ( .A(n5225), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7475) );
  XNOR2_X1 U8650 ( .A(n7476), .B(n7475), .ZN(ADD_1068_U4) );
  INV_X1 U8651 ( .A(n8564), .ZN(n7492) );
  INV_X1 U8652 ( .A(n9975), .ZN(n9971) );
  INV_X1 U8653 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10562) );
  OAI222_X1 U8654 ( .A1(n10340), .A2(n7492), .B1(n9971), .B2(P1_U3086), .C1(
        n10562), .C2(n10337), .ZN(P1_U3337) );
  AOI22_X1 U8655 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7885), .B1(n7881), .B2(
        n7872), .ZN(n7479) );
  AOI211_X1 U8656 ( .C1(n7480), .C2(n7479), .A(n7880), .B(n10862), .ZN(n7489)
         );
  INV_X1 U8657 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7481) );
  MUX2_X1 U8658 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7481), .S(n7881), .Z(n7485)
         );
  OAI21_X1 U8659 ( .B1(n7483), .B2(n7368), .A(n7482), .ZN(n7484) );
  NAND2_X1 U8660 ( .A1(n7485), .A2(n7484), .ZN(n7884) );
  OAI211_X1 U8661 ( .C1(n7485), .C2(n7484), .A(n10871), .B(n7884), .ZN(n7487)
         );
  AND2_X1 U8662 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7968) );
  AOI21_X1 U8663 ( .B1(n10861), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7968), .ZN(
        n7486) );
  OAI211_X1 U8664 ( .C1(n10849), .C2(n7885), .A(n7487), .B(n7486), .ZN(n7488)
         );
  OR2_X1 U8665 ( .A1(n7489), .A2(n7488), .ZN(P1_U3254) );
  INV_X1 U8666 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7493) );
  XNOR2_X1 U8667 ( .A(n7491), .B(n7490), .ZN(n8565) );
  INV_X1 U8668 ( .A(n8565), .ZN(n8352) );
  OAI222_X1 U8669 ( .A1(n9516), .A2(n7493), .B1(P2_U3151), .B2(n8352), .C1(
        n7492), .C2(n9518), .ZN(P2_U3277) );
  INV_X1 U8670 ( .A(n7495), .ZN(n7496) );
  NAND2_X1 U8671 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7670), .ZN(n7497) );
  OAI21_X1 U8672 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7670), .A(n7497), .ZN(
        n7498) );
  AOI21_X1 U8673 ( .B1(n5610), .B2(n7498), .A(n7669), .ZN(n7522) );
  INV_X1 U8674 ( .A(n7499), .ZN(n7501) );
  AOI21_X1 U8675 ( .B1(n7502), .B2(n7501), .A(n7500), .ZN(n10351) );
  INV_X1 U8676 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7504) );
  INV_X1 U8677 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7503) );
  MUX2_X1 U8678 ( .A(n7504), .B(n7503), .S(n8381), .Z(n7505) );
  XNOR2_X1 U8679 ( .A(n7505), .B(n7512), .ZN(n10350) );
  INV_X1 U8680 ( .A(n7505), .ZN(n7506) );
  OAI22_X1 U8681 ( .A1(n10351), .A2(n10350), .B1(n10356), .B2(n7506), .ZN(
        n7508) );
  MUX2_X1 U8682 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8381), .Z(n7665) );
  INV_X1 U8683 ( .A(n7670), .ZN(n7765) );
  XNOR2_X1 U8684 ( .A(n7665), .B(n7765), .ZN(n7507) );
  NAND2_X1 U8685 ( .A1(n7508), .A2(n7507), .ZN(n7666) );
  OAI21_X1 U8686 ( .B1(n7508), .B2(n7507), .A(n7666), .ZN(n7509) );
  NAND2_X1 U8687 ( .A1(n7509), .A2(n10352), .ZN(n7521) );
  INV_X1 U8688 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U8689 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7773) );
  OAI21_X1 U8690 ( .B1(n9158), .B2(n7510), .A(n7773), .ZN(n7519) );
  NAND2_X1 U8691 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7670), .ZN(n7514) );
  OAI21_X1 U8692 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7670), .A(n7514), .ZN(
        n7515) );
  AOI21_X1 U8693 ( .B1(n7516), .B2(n7515), .A(n7660), .ZN(n7517) );
  NOR2_X1 U8694 ( .A1(n7517), .A2(n10346), .ZN(n7518) );
  AOI211_X1 U8695 ( .C1(n9166), .C2(n7765), .A(n7519), .B(n7518), .ZN(n7520)
         );
  OAI211_X1 U8696 ( .C1(n7522), .C2(n10348), .A(n7521), .B(n7520), .ZN(
        P2_U3190) );
  XNOR2_X1 U8697 ( .A(n10880), .B(n5886), .ZN(n9800) );
  INV_X1 U8698 ( .A(n9800), .ZN(n7530) );
  NAND2_X1 U8699 ( .A1(n6953), .A2(n6947), .ZN(n7622) );
  XNOR2_X1 U8700 ( .A(n7530), .B(n7622), .ZN(n10878) );
  NAND3_X1 U8701 ( .A1(n7526), .A2(n7525), .A3(n7524), .ZN(n7535) );
  INV_X1 U8702 ( .A(n7637), .ZN(n7527) );
  NAND2_X1 U8703 ( .A1(n10218), .A2(n7527), .ZN(n10923) );
  AOI22_X1 U8704 ( .A1(n10969), .A2(n5839), .B1(n6953), .B2(n10967), .ZN(n7533) );
  NAND2_X1 U8705 ( .A1(n7530), .A2(n7529), .ZN(n7606) );
  OAI21_X1 U8706 ( .B1(n7530), .B2(n7529), .A(n7606), .ZN(n7531) );
  NAND2_X1 U8707 ( .A1(n7531), .A2(n10972), .ZN(n7532) );
  OAI211_X1 U8708 ( .C1(n10878), .C2(n10905), .A(n7533), .B(n7532), .ZN(n10881) );
  NAND2_X1 U8709 ( .A1(n10881), .A2(n10218), .ZN(n7542) );
  NOR2_X2 U8710 ( .A1(n7535), .A2(n6328), .ZN(n11035) );
  NAND2_X1 U8711 ( .A1(n7523), .A2(n6947), .ZN(n7536) );
  NAND2_X1 U8712 ( .A1(n7536), .A2(n11006), .ZN(n7537) );
  OR2_X1 U8713 ( .A1(n7537), .A2(n7749), .ZN(n10879) );
  INV_X1 U8714 ( .A(n10879), .ZN(n7538) );
  INV_X1 U8715 ( .A(n10227), .ZN(n11026) );
  AOI22_X1 U8716 ( .A1(n11035), .A2(n7538), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n11026), .ZN(n7539) );
  OAI21_X1 U8717 ( .B1(n6791), .B2(n10218), .A(n7539), .ZN(n7540) );
  AOI21_X1 U8718 ( .B1(n10235), .B2(n7523), .A(n7540), .ZN(n7541) );
  OAI211_X1 U8719 ( .C1(n10878), .C2(n10923), .A(n7542), .B(n7541), .ZN(
        P1_U3292) );
  XOR2_X1 U8720 ( .A(n7544), .B(n7543), .Z(n7550) );
  INV_X1 U8721 ( .A(n9904), .ZN(n7966) );
  AOI22_X1 U8722 ( .A1(n9623), .A2(n9906), .B1(n9624), .B2(n7614), .ZN(n7547)
         );
  INV_X1 U8723 ( .A(n7545), .ZN(n7546) );
  OAI211_X1 U8724 ( .C1(n7966), .C2(n9605), .A(n7547), .B(n7546), .ZN(n7548)
         );
  AOI21_X1 U8725 ( .B1(n7712), .B2(n9625), .A(n7548), .ZN(n7549) );
  OAI21_X1 U8726 ( .B1(n7550), .B2(n9616), .A(n7549), .ZN(P1_U3231) );
  NAND2_X1 U8727 ( .A1(n8540), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7557) );
  INV_X1 U8728 ( .A(n7551), .ZN(n7650) );
  NAND2_X1 U8729 ( .A1(n7552), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7553) );
  NAND2_X1 U8730 ( .A1(n7650), .A2(n7553), .ZN(n7738) );
  NAND2_X1 U8731 ( .A1(n8643), .A2(n7738), .ZN(n7556) );
  NAND2_X1 U8732 ( .A1(n5107), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U8733 ( .A1(n8597), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7554) );
  NAND4_X1 U8734 ( .A1(n7557), .A2(n7556), .A3(n7555), .A4(n7554), .ZN(n9067)
         );
  NAND2_X1 U8735 ( .A1(n7558), .A2(n8110), .ZN(n7560) );
  NAND2_X1 U8736 ( .A1(n8392), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7559) );
  OAI211_X1 U8737 ( .C1(n8884), .C2(n7561), .A(n7560), .B(n7559), .ZN(n7733)
         );
  NAND2_X1 U8738 ( .A1(n7737), .A2(n7733), .ZN(n8499) );
  INV_X1 U8739 ( .A(n7733), .ZN(n10988) );
  NAND2_X1 U8740 ( .A1(n9068), .A2(n10988), .ZN(n8484) );
  NAND2_X1 U8741 ( .A1(n9069), .A2(n7602), .ZN(n7564) );
  XOR2_X1 U8742 ( .A(n8746), .B(n7735), .Z(n7565) );
  INV_X1 U8743 ( .A(n9358), .ZN(n9287) );
  OAI222_X1 U8744 ( .A1(n9289), .A2(n7827), .B1(n9291), .B2(n7567), .C1(n7565), 
        .C2(n9287), .ZN(n10989) );
  INV_X1 U8745 ( .A(n10989), .ZN(n7577) );
  NAND2_X1 U8746 ( .A1(n7566), .A2(n8473), .ZN(n7590) );
  NAND2_X1 U8747 ( .A1(n7567), .A2(n7602), .ZN(n8472) );
  NAND2_X1 U8748 ( .A1(n9069), .A2(n10953), .ZN(n8485) );
  AND2_X1 U8749 ( .A1(n8472), .A2(n8485), .ZN(n8745) );
  NAND2_X1 U8750 ( .A1(n7569), .A2(n8472), .ZN(n7568) );
  INV_X1 U8751 ( .A(n8746), .ZN(n7570) );
  NAND3_X1 U8752 ( .A1(n7569), .A2(n8472), .A3(n7570), .ZN(n7571) );
  NAND2_X1 U8753 ( .A1(n7729), .A2(n7571), .ZN(n10991) );
  NOR2_X1 U8754 ( .A1(n9354), .A2(n10988), .ZN(n7575) );
  INV_X1 U8755 ( .A(n7572), .ZN(n7581) );
  OAI22_X1 U8756 ( .A1(n11111), .A2(n7573), .B1(n7581), .B2(n11102), .ZN(n7574) );
  AOI211_X1 U8757 ( .C1(n10991), .C2(n11104), .A(n7575), .B(n7574), .ZN(n7576)
         );
  OAI21_X1 U8758 ( .B1(n7577), .B2(n9352), .A(n7576), .ZN(P2_U3227) );
  OAI21_X1 U8759 ( .B1(n7827), .B2(n9050), .A(n7578), .ZN(n7579) );
  AOI21_X1 U8760 ( .B1(n9048), .B2(n9069), .A(n7579), .ZN(n7580) );
  OAI21_X1 U8761 ( .B1(n7581), .B2(n11079), .A(n7580), .ZN(n7588) );
  XNOR2_X1 U8762 ( .A(n7733), .B(n7035), .ZN(n7644) );
  XOR2_X1 U8763 ( .A(n9068), .B(n7644), .Z(n7586) );
  AOI211_X1 U8764 ( .C1(n7586), .C2(n7585), .A(n11072), .B(n5196), .ZN(n7587)
         );
  AOI211_X1 U8765 ( .C1(n7733), .C2(n11077), .A(n7588), .B(n7587), .ZN(n7589)
         );
  INV_X1 U8766 ( .A(n7589), .ZN(P2_U3179) );
  OR2_X1 U8767 ( .A1(n7590), .A2(n8745), .ZN(n7591) );
  NAND2_X1 U8768 ( .A1(n7569), .A2(n7591), .ZN(n7597) );
  INV_X1 U8769 ( .A(n7597), .ZN(n10955) );
  NAND2_X1 U8770 ( .A1(n11111), .A2(n7592), .ZN(n8892) );
  INV_X1 U8771 ( .A(n8745), .ZN(n7593) );
  XNOR2_X1 U8772 ( .A(n7594), .B(n7593), .ZN(n7595) );
  NAND2_X1 U8773 ( .A1(n7595), .A2(n9358), .ZN(n7600) );
  INV_X1 U8774 ( .A(n8883), .ZN(n7596) );
  NAND2_X1 U8775 ( .A1(n7597), .A2(n7596), .ZN(n7599) );
  AOI22_X1 U8776 ( .A1(n9363), .A2(n9070), .B1(n9068), .B2(n7120), .ZN(n7598)
         );
  AND3_X1 U8777 ( .A1(n7600), .A2(n7599), .A3(n7598), .ZN(n10952) );
  MUX2_X1 U8778 ( .A(n7168), .B(n10952), .S(n11111), .Z(n7604) );
  AOI22_X1 U8779 ( .A1(n11106), .A2(n7602), .B1(n11086), .B2(n7601), .ZN(n7603) );
  OAI211_X1 U8780 ( .C1(n10955), .C2(n8892), .A(n7604), .B(n7603), .ZN(
        P2_U3228) );
  NAND2_X1 U8781 ( .A1(n7623), .A2(n7523), .ZN(n7605) );
  NAND2_X1 U8782 ( .A1(n7606), .A2(n7605), .ZN(n9841) );
  INV_X1 U8783 ( .A(n5839), .ZN(n10907) );
  NAND2_X1 U8784 ( .A1(n5839), .A2(n10888), .ZN(n9649) );
  NAND2_X1 U8785 ( .A1(n10909), .A2(n9649), .ZN(n9648) );
  INV_X1 U8786 ( .A(n9648), .ZN(n9798) );
  NAND2_X1 U8787 ( .A1(n9841), .A2(n9798), .ZN(n10910) );
  NAND2_X1 U8788 ( .A1(n7628), .A2(n7617), .ZN(n9844) );
  NAND3_X1 U8789 ( .A1(n10910), .A2(n9844), .A3(n10909), .ZN(n7607) );
  NAND2_X1 U8790 ( .A1(n10968), .A2(n10946), .ZN(n9842) );
  INV_X1 U8791 ( .A(n7617), .ZN(n10921) );
  NAND2_X1 U8792 ( .A1(n9909), .A2(n10921), .ZN(n9650) );
  NAND3_X1 U8793 ( .A1(n7607), .A2(n9842), .A3(n9650), .ZN(n9654) );
  INV_X1 U8794 ( .A(n10968), .ZN(n10906) );
  NAND2_X1 U8795 ( .A1(n10906), .A2(n7692), .ZN(n9651) );
  INV_X1 U8796 ( .A(n9908), .ZN(n7608) );
  NAND2_X1 U8797 ( .A1(n7608), .A2(n7634), .ZN(n7633) );
  AND2_X1 U8798 ( .A1(n9651), .A2(n7633), .ZN(n9655) );
  NAND2_X1 U8799 ( .A1(n9654), .A2(n9655), .ZN(n7609) );
  NAND2_X1 U8800 ( .A1(n9908), .A2(n10978), .ZN(n9846) );
  NAND2_X1 U8801 ( .A1(n7609), .A2(n9846), .ZN(n7786) );
  NAND2_X1 U8802 ( .A1(n11011), .A2(n7783), .ZN(n9851) );
  NAND2_X1 U8803 ( .A1(n7786), .A2(n9851), .ZN(n11012) );
  INV_X1 U8804 ( .A(n9907), .ZN(n7636) );
  NAND2_X1 U8805 ( .A1(n7636), .A2(n7618), .ZN(n9678) );
  NAND2_X1 U8806 ( .A1(n9907), .A2(n11030), .ZN(n9670) );
  NAND2_X1 U8807 ( .A1(n9678), .A2(n9670), .ZN(n11013) );
  INV_X1 U8808 ( .A(n7783), .ZN(n10997) );
  NAND2_X1 U8809 ( .A1(n10970), .A2(n10997), .ZN(n9660) );
  INV_X1 U8810 ( .A(n9660), .ZN(n11014) );
  NOR2_X1 U8811 ( .A1(n11013), .A2(n11014), .ZN(n7610) );
  NAND2_X1 U8812 ( .A1(n11012), .A2(n7610), .ZN(n11017) );
  INV_X1 U8813 ( .A(n9906), .ZN(n11009) );
  NAND2_X1 U8814 ( .A1(n11009), .A2(n9543), .ZN(n7717) );
  INV_X1 U8815 ( .A(n9543), .ZN(n11041) );
  NAND2_X1 U8816 ( .A1(n11041), .A2(n9906), .ZN(n7715) );
  NAND3_X1 U8817 ( .A1(n11017), .A2(n9668), .A3(n9678), .ZN(n7611) );
  NAND2_X1 U8818 ( .A1(n7611), .A2(n7715), .ZN(n7612) );
  OR2_X1 U8819 ( .A1(n7722), .A2(n7712), .ZN(n9669) );
  NAND2_X1 U8820 ( .A1(n7712), .A2(n7722), .ZN(n9677) );
  NAND2_X1 U8821 ( .A1(n9669), .A2(n9677), .ZN(n7713) );
  XNOR2_X1 U8822 ( .A(n7612), .B(n7713), .ZN(n7613) );
  AOI22_X1 U8823 ( .A1(n7613), .A2(n10972), .B1(n10967), .B2(n9906), .ZN(
        n11049) );
  INV_X1 U8824 ( .A(n7614), .ZN(n7615) );
  OAI22_X1 U8825 ( .A1(n10218), .A2(n7616), .B1(n7615), .B2(n10227), .ZN(n7621) );
  NAND2_X1 U8826 ( .A1(n7749), .A2(n10888), .ZN(n10902) );
  OR2_X1 U8827 ( .A1(n10902), .A2(n7617), .ZN(n10903) );
  INV_X1 U8828 ( .A(n11006), .ZN(n11042) );
  AOI211_X1 U8829 ( .C1(n7712), .C2(n7704), .A(n11042), .B(n7723), .ZN(n7619)
         );
  AOI21_X1 U8830 ( .B1(n10969), .B2(n9904), .A(n7619), .ZN(n11048) );
  INV_X1 U8831 ( .A(n11035), .ZN(n10231) );
  NOR2_X1 U8832 ( .A1(n11048), .A2(n10231), .ZN(n7620) );
  AOI211_X1 U8833 ( .C1(n10235), .C2(n7712), .A(n7621), .B(n7620), .ZN(n7640)
         );
  NAND2_X1 U8834 ( .A1(n9800), .A2(n7622), .ZN(n7625) );
  NAND2_X1 U8835 ( .A1(n7623), .A2(n10880), .ZN(n7624) );
  NAND2_X1 U8836 ( .A1(n7625), .A2(n7624), .ZN(n7745) );
  NAND2_X1 U8837 ( .A1(n7745), .A2(n9648), .ZN(n7627) );
  NAND2_X1 U8838 ( .A1(n10907), .A2(n10888), .ZN(n7626) );
  NAND2_X1 U8839 ( .A1(n7627), .A2(n7626), .ZN(n10901) );
  NAND2_X1 U8840 ( .A1(n10901), .A2(n10908), .ZN(n7630) );
  NAND2_X1 U8841 ( .A1(n7628), .A2(n10921), .ZN(n7629) );
  NAND2_X1 U8842 ( .A1(n7630), .A2(n7629), .ZN(n7688) );
  NAND2_X1 U8843 ( .A1(n9651), .A2(n9842), .ZN(n9799) );
  NAND2_X1 U8844 ( .A1(n7688), .A2(n9799), .ZN(n7632) );
  NAND2_X1 U8845 ( .A1(n10906), .A2(n10946), .ZN(n7631) );
  NOR2_X1 U8846 ( .A1(n9908), .A2(n7634), .ZN(n7635) );
  OAI22_X2 U8847 ( .A1(n7781), .A2(n9658), .B1(n7783), .B2(n10970), .ZN(n11003) );
  AOI22_X2 U8848 ( .A1(n11003), .A2(n11013), .B1(n11030), .B2(n7636), .ZN(
        n7699) );
  XNOR2_X1 U8849 ( .A(n7714), .B(n7713), .ZN(n11052) );
  AND2_X1 U8850 ( .A1(n10905), .A2(n7637), .ZN(n7638) );
  NAND2_X1 U8851 ( .A1(n11052), .A2(n10982), .ZN(n7639) );
  OAI211_X1 U8852 ( .C1(n11028), .C2(n11049), .A(n7640), .B(n7639), .ZN(
        P1_U3284) );
  NAND2_X1 U8853 ( .A1(n7641), .A2(n8110), .ZN(n7643) );
  AOI22_X1 U8854 ( .A1(n8392), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8578), .B2(
        n7512), .ZN(n7642) );
  NAND2_X1 U8855 ( .A1(n7643), .A2(n7642), .ZN(n7759) );
  INV_X1 U8856 ( .A(n7644), .ZN(n7645) );
  XNOR2_X1 U8857 ( .A(n7759), .B(n5099), .ZN(n7762) );
  XNOR2_X1 U8858 ( .A(n7762), .B(n9067), .ZN(n7646) );
  OAI21_X1 U8859 ( .B1(n7647), .B2(n7646), .A(n7763), .ZN(n7648) );
  NAND2_X1 U8860 ( .A1(n7648), .A2(n9011), .ZN(n7659) );
  NAND2_X1 U8861 ( .A1(n8540), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7655) );
  INV_X1 U8862 ( .A(n7649), .ZN(n7810) );
  NAND2_X1 U8863 ( .A1(n7650), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U8864 ( .A1(n7810), .A2(n7651), .ZN(n7828) );
  NAND2_X1 U8865 ( .A1(n8643), .A2(n7828), .ZN(n7654) );
  NAND2_X1 U8866 ( .A1(n5107), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U8867 ( .A1(n8597), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7652) );
  NAND4_X1 U8868 ( .A1(n7655), .A2(n7654), .A3(n7653), .A4(n7652), .ZN(n9066)
         );
  NAND2_X1 U8869 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3151), .ZN(n10354) );
  NAND2_X1 U8870 ( .A1(n9048), .A2(n9068), .ZN(n7656) );
  OAI211_X1 U8871 ( .C1(n7922), .C2(n9050), .A(n10354), .B(n7656), .ZN(n7657)
         );
  AOI21_X1 U8872 ( .B1(n9053), .B2(n7738), .A(n7657), .ZN(n7658) );
  OAI211_X1 U8873 ( .C1(n7823), .C2(n9056), .A(n7659), .B(n7658), .ZN(P2_U3153) );
  XNOR2_X1 U8874 ( .A(n7845), .B(n7852), .ZN(n7662) );
  INV_X1 U8875 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7661) );
  NOR2_X1 U8876 ( .A1(n7661), .A2(n7662), .ZN(n7846) );
  AOI21_X1 U8877 ( .B1(n7662), .B2(n7661), .A(n7846), .ZN(n7681) );
  MUX2_X1 U8878 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8381), .Z(n7664) );
  INV_X1 U8879 ( .A(n7852), .ZN(n7663) );
  NOR2_X1 U8880 ( .A1(n7664), .A2(n7663), .ZN(n7834) );
  AND2_X1 U8881 ( .A1(n7664), .A2(n7663), .ZN(n7833) );
  NOR2_X1 U8882 ( .A1(n7834), .A2(n7833), .ZN(n7668) );
  OR2_X1 U8883 ( .A1(n7665), .A2(n7670), .ZN(n7667) );
  NAND2_X1 U8884 ( .A1(n7667), .A2(n7666), .ZN(n7835) );
  XNOR2_X1 U8885 ( .A(n7668), .B(n7835), .ZN(n7679) );
  INV_X1 U8886 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7672) );
  XNOR2_X1 U8887 ( .A(n7851), .B(n7852), .ZN(n7671) );
  NOR2_X1 U8888 ( .A1(n7672), .A2(n7671), .ZN(n7853) );
  AOI21_X1 U8889 ( .B1(n7672), .B2(n7671), .A(n7853), .ZN(n7677) );
  INV_X1 U8890 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7673) );
  NOR2_X1 U8891 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7673), .ZN(n7816) );
  INV_X1 U8892 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7674) );
  NOR2_X1 U8893 ( .A1(n9158), .A2(n7674), .ZN(n7675) );
  AOI211_X1 U8894 ( .C1(n9166), .C2(n7852), .A(n7816), .B(n7675), .ZN(n7676)
         );
  OAI21_X1 U8895 ( .B1(n7677), .B2(n10348), .A(n7676), .ZN(n7678) );
  AOI21_X1 U8896 ( .B1(n10352), .B2(n7679), .A(n7678), .ZN(n7680) );
  OAI21_X1 U8897 ( .B1(n7681), .B2(n10346), .A(n7680), .ZN(P2_U3191) );
  NAND2_X1 U8898 ( .A1(n10910), .A2(n10909), .ZN(n7682) );
  INV_X1 U8899 ( .A(n10908), .ZN(n9796) );
  NAND2_X1 U8900 ( .A1(n7682), .A2(n9796), .ZN(n10912) );
  NAND2_X1 U8901 ( .A1(n10912), .A2(n9844), .ZN(n7684) );
  INV_X1 U8902 ( .A(n9799), .ZN(n7683) );
  XNOR2_X1 U8903 ( .A(n7684), .B(n7683), .ZN(n7685) );
  NAND2_X1 U8904 ( .A1(n7685), .A2(n10972), .ZN(n7687) );
  AOI22_X1 U8905 ( .A1(n10967), .A2(n9909), .B1(n9908), .B2(n10969), .ZN(n7686) );
  AND2_X1 U8906 ( .A1(n7687), .A2(n7686), .ZN(n10950) );
  XNOR2_X1 U8907 ( .A(n7688), .B(n9799), .ZN(n10948) );
  NAND2_X1 U8908 ( .A1(n10903), .A2(n7692), .ZN(n7689) );
  NAND2_X1 U8909 ( .A1(n7689), .A2(n11006), .ZN(n7690) );
  OR2_X1 U8910 ( .A1(n7690), .A2(n10964), .ZN(n10945) );
  AOI22_X1 U8911 ( .A1(n10180), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7691), .B2(
        n11026), .ZN(n7694) );
  NAND2_X1 U8912 ( .A1(n10235), .A2(n7692), .ZN(n7693) );
  OAI211_X1 U8913 ( .C1(n10945), .C2(n10231), .A(n7694), .B(n7693), .ZN(n7695)
         );
  AOI21_X1 U8914 ( .B1(n10948), .B2(n10982), .A(n7695), .ZN(n7696) );
  OAI21_X1 U8915 ( .B1(n10950), .B2(n10180), .A(n7696), .ZN(P1_U3289) );
  INV_X1 U8916 ( .A(n8577), .ZN(n7697) );
  OAI222_X1 U8917 ( .A1(n10337), .A2(n10695), .B1(n10340), .B2(n7697), .C1(
        P1_U3086), .C2(n10179), .ZN(P1_U3336) );
  OAI222_X1 U8918 ( .A1(n9516), .A2(n7698), .B1(n9518), .B2(n7697), .C1(
        P2_U3151), .C2(n8779), .ZN(P2_U3276) );
  XNOR2_X1 U8919 ( .A(n7699), .B(n9668), .ZN(n11046) );
  INV_X1 U8920 ( .A(n11046), .ZN(n7711) );
  NAND2_X1 U8921 ( .A1(n11017), .A2(n9678), .ZN(n7700) );
  XNOR2_X1 U8922 ( .A(n7700), .B(n9668), .ZN(n7701) );
  NAND2_X1 U8923 ( .A1(n7701), .A2(n10972), .ZN(n7703) );
  AOI22_X1 U8924 ( .A1(n10969), .A2(n9905), .B1(n9907), .B2(n10967), .ZN(n7702) );
  NAND2_X1 U8925 ( .A1(n7703), .A2(n7702), .ZN(n11044) );
  INV_X1 U8926 ( .A(n11005), .ZN(n7705) );
  OAI21_X1 U8927 ( .B1(n7705), .B2(n11041), .A(n7704), .ZN(n11043) );
  AND2_X1 U8928 ( .A1(n11035), .A2(n11006), .ZN(n10153) );
  INV_X1 U8929 ( .A(n10153), .ZN(n7708) );
  AOI22_X1 U8930 ( .A1(n10180), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9542), .B2(
        n11026), .ZN(n7707) );
  NAND2_X1 U8931 ( .A1(n10235), .A2(n9543), .ZN(n7706) );
  OAI211_X1 U8932 ( .C1(n11043), .C2(n7708), .A(n7707), .B(n7706), .ZN(n7709)
         );
  AOI21_X1 U8933 ( .B1(n11044), .B2(n10218), .A(n7709), .ZN(n7710) );
  OAI21_X1 U8934 ( .B1(n7711), .B2(n10220), .A(n7710), .ZN(P1_U3285) );
  INV_X1 U8935 ( .A(n7712), .ZN(n11050) );
  OR2_X1 U8936 ( .A1(n7864), .A2(n7966), .ZN(n9853) );
  NAND2_X1 U8937 ( .A1(n7864), .A2(n7966), .ZN(n9672) );
  XNOR2_X1 U8938 ( .A(n7866), .B(n7865), .ZN(n11057) );
  INV_X1 U8939 ( .A(n11057), .ZN(n7728) );
  INV_X1 U8940 ( .A(n9903), .ZN(n7902) );
  NAND2_X1 U8941 ( .A1(n9669), .A2(n7715), .ZN(n9679) );
  NAND2_X1 U8942 ( .A1(n9660), .A2(n9670), .ZN(n7716) );
  NAND2_X1 U8943 ( .A1(n9677), .A2(n7717), .ZN(n9671) );
  INV_X1 U8944 ( .A(n9678), .ZN(n7718) );
  OR2_X1 U8945 ( .A1(n9671), .A2(n7718), .ZN(n9802) );
  NAND2_X1 U8946 ( .A1(n9679), .A2(n9677), .ZN(n7719) );
  AOI21_X1 U8947 ( .B1(n7720), .B2(n5683), .A(n7900), .ZN(n7721) );
  OAI222_X1 U8948 ( .A1(n11010), .A2(n7722), .B1(n11008), .B2(n7902), .C1(
        n11016), .C2(n7721), .ZN(n11055) );
  NAND2_X1 U8949 ( .A1(n7723), .A2(n5681), .ZN(n7873) );
  OAI211_X1 U8950 ( .C1(n7723), .C2(n5681), .A(n7873), .B(n11006), .ZN(n11054)
         );
  AOI22_X1 U8951 ( .A1(n10180), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7797), .B2(
        n11026), .ZN(n7725) );
  NAND2_X1 U8952 ( .A1(n10235), .A2(n7864), .ZN(n7724) );
  OAI211_X1 U8953 ( .C1(n11054), .C2(n10231), .A(n7725), .B(n7724), .ZN(n7726)
         );
  AOI21_X1 U8954 ( .B1(n11055), .B2(n10218), .A(n7726), .ZN(n7727) );
  OAI21_X1 U8955 ( .B1(n7728), .B2(n10220), .A(n7727), .ZN(P1_U3283) );
  NAND2_X1 U8956 ( .A1(n7827), .A2(n7759), .ZN(n8494) );
  NAND2_X1 U8957 ( .A1(n7823), .A2(n9067), .ZN(n7923) );
  NAND2_X1 U8958 ( .A1(n8494), .A2(n7923), .ZN(n8750) );
  INV_X1 U8959 ( .A(n8750), .ZN(n7730) );
  NAND2_X1 U8960 ( .A1(n7731), .A2(n8750), .ZN(n7732) );
  AND2_X1 U8961 ( .A1(n7924), .A2(n7732), .ZN(n7755) );
  INV_X1 U8962 ( .A(n7755), .ZN(n7744) );
  AND2_X1 U8963 ( .A1(n9068), .A2(n7733), .ZN(n7734) );
  XOR2_X1 U8964 ( .A(n7822), .B(n8750), .Z(n7736) );
  OAI222_X1 U8965 ( .A1(n9289), .A2(n7922), .B1(n9291), .B2(n7737), .C1(n9287), 
        .C2(n7736), .ZN(n7754) );
  NAND2_X1 U8966 ( .A1(n7754), .A2(n11111), .ZN(n7743) );
  INV_X1 U8967 ( .A(n7738), .ZN(n7739) );
  OAI22_X1 U8968 ( .A1(n11111), .A2(n7504), .B1(n7739), .B2(n11102), .ZN(n7741) );
  NOR2_X1 U8969 ( .A1(n9354), .A2(n7823), .ZN(n7740) );
  NOR2_X1 U8970 ( .A1(n7741), .A2(n7740), .ZN(n7742) );
  OAI211_X1 U8971 ( .C1(n7744), .C2(n7361), .A(n7743), .B(n7742), .ZN(P2_U3226) );
  XNOR2_X1 U8972 ( .A(n7745), .B(n9798), .ZN(n10886) );
  OAI21_X1 U8973 ( .B1(n9798), .B2(n9841), .A(n10910), .ZN(n7746) );
  NAND2_X1 U8974 ( .A1(n7746), .A2(n10972), .ZN(n7748) );
  AOI22_X1 U8975 ( .A1(n10967), .A2(n5886), .B1(n9909), .B2(n10969), .ZN(n7747) );
  NAND2_X1 U8976 ( .A1(n7748), .A2(n7747), .ZN(n10891) );
  OAI211_X1 U8977 ( .C1(n7749), .C2(n10888), .A(n10902), .B(n11006), .ZN(
        n10887) );
  OAI22_X1 U8978 ( .A1(n10887), .A2(n6328), .B1(n10227), .B2(n7750), .ZN(n7751) );
  OAI21_X1 U8979 ( .B1(n10891), .B2(n7751), .A(n10218), .ZN(n7753) );
  AOI22_X1 U8980 ( .A1(n10235), .A2(n7334), .B1(n11028), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n7752) );
  OAI211_X1 U8981 ( .C1(n10886), .C2(n10220), .A(n7753), .B(n7752), .ZN(
        P1_U3291) );
  AOI21_X1 U8982 ( .B1(n7755), .B2(n11119), .A(n7754), .ZN(n7761) );
  INV_X1 U8983 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7756) );
  OAI22_X1 U8984 ( .A1(n9503), .A2(n7823), .B1(n11131), .B2(n7756), .ZN(n7757)
         );
  INV_X1 U8985 ( .A(n7757), .ZN(n7758) );
  OAI21_X1 U8986 ( .B1(n7761), .B2(n11128), .A(n7758), .ZN(P2_U3411) );
  AOI22_X1 U8987 ( .A1(n8018), .A2(n7759), .B1(n11126), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7760) );
  OAI21_X1 U8988 ( .B1(n7761), .B2(n11126), .A(n7760), .ZN(P2_U3466) );
  NAND2_X1 U8989 ( .A1(n7764), .A2(n8689), .ZN(n7767) );
  AOI22_X1 U8990 ( .A1(n8392), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8578), .B2(
        n7765), .ZN(n7766) );
  NAND2_X1 U8991 ( .A1(n7767), .A2(n7766), .ZN(n7919) );
  XOR2_X1 U8992 ( .A(n5099), .B(n7919), .Z(n7803) );
  XNOR2_X1 U8993 ( .A(n7803), .B(n9066), .ZN(n7768) );
  XNOR2_X1 U8994 ( .A(n7806), .B(n7768), .ZN(n7780) );
  INV_X1 U8995 ( .A(n7828), .ZN(n7777) );
  NAND2_X1 U8996 ( .A1(n7223), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7772) );
  XNOR2_X1 U8997 ( .A(n7810), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U8998 ( .A1(n8643), .A2(n7926), .ZN(n7771) );
  NAND2_X1 U8999 ( .A1(n5107), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U9000 ( .A1(n8597), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7769) );
  NAND4_X1 U9001 ( .A1(n7772), .A2(n7771), .A3(n7770), .A4(n7769), .ZN(n9065)
         );
  INV_X1 U9002 ( .A(n7773), .ZN(n7774) );
  AOI21_X1 U9003 ( .B1(n9034), .B2(n9065), .A(n7774), .ZN(n7776) );
  NAND2_X1 U9004 ( .A1(n9048), .A2(n9067), .ZN(n7775) );
  OAI211_X1 U9005 ( .C1(n11079), .C2(n7777), .A(n7776), .B(n7775), .ZN(n7778)
         );
  AOI21_X1 U9006 ( .B1(n7919), .B2(n11077), .A(n7778), .ZN(n7779) );
  OAI21_X1 U9007 ( .B1(n7780), .B2(n11072), .A(n7779), .ZN(P2_U3161) );
  XNOR2_X1 U9008 ( .A(n7781), .B(n9658), .ZN(n10995) );
  OAI211_X1 U9009 ( .C1(n10962), .C2(n10997), .A(n11006), .B(n11004), .ZN(
        n10996) );
  AOI22_X1 U9010 ( .A1(n10235), .A2(n7783), .B1(n11026), .B2(n7782), .ZN(n7784) );
  OAI21_X1 U9011 ( .B1(n10996), .B2(n10231), .A(n7784), .ZN(n7791) );
  INV_X1 U9012 ( .A(n9658), .ZN(n7785) );
  XNOR2_X1 U9013 ( .A(n7786), .B(n7785), .ZN(n7787) );
  NAND2_X1 U9014 ( .A1(n7787), .A2(n10972), .ZN(n7789) );
  AOI22_X1 U9015 ( .A1(n10967), .A2(n9908), .B1(n9907), .B2(n10969), .ZN(n7788) );
  NAND2_X1 U9016 ( .A1(n7789), .A2(n7788), .ZN(n10999) );
  MUX2_X1 U9017 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10999), .S(n10218), .Z(n7790) );
  AOI211_X1 U9018 ( .C1(n10982), .C2(n10995), .A(n7791), .B(n7790), .ZN(n7792)
         );
  INV_X1 U9019 ( .A(n7792), .ZN(P1_U3287) );
  NAND2_X1 U9020 ( .A1(n5094), .A2(n7794), .ZN(n7796) );
  XNOR2_X1 U9021 ( .A(n7796), .B(n7795), .ZN(n7802) );
  AOI22_X1 U9022 ( .A1(n9623), .A2(n9905), .B1(n9624), .B2(n7797), .ZN(n7799)
         );
  OAI211_X1 U9023 ( .C1(n7902), .C2(n9605), .A(n7799), .B(n7798), .ZN(n7800)
         );
  AOI21_X1 U9024 ( .B1(n7864), .B2(n9625), .A(n7800), .ZN(n7801) );
  OAI21_X1 U9025 ( .B1(n7802), .B2(n9616), .A(n7801), .ZN(P1_U3217) );
  NOR2_X1 U9026 ( .A1(n7803), .A2(n9066), .ZN(n7805) );
  INV_X1 U9027 ( .A(n7803), .ZN(n7804) );
  NAND2_X1 U9028 ( .A1(n7807), .A2(n8689), .ZN(n7809) );
  AOI22_X1 U9029 ( .A1(n8392), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8578), .B2(
        n7852), .ZN(n7808) );
  NAND2_X2 U9030 ( .A1(n7809), .A2(n7808), .ZN(n7976) );
  XNOR2_X1 U9031 ( .A(n7976), .B(n5099), .ZN(n8070) );
  XNOR2_X1 U9032 ( .A(n8070), .B(n9065), .ZN(n8072) );
  XNOR2_X1 U9033 ( .A(n8073), .B(n8072), .ZN(n7821) );
  INV_X1 U9034 ( .A(n9048), .ZN(n9037) );
  NAND2_X1 U9035 ( .A1(n9053), .A2(n7926), .ZN(n7818) );
  NAND2_X1 U9036 ( .A1(n7223), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7815) );
  OAI21_X1 U9037 ( .B1(n7810), .B2(P2_REG3_REG_9__SCAN_IN), .A(
        P2_REG3_REG_10__SCAN_IN), .ZN(n7811) );
  NAND2_X1 U9038 ( .A1(n7811), .A2(n7942), .ZN(n8077) );
  NAND2_X1 U9039 ( .A1(n8643), .A2(n8077), .ZN(n7814) );
  NAND2_X1 U9040 ( .A1(n8187), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U9041 ( .A1(n7194), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7812) );
  NAND4_X1 U9042 ( .A1(n7815), .A2(n7814), .A3(n7813), .A4(n7812), .ZN(n9064)
         );
  AOI21_X1 U9043 ( .B1(n9034), .B2(n9064), .A(n7816), .ZN(n7817) );
  OAI211_X1 U9044 ( .C1(n7922), .C2(n9037), .A(n7818), .B(n7817), .ZN(n7819)
         );
  AOI21_X1 U9045 ( .B1(n7976), .B2(n11077), .A(n7819), .ZN(n7820) );
  OAI21_X1 U9046 ( .B1(n7821), .B2(n11072), .A(n7820), .ZN(P2_U3171) );
  NAND2_X1 U9047 ( .A1(n7822), .A2(n8750), .ZN(n7825) );
  NAND2_X1 U9048 ( .A1(n7827), .A2(n7823), .ZN(n7824) );
  NAND2_X1 U9049 ( .A1(n7825), .A2(n7824), .ZN(n7918) );
  OR2_X1 U9050 ( .A1(n7922), .A2(n7919), .ZN(n8490) );
  NAND2_X1 U9051 ( .A1(n7919), .A2(n7922), .ZN(n8495) );
  NAND2_X1 U9052 ( .A1(n8490), .A2(n8495), .ZN(n8749) );
  XOR2_X1 U9053 ( .A(n7918), .B(n8749), .Z(n7826) );
  OAI222_X1 U9054 ( .A1(n9291), .A2(n7827), .B1(n9289), .B2(n8081), .C1(n9287), 
        .C2(n7826), .ZN(n7909) );
  AOI21_X1 U9055 ( .B1(n11086), .B2(n7828), .A(n7909), .ZN(n7832) );
  AOI22_X1 U9056 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n9352), .B1(n11106), .B2(
        n7919), .ZN(n7831) );
  NAND2_X1 U9057 ( .A1(n7924), .A2(n7923), .ZN(n7829) );
  XNOR2_X1 U9058 ( .A(n7829), .B(n8749), .ZN(n7910) );
  NAND2_X1 U9059 ( .A1(n7910), .A2(n11104), .ZN(n7830) );
  OAI211_X1 U9060 ( .C1(n7832), .C2(n9352), .A(n7831), .B(n7830), .ZN(P2_U3225) );
  INV_X1 U9061 ( .A(n7833), .ZN(n7836) );
  AOI21_X1 U9062 ( .B1(n7836), .B2(n7835), .A(n7834), .ZN(n8063) );
  MUX2_X1 U9063 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8381), .Z(n7837) );
  AND2_X1 U9064 ( .A1(n7837), .A2(n8054), .ZN(n8061) );
  INV_X1 U9065 ( .A(n8061), .ZN(n7840) );
  INV_X1 U9066 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7838) );
  MUX2_X1 U9067 ( .A(n5594), .B(n7838), .S(n8381), .Z(n7839) );
  INV_X1 U9068 ( .A(n8054), .ZN(n7937) );
  NAND2_X1 U9069 ( .A1(n7839), .A2(n7937), .ZN(n8062) );
  NAND2_X1 U9070 ( .A1(n7840), .A2(n8062), .ZN(n7841) );
  XNOR2_X1 U9071 ( .A(n8063), .B(n7841), .ZN(n7862) );
  INV_X1 U9072 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U9073 ( .A1(n9166), .A2(n7937), .ZN(n7843) );
  INV_X1 U9074 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10640) );
  NOR2_X1 U9075 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10640), .ZN(n8078) );
  INV_X1 U9076 ( .A(n8078), .ZN(n7842) );
  OAI211_X1 U9077 ( .C1(n7844), .C2(n9158), .A(n7843), .B(n7842), .ZN(n7861)
         );
  NOR2_X1 U9078 ( .A1(n7852), .A2(n7845), .ZN(n7847) );
  NAND2_X1 U9079 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n8054), .ZN(n7848) );
  OAI21_X1 U9080 ( .B1(n8054), .B2(P2_REG1_REG_10__SCAN_IN), .A(n7848), .ZN(
        n7849) );
  AOI21_X1 U9081 ( .B1(n7850), .B2(n7849), .A(n8053), .ZN(n7859) );
  NOR2_X1 U9082 ( .A1(n7852), .A2(n7851), .ZN(n7854) );
  NAND2_X1 U9083 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n8054), .ZN(n7855) );
  OAI21_X1 U9084 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n8054), .A(n7855), .ZN(
        n7856) );
  AOI21_X1 U9085 ( .B1(n7857), .B2(n7856), .A(n8051), .ZN(n7858) );
  OAI22_X1 U9086 ( .A1(n7859), .A2(n10346), .B1(n7858), .B2(n10348), .ZN(n7860) );
  AOI211_X1 U9087 ( .C1(n10352), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7863)
         );
  INV_X1 U9088 ( .A(n7863), .ZN(P2_U3192) );
  NOR2_X1 U9089 ( .A1(n7898), .A2(n7902), .ZN(n9676) );
  AND2_X1 U9090 ( .A1(n7898), .A2(n7902), .ZN(n9684) );
  NOR2_X1 U9091 ( .A1(n9676), .A2(n9684), .ZN(n7899) );
  XNOR2_X1 U9092 ( .A(n7897), .B(n7899), .ZN(n11091) );
  INV_X1 U9093 ( .A(n9672), .ZN(n9680) );
  NOR2_X1 U9094 ( .A1(n7900), .A2(n9680), .ZN(n7867) );
  INV_X1 U9095 ( .A(n7899), .ZN(n9806) );
  XNOR2_X1 U9096 ( .A(n7867), .B(n9806), .ZN(n7869) );
  INV_X1 U9097 ( .A(n9902), .ZN(n8040) );
  OAI22_X1 U9098 ( .A1(n8040), .A2(n11008), .B1(n7966), .B2(n11010), .ZN(n7868) );
  AOI21_X1 U9099 ( .B1(n7869), .B2(n10972), .A(n7868), .ZN(n7870) );
  OAI21_X1 U9100 ( .B1(n11091), .B2(n10905), .A(n7870), .ZN(n11094) );
  NAND2_X1 U9101 ( .A1(n11094), .A2(n10218), .ZN(n7878) );
  INV_X1 U9102 ( .A(n7871), .ZN(n7965) );
  OAI22_X1 U9103 ( .A1(n10218), .A2(n7872), .B1(n7965), .B2(n10227), .ZN(n7876) );
  INV_X1 U9104 ( .A(n7873), .ZN(n7874) );
  INV_X1 U9105 ( .A(n7898), .ZN(n11093) );
  OAI211_X1 U9106 ( .C1(n7874), .C2(n11093), .A(n11006), .B(n7903), .ZN(n11092) );
  NOR2_X1 U9107 ( .A1(n11092), .A2(n10231), .ZN(n7875) );
  AOI211_X1 U9108 ( .C1(n10235), .C2(n7898), .A(n7876), .B(n7875), .ZN(n7877)
         );
  OAI211_X1 U9109 ( .C1(n11091), .C2(n10923), .A(n7878), .B(n7877), .ZN(
        P1_U3282) );
  NOR2_X1 U9110 ( .A1(n7886), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7879) );
  AOI21_X1 U9111 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7886), .A(n7879), .ZN(
        n10845) );
  NAND2_X1 U9112 ( .A1(n10845), .A2(n10844), .ZN(n10843) );
  AOI22_X1 U9113 ( .A1(n8093), .A2(n8045), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n7894), .ZN(n7882) );
  AOI211_X1 U9114 ( .C1(n7883), .C2(n7882), .A(n8092), .B(n10862), .ZN(n7896)
         );
  INV_X1 U9115 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7988) );
  AOI22_X1 U9116 ( .A1(n7886), .A2(n7988), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n10850), .ZN(n10848) );
  OAI21_X1 U9117 ( .B1(n7885), .B2(n7481), .A(n7884), .ZN(n10847) );
  NOR2_X1 U9118 ( .A1(n10848), .A2(n10847), .ZN(n10846) );
  NOR2_X1 U9119 ( .A1(n7886), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7887) );
  NOR2_X1 U9120 ( .A1(n10846), .A2(n7887), .ZN(n7890) );
  INV_X1 U9121 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11117) );
  NAND2_X1 U9122 ( .A1(n7894), .A2(n11117), .ZN(n7888) );
  NAND2_X1 U9123 ( .A1(n8093), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8086) );
  AND2_X1 U9124 ( .A1(n7888), .A2(n8086), .ZN(n7889) );
  NAND2_X1 U9125 ( .A1(n7889), .A2(n7890), .ZN(n8085) );
  OAI211_X1 U9126 ( .C1(n7890), .C2(n7889), .A(n10871), .B(n8085), .ZN(n7893)
         );
  NAND2_X1 U9127 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n8212) );
  INV_X1 U9128 ( .A(n8212), .ZN(n7891) );
  AOI21_X1 U9129 ( .B1(n10861), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7891), .ZN(
        n7892) );
  OAI211_X1 U9130 ( .C1(n10849), .C2(n7894), .A(n7893), .B(n7892), .ZN(n7895)
         );
  OR2_X1 U9131 ( .A1(n7896), .A2(n7895), .ZN(P1_U3256) );
  NAND2_X1 U9132 ( .A1(n8043), .A2(n8040), .ZN(n9687) );
  XNOR2_X1 U9133 ( .A(n8039), .B(n9795), .ZN(n7986) );
  INV_X1 U9134 ( .A(n9901), .ZN(n8272) );
  XNOR2_X1 U9135 ( .A(n8035), .B(n9795), .ZN(n7901) );
  OAI222_X1 U9136 ( .A1(n11008), .A2(n8272), .B1(n11010), .B2(n7902), .C1(
        n11016), .C2(n7901), .ZN(n7983) );
  INV_X1 U9137 ( .A(n8043), .ZN(n8041) );
  AOI211_X1 U9138 ( .C1(n8043), .C2(n7903), .A(n11042), .B(n8046), .ZN(n7984)
         );
  NAND2_X1 U9139 ( .A1(n7984), .A2(n11035), .ZN(n7905) );
  AOI22_X1 U9140 ( .A1(n10180), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8030), .B2(
        n11026), .ZN(n7904) );
  OAI211_X1 U9141 ( .C1(n8041), .C2(n11031), .A(n7905), .B(n7904), .ZN(n7906)
         );
  AOI21_X1 U9142 ( .B1(n7983), .B2(n10218), .A(n7906), .ZN(n7907) );
  OAI21_X1 U9143 ( .B1(n7986), .B2(n10220), .A(n7907), .ZN(P1_U3281) );
  INV_X1 U9144 ( .A(n8594), .ZN(n7933) );
  OAI222_X1 U9145 ( .A1(n10340), .A2(n7933), .B1(n7908), .B2(P1_U3086), .C1(
        n10694), .C2(n10337), .ZN(P1_U3335) );
  AOI21_X1 U9146 ( .B1(n11119), .B2(n7910), .A(n7909), .ZN(n7917) );
  INV_X1 U9147 ( .A(n9503), .ZN(n8022) );
  INV_X1 U9148 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7911) );
  NOR2_X1 U9149 ( .A1(n11131), .A2(n7911), .ZN(n7912) );
  AOI21_X1 U9150 ( .B1(n8022), .B2(n7919), .A(n7912), .ZN(n7913) );
  OAI21_X1 U9151 ( .B1(n7917), .B2(n11128), .A(n7913), .ZN(P2_U3414) );
  INV_X1 U9152 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7914) );
  NOR2_X1 U9153 ( .A1(n11127), .A2(n7914), .ZN(n7915) );
  AOI21_X1 U9154 ( .B1(n8018), .B2(n7919), .A(n7915), .ZN(n7916) );
  OAI21_X1 U9155 ( .B1(n7917), .B2(n11126), .A(n7916), .ZN(P2_U3467) );
  INV_X1 U9156 ( .A(n9064), .ZN(n7940) );
  OR2_X2 U9157 ( .A1(n7976), .A2(n8081), .ZN(n8506) );
  NAND2_X1 U9158 ( .A1(n7976), .A2(n8081), .ZN(n8496) );
  OR2_X1 U9159 ( .A1(n9066), .A2(n7919), .ZN(n7920) );
  XOR2_X1 U9160 ( .A(n8751), .B(n7935), .Z(n7921) );
  OAI222_X1 U9161 ( .A1(n9291), .A2(n7922), .B1(n9289), .B2(n7940), .C1(n9287), 
        .C2(n7921), .ZN(n7971) );
  INV_X1 U9162 ( .A(n7971), .ZN(n7931) );
  AND2_X1 U9163 ( .A1(n8490), .A2(n7923), .ZN(n8507) );
  NAND2_X1 U9164 ( .A1(n7952), .A2(n8495), .ZN(n7925) );
  XOR2_X1 U9165 ( .A(n8751), .B(n7925), .Z(n7972) );
  INV_X1 U9166 ( .A(n7976), .ZN(n7928) );
  AOI22_X1 U9167 ( .A1(n9352), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7926), .B2(
        n11086), .ZN(n7927) );
  OAI21_X1 U9168 ( .B1(n7928), .B2(n9354), .A(n7927), .ZN(n7929) );
  AOI21_X1 U9169 ( .B1(n7972), .B2(n11104), .A(n7929), .ZN(n7930) );
  OAI21_X1 U9170 ( .B1(n7931), .B2(n9352), .A(n7930), .ZN(P2_U3224) );
  OAI222_X1 U9171 ( .A1(n9516), .A2(n7934), .B1(n9518), .B2(n7933), .C1(n7932), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  NAND2_X1 U9172 ( .A1(n7936), .A2(n8689), .ZN(n7939) );
  AOI22_X1 U9173 ( .A1(n8392), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8578), .B2(
        n7937), .ZN(n7938) );
  NAND2_X1 U9174 ( .A1(n7939), .A2(n7938), .ZN(n11060) );
  OR2_X1 U9175 ( .A1(n11060), .A2(n7940), .ZN(n8505) );
  NAND2_X1 U9176 ( .A1(n11060), .A2(n7940), .ZN(n8509) );
  NAND2_X1 U9177 ( .A1(n8505), .A2(n8509), .ZN(n8753) );
  XNOR2_X1 U9178 ( .A(n8006), .B(n8753), .ZN(n7941) );
  NAND2_X1 U9179 ( .A1(n7941), .A2(n9358), .ZN(n7949) );
  NAND2_X1 U9180 ( .A1(n7223), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7947) );
  NAND2_X1 U9181 ( .A1(n7942), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7943) );
  AND2_X1 U9182 ( .A1(n8009), .A2(n7943), .ZN(n11080) );
  INV_X1 U9183 ( .A(n11080), .ZN(n11087) );
  NAND2_X1 U9184 ( .A1(n8643), .A2(n11087), .ZN(n7946) );
  NAND2_X1 U9185 ( .A1(n7226), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U9186 ( .A1(n7194), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7944) );
  NAND4_X1 U9187 ( .A1(n7947), .A2(n7946), .A3(n7945), .A4(n7944), .ZN(n9063)
         );
  AOI22_X1 U9188 ( .A1(n7120), .A2(n9063), .B1(n9065), .B2(n9363), .ZN(n7948)
         );
  NAND2_X1 U9189 ( .A1(n7949), .A2(n7948), .ZN(n11062) );
  INV_X1 U9190 ( .A(n11062), .ZN(n7958) );
  INV_X1 U9191 ( .A(n8751), .ZN(n7950) );
  AND2_X1 U9192 ( .A1(n7950), .A2(n8495), .ZN(n7951) );
  NAND2_X1 U9193 ( .A1(n7952), .A2(n7951), .ZN(n8000) );
  NAND2_X1 U9194 ( .A1(n8000), .A2(n8506), .ZN(n7953) );
  XNOR2_X1 U9195 ( .A(n7953), .B(n8753), .ZN(n11059) );
  INV_X1 U9196 ( .A(n11060), .ZN(n7955) );
  AOI22_X1 U9197 ( .A1(n9352), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11086), .B2(
        n8077), .ZN(n7954) );
  OAI21_X1 U9198 ( .B1(n7955), .B2(n9354), .A(n7954), .ZN(n7956) );
  AOI21_X1 U9199 ( .B1(n11059), .B2(n11104), .A(n7956), .ZN(n7957) );
  OAI21_X1 U9200 ( .B1(n7958), .B2(n9352), .A(n7957), .ZN(P2_U3223) );
  INV_X1 U9201 ( .A(n8614), .ZN(n7979) );
  OAI222_X1 U9202 ( .A1(n10340), .A2(n7979), .B1(n9822), .B2(P1_U3086), .C1(
        n10485), .C2(n10337), .ZN(P1_U3334) );
  INV_X1 U9203 ( .A(n7960), .ZN(n7962) );
  NOR2_X1 U9204 ( .A1(n7962), .A2(n7961), .ZN(n7963) );
  XNOR2_X1 U9205 ( .A(n7959), .B(n7963), .ZN(n7964) );
  NAND2_X1 U9206 ( .A1(n7964), .A2(n9633), .ZN(n7970) );
  OAI22_X1 U9207 ( .A1(n7966), .A2(n9637), .B1(n9636), .B2(n7965), .ZN(n7967)
         );
  AOI211_X1 U9208 ( .C1(n9640), .C2(n9902), .A(n7968), .B(n7967), .ZN(n7969)
         );
  OAI211_X1 U9209 ( .C1(n11093), .C2(n9643), .A(n7970), .B(n7969), .ZN(
        P1_U3236) );
  AOI21_X1 U9210 ( .B1(n7972), .B2(n11119), .A(n7971), .ZN(n7978) );
  AOI22_X1 U9211 ( .A1(n7976), .A2(n8018), .B1(n11126), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7973) );
  OAI21_X1 U9212 ( .B1(n7978), .B2(n11126), .A(n7973), .ZN(P2_U3468) );
  INV_X1 U9213 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7974) );
  NOR2_X1 U9214 ( .A1(n11131), .A2(n7974), .ZN(n7975) );
  AOI21_X1 U9215 ( .B1(n8022), .B2(n7976), .A(n7975), .ZN(n7977) );
  OAI21_X1 U9216 ( .B1(n7978), .B2(n11128), .A(n7977), .ZN(P2_U3417) );
  INV_X1 U9217 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7980) );
  OAI222_X1 U9218 ( .A1(n9516), .A2(n7980), .B1(n9518), .B2(n7979), .C1(n8451), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  AND2_X2 U9219 ( .A1(n7982), .A2(n7981), .ZN(n11147) );
  INV_X1 U9220 ( .A(n11141), .ZN(n10308) );
  AOI211_X1 U9221 ( .C1(n10308), .C2(n8043), .A(n7984), .B(n7983), .ZN(n7985)
         );
  OAI21_X1 U9222 ( .B1(n7986), .B2(n10885), .A(n7985), .ZN(n7989) );
  NAND2_X1 U9223 ( .A1(n7989), .A2(n11147), .ZN(n7987) );
  OAI21_X1 U9224 ( .B1(n11147), .B2(n7988), .A(n7987), .ZN(P1_U3534) );
  NAND2_X1 U9225 ( .A1(n7989), .A2(n11150), .ZN(n7990) );
  OAI21_X1 U9226 ( .B1(n11150), .B2(n6154), .A(n7990), .ZN(P1_U3489) );
  INV_X1 U9227 ( .A(n8633), .ZN(n7993) );
  NAND2_X1 U9228 ( .A1(n9513), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7992) );
  OR2_X1 U9229 ( .A1(n7991), .A2(P2_U3151), .ZN(n8792) );
  OAI211_X1 U9230 ( .C1(n7993), .C2(n9518), .A(n7992), .B(n8792), .ZN(P2_U3272) );
  NAND2_X1 U9231 ( .A1(n8633), .A2(n7994), .ZN(n7996) );
  OR2_X1 U9232 ( .A1(n7995), .A2(P1_U3086), .ZN(n9896) );
  OAI211_X1 U9233 ( .C1(n6424), .C2(n10337), .A(n7996), .B(n9896), .ZN(
        P1_U3332) );
  INV_X1 U9234 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7998) );
  INV_X1 U9235 ( .A(n8618), .ZN(n8380) );
  OAI222_X1 U9236 ( .A1(n9516), .A2(n7998), .B1(n9518), .B2(n8380), .C1(
        P2_U3151), .C2(n7997), .ZN(P2_U3273) );
  AND2_X1 U9237 ( .A1(n8506), .A2(n8505), .ZN(n7999) );
  NAND2_X1 U9238 ( .A1(n8000), .A2(n7999), .ZN(n8001) );
  NAND2_X1 U9239 ( .A1(n8002), .A2(n8689), .ZN(n8004) );
  AOI22_X1 U9240 ( .A1(n8392), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8578), .B2(
        n8236), .ZN(n8003) );
  INV_X1 U9241 ( .A(n9063), .ZN(n8254) );
  OR2_X1 U9242 ( .A1(n11085), .A2(n8254), .ZN(n8514) );
  NAND2_X1 U9243 ( .A1(n11085), .A2(n8254), .ZN(n8512) );
  OAI21_X1 U9244 ( .B1(n8005), .B2(n8755), .A(n8134), .ZN(n11082) );
  NAND2_X1 U9245 ( .A1(n8006), .A2(n8753), .ZN(n8008) );
  OR2_X1 U9246 ( .A1(n11060), .A2(n9064), .ZN(n8007) );
  XNOR2_X1 U9247 ( .A(n8116), .B(n8755), .ZN(n8017) );
  NAND2_X1 U9248 ( .A1(n7223), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U9249 ( .A1(n8009), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U9250 ( .A1(n8108), .A2(n8010), .ZN(n11099) );
  NAND2_X1 U9251 ( .A1(n8643), .A2(n11099), .ZN(n8013) );
  NAND2_X1 U9252 ( .A1(n7226), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U9253 ( .A1(n8597), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8011) );
  NAND4_X1 U9254 ( .A1(n8014), .A2(n8013), .A3(n8012), .A4(n8011), .ZN(n9062)
         );
  NAND2_X1 U9255 ( .A1(n9062), .A2(n7120), .ZN(n8016) );
  NAND2_X1 U9256 ( .A1(n9064), .A2(n9363), .ZN(n8015) );
  AND2_X1 U9257 ( .A1(n8016), .A2(n8015), .ZN(n11068) );
  OAI21_X1 U9258 ( .B1(n8017), .B2(n9287), .A(n11068), .ZN(n11081) );
  AOI21_X1 U9259 ( .B1(n11119), .B2(n11082), .A(n11081), .ZN(n8024) );
  AOI22_X1 U9260 ( .A1(n11085), .A2(n8018), .B1(n11126), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n8019) );
  OAI21_X1 U9261 ( .B1(n8024), .B2(n11126), .A(n8019), .ZN(P2_U3470) );
  INV_X1 U9262 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8020) );
  NOR2_X1 U9263 ( .A1(n11131), .A2(n8020), .ZN(n8021) );
  AOI21_X1 U9264 ( .B1(n11085), .B2(n8022), .A(n8021), .ZN(n8023) );
  OAI21_X1 U9265 ( .B1(n8024), .B2(n11128), .A(n8023), .ZN(P2_U3423) );
  INV_X1 U9266 ( .A(n8026), .ZN(n8027) );
  AOI21_X1 U9267 ( .B1(n8029), .B2(n8028), .A(n8027), .ZN(n8034) );
  AOI22_X1 U9268 ( .A1(n9623), .A2(n9903), .B1(n9624), .B2(n8030), .ZN(n8031)
         );
  NAND2_X1 U9269 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n10856) );
  OAI211_X1 U9270 ( .C1(n8272), .C2(n9605), .A(n8031), .B(n10856), .ZN(n8032)
         );
  AOI21_X1 U9271 ( .B1(n8043), .B2(n9625), .A(n8032), .ZN(n8033) );
  OAI21_X1 U9272 ( .B1(n8034), .B2(n9616), .A(n8033), .ZN(P1_U3224) );
  AND2_X1 U9273 ( .A1(n8036), .A2(n9693), .ZN(n8037) );
  OR2_X1 U9274 ( .A1(n8220), .A2(n8272), .ZN(n9860) );
  NAND2_X1 U9275 ( .A1(n8220), .A2(n8272), .ZN(n9694) );
  NAND3_X1 U9276 ( .A1(n8036), .A2(n9810), .A3(n9693), .ZN(n8156) );
  OAI21_X1 U9277 ( .B1(n8037), .B2(n9810), .A(n8156), .ZN(n8038) );
  AOI222_X1 U9278 ( .A1(n10972), .A2(n8038), .B1(n9900), .B2(n10969), .C1(
        n9902), .C2(n10967), .ZN(n11113) );
  XOR2_X1 U9279 ( .A(n8155), .B(n9810), .Z(n11116) );
  NAND2_X1 U9280 ( .A1(n11116), .A2(n10982), .ZN(n8050) );
  INV_X1 U9281 ( .A(n8211), .ZN(n8044) );
  OAI22_X1 U9282 ( .A1(n10218), .A2(n8045), .B1(n8044), .B2(n10227), .ZN(n8048) );
  INV_X1 U9283 ( .A(n8159), .ZN(n8277) );
  OAI211_X1 U9284 ( .C1(n11114), .C2(n8046), .A(n8277), .B(n11006), .ZN(n11112) );
  NOR2_X1 U9285 ( .A1(n11112), .A2(n10231), .ZN(n8047) );
  AOI211_X1 U9286 ( .C1(n10235), .C2(n8220), .A(n8048), .B(n8047), .ZN(n8049)
         );
  OAI211_X1 U9287 ( .C1(n11028), .C2(n11113), .A(n8050), .B(n8049), .ZN(
        P1_U3280) );
  INV_X1 U9288 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11090) );
  AOI21_X1 U9289 ( .B1(n11090), .B2(n8052), .A(n8237), .ZN(n8069) );
  INV_X1 U9290 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8055) );
  AOI21_X1 U9291 ( .B1(n8056), .B2(n8055), .A(n8224), .ZN(n8057) );
  INV_X1 U9292 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10572) );
  OR2_X1 U9293 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10572), .ZN(n11066) );
  OAI21_X1 U9294 ( .B1(n10346), .B2(n8057), .A(n11066), .ZN(n8060) );
  INV_X1 U9295 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8058) );
  NOR2_X1 U9296 ( .A1(n9158), .A2(n8058), .ZN(n8059) );
  AOI211_X1 U9297 ( .C1(n9166), .C2(n8236), .A(n8060), .B(n8059), .ZN(n8068)
         );
  AOI21_X1 U9298 ( .B1(n8063), .B2(n8062), .A(n8061), .ZN(n8065) );
  MUX2_X1 U9299 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8381), .Z(n8226) );
  XNOR2_X1 U9300 ( .A(n8226), .B(n8236), .ZN(n8064) );
  NAND2_X1 U9301 ( .A1(n8065), .A2(n8064), .ZN(n8227) );
  OAI21_X1 U9302 ( .B1(n8065), .B2(n8064), .A(n8227), .ZN(n8066) );
  NAND2_X1 U9303 ( .A1(n8066), .A2(n10352), .ZN(n8067) );
  OAI211_X1 U9304 ( .C1(n8069), .C2(n10348), .A(n8068), .B(n8067), .ZN(
        P2_U3193) );
  INV_X1 U9305 ( .A(n8070), .ZN(n8071) );
  XNOR2_X1 U9306 ( .A(n11060), .B(n5099), .ZN(n8074) );
  OAI21_X1 U9307 ( .B1(n8075), .B2(n8074), .A(n8246), .ZN(n8076) );
  NOR2_X1 U9308 ( .A1(n8076), .A2(n9064), .ZN(n11071) );
  AOI21_X1 U9309 ( .B1(n9064), .B2(n8076), .A(n11071), .ZN(n8084) );
  NAND2_X1 U9310 ( .A1(n9053), .A2(n8077), .ZN(n8080) );
  AOI21_X1 U9311 ( .B1(n9034), .B2(n9063), .A(n8078), .ZN(n8079) );
  OAI211_X1 U9312 ( .C1(n8081), .C2(n9037), .A(n8080), .B(n8079), .ZN(n8082)
         );
  AOI21_X1 U9313 ( .B1(n11060), .B2(n11077), .A(n8082), .ZN(n8083) );
  OAI21_X1 U9314 ( .B1(n8084), .B2(n11072), .A(n8083), .ZN(P2_U3157) );
  NAND2_X1 U9315 ( .A1(n8086), .A2(n8085), .ZN(n8091) );
  NAND2_X1 U9316 ( .A1(n8103), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8087) );
  OAI21_X1 U9317 ( .B1(n8103), .B2(P1_REG1_REG_14__SCAN_IN), .A(n8087), .ZN(
        n8090) );
  INV_X1 U9318 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U9319 ( .A1(n8103), .A2(n8089), .ZN(n8088) );
  OAI211_X1 U9320 ( .C1(n8089), .C2(n8103), .A(n8088), .B(n8091), .ZN(n8149)
         );
  OAI211_X1 U9321 ( .C1(n8091), .C2(n8090), .A(n10871), .B(n8149), .ZN(n8102)
         );
  NAND2_X1 U9322 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n8206) );
  INV_X1 U9323 ( .A(n8206), .ZN(n8100) );
  NAND2_X1 U9324 ( .A1(n8103), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8094) );
  OAI21_X1 U9325 ( .B1(n8103), .B2(P1_REG2_REG_14__SCAN_IN), .A(n8094), .ZN(
        n8095) );
  INV_X1 U9326 ( .A(n8095), .ZN(n8097) );
  INV_X1 U9327 ( .A(n8142), .ZN(n8096) );
  AOI211_X1 U9328 ( .C1(n8098), .C2(n8097), .A(n8096), .B(n10862), .ZN(n8099)
         );
  AOI211_X1 U9329 ( .C1(n10861), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n8100), .B(
        n8099), .ZN(n8101) );
  OAI211_X1 U9330 ( .C1(n10849), .C2(n8103), .A(n8102), .B(n8101), .ZN(
        P1_U3257) );
  INV_X1 U9331 ( .A(n8436), .ZN(n8105) );
  OAI222_X1 U9332 ( .A1(n9516), .A2(n8106), .B1(n9518), .B2(n8105), .C1(n8104), 
        .C2(P2_U3151), .ZN(P2_U3270) );
  INV_X1 U9333 ( .A(n8107), .ZN(n8125) );
  NAND2_X1 U9334 ( .A1(n8108), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U9335 ( .A1(n8125), .A2(n8109), .ZN(n9004) );
  NAND2_X1 U9336 ( .A1(n8111), .A2(n8689), .ZN(n8113) );
  AOI22_X1 U9337 ( .A1(n8392), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8578), .B2(
        n9087), .ZN(n8112) );
  NAND2_X1 U9338 ( .A1(n8113), .A2(n8112), .ZN(n11122) );
  INV_X1 U9339 ( .A(n11122), .ZN(n8174) );
  NOR2_X1 U9340 ( .A1(n8174), .A2(n9233), .ZN(n8133) );
  NOR2_X1 U9341 ( .A1(n11085), .A2(n9063), .ZN(n8115) );
  NAND2_X1 U9342 ( .A1(n11085), .A2(n9063), .ZN(n8114) );
  NAND2_X1 U9343 ( .A1(n8117), .A2(n8689), .ZN(n8119) );
  AOI22_X1 U9344 ( .A1(n8392), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8578), .B2(
        n8323), .ZN(n8118) );
  XNOR2_X1 U9345 ( .A(n11107), .B(n9007), .ZN(n8758) );
  NAND2_X1 U9346 ( .A1(n8540), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U9347 ( .A1(n8187), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8122) );
  NAND2_X1 U9348 ( .A1(n8643), .A2(n9004), .ZN(n8121) );
  NAND2_X1 U9349 ( .A1(n8597), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8120) );
  OR2_X1 U9350 ( .A1(n11122), .A2(n8803), .ZN(n8527) );
  AND2_X1 U9351 ( .A1(n11122), .A2(n8803), .ZN(n8525) );
  OR2_X1 U9352 ( .A1(n5432), .A2(n8525), .ZN(n8759) );
  INV_X1 U9353 ( .A(n8759), .ZN(n8137) );
  XNOR2_X1 U9354 ( .A(n8176), .B(n8137), .ZN(n8124) );
  NAND2_X1 U9355 ( .A1(n8124), .A2(n9358), .ZN(n8132) );
  NAND2_X1 U9356 ( .A1(n8540), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8130) );
  NAND2_X1 U9357 ( .A1(n8125), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U9358 ( .A1(n8185), .A2(n8126), .ZN(n8195) );
  NAND2_X1 U9359 ( .A1(n8643), .A2(n8195), .ZN(n8129) );
  NAND2_X1 U9360 ( .A1(n7226), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U9361 ( .A1(n8597), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8127) );
  NAND4_X1 U9362 ( .A1(n8130), .A2(n8129), .A3(n8128), .A4(n8127), .ZN(n9362)
         );
  AOI22_X1 U9363 ( .A1(n9363), .A2(n9062), .B1(n9362), .B2(n7120), .ZN(n8131)
         );
  NAND2_X1 U9364 ( .A1(n8132), .A2(n8131), .ZN(n11124) );
  AOI211_X1 U9365 ( .C1(n11086), .C2(n9004), .A(n8133), .B(n11124), .ZN(n8139)
         );
  NAND2_X1 U9366 ( .A1(n11107), .A2(n9007), .ZN(n8136) );
  XNOR2_X1 U9367 ( .A(n8197), .B(n8137), .ZN(n11120) );
  AOI22_X1 U9368 ( .A1(n11120), .A2(n11104), .B1(P2_REG2_REG_13__SCAN_IN), 
        .B2(n9352), .ZN(n8138) );
  OAI21_X1 U9369 ( .B1(n8139), .B2(n9352), .A(n8138), .ZN(P2_U3220) );
  INV_X1 U9370 ( .A(n8636), .ZN(n8798) );
  OAI222_X1 U9371 ( .A1(n10337), .A2(n10688), .B1(P1_U3086), .B2(n8140), .C1(
        n10340), .C2(n8798), .ZN(P1_U3331) );
  NAND2_X1 U9372 ( .A1(n8147), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U9373 ( .A1(n8142), .A2(n8141), .ZN(n8144) );
  INV_X1 U9374 ( .A(n9922), .ZN(n8143) );
  OAI21_X1 U9375 ( .B1(n9911), .B2(n8144), .A(n8143), .ZN(n8145) );
  NOR2_X1 U9376 ( .A1(n6235), .A2(n8145), .ZN(n9921) );
  AOI211_X1 U9377 ( .C1(n6235), .C2(n8145), .A(n9921), .B(n10862), .ZN(n8146)
         );
  INV_X1 U9378 ( .A(n8146), .ZN(n8153) );
  AND2_X1 U9379 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U9380 ( .A1(n8147), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U9381 ( .A1(n8149), .A2(n8148), .ZN(n9912) );
  XNOR2_X1 U9382 ( .A(n9912), .B(n8154), .ZN(n9914) );
  XNOR2_X1 U9383 ( .A(n9914), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n8150) );
  NOR2_X1 U9384 ( .A1(n10851), .A2(n8150), .ZN(n8151) );
  AOI211_X1 U9385 ( .C1(n10861), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n9639), .B(
        n8151), .ZN(n8152) );
  OAI211_X1 U9386 ( .C1(n10849), .C2(n8154), .A(n8153), .B(n8152), .ZN(
        P1_U3258) );
  XNOR2_X1 U9387 ( .A(n10307), .B(n9900), .ZN(n9808) );
  INV_X1 U9388 ( .A(n10307), .ZN(n8280) );
  INV_X1 U9389 ( .A(n9900), .ZN(n9688) );
  NAND2_X1 U9390 ( .A1(n8259), .A2(n8271), .ZN(n9701) );
  NAND2_X1 U9391 ( .A1(n9700), .A2(n9701), .ZN(n8260) );
  INV_X1 U9392 ( .A(n8260), .ZN(n9811) );
  XNOR2_X1 U9393 ( .A(n8261), .B(n9811), .ZN(n11136) );
  INV_X1 U9394 ( .A(n11136), .ZN(n8164) );
  AOI22_X1 U9395 ( .A1(n8259), .A2(n10235), .B1(P1_REG2_REG_15__SCAN_IN), .B2(
        n11028), .ZN(n8163) );
  NAND2_X1 U9396 ( .A1(n8156), .A2(n9694), .ZN(n8270) );
  INV_X1 U9397 ( .A(n9808), .ZN(n8157) );
  OR2_X1 U9398 ( .A1(n10307), .A2(n9688), .ZN(n9689) );
  XNOR2_X1 U9399 ( .A(n8264), .B(n8260), .ZN(n8158) );
  AOI222_X1 U9400 ( .A1(n10972), .A2(n8158), .B1(n10222), .B2(n10969), .C1(
        n9900), .C2(n10967), .ZN(n11133) );
  INV_X1 U9401 ( .A(n11133), .ZN(n8161) );
  OAI211_X1 U9402 ( .C1(n5180), .C2(n11134), .A(n8262), .B(n11006), .ZN(n11132) );
  OAI22_X1 U9403 ( .A1(n11132), .A2(n6328), .B1(n9635), .B2(n10227), .ZN(n8160) );
  OAI21_X1 U9404 ( .B1(n8161), .B2(n8160), .A(n10218), .ZN(n8162) );
  OAI211_X1 U9405 ( .C1(n8164), .C2(n10220), .A(n8163), .B(n8162), .ZN(
        P1_U3278) );
  INV_X1 U9406 ( .A(n11107), .ZN(n8258) );
  INV_X1 U9407 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8169) );
  NAND3_X1 U9408 ( .A1(n8134), .A2(n8758), .A3(n8512), .ZN(n8165) );
  NAND2_X1 U9409 ( .A1(n8166), .A2(n8165), .ZN(n11105) );
  XNOR2_X1 U9410 ( .A(n8167), .B(n8758), .ZN(n8168) );
  OAI222_X1 U9411 ( .A1(n9289), .A2(n8803), .B1(n9291), .B2(n8254), .C1(n9287), 
        .C2(n8168), .ZN(n11100) );
  AOI21_X1 U9412 ( .B1(n11119), .B2(n11105), .A(n11100), .ZN(n8171) );
  MUX2_X1 U9413 ( .A(n8169), .B(n8171), .S(n11127), .Z(n8170) );
  OAI21_X1 U9414 ( .B1(n8258), .B2(n9445), .A(n8170), .ZN(P2_U3471) );
  INV_X1 U9415 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8172) );
  MUX2_X1 U9416 ( .A(n8172), .B(n8171), .S(n11131), .Z(n8173) );
  OAI21_X1 U9417 ( .B1(n8258), .B2(n9503), .A(n8173), .ZN(P2_U3426) );
  INV_X1 U9418 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8201) );
  INV_X1 U9419 ( .A(n8803), .ZN(n9061) );
  NAND2_X1 U9420 ( .A1(n8175), .A2(n8174), .ZN(n8178) );
  NAND2_X1 U9421 ( .A1(n8179), .A2(n8689), .ZN(n8181) );
  INV_X1 U9422 ( .A(n8330), .ZN(n9104) );
  AOI22_X1 U9423 ( .A1(n8392), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8578), .B2(
        n9104), .ZN(n8180) );
  XNOR2_X1 U9424 ( .A(n8916), .B(n9362), .ZN(n8760) );
  INV_X1 U9425 ( .A(n8760), .ZN(n8182) );
  NAND2_X1 U9426 ( .A1(n8183), .A2(n8760), .ZN(n8184) );
  NAND3_X1 U9427 ( .A1(n8856), .A2(n9358), .A3(n8184), .ZN(n8194) );
  NAND2_X1 U9428 ( .A1(n8540), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U9429 ( .A1(n8185), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U9430 ( .A1(n8542), .A2(n8186), .ZN(n9366) );
  NAND2_X1 U9431 ( .A1(n8643), .A2(n9366), .ZN(n8190) );
  INV_X1 U9432 ( .A(n7044), .ZN(n8187) );
  NAND2_X1 U9433 ( .A1(n7226), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U9434 ( .A1(n7194), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8188) );
  NAND4_X1 U9435 ( .A1(n8191), .A2(n8190), .A3(n8189), .A4(n8188), .ZN(n9060)
         );
  NAND2_X1 U9436 ( .A1(n9060), .A2(n7120), .ZN(n8192) );
  OAI21_X1 U9437 ( .B1(n8803), .B2(n9291), .A(n8192), .ZN(n8912) );
  INV_X1 U9438 ( .A(n8912), .ZN(n8193) );
  NAND2_X1 U9439 ( .A1(n8194), .A2(n8193), .ZN(n9450) );
  INV_X1 U9440 ( .A(n8916), .ZN(n9448) );
  INV_X1 U9441 ( .A(n8195), .ZN(n8914) );
  OAI22_X1 U9442 ( .A1(n9448), .A2(n9233), .B1(n8914), .B2(n11102), .ZN(n8196)
         );
  OAI21_X1 U9443 ( .B1(n9450), .B2(n8196), .A(n11111), .ZN(n8200) );
  OR2_X1 U9444 ( .A1(n8198), .A2(n8760), .ZN(n9446) );
  NAND3_X1 U9445 ( .A1(n9446), .A2(n8701), .A3(n11104), .ZN(n8199) );
  OAI211_X1 U9446 ( .C1(n11111), .C2(n8201), .A(n8200), .B(n8199), .ZN(
        P2_U3219) );
  NAND2_X1 U9447 ( .A1(n8203), .A2(n8202), .ZN(n8205) );
  XNOR2_X1 U9448 ( .A(n8205), .B(n8204), .ZN(n8210) );
  AOI22_X1 U9449 ( .A1(n9623), .A2(n9901), .B1(n9624), .B2(n8278), .ZN(n8207)
         );
  OAI211_X1 U9450 ( .C1(n8271), .C2(n9605), .A(n8207), .B(n8206), .ZN(n8208)
         );
  AOI21_X1 U9451 ( .B1(n10307), .B2(n9625), .A(n8208), .ZN(n8209) );
  OAI21_X1 U9452 ( .B1(n8210), .B2(n9616), .A(n8209), .ZN(P1_U3215) );
  AOI22_X1 U9453 ( .A1(n9623), .A2(n9902), .B1(n9624), .B2(n8211), .ZN(n8213)
         );
  OAI211_X1 U9454 ( .C1(n9688), .C2(n9605), .A(n8213), .B(n8212), .ZN(n8219)
         );
  INV_X1 U9455 ( .A(n8215), .ZN(n8216) );
  AOI211_X1 U9456 ( .C1(n8217), .C2(n8214), .A(n9616), .B(n8216), .ZN(n8218)
         );
  AOI211_X1 U9457 ( .C1(n8220), .C2(n9625), .A(n8219), .B(n8218), .ZN(n8221)
         );
  INV_X1 U9458 ( .A(n8221), .ZN(P1_U3234) );
  NOR2_X1 U9459 ( .A1(n8236), .A2(n8222), .ZN(n8223) );
  MUX2_X1 U9460 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8169), .S(n8323), .Z(n8225)
         );
  AOI21_X1 U9461 ( .B1(n5187), .B2(n8225), .A(n8289), .ZN(n8245) );
  INV_X1 U9462 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8234) );
  MUX2_X1 U9463 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8381), .Z(n8309) );
  XNOR2_X1 U9464 ( .A(n8309), .B(n8323), .ZN(n8230) );
  OR2_X1 U9465 ( .A1(n8226), .A2(n5591), .ZN(n8228) );
  NAND2_X1 U9466 ( .A1(n8228), .A2(n8227), .ZN(n8229) );
  NAND2_X1 U9467 ( .A1(n8230), .A2(n8229), .ZN(n8310) );
  OAI21_X1 U9468 ( .B1(n8230), .B2(n8229), .A(n8310), .ZN(n8231) );
  NAND2_X1 U9469 ( .A1(n8231), .A2(n10352), .ZN(n8233) );
  INV_X1 U9470 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10376) );
  NOR2_X1 U9471 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10376), .ZN(n8252) );
  INV_X1 U9472 ( .A(n8252), .ZN(n8232) );
  OAI211_X1 U9473 ( .C1(n8234), .C2(n9158), .A(n8233), .B(n8232), .ZN(n8243)
         );
  NOR2_X1 U9474 ( .A1(n8236), .A2(n8235), .ZN(n8238) );
  INV_X1 U9475 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U9476 ( .A1(n8323), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11110), .B2(
        n8308), .ZN(n8239) );
  AOI21_X1 U9477 ( .B1(n8240), .B2(n8239), .A(n8325), .ZN(n8241) );
  NOR2_X1 U9478 ( .A1(n8241), .A2(n10348), .ZN(n8242) );
  AOI211_X1 U9479 ( .C1(n9166), .C2(n8323), .A(n8243), .B(n8242), .ZN(n8244)
         );
  OAI21_X1 U9480 ( .B1(n8245), .B2(n10346), .A(n8244), .ZN(P2_U3194) );
  XNOR2_X1 U9481 ( .A(n11085), .B(n5099), .ZN(n8247) );
  INV_X1 U9482 ( .A(n8247), .ZN(n8248) );
  INV_X1 U9483 ( .A(n8246), .ZN(n11070) );
  XNOR2_X1 U9484 ( .A(n8247), .B(n9063), .ZN(n11069) );
  OAI21_X1 U9485 ( .B1(n8248), .B2(n9063), .A(n11074), .ZN(n8250) );
  XNOR2_X1 U9486 ( .A(n11107), .B(n5099), .ZN(n8800) );
  XOR2_X1 U9487 ( .A(n9062), .B(n8800), .Z(n8249) );
  AOI21_X1 U9488 ( .B1(n8250), .B2(n8249), .A(n11072), .ZN(n8251) );
  NAND2_X1 U9489 ( .A1(n8251), .A2(n8802), .ZN(n8257) );
  AOI21_X1 U9490 ( .B1(n9061), .B2(n9034), .A(n8252), .ZN(n8253) );
  OAI21_X1 U9491 ( .B1(n8254), .B2(n9037), .A(n8253), .ZN(n8255) );
  AOI21_X1 U9492 ( .B1(n11099), .B2(n9053), .A(n8255), .ZN(n8256) );
  OAI211_X1 U9493 ( .C1(n8258), .C2(n9056), .A(n8257), .B(n8256), .ZN(P2_U3164) );
  INV_X1 U9494 ( .A(n10222), .ZN(n10013) );
  OR2_X1 U9495 ( .A1(n10303), .A2(n10013), .ZN(n9868) );
  NAND2_X1 U9496 ( .A1(n10303), .A2(n10013), .ZN(n9864) );
  XNOR2_X1 U9497 ( .A(n10015), .B(n10014), .ZN(n10306) );
  AOI211_X1 U9498 ( .C1(n10303), .C2(n8262), .A(n11042), .B(n5181), .ZN(n10302) );
  INV_X1 U9499 ( .A(n10303), .ZN(n10012) );
  AOI22_X1 U9500 ( .A1(n10180), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n11026), 
        .B2(n9566), .ZN(n8263) );
  OAI21_X1 U9501 ( .B1(n10012), .B2(n11031), .A(n8263), .ZN(n8268) );
  OAI21_X1 U9502 ( .B1(n8265), .B2(n10014), .A(n9758), .ZN(n8266) );
  AOI222_X1 U9503 ( .A1(n10972), .A2(n8266), .B1(n10016), .B2(n10969), .C1(
        n9899), .C2(n10967), .ZN(n10305) );
  NOR2_X1 U9504 ( .A1(n10305), .A2(n10180), .ZN(n8267) );
  AOI211_X1 U9505 ( .C1(n10302), .C2(n11035), .A(n8268), .B(n8267), .ZN(n8269)
         );
  OAI21_X1 U9506 ( .B1(n10306), .B2(n10220), .A(n8269), .ZN(P1_U3277) );
  XNOR2_X1 U9507 ( .A(n8270), .B(n9808), .ZN(n8276) );
  OAI22_X1 U9508 ( .A1(n8272), .A2(n11010), .B1(n8271), .B2(n11008), .ZN(n8275) );
  XNOR2_X1 U9509 ( .A(n8273), .B(n9808), .ZN(n10312) );
  NOR2_X1 U9510 ( .A1(n10312), .A2(n10905), .ZN(n8274) );
  AOI211_X1 U9511 ( .C1(n10972), .C2(n8276), .A(n8275), .B(n8274), .ZN(n10311)
         );
  AOI21_X1 U9512 ( .B1(n10307), .B2(n8277), .A(n5180), .ZN(n10309) );
  AOI22_X1 U9513 ( .A1(n10180), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8278), .B2(
        n11026), .ZN(n8279) );
  OAI21_X1 U9514 ( .B1(n8280), .B2(n11031), .A(n8279), .ZN(n8282) );
  NOR2_X1 U9515 ( .A1(n10312), .A2(n10923), .ZN(n8281) );
  AOI211_X1 U9516 ( .C1(n10309), .C2(n10153), .A(n8282), .B(n8281), .ZN(n8283)
         );
  OAI21_X1 U9517 ( .B1(n10311), .B2(n10180), .A(n8283), .ZN(P1_U3279) );
  INV_X1 U9518 ( .A(n8426), .ZN(n8284) );
  OAI222_X1 U9519 ( .A1(n10337), .A2(n10685), .B1(n10340), .B2(n8284), .C1(
        n6576), .C2(P1_U3086), .ZN(P1_U3329) );
  OAI222_X1 U9520 ( .A1(P2_U3151), .A2(n8285), .B1(n9518), .B2(n8284), .C1(
        n9516), .C2(n6507), .ZN(P2_U3269) );
  INV_X1 U9521 ( .A(n8416), .ZN(n8382) );
  OAI222_X1 U9522 ( .A1(n10337), .A2(n10570), .B1(n10340), .B2(n8382), .C1(
        P1_U3086), .C2(n10823), .ZN(P1_U3328) );
  INV_X1 U9523 ( .A(n8406), .ZN(n10339) );
  AOI21_X1 U9524 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9513), .A(n8286), .ZN(
        n8287) );
  OAI21_X1 U9525 ( .B1(n10339), .B2(n9518), .A(n8287), .ZN(P2_U3267) );
  AND2_X1 U9526 ( .A1(n8288), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U9527 ( .A1(n8288), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U9528 ( .A1(n8288), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U9529 ( .A1(n8288), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U9530 ( .A1(n8288), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U9531 ( .A1(n8288), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U9532 ( .A1(n8288), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U9533 ( .A1(n8288), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U9534 ( .A1(n8288), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U9535 ( .A1(n8288), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U9536 ( .A1(n8288), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U9537 ( .A1(n8288), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U9538 ( .A1(n8288), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U9539 ( .A1(n8288), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U9540 ( .A1(n8288), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U9541 ( .A1(n8288), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U9542 ( .A1(n8288), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U9543 ( .A1(n8288), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U9544 ( .A1(n8288), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U9545 ( .A1(n8288), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U9546 ( .A1(n8288), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U9547 ( .A1(n8288), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U9548 ( .A1(n8288), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U9549 ( .A1(n8288), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U9550 ( .A1(n8288), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U9551 ( .A1(n8288), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U9552 ( .A1(n8288), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U9553 ( .A1(n8288), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U9554 ( .A1(n8288), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U9555 ( .A1(n8288), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  OR2_X1 U9556 ( .A1(n8323), .A2(n8169), .ZN(n8291) );
  INV_X1 U9557 ( .A(n8289), .ZN(n8290) );
  NAND2_X1 U9558 ( .A1(n8291), .A2(n8290), .ZN(n8292) );
  XNOR2_X1 U9559 ( .A(n8292), .B(n9087), .ZN(n9078) );
  NAND2_X1 U9560 ( .A1(n8292), .A2(n8326), .ZN(n8293) );
  OR2_X1 U9561 ( .A1(n8330), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U9562 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8330), .ZN(n8294) );
  NAND2_X1 U9563 ( .A1(n8295), .A2(n8294), .ZN(n9095) );
  NOR2_X1 U9564 ( .A1(n8534), .A2(n8296), .ZN(n8297) );
  INV_X1 U9565 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9443) );
  XNOR2_X1 U9566 ( .A(n8534), .B(n8296), .ZN(n9116) );
  NOR2_X1 U9567 ( .A1(n9443), .A2(n9116), .ZN(n9119) );
  INV_X1 U9568 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9438) );
  AOI22_X1 U9569 ( .A1(n9145), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9438), .B2(
        n8335), .ZN(n9140) );
  NOR2_X1 U9570 ( .A1(n9165), .A2(n8298), .ZN(n8299) );
  INV_X1 U9571 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U9572 ( .A1(n8352), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8346) );
  OAI21_X1 U9573 ( .B1(n8352), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8346), .ZN(
        n8300) );
  AOI21_X1 U9574 ( .B1(n8301), .B2(n8300), .A(n5175), .ZN(n8345) );
  MUX2_X1 U9575 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8381), .Z(n8317) );
  XNOR2_X1 U9576 ( .A(n8317), .B(n9165), .ZN(n9153) );
  MUX2_X1 U9577 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8381), .Z(n8302) );
  OR2_X1 U9578 ( .A1(n8302), .A2(n8335), .ZN(n8315) );
  XNOR2_X1 U9579 ( .A(n8302), .B(n9145), .ZN(n9134) );
  MUX2_X1 U9580 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8381), .Z(n8303) );
  OR2_X1 U9581 ( .A1(n8303), .A2(n9124), .ZN(n8314) );
  XNOR2_X1 U9582 ( .A(n8303), .B(n8534), .ZN(n9115) );
  MUX2_X1 U9583 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8381), .Z(n8304) );
  OR2_X1 U9584 ( .A1(n8304), .A2(n8330), .ZN(n8313) );
  XNOR2_X1 U9585 ( .A(n8304), .B(n9104), .ZN(n9098) );
  INV_X1 U9586 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8306) );
  INV_X1 U9587 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8305) );
  MUX2_X1 U9588 ( .A(n8306), .B(n8305), .S(n8381), .Z(n8307) );
  NAND2_X1 U9589 ( .A1(n8307), .A2(n9087), .ZN(n8312) );
  XNOR2_X1 U9590 ( .A(n8307), .B(n8326), .ZN(n9085) );
  OR2_X1 U9591 ( .A1(n8309), .A2(n8308), .ZN(n8311) );
  NAND2_X1 U9592 ( .A1(n8311), .A2(n8310), .ZN(n9084) );
  NAND2_X1 U9593 ( .A1(n9085), .A2(n9084), .ZN(n9083) );
  NAND2_X1 U9594 ( .A1(n8312), .A2(n9083), .ZN(n9099) );
  NAND2_X1 U9595 ( .A1(n9098), .A2(n9099), .ZN(n9097) );
  NAND2_X1 U9596 ( .A1(n8313), .A2(n9097), .ZN(n9114) );
  NAND2_X1 U9597 ( .A1(n9115), .A2(n9114), .ZN(n9113) );
  NAND2_X1 U9598 ( .A1(n8314), .A2(n9113), .ZN(n9133) );
  NAND2_X1 U9599 ( .A1(n9134), .A2(n9133), .ZN(n9132) );
  NAND2_X1 U9600 ( .A1(n8315), .A2(n9132), .ZN(n9152) );
  NAND2_X1 U9601 ( .A1(n9153), .A2(n9152), .ZN(n9151) );
  OAI21_X1 U9602 ( .B1(n8317), .B2(n8316), .A(n9151), .ZN(n8320) );
  INV_X1 U9603 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9322) );
  INV_X1 U9604 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8318) );
  MUX2_X1 U9605 ( .A(n9322), .B(n8318), .S(n8381), .Z(n8319) );
  NOR2_X1 U9606 ( .A1(n8320), .A2(n8319), .ZN(n8350) );
  INV_X1 U9607 ( .A(n8350), .ZN(n8321) );
  NAND2_X1 U9608 ( .A1(n8320), .A2(n8319), .ZN(n8351) );
  NAND2_X1 U9609 ( .A1(n8321), .A2(n8351), .ZN(n8338) );
  OAI21_X1 U9610 ( .B1(n8338), .B2(n9073), .A(n10357), .ZN(n8343) );
  INV_X1 U9611 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8322) );
  NOR2_X1 U9612 ( .A1(n9158), .A2(n8322), .ZN(n8342) );
  INV_X1 U9613 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9150) );
  NOR2_X1 U9614 ( .A1(n8323), .A2(n11110), .ZN(n8324) );
  INV_X1 U9615 ( .A(n8327), .ZN(n8328) );
  NAND2_X1 U9616 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8330), .ZN(n8329) );
  OAI21_X1 U9617 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8330), .A(n8329), .ZN(
        n9092) );
  NOR2_X1 U9618 ( .A1(n9093), .A2(n9092), .ZN(n9091) );
  NOR2_X1 U9619 ( .A1(n8534), .A2(n8332), .ZN(n8333) );
  INV_X1 U9620 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9368) );
  INV_X1 U9621 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8334) );
  AOI22_X1 U9622 ( .A1(n9145), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8334), .B2(
        n8335), .ZN(n9131) );
  XNOR2_X1 U9623 ( .A(n8336), .B(n9165), .ZN(n9149) );
  NOR2_X1 U9624 ( .A1(n9150), .A2(n9149), .ZN(n9148) );
  XOR2_X1 U9625 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n8565), .Z(n8356) );
  XOR2_X1 U9626 ( .A(n8337), .B(n8356), .Z(n8340) );
  NAND3_X1 U9627 ( .A1(n8338), .A2(n10352), .A3(n8352), .ZN(n8339) );
  NAND2_X1 U9628 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9024) );
  OAI211_X1 U9629 ( .C1(n10348), .C2(n8340), .A(n8339), .B(n9024), .ZN(n8341)
         );
  OAI21_X1 U9630 ( .B1(n8345), .B2(n10346), .A(n8344), .ZN(P2_U3200) );
  INV_X1 U9631 ( .A(n8346), .ZN(n8347) );
  XNOR2_X1 U9632 ( .A(n8779), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8349) );
  INV_X1 U9633 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8348) );
  MUX2_X1 U9634 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8348), .S(n8579), .Z(n8362)
         );
  MUX2_X1 U9635 ( .A(n8362), .B(n8349), .S(n8381), .Z(n8354) );
  AOI21_X1 U9636 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8353) );
  XOR2_X1 U9637 ( .A(n8354), .B(n8353), .Z(n8367) );
  NAND2_X1 U9638 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U9639 ( .A1(n10360), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8355) );
  OAI211_X1 U9640 ( .C1(n10357), .C2(n8779), .A(n8938), .B(n8355), .ZN(n8366)
         );
  INV_X1 U9641 ( .A(n9148), .ZN(n8357) );
  NAND2_X1 U9642 ( .A1(n8358), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8360) );
  AOI22_X1 U9643 ( .A1(n8360), .A2(n8565), .B1(n9322), .B2(n8359), .ZN(n8363)
         );
  INV_X1 U9644 ( .A(n8362), .ZN(n8361) );
  OAI21_X1 U9645 ( .B1(n8364), .B2(n8363), .A(n8361), .ZN(n8365) );
  INV_X1 U9646 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U9647 ( .A1(n8369), .A2(n9633), .ZN(n8371) );
  AOI22_X1 U9648 ( .A1(n9640), .A2(n5886), .B1(n6947), .B2(n9625), .ZN(n8370)
         );
  OAI211_X1 U9649 ( .C1(n8373), .C2(n8372), .A(n8371), .B(n8370), .ZN(P1_U3232) );
  NOR2_X1 U9650 ( .A1(n9797), .A2(n8374), .ZN(n8375) );
  AOI211_X1 U9651 ( .C1(n11026), .C2(P1_REG3_REG_0__SCAN_IN), .A(n8376), .B(
        n8375), .ZN(n8379) );
  NAND2_X1 U9652 ( .A1(n11028), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n8378) );
  OAI21_X1 U9653 ( .B1(n10235), .B2(n10153), .A(n6947), .ZN(n8377) );
  OAI211_X1 U9654 ( .C1(n8379), .C2(n10180), .A(n8378), .B(n8377), .ZN(
        P1_U3293) );
  INV_X1 U9655 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10568) );
  OAI222_X1 U9656 ( .A1(n10337), .A2(n10568), .B1(n10340), .B2(n8380), .C1(
        P1_U3086), .C2(n6594), .ZN(P1_U3333) );
  OAI222_X1 U9657 ( .A1(n9516), .A2(n8383), .B1(n9518), .B2(n8382), .C1(
        P2_U3151), .C2(n8381), .ZN(P2_U3268) );
  MUX2_X1 U9658 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n8684), .Z(n8388) );
  INV_X1 U9659 ( .A(n8388), .ZN(n8389) );
  MUX2_X1 U9660 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n8684), .Z(n8681) );
  XNOR2_X1 U9661 ( .A(n8681), .B(SI_30_), .ZN(n8682) );
  NAND2_X1 U9662 ( .A1(n9734), .A2(n8689), .ZN(n8394) );
  NAND2_X1 U9663 ( .A1(n8392), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8393) );
  INV_X1 U9664 ( .A(n8395), .ZN(n8396) );
  NAND2_X1 U9665 ( .A1(n8396), .A2(n10589), .ZN(n8397) );
  NAND2_X1 U9666 ( .A1(n8398), .A2(n8397), .ZN(n10336) );
  NAND2_X1 U9667 ( .A1(n8392), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U9668 ( .A1(n5107), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8404) );
  NAND2_X1 U9669 ( .A1(n8540), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U9670 ( .A1(n8597), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8402) );
  AND2_X1 U9671 ( .A1(n8737), .A2(n8679), .ZN(n8405) );
  NAND2_X1 U9672 ( .A1(n8406), .A2(n8689), .ZN(n8408) );
  NAND2_X1 U9673 ( .A1(n8392), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8407) );
  INV_X1 U9674 ( .A(n8877), .ZN(n9385) );
  NAND2_X1 U9675 ( .A1(n8540), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U9676 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n8420), .ZN(n8409) );
  NAND2_X1 U9677 ( .A1(n8410), .A2(n8409), .ZN(n9187) );
  NAND2_X1 U9678 ( .A1(n8643), .A2(n9187), .ZN(n8413) );
  NAND2_X1 U9679 ( .A1(n5107), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8412) );
  NAND2_X1 U9680 ( .A1(n8597), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8411) );
  NAND4_X1 U9681 ( .A1(n8414), .A2(n8413), .A3(n8412), .A4(n8411), .ZN(n9058)
         );
  NAND2_X1 U9682 ( .A1(n9058), .A2(n8670), .ZN(n8415) );
  NAND2_X1 U9683 ( .A1(n8416), .A2(n8689), .ZN(n8418) );
  NAND2_X1 U9684 ( .A1(n8392), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8417) );
  NAND2_X1 U9685 ( .A1(n8540), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8425) );
  INV_X1 U9686 ( .A(n8419), .ZN(n8429) );
  NAND2_X1 U9687 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(n8429), .ZN(n8421) );
  NAND2_X1 U9688 ( .A1(n8421), .A2(n8420), .ZN(n9200) );
  NAND2_X1 U9689 ( .A1(n8643), .A2(n9200), .ZN(n8424) );
  NAND2_X1 U9690 ( .A1(n5107), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U9691 ( .A1(n8597), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8422) );
  NAND4_X1 U9692 ( .A1(n8425), .A2(n8424), .A3(n8423), .A4(n8422), .ZN(n9180)
         );
  MUX2_X1 U9693 ( .A(n8724), .B(n8723), .S(n8679), .Z(n8668) );
  INV_X1 U9694 ( .A(n9198), .ZN(n9191) );
  NAND2_X1 U9695 ( .A1(n8392), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8427) );
  NAND2_X1 U9696 ( .A1(n8441), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U9697 ( .A1(n8430), .A2(n8429), .ZN(n9212) );
  NAND2_X1 U9698 ( .A1(n9212), .A2(n8643), .ZN(n8435) );
  INV_X1 U9699 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U9700 ( .A1(n8540), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8432) );
  NAND2_X1 U9701 ( .A1(n8597), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8431) );
  OAI211_X1 U9702 ( .C1(n9213), .C2(n5106), .A(n8432), .B(n8431), .ZN(n8433)
         );
  INV_X1 U9703 ( .A(n8433), .ZN(n8434) );
  NAND2_X1 U9704 ( .A1(n8435), .A2(n8434), .ZN(n9059) );
  INV_X1 U9705 ( .A(n9216), .ZN(n9205) );
  NAND2_X1 U9706 ( .A1(n8436), .A2(n8689), .ZN(n8438) );
  NAND2_X1 U9707 ( .A1(n8392), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8437) );
  OR2_X1 U9708 ( .A1(n8639), .A2(n8439), .ZN(n8440) );
  NAND2_X1 U9709 ( .A1(n8441), .A2(n8440), .ZN(n9227) );
  NAND2_X1 U9710 ( .A1(n9227), .A2(n8643), .ZN(n8447) );
  INV_X1 U9711 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8444) );
  NAND2_X1 U9712 ( .A1(n8540), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U9713 ( .A1(n8597), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8442) );
  OAI211_X1 U9714 ( .C1(n5106), .C2(n8444), .A(n8443), .B(n8442), .ZN(n8445)
         );
  INV_X1 U9715 ( .A(n8445), .ZN(n8446) );
  NAND2_X1 U9716 ( .A1(n8447), .A2(n8446), .ZN(n9207) );
  NAND2_X1 U9717 ( .A1(n9220), .A2(n9237), .ZN(n8721) );
  MUX2_X1 U9718 ( .A(n8721), .B(n8655), .S(n8679), .Z(n8663) );
  AND2_X1 U9719 ( .A1(n8472), .A2(n8499), .ZN(n8476) );
  INV_X1 U9720 ( .A(n8448), .ZN(n8450) );
  OAI211_X1 U9721 ( .C1(n8452), .C2(n8451), .A(n8450), .B(n8449), .ZN(n8453)
         );
  OAI21_X1 U9722 ( .B1(n8455), .B2(n8454), .A(n8453), .ZN(n8460) );
  INV_X1 U9723 ( .A(n8456), .ZN(n8458) );
  NAND2_X1 U9724 ( .A1(n8744), .A2(n8741), .ZN(n8457) );
  NAND2_X1 U9725 ( .A1(n8458), .A2(n8457), .ZN(n8459) );
  MUX2_X1 U9726 ( .A(n8460), .B(n8459), .S(n8679), .Z(n8469) );
  NAND2_X1 U9727 ( .A1(n8462), .A2(n8461), .ZN(n8465) );
  NAND2_X1 U9728 ( .A1(n8471), .A2(n8463), .ZN(n8464) );
  MUX2_X1 U9729 ( .A(n8465), .B(n8464), .S(n8679), .Z(n8466) );
  INV_X1 U9730 ( .A(n8466), .ZN(n8467) );
  OAI21_X1 U9731 ( .B1(n8469), .B2(n8468), .A(n8467), .ZN(n8470) );
  NAND2_X1 U9732 ( .A1(n8470), .A2(n8747), .ZN(n8480) );
  INV_X1 U9733 ( .A(n8471), .ZN(n8474) );
  OAI211_X1 U9734 ( .C1(n8480), .C2(n8474), .A(n8473), .B(n8472), .ZN(n8475)
         );
  MUX2_X1 U9735 ( .A(n8476), .B(n8475), .S(n8670), .Z(n8482) );
  AND3_X1 U9736 ( .A1(n8485), .A2(n8477), .A3(n8679), .ZN(n8478) );
  OAI21_X1 U9737 ( .B1(n8480), .B2(n8479), .A(n8478), .ZN(n8481) );
  NAND2_X1 U9738 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  NAND2_X1 U9739 ( .A1(n8483), .A2(n8484), .ZN(n8488) );
  NAND2_X1 U9740 ( .A1(n8485), .A2(n8484), .ZN(n8486) );
  NAND2_X1 U9741 ( .A1(n8486), .A2(n8670), .ZN(n8487) );
  NAND2_X1 U9742 ( .A1(n8488), .A2(n8487), .ZN(n8493) );
  AND2_X1 U9743 ( .A1(n8496), .A2(n8495), .ZN(n8489) );
  MUX2_X1 U9744 ( .A(n8490), .B(n8489), .S(n8670), .Z(n8491) );
  NAND2_X1 U9745 ( .A1(n8491), .A2(n8506), .ZN(n8508) );
  NOR2_X1 U9746 ( .A1(n8508), .A2(n8750), .ZN(n8492) );
  NAND2_X1 U9747 ( .A1(n8493), .A2(n8492), .ZN(n8502) );
  AND2_X1 U9748 ( .A1(n8495), .A2(n8494), .ZN(n8497) );
  OAI211_X1 U9749 ( .C1(n8508), .C2(n8497), .A(n8509), .B(n8496), .ZN(n8498)
         );
  NAND2_X1 U9750 ( .A1(n8498), .A2(n8679), .ZN(n8501) );
  NOR2_X1 U9751 ( .A1(n8499), .A2(n8679), .ZN(n8500) );
  AOI21_X1 U9752 ( .B1(n8502), .B2(n8501), .A(n8500), .ZN(n8511) );
  INV_X1 U9753 ( .A(n8511), .ZN(n8504) );
  NAND2_X1 U9754 ( .A1(n8514), .A2(n8505), .ZN(n8503) );
  OAI21_X1 U9755 ( .B1(n8504), .B2(n8503), .A(n8512), .ZN(n8517) );
  OAI211_X1 U9756 ( .C1(n8508), .C2(n8507), .A(n8506), .B(n8505), .ZN(n8510)
         );
  OAI21_X1 U9757 ( .B1(n8511), .B2(n8510), .A(n8509), .ZN(n8515) );
  INV_X1 U9758 ( .A(n8512), .ZN(n8513) );
  AOI21_X1 U9759 ( .B1(n8515), .B2(n8514), .A(n8513), .ZN(n8516) );
  MUX2_X1 U9760 ( .A(n8517), .B(n8516), .S(n8670), .Z(n8519) );
  NAND2_X1 U9761 ( .A1(n8519), .A2(n8518), .ZN(n8524) );
  NOR2_X1 U9762 ( .A1(n11107), .A2(n8679), .ZN(n8521) );
  AND2_X1 U9763 ( .A1(n11107), .A2(n8679), .ZN(n8520) );
  MUX2_X1 U9764 ( .A(n8521), .B(n8520), .S(n9007), .Z(n8522) );
  NOR2_X1 U9765 ( .A1(n8759), .A2(n8522), .ZN(n8523) );
  NAND2_X1 U9766 ( .A1(n8524), .A2(n8523), .ZN(n8529) );
  INV_X1 U9767 ( .A(n8525), .ZN(n8526) );
  MUX2_X1 U9768 ( .A(n8527), .B(n8526), .S(n8670), .Z(n8528) );
  NAND3_X1 U9769 ( .A1(n8529), .A2(n8760), .A3(n8528), .ZN(n8532) );
  INV_X1 U9770 ( .A(n9362), .ZN(n8804) );
  NAND2_X1 U9771 ( .A1(n8916), .A2(n8804), .ZN(n8530) );
  OR2_X1 U9772 ( .A1(n8916), .A2(n8804), .ZN(n8700) );
  MUX2_X1 U9773 ( .A(n8530), .B(n8700), .S(n8670), .Z(n8531) );
  NAND2_X1 U9774 ( .A1(n8532), .A2(n8531), .ZN(n8549) );
  NAND2_X1 U9775 ( .A1(n8533), .A2(n8689), .ZN(n8536) );
  AOI22_X1 U9776 ( .A1(n8392), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8578), .B2(
        n8534), .ZN(n8535) );
  INV_X1 U9777 ( .A(n9060), .ZN(n8813) );
  OR2_X1 U9778 ( .A1(n9370), .A2(n8813), .ZN(n9342) );
  NAND2_X1 U9779 ( .A1(n9370), .A2(n8813), .ZN(n8702) );
  NAND2_X1 U9780 ( .A1(n9342), .A2(n8702), .ZN(n9371) );
  INV_X1 U9781 ( .A(n9371), .ZN(n8762) );
  NAND2_X1 U9782 ( .A1(n8537), .A2(n8689), .ZN(n8539) );
  AOI22_X1 U9783 ( .A1(n8392), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8578), .B2(
        n9145), .ZN(n8538) );
  NAND2_X1 U9784 ( .A1(n8540), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8547) );
  INV_X1 U9785 ( .A(n8541), .ZN(n8556) );
  NAND2_X1 U9786 ( .A1(n8542), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U9787 ( .A1(n8556), .A2(n8543), .ZN(n9351) );
  NAND2_X1 U9788 ( .A1(n8643), .A2(n9351), .ZN(n8546) );
  NAND2_X1 U9789 ( .A1(n8187), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U9790 ( .A1(n8597), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8544) );
  NAND4_X1 U9791 ( .A1(n8547), .A2(n8546), .A3(n8545), .A4(n8544), .ZN(n9361)
         );
  INV_X1 U9792 ( .A(n9361), .ZN(n9051) );
  NAND2_X1 U9793 ( .A1(n8964), .A2(n9051), .ZN(n8739) );
  OAI21_X1 U9794 ( .B1(n8702), .B2(n8670), .A(n8739), .ZN(n8548) );
  AOI21_X1 U9795 ( .B1(n8549), .B2(n8762), .A(n8548), .ZN(n8551) );
  INV_X1 U9796 ( .A(n8740), .ZN(n8550) );
  AND2_X1 U9797 ( .A1(n8740), .A2(n9342), .ZN(n8703) );
  OAI22_X1 U9798 ( .A1(n8551), .A2(n8550), .B1(n8679), .B2(n8703), .ZN(n8563)
         );
  NAND2_X1 U9799 ( .A1(n8552), .A2(n8689), .ZN(n8554) );
  AOI22_X1 U9800 ( .A1(n8392), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8578), .B2(
        n9165), .ZN(n8553) );
  NAND2_X1 U9801 ( .A1(n8540), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8561) );
  INV_X1 U9802 ( .A(n8555), .ZN(n8568) );
  NAND2_X1 U9803 ( .A1(n8556), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U9804 ( .A1(n8568), .A2(n8557), .ZN(n9337) );
  NAND2_X1 U9805 ( .A1(n8643), .A2(n9337), .ZN(n8560) );
  NAND2_X1 U9806 ( .A1(n8187), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U9807 ( .A1(n7194), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8558) );
  NAND4_X1 U9808 ( .A1(n8561), .A2(n8560), .A3(n8559), .A4(n8558), .ZN(n9316)
         );
  INV_X1 U9809 ( .A(n9316), .ZN(n8562) );
  OR2_X1 U9810 ( .A1(n9336), .A2(n8562), .ZN(n8589) );
  NAND2_X1 U9811 ( .A1(n9336), .A2(n8562), .ZN(n8705) );
  NAND2_X1 U9812 ( .A1(n8589), .A2(n8705), .ZN(n8859) );
  NAND2_X1 U9813 ( .A1(n8563), .A2(n9334), .ZN(n8576) );
  NAND2_X1 U9814 ( .A1(n8564), .A2(n8689), .ZN(n8567) );
  AOI22_X1 U9815 ( .A1(n8392), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8578), .B2(
        n8565), .ZN(n8566) );
  NAND2_X1 U9816 ( .A1(n8540), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U9817 ( .A1(n8568), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U9818 ( .A1(n8582), .A2(n8569), .ZN(n9320) );
  NAND2_X1 U9819 ( .A1(n8643), .A2(n9320), .ZN(n8572) );
  NAND2_X1 U9820 ( .A1(n7226), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U9821 ( .A1(n7194), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8570) );
  NAND4_X1 U9822 ( .A1(n8573), .A2(n8572), .A3(n8571), .A4(n8570), .ZN(n9303)
         );
  INV_X1 U9823 ( .A(n9303), .ZN(n8940) );
  NAND2_X1 U9824 ( .A1(n9428), .A2(n8940), .ZN(n8574) );
  INV_X1 U9825 ( .A(n9324), .ZN(n8765) );
  MUX2_X1 U9826 ( .A(n8589), .B(n8705), .S(n8679), .Z(n8575) );
  NAND3_X1 U9827 ( .A1(n8576), .A2(n8765), .A3(n8575), .ZN(n8593) );
  NAND2_X1 U9828 ( .A1(n8577), .A2(n8689), .ZN(n8581) );
  AOI22_X1 U9829 ( .A1(n8392), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8579), .B2(
        n8578), .ZN(n8580) );
  NAND2_X1 U9830 ( .A1(n8582), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U9831 ( .A1(n8599), .A2(n8583), .ZN(n9309) );
  NAND2_X1 U9832 ( .A1(n9309), .A2(n8643), .ZN(n8587) );
  NAND2_X1 U9833 ( .A1(n5107), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U9834 ( .A1(n8540), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U9835 ( .A1(n8597), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U9836 ( .A1(n8934), .A2(n9290), .ZN(n9292) );
  INV_X1 U9837 ( .A(n8739), .ZN(n8588) );
  AND2_X1 U9838 ( .A1(n8589), .A2(n8588), .ZN(n8591) );
  XNOR2_X1 U9839 ( .A(n8707), .B(n8670), .ZN(n8590) );
  OAI21_X1 U9840 ( .B1(n9324), .B2(n8591), .A(n8590), .ZN(n8592) );
  NAND3_X1 U9841 ( .A1(n8593), .A2(n5533), .A3(n8592), .ZN(n8605) );
  NAND2_X1 U9842 ( .A1(n8594), .A2(n8689), .ZN(n8596) );
  NAND2_X1 U9843 ( .A1(n8392), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8595) );
  INV_X1 U9844 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9484) );
  INV_X1 U9845 ( .A(n8598), .ZN(n8609) );
  NAND2_X1 U9846 ( .A1(n8599), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U9847 ( .A1(n8609), .A2(n8600), .ZN(n9296) );
  NAND2_X1 U9848 ( .A1(n9296), .A2(n8643), .ZN(n8602) );
  AOI22_X1 U9849 ( .A1(n8540), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5107), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n8601) );
  OAI211_X1 U9850 ( .C1(n7248), .C2(n9484), .A(n8602), .B(n8601), .ZN(n9304)
         );
  INV_X1 U9851 ( .A(n9304), .ZN(n8826) );
  NAND2_X1 U9852 ( .A1(n9273), .A2(n8708), .ZN(n8603) );
  NAND2_X1 U9853 ( .A1(n8603), .A2(n8670), .ZN(n8604) );
  NAND2_X1 U9854 ( .A1(n8605), .A2(n8604), .ZN(n8607) );
  NAND2_X1 U9855 ( .A1(n9295), .A2(n8826), .ZN(n8738) );
  AND2_X1 U9856 ( .A1(n8738), .A2(n9292), .ZN(n9272) );
  NOR2_X1 U9857 ( .A1(n9272), .A2(n8670), .ZN(n8606) );
  AOI21_X1 U9858 ( .B1(n8607), .B2(n8738), .A(n8606), .ZN(n8632) );
  INV_X1 U9859 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8613) );
  INV_X1 U9860 ( .A(n8608), .ZN(n8621) );
  NAND2_X1 U9861 ( .A1(n8609), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U9862 ( .A1(n8621), .A2(n8610), .ZN(n8946) );
  NAND2_X1 U9863 ( .A1(n8946), .A2(n8643), .ZN(n8612) );
  AOI22_X1 U9864 ( .A1(n8540), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5107), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n8611) );
  OAI211_X1 U9865 ( .C1(n7248), .C2(n8613), .A(n8612), .B(n8611), .ZN(n9261)
         );
  NAND2_X1 U9866 ( .A1(n8614), .A2(n8689), .ZN(n8616) );
  NAND2_X1 U9867 ( .A1(n8392), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8615) );
  MUX2_X1 U9868 ( .A(n9261), .B(n8628), .S(n8679), .Z(n8629) );
  INV_X1 U9869 ( .A(n8865), .ZN(n8617) );
  OAI22_X1 U9870 ( .A1(n8629), .A2(n8617), .B1(n8670), .B2(n9273), .ZN(n8631)
         );
  NAND2_X1 U9871 ( .A1(n8618), .A2(n8689), .ZN(n8620) );
  NAND2_X1 U9872 ( .A1(n8392), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U9873 ( .A1(n8621), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U9874 ( .A1(n8623), .A2(n8622), .ZN(n9266) );
  INV_X1 U9875 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U9876 ( .A1(n8540), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U9877 ( .A1(n8597), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8624) );
  OAI211_X1 U9878 ( .C1(n5106), .C2(n8626), .A(n8625), .B(n8624), .ZN(n8627)
         );
  AOI21_X1 U9879 ( .B1(n9266), .B2(n8643), .A(n8627), .ZN(n8947) );
  NOR2_X1 U9880 ( .A1(n9411), .A2(n8947), .ZN(n8712) );
  NAND2_X1 U9881 ( .A1(n9411), .A2(n8947), .ZN(n8715) );
  INV_X1 U9882 ( .A(n8715), .ZN(n8651) );
  OR2_X1 U9883 ( .A1(n8712), .A2(n8651), .ZN(n9264) );
  INV_X1 U9884 ( .A(n9264), .ZN(n8767) );
  NAND2_X1 U9885 ( .A1(n8628), .A2(n9261), .ZN(n8864) );
  NAND2_X1 U9886 ( .A1(n8629), .A2(n8864), .ZN(n8630) );
  OAI211_X1 U9887 ( .C1(n8632), .C2(n8631), .A(n8767), .B(n8630), .ZN(n8654)
         );
  NAND2_X1 U9888 ( .A1(n8633), .A2(n8689), .ZN(n8635) );
  NAND2_X1 U9889 ( .A1(n8392), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U9890 ( .A1(n9253), .A2(n9238), .ZN(n8656) );
  NAND2_X1 U9891 ( .A1(n8636), .A2(n8689), .ZN(n8638) );
  NAND2_X1 U9892 ( .A1(n8392), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8637) );
  INV_X1 U9893 ( .A(n8639), .ZN(n8642) );
  NAND2_X1 U9894 ( .A1(n8640), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U9895 ( .A1(n8642), .A2(n8641), .ZN(n9240) );
  NAND2_X1 U9896 ( .A1(n9240), .A2(n8643), .ZN(n8649) );
  INV_X1 U9897 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U9898 ( .A1(n8540), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U9899 ( .A1(n8597), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8644) );
  OAI211_X1 U9900 ( .C1(n8646), .C2(n5106), .A(n8645), .B(n8644), .ZN(n8647)
         );
  INV_X1 U9901 ( .A(n8647), .ZN(n8648) );
  NAND2_X1 U9902 ( .A1(n8649), .A2(n8648), .ZN(n9248) );
  INV_X1 U9903 ( .A(n8872), .ZN(n8650) );
  MUX2_X1 U9904 ( .A(n8651), .B(n8712), .S(n8679), .Z(n8652) );
  INV_X1 U9905 ( .A(n8652), .ZN(n8653) );
  NAND4_X1 U9906 ( .A1(n8654), .A2(n9251), .A3(n9242), .A4(n8653), .ZN(n8661)
         );
  MUX2_X1 U9907 ( .A(n8717), .B(n8656), .S(n8679), .Z(n8657) );
  NAND2_X1 U9908 ( .A1(n9242), .A2(n8657), .ZN(n8659) );
  INV_X1 U9909 ( .A(n9248), .ZN(n9225) );
  NAND2_X1 U9910 ( .A1(n9232), .A2(n9225), .ZN(n8718) );
  OR2_X1 U9911 ( .A1(n9232), .A2(n9225), .ZN(n8719) );
  MUX2_X1 U9912 ( .A(n8718), .B(n8719), .S(n8679), .Z(n8658) );
  NAND2_X1 U9913 ( .A1(n8659), .A2(n8658), .ZN(n8660) );
  NAND3_X1 U9914 ( .A1(n8661), .A2(n9221), .A3(n8660), .ZN(n8662) );
  NAND3_X1 U9915 ( .A1(n9205), .A2(n8663), .A3(n8662), .ZN(n8666) );
  NAND2_X1 U9916 ( .A1(n9392), .A2(n9224), .ZN(n8664) );
  MUX2_X1 U9917 ( .A(n8722), .B(n8664), .S(n8679), .Z(n8665) );
  NAND3_X1 U9918 ( .A1(n9191), .A2(n8666), .A3(n8665), .ZN(n8667) );
  AND2_X1 U9919 ( .A1(n8668), .A2(n8667), .ZN(n8673) );
  NAND2_X1 U9920 ( .A1(n9058), .A2(n8679), .ZN(n9194) );
  INV_X1 U9921 ( .A(n9194), .ZN(n8669) );
  AOI21_X1 U9922 ( .B1(n8877), .B2(n8670), .A(n8669), .ZN(n8671) );
  OAI21_X1 U9923 ( .B1(n8674), .B2(n8673), .A(n8671), .ZN(n8676) );
  INV_X1 U9924 ( .A(n8737), .ZN(n8672) );
  NAND2_X1 U9925 ( .A1(n8676), .A2(n8675), .ZN(n8680) );
  INV_X1 U9926 ( .A(n8680), .ZN(n8678) );
  AOI21_X1 U9927 ( .B1(n8678), .B2(n8736), .A(n8677), .ZN(n8699) );
  INV_X1 U9928 ( .A(n8732), .ZN(n8772) );
  AOI211_X1 U9929 ( .C1(n8680), .C2(n8736), .A(n8679), .B(n8772), .ZN(n8698)
         );
  MUX2_X1 U9930 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8684), .Z(n8686) );
  INV_X1 U9931 ( .A(SI_31_), .ZN(n8685) );
  XNOR2_X1 U9932 ( .A(n8686), .B(n8685), .ZN(n8687) );
  NAND2_X1 U9933 ( .A1(n9645), .A2(n8689), .ZN(n8691) );
  NAND2_X1 U9934 ( .A1(n8392), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U9935 ( .A1(n8540), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U9936 ( .A1(n5107), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U9937 ( .A1(n8597), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8692) );
  NAND4_X1 U9938 ( .A1(n8695), .A2(n8694), .A3(n8693), .A4(n8692), .ZN(n9172)
         );
  INV_X1 U9939 ( .A(n9172), .ZN(n8696) );
  OR2_X1 U9940 ( .A1(n8728), .A2(n8696), .ZN(n8697) );
  NAND2_X1 U9941 ( .A1(n9175), .A2(n8886), .ZN(n8730) );
  NAND2_X1 U9942 ( .A1(n8697), .A2(n8730), .ZN(n8773) );
  NAND2_X1 U9943 ( .A1(n8701), .A2(n8700), .ZN(n9372) );
  NAND2_X1 U9944 ( .A1(n9372), .A2(n8702), .ZN(n9343) );
  NAND2_X1 U9945 ( .A1(n9343), .A2(n8703), .ZN(n8704) );
  NAND2_X1 U9946 ( .A1(n8704), .A2(n8739), .ZN(n9335) );
  NAND2_X1 U9947 ( .A1(n9335), .A2(n9334), .ZN(n8706) );
  NAND2_X1 U9948 ( .A1(n8706), .A2(n8705), .ZN(n9325) );
  NAND2_X1 U9949 ( .A1(n8865), .A2(n8864), .ZN(n9277) );
  AND2_X1 U9950 ( .A1(n9272), .A2(n9277), .ZN(n8711) );
  INV_X1 U9951 ( .A(n9273), .ZN(n8709) );
  AND2_X1 U9952 ( .A1(n9277), .A2(n8709), .ZN(n8710) );
  INV_X1 U9953 ( .A(n9261), .ZN(n9288) );
  OR2_X1 U9954 ( .A1(n8628), .A2(n9288), .ZN(n9263) );
  INV_X1 U9955 ( .A(n8712), .ZN(n8713) );
  AND2_X1 U9956 ( .A1(n9263), .A2(n8713), .ZN(n8714) );
  NAND2_X1 U9957 ( .A1(n9275), .A2(n8714), .ZN(n8716) );
  NAND2_X1 U9958 ( .A1(n8716), .A2(n8715), .ZN(n9252) );
  OAI21_X2 U9959 ( .B1(n9252), .B2(n9246), .A(n8717), .ZN(n9241) );
  NAND2_X1 U9960 ( .A1(n9241), .A2(n8718), .ZN(n8720) );
  INV_X1 U9961 ( .A(n8723), .ZN(n8725) );
  NAND2_X1 U9962 ( .A1(n9184), .A2(n9183), .ZN(n9186) );
  INV_X1 U9963 ( .A(n9058), .ZN(n8876) );
  NAND2_X1 U9964 ( .A1(n8877), .A2(n8876), .ZN(n8726) );
  NAND2_X1 U9965 ( .A1(n9186), .A2(n8726), .ZN(n8882) );
  NAND2_X1 U9966 ( .A1(n8882), .A2(n8737), .ZN(n8731) );
  NOR2_X1 U9967 ( .A1(n9175), .A2(n9172), .ZN(n8727) );
  OR2_X1 U9968 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  NAND4_X1 U9969 ( .A1(n8731), .A2(n8736), .A3(n8730), .A4(n8729), .ZN(n8734)
         );
  NAND2_X1 U9970 ( .A1(n8728), .A2(n8772), .ZN(n8733) );
  NAND2_X1 U9971 ( .A1(n8735), .A2(n8774), .ZN(n8777) );
  NAND2_X1 U9972 ( .A1(n8740), .A2(n8739), .ZN(n9348) );
  INV_X1 U9973 ( .A(n9348), .ZN(n8857) );
  AND4_X1 U9974 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(n8748)
         );
  NAND4_X1 U9975 ( .A1(n8748), .A2(n8747), .A3(n8746), .A4(n8745), .ZN(n8752)
         );
  NOR4_X1 U9976 ( .A1(n8752), .A2(n8751), .A3(n8750), .A4(n8749), .ZN(n8756)
         );
  INV_X1 U9977 ( .A(n8753), .ZN(n8754) );
  NAND3_X1 U9978 ( .A1(n8756), .A2(n8755), .A3(n8754), .ZN(n8757) );
  NOR3_X1 U9979 ( .A1(n8759), .A2(n8758), .A3(n8757), .ZN(n8761) );
  NAND4_X1 U9980 ( .A1(n8857), .A2(n8762), .A3(n8761), .A4(n8760), .ZN(n8763)
         );
  NOR2_X1 U9981 ( .A1(n8859), .A2(n8763), .ZN(n8764) );
  AND4_X1 U9982 ( .A1(n9293), .A2(n5533), .A3(n8765), .A4(n8764), .ZN(n8766)
         );
  AND4_X1 U9983 ( .A1(n9251), .A2(n8767), .A3(n8766), .A4(n9277), .ZN(n8768)
         );
  NAND3_X1 U9984 ( .A1(n9221), .A2(n8768), .A3(n9242), .ZN(n8769) );
  NOR3_X1 U9985 ( .A1(n9198), .A2(n9216), .A3(n8769), .ZN(n8770) );
  NAND2_X1 U9986 ( .A1(n9183), .A2(n8770), .ZN(n8771) );
  NAND3_X1 U9987 ( .A1(n8781), .A2(n8780), .A3(n8779), .ZN(n8782) );
  NOR3_X1 U9988 ( .A1(n8787), .A2(n8786), .A3(n8785), .ZN(n8795) );
  NOR4_X1 U9989 ( .A1(n8790), .A2(n9508), .A3(n8789), .A4(n8788), .ZN(n8794)
         );
  OAI21_X1 U9990 ( .B1(n8792), .B2(n8791), .A(P2_B_REG_SCAN_IN), .ZN(n8793) );
  OAI22_X1 U9991 ( .A1(n8796), .A2(n8795), .B1(n8794), .B2(n8793), .ZN(
        P2_U3296) );
  OAI222_X1 U9992 ( .A1(n9516), .A2(n8799), .B1(n9518), .B2(n8798), .C1(n8797), 
        .C2(P2_U3151), .ZN(P2_U3271) );
  XNOR2_X1 U9993 ( .A(n9336), .B(n5099), .ZN(n8818) );
  XNOR2_X1 U9994 ( .A(n11122), .B(n5099), .ZN(n8808) );
  NAND2_X1 U9995 ( .A1(n8808), .A2(n8803), .ZN(n9001) );
  XNOR2_X1 U9996 ( .A(n8916), .B(n5099), .ZN(n8807) );
  NAND2_X1 U9997 ( .A1(n8807), .A2(n8804), .ZN(n8806) );
  AND2_X1 U9998 ( .A1(n9001), .A2(n8806), .ZN(n9041) );
  XNOR2_X1 U9999 ( .A(n9370), .B(n5099), .ZN(n8814) );
  XOR2_X1 U10000 ( .A(n9060), .B(n8814), .Z(n9044) );
  INV_X1 U10001 ( .A(n9044), .ZN(n8805) );
  INV_X1 U10002 ( .A(n8806), .ZN(n8812) );
  XOR2_X1 U10003 ( .A(n9362), .B(n8807), .Z(n8911) );
  INV_X1 U10004 ( .A(n8911), .ZN(n8810) );
  INV_X1 U10005 ( .A(n8808), .ZN(n8809) );
  NAND2_X1 U10006 ( .A1(n8809), .A2(n9061), .ZN(n9002) );
  AND2_X1 U10007 ( .A1(n8810), .A2(n9002), .ZN(n8811) );
  XNOR2_X1 U10008 ( .A(n8964), .B(n5099), .ZN(n8815) );
  XNOR2_X1 U10009 ( .A(n8815), .B(n9361), .ZN(n8966) );
  NAND2_X1 U10010 ( .A1(n8967), .A2(n8966), .ZN(n8965) );
  INV_X1 U10011 ( .A(n8815), .ZN(n8816) );
  NAND2_X1 U10012 ( .A1(n8816), .A2(n9361), .ZN(n8817) );
  NAND2_X1 U10013 ( .A1(n8965), .A2(n8817), .ZN(n8975) );
  INV_X1 U10014 ( .A(n8975), .ZN(n8820) );
  XOR2_X1 U10015 ( .A(n9316), .B(n8818), .Z(n8976) );
  INV_X1 U10016 ( .A(n8976), .ZN(n8819) );
  XNOR2_X1 U10017 ( .A(n9428), .B(n5099), .ZN(n8821) );
  XOR2_X1 U10018 ( .A(n9303), .B(n8821), .Z(n9020) );
  INV_X1 U10019 ( .A(n8821), .ZN(n8822) );
  NAND2_X1 U10020 ( .A1(n8822), .A2(n9303), .ZN(n8823) );
  INV_X1 U10021 ( .A(n8936), .ZN(n8824) );
  INV_X1 U10022 ( .A(n9290), .ZN(n9317) );
  NAND2_X1 U10023 ( .A1(n8824), .A2(n9317), .ZN(n8825) );
  XNOR2_X1 U10024 ( .A(n9295), .B(n5099), .ZN(n8827) );
  XOR2_X1 U10025 ( .A(n9304), .B(n8827), .Z(n8995) );
  NAND2_X1 U10026 ( .A1(n8827), .A2(n8826), .ZN(n8828) );
  XNOR2_X1 U10027 ( .A(n8829), .B(n9261), .ZN(n8945) );
  XNOR2_X1 U10028 ( .A(n9411), .B(n5099), .ZN(n8830) );
  XOR2_X1 U10029 ( .A(n8947), .B(n8830), .Z(n9013) );
  INV_X1 U10030 ( .A(n8830), .ZN(n8831) );
  INV_X1 U10031 ( .A(n8947), .ZN(n9247) );
  NAND2_X1 U10032 ( .A1(n8831), .A2(n9247), .ZN(n8832) );
  NAND2_X1 U10033 ( .A1(n9012), .A2(n8832), .ZN(n8833) );
  XNOR2_X1 U10034 ( .A(n9253), .B(n5099), .ZN(n8834) );
  NAND2_X1 U10035 ( .A1(n8919), .A2(n9238), .ZN(n8984) );
  INV_X1 U10036 ( .A(n8833), .ZN(n8835) );
  NAND2_X1 U10037 ( .A1(n8835), .A2(n8834), .ZN(n8983) );
  XNOR2_X1 U10038 ( .A(n9232), .B(n5099), .ZN(n8838) );
  NAND2_X1 U10039 ( .A1(n8838), .A2(n9225), .ZN(n8837) );
  NAND2_X2 U10040 ( .A1(n8984), .A2(n8836), .ZN(n8956) );
  INV_X1 U10041 ( .A(n8837), .ZN(n8839) );
  XNOR2_X1 U10042 ( .A(n8838), .B(n9248), .ZN(n8986) );
  XNOR2_X1 U10043 ( .A(n9220), .B(n5099), .ZN(n8841) );
  XNOR2_X1 U10044 ( .A(n8841), .B(n9207), .ZN(n8958) );
  NAND2_X1 U10045 ( .A1(n8841), .A2(n9237), .ZN(n9030) );
  XNOR2_X1 U10046 ( .A(n9392), .B(n5099), .ZN(n8846) );
  NAND2_X1 U10047 ( .A1(n8846), .A2(n9224), .ZN(n8845) );
  AND2_X1 U10048 ( .A1(n9030), .A2(n8845), .ZN(n8899) );
  XNOR2_X1 U10049 ( .A(n8896), .B(n8842), .ZN(n8843) );
  NAND2_X1 U10050 ( .A1(n8843), .A2(n9180), .ZN(n8848) );
  OAI21_X1 U10051 ( .B1(n8843), .B2(n9180), .A(n8848), .ZN(n8900) );
  INV_X1 U10052 ( .A(n8900), .ZN(n8844) );
  INV_X1 U10053 ( .A(n8845), .ZN(n8847) );
  XNOR2_X1 U10054 ( .A(n8846), .B(n9059), .ZN(n9033) );
  XNOR2_X1 U10055 ( .A(n9183), .B(n5099), .ZN(n8849) );
  NAND2_X1 U10056 ( .A1(n9053), .A2(n9187), .ZN(n8851) );
  AOI22_X1 U10057 ( .A1(n9048), .A2(n9180), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8850) );
  OAI211_X1 U10058 ( .C1(n9057), .C2(n9050), .A(n8851), .B(n8850), .ZN(n8852)
         );
  AOI21_X1 U10059 ( .B1(n8877), .B2(n11077), .A(n8852), .ZN(n8853) );
  OAI21_X1 U10060 ( .B1(n8854), .B2(n11072), .A(n8853), .ZN(P2_U3160) );
  NAND2_X1 U10061 ( .A1(n8916), .A2(n9362), .ZN(n8855) );
  AND2_X1 U10062 ( .A1(n9371), .A2(n9348), .ZN(n8858) );
  NAND2_X1 U10063 ( .A1(n9370), .A2(n9060), .ZN(n9345) );
  NAND2_X1 U10064 ( .A1(n8964), .A2(n9361), .ZN(n9329) );
  NAND2_X1 U10065 ( .A1(n9346), .A2(n9329), .ZN(n8860) );
  NAND2_X1 U10066 ( .A1(n8860), .A2(n8859), .ZN(n9331) );
  NAND2_X1 U10067 ( .A1(n9336), .A2(n9316), .ZN(n8861) );
  NAND2_X1 U10068 ( .A1(n9331), .A2(n8861), .ZN(n9315) );
  NAND2_X1 U10069 ( .A1(n9315), .A2(n9324), .ZN(n9314) );
  NAND2_X1 U10070 ( .A1(n9428), .A2(n9303), .ZN(n8862) );
  NAND2_X1 U10071 ( .A1(n9314), .A2(n8862), .ZN(n9302) );
  NAND2_X1 U10072 ( .A1(n8934), .A2(n9317), .ZN(n8863) );
  NAND2_X1 U10073 ( .A1(n9278), .A2(n8864), .ZN(n8866) );
  NAND2_X1 U10074 ( .A1(n8866), .A2(n8865), .ZN(n9259) );
  NAND2_X1 U10075 ( .A1(n9411), .A2(n9247), .ZN(n8867) );
  NAND2_X1 U10076 ( .A1(n9259), .A2(n8867), .ZN(n8869) );
  OR2_X1 U10077 ( .A1(n9411), .A2(n9247), .ZN(n8868) );
  NAND2_X1 U10078 ( .A1(n9253), .A2(n9260), .ZN(n9234) );
  INV_X1 U10079 ( .A(n8870), .ZN(n8871) );
  NAND2_X1 U10080 ( .A1(n9220), .A2(n9207), .ZN(n8873) );
  NAND2_X1 U10081 ( .A1(n8874), .A2(n8873), .ZN(n9206) );
  NAND2_X1 U10082 ( .A1(n9385), .A2(n8876), .ZN(n8878) );
  XNOR2_X1 U10083 ( .A(n8879), .B(n8881), .ZN(n8880) );
  NAND2_X1 U10084 ( .A1(n8880), .A2(n9358), .ZN(n8889) );
  INV_X1 U10085 ( .A(n9193), .ZN(n8887) );
  NAND2_X1 U10086 ( .A1(n8884), .A2(P2_B_REG_SCAN_IN), .ZN(n8885) );
  NAND2_X1 U10087 ( .A1(n7120), .A2(n8885), .ZN(n9170) );
  OAI22_X1 U10088 ( .A1(n8887), .A2(n9194), .B1(n8886), .B2(n9170), .ZN(n8888)
         );
  INV_X1 U10089 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U10090 ( .A1(n11086), .A2(n8890), .ZN(n9169) );
  OAI21_X1 U10091 ( .B1(n11111), .B2(n8891), .A(n9169), .ZN(n8894) );
  NOR2_X1 U10092 ( .A1(n9379), .A2(n8892), .ZN(n8893) );
  OAI21_X1 U10093 ( .B1(n9382), .B2(n9352), .A(n8895), .ZN(P2_U3204) );
  INV_X1 U10094 ( .A(n8896), .ZN(n9464) );
  INV_X1 U10095 ( .A(n8897), .ZN(n8898) );
  AOI21_X1 U10096 ( .B1(n8901), .B2(n8900), .A(n11072), .ZN(n8903) );
  NAND2_X1 U10097 ( .A1(n8903), .A2(n8902), .ZN(n8907) );
  AOI22_X1 U10098 ( .A1(n9034), .A2(n9058), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8904) );
  OAI21_X1 U10099 ( .B1(n9224), .B2(n9037), .A(n8904), .ZN(n8905) );
  AOI21_X1 U10100 ( .B1(n9200), .B2(n9053), .A(n8905), .ZN(n8906) );
  OAI211_X1 U10101 ( .C1(n9464), .C2(n9056), .A(n8907), .B(n8906), .ZN(
        P2_U3154) );
  NAND2_X1 U10102 ( .A1(n8908), .A2(n9001), .ZN(n8909) );
  NAND2_X1 U10103 ( .A1(n8909), .A2(n9002), .ZN(n8910) );
  XOR2_X1 U10104 ( .A(n8911), .B(n8910), .Z(n8918) );
  NAND2_X1 U10105 ( .A1(n8912), .A2(n8950), .ZN(n8913) );
  NAND2_X1 U10106 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9100) );
  OAI211_X1 U10107 ( .C1(n8914), .C2(n11079), .A(n8913), .B(n9100), .ZN(n8915)
         );
  AOI21_X1 U10108 ( .B1(n8916), .B2(n11077), .A(n8915), .ZN(n8917) );
  OAI21_X1 U10109 ( .B1(n8918), .B2(n11072), .A(n8917), .ZN(P2_U3155) );
  XNOR2_X1 U10110 ( .A(n8919), .B(n9260), .ZN(n8924) );
  AOI22_X1 U10111 ( .A1(n9248), .A2(n9034), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8921) );
  NAND2_X1 U10112 ( .A1(n9053), .A2(n9254), .ZN(n8920) );
  OAI211_X1 U10113 ( .C1(n8947), .C2(n9037), .A(n8921), .B(n8920), .ZN(n8922)
         );
  AOI21_X1 U10114 ( .B1(n9253), .B2(n11077), .A(n8922), .ZN(n8923) );
  OAI21_X1 U10115 ( .B1(n8924), .B2(n11072), .A(n8923), .ZN(P2_U3156) );
  OAI211_X1 U10116 ( .C1(n8927), .C2(n8926), .A(n8925), .B(n9011), .ZN(n8933)
         );
  INV_X1 U10117 ( .A(n8928), .ZN(n8929) );
  AOI21_X1 U10118 ( .B1(n11077), .B2(n10930), .A(n8929), .ZN(n8932) );
  AOI22_X1 U10119 ( .A1(n9034), .A2(n9070), .B1(n9048), .B2(n9072), .ZN(n8931)
         );
  OR2_X1 U10120 ( .A1(n11079), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8930) );
  NAND4_X1 U10121 ( .A1(n8933), .A2(n8932), .A3(n8931), .A4(n8930), .ZN(
        P2_U3158) );
  INV_X1 U10122 ( .A(n8934), .ZN(n9490) );
  OAI211_X1 U10123 ( .C1(n8937), .C2(n8936), .A(n8935), .B(n9011), .ZN(n8943)
         );
  NAND2_X1 U10124 ( .A1(n9304), .A2(n9034), .ZN(n8939) );
  OAI211_X1 U10125 ( .C1(n9037), .C2(n8940), .A(n8939), .B(n8938), .ZN(n8941)
         );
  AOI21_X1 U10126 ( .B1(n9053), .B2(n9309), .A(n8941), .ZN(n8942) );
  OAI211_X1 U10127 ( .C1(n9490), .C2(n9056), .A(n8943), .B(n8942), .ZN(
        P2_U3159) );
  XOR2_X1 U10128 ( .A(n8945), .B(n8944), .Z(n8954) );
  INV_X1 U10129 ( .A(n8946), .ZN(n9281) );
  OR2_X1 U10130 ( .A1(n8947), .A2(n9289), .ZN(n8949) );
  NAND2_X1 U10131 ( .A1(n9304), .A2(n9363), .ZN(n8948) );
  NAND2_X1 U10132 ( .A1(n8949), .A2(n8948), .ZN(n9279) );
  AOI22_X1 U10133 ( .A1(n9279), .A2(n8950), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8951) );
  OAI21_X1 U10134 ( .B1(n9281), .B2(n11079), .A(n8951), .ZN(n8952) );
  AOI21_X1 U10135 ( .B1(n8628), .B2(n11077), .A(n8952), .ZN(n8953) );
  OAI21_X1 U10136 ( .B1(n8954), .B2(n11072), .A(n8953), .ZN(P2_U3163) );
  XOR2_X1 U10137 ( .A(n8958), .B(n8957), .Z(n8963) );
  AOI22_X1 U10138 ( .A1(n9248), .A2(n9048), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8960) );
  NAND2_X1 U10139 ( .A1(n9227), .A2(n9053), .ZN(n8959) );
  OAI211_X1 U10140 ( .C1(n9224), .C2(n9050), .A(n8960), .B(n8959), .ZN(n8961)
         );
  AOI21_X1 U10141 ( .B1(n9220), .B2(n11077), .A(n8961), .ZN(n8962) );
  OAI21_X1 U10142 ( .B1(n8963), .B2(n11072), .A(n8962), .ZN(P2_U3165) );
  INV_X1 U10143 ( .A(n8964), .ZN(n9499) );
  OAI211_X1 U10144 ( .C1(n8967), .C2(n8966), .A(n8965), .B(n9011), .ZN(n8972)
         );
  NAND2_X1 U10145 ( .A1(n9060), .A2(n9363), .ZN(n8969) );
  NAND2_X1 U10146 ( .A1(n9316), .A2(n7120), .ZN(n8968) );
  AND2_X1 U10147 ( .A1(n8969), .A2(n8968), .ZN(n9349) );
  NAND2_X1 U10148 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9136) );
  OAI21_X1 U10149 ( .B1(n9349), .B2(n11067), .A(n9136), .ZN(n8970) );
  AOI21_X1 U10150 ( .B1(n9351), .B2(n9053), .A(n8970), .ZN(n8971) );
  OAI211_X1 U10151 ( .C1(n9499), .C2(n9056), .A(n8972), .B(n8971), .ZN(
        P2_U3166) );
  INV_X1 U10152 ( .A(n8973), .ZN(n8974) );
  AOI21_X1 U10153 ( .B1(n8976), .B2(n8975), .A(n8974), .ZN(n8982) );
  NAND2_X1 U10154 ( .A1(n9361), .A2(n9363), .ZN(n8978) );
  NAND2_X1 U10155 ( .A1(n9303), .A2(n7120), .ZN(n8977) );
  AND2_X1 U10156 ( .A1(n8978), .A2(n8977), .ZN(n9332) );
  NAND2_X1 U10157 ( .A1(n9053), .A2(n9337), .ZN(n8979) );
  NAND2_X1 U10158 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9155) );
  OAI211_X1 U10159 ( .C1(n9332), .C2(n11067), .A(n8979), .B(n9155), .ZN(n8980)
         );
  AOI21_X1 U10160 ( .B1(n9336), .B2(n11077), .A(n8980), .ZN(n8981) );
  OAI21_X1 U10161 ( .B1(n8982), .B2(n11072), .A(n8981), .ZN(P2_U3168) );
  NAND2_X1 U10162 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  XOR2_X1 U10163 ( .A(n8986), .B(n8985), .Z(n8991) );
  AOI22_X1 U10164 ( .A1(n9260), .A2(n9048), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8988) );
  NAND2_X1 U10165 ( .A1(n9240), .A2(n9053), .ZN(n8987) );
  OAI211_X1 U10166 ( .C1(n9237), .C2(n9050), .A(n8988), .B(n8987), .ZN(n8989)
         );
  AOI21_X1 U10167 ( .B1(n9232), .B2(n11077), .A(n8989), .ZN(n8990) );
  OAI21_X1 U10168 ( .B1(n8991), .B2(n11072), .A(n8990), .ZN(P2_U3169) );
  INV_X1 U10169 ( .A(n8992), .ZN(n8993) );
  AOI21_X1 U10170 ( .B1(n8995), .B2(n8994), .A(n8993), .ZN(n9000) );
  NAND2_X1 U10171 ( .A1(n9053), .A2(n9296), .ZN(n8997) );
  AOI22_X1 U10172 ( .A1(n9261), .A2(n9034), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8996) );
  OAI211_X1 U10173 ( .C1(n9290), .C2(n9037), .A(n8997), .B(n8996), .ZN(n8998)
         );
  AOI21_X1 U10174 ( .B1(n9295), .B2(n11077), .A(n8998), .ZN(n8999) );
  OAI21_X1 U10175 ( .B1(n9000), .B2(n11072), .A(n8999), .ZN(P2_U3173) );
  NAND2_X1 U10176 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  XOR2_X1 U10177 ( .A(n9003), .B(n8908), .Z(n9010) );
  NAND2_X1 U10178 ( .A1(n9053), .A2(n9004), .ZN(n9006) );
  INV_X1 U10179 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10576) );
  NOR2_X1 U10180 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10576), .ZN(n9081) );
  AOI21_X1 U10181 ( .B1(n9034), .B2(n9362), .A(n9081), .ZN(n9005) );
  OAI211_X1 U10182 ( .C1(n9007), .C2(n9037), .A(n9006), .B(n9005), .ZN(n9008)
         );
  AOI21_X1 U10183 ( .B1(n11122), .B2(n11077), .A(n9008), .ZN(n9009) );
  OAI21_X1 U10184 ( .B1(n9010), .B2(n11072), .A(n9009), .ZN(P2_U3174) );
  INV_X1 U10185 ( .A(n9411), .ZN(n9019) );
  OAI211_X1 U10186 ( .C1(n9014), .C2(n9013), .A(n9012), .B(n9011), .ZN(n9018)
         );
  AOI22_X1 U10187 ( .A1(n9261), .A2(n9048), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n9015) );
  OAI21_X1 U10188 ( .B1(n9238), .B2(n9050), .A(n9015), .ZN(n9016) );
  AOI21_X1 U10189 ( .B1(n9266), .B2(n9053), .A(n9016), .ZN(n9017) );
  OAI211_X1 U10190 ( .C1(n9019), .C2(n9056), .A(n9018), .B(n9017), .ZN(
        P2_U3175) );
  INV_X1 U10191 ( .A(n9428), .ZN(n9029) );
  AOI21_X1 U10192 ( .B1(n9021), .B2(n9020), .A(n11072), .ZN(n9023) );
  NAND2_X1 U10193 ( .A1(n9023), .A2(n9022), .ZN(n9028) );
  NAND2_X1 U10194 ( .A1(n9048), .A2(n9316), .ZN(n9025) );
  OAI211_X1 U10195 ( .C1(n9290), .C2(n9050), .A(n9025), .B(n9024), .ZN(n9026)
         );
  AOI21_X1 U10196 ( .B1(n9053), .B2(n9320), .A(n9026), .ZN(n9027) );
  OAI211_X1 U10197 ( .C1(n9029), .C2(n9056), .A(n9028), .B(n9027), .ZN(
        P2_U3178) );
  NAND2_X1 U10198 ( .A1(n9031), .A2(n9030), .ZN(n9032) );
  XOR2_X1 U10199 ( .A(n9033), .B(n9032), .Z(n9040) );
  AOI22_X1 U10200 ( .A1(n9034), .A2(n9180), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n9036) );
  NAND2_X1 U10201 ( .A1(n9212), .A2(n9053), .ZN(n9035) );
  OAI211_X1 U10202 ( .C1(n9237), .C2(n9037), .A(n9036), .B(n9035), .ZN(n9038)
         );
  AOI21_X1 U10203 ( .B1(n9392), .B2(n11077), .A(n9038), .ZN(n9039) );
  OAI21_X1 U10204 ( .B1(n9040), .B2(n11072), .A(n9039), .ZN(P2_U3180) );
  INV_X1 U10205 ( .A(n9370), .ZN(n9504) );
  NAND2_X1 U10206 ( .A1(n8908), .A2(n9041), .ZN(n9043) );
  AND2_X1 U10207 ( .A1(n9043), .A2(n9042), .ZN(n9045) );
  AOI21_X1 U10208 ( .B1(n9045), .B2(n9044), .A(n11072), .ZN(n9047) );
  NAND2_X1 U10209 ( .A1(n9047), .A2(n9046), .ZN(n9055) );
  INV_X1 U10210 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10673) );
  NOR2_X1 U10211 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10673), .ZN(n9120) );
  AOI21_X1 U10212 ( .B1(n9048), .B2(n9362), .A(n9120), .ZN(n9049) );
  OAI21_X1 U10213 ( .B1(n9051), .B2(n9050), .A(n9049), .ZN(n9052) );
  AOI21_X1 U10214 ( .B1(n9053), .B2(n9366), .A(n9052), .ZN(n9054) );
  OAI211_X1 U10215 ( .C1(n9504), .C2(n9056), .A(n9055), .B(n9054), .ZN(
        P2_U3181) );
  MUX2_X1 U10216 ( .A(n9172), .B(P2_DATAO_REG_31__SCAN_IN), .S(n9073), .Z(
        P2_U3522) );
  MUX2_X1 U10217 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n5438), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10218 ( .A(n9058), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9073), .Z(
        P2_U3519) );
  MUX2_X1 U10219 ( .A(n9180), .B(P2_DATAO_REG_27__SCAN_IN), .S(n9073), .Z(
        P2_U3518) );
  MUX2_X1 U10220 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9059), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10221 ( .A(n9207), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9073), .Z(
        P2_U3516) );
  MUX2_X1 U10222 ( .A(n9248), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9073), .Z(
        P2_U3515) );
  MUX2_X1 U10223 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9247), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10224 ( .A(n9261), .B(P2_DATAO_REG_21__SCAN_IN), .S(n9073), .Z(
        P2_U3512) );
  MUX2_X1 U10225 ( .A(n9304), .B(P2_DATAO_REG_20__SCAN_IN), .S(n9073), .Z(
        P2_U3511) );
  MUX2_X1 U10226 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9317), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10227 ( .A(n9303), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9073), .Z(
        P2_U3509) );
  MUX2_X1 U10228 ( .A(n9316), .B(P2_DATAO_REG_17__SCAN_IN), .S(n9073), .Z(
        P2_U3508) );
  MUX2_X1 U10229 ( .A(n9361), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9073), .Z(
        P2_U3507) );
  MUX2_X1 U10230 ( .A(n9060), .B(P2_DATAO_REG_15__SCAN_IN), .S(n9073), .Z(
        P2_U3506) );
  MUX2_X1 U10231 ( .A(n9362), .B(P2_DATAO_REG_14__SCAN_IN), .S(n9073), .Z(
        P2_U3505) );
  MUX2_X1 U10232 ( .A(n9061), .B(P2_DATAO_REG_13__SCAN_IN), .S(n9073), .Z(
        P2_U3504) );
  MUX2_X1 U10233 ( .A(n9062), .B(P2_DATAO_REG_12__SCAN_IN), .S(n9073), .Z(
        P2_U3503) );
  MUX2_X1 U10234 ( .A(n9063), .B(P2_DATAO_REG_11__SCAN_IN), .S(n9073), .Z(
        P2_U3502) );
  MUX2_X1 U10235 ( .A(n9064), .B(P2_DATAO_REG_10__SCAN_IN), .S(n9073), .Z(
        P2_U3501) );
  MUX2_X1 U10236 ( .A(n9065), .B(P2_DATAO_REG_9__SCAN_IN), .S(n9073), .Z(
        P2_U3500) );
  MUX2_X1 U10237 ( .A(n9066), .B(P2_DATAO_REG_8__SCAN_IN), .S(n9073), .Z(
        P2_U3499) );
  MUX2_X1 U10238 ( .A(n9067), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9073), .Z(
        P2_U3498) );
  MUX2_X1 U10239 ( .A(n9068), .B(P2_DATAO_REG_6__SCAN_IN), .S(n9073), .Z(
        P2_U3497) );
  MUX2_X1 U10240 ( .A(n9069), .B(P2_DATAO_REG_5__SCAN_IN), .S(n9073), .Z(
        P2_U3496) );
  MUX2_X1 U10241 ( .A(n9070), .B(P2_DATAO_REG_4__SCAN_IN), .S(n9073), .Z(
        P2_U3495) );
  MUX2_X1 U10242 ( .A(n9071), .B(P2_DATAO_REG_3__SCAN_IN), .S(n9073), .Z(
        P2_U3494) );
  MUX2_X1 U10243 ( .A(n9072), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9073), .Z(
        P2_U3493) );
  MUX2_X1 U10244 ( .A(n9074), .B(P2_DATAO_REG_0__SCAN_IN), .S(n9073), .Z(
        P2_U3491) );
  AOI21_X1 U10245 ( .B1(n9076), .B2(n8306), .A(n9075), .ZN(n9090) );
  OAI21_X1 U10246 ( .B1(n9078), .B2(P2_REG1_REG_13__SCAN_IN), .A(n9077), .ZN(
        n9082) );
  INV_X1 U10247 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9079) );
  NOR2_X1 U10248 ( .A1(n9158), .A2(n9079), .ZN(n9080) );
  AOI211_X1 U10249 ( .C1(n9117), .C2(n9082), .A(n9081), .B(n9080), .ZN(n9089)
         );
  OAI21_X1 U10250 ( .B1(n9085), .B2(n9084), .A(n9083), .ZN(n9086) );
  AOI22_X1 U10251 ( .A1(n9166), .A2(n9087), .B1(n10352), .B2(n9086), .ZN(n9088) );
  OAI211_X1 U10252 ( .C1(n9090), .C2(n10348), .A(n9089), .B(n9088), .ZN(
        P2_U3195) );
  AOI21_X1 U10253 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9110) );
  AOI21_X1 U10254 ( .B1(n9096), .B2(n9095), .A(n9094), .ZN(n9107) );
  OAI21_X1 U10255 ( .B1(n9099), .B2(n9098), .A(n9097), .ZN(n9103) );
  INV_X1 U10256 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9101) );
  OAI21_X1 U10257 ( .B1(n9158), .B2(n9101), .A(n9100), .ZN(n9102) );
  AOI21_X1 U10258 ( .B1(n10352), .B2(n9103), .A(n9102), .ZN(n9106) );
  NAND2_X1 U10259 ( .A1(n9166), .A2(n9104), .ZN(n9105) );
  OAI211_X1 U10260 ( .C1(n9107), .C2(n10346), .A(n9106), .B(n9105), .ZN(n9108)
         );
  INV_X1 U10261 ( .A(n9108), .ZN(n9109) );
  OAI21_X1 U10262 ( .B1(n9110), .B2(n10348), .A(n9109), .ZN(P2_U3196) );
  AOI21_X1 U10263 ( .B1(n9368), .B2(n9112), .A(n9111), .ZN(n9129) );
  OAI21_X1 U10264 ( .B1(n9115), .B2(n9114), .A(n9113), .ZN(n9127) );
  INV_X1 U10265 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9123) );
  AND2_X1 U10266 ( .A1(n9116), .A2(n9443), .ZN(n9118) );
  OAI21_X1 U10267 ( .B1(n9119), .B2(n9118), .A(n9117), .ZN(n9122) );
  INV_X1 U10268 ( .A(n9120), .ZN(n9121) );
  OAI211_X1 U10269 ( .C1(n9123), .C2(n9158), .A(n9122), .B(n9121), .ZN(n9126)
         );
  NOR2_X1 U10270 ( .A1(n10357), .A2(n9124), .ZN(n9125) );
  AOI211_X1 U10271 ( .C1(n10352), .C2(n9127), .A(n9126), .B(n9125), .ZN(n9128)
         );
  OAI21_X1 U10272 ( .B1(n9129), .B2(n10348), .A(n9128), .ZN(P2_U3197) );
  AOI21_X1 U10273 ( .B1(n5144), .B2(n9131), .A(n9130), .ZN(n9147) );
  INV_X1 U10274 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9138) );
  OAI21_X1 U10275 ( .B1(n9134), .B2(n9133), .A(n9132), .ZN(n9135) );
  NAND2_X1 U10276 ( .A1(n9135), .A2(n10352), .ZN(n9137) );
  OAI211_X1 U10277 ( .C1(n9158), .C2(n9138), .A(n9137), .B(n9136), .ZN(n9144)
         );
  AOI21_X1 U10278 ( .B1(n9141), .B2(n9140), .A(n9139), .ZN(n9142) );
  NOR2_X1 U10279 ( .A1(n9142), .A2(n10346), .ZN(n9143) );
  AOI211_X1 U10280 ( .C1(n9166), .C2(n9145), .A(n9144), .B(n9143), .ZN(n9146)
         );
  OAI21_X1 U10281 ( .B1(n9147), .B2(n10348), .A(n9146), .ZN(P2_U3198) );
  AOI21_X1 U10282 ( .B1(n9150), .B2(n9149), .A(n9148), .ZN(n9168) );
  INV_X1 U10283 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9157) );
  OAI21_X1 U10284 ( .B1(n9153), .B2(n9152), .A(n9151), .ZN(n9154) );
  NAND2_X1 U10285 ( .A1(n9154), .A2(n10352), .ZN(n9156) );
  OAI211_X1 U10286 ( .C1(n9158), .C2(n9157), .A(n9156), .B(n9155), .ZN(n9164)
         );
  INV_X1 U10287 ( .A(n9159), .ZN(n9162) );
  NAND2_X1 U10288 ( .A1(n9160), .A2(n9434), .ZN(n9161) );
  AOI211_X1 U10289 ( .C1(n9166), .C2(n9165), .A(n9164), .B(n9163), .ZN(n9167)
         );
  OAI21_X1 U10290 ( .B1(n9168), .B2(n10348), .A(n9167), .ZN(P2_U3199) );
  AND2_X1 U10291 ( .A1(n11111), .A2(n9169), .ZN(n9173) );
  INV_X1 U10292 ( .A(n9170), .ZN(n9171) );
  NAND2_X1 U10293 ( .A1(n9172), .A2(n9171), .ZN(n9453) );
  NAND2_X1 U10294 ( .A1(n9173), .A2(n9453), .ZN(n9176) );
  OAI21_X1 U10295 ( .B1(n11111), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9176), .ZN(
        n9174) );
  OAI21_X1 U10296 ( .B1(n9455), .B2(n9354), .A(n9174), .ZN(P2_U3202) );
  OAI21_X1 U10297 ( .B1(n11111), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9176), .ZN(
        n9177) );
  OAI21_X1 U10298 ( .B1(n9458), .B2(n9354), .A(n9177), .ZN(P2_U3203) );
  XNOR2_X1 U10299 ( .A(n9178), .B(n9183), .ZN(n9179) );
  NAND2_X1 U10300 ( .A1(n9179), .A2(n9358), .ZN(n9182) );
  AOI22_X1 U10301 ( .A1(n5438), .A2(n7120), .B1(n9363), .B2(n9180), .ZN(n9181)
         );
  OR2_X1 U10302 ( .A1(n9184), .A2(n9183), .ZN(n9185) );
  NAND2_X1 U10303 ( .A1(n9186), .A2(n9185), .ZN(n9383) );
  AOI22_X1 U10304 ( .A1(n9352), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n11086), 
        .B2(n9187), .ZN(n9188) );
  OAI21_X1 U10305 ( .B1(n9385), .B2(n9354), .A(n9188), .ZN(n9189) );
  AOI21_X1 U10306 ( .B1(n9383), .B2(n11104), .A(n9189), .ZN(n9190) );
  OAI21_X1 U10307 ( .B1(n5147), .B2(n9352), .A(n9190), .ZN(P2_U3205) );
  XNOR2_X1 U10308 ( .A(n9192), .B(n9191), .ZN(n9197) );
  INV_X1 U10309 ( .A(n9388), .ZN(n9204) );
  XNOR2_X1 U10310 ( .A(n9199), .B(n9198), .ZN(n9389) );
  AOI22_X1 U10311 ( .A1(n9352), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n11086), 
        .B2(n9200), .ZN(n9201) );
  OAI21_X1 U10312 ( .B1(n9464), .B2(n9354), .A(n9201), .ZN(n9202) );
  AOI21_X1 U10313 ( .B1(n9389), .B2(n11104), .A(n9202), .ZN(n9203) );
  OAI21_X1 U10314 ( .B1(n9204), .B2(n9352), .A(n9203), .ZN(P2_U3206) );
  XNOR2_X1 U10315 ( .A(n9206), .B(n9205), .ZN(n9211) );
  NAND2_X1 U10316 ( .A1(n9207), .A2(n9363), .ZN(n9208) );
  OAI21_X1 U10317 ( .B1(n9209), .B2(n9289), .A(n9208), .ZN(n9210) );
  INV_X1 U10318 ( .A(n9212), .ZN(n9214) );
  OAI22_X1 U10319 ( .A1(n9214), .A2(n11102), .B1(n11111), .B2(n9213), .ZN(
        n9215) );
  AOI21_X1 U10320 ( .B1(n9392), .B2(n11106), .A(n9215), .ZN(n9219) );
  NAND2_X1 U10321 ( .A1(n9217), .A2(n9216), .ZN(n9393) );
  NAND3_X1 U10322 ( .A1(n9394), .A2(n9393), .A3(n11104), .ZN(n9218) );
  OAI211_X1 U10323 ( .C1(n9396), .C2(n9352), .A(n9219), .B(n9218), .ZN(
        P2_U3207) );
  INV_X1 U10324 ( .A(n9220), .ZN(n9472) );
  NOR2_X1 U10325 ( .A1(n9472), .A2(n9233), .ZN(n9226) );
  XNOR2_X1 U10326 ( .A(n9222), .B(n9221), .ZN(n9223) );
  OAI222_X1 U10327 ( .A1(n9291), .A2(n9225), .B1(n9289), .B2(n9224), .C1(n9287), .C2(n9223), .ZN(n9399) );
  AOI211_X1 U10328 ( .C1(n11086), .C2(n9227), .A(n9226), .B(n9399), .ZN(n9231)
         );
  XNOR2_X1 U10329 ( .A(n9229), .B(n9228), .ZN(n9400) );
  AOI22_X1 U10330 ( .A1(n9400), .A2(n11104), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n9352), .ZN(n9230) );
  OAI21_X1 U10331 ( .B1(n9231), .B2(n9352), .A(n9230), .ZN(P2_U3208) );
  INV_X1 U10332 ( .A(n9232), .ZN(n9476) );
  NOR2_X1 U10333 ( .A1(n9476), .A2(n9233), .ZN(n9239) );
  NAND2_X1 U10334 ( .A1(n9245), .A2(n9234), .ZN(n9235) );
  XOR2_X1 U10335 ( .A(n9242), .B(n9235), .Z(n9236) );
  OAI222_X1 U10336 ( .A1(n9291), .A2(n9238), .B1(n9289), .B2(n9237), .C1(n9287), .C2(n9236), .ZN(n9403) );
  AOI211_X1 U10337 ( .C1(n11086), .C2(n9240), .A(n9239), .B(n9403), .ZN(n9244)
         );
  XOR2_X1 U10338 ( .A(n9242), .B(n9241), .Z(n9404) );
  AOI22_X1 U10339 ( .A1(n9404), .A2(n11104), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n9352), .ZN(n9243) );
  OAI21_X1 U10340 ( .B1(n9244), .B2(n9352), .A(n9243), .ZN(P2_U3209) );
  OAI211_X1 U10341 ( .C1(n5172), .C2(n9246), .A(n9358), .B(n9245), .ZN(n9250)
         );
  AOI22_X1 U10342 ( .A1(n9248), .A2(n7120), .B1(n9247), .B2(n9363), .ZN(n9249)
         );
  NAND2_X1 U10343 ( .A1(n9250), .A2(n9249), .ZN(n9407) );
  INV_X1 U10344 ( .A(n9407), .ZN(n9258) );
  XNOR2_X1 U10345 ( .A(n9252), .B(n9251), .ZN(n9408) );
  INV_X1 U10346 ( .A(n9253), .ZN(n9480) );
  AOI22_X1 U10347 ( .A1(n9254), .A2(n11086), .B1(n9352), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n9255) );
  OAI21_X1 U10348 ( .B1(n9480), .B2(n9354), .A(n9255), .ZN(n9256) );
  AOI21_X1 U10349 ( .B1(n9408), .B2(n11104), .A(n9256), .ZN(n9257) );
  OAI21_X1 U10350 ( .B1(n9258), .B2(n9352), .A(n9257), .ZN(P2_U3210) );
  XNOR2_X1 U10351 ( .A(n9259), .B(n9264), .ZN(n9262) );
  AOI222_X1 U10352 ( .A1(n9358), .A2(n9262), .B1(n9261), .B2(n9363), .C1(n9260), .C2(n7120), .ZN(n9414) );
  NAND2_X1 U10353 ( .A1(n9275), .A2(n9263), .ZN(n9265) );
  XNOR2_X1 U10354 ( .A(n9265), .B(n9264), .ZN(n9412) );
  NAND2_X1 U10355 ( .A1(n9411), .A2(n11106), .ZN(n9268) );
  AOI22_X1 U10356 ( .A1(n9352), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9266), .B2(
        n11086), .ZN(n9267) );
  NAND2_X1 U10357 ( .A1(n9268), .A2(n9267), .ZN(n9269) );
  AOI21_X1 U10358 ( .B1(n9412), .B2(n11104), .A(n9269), .ZN(n9270) );
  OAI21_X1 U10359 ( .B1(n9414), .B2(n9352), .A(n9270), .ZN(P2_U3211) );
  NAND2_X1 U10360 ( .A1(n9271), .A2(n9272), .ZN(n9274) );
  NAND2_X1 U10361 ( .A1(n9274), .A2(n9273), .ZN(n9276) );
  OAI21_X1 U10362 ( .B1(n9276), .B2(n9277), .A(n9275), .ZN(n9417) );
  XOR2_X1 U10363 ( .A(n9278), .B(n9277), .Z(n9280) );
  AOI21_X1 U10364 ( .B1(n9280), .B2(n9358), .A(n9279), .ZN(n9416) );
  OAI21_X1 U10365 ( .B1(n9281), .B2(n11102), .A(n9416), .ZN(n9282) );
  NAND2_X1 U10366 ( .A1(n9282), .A2(n11111), .ZN(n9284) );
  AOI22_X1 U10367 ( .A1(n8628), .A2(n11106), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n9352), .ZN(n9283) );
  OAI211_X1 U10368 ( .C1(n9417), .C2(n7361), .A(n9284), .B(n9283), .ZN(
        P2_U3212) );
  AOI21_X1 U10369 ( .B1(n9293), .B2(n9285), .A(n5153), .ZN(n9286) );
  OAI222_X1 U10370 ( .A1(n9291), .A2(n9290), .B1(n9289), .B2(n9288), .C1(n9287), .C2(n9286), .ZN(n9418) );
  INV_X1 U10371 ( .A(n9418), .ZN(n9300) );
  NAND2_X1 U10372 ( .A1(n9271), .A2(n9292), .ZN(n9294) );
  XNOR2_X1 U10373 ( .A(n9294), .B(n9293), .ZN(n9419) );
  INV_X1 U10374 ( .A(n9295), .ZN(n9486) );
  AOI22_X1 U10375 ( .A1(n9352), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n11086), 
        .B2(n9296), .ZN(n9297) );
  OAI21_X1 U10376 ( .B1(n9486), .B2(n9354), .A(n9297), .ZN(n9298) );
  AOI21_X1 U10377 ( .B1(n9419), .B2(n11104), .A(n9298), .ZN(n9299) );
  OAI21_X1 U10378 ( .B1(n9300), .B2(n9352), .A(n9299), .ZN(P2_U3213) );
  OAI211_X1 U10379 ( .C1(n9302), .C2(n9307), .A(n9301), .B(n9358), .ZN(n9306)
         );
  AOI22_X1 U10380 ( .A1(n9304), .A2(n7120), .B1(n9363), .B2(n9303), .ZN(n9305)
         );
  NAND2_X1 U10381 ( .A1(n9306), .A2(n9305), .ZN(n9422) );
  INV_X1 U10382 ( .A(n9422), .ZN(n9313) );
  XNOR2_X1 U10383 ( .A(n9308), .B(n9307), .ZN(n9423) );
  AOI22_X1 U10384 ( .A1(n9352), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n11086), 
        .B2(n9309), .ZN(n9310) );
  OAI21_X1 U10385 ( .B1(n9490), .B2(n9354), .A(n9310), .ZN(n9311) );
  AOI21_X1 U10386 ( .B1(n9423), .B2(n11104), .A(n9311), .ZN(n9312) );
  OAI21_X1 U10387 ( .B1(n9313), .B2(n9352), .A(n9312), .ZN(P2_U3214) );
  OAI211_X1 U10388 ( .C1(n9315), .C2(n9324), .A(n9314), .B(n9358), .ZN(n9319)
         );
  AOI22_X1 U10389 ( .A1(n9317), .A2(n7120), .B1(n9363), .B2(n9316), .ZN(n9318)
         );
  NAND2_X1 U10390 ( .A1(n9319), .A2(n9318), .ZN(n9431) );
  INV_X1 U10391 ( .A(n9431), .ZN(n9328) );
  INV_X1 U10392 ( .A(n9320), .ZN(n9321) );
  OAI22_X1 U10393 ( .A1(n11111), .A2(n9322), .B1(n9321), .B2(n11102), .ZN(
        n9323) );
  AOI21_X1 U10394 ( .B1(n9428), .B2(n11106), .A(n9323), .ZN(n9327) );
  NAND2_X1 U10395 ( .A1(n9325), .A2(n9324), .ZN(n9426) );
  NAND3_X1 U10396 ( .A1(n9427), .A2(n9426), .A3(n11104), .ZN(n9326) );
  OAI211_X1 U10397 ( .C1(n9328), .C2(n9352), .A(n9327), .B(n9326), .ZN(
        P2_U3215) );
  NAND3_X1 U10398 ( .A1(n9346), .A2(n9334), .A3(n9329), .ZN(n9330) );
  NAND3_X1 U10399 ( .A1(n9331), .A2(n9358), .A3(n9330), .ZN(n9333) );
  NAND2_X1 U10400 ( .A1(n9333), .A2(n9332), .ZN(n9432) );
  INV_X1 U10401 ( .A(n9432), .ZN(n9341) );
  XNOR2_X1 U10402 ( .A(n9335), .B(n9334), .ZN(n9433) );
  INV_X1 U10403 ( .A(n9336), .ZN(n9495) );
  AOI22_X1 U10404 ( .A1(n9352), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n11086), 
        .B2(n9337), .ZN(n9338) );
  OAI21_X1 U10405 ( .B1(n9495), .B2(n9354), .A(n9338), .ZN(n9339) );
  AOI21_X1 U10406 ( .B1(n9433), .B2(n11104), .A(n9339), .ZN(n9340) );
  OAI21_X1 U10407 ( .B1(n9341), .B2(n9352), .A(n9340), .ZN(P2_U3216) );
  NAND2_X1 U10408 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  XNOR2_X1 U10409 ( .A(n9344), .B(n9348), .ZN(n9437) );
  INV_X1 U10410 ( .A(n9437), .ZN(n9357) );
  NAND2_X1 U10411 ( .A1(n9360), .A2(n9371), .ZN(n9359) );
  NAND2_X1 U10412 ( .A1(n9359), .A2(n9345), .ZN(n9347) );
  OAI211_X1 U10413 ( .C1(n9348), .C2(n9347), .A(n9346), .B(n9358), .ZN(n9350)
         );
  NAND2_X1 U10414 ( .A1(n9350), .A2(n9349), .ZN(n9436) );
  AOI22_X1 U10415 ( .A1(n9352), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n11086), 
        .B2(n9351), .ZN(n9353) );
  OAI21_X1 U10416 ( .B1(n9499), .B2(n9354), .A(n9353), .ZN(n9355) );
  AOI21_X1 U10417 ( .B1(n9436), .B2(n11111), .A(n9355), .ZN(n9356) );
  OAI21_X1 U10418 ( .B1(n9357), .B2(n7361), .A(n9356), .ZN(P2_U3217) );
  OAI211_X1 U10419 ( .C1(n9360), .C2(n9371), .A(n9359), .B(n9358), .ZN(n9365)
         );
  AOI22_X1 U10420 ( .A1(n9363), .A2(n9362), .B1(n9361), .B2(n7120), .ZN(n9364)
         );
  INV_X1 U10421 ( .A(n9366), .ZN(n9367) );
  OAI22_X1 U10422 ( .A1(n11111), .A2(n9368), .B1(n9367), .B2(n11102), .ZN(
        n9369) );
  AOI21_X1 U10423 ( .B1(n9370), .B2(n11106), .A(n9369), .ZN(n9374) );
  XNOR2_X1 U10424 ( .A(n9372), .B(n9371), .ZN(n9440) );
  NAND2_X1 U10425 ( .A1(n9440), .A2(n11104), .ZN(n9373) );
  OAI211_X1 U10426 ( .C1(n9442), .C2(n9352), .A(n9374), .B(n9373), .ZN(
        P2_U3218) );
  NOR2_X1 U10427 ( .A1(n11126), .A2(n9453), .ZN(n9376) );
  AOI21_X1 U10428 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n11126), .A(n9376), .ZN(
        n9375) );
  OAI21_X1 U10429 ( .B1(n9455), .B2(n9445), .A(n9375), .ZN(P2_U3490) );
  AOI21_X1 U10430 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n11126), .A(n9376), .ZN(
        n9377) );
  OAI21_X1 U10431 ( .B1(n9458), .B2(n9445), .A(n9377), .ZN(P2_U3489) );
  NAND2_X1 U10432 ( .A1(n9382), .A2(n9381), .ZN(n9459) );
  MUX2_X1 U10433 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9459), .S(n11127), .Z(
        P2_U3488) );
  NAND2_X1 U10434 ( .A1(n9383), .A2(n11119), .ZN(n9384) );
  OAI21_X1 U10435 ( .B1(n9385), .B2(n10987), .A(n9384), .ZN(n9386) );
  INV_X1 U10436 ( .A(n9386), .ZN(n9387) );
  MUX2_X1 U10437 ( .A(n9460), .B(P2_REG1_REG_28__SCAN_IN), .S(n11126), .Z(
        P2_U3487) );
  INV_X1 U10438 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9390) );
  AOI21_X1 U10439 ( .B1(n11119), .B2(n9389), .A(n9388), .ZN(n9461) );
  MUX2_X1 U10440 ( .A(n9390), .B(n9461), .S(n11127), .Z(n9391) );
  OAI21_X1 U10441 ( .B1(n9464), .B2(n9445), .A(n9391), .ZN(P2_U3486) );
  INV_X1 U10442 ( .A(n9392), .ZN(n9468) );
  INV_X1 U10443 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9397) );
  NAND3_X1 U10444 ( .A1(n9394), .A2(n9393), .A3(n11119), .ZN(n9395) );
  MUX2_X1 U10445 ( .A(n9397), .B(n9465), .S(n11127), .Z(n9398) );
  OAI21_X1 U10446 ( .B1(n9468), .B2(n9445), .A(n9398), .ZN(P2_U3485) );
  INV_X1 U10447 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9401) );
  AOI21_X1 U10448 ( .B1(n11119), .B2(n9400), .A(n9399), .ZN(n9469) );
  MUX2_X1 U10449 ( .A(n9401), .B(n9469), .S(n11127), .Z(n9402) );
  OAI21_X1 U10450 ( .B1(n9472), .B2(n9445), .A(n9402), .ZN(P2_U3484) );
  INV_X1 U10451 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9405) );
  AOI21_X1 U10452 ( .B1(n9404), .B2(n11119), .A(n9403), .ZN(n9473) );
  MUX2_X1 U10453 ( .A(n9405), .B(n9473), .S(n11127), .Z(n9406) );
  OAI21_X1 U10454 ( .B1(n9476), .B2(n9445), .A(n9406), .ZN(P2_U3483) );
  INV_X1 U10455 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9409) );
  AOI21_X1 U10456 ( .B1(n9408), .B2(n11119), .A(n9407), .ZN(n9477) );
  MUX2_X1 U10457 ( .A(n9409), .B(n9477), .S(n11127), .Z(n9410) );
  OAI21_X1 U10458 ( .B1(n9480), .B2(n9445), .A(n9410), .ZN(P2_U3482) );
  AOI22_X1 U10459 ( .A1(n9412), .A2(n11119), .B1(n11121), .B2(n9411), .ZN(
        n9413) );
  NAND2_X1 U10460 ( .A1(n9414), .A2(n9413), .ZN(n9481) );
  MUX2_X1 U10461 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9481), .S(n11127), .Z(
        P2_U3481) );
  INV_X1 U10462 ( .A(n11119), .ZN(n10938) );
  NAND2_X1 U10463 ( .A1(n8628), .A2(n11121), .ZN(n9415) );
  OAI211_X1 U10464 ( .C1(n10938), .C2(n9417), .A(n9416), .B(n9415), .ZN(n9482)
         );
  MUX2_X1 U10465 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9482), .S(n11127), .Z(
        P2_U3480) );
  INV_X1 U10466 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9420) );
  AOI21_X1 U10467 ( .B1(n9419), .B2(n11119), .A(n9418), .ZN(n9483) );
  MUX2_X1 U10468 ( .A(n9420), .B(n9483), .S(n11127), .Z(n9421) );
  OAI21_X1 U10469 ( .B1(n9486), .B2(n9445), .A(n9421), .ZN(P2_U3479) );
  INV_X1 U10470 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9424) );
  AOI21_X1 U10471 ( .B1(n11119), .B2(n9423), .A(n9422), .ZN(n9487) );
  MUX2_X1 U10472 ( .A(n9424), .B(n9487), .S(n11127), .Z(n9425) );
  OAI21_X1 U10473 ( .B1(n9490), .B2(n9445), .A(n9425), .ZN(P2_U3478) );
  AND3_X1 U10474 ( .A1(n9427), .A2(n11119), .A3(n9426), .ZN(n9430) );
  AND2_X1 U10475 ( .A1(n9428), .A2(n11121), .ZN(n9429) );
  MUX2_X1 U10476 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9491), .S(n11127), .Z(
        P2_U3477) );
  AOI21_X1 U10477 ( .B1(n9433), .B2(n11119), .A(n9432), .ZN(n9492) );
  MUX2_X1 U10478 ( .A(n9434), .B(n9492), .S(n11127), .Z(n9435) );
  OAI21_X1 U10479 ( .B1(n9495), .B2(n9445), .A(n9435), .ZN(P2_U3476) );
  AOI21_X1 U10480 ( .B1(n11119), .B2(n9437), .A(n9436), .ZN(n9496) );
  MUX2_X1 U10481 ( .A(n9438), .B(n9496), .S(n11127), .Z(n9439) );
  OAI21_X1 U10482 ( .B1(n9499), .B2(n9445), .A(n9439), .ZN(P2_U3475) );
  NAND2_X1 U10483 ( .A1(n9440), .A2(n11119), .ZN(n9441) );
  MUX2_X1 U10484 ( .A(n9443), .B(n9500), .S(n11127), .Z(n9444) );
  OAI21_X1 U10485 ( .B1(n9504), .B2(n9445), .A(n9444), .ZN(P2_U3474) );
  INV_X1 U10486 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9451) );
  NAND3_X1 U10487 ( .A1(n9446), .A2(n8701), .A3(n11119), .ZN(n9447) );
  OAI21_X1 U10488 ( .B1(n9448), .B2(n10987), .A(n9447), .ZN(n9449) );
  NOR2_X1 U10489 ( .A1(n9450), .A2(n9449), .ZN(n9505) );
  MUX2_X1 U10490 ( .A(n9451), .B(n9505), .S(n11127), .Z(n9452) );
  INV_X1 U10491 ( .A(n9452), .ZN(P2_U3473) );
  NOR2_X1 U10492 ( .A1(n11128), .A2(n9453), .ZN(n9456) );
  AOI21_X1 U10493 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(n11128), .A(n9456), .ZN(
        n9454) );
  OAI21_X1 U10494 ( .B1(n9455), .B2(n9503), .A(n9454), .ZN(P2_U3458) );
  AOI21_X1 U10495 ( .B1(P2_REG0_REG_30__SCAN_IN), .B2(n11128), .A(n9456), .ZN(
        n9457) );
  OAI21_X1 U10496 ( .B1(n9458), .B2(n9503), .A(n9457), .ZN(P2_U3457) );
  MUX2_X1 U10497 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9459), .S(n11131), .Z(
        P2_U3456) );
  MUX2_X1 U10498 ( .A(n9460), .B(P2_REG0_REG_28__SCAN_IN), .S(n11128), .Z(
        P2_U3455) );
  INV_X1 U10499 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9462) );
  MUX2_X1 U10500 ( .A(n9462), .B(n9461), .S(n11131), .Z(n9463) );
  OAI21_X1 U10501 ( .B1(n9464), .B2(n9503), .A(n9463), .ZN(P2_U3454) );
  INV_X1 U10502 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9466) );
  MUX2_X1 U10503 ( .A(n9466), .B(n9465), .S(n11131), .Z(n9467) );
  OAI21_X1 U10504 ( .B1(n9468), .B2(n9503), .A(n9467), .ZN(P2_U3453) );
  INV_X1 U10505 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9470) );
  MUX2_X1 U10506 ( .A(n9470), .B(n9469), .S(n11131), .Z(n9471) );
  OAI21_X1 U10507 ( .B1(n9472), .B2(n9503), .A(n9471), .ZN(P2_U3452) );
  INV_X1 U10508 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9474) );
  MUX2_X1 U10509 ( .A(n9474), .B(n9473), .S(n11131), .Z(n9475) );
  OAI21_X1 U10510 ( .B1(n9476), .B2(n9503), .A(n9475), .ZN(P2_U3451) );
  INV_X1 U10511 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9478) );
  MUX2_X1 U10512 ( .A(n9478), .B(n9477), .S(n11131), .Z(n9479) );
  OAI21_X1 U10513 ( .B1(n9480), .B2(n9503), .A(n9479), .ZN(P2_U3450) );
  MUX2_X1 U10514 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9481), .S(n11131), .Z(
        P2_U3449) );
  MUX2_X1 U10515 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9482), .S(n11131), .Z(
        P2_U3448) );
  MUX2_X1 U10516 ( .A(n9484), .B(n9483), .S(n11131), .Z(n9485) );
  OAI21_X1 U10517 ( .B1(n9486), .B2(n9503), .A(n9485), .ZN(P2_U3447) );
  INV_X1 U10518 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9488) );
  MUX2_X1 U10519 ( .A(n9488), .B(n9487), .S(n11131), .Z(n9489) );
  OAI21_X1 U10520 ( .B1(n9490), .B2(n9503), .A(n9489), .ZN(P2_U3446) );
  MUX2_X1 U10521 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9491), .S(n11131), .Z(
        P2_U3444) );
  INV_X1 U10522 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U10523 ( .A(n9493), .B(n9492), .S(n11131), .Z(n9494) );
  OAI21_X1 U10524 ( .B1(n9495), .B2(n9503), .A(n9494), .ZN(P2_U3441) );
  INV_X1 U10525 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9497) );
  MUX2_X1 U10526 ( .A(n9497), .B(n9496), .S(n11131), .Z(n9498) );
  OAI21_X1 U10527 ( .B1(n9499), .B2(n9503), .A(n9498), .ZN(P2_U3438) );
  INV_X1 U10528 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9501) );
  MUX2_X1 U10529 ( .A(n9501), .B(n9500), .S(n11131), .Z(n9502) );
  OAI21_X1 U10530 ( .B1(n9504), .B2(n9503), .A(n9502), .ZN(P2_U3435) );
  INV_X1 U10531 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9506) );
  MUX2_X1 U10532 ( .A(n9506), .B(n9505), .S(n11131), .Z(n9507) );
  INV_X1 U10533 ( .A(n9507), .ZN(P2_U3432) );
  MUX2_X1 U10534 ( .A(n9509), .B(P2_D_REG_1__SCAN_IN), .S(n9508), .Z(P2_U3377)
         );
  INV_X1 U10535 ( .A(n9645), .ZN(n10333) );
  NOR4_X1 U10536 ( .A1(n6770), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9510), .A4(
        P2_U3151), .ZN(n9511) );
  AOI21_X1 U10537 ( .B1(n9513), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9511), .ZN(
        n9512) );
  OAI21_X1 U10538 ( .B1(n10333), .B2(n9518), .A(n9512), .ZN(P2_U3264) );
  INV_X1 U10539 ( .A(n9734), .ZN(n10335) );
  AOI22_X1 U10540 ( .A1(n9514), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9513), .ZN(n9515) );
  OAI21_X1 U10541 ( .B1(n10335), .B2(n9518), .A(n9515), .ZN(P2_U3265) );
  INV_X1 U10542 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9517) );
  MUX2_X1 U10543 ( .A(n9520), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10544 ( .A(n9583), .ZN(n9524) );
  OAI21_X1 U10545 ( .B1(n9600), .B2(n9522), .A(n9521), .ZN(n9523) );
  AOI21_X1 U10546 ( .B1(n9524), .B2(n9523), .A(n9616), .ZN(n9528) );
  INV_X1 U10547 ( .A(n10273), .ZN(n10126) );
  AOI22_X1 U10548 ( .A1(n9640), .A2(n10133), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9526) );
  AOI22_X1 U10549 ( .A1(n9623), .A2(n10132), .B1(n9624), .B2(n10124), .ZN(
        n9525) );
  OAI211_X1 U10550 ( .C1(n10126), .C2(n9643), .A(n9526), .B(n9525), .ZN(n9527)
         );
  OR2_X1 U10551 ( .A1(n9528), .A2(n9527), .ZN(P1_U3216) );
  AOI21_X1 U10552 ( .B1(n9531), .B2(n9529), .A(n9530), .ZN(n9535) );
  INV_X1 U10553 ( .A(n10197), .ZN(n10161) );
  AOI22_X1 U10554 ( .A1(n9623), .A2(n10223), .B1(n9624), .B2(n10188), .ZN(
        n9532) );
  NAND2_X1 U10555 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9982) );
  OAI211_X1 U10556 ( .C1(n10161), .C2(n9605), .A(n9532), .B(n9982), .ZN(n9533)
         );
  AOI21_X1 U10557 ( .B1(n10293), .B2(n9625), .A(n9533), .ZN(n9534) );
  OAI21_X1 U10558 ( .B1(n9535), .B2(n9616), .A(n9534), .ZN(P1_U3219) );
  XNOR2_X1 U10559 ( .A(n9538), .B(n9537), .ZN(n9539) );
  XNOR2_X1 U10560 ( .A(n9536), .B(n9539), .ZN(n9540) );
  NAND2_X1 U10561 ( .A1(n9540), .A2(n9633), .ZN(n9547) );
  AOI21_X1 U10562 ( .B1(n9640), .B2(n9905), .A(n9541), .ZN(n9546) );
  AOI22_X1 U10563 ( .A1(n9623), .A2(n9907), .B1(n9624), .B2(n9542), .ZN(n9545)
         );
  NAND2_X1 U10564 ( .A1(n9625), .A2(n9543), .ZN(n9544) );
  NAND4_X1 U10565 ( .A1(n9547), .A2(n9546), .A3(n9545), .A4(n9544), .ZN(
        P1_U3221) );
  INV_X1 U10566 ( .A(n9548), .ZN(n9552) );
  OAI21_X1 U10567 ( .B1(n9590), .B2(n9550), .A(n9549), .ZN(n9551) );
  NAND3_X1 U10568 ( .A1(n9552), .A2(n9633), .A3(n9551), .ZN(n9556) );
  AOI22_X1 U10569 ( .A1(n9623), .A2(n10197), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9555) );
  AOI22_X1 U10570 ( .A1(n9640), .A2(n10132), .B1(n9624), .B2(n10165), .ZN(
        n9554) );
  NAND2_X1 U10571 ( .A1(n10284), .A2(n9625), .ZN(n9553) );
  NAND4_X1 U10572 ( .A1(n9556), .A2(n9555), .A3(n9554), .A4(n9553), .ZN(
        P1_U3223) );
  OAI21_X1 U10573 ( .B1(n9558), .B2(n9557), .A(n9619), .ZN(n9559) );
  NAND2_X1 U10574 ( .A1(n9559), .A2(n9633), .ZN(n9563) );
  AOI22_X1 U10575 ( .A1(n9640), .A2(n10060), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9562) );
  AOI22_X1 U10576 ( .A1(n9623), .A2(n10133), .B1(n9624), .B2(n10090), .ZN(
        n9561) );
  NAND2_X1 U10577 ( .A1(n10263), .A2(n9625), .ZN(n9560) );
  NAND4_X1 U10578 ( .A1(n9563), .A2(n9562), .A3(n9561), .A4(n9560), .ZN(
        P1_U3225) );
  XOR2_X1 U10579 ( .A(n9564), .B(n9565), .Z(n9570) );
  INV_X1 U10580 ( .A(n10016), .ZN(n10208) );
  AOI22_X1 U10581 ( .A1(n9623), .A2(n9899), .B1(n9624), .B2(n9566), .ZN(n9567)
         );
  NAND2_X1 U10582 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n9920) );
  OAI211_X1 U10583 ( .C1(n10208), .C2(n9605), .A(n9567), .B(n9920), .ZN(n9568)
         );
  AOI21_X1 U10584 ( .B1(n10303), .B2(n9625), .A(n9568), .ZN(n9569) );
  OAI21_X1 U10585 ( .B1(n9570), .B2(n9616), .A(n9569), .ZN(P1_U3226) );
  INV_X1 U10586 ( .A(n10234), .ZN(n11142) );
  XNOR2_X1 U10587 ( .A(n9572), .B(n9571), .ZN(n9573) );
  XNOR2_X1 U10588 ( .A(n9574), .B(n9573), .ZN(n9575) );
  NAND2_X1 U10589 ( .A1(n9575), .A2(n9633), .ZN(n9579) );
  AND2_X1 U10590 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9950) );
  INV_X1 U10591 ( .A(n9576), .ZN(n10228) );
  OAI22_X1 U10592 ( .A1(n10013), .A2(n9637), .B1(n9636), .B2(n10228), .ZN(
        n9577) );
  AOI211_X1 U10593 ( .C1(n9640), .C2(n10223), .A(n9950), .B(n9577), .ZN(n9578)
         );
  OAI211_X1 U10594 ( .C1(n11142), .C2(n9643), .A(n9579), .B(n9578), .ZN(
        P1_U3228) );
  INV_X1 U10595 ( .A(n9580), .ZN(n9585) );
  NOR3_X1 U10596 ( .A1(n9583), .A2(n9582), .A3(n9581), .ZN(n9584) );
  OAI21_X1 U10597 ( .B1(n9585), .B2(n9584), .A(n9633), .ZN(n9589) );
  AOI22_X1 U10598 ( .A1(n9640), .A2(n9898), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9588) );
  AOI22_X1 U10599 ( .A1(n9623), .A2(n10147), .B1(n9624), .B2(n10109), .ZN(
        n9587) );
  NAND2_X1 U10600 ( .A1(n10268), .A2(n9625), .ZN(n9586) );
  NAND4_X1 U10601 ( .A1(n9589), .A2(n9588), .A3(n9587), .A4(n9586), .ZN(
        P1_U3229) );
  AOI21_X1 U10602 ( .B1(n9592), .B2(n9591), .A(n9590), .ZN(n9598) );
  INV_X1 U10603 ( .A(n10148), .ZN(n10178) );
  OAI22_X1 U10604 ( .A1(n9605), .A2(n10178), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9593), .ZN(n9596) );
  INV_X1 U10605 ( .A(n10017), .ZN(n10209) );
  INV_X1 U10606 ( .A(n9594), .ZN(n10172) );
  OAI22_X1 U10607 ( .A1(n10209), .A2(n9637), .B1(n9636), .B2(n10172), .ZN(
        n9595) );
  AOI211_X1 U10608 ( .C1(n10289), .C2(n9625), .A(n9596), .B(n9595), .ZN(n9597)
         );
  OAI21_X1 U10609 ( .B1(n9598), .B2(n9616), .A(n9597), .ZN(P1_U3233) );
  NOR2_X1 U10610 ( .A1(n9600), .A2(n9599), .ZN(n9601) );
  XOR2_X1 U10611 ( .A(n9602), .B(n9601), .Z(n9609) );
  OAI22_X1 U10612 ( .A1(n9637), .A2(n10178), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9603), .ZN(n9607) );
  INV_X1 U10613 ( .A(n10147), .ZN(n10116) );
  INV_X1 U10614 ( .A(n10141), .ZN(n9604) );
  OAI22_X1 U10615 ( .A1(n10116), .A2(n9605), .B1(n9636), .B2(n9604), .ZN(n9606) );
  AOI211_X1 U10616 ( .C1(n10277), .C2(n9625), .A(n9607), .B(n9606), .ZN(n9608)
         );
  OAI21_X1 U10617 ( .B1(n9609), .B2(n9616), .A(n9608), .ZN(P1_U3235) );
  XNOR2_X1 U10618 ( .A(n9611), .B(n5643), .ZN(n9612) );
  XNOR2_X1 U10619 ( .A(n9610), .B(n9612), .ZN(n9617) );
  AOI22_X1 U10620 ( .A1(n9640), .A2(n10017), .B1(n9624), .B2(n10213), .ZN(
        n9613) );
  NAND2_X1 U10621 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9960) );
  OAI211_X1 U10622 ( .C1(n10208), .C2(n9637), .A(n9613), .B(n9960), .ZN(n9614)
         );
  AOI21_X1 U10623 ( .B1(n10299), .B2(n9625), .A(n9614), .ZN(n9615) );
  OAI21_X1 U10624 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(P1_U3238) );
  AND2_X1 U10625 ( .A1(n9619), .A2(n9618), .ZN(n9622) );
  OAI211_X1 U10626 ( .C1(n9622), .C2(n9621), .A(n9633), .B(n9620), .ZN(n9629)
         );
  AOI22_X1 U10627 ( .A1(n9623), .A2(n9898), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9628) );
  AOI22_X1 U10628 ( .A1(n9640), .A2(n10051), .B1(n9624), .B2(n10082), .ZN(
        n9627) );
  NAND2_X1 U10629 ( .A1(n10259), .A2(n9625), .ZN(n9626) );
  NAND4_X1 U10630 ( .A1(n9629), .A2(n9628), .A3(n9627), .A4(n9626), .ZN(
        P1_U3240) );
  NAND2_X1 U10631 ( .A1(n5191), .A2(n9630), .ZN(n9632) );
  XNOR2_X1 U10632 ( .A(n9632), .B(n9631), .ZN(n9634) );
  NAND2_X1 U10633 ( .A1(n9634), .A2(n9633), .ZN(n9642) );
  OAI22_X1 U10634 ( .A1(n9688), .A2(n9637), .B1(n9636), .B2(n9635), .ZN(n9638)
         );
  AOI211_X1 U10635 ( .C1(n9640), .C2(n10222), .A(n9639), .B(n9638), .ZN(n9641)
         );
  OAI211_X1 U10636 ( .C1(n11134), .C2(n9643), .A(n9642), .B(n9641), .ZN(
        P1_U3241) );
  NAND2_X1 U10637 ( .A1(n9645), .A2(n9644), .ZN(n9647) );
  NAND2_X1 U10638 ( .A1(n5979), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9646) );
  NAND2_X1 U10639 ( .A1(n10239), .A2(n9991), .ZN(n9785) );
  NOR2_X1 U10640 ( .A1(n9841), .A2(n9648), .ZN(n9652) );
  NAND2_X1 U10641 ( .A1(n9650), .A2(n9649), .ZN(n9838) );
  OAI211_X1 U10642 ( .C1(n9652), .C2(n9838), .A(n9651), .B(n9844), .ZN(n9653)
         );
  AND2_X1 U10643 ( .A1(n9653), .A2(n9842), .ZN(n10965) );
  MUX2_X1 U10644 ( .A(n9654), .B(n10965), .S(n9742), .Z(n9659) );
  INV_X1 U10645 ( .A(n9655), .ZN(n9847) );
  NAND2_X1 U10646 ( .A1(n9847), .A2(n9846), .ZN(n9656) );
  MUX2_X1 U10647 ( .A(n9656), .B(n9846), .S(n9742), .Z(n9657) );
  OAI211_X1 U10648 ( .C1(n9659), .C2(n10966), .A(n9658), .B(n9657), .ZN(n9663)
         );
  INV_X1 U10649 ( .A(n11013), .ZN(n9662) );
  MUX2_X1 U10650 ( .A(n9851), .B(n9660), .S(n9747), .Z(n9661) );
  INV_X1 U10651 ( .A(n9679), .ZN(n9664) );
  NAND2_X1 U10652 ( .A1(n9664), .A2(n9853), .ZN(n9667) );
  INV_X1 U10653 ( .A(n9671), .ZN(n9665) );
  NAND2_X1 U10654 ( .A1(n9665), .A2(n9672), .ZN(n9666) );
  OAI21_X1 U10655 ( .B1(n9671), .B2(n9670), .A(n9669), .ZN(n9673) );
  NAND2_X1 U10656 ( .A1(n9673), .A2(n9672), .ZN(n9674) );
  NAND2_X1 U10657 ( .A1(n9674), .A2(n9853), .ZN(n9675) );
  NOR2_X1 U10658 ( .A1(n9676), .A2(n9675), .ZN(n9682) );
  OAI21_X1 U10659 ( .B1(n9679), .B2(n9678), .A(n9677), .ZN(n9681) );
  INV_X1 U10660 ( .A(n9684), .ZN(n9685) );
  NAND2_X1 U10661 ( .A1(n9687), .A2(n9685), .ZN(n9686) );
  NAND2_X1 U10662 ( .A1(n9694), .A2(n9687), .ZN(n9861) );
  OAI21_X1 U10663 ( .B1(n9696), .B2(n9861), .A(n9860), .ZN(n9690) );
  NAND2_X1 U10664 ( .A1(n10307), .A2(n9688), .ZN(n9698) );
  NAND2_X1 U10665 ( .A1(n9700), .A2(n9689), .ZN(n9697) );
  AOI21_X1 U10666 ( .B1(n9690), .B2(n9698), .A(n9697), .ZN(n9692) );
  NAND2_X1 U10667 ( .A1(n9864), .A2(n9701), .ZN(n9691) );
  OAI21_X1 U10668 ( .B1(n9692), .B2(n9691), .A(n9868), .ZN(n9707) );
  NAND2_X1 U10669 ( .A1(n9860), .A2(n9693), .ZN(n9695) );
  OAI21_X1 U10670 ( .B1(n9696), .B2(n9695), .A(n9694), .ZN(n9703) );
  INV_X1 U10671 ( .A(n9698), .ZN(n9699) );
  NAND2_X1 U10672 ( .A1(n9700), .A2(n9699), .ZN(n9702) );
  NAND2_X1 U10673 ( .A1(n9702), .A2(n9701), .ZN(n9863) );
  AOI21_X1 U10674 ( .B1(n9703), .B2(n5330), .A(n9863), .ZN(n9705) );
  INV_X1 U10675 ( .A(n9868), .ZN(n9704) );
  OAI21_X1 U10676 ( .B1(n9705), .B2(n9704), .A(n9864), .ZN(n9706) );
  MUX2_X1 U10677 ( .A(n9707), .B(n9706), .S(n9742), .Z(n9708) );
  OR2_X1 U10678 ( .A1(n10234), .A2(n10208), .ZN(n9869) );
  NAND2_X1 U10679 ( .A1(n10234), .A2(n10208), .ZN(n9759) );
  NAND2_X1 U10680 ( .A1(n9869), .A2(n9759), .ZN(n10226) );
  NOR2_X1 U10681 ( .A1(n9708), .A2(n10226), .ZN(n9711) );
  NAND2_X1 U10682 ( .A1(n9794), .A2(n9869), .ZN(n9710) );
  NAND2_X1 U10683 ( .A1(n10299), .A2(n9709), .ZN(n10192) );
  NAND2_X1 U10684 ( .A1(n10192), .A2(n9759), .ZN(n9832) );
  OR2_X1 U10685 ( .A1(n10293), .A2(n10209), .ZN(n9761) );
  NAND2_X1 U10686 ( .A1(n10293), .A2(n10209), .ZN(n9763) );
  INV_X1 U10687 ( .A(n9763), .ZN(n9877) );
  OR2_X1 U10688 ( .A1(n10289), .A2(n10161), .ZN(n9793) );
  NAND2_X1 U10689 ( .A1(n9793), .A2(n9761), .ZN(n9873) );
  NAND2_X1 U10690 ( .A1(n10289), .A2(n10161), .ZN(n10156) );
  NAND2_X1 U10691 ( .A1(n10156), .A2(n9763), .ZN(n9712) );
  MUX2_X1 U10692 ( .A(n9873), .B(n9712), .S(n9747), .Z(n9714) );
  OR2_X1 U10693 ( .A1(n10284), .A2(n10178), .ZN(n9874) );
  NAND2_X1 U10694 ( .A1(n10284), .A2(n10178), .ZN(n9766) );
  NAND2_X1 U10695 ( .A1(n9874), .A2(n9766), .ZN(n10158) );
  MUX2_X1 U10696 ( .A(n9793), .B(n10156), .S(n9742), .Z(n9713) );
  MUX2_X1 U10697 ( .A(n9874), .B(n9766), .S(n9747), .Z(n9715) );
  INV_X1 U10698 ( .A(n10132), .ZN(n10162) );
  NAND2_X1 U10699 ( .A1(n10277), .A2(n10162), .ZN(n9717) );
  AOI21_X1 U10700 ( .B1(n9716), .B2(n9715), .A(n10021), .ZN(n9719) );
  NOR2_X1 U10701 ( .A1(n10273), .A2(n10116), .ZN(n9792) );
  INV_X1 U10702 ( .A(n10001), .ZN(n10128) );
  OR2_X1 U10703 ( .A1(n9792), .A2(n10128), .ZN(n9752) );
  AND2_X1 U10704 ( .A1(n10273), .A2(n10116), .ZN(n9791) );
  INV_X1 U10705 ( .A(n9791), .ZN(n10003) );
  NAND2_X1 U10706 ( .A1(n10003), .A2(n9717), .ZN(n9768) );
  MUX2_X1 U10707 ( .A(n9752), .B(n9768), .S(n9747), .Z(n9718) );
  NOR2_X1 U10708 ( .A1(n9719), .A2(n9718), .ZN(n9721) );
  MUX2_X1 U10709 ( .A(n9791), .B(n9792), .S(n9747), .Z(n9720) );
  INV_X1 U10710 ( .A(n10133), .ZN(n10097) );
  NAND2_X1 U10711 ( .A1(n10268), .A2(n10097), .ZN(n9754) );
  NAND2_X1 U10712 ( .A1(n10004), .A2(n9754), .ZN(n10114) );
  NOR3_X1 U10713 ( .A1(n9721), .A2(n9720), .A3(n10114), .ZN(n9722) );
  NAND2_X1 U10714 ( .A1(n10263), .A2(n10115), .ZN(n9723) );
  INV_X1 U10715 ( .A(n10094), .ZN(n10088) );
  INV_X1 U10716 ( .A(n9754), .ZN(n9769) );
  INV_X1 U10717 ( .A(n10060), .ZN(n10096) );
  NAND2_X1 U10718 ( .A1(n10259), .A2(n10096), .ZN(n10005) );
  NAND2_X1 U10719 ( .A1(n10254), .A2(n10080), .ZN(n9774) );
  NAND2_X1 U10720 ( .A1(n10005), .A2(n9723), .ZN(n9770) );
  NAND2_X1 U10721 ( .A1(n9751), .A2(n9770), .ZN(n9724) );
  MUX2_X1 U10722 ( .A(n9724), .B(n9751), .S(n9747), .Z(n9725) );
  INV_X1 U10723 ( .A(n10059), .ZN(n10029) );
  NAND2_X1 U10724 ( .A1(n10248), .A2(n10029), .ZN(n10007) );
  MUX2_X1 U10725 ( .A(n10047), .B(n9774), .S(n9747), .Z(n9726) );
  NAND3_X1 U10726 ( .A1(n9727), .A2(n10049), .A3(n9726), .ZN(n9729) );
  MUX2_X1 U10727 ( .A(n9749), .B(n10007), .S(n9742), .Z(n9728) );
  AND2_X1 U10728 ( .A1(n9729), .A2(n9728), .ZN(n9741) );
  NAND2_X1 U10729 ( .A1(n5979), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9731) );
  INV_X1 U10730 ( .A(n10052), .ZN(n9733) );
  NAND2_X1 U10731 ( .A1(n10245), .A2(n9733), .ZN(n9779) );
  NAND2_X1 U10732 ( .A1(n9734), .A2(n6143), .ZN(n9736) );
  NAND2_X1 U10733 ( .A1(n5979), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9735) );
  INV_X1 U10734 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9995) );
  NAND2_X1 U10735 ( .A1(n6121), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9739) );
  INV_X1 U10736 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9737) );
  OR2_X1 U10737 ( .A1(n5954), .A2(n9737), .ZN(n9738) );
  OAI211_X1 U10738 ( .C1(n6645), .C2(n9995), .A(n9739), .B(n9738), .ZN(n10010)
         );
  INV_X1 U10739 ( .A(n10010), .ZN(n9790) );
  NOR2_X1 U10740 ( .A1(n9789), .A2(n9790), .ZN(n9880) );
  NAND2_X1 U10741 ( .A1(n9880), .A2(n9991), .ZN(n9784) );
  MUX2_X1 U10742 ( .A(n9750), .B(n9779), .S(n9742), .Z(n9740) );
  AOI21_X1 U10743 ( .B1(n9991), .B2(n10010), .A(n10242), .ZN(n9782) );
  AOI21_X1 U10744 ( .B1(n9782), .B2(n9747), .A(n9743), .ZN(n9744) );
  INV_X1 U10745 ( .A(n10239), .ZN(n9746) );
  INV_X1 U10746 ( .A(n9991), .ZN(n9745) );
  AOI21_X1 U10747 ( .B1(n9784), .B2(n9818), .A(n9747), .ZN(n9748) );
  AOI211_X1 U10748 ( .C1(n6328), .C2(n9743), .A(n9893), .B(n9829), .ZN(n9891)
         );
  NAND2_X1 U10749 ( .A1(n9750), .A2(n9749), .ZN(n9780) );
  AND2_X1 U10750 ( .A1(n10047), .A2(n9751), .ZN(n9778) );
  INV_X1 U10751 ( .A(n9778), .ZN(n9757) );
  NAND2_X1 U10752 ( .A1(n9752), .A2(n10003), .ZN(n9753) );
  NAND2_X1 U10753 ( .A1(n9753), .A2(n10004), .ZN(n9755) );
  NAND2_X1 U10754 ( .A1(n9755), .A2(n9754), .ZN(n9756) );
  NAND2_X1 U10755 ( .A1(n10076), .A2(n9756), .ZN(n9772) );
  INV_X1 U10756 ( .A(n9879), .ZN(n9783) );
  INV_X1 U10757 ( .A(n9759), .ZN(n9760) );
  INV_X1 U10758 ( .A(n9794), .ZN(n9870) );
  INV_X1 U10759 ( .A(n10192), .ZN(n9762) );
  NAND2_X1 U10760 ( .A1(n10194), .A2(n9763), .ZN(n10175) );
  INV_X1 U10761 ( .A(n9874), .ZN(n9764) );
  INV_X1 U10762 ( .A(n10156), .ZN(n9765) );
  NAND2_X1 U10763 ( .A1(n9874), .A2(n9765), .ZN(n9767) );
  NAND2_X1 U10764 ( .A1(n9767), .A2(n9766), .ZN(n9999) );
  NOR3_X1 U10765 ( .A1(n9769), .A2(n9768), .A3(n9999), .ZN(n9773) );
  INV_X1 U10766 ( .A(n9770), .ZN(n9771) );
  OAI21_X1 U10767 ( .B1(n9773), .B2(n9772), .A(n9771), .ZN(n9777) );
  INV_X1 U10768 ( .A(n9774), .ZN(n9776) );
  INV_X1 U10769 ( .A(n10007), .ZN(n9775) );
  AOI211_X1 U10770 ( .C1(n9778), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9781)
         );
  OAI21_X1 U10771 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9883) );
  AOI211_X1 U10772 ( .C1(n9783), .C2(n10000), .A(n9883), .B(n9782), .ZN(n9786)
         );
  OAI21_X1 U10773 ( .B1(n9786), .B2(n5255), .A(n9785), .ZN(n9788) );
  NAND3_X1 U10774 ( .A1(n9788), .A2(n9787), .A3(n9818), .ZN(n9820) );
  AOI21_X1 U10775 ( .B1(n9790), .B2(n9789), .A(n9743), .ZN(n9886) );
  INV_X1 U10776 ( .A(n10049), .ZN(n9817) );
  NOR2_X1 U10777 ( .A1(n9792), .A2(n9791), .ZN(n10002) );
  INV_X1 U10778 ( .A(n10002), .ZN(n10127) );
  NAND2_X1 U10779 ( .A1(n9794), .A2(n10192), .ZN(n10206) );
  INV_X1 U10780 ( .A(n9795), .ZN(n9807) );
  NAND4_X1 U10781 ( .A1(n9798), .A2(n9797), .A3(n9796), .A4(n9822), .ZN(n9801)
         );
  NOR4_X1 U10782 ( .A1(n9801), .A2(n9800), .A3(n9799), .A4(n10966), .ZN(n9804)
         );
  INV_X1 U10783 ( .A(n9802), .ZN(n9803) );
  NAND4_X1 U10784 ( .A1(n9804), .A2(n9849), .A3(n9803), .A4(n9851), .ZN(n9805)
         );
  NOR4_X1 U10785 ( .A1(n9807), .A2(n9806), .A3(n5683), .A4(n9805), .ZN(n9809)
         );
  NAND4_X1 U10786 ( .A1(n9811), .A2(n9810), .A3(n9809), .A4(n9808), .ZN(n9812)
         );
  NOR4_X1 U10787 ( .A1(n10206), .A2(n10226), .A3(n5328), .A4(n9812), .ZN(n9813) );
  NAND4_X1 U10788 ( .A1(n5705), .A2(n10191), .A3(n10176), .A4(n9813), .ZN(
        n9814) );
  NOR4_X1 U10789 ( .A1(n10127), .A2(n10114), .A3(n10021), .A4(n9814), .ZN(
        n9815) );
  NAND4_X1 U10790 ( .A1(n10057), .A2(n10075), .A3(n10088), .A4(n9815), .ZN(
        n9816) );
  NOR4_X1 U10791 ( .A1(n9880), .A2(n10031), .A3(n9817), .A4(n9816), .ZN(n9819)
         );
  NAND3_X1 U10792 ( .A1(n9886), .A2(n9819), .A3(n9818), .ZN(n9823) );
  AOI21_X1 U10793 ( .B1(n9820), .B2(n9823), .A(n6328), .ZN(n9821) );
  INV_X1 U10794 ( .A(n9821), .ZN(n9831) );
  NAND2_X1 U10795 ( .A1(n6328), .A2(n9822), .ZN(n9825) );
  INV_X1 U10796 ( .A(n9823), .ZN(n9824) );
  AOI21_X1 U10797 ( .B1(n9826), .B2(n9825), .A(n9824), .ZN(n9828) );
  NAND2_X1 U10798 ( .A1(n9831), .A2(n9830), .ZN(n9890) );
  INV_X1 U10799 ( .A(n9832), .ZN(n9872) );
  INV_X1 U10800 ( .A(n9833), .ZN(n9836) );
  NAND2_X1 U10801 ( .A1(n5886), .A2(n10880), .ZN(n9834) );
  NAND3_X1 U10802 ( .A1(n9836), .A2(n9835), .A3(n9834), .ZN(n9837) );
  NAND2_X1 U10803 ( .A1(n10909), .A2(n9837), .ZN(n9840) );
  INV_X1 U10804 ( .A(n9838), .ZN(n9839) );
  OAI21_X1 U10805 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n9845) );
  INV_X1 U10806 ( .A(n9842), .ZN(n9843) );
  AOI21_X1 U10807 ( .B1(n9845), .B2(n9844), .A(n9843), .ZN(n9848) );
  OAI21_X1 U10808 ( .B1(n9848), .B2(n9847), .A(n9846), .ZN(n9852) );
  INV_X1 U10809 ( .A(n9849), .ZN(n9850) );
  AOI21_X1 U10810 ( .B1(n9852), .B2(n9851), .A(n9850), .ZN(n9855) );
  OAI21_X1 U10811 ( .B1(n9855), .B2(n9854), .A(n9853), .ZN(n9859) );
  INV_X1 U10812 ( .A(n9856), .ZN(n9858) );
  AOI21_X1 U10813 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9862) );
  OAI211_X1 U10814 ( .C1(n9862), .C2(n9861), .A(n5330), .B(n9860), .ZN(n9866)
         );
  INV_X1 U10815 ( .A(n9863), .ZN(n9865) );
  NAND3_X1 U10816 ( .A1(n9866), .A2(n9865), .A3(n9864), .ZN(n9867) );
  NAND3_X1 U10817 ( .A1(n9869), .A2(n9868), .A3(n9867), .ZN(n9871) );
  AOI21_X1 U10818 ( .B1(n9872), .B2(n9871), .A(n9870), .ZN(n9876) );
  INV_X1 U10819 ( .A(n9873), .ZN(n9875) );
  OAI211_X1 U10820 ( .C1(n9877), .C2(n9876), .A(n9875), .B(n9874), .ZN(n9878)
         );
  NOR2_X1 U10821 ( .A1(n9879), .A2(n9878), .ZN(n9882) );
  INV_X1 U10822 ( .A(n9880), .ZN(n9881) );
  OAI21_X1 U10823 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9885) );
  AOI21_X1 U10824 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9887) );
  XNOR2_X1 U10825 ( .A(n9887), .B(n6328), .ZN(n9888) );
  NAND2_X1 U10826 ( .A1(n9888), .A2(n7908), .ZN(n9889) );
  NOR2_X1 U10827 ( .A1(n9892), .A2(n10826), .ZN(n9895) );
  OAI21_X1 U10828 ( .B1(n9896), .B2(n9893), .A(P1_B_REG_SCAN_IN), .ZN(n9894)
         );
  OAI22_X1 U10829 ( .A1(n9897), .A2(n9896), .B1(n9895), .B2(n9894), .ZN(
        P1_U3242) );
  MUX2_X1 U10830 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n10010), .S(n9910), .Z(
        P1_U3584) );
  MUX2_X1 U10831 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n10052), .S(n9910), .Z(
        P1_U3583) );
  MUX2_X1 U10832 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10059), .S(n9910), .Z(
        P1_U3582) );
  MUX2_X1 U10833 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10051), .S(n9910), .Z(
        P1_U3581) );
  MUX2_X1 U10834 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9898), .S(n9910), .Z(
        P1_U3579) );
  MUX2_X1 U10835 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10133), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10836 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10132), .S(n9910), .Z(
        P1_U3576) );
  MUX2_X1 U10837 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10148), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10838 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10197), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10839 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10017), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10840 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10223), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10841 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n10016), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10842 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10222), .S(n9910), .Z(
        P1_U3570) );
  MUX2_X1 U10843 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9899), .S(n9910), .Z(
        P1_U3569) );
  MUX2_X1 U10844 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9900), .S(n9910), .Z(
        P1_U3568) );
  MUX2_X1 U10845 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9901), .S(n9910), .Z(
        P1_U3567) );
  MUX2_X1 U10846 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9902), .S(n9910), .Z(
        P1_U3566) );
  MUX2_X1 U10847 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9903), .S(n9910), .Z(
        P1_U3565) );
  MUX2_X1 U10848 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9904), .S(n9910), .Z(
        P1_U3564) );
  MUX2_X1 U10849 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9905), .S(n9910), .Z(
        P1_U3563) );
  MUX2_X1 U10850 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9906), .S(n9910), .Z(
        P1_U3562) );
  MUX2_X1 U10851 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9907), .S(n9910), .Z(
        P1_U3561) );
  MUX2_X1 U10852 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n10970), .S(n9910), .Z(
        P1_U3560) );
  MUX2_X1 U10853 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9908), .S(n9910), .Z(
        P1_U3559) );
  MUX2_X1 U10854 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n10968), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10855 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9909), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10856 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n5839), .S(n9910), .Z(
        P1_U3556) );
  MUX2_X1 U10857 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5886), .S(n9910), .Z(
        P1_U3555) );
  MUX2_X1 U10858 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6953), .S(n9910), .Z(
        P1_U3554) );
  AND2_X1 U10859 ( .A1(n9912), .A2(n9911), .ZN(n9913) );
  AOI21_X1 U10860 ( .B1(n9914), .B2(P1_REG1_REG_15__SCAN_IN), .A(n9913), .ZN(
        n9916) );
  INV_X1 U10861 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9918) );
  MUX2_X1 U10862 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9918), .S(n9932), .Z(n9915) );
  NAND2_X1 U10863 ( .A1(n9916), .A2(n9915), .ZN(n9933) );
  INV_X1 U10864 ( .A(n9933), .ZN(n9941) );
  NOR2_X1 U10865 ( .A1(n9932), .A2(n9918), .ZN(n9917) );
  AOI211_X1 U10866 ( .C1(n9918), .C2(n9932), .A(n9917), .B(n9916), .ZN(n9919)
         );
  OAI21_X1 U10867 ( .B1(n9941), .B2(n9919), .A(n10871), .ZN(n9930) );
  INV_X1 U10868 ( .A(n9920), .ZN(n9928) );
  NAND2_X1 U10869 ( .A1(n9932), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9944) );
  OR2_X1 U10870 ( .A1(n9932), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U10871 ( .A1(n9944), .A2(n9923), .ZN(n9925) );
  INV_X1 U10872 ( .A(n9945), .ZN(n9924) );
  AOI211_X1 U10873 ( .C1(n9926), .C2(n9925), .A(n9924), .B(n10862), .ZN(n9927)
         );
  AOI211_X1 U10874 ( .C1(n10861), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9928), .B(
        n9927), .ZN(n9929) );
  OAI211_X1 U10875 ( .C1(n10849), .C2(n9931), .A(n9930), .B(n9929), .ZN(
        P1_U3259) );
  OR2_X1 U10876 ( .A1(n9932), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U10877 ( .A1(n9933), .A2(n9938), .ZN(n9937) );
  INV_X1 U10878 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9934) );
  OR2_X1 U10879 ( .A1(n9962), .A2(n9934), .ZN(n9936) );
  NAND2_X1 U10880 ( .A1(n9962), .A2(n9934), .ZN(n9935) );
  NAND2_X1 U10881 ( .A1(n9936), .A2(n9935), .ZN(n9939) );
  NAND2_X1 U10882 ( .A1(n9937), .A2(n9939), .ZN(n9957) );
  INV_X1 U10883 ( .A(n9957), .ZN(n9943) );
  INV_X1 U10884 ( .A(n9938), .ZN(n9940) );
  NOR3_X1 U10885 ( .A1(n9941), .A2(n9940), .A3(n9939), .ZN(n9942) );
  OAI21_X1 U10886 ( .B1(n9943), .B2(n9942), .A(n10871), .ZN(n9952) );
  NOR2_X1 U10887 ( .A1(n9953), .A2(n10229), .ZN(n9946) );
  AOI21_X1 U10888 ( .B1(n10229), .B2(n9953), .A(n9946), .ZN(n9947) );
  AOI221_X1 U10889 ( .B1(n9948), .B2(n9961), .C1(n9947), .C2(n9961), .A(n10862), .ZN(n9949) );
  AOI211_X1 U10890 ( .C1(n10861), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9950), .B(
        n9949), .ZN(n9951) );
  OAI211_X1 U10891 ( .C1(n10849), .C2(n9953), .A(n9952), .B(n9951), .ZN(
        P1_U3260) );
  INV_X1 U10892 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9954) );
  XNOR2_X1 U10893 ( .A(n9975), .B(n9954), .ZN(n9959) );
  OR2_X1 U10894 ( .A1(n9962), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9955) );
  AND2_X1 U10895 ( .A1(n9957), .A2(n9955), .ZN(n9958) );
  AND2_X1 U10896 ( .A1(n9959), .A2(n9955), .ZN(n9956) );
  NAND2_X1 U10897 ( .A1(n9957), .A2(n9956), .ZN(n9977) );
  OAI211_X1 U10898 ( .C1(n9959), .C2(n9958), .A(n10871), .B(n9977), .ZN(n9970)
         );
  INV_X1 U10899 ( .A(n9960), .ZN(n9968) );
  OAI21_X1 U10900 ( .B1(n9962), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9961), .ZN(
        n9966) );
  NOR2_X1 U10901 ( .A1(n9975), .A2(n9963), .ZN(n9964) );
  AOI21_X1 U10902 ( .B1(n9975), .B2(n9963), .A(n9964), .ZN(n9965) );
  AOI211_X1 U10903 ( .C1(n9966), .C2(n9965), .A(n9972), .B(n10862), .ZN(n9967)
         );
  AOI211_X1 U10904 ( .C1(n10861), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9968), .B(
        n9967), .ZN(n9969) );
  OAI211_X1 U10905 ( .C1(n10849), .C2(n9971), .A(n9970), .B(n9969), .ZN(
        P1_U3261) );
  AOI21_X1 U10906 ( .B1(n9975), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9972), .ZN(
        n9974) );
  MUX2_X1 U10907 ( .A(n6333), .B(P1_REG2_REG_19__SCAN_IN), .S(n10179), .Z(
        n9973) );
  XNOR2_X1 U10908 ( .A(n9974), .B(n9973), .ZN(n9985) );
  NAND2_X1 U10909 ( .A1(n9975), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U10910 ( .A1(n9977), .A2(n9976), .ZN(n9979) );
  XNOR2_X1 U10911 ( .A(n10179), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9978) );
  XNOR2_X1 U10912 ( .A(n9979), .B(n9978), .ZN(n9980) );
  NOR2_X1 U10913 ( .A1(n10851), .A2(n9980), .ZN(n9984) );
  NAND2_X1 U10914 ( .A1(n10861), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9981) );
  OAI211_X1 U10915 ( .C1(n10849), .C2(n10179), .A(n9982), .B(n9981), .ZN(n9983) );
  AOI211_X1 U10916 ( .C1(n9985), .C2(n10855), .A(n9984), .B(n9983), .ZN(n9986)
         );
  INV_X1 U10917 ( .A(n9986), .ZN(P1_U3262) );
  NAND2_X1 U10918 ( .A1(n10210), .A2(n10216), .ZN(n10211) );
  INV_X1 U10919 ( .A(n10284), .ZN(n10168) );
  INV_X1 U10920 ( .A(n10277), .ZN(n10143) );
  XNOR2_X1 U10921 ( .A(n10239), .B(n9987), .ZN(n9988) );
  NAND2_X1 U10922 ( .A1(n9988), .A2(n11006), .ZN(n10238) );
  NAND2_X1 U10923 ( .A1(n9989), .A2(P1_B_REG_SCAN_IN), .ZN(n9990) );
  AND2_X1 U10924 ( .A1(n10969), .A2(n9990), .ZN(n10009) );
  NAND2_X1 U10925 ( .A1(n9991), .A2(n10009), .ZN(n10240) );
  NOR2_X1 U10926 ( .A1(n10180), .A2(n10240), .ZN(n9996) );
  NOR2_X1 U10927 ( .A1(n10239), .A2(n11031), .ZN(n9992) );
  AOI211_X1 U10928 ( .C1(n11028), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9996), .B(
        n9992), .ZN(n9993) );
  OAI21_X1 U10929 ( .B1(n10238), .B2(n10231), .A(n9993), .ZN(P1_U3263) );
  XNOR2_X1 U10930 ( .A(n9789), .B(n10033), .ZN(n9994) );
  NAND2_X1 U10931 ( .A1(n9994), .A2(n11006), .ZN(n10241) );
  NOR2_X1 U10932 ( .A1(n10218), .A2(n9995), .ZN(n9997) );
  AOI211_X1 U10933 ( .C1(n9789), .C2(n10235), .A(n9997), .B(n9996), .ZN(n9998)
         );
  OAI21_X1 U10934 ( .B1(n10241), .B2(n10231), .A(n9998), .ZN(P1_U3264) );
  NAND3_X1 U10935 ( .A1(n10144), .A2(n10002), .A3(n10001), .ZN(n10130) );
  INV_X1 U10936 ( .A(n10005), .ZN(n10006) );
  NAND3_X1 U10937 ( .A1(n10056), .A2(n10049), .A3(n10047), .ZN(n10048) );
  NAND2_X1 U10938 ( .A1(n10048), .A2(n10007), .ZN(n10008) );
  AOI22_X1 U10939 ( .A1(n10967), .A2(n10059), .B1(n10010), .B2(n10009), .ZN(
        n10011) );
  NAND2_X1 U10940 ( .A1(n10203), .A2(n10206), .ZN(n10202) );
  NAND2_X1 U10941 ( .A1(n10293), .A2(n10017), .ZN(n10018) );
  INV_X1 U10942 ( .A(n10293), .ZN(n10190) );
  NAND2_X1 U10943 ( .A1(n10168), .A2(n10178), .ZN(n10019) );
  NOR2_X1 U10944 ( .A1(n10277), .A2(n10132), .ZN(n10020) );
  AOI21_X1 U10945 ( .B1(n10138), .B2(n10021), .A(n10020), .ZN(n10122) );
  NAND2_X1 U10946 ( .A1(n10126), .A2(n10116), .ZN(n10022) );
  NAND2_X1 U10947 ( .A1(n10122), .A2(n10022), .ZN(n10024) );
  NAND2_X1 U10948 ( .A1(n10273), .A2(n10147), .ZN(n10023) );
  NAND2_X1 U10949 ( .A1(n10024), .A2(n10023), .ZN(n10107) );
  NOR2_X1 U10950 ( .A1(n10111), .A2(n10097), .ZN(n10026) );
  NAND2_X1 U10951 ( .A1(n10111), .A2(n10097), .ZN(n10025) );
  OAI21_X2 U10952 ( .B1(n10107), .B2(n10026), .A(n10025), .ZN(n10089) );
  AOI21_X1 U10953 ( .B1(n10089), .B2(n10094), .A(n5762), .ZN(n10074) );
  NAND2_X1 U10954 ( .A1(n10259), .A2(n10060), .ZN(n10028) );
  NOR2_X1 U10955 ( .A1(n10248), .A2(n10059), .ZN(n10030) );
  INV_X1 U10956 ( .A(n10248), .ZN(n10046) );
  OAI22_X1 U10957 ( .A1(n10041), .A2(n10030), .B1(n10046), .B2(n10029), .ZN(
        n10032) );
  XNOR2_X1 U10958 ( .A(n10032), .B(n5269), .ZN(n10243) );
  NAND2_X1 U10959 ( .A1(n10243), .A2(n10982), .ZN(n10040) );
  AOI211_X1 U10960 ( .C1(n10245), .C2(n10042), .A(n11042), .B(n10033), .ZN(
        n10244) );
  INV_X1 U10961 ( .A(n10245), .ZN(n10034) );
  NOR2_X1 U10962 ( .A1(n10034), .A2(n11031), .ZN(n10038) );
  OAI22_X1 U10963 ( .A1(n10218), .A2(n10036), .B1(n10035), .B2(n10227), .ZN(
        n10037) );
  AOI211_X1 U10964 ( .C1(n10244), .C2(n11035), .A(n10038), .B(n10037), .ZN(
        n10039) );
  OAI211_X1 U10965 ( .C1(n5173), .C2(n10180), .A(n10040), .B(n10039), .ZN(
        P1_U3356) );
  XNOR2_X1 U10966 ( .A(n10041), .B(n10049), .ZN(n10251) );
  INV_X1 U10967 ( .A(n10042), .ZN(n10043) );
  AOI211_X1 U10968 ( .C1(n10248), .C2(n10063), .A(n11042), .B(n10043), .ZN(
        n10247) );
  AOI22_X1 U10969 ( .A1(n10180), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n10044), 
        .B2(n11026), .ZN(n10045) );
  OAI21_X1 U10970 ( .B1(n10046), .B2(n11031), .A(n10045), .ZN(n10054) );
  OAI21_X1 U10971 ( .B1(n10050), .B2(n10049), .A(n10048), .ZN(n10053) );
  OAI211_X1 U10972 ( .C1(n10058), .C2(n10057), .A(n10056), .B(n10972), .ZN(
        n10062) );
  AOI22_X1 U10973 ( .A1(n10967), .A2(n10060), .B1(n10059), .B2(n10969), .ZN(
        n10061) );
  NAND2_X1 U10974 ( .A1(n10062), .A2(n10061), .ZN(n10252) );
  INV_X1 U10975 ( .A(n10063), .ZN(n10064) );
  AOI211_X1 U10976 ( .C1(n10254), .C2(n10065), .A(n11042), .B(n10064), .ZN(
        n10253) );
  NAND2_X1 U10977 ( .A1(n10253), .A2(n11035), .ZN(n10068) );
  AOI22_X1 U10978 ( .A1(n11028), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10066), 
        .B2(n11026), .ZN(n10067) );
  OAI211_X1 U10979 ( .C1(n10069), .C2(n11031), .A(n10068), .B(n10067), .ZN(
        n10070) );
  AOI21_X1 U10980 ( .B1(n10252), .B2(n10218), .A(n10070), .ZN(n10071) );
  OAI21_X1 U10981 ( .B1(n10256), .B2(n10220), .A(n10071), .ZN(P1_U3266) );
  OAI21_X1 U10982 ( .B1(n10074), .B2(n10073), .A(n10072), .ZN(n10261) );
  AOI21_X1 U10983 ( .B1(n5337), .B2(n10076), .A(n10075), .ZN(n10077) );
  NOR2_X1 U10984 ( .A1(n10078), .A2(n10077), .ZN(n10079) );
  OAI222_X1 U10985 ( .A1(n11008), .A2(n10080), .B1(n11010), .B2(n10115), .C1(
        n11016), .C2(n10079), .ZN(n10257) );
  INV_X1 U10986 ( .A(n10259), .ZN(n10085) );
  AOI211_X1 U10987 ( .C1(n10259), .C2(n10100), .A(n11042), .B(n10081), .ZN(
        n10258) );
  NAND2_X1 U10988 ( .A1(n10258), .A2(n11035), .ZN(n10084) );
  AOI22_X1 U10989 ( .A1(n11028), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n10082), 
        .B2(n11026), .ZN(n10083) );
  OAI211_X1 U10990 ( .C1(n10085), .C2(n11031), .A(n10084), .B(n10083), .ZN(
        n10086) );
  AOI21_X1 U10991 ( .B1(n10257), .B2(n10218), .A(n10086), .ZN(n10087) );
  OAI21_X1 U10992 ( .B1(n10261), .B2(n10220), .A(n10087), .ZN(P1_U3267) );
  XNOR2_X1 U10993 ( .A(n10089), .B(n10088), .ZN(n10266) );
  INV_X1 U10994 ( .A(n10090), .ZN(n10091) );
  OAI22_X1 U10995 ( .A1(n10218), .A2(n10092), .B1(n10091), .B2(n10227), .ZN(
        n10105) );
  AOI211_X1 U10996 ( .C1(n10095), .C2(n10094), .A(n11016), .B(n10093), .ZN(
        n10099) );
  OAI22_X1 U10997 ( .A1(n10097), .A2(n11010), .B1(n10096), .B2(n11008), .ZN(
        n10098) );
  NOR2_X1 U10998 ( .A1(n10099), .A2(n10098), .ZN(n10265) );
  INV_X1 U10999 ( .A(n10100), .ZN(n10101) );
  AOI211_X1 U11000 ( .C1(n10263), .C2(n10102), .A(n11042), .B(n10101), .ZN(
        n10262) );
  NAND2_X1 U11001 ( .A1(n10262), .A2(n10179), .ZN(n10103) );
  AOI21_X1 U11002 ( .B1(n10265), .B2(n10103), .A(n10180), .ZN(n10104) );
  AOI211_X1 U11003 ( .C1(n10235), .C2(n10263), .A(n10105), .B(n10104), .ZN(
        n10106) );
  OAI21_X1 U11004 ( .B1(n10266), .B2(n10220), .A(n10106), .ZN(P1_U3268) );
  XNOR2_X1 U11005 ( .A(n10107), .B(n10114), .ZN(n10271) );
  AOI211_X1 U11006 ( .C1(n10268), .C2(n10123), .A(n11042), .B(n10108), .ZN(
        n10267) );
  AOI22_X1 U11007 ( .A1(n11028), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n10109), 
        .B2(n11026), .ZN(n10110) );
  OAI21_X1 U11008 ( .B1(n10111), .B2(n11031), .A(n10110), .ZN(n10120) );
  AOI211_X1 U11009 ( .C1(n10114), .C2(n10113), .A(n11016), .B(n10112), .ZN(
        n10118) );
  OAI22_X1 U11010 ( .A1(n10116), .A2(n11010), .B1(n10115), .B2(n11008), .ZN(
        n10117) );
  NOR2_X1 U11011 ( .A1(n10118), .A2(n10117), .ZN(n10270) );
  NOR2_X1 U11012 ( .A1(n10270), .A2(n10180), .ZN(n10119) );
  AOI211_X1 U11013 ( .C1(n10267), .C2(n11035), .A(n10120), .B(n10119), .ZN(
        n10121) );
  OAI21_X1 U11014 ( .B1(n10271), .B2(n10220), .A(n10121), .ZN(P1_U3269) );
  XNOR2_X1 U11015 ( .A(n10122), .B(n10127), .ZN(n10276) );
  AOI211_X1 U11016 ( .C1(n10273), .C2(n10139), .A(n11042), .B(n5350), .ZN(
        n10272) );
  AOI22_X1 U11017 ( .A1(n11028), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10124), 
        .B2(n11026), .ZN(n10125) );
  OAI21_X1 U11018 ( .B1(n10126), .B2(n11031), .A(n10125), .ZN(n10136) );
  INV_X1 U11019 ( .A(n10144), .ZN(n10129) );
  OAI21_X1 U11020 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(n10131) );
  NAND2_X1 U11021 ( .A1(n10131), .A2(n10130), .ZN(n10134) );
  AOI222_X1 U11022 ( .A1(n10972), .A2(n10134), .B1(n10133), .B2(n10969), .C1(
        n10132), .C2(n10967), .ZN(n10275) );
  NOR2_X1 U11023 ( .A1(n10275), .A2(n11028), .ZN(n10135) );
  AOI211_X1 U11024 ( .C1(n10272), .C2(n11035), .A(n10136), .B(n10135), .ZN(
        n10137) );
  OAI21_X1 U11025 ( .B1(n10276), .B2(n10220), .A(n10137), .ZN(P1_U3270) );
  XNOR2_X1 U11026 ( .A(n10138), .B(n10145), .ZN(n10281) );
  INV_X1 U11027 ( .A(n10163), .ZN(n10140) );
  AOI21_X1 U11028 ( .B1(n10277), .B2(n10140), .A(n5351), .ZN(n10278) );
  AOI22_X1 U11029 ( .A1(n11028), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10141), 
        .B2(n11026), .ZN(n10142) );
  OAI21_X1 U11030 ( .B1(n10143), .B2(n11031), .A(n10142), .ZN(n10152) );
  OAI211_X1 U11031 ( .C1(n10146), .C2(n10145), .A(n10144), .B(n10972), .ZN(
        n10150) );
  AOI22_X1 U11032 ( .A1(n10967), .A2(n10148), .B1(n10147), .B2(n10969), .ZN(
        n10149) );
  AND2_X1 U11033 ( .A1(n10150), .A2(n10149), .ZN(n10280) );
  NOR2_X1 U11034 ( .A1(n10280), .A2(n10180), .ZN(n10151) );
  AOI211_X1 U11035 ( .C1(n10278), .C2(n10153), .A(n10152), .B(n10151), .ZN(
        n10154) );
  OAI21_X1 U11036 ( .B1(n10281), .B2(n10220), .A(n10154), .ZN(P1_U3271) );
  XNOR2_X1 U11037 ( .A(n10155), .B(n5705), .ZN(n10286) );
  NAND2_X1 U11038 ( .A1(n10157), .A2(n10156), .ZN(n10159) );
  XNOR2_X1 U11039 ( .A(n10159), .B(n10158), .ZN(n10160) );
  OAI222_X1 U11040 ( .A1(n11008), .A2(n10162), .B1(n11010), .B2(n10161), .C1(
        n10160), .C2(n11016), .ZN(n10282) );
  INV_X1 U11041 ( .A(n10174), .ZN(n10164) );
  AOI211_X1 U11042 ( .C1(n10284), .C2(n10164), .A(n11042), .B(n10163), .ZN(
        n10283) );
  NAND2_X1 U11043 ( .A1(n10283), .A2(n11035), .ZN(n10167) );
  AOI22_X1 U11044 ( .A1(n11028), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10165), 
        .B2(n11026), .ZN(n10166) );
  OAI211_X1 U11045 ( .C1(n10168), .C2(n11031), .A(n10167), .B(n10166), .ZN(
        n10169) );
  AOI21_X1 U11046 ( .B1(n10282), .B2(n10218), .A(n10169), .ZN(n10170) );
  OAI21_X1 U11047 ( .B1(n10286), .B2(n10220), .A(n10170), .ZN(P1_U3272) );
  XOR2_X1 U11048 ( .A(n10176), .B(n10171), .Z(n10291) );
  OAI22_X1 U11049 ( .A1(n10218), .A2(n10173), .B1(n10172), .B2(n10227), .ZN(
        n10183) );
  AOI211_X1 U11050 ( .C1(n10289), .C2(n10186), .A(n11042), .B(n10174), .ZN(
        n10288) );
  XOR2_X1 U11051 ( .A(n10176), .B(n10175), .Z(n10177) );
  OAI222_X1 U11052 ( .A1(n11008), .A2(n10178), .B1(n11010), .B2(n10209), .C1(
        n10177), .C2(n11016), .ZN(n10287) );
  AOI21_X1 U11053 ( .B1(n10288), .B2(n10179), .A(n10287), .ZN(n10181) );
  NOR2_X1 U11054 ( .A1(n10181), .A2(n10180), .ZN(n10182) );
  AOI211_X1 U11055 ( .C1(n10235), .C2(n10289), .A(n10183), .B(n10182), .ZN(
        n10184) );
  OAI21_X1 U11056 ( .B1(n10291), .B2(n10220), .A(n10184), .ZN(P1_U3273) );
  XNOR2_X1 U11057 ( .A(n10185), .B(n10191), .ZN(n10296) );
  INV_X1 U11058 ( .A(n10186), .ZN(n10187) );
  AOI211_X1 U11059 ( .C1(n10293), .C2(n10211), .A(n11042), .B(n10187), .ZN(
        n10292) );
  AOI22_X1 U11060 ( .A1(n11028), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n11026), 
        .B2(n10188), .ZN(n10189) );
  OAI21_X1 U11061 ( .B1(n10190), .B2(n11031), .A(n10189), .ZN(n10200) );
  INV_X1 U11062 ( .A(n10191), .ZN(n10193) );
  NAND2_X1 U11063 ( .A1(n10193), .A2(n10192), .ZN(n10195) );
  OAI21_X1 U11064 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10198) );
  AOI222_X1 U11065 ( .A1(n10972), .A2(n10198), .B1(n10223), .B2(n10967), .C1(
        n10197), .C2(n10969), .ZN(n10295) );
  NOR2_X1 U11066 ( .A1(n10295), .A2(n11028), .ZN(n10199) );
  AOI211_X1 U11067 ( .C1(n10292), .C2(n11035), .A(n10200), .B(n10199), .ZN(
        n10201) );
  OAI21_X1 U11068 ( .B1(n10296), .B2(n10220), .A(n10201), .ZN(P1_U3274) );
  OAI21_X1 U11069 ( .B1(n10203), .B2(n10206), .A(n10202), .ZN(n10204) );
  INV_X1 U11070 ( .A(n10204), .ZN(n10301) );
  XOR2_X1 U11071 ( .A(n10206), .B(n10205), .Z(n10207) );
  OAI222_X1 U11072 ( .A1(n11008), .A2(n10209), .B1(n11010), .B2(n10208), .C1(
        n11016), .C2(n10207), .ZN(n10297) );
  INV_X1 U11073 ( .A(n10210), .ZN(n10230) );
  INV_X1 U11074 ( .A(n10211), .ZN(n10212) );
  AOI211_X1 U11075 ( .C1(n10299), .C2(n10230), .A(n11042), .B(n10212), .ZN(
        n10298) );
  NAND2_X1 U11076 ( .A1(n10298), .A2(n11035), .ZN(n10215) );
  AOI22_X1 U11077 ( .A1(n11028), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10213), 
        .B2(n11026), .ZN(n10214) );
  OAI211_X1 U11078 ( .C1(n10216), .C2(n11031), .A(n10215), .B(n10214), .ZN(
        n10217) );
  AOI21_X1 U11079 ( .B1(n10297), .B2(n10218), .A(n10217), .ZN(n10219) );
  OAI21_X1 U11080 ( .B1(n10301), .B2(n10220), .A(n10219), .ZN(P1_U3275) );
  XOR2_X1 U11081 ( .A(n10226), .B(n10221), .Z(n10224) );
  AOI222_X1 U11082 ( .A1(n10972), .A2(n10224), .B1(n10223), .B2(n10969), .C1(
        n10222), .C2(n10967), .ZN(n11140) );
  XOR2_X1 U11083 ( .A(n10225), .B(n10226), .Z(n11145) );
  NAND2_X1 U11084 ( .A1(n11145), .A2(n10982), .ZN(n10237) );
  OAI22_X1 U11085 ( .A1(n10218), .A2(n10229), .B1(n10228), .B2(n10227), .ZN(
        n10233) );
  OAI211_X1 U11086 ( .C1(n11142), .C2(n5181), .A(n10230), .B(n11006), .ZN(
        n11139) );
  NOR2_X1 U11087 ( .A1(n11139), .A2(n10231), .ZN(n10232) );
  AOI211_X1 U11088 ( .C1(n10235), .C2(n10234), .A(n10233), .B(n10232), .ZN(
        n10236) );
  OAI211_X1 U11089 ( .C1(n11028), .C2(n11140), .A(n10237), .B(n10236), .ZN(
        P1_U3276) );
  OAI211_X1 U11090 ( .C1(n10239), .C2(n11141), .A(n10238), .B(n10240), .ZN(
        n10314) );
  MUX2_X1 U11091 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10314), .S(n11147), .Z(
        P1_U3553) );
  OAI211_X1 U11092 ( .C1(n10242), .C2(n11141), .A(n10241), .B(n10240), .ZN(
        n10315) );
  MUX2_X1 U11093 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10315), .S(n11147), .Z(
        P1_U3552) );
  NAND2_X1 U11094 ( .A1(n10243), .A2(n11144), .ZN(n10246) );
  MUX2_X1 U11095 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10316), .S(n11147), .Z(
        P1_U3551) );
  AOI21_X1 U11096 ( .B1(n10308), .B2(n10248), .A(n10247), .ZN(n10249) );
  OAI211_X1 U11097 ( .C1(n10251), .C2(n10885), .A(n10250), .B(n10249), .ZN(
        n10317) );
  MUX2_X1 U11098 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10317), .S(n11147), .Z(
        P1_U3550) );
  AOI211_X1 U11099 ( .C1(n10308), .C2(n10254), .A(n10253), .B(n10252), .ZN(
        n10255) );
  OAI21_X1 U11100 ( .B1(n10256), .B2(n10885), .A(n10255), .ZN(n10318) );
  MUX2_X1 U11101 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10318), .S(n11147), .Z(
        P1_U3549) );
  AOI211_X1 U11102 ( .C1(n10308), .C2(n10259), .A(n10258), .B(n10257), .ZN(
        n10260) );
  OAI21_X1 U11103 ( .B1(n10261), .B2(n10885), .A(n10260), .ZN(n10319) );
  MUX2_X1 U11104 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10319), .S(n11147), .Z(
        P1_U3548) );
  AOI21_X1 U11105 ( .B1(n10308), .B2(n10263), .A(n10262), .ZN(n10264) );
  OAI211_X1 U11106 ( .C1(n10266), .C2(n10885), .A(n10265), .B(n10264), .ZN(
        n10320) );
  MUX2_X1 U11107 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10320), .S(n11147), .Z(
        P1_U3547) );
  AOI21_X1 U11108 ( .B1(n10308), .B2(n10268), .A(n10267), .ZN(n10269) );
  OAI211_X1 U11109 ( .C1(n10271), .C2(n10885), .A(n10270), .B(n10269), .ZN(
        n10321) );
  MUX2_X1 U11110 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10321), .S(n11147), .Z(
        P1_U3546) );
  AOI21_X1 U11111 ( .B1(n10308), .B2(n10273), .A(n10272), .ZN(n10274) );
  OAI211_X1 U11112 ( .C1(n10276), .C2(n10885), .A(n10275), .B(n10274), .ZN(
        n10322) );
  MUX2_X1 U11113 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10322), .S(n11147), .Z(
        P1_U3545) );
  AOI22_X1 U11114 ( .A1(n10278), .A2(n11006), .B1(n10308), .B2(n10277), .ZN(
        n10279) );
  OAI211_X1 U11115 ( .C1(n10281), .C2(n10885), .A(n10280), .B(n10279), .ZN(
        n10323) );
  MUX2_X1 U11116 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10323), .S(n11147), .Z(
        P1_U3544) );
  AOI211_X1 U11117 ( .C1(n10308), .C2(n10284), .A(n10283), .B(n10282), .ZN(
        n10285) );
  OAI21_X1 U11118 ( .B1(n10286), .B2(n10885), .A(n10285), .ZN(n10324) );
  MUX2_X1 U11119 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10324), .S(n11147), .Z(
        P1_U3543) );
  AOI211_X1 U11120 ( .C1(n10308), .C2(n10289), .A(n10288), .B(n10287), .ZN(
        n10290) );
  OAI21_X1 U11121 ( .B1(n10291), .B2(n10885), .A(n10290), .ZN(n10325) );
  MUX2_X1 U11122 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10325), .S(n11147), .Z(
        P1_U3542) );
  AOI21_X1 U11123 ( .B1(n10308), .B2(n10293), .A(n10292), .ZN(n10294) );
  OAI211_X1 U11124 ( .C1(n10296), .C2(n10885), .A(n10295), .B(n10294), .ZN(
        n10326) );
  MUX2_X1 U11125 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10326), .S(n11147), .Z(
        P1_U3541) );
  AOI211_X1 U11126 ( .C1(n10308), .C2(n10299), .A(n10298), .B(n10297), .ZN(
        n10300) );
  OAI21_X1 U11127 ( .B1(n10301), .B2(n10885), .A(n10300), .ZN(n10327) );
  MUX2_X1 U11128 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10327), .S(n11147), .Z(
        P1_U3540) );
  AOI21_X1 U11129 ( .B1(n10308), .B2(n10303), .A(n10302), .ZN(n10304) );
  OAI211_X1 U11130 ( .C1(n10306), .C2(n10885), .A(n10305), .B(n10304), .ZN(
        n10328) );
  MUX2_X1 U11131 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10328), .S(n11147), .Z(
        P1_U3538) );
  AOI22_X1 U11132 ( .A1(n10309), .A2(n11006), .B1(n10308), .B2(n10307), .ZN(
        n10310) );
  OAI211_X1 U11133 ( .C1(n10312), .C2(n10877), .A(n10311), .B(n10310), .ZN(
        n10329) );
  MUX2_X1 U11134 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10329), .S(n11147), .Z(
        P1_U3536) );
  MUX2_X1 U11135 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10313), .S(n11147), .Z(
        P1_U3522) );
  MUX2_X1 U11136 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10314), .S(n11150), .Z(
        P1_U3521) );
  MUX2_X1 U11137 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10315), .S(n11150), .Z(
        P1_U3520) );
  MUX2_X1 U11138 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10316), .S(n11150), .Z(
        P1_U3519) );
  MUX2_X1 U11139 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10317), .S(n11150), .Z(
        P1_U3518) );
  MUX2_X1 U11140 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10318), .S(n11150), .Z(
        P1_U3517) );
  MUX2_X1 U11141 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10319), .S(n11150), .Z(
        P1_U3516) );
  MUX2_X1 U11142 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10320), .S(n11150), .Z(
        P1_U3515) );
  MUX2_X1 U11143 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10321), .S(n11150), .Z(
        P1_U3514) );
  MUX2_X1 U11144 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10322), .S(n11150), .Z(
        P1_U3513) );
  MUX2_X1 U11145 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10323), .S(n11150), .Z(
        P1_U3512) );
  MUX2_X1 U11146 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10324), .S(n11150), .Z(
        P1_U3511) );
  MUX2_X1 U11147 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10325), .S(n11150), .Z(
        P1_U3510) );
  MUX2_X1 U11148 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10326), .S(n11150), .Z(
        P1_U3509) );
  MUX2_X1 U11149 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10327), .S(n11150), .Z(
        P1_U3507) );
  MUX2_X1 U11150 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10328), .S(n11150), .Z(
        P1_U3501) );
  MUX2_X1 U11151 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10329), .S(n11150), .Z(
        P1_U3495) );
  NOR4_X1 U11152 ( .A1(n5776), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n5789), .ZN(n10330) );
  AOI21_X1 U11153 ( .B1(n10331), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10330), 
        .ZN(n10332) );
  OAI21_X1 U11154 ( .B1(n10333), .B2(n10340), .A(n10332), .ZN(P1_U3324) );
  INV_X1 U11155 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10675) );
  OAI222_X1 U11156 ( .A1(n10337), .A2(n10675), .B1(n10340), .B2(n10335), .C1(
        P1_U3086), .C2(n10334), .ZN(P1_U3325) );
  INV_X1 U11157 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10681) );
  OAI222_X1 U11158 ( .A1(n10340), .A2(n10336), .B1(n5780), .B2(P1_U3086), .C1(
        n10681), .C2(n10337), .ZN(P1_U3326) );
  OAI222_X1 U11159 ( .A1(n10340), .A2(n10339), .B1(n10338), .B2(P1_U3086), 
        .C1(n10373), .C2(n10337), .ZN(P1_U3327) );
  MUX2_X1 U11160 ( .A(n10341), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11161 ( .A(n10343), .ZN(n10342) );
  INV_X1 U11162 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10761) );
  NOR2_X1 U11163 ( .A1(n10342), .A2(n10761), .ZN(P1_U3323) );
  INV_X1 U11164 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10545) );
  NOR2_X1 U11165 ( .A1(n10342), .A2(n10545), .ZN(P1_U3322) );
  INV_X1 U11166 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10758) );
  NOR2_X1 U11167 ( .A1(n10342), .A2(n10758), .ZN(P1_U3321) );
  INV_X1 U11168 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10759) );
  NOR2_X1 U11169 ( .A1(n10342), .A2(n10759), .ZN(P1_U3320) );
  AND2_X1 U11170 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10343), .ZN(P1_U3319) );
  AND2_X1 U11171 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10343), .ZN(P1_U3318) );
  AND2_X1 U11172 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10343), .ZN(P1_U3317) );
  AND2_X1 U11173 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10343), .ZN(P1_U3316) );
  AND2_X1 U11174 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10343), .ZN(P1_U3315) );
  AND2_X1 U11175 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10343), .ZN(P1_U3314) );
  AND2_X1 U11176 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10343), .ZN(P1_U3313) );
  AND2_X1 U11177 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10343), .ZN(P1_U3312) );
  AND2_X1 U11178 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10343), .ZN(P1_U3311) );
  AND2_X1 U11179 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10343), .ZN(P1_U3310) );
  AND2_X1 U11180 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10343), .ZN(P1_U3309) );
  AND2_X1 U11181 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10343), .ZN(P1_U3308) );
  AND2_X1 U11182 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10343), .ZN(P1_U3307) );
  AND2_X1 U11183 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10343), .ZN(P1_U3306) );
  AND2_X1 U11184 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10343), .ZN(P1_U3305) );
  AND2_X1 U11185 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10343), .ZN(P1_U3304) );
  AND2_X1 U11186 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10343), .ZN(P1_U3303) );
  AND2_X1 U11187 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10343), .ZN(P1_U3302) );
  AND2_X1 U11188 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10343), .ZN(P1_U3301) );
  AND2_X1 U11189 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10343), .ZN(P1_U3300) );
  AND2_X1 U11190 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10343), .ZN(P1_U3299) );
  AND2_X1 U11191 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10343), .ZN(P1_U3298) );
  AND2_X1 U11192 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10343), .ZN(P1_U3297) );
  AND2_X1 U11193 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10343), .ZN(P1_U3296) );
  AND2_X1 U11194 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10343), .ZN(P1_U3295) );
  AND2_X1 U11195 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10343), .ZN(P1_U3294) );
  XOR2_X1 U11196 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10344), .Z(n10349) );
  XOR2_X1 U11197 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10345), .Z(n10347) );
  OAI22_X1 U11198 ( .A1(n10349), .A2(n10348), .B1(n10347), .B2(n10346), .ZN(
        n10359) );
  XNOR2_X1 U11199 ( .A(n10351), .B(n10350), .ZN(n10353) );
  NAND2_X1 U11200 ( .A1(n10353), .A2(n10352), .ZN(n10355) );
  OAI211_X1 U11201 ( .C1(n10357), .C2(n10356), .A(n10355), .B(n10354), .ZN(
        n10358) );
  AOI211_X1 U11202 ( .C1(n10360), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10359), .B(
        n10358), .ZN(n10766) );
  OAI22_X1 U11203 ( .A1(n10362), .A2(keyinput_123), .B1(keyinput_122), .B2(
        P1_D_REG_0__SCAN_IN), .ZN(n10361) );
  AOI221_X1 U11204 ( .B1(n10362), .B2(keyinput_123), .C1(P1_D_REG_0__SCAN_IN), 
        .C2(keyinput_122), .A(n10361), .ZN(n10550) );
  XOR2_X1 U11205 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .Z(n10364) );
  XNOR2_X1 U11206 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_106), .ZN(n10363)
         );
  OAI211_X1 U11207 ( .C1(P1_IR_REG_14__SCAN_IN), .C2(keyinput_104), .A(n10364), 
        .B(n10363), .ZN(n10368) );
  XNOR2_X1 U11208 ( .A(n10365), .B(keyinput_105), .ZN(n10367) );
  XNOR2_X1 U11209 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_102), .ZN(n10366)
         );
  OR3_X1 U11210 ( .A1(n10368), .A2(n10367), .A3(n10366), .ZN(n10369) );
  AOI21_X1 U11211 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_104), .A(n10369), 
        .ZN(n10526) );
  INV_X1 U11212 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10719) );
  INV_X1 U11213 ( .A(keyinput_101), .ZN(n10522) );
  OAI22_X1 U11214 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_91), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput_90), .ZN(n10370) );
  AOI221_X1 U11215 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_91), .C1(
        keyinput_90), .C2(P1_IR_REG_0__SCAN_IN), .A(n10370), .ZN(n10512) );
  OAI22_X1 U11216 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_87), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_88), .ZN(n10371) );
  AOI221_X1 U11217 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_87), .C1(
        keyinput_88), .C2(P2_DATAO_REG_8__SCAN_IN), .A(n10371), .ZN(n10505) );
  INV_X1 U11218 ( .A(keyinput_77), .ZN(n10491) );
  INV_X1 U11219 ( .A(keyinput_73), .ZN(n10482) );
  INV_X1 U11220 ( .A(keyinput_72), .ZN(n10481) );
  INV_X1 U11221 ( .A(keyinput_71), .ZN(n10480) );
  AOI22_X1 U11222 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_69), .B1(
        n10373), .B2(keyinput_68), .ZN(n10372) );
  OAI221_X1 U11223 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_69), .C1(
        n10373), .C2(keyinput_68), .A(n10372), .ZN(n10478) );
  INV_X1 U11224 ( .A(keyinput_67), .ZN(n10476) );
  OAI22_X1 U11225 ( .A1(n10673), .A2(keyinput_63), .B1(keyinput_64), .B2(
        P2_B_REG_SCAN_IN), .ZN(n10374) );
  AOI221_X1 U11226 ( .B1(n10673), .B2(keyinput_63), .C1(P2_B_REG_SCAN_IN), 
        .C2(keyinput_64), .A(n10374), .ZN(n10474) );
  INV_X1 U11227 ( .A(keyinput_51), .ZN(n10453) );
  INV_X1 U11228 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10660) );
  INV_X1 U11229 ( .A(keyinput_50), .ZN(n10452) );
  INV_X1 U11230 ( .A(keyinput_49), .ZN(n10451) );
  INV_X1 U11231 ( .A(keyinput_48), .ZN(n10450) );
  INV_X1 U11232 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U11233 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_45), .B1(n10376), .B2(keyinput_46), .ZN(n10375) );
  OAI221_X1 U11234 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(
        n10376), .C2(keyinput_46), .A(n10375), .ZN(n10447) );
  INV_X1 U11235 ( .A(keyinput_44), .ZN(n10445) );
  XNOR2_X1 U11236 ( .A(n10640), .B(keyinput_39), .ZN(n10443) );
  OAI22_X1 U11237 ( .A1(n10619), .A2(keyinput_23), .B1(n10618), .B2(
        keyinput_24), .ZN(n10377) );
  AOI221_X1 U11238 ( .B1(n10619), .B2(keyinput_23), .C1(keyinput_24), .C2(
        n10618), .A(n10377), .ZN(n10420) );
  INV_X1 U11239 ( .A(keyinput_19), .ZN(n10412) );
  INV_X1 U11240 ( .A(SI_13_), .ZN(n10613) );
  AOI22_X1 U11241 ( .A1(SI_16_), .A2(keyinput_16), .B1(n10379), .B2(
        keyinput_17), .ZN(n10378) );
  OAI221_X1 U11242 ( .B1(SI_16_), .B2(keyinput_16), .C1(n10379), .C2(
        keyinput_17), .A(n10378), .ZN(n10410) );
  INV_X1 U11243 ( .A(keyinput_2), .ZN(n10384) );
  INV_X1 U11244 ( .A(keyinput_3), .ZN(n10383) );
  INV_X1 U11245 ( .A(SI_30_), .ZN(n10380) );
  OAI22_X1 U11246 ( .A1(n10380), .A2(keyinput_2), .B1(keyinput_3), .B2(SI_29_), 
        .ZN(n10381) );
  INV_X1 U11247 ( .A(n10381), .ZN(n10382) );
  INV_X1 U11248 ( .A(n10385), .ZN(n10390) );
  AOI22_X1 U11249 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n10386) );
  OAI221_X1 U11250 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n10386), .ZN(n10389) );
  INV_X1 U11251 ( .A(SI_28_), .ZN(n10591) );
  AOI22_X1 U11252 ( .A1(SI_27_), .A2(keyinput_5), .B1(n10591), .B2(keyinput_4), 
        .ZN(n10387) );
  OAI221_X1 U11253 ( .B1(SI_27_), .B2(keyinput_5), .C1(n10591), .C2(keyinput_4), .A(n10387), .ZN(n10388) );
  AOI21_X1 U11254 ( .B1(n10390), .B2(n10389), .A(n10388), .ZN(n10398) );
  INV_X1 U11255 ( .A(keyinput_6), .ZN(n10391) );
  NAND2_X1 U11256 ( .A1(n10393), .A2(n10392), .ZN(n10397) );
  INV_X1 U11257 ( .A(SI_25_), .ZN(n10586) );
  AOI22_X1 U11258 ( .A1(n10585), .A2(keyinput_8), .B1(n10586), .B2(keyinput_7), 
        .ZN(n10394) );
  OAI221_X1 U11259 ( .B1(n10585), .B2(keyinput_8), .C1(n10586), .C2(keyinput_7), .A(n10394), .ZN(n10395) );
  OAI22_X1 U11260 ( .A1(n10599), .A2(keyinput_9), .B1(keyinput_11), .B2(SI_21_), .ZN(n10399) );
  AOI221_X1 U11261 ( .B1(n10599), .B2(keyinput_9), .C1(SI_21_), .C2(
        keyinput_11), .A(n10399), .ZN(n10402) );
  OAI22_X1 U11262 ( .A1(SI_22_), .A2(keyinput_10), .B1(keyinput_12), .B2(
        SI_20_), .ZN(n10400) );
  AOI221_X1 U11263 ( .B1(SI_22_), .B2(keyinput_10), .C1(SI_20_), .C2(
        keyinput_12), .A(n10400), .ZN(n10401) );
  OAI22_X1 U11264 ( .A1(SI_19_), .A2(keyinput_13), .B1(SI_18_), .B2(
        keyinput_14), .ZN(n10405) );
  AOI221_X1 U11265 ( .B1(SI_19_), .B2(keyinput_13), .C1(keyinput_14), .C2(
        SI_18_), .A(n10405), .ZN(n10407) );
  NOR2_X1 U11266 ( .A1(n10606), .A2(keyinput_15), .ZN(n10406) );
  AOI221_X1 U11267 ( .B1(n10408), .B2(n10407), .C1(keyinput_15), .C2(n10606), 
        .A(n10406), .ZN(n10409) );
  OAI22_X1 U11268 ( .A1(n10410), .A2(n10409), .B1(keyinput_18), .B2(SI_14_), 
        .ZN(n10411) );
  AOI22_X1 U11269 ( .A1(SI_12_), .A2(keyinput_20), .B1(n10414), .B2(
        keyinput_22), .ZN(n10413) );
  OAI221_X1 U11270 ( .B1(SI_12_), .B2(keyinput_20), .C1(n10414), .C2(
        keyinput_22), .A(n10413), .ZN(n10415) );
  XOR2_X1 U11271 ( .A(SI_5_), .B(keyinput_27), .Z(n10418) );
  INV_X1 U11272 ( .A(SI_7_), .ZN(n10620) );
  AOI22_X1 U11273 ( .A1(SI_6_), .A2(keyinput_26), .B1(n10620), .B2(keyinput_25), .ZN(n10416) );
  OAI221_X1 U11274 ( .B1(SI_6_), .B2(keyinput_26), .C1(n10620), .C2(
        keyinput_25), .A(n10416), .ZN(n10417) );
  AOI211_X1 U11275 ( .C1(n10420), .C2(n10419), .A(n10418), .B(n10417), .ZN(
        n10436) );
  XOR2_X1 U11276 ( .A(SI_4_), .B(keyinput_28), .Z(n10435) );
  INV_X1 U11277 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10422) );
  OAI22_X1 U11278 ( .A1(n10422), .A2(keyinput_38), .B1(n10626), .B2(
        keyinput_37), .ZN(n10421) );
  AOI221_X1 U11279 ( .B1(n10422), .B2(keyinput_38), .C1(keyinput_37), .C2(
        n10626), .A(n10421), .ZN(n10434) );
  AOI22_X1 U11280 ( .A1(SI_0_), .A2(keyinput_32), .B1(n5228), .B2(keyinput_33), 
        .ZN(n10423) );
  OAI221_X1 U11281 ( .B1(SI_0_), .B2(keyinput_32), .C1(n5228), .C2(keyinput_33), .A(n10423), .ZN(n10432) );
  AOI22_X1 U11282 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_35), .B1(n10425), 
        .B2(keyinput_36), .ZN(n10424) );
  OAI221_X1 U11283 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .C1(n10425), .C2(keyinput_36), .A(n10424), .ZN(n10431) );
  XNOR2_X1 U11284 ( .A(SI_1_), .B(keyinput_31), .ZN(n10429) );
  XNOR2_X1 U11285 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_34), .ZN(n10428) );
  XNOR2_X1 U11286 ( .A(SI_2_), .B(keyinput_30), .ZN(n10427) );
  XNOR2_X1 U11287 ( .A(SI_3_), .B(keyinput_29), .ZN(n10426) );
  NAND4_X1 U11288 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10430) );
  NOR3_X1 U11289 ( .A1(n10432), .A2(n10431), .A3(n10430), .ZN(n10433) );
  OAI211_X1 U11290 ( .C1(n10436), .C2(n10435), .A(n10434), .B(n10433), .ZN(
        n10442) );
  INV_X1 U11291 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U11292 ( .A1(n7021), .A2(keyinput_43), .B1(n10438), .B2(keyinput_41), .ZN(n10437) );
  OAI221_X1 U11293 ( .B1(n7021), .B2(keyinput_43), .C1(n10438), .C2(
        keyinput_41), .A(n10437), .ZN(n10441) );
  AOI22_X1 U11294 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_40), .B1(n7262), 
        .B2(keyinput_42), .ZN(n10439) );
  OAI221_X1 U11295 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(n7262), 
        .C2(keyinput_42), .A(n10439), .ZN(n10440) );
  AOI211_X1 U11296 ( .C1(n10443), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        n10444) );
  AOI221_X1 U11297 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n10445), .C1(n10649), 
        .C2(keyinput_44), .A(n10444), .ZN(n10446) );
  OAI22_X1 U11298 ( .A1(n10447), .A2(n10446), .B1(keyinput_47), .B2(
        P2_REG3_REG_25__SCAN_IN), .ZN(n10448) );
  AOI21_X1 U11299 ( .B1(keyinput_47), .B2(P2_REG3_REG_25__SCAN_IN), .A(n10448), 
        .ZN(n10449) );
  AOI22_X1 U11300 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_53), .B1(n10577), 
        .B2(keyinput_57), .ZN(n10454) );
  OAI221_X1 U11301 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .C1(n10577), .C2(keyinput_57), .A(n10454), .ZN(n10462) );
  AOI22_X1 U11302 ( .A1(n10456), .A2(keyinput_54), .B1(n10576), .B2(
        keyinput_56), .ZN(n10455) );
  OAI221_X1 U11303 ( .B1(n10456), .B2(keyinput_54), .C1(n10576), .C2(
        keyinput_56), .A(n10455), .ZN(n10461) );
  INV_X1 U11304 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10459) );
  INV_X1 U11305 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U11306 ( .A1(n10459), .A2(keyinput_55), .B1(keyinput_52), .B2(
        n10458), .ZN(n10457) );
  OAI221_X1 U11307 ( .B1(n10459), .B2(keyinput_55), .C1(n10458), .C2(
        keyinput_52), .A(n10457), .ZN(n10460) );
  AOI22_X1 U11308 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(n10572), 
        .B2(keyinput_58), .ZN(n10464) );
  OAI221_X1 U11309 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(n10572), .C2(keyinput_58), .A(n10464), .ZN(n10468) );
  OAI22_X1 U11310 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_62), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .ZN(n10465) );
  AOI221_X1 U11311 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_62), .C1(
        keyinput_60), .C2(P2_REG3_REG_18__SCAN_IN), .A(n10465), .ZN(n10467) );
  XNOR2_X1 U11312 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n10466)
         );
  OAI211_X1 U11313 ( .C1(n10469), .C2(n10468), .A(n10467), .B(n10466), .ZN(
        n10473) );
  INV_X1 U11314 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U11315 ( .A1(n10675), .A2(keyinput_66), .B1(keyinput_65), .B2(
        n10471), .ZN(n10470) );
  OAI221_X1 U11316 ( .B1(n10675), .B2(keyinput_66), .C1(n10471), .C2(
        keyinput_65), .A(n10470), .ZN(n10472) );
  AOI21_X1 U11317 ( .B1(n10474), .B2(n10473), .A(n10472), .ZN(n10475) );
  AOI221_X1 U11318 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_67), .C1(
        n10681), .C2(n10476), .A(n10475), .ZN(n10477) );
  OAI22_X1 U11319 ( .A1(keyinput_70), .A2(n10685), .B1(n10478), .B2(n10477), 
        .ZN(n10479) );
  AOI22_X1 U11320 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput_76), .B1(
        n10568), .B2(keyinput_74), .ZN(n10483) );
  OAI221_X1 U11321 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_76), .C1(
        n10568), .C2(keyinput_74), .A(n10483), .ZN(n10484) );
  INV_X1 U11322 ( .A(n10484), .ZN(n10487) );
  OAI221_X1 U11323 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(n10491), .C1(n10695), 
        .C2(keyinput_77), .A(n10490), .ZN(n10503) );
  AOI22_X1 U11324 ( .A1(n10557), .A2(keyinput_82), .B1(n10562), .B2(
        keyinput_78), .ZN(n10492) );
  OAI221_X1 U11325 ( .B1(n10557), .B2(keyinput_82), .C1(n10562), .C2(
        keyinput_78), .A(n10492), .ZN(n10499) );
  AOI22_X1 U11326 ( .A1(n10555), .A2(keyinput_79), .B1(keyinput_81), .B2(
        n10554), .ZN(n10493) );
  OAI221_X1 U11327 ( .B1(n10555), .B2(keyinput_79), .C1(n10554), .C2(
        keyinput_81), .A(n10493), .ZN(n10498) );
  AOI22_X1 U11328 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_85), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_83), .ZN(n10494) );
  OAI221_X1 U11329 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_85), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_83), .A(n10494), .ZN(n10497)
         );
  AOI22_X1 U11330 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_84), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_80), .ZN(n10495) );
  OAI221_X1 U11331 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_84), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_80), .A(n10495), .ZN(n10496)
         );
  NOR4_X1 U11332 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10502) );
  AOI22_X1 U11333 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(keyinput_93), .B1(n10508), 
        .B2(keyinput_92), .ZN(n10507) );
  OAI221_X1 U11334 ( .B1(P1_IR_REG_3__SCAN_IN), .B2(keyinput_93), .C1(n10508), 
        .C2(keyinput_92), .A(n10507), .ZN(n10511) );
  AOI22_X1 U11335 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_94), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_95), .ZN(n10509) );
  OAI221_X1 U11336 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_94), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_95), .A(n10509), .ZN(n10510) );
  INV_X1 U11337 ( .A(keyinput_96), .ZN(n10513) );
  MUX2_X1 U11338 ( .A(keyinput_96), .B(n10513), .S(P1_IR_REG_6__SCAN_IN), .Z(
        n10514) );
  NOR2_X1 U11339 ( .A1(n10515), .A2(n10514), .ZN(n10521) );
  AOI22_X1 U11340 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_98), .B1(n10517), 
        .B2(keyinput_97), .ZN(n10516) );
  OAI221_X1 U11341 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_98), .C1(n10517), 
        .C2(keyinput_97), .A(n10516), .ZN(n10520) );
  OAI22_X1 U11342 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_100), .B1(
        keyinput_99), .B2(P1_IR_REG_9__SCAN_IN), .ZN(n10518) );
  AOI221_X1 U11343 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_100), .C1(
        P1_IR_REG_9__SCAN_IN), .C2(keyinput_99), .A(n10518), .ZN(n10519) );
  XNOR2_X1 U11344 ( .A(n10729), .B(keyinput_107), .ZN(n10525) );
  AOI22_X1 U11345 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_109), .B1(n10730), 
        .B2(keyinput_108), .ZN(n10523) );
  OAI221_X1 U11346 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_109), .C1(n10730), .C2(keyinput_108), .A(n10523), .ZN(n10524) );
  AOI22_X1 U11347 ( .A1(n10735), .A2(keyinput_110), .B1(n5366), .B2(
        keyinput_113), .ZN(n10527) );
  OAI221_X1 U11348 ( .B1(n10735), .B2(keyinput_110), .C1(n5366), .C2(
        keyinput_113), .A(n10527), .ZN(n10532) );
  XOR2_X1 U11349 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_114), .Z(n10530) );
  XNOR2_X1 U11350 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_112), .ZN(n10529)
         );
  XNOR2_X1 U11351 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_111), .ZN(n10528)
         );
  NAND3_X1 U11352 ( .A1(n10530), .A2(n10529), .A3(n10528), .ZN(n10531) );
  XNOR2_X1 U11353 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_115), .ZN(n10535)
         );
  INV_X1 U11354 ( .A(keyinput_116), .ZN(n10533) );
  MUX2_X1 U11355 ( .A(keyinput_116), .B(n10533), .S(P1_IR_REG_26__SCAN_IN), 
        .Z(n10534) );
  AOI21_X1 U11356 ( .B1(n10536), .B2(n10535), .A(n10534), .ZN(n10539) );
  XOR2_X1 U11357 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_117), .Z(n10538) );
  XOR2_X1 U11358 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_118), .Z(n10537) );
  XNOR2_X1 U11359 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_119), .ZN(n10542)
         );
  XOR2_X1 U11360 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_120), .Z(n10541) );
  XNOR2_X1 U11361 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_121), .ZN(n10540)
         );
  OAI211_X1 U11362 ( .C1(n10543), .C2(n10542), .A(n10541), .B(n10540), .ZN(
        n10549) );
  AOI22_X1 U11363 ( .A1(n10545), .A2(keyinput_125), .B1(n10761), .B2(
        keyinput_124), .ZN(n10544) );
  OAI221_X1 U11364 ( .B1(n10545), .B2(keyinput_125), .C1(n10761), .C2(
        keyinput_124), .A(n10544), .ZN(n10548) );
  AOI22_X1 U11365 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput_127), .B1(n10758), 
        .B2(keyinput_126), .ZN(n10546) );
  OAI221_X1 U11366 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput_127), .C1(n10758), 
        .C2(keyinput_126), .A(n10546), .ZN(n10547) );
  AOI211_X1 U11367 ( .C1(n10550), .C2(n10549), .A(n10548), .B(n10547), .ZN(
        n10764) );
  INV_X1 U11368 ( .A(keyinput_229), .ZN(n10720) );
  AOI22_X1 U11369 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_216), .B1(
        n10552), .B2(keyinput_215), .ZN(n10551) );
  OAI221_X1 U11370 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_216), .C1(
        n10552), .C2(keyinput_215), .A(n10551), .ZN(n10698) );
  OAI22_X1 U11371 ( .A1(n10555), .A2(keyinput_207), .B1(n10554), .B2(
        keyinput_209), .ZN(n10553) );
  AOI221_X1 U11372 ( .B1(n10555), .B2(keyinput_207), .C1(keyinput_209), .C2(
        n10554), .A(n10553), .ZN(n10566) );
  OAI22_X1 U11373 ( .A1(n10558), .A2(keyinput_208), .B1(n10557), .B2(
        keyinput_210), .ZN(n10556) );
  AOI221_X1 U11374 ( .B1(n10558), .B2(keyinput_208), .C1(keyinput_210), .C2(
        n10557), .A(n10556), .ZN(n10565) );
  OAI22_X1 U11375 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_212), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_213), .ZN(n10559) );
  AOI221_X1 U11376 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_212), .C1(
        keyinput_213), .C2(P2_DATAO_REG_11__SCAN_IN), .A(n10559), .ZN(n10564)
         );
  OAI22_X1 U11377 ( .A1(n10562), .A2(keyinput_206), .B1(n10561), .B2(
        keyinput_211), .ZN(n10560) );
  AOI221_X1 U11378 ( .B1(n10562), .B2(keyinput_206), .C1(keyinput_211), .C2(
        n10561), .A(n10560), .ZN(n10563) );
  INV_X1 U11379 ( .A(keyinput_205), .ZN(n10696) );
  OAI22_X1 U11380 ( .A1(n10568), .A2(keyinput_202), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_203), .ZN(n10567) );
  AOI221_X1 U11381 ( .B1(n10568), .B2(keyinput_202), .C1(keyinput_203), .C2(
        P2_DATAO_REG_21__SCAN_IN), .A(n10567), .ZN(n10692) );
  INV_X1 U11382 ( .A(keyinput_201), .ZN(n10690) );
  INV_X1 U11383 ( .A(keyinput_200), .ZN(n10689) );
  INV_X1 U11384 ( .A(keyinput_199), .ZN(n10686) );
  OAI22_X1 U11385 ( .A1(n10570), .A2(keyinput_197), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_196), .ZN(n10569) );
  AOI221_X1 U11386 ( .B1(n10570), .B2(keyinput_197), .C1(keyinput_196), .C2(
        P2_DATAO_REG_28__SCAN_IN), .A(n10569), .ZN(n10683) );
  INV_X1 U11387 ( .A(keyinput_195), .ZN(n10680) );
  OAI22_X1 U11388 ( .A1(n10572), .A2(keyinput_186), .B1(keyinput_187), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10571) );
  AOI221_X1 U11389 ( .B1(n10572), .B2(keyinput_186), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_187), .A(n10571), .ZN(n10670) );
  OAI22_X1 U11390 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_183), .B1(
        keyinput_180), .B2(P2_REG3_REG_4__SCAN_IN), .ZN(n10573) );
  AOI221_X1 U11391 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_183), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_180), .A(n10573), .ZN(n10664) );
  OAI22_X1 U11392 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_181), .B1(
        keyinput_182), .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n10574) );
  AOI221_X1 U11393 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_181), .C1(
        P2_REG3_REG_0__SCAN_IN), .C2(keyinput_182), .A(n10574), .ZN(n10663) );
  OAI22_X1 U11394 ( .A1(n10577), .A2(keyinput_185), .B1(n10576), .B2(
        keyinput_184), .ZN(n10575) );
  AOI221_X1 U11395 ( .B1(n10577), .B2(keyinput_185), .C1(keyinput_184), .C2(
        n10576), .A(n10575), .ZN(n10662) );
  INV_X1 U11396 ( .A(keyinput_179), .ZN(n10661) );
  INV_X1 U11397 ( .A(keyinput_178), .ZN(n10659) );
  INV_X1 U11398 ( .A(keyinput_177), .ZN(n10657) );
  INV_X1 U11399 ( .A(keyinput_176), .ZN(n10654) );
  OAI22_X1 U11400 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_173), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_174), .ZN(n10578) );
  AOI221_X1 U11401 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_173), .C1(
        keyinput_174), .C2(P2_REG3_REG_12__SCAN_IN), .A(n10578), .ZN(n10651)
         );
  INV_X1 U11402 ( .A(keyinput_172), .ZN(n10648) );
  XNOR2_X1 U11403 ( .A(SI_4_), .B(keyinput_156), .ZN(n10639) );
  OAI22_X1 U11404 ( .A1(SI_11_), .A2(keyinput_149), .B1(SI_10_), .B2(
        keyinput_150), .ZN(n10579) );
  AOI221_X1 U11405 ( .B1(SI_11_), .B2(keyinput_149), .C1(keyinput_150), .C2(
        SI_10_), .A(n10579), .ZN(n10616) );
  INV_X1 U11406 ( .A(keyinput_147), .ZN(n10614) );
  OAI22_X1 U11407 ( .A1(SI_16_), .A2(keyinput_144), .B1(keyinput_145), .B2(
        SI_15_), .ZN(n10580) );
  AOI221_X1 U11408 ( .B1(SI_16_), .B2(keyinput_144), .C1(SI_15_), .C2(
        keyinput_145), .A(n10580), .ZN(n10610) );
  AOI22_X1 U11409 ( .A1(n10583), .A2(keyinput_142), .B1(n10582), .B2(
        keyinput_141), .ZN(n10581) );
  OAI221_X1 U11410 ( .B1(n10583), .B2(keyinput_142), .C1(n10582), .C2(
        keyinput_141), .A(n10581), .ZN(n10608) );
  OAI22_X1 U11411 ( .A1(n10586), .A2(keyinput_135), .B1(n10585), .B2(
        keyinput_136), .ZN(n10584) );
  AOI221_X1 U11412 ( .B1(n10586), .B2(keyinput_135), .C1(keyinput_136), .C2(
        n10585), .A(n10584), .ZN(n10604) );
  INV_X1 U11413 ( .A(keyinput_134), .ZN(n10596) );
  OAI22_X1 U11414 ( .A1(SI_31_), .A2(keyinput_129), .B1(keyinput_128), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n10587) );
  AOI221_X1 U11415 ( .B1(SI_31_), .B2(keyinput_129), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_128), .A(n10587), .ZN(n10594) );
  OAI221_X1 U11416 ( .B1(SI_30_), .B2(keyinput_130), .C1(n10589), .C2(
        keyinput_131), .A(n10588), .ZN(n10593) );
  OAI22_X1 U11417 ( .A1(n10591), .A2(keyinput_132), .B1(SI_27_), .B2(
        keyinput_133), .ZN(n10590) );
  AOI221_X1 U11418 ( .B1(n10591), .B2(keyinput_132), .C1(keyinput_133), .C2(
        SI_27_), .A(n10590), .ZN(n10592) );
  OAI21_X1 U11419 ( .B1(n10594), .B2(n10593), .A(n10592), .ZN(n10595) );
  OAI221_X1 U11420 ( .B1(SI_26_), .B2(keyinput_134), .C1(n10597), .C2(n10596), 
        .A(n10595), .ZN(n10603) );
  AOI22_X1 U11421 ( .A1(SI_21_), .A2(keyinput_139), .B1(n10599), .B2(
        keyinput_137), .ZN(n10598) );
  OAI221_X1 U11422 ( .B1(SI_21_), .B2(keyinput_139), .C1(n10599), .C2(
        keyinput_137), .A(n10598), .ZN(n10602) );
  AOI22_X1 U11423 ( .A1(SI_20_), .A2(keyinput_140), .B1(SI_22_), .B2(
        keyinput_138), .ZN(n10600) );
  OAI221_X1 U11424 ( .B1(SI_20_), .B2(keyinput_140), .C1(SI_22_), .C2(
        keyinput_138), .A(n10600), .ZN(n10601) );
  AOI211_X1 U11425 ( .C1(n10604), .C2(n10603), .A(n10602), .B(n10601), .ZN(
        n10607) );
  NAND2_X1 U11426 ( .A1(n10606), .A2(keyinput_143), .ZN(n10605) );
  OAI221_X1 U11427 ( .B1(n10608), .B2(n10607), .C1(n10606), .C2(keyinput_143), 
        .A(n10605), .ZN(n10609) );
  AOI22_X1 U11428 ( .A1(n10610), .A2(n10609), .B1(keyinput_146), .B2(SI_14_), 
        .ZN(n10611) );
  OAI21_X1 U11429 ( .B1(keyinput_146), .B2(SI_14_), .A(n10611), .ZN(n10612) );
  OAI221_X1 U11430 ( .B1(SI_13_), .B2(n10614), .C1(n10613), .C2(keyinput_147), 
        .A(n10612), .ZN(n10615) );
  AOI22_X1 U11431 ( .A1(n10619), .A2(keyinput_151), .B1(keyinput_152), .B2(
        n10618), .ZN(n10617) );
  OAI221_X1 U11432 ( .B1(n10619), .B2(keyinput_151), .C1(n10618), .C2(
        keyinput_152), .A(n10617), .ZN(n10624) );
  XNOR2_X1 U11433 ( .A(n10620), .B(keyinput_153), .ZN(n10623) );
  OAI22_X1 U11434 ( .A1(SI_6_), .A2(keyinput_154), .B1(SI_5_), .B2(
        keyinput_155), .ZN(n10621) );
  AOI221_X1 U11435 ( .B1(SI_6_), .B2(keyinput_154), .C1(keyinput_155), .C2(
        SI_5_), .A(n10621), .ZN(n10622) );
  AOI22_X1 U11436 ( .A1(P2_U3151), .A2(keyinput_162), .B1(keyinput_165), .B2(
        n10626), .ZN(n10625) );
  OAI221_X1 U11437 ( .B1(P2_U3151), .B2(keyinput_162), .C1(n10626), .C2(
        keyinput_165), .A(n10625), .ZN(n10638) );
  INV_X1 U11438 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10628) );
  OAI22_X1 U11439 ( .A1(n10628), .A2(keyinput_163), .B1(keyinput_161), .B2(
        P2_RD_REG_SCAN_IN), .ZN(n10627) );
  AOI221_X1 U11440 ( .B1(n10628), .B2(keyinput_163), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_161), .A(n10627), .ZN(n10636) );
  OAI22_X1 U11441 ( .A1(SI_3_), .A2(keyinput_157), .B1(keyinput_159), .B2(
        SI_1_), .ZN(n10629) );
  AOI221_X1 U11442 ( .B1(SI_3_), .B2(keyinput_157), .C1(SI_1_), .C2(
        keyinput_159), .A(n10629), .ZN(n10635) );
  OAI22_X1 U11443 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_164), .B1(SI_2_), .B2(keyinput_158), .ZN(n10630) );
  AOI221_X1 U11444 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_164), .C1(
        keyinput_158), .C2(SI_2_), .A(n10630), .ZN(n10634) );
  XOR2_X1 U11445 ( .A(SI_0_), .B(keyinput_160), .Z(n10632) );
  XNOR2_X1 U11446 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .ZN(n10631)
         );
  NOR2_X1 U11447 ( .A1(n10632), .A2(n10631), .ZN(n10633) );
  NAND4_X1 U11448 ( .A1(n10636), .A2(n10635), .A3(n10634), .A4(n10633), .ZN(
        n10637) );
  XOR2_X1 U11449 ( .A(n10640), .B(keyinput_167), .Z(n10645) );
  OAI22_X1 U11450 ( .A1(n7262), .A2(keyinput_170), .B1(n7193), .B2(
        keyinput_168), .ZN(n10641) );
  AOI221_X1 U11451 ( .B1(n7262), .B2(keyinput_170), .C1(keyinput_168), .C2(
        n7193), .A(n10641), .ZN(n10644) );
  OAI22_X1 U11452 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_169), .B1(
        keyinput_171), .B2(P2_REG3_REG_8__SCAN_IN), .ZN(n10642) );
  AOI221_X1 U11453 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_169), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_171), .A(n10642), .ZN(n10643) );
  OAI211_X1 U11454 ( .C1(n10646), .C2(n10645), .A(n10644), .B(n10643), .ZN(
        n10647) );
  OAI221_X1 U11455 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_172), .C1(
        n10649), .C2(n10648), .A(n10647), .ZN(n10650) );
  AOI22_X1 U11456 ( .A1(n10651), .A2(n10650), .B1(keyinput_175), .B2(
        P2_REG3_REG_25__SCAN_IN), .ZN(n10652) );
  OAI21_X1 U11457 ( .B1(keyinput_175), .B2(P2_REG3_REG_25__SCAN_IN), .A(n10652), .ZN(n10653) );
  OAI221_X1 U11458 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_176), .C1(
        n10655), .C2(n10654), .A(n10653), .ZN(n10656) );
  XNOR2_X1 U11459 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n10668)
         );
  AOI22_X1 U11460 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_190), .B1(
        n10666), .B2(keyinput_188), .ZN(n10665) );
  OAI221_X1 U11461 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_190), .C1(
        n10666), .C2(keyinput_188), .A(n10665), .ZN(n10667) );
  AOI211_X1 U11462 ( .C1(n10670), .C2(n10669), .A(n10668), .B(n10667), .ZN(
        n10678) );
  INV_X1 U11463 ( .A(P2_B_REG_SCAN_IN), .ZN(n10672) );
  AOI22_X1 U11464 ( .A1(n10673), .A2(keyinput_191), .B1(n10672), .B2(
        keyinput_192), .ZN(n10671) );
  OAI221_X1 U11465 ( .B1(n10673), .B2(keyinput_191), .C1(n10672), .C2(
        keyinput_192), .A(n10671), .ZN(n10677) );
  OAI22_X1 U11466 ( .A1(n10675), .A2(keyinput_194), .B1(keyinput_193), .B2(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n10674) );
  AOI221_X1 U11467 ( .B1(n10675), .B2(keyinput_194), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_193), .A(n10674), .ZN(n10676)
         );
  OAI21_X1 U11468 ( .B1(n10678), .B2(n10677), .A(n10676), .ZN(n10679) );
  OAI221_X1 U11469 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_195), .C1(
        n10681), .C2(n10680), .A(n10679), .ZN(n10682) );
  AOI22_X1 U11470 ( .A1(keyinput_198), .A2(n10685), .B1(n10683), .B2(n10682), 
        .ZN(n10684) );
  OAI211_X1 U11471 ( .C1(n10694), .C2(keyinput_204), .A(n10692), .B(n10691), 
        .ZN(n10693) );
  OAI22_X1 U11472 ( .A1(n10698), .A2(n10697), .B1(keyinput_217), .B2(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n10699) );
  AOI21_X1 U11473 ( .B1(keyinput_217), .B2(P2_DATAO_REG_7__SCAN_IN), .A(n10699), .ZN(n10708) );
  INV_X1 U11474 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U11475 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_218), .B1(n10701), 
        .B2(keyinput_219), .ZN(n10700) );
  OAI221_X1 U11476 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_218), .C1(n10701), 
        .C2(keyinput_219), .A(n10700), .ZN(n10707) );
  INV_X1 U11477 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10703) );
  OAI22_X1 U11478 ( .A1(n10703), .A2(keyinput_223), .B1(keyinput_222), .B2(
        P1_IR_REG_4__SCAN_IN), .ZN(n10702) );
  AOI221_X1 U11479 ( .B1(n10703), .B2(keyinput_223), .C1(P1_IR_REG_4__SCAN_IN), 
        .C2(keyinput_222), .A(n10702), .ZN(n10706) );
  OAI22_X1 U11480 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_220), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput_221), .ZN(n10704) );
  AOI221_X1 U11481 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_220), .C1(
        keyinput_221), .C2(P1_IR_REG_3__SCAN_IN), .A(n10704), .ZN(n10705) );
  OAI211_X1 U11482 ( .C1(n10708), .C2(n10707), .A(n10706), .B(n10705), .ZN(
        n10711) );
  INV_X1 U11483 ( .A(keyinput_224), .ZN(n10709) );
  MUX2_X1 U11484 ( .A(n10709), .B(keyinput_224), .S(P1_IR_REG_6__SCAN_IN), .Z(
        n10710) );
  NAND2_X1 U11485 ( .A1(n10711), .A2(n10710), .ZN(n10718) );
  OAI22_X1 U11486 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_225), .B1(
        keyinput_226), .B2(P1_IR_REG_8__SCAN_IN), .ZN(n10712) );
  AOI221_X1 U11487 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_225), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_226), .A(n10712), .ZN(n10717) );
  AOI22_X1 U11488 ( .A1(n10715), .A2(keyinput_227), .B1(n10714), .B2(
        keyinput_228), .ZN(n10713) );
  OAI221_X1 U11489 ( .B1(n10715), .B2(keyinput_227), .C1(n10714), .C2(
        keyinput_228), .A(n10713), .ZN(n10716) );
  XNOR2_X1 U11490 ( .A(n10721), .B(keyinput_234), .ZN(n10723) );
  XOR2_X1 U11491 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_232), .Z(n10722) );
  AOI211_X1 U11492 ( .C1(P1_IR_REG_12__SCAN_IN), .C2(keyinput_230), .A(n10723), 
        .B(n10722), .ZN(n10726) );
  XNOR2_X1 U11493 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_233), .ZN(n10725)
         );
  XNOR2_X1 U11494 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_231), .ZN(n10724)
         );
  AND3_X1 U11495 ( .A1(n10726), .A2(n10725), .A3(n10724), .ZN(n10727) );
  OAI21_X1 U11496 ( .B1(keyinput_230), .B2(P1_IR_REG_12__SCAN_IN), .A(n10727), 
        .ZN(n10733) );
  OAI22_X1 U11497 ( .A1(n10729), .A2(keyinput_235), .B1(P1_IR_REG_19__SCAN_IN), 
        .B2(keyinput_237), .ZN(n10728) );
  AOI221_X1 U11498 ( .B1(n10729), .B2(keyinput_235), .C1(keyinput_237), .C2(
        P1_IR_REG_19__SCAN_IN), .A(n10728), .ZN(n10732) );
  XOR2_X1 U11499 ( .A(n10730), .B(keyinput_236), .Z(n10731) );
  OAI22_X1 U11500 ( .A1(n10735), .A2(keyinput_238), .B1(n5798), .B2(
        keyinput_242), .ZN(n10734) );
  AOI221_X1 U11501 ( .B1(n10735), .B2(keyinput_238), .C1(keyinput_242), .C2(
        n5798), .A(n10734), .ZN(n10742) );
  XNOR2_X1 U11502 ( .A(n10736), .B(keyinput_240), .ZN(n10740) );
  XNOR2_X1 U11503 ( .A(n10737), .B(keyinput_239), .ZN(n10739) );
  XNOR2_X1 U11504 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_241), .ZN(n10738)
         );
  NOR3_X1 U11505 ( .A1(n10740), .A2(n10739), .A3(n10738), .ZN(n10741) );
  XNOR2_X1 U11506 ( .A(n10743), .B(keyinput_243), .ZN(n10746) );
  INV_X1 U11507 ( .A(keyinput_244), .ZN(n10744) );
  MUX2_X1 U11508 ( .A(keyinput_244), .B(n10744), .S(P1_IR_REG_26__SCAN_IN), 
        .Z(n10745) );
  OAI21_X1 U11509 ( .B1(n10747), .B2(n10746), .A(n10745), .ZN(n10751) );
  XNOR2_X1 U11510 ( .A(n10748), .B(keyinput_245), .ZN(n10750) );
  XNOR2_X1 U11511 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_246), .ZN(n10749)
         );
  XOR2_X1 U11512 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_247), .Z(n10754) );
  XOR2_X1 U11513 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .Z(n10753) );
  XNOR2_X1 U11514 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_248), .ZN(n10752)
         );
  AOI22_X1 U11515 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_251), .B1(
        P1_D_REG_0__SCAN_IN), .B2(keyinput_250), .ZN(n10755) );
  OAI221_X1 U11516 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_251), .C1(
        P1_D_REG_0__SCAN_IN), .C2(keyinput_250), .A(n10755), .ZN(n10756) );
  AOI22_X1 U11517 ( .A1(n10759), .A2(keyinput_255), .B1(n10758), .B2(
        keyinput_254), .ZN(n10757) );
  OAI221_X1 U11518 ( .B1(n10759), .B2(keyinput_255), .C1(n10758), .C2(
        keyinput_254), .A(n10757), .ZN(n10763) );
  AOI22_X1 U11519 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_253), .B1(n10761), 
        .B2(keyinput_252), .ZN(n10760) );
  OAI221_X1 U11520 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_253), .C1(n10761), 
        .C2(keyinput_252), .A(n10760), .ZN(n10762) );
  XNOR2_X1 U11521 ( .A(n10766), .B(n10765), .ZN(P2_U3189) );
  XOR2_X1 U11522 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI222_X1 U11523 ( .A1(n10771), .A2(n10770), .B1(n10771), .B2(n10769), .C1(
        n10768), .C2(n10767), .ZN(ADD_1068_U5) );
  AOI21_X1 U11524 ( .B1(n10774), .B2(n10773), .A(n10772), .ZN(ADD_1068_U54) );
  AOI21_X1 U11525 ( .B1(n10777), .B2(n10776), .A(n10775), .ZN(ADD_1068_U53) );
  OAI21_X1 U11526 ( .B1(n10780), .B2(n10779), .A(n10778), .ZN(ADD_1068_U52) );
  OAI21_X1 U11527 ( .B1(n10783), .B2(n10782), .A(n10781), .ZN(ADD_1068_U51) );
  OAI21_X1 U11528 ( .B1(n10786), .B2(n10785), .A(n10784), .ZN(ADD_1068_U50) );
  OAI21_X1 U11529 ( .B1(n10789), .B2(n10788), .A(n10787), .ZN(ADD_1068_U49) );
  OAI21_X1 U11530 ( .B1(n10792), .B2(n10791), .A(n10790), .ZN(ADD_1068_U48) );
  OAI21_X1 U11531 ( .B1(n10795), .B2(n10794), .A(n10793), .ZN(ADD_1068_U47) );
  OAI21_X1 U11532 ( .B1(n10798), .B2(n10797), .A(n10796), .ZN(ADD_1068_U63) );
  OAI21_X1 U11533 ( .B1(n10801), .B2(n10800), .A(n10799), .ZN(ADD_1068_U62) );
  OAI21_X1 U11534 ( .B1(n10804), .B2(n10803), .A(n10802), .ZN(ADD_1068_U61) );
  OAI21_X1 U11535 ( .B1(n10807), .B2(n10806), .A(n10805), .ZN(ADD_1068_U60) );
  OAI21_X1 U11536 ( .B1(n10810), .B2(n10809), .A(n10808), .ZN(ADD_1068_U59) );
  OAI21_X1 U11537 ( .B1(n10813), .B2(n10812), .A(n10811), .ZN(ADD_1068_U58) );
  OAI21_X1 U11538 ( .B1(n10816), .B2(n10815), .A(n10814), .ZN(ADD_1068_U57) );
  OAI21_X1 U11539 ( .B1(n10819), .B2(n10818), .A(n10817), .ZN(ADD_1068_U56) );
  OAI21_X1 U11540 ( .B1(n10822), .B2(n10821), .A(n10820), .ZN(ADD_1068_U55) );
  NAND2_X1 U11541 ( .A1(n10823), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10824) );
  OAI21_X1 U11542 ( .B1(n10826), .B2(n10825), .A(n10824), .ZN(n10827) );
  XOR2_X1 U11543 ( .A(n10827), .B(n5360), .Z(n10829) );
  AOI22_X1 U11544 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10861), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10828) );
  OAI21_X1 U11545 ( .B1(n10830), .B2(n10829), .A(n10828), .ZN(P1_U3243) );
  AOI22_X1 U11546 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10861), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10842) );
  AOI211_X1 U11547 ( .C1(n10833), .C2(n10832), .A(n10831), .B(n10862), .ZN(
        n10834) );
  AOI21_X1 U11548 ( .B1(n10869), .B2(n10835), .A(n10834), .ZN(n10841) );
  INV_X1 U11549 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10836) );
  NOR2_X1 U11550 ( .A1(n5360), .A2(n10836), .ZN(n10839) );
  OAI211_X1 U11551 ( .C1(n10839), .C2(n10838), .A(n10871), .B(n10837), .ZN(
        n10840) );
  NAND3_X1 U11552 ( .A1(n10842), .A2(n10841), .A3(n10840), .ZN(P1_U3244) );
  INV_X1 U11553 ( .A(n10861), .ZN(n10859) );
  INV_X1 U11554 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10858) );
  OAI21_X1 U11555 ( .B1(n10845), .B2(n10844), .A(n10843), .ZN(n10854) );
  AOI21_X1 U11556 ( .B1(n10848), .B2(n10847), .A(n10846), .ZN(n10852) );
  OAI22_X1 U11557 ( .A1(n10852), .A2(n10851), .B1(n10850), .B2(n10849), .ZN(
        n10853) );
  AOI21_X1 U11558 ( .B1(n10855), .B2(n10854), .A(n10853), .ZN(n10857) );
  OAI211_X1 U11559 ( .C1(n10859), .C2(n10858), .A(n10857), .B(n10856), .ZN(
        P1_U3255) );
  XOR2_X1 U11560 ( .A(n5228), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  AOI21_X1 U11561 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n10861), .A(n10860), .ZN(
        n10876) );
  AOI211_X1 U11562 ( .C1(n10865), .C2(n10864), .A(n10863), .B(n10862), .ZN(
        n10867) );
  AOI211_X1 U11563 ( .C1(n10869), .C2(n10868), .A(n10867), .B(n10866), .ZN(
        n10875) );
  OAI211_X1 U11564 ( .C1(n10873), .C2(n10872), .A(n10871), .B(n10870), .ZN(
        n10874) );
  NAND3_X1 U11565 ( .A1(n10876), .A2(n10875), .A3(n10874), .ZN(P1_U3247) );
  INV_X1 U11566 ( .A(n10877), .ZN(n11097) );
  INV_X1 U11567 ( .A(n10878), .ZN(n10883) );
  OAI21_X1 U11568 ( .B1(n10880), .B2(n11141), .A(n10879), .ZN(n10882) );
  AOI211_X1 U11569 ( .C1(n11097), .C2(n10883), .A(n10882), .B(n10881), .ZN(
        n10884) );
  AOI22_X1 U11570 ( .A1(n11147), .A2(n10884), .B1(n6803), .B2(n11146), .ZN(
        P1_U3523) );
  AOI22_X1 U11571 ( .A1(n11150), .A2(n10884), .B1(n5875), .B2(n11148), .ZN(
        P1_U3456) );
  NOR2_X1 U11572 ( .A1(n10886), .A2(n10885), .ZN(n10890) );
  OAI21_X1 U11573 ( .B1(n10888), .B2(n11141), .A(n10887), .ZN(n10889) );
  NOR3_X1 U11574 ( .A1(n10891), .A2(n10890), .A3(n10889), .ZN(n10892) );
  AOI22_X1 U11575 ( .A1(n11147), .A2(n10892), .B1(n6802), .B2(n11146), .ZN(
        P1_U3524) );
  AOI22_X1 U11576 ( .A1(n11150), .A2(n10892), .B1(n5778), .B2(n11148), .ZN(
        P1_U3459) );
  INV_X1 U11577 ( .A(n10893), .ZN(n10897) );
  OR2_X1 U11578 ( .A1(n10894), .A2(n10938), .ZN(n10895) );
  AND3_X1 U11579 ( .A1(n10897), .A2(n10896), .A3(n10895), .ZN(n10900) );
  AOI22_X1 U11580 ( .A1(n11127), .A2(n10900), .B1(n10898), .B2(n11126), .ZN(
        P2_U3461) );
  INV_X1 U11581 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U11582 ( .A1(n11131), .A2(n10900), .B1(n10899), .B2(n11128), .ZN(
        P2_U3396) );
  XNOR2_X1 U11583 ( .A(n10901), .B(n10908), .ZN(n10926) );
  INV_X1 U11584 ( .A(n10902), .ZN(n10904) );
  OAI211_X1 U11585 ( .C1(n10904), .C2(n10921), .A(n11006), .B(n10903), .ZN(
        n10924) );
  OAI21_X1 U11586 ( .B1(n10921), .B2(n11141), .A(n10924), .ZN(n10916) );
  INV_X1 U11587 ( .A(n10905), .ZN(n11021) );
  OAI22_X1 U11588 ( .A1(n10907), .A2(n11010), .B1(n10906), .B2(n11008), .ZN(
        n10914) );
  NAND3_X1 U11589 ( .A1(n10910), .A2(n10909), .A3(n10908), .ZN(n10911) );
  AOI21_X1 U11590 ( .B1(n10912), .B2(n10911), .A(n11016), .ZN(n10913) );
  AOI211_X1 U11591 ( .C1(n11021), .C2(n10926), .A(n10914), .B(n10913), .ZN(
        n10929) );
  INV_X1 U11592 ( .A(n10929), .ZN(n10915) );
  AOI211_X1 U11593 ( .C1(n11097), .C2(n10926), .A(n10916), .B(n10915), .ZN(
        n10918) );
  INV_X1 U11594 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U11595 ( .A1(n11147), .A2(n10918), .B1(n10917), .B2(n11146), .ZN(
        P1_U3525) );
  AOI22_X1 U11596 ( .A1(n11150), .A2(n10918), .B1(n5895), .B2(n11148), .ZN(
        P1_U3462) );
  AOI22_X1 U11597 ( .A1(n11028), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n11026), 
        .B2(n10919), .ZN(n10920) );
  OAI21_X1 U11598 ( .B1(n11031), .B2(n10921), .A(n10920), .ZN(n10922) );
  INV_X1 U11599 ( .A(n10922), .ZN(n10928) );
  INV_X1 U11600 ( .A(n10923), .ZN(n11036) );
  INV_X1 U11601 ( .A(n10924), .ZN(n10925) );
  AOI22_X1 U11602 ( .A1(n10926), .A2(n11036), .B1(n11035), .B2(n10925), .ZN(
        n10927) );
  OAI211_X1 U11603 ( .C1(n10180), .C2(n10929), .A(n10928), .B(n10927), .ZN(
        P1_U3290) );
  AOI22_X1 U11604 ( .A1(n10931), .A2(n11119), .B1(n11121), .B2(n10930), .ZN(
        n10932) );
  AND2_X1 U11605 ( .A1(n10933), .A2(n10932), .ZN(n10936) );
  AOI22_X1 U11606 ( .A1(n11127), .A2(n10936), .B1(n10934), .B2(n11126), .ZN(
        P2_U3462) );
  INV_X1 U11607 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U11608 ( .A1(n11131), .A2(n10936), .B1(n10935), .B2(n11128), .ZN(
        P2_U3399) );
  OAI22_X1 U11609 ( .A1(n10939), .A2(n10938), .B1(n10937), .B2(n10987), .ZN(
        n10941) );
  NOR2_X1 U11610 ( .A1(n10941), .A2(n10940), .ZN(n10944) );
  AOI22_X1 U11611 ( .A1(n11127), .A2(n10944), .B1(n10942), .B2(n11126), .ZN(
        P2_U3463) );
  INV_X1 U11612 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U11613 ( .A1(n11131), .A2(n10944), .B1(n10943), .B2(n11128), .ZN(
        P2_U3402) );
  OAI21_X1 U11614 ( .B1(n10946), .B2(n11141), .A(n10945), .ZN(n10947) );
  AOI21_X1 U11615 ( .B1(n10948), .B2(n11144), .A(n10947), .ZN(n10949) );
  AND2_X1 U11616 ( .A1(n10950), .A2(n10949), .ZN(n10951) );
  AOI22_X1 U11617 ( .A1(n11147), .A2(n10951), .B1(n6808), .B2(n11146), .ZN(
        P1_U3526) );
  AOI22_X1 U11618 ( .A1(n11150), .A2(n10951), .B1(n5921), .B2(n11148), .ZN(
        P1_U3465) );
  INV_X1 U11619 ( .A(n10952), .ZN(n10957) );
  OAI22_X1 U11620 ( .A1(n10955), .A2(n10954), .B1(n10953), .B2(n10987), .ZN(
        n10956) );
  NOR2_X1 U11621 ( .A1(n10957), .A2(n10956), .ZN(n10960) );
  AOI22_X1 U11622 ( .A1(n11127), .A2(n10960), .B1(n10958), .B2(n11126), .ZN(
        P2_U3464) );
  INV_X1 U11623 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U11624 ( .A1(n11131), .A2(n10960), .B1(n10959), .B2(n11128), .ZN(
        P2_U3405) );
  XNOR2_X1 U11625 ( .A(n10961), .B(n10966), .ZN(n10983) );
  INV_X1 U11626 ( .A(n10962), .ZN(n10963) );
  OAI211_X1 U11627 ( .C1(n10978), .C2(n10964), .A(n10963), .B(n11006), .ZN(
        n10980) );
  OAI21_X1 U11628 ( .B1(n10978), .B2(n11141), .A(n10980), .ZN(n10974) );
  XOR2_X1 U11629 ( .A(n10966), .B(n10965), .Z(n10971) );
  AOI222_X1 U11630 ( .A1(n10972), .A2(n10971), .B1(n10970), .B2(n10969), .C1(
        n10968), .C2(n10967), .ZN(n10986) );
  INV_X1 U11631 ( .A(n10986), .ZN(n10973) );
  AOI211_X1 U11632 ( .C1(n11144), .C2(n10983), .A(n10974), .B(n10973), .ZN(
        n10975) );
  AOI22_X1 U11633 ( .A1(n11147), .A2(n10975), .B1(n6809), .B2(n11146), .ZN(
        P1_U3527) );
  AOI22_X1 U11634 ( .A1(n11150), .A2(n10975), .B1(n5955), .B2(n11148), .ZN(
        P1_U3468) );
  AOI22_X1 U11635 ( .A1(n11028), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n10976), 
        .B2(n11026), .ZN(n10977) );
  OAI21_X1 U11636 ( .B1(n11031), .B2(n10978), .A(n10977), .ZN(n10979) );
  INV_X1 U11637 ( .A(n10979), .ZN(n10985) );
  INV_X1 U11638 ( .A(n10980), .ZN(n10981) );
  AOI22_X1 U11639 ( .A1(n10983), .A2(n10982), .B1(n11035), .B2(n10981), .ZN(
        n10984) );
  OAI211_X1 U11640 ( .C1(n10180), .C2(n10986), .A(n10985), .B(n10984), .ZN(
        P1_U3288) );
  NOR2_X1 U11641 ( .A1(n10988), .A2(n10987), .ZN(n10990) );
  AOI211_X1 U11642 ( .C1(n11119), .C2(n10991), .A(n10990), .B(n10989), .ZN(
        n10994) );
  AOI22_X1 U11643 ( .A1(n11127), .A2(n10994), .B1(n10992), .B2(n11126), .ZN(
        P2_U3465) );
  INV_X1 U11644 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10993) );
  AOI22_X1 U11645 ( .A1(n11131), .A2(n10994), .B1(n10993), .B2(n11128), .ZN(
        P2_U3408) );
  AND2_X1 U11646 ( .A1(n10995), .A2(n11144), .ZN(n11000) );
  OAI21_X1 U11647 ( .B1(n10997), .B2(n11141), .A(n10996), .ZN(n10998) );
  NOR3_X1 U11648 ( .A1(n11000), .A2(n10999), .A3(n10998), .ZN(n11002) );
  AOI22_X1 U11649 ( .A1(n11147), .A2(n11002), .B1(n11001), .B2(n11146), .ZN(
        P1_U3528) );
  AOI22_X1 U11650 ( .A1(n11150), .A2(n11002), .B1(n5974), .B2(n11148), .ZN(
        P1_U3471) );
  XNOR2_X1 U11651 ( .A(n11003), .B(n11013), .ZN(n11037) );
  INV_X1 U11652 ( .A(n11004), .ZN(n11007) );
  OAI211_X1 U11653 ( .C1(n11007), .C2(n11030), .A(n11006), .B(n11005), .ZN(
        n11033) );
  OAI21_X1 U11654 ( .B1(n11030), .B2(n11141), .A(n11033), .ZN(n11023) );
  OAI22_X1 U11655 ( .A1(n11011), .A2(n11010), .B1(n11009), .B2(n11008), .ZN(
        n11020) );
  INV_X1 U11656 ( .A(n11012), .ZN(n11015) );
  OAI21_X1 U11657 ( .B1(n11015), .B2(n11014), .A(n11013), .ZN(n11018) );
  AOI21_X1 U11658 ( .B1(n11018), .B2(n11017), .A(n11016), .ZN(n11019) );
  AOI211_X1 U11659 ( .C1(n11021), .C2(n11037), .A(n11020), .B(n11019), .ZN(
        n11040) );
  INV_X1 U11660 ( .A(n11040), .ZN(n11022) );
  AOI211_X1 U11661 ( .C1(n11097), .C2(n11037), .A(n11023), .B(n11022), .ZN(
        n11025) );
  AOI22_X1 U11662 ( .A1(n11147), .A2(n11025), .B1(n11024), .B2(n11146), .ZN(
        P1_U3529) );
  AOI22_X1 U11663 ( .A1(n11150), .A2(n11025), .B1(n6008), .B2(n11148), .ZN(
        P1_U3474) );
  AOI22_X1 U11664 ( .A1(n11028), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n11027), 
        .B2(n11026), .ZN(n11029) );
  OAI21_X1 U11665 ( .B1(n11031), .B2(n11030), .A(n11029), .ZN(n11032) );
  INV_X1 U11666 ( .A(n11032), .ZN(n11039) );
  INV_X1 U11667 ( .A(n11033), .ZN(n11034) );
  AOI22_X1 U11668 ( .A1(n11037), .A2(n11036), .B1(n11035), .B2(n11034), .ZN(
        n11038) );
  OAI211_X1 U11669 ( .C1(n10180), .C2(n11040), .A(n11039), .B(n11038), .ZN(
        P1_U3286) );
  OAI22_X1 U11670 ( .A1(n11043), .A2(n11042), .B1(n11041), .B2(n11141), .ZN(
        n11045) );
  AOI211_X1 U11671 ( .C1(n11046), .C2(n11144), .A(n11045), .B(n11044), .ZN(
        n11047) );
  AOI22_X1 U11672 ( .A1(n11147), .A2(n11047), .B1(n7099), .B2(n11146), .ZN(
        P1_U3530) );
  AOI22_X1 U11673 ( .A1(n11150), .A2(n11047), .B1(n6031), .B2(n11148), .ZN(
        P1_U3477) );
  OAI211_X1 U11674 ( .C1(n11050), .C2(n11141), .A(n11049), .B(n11048), .ZN(
        n11051) );
  AOI21_X1 U11675 ( .B1(n11052), .B2(n11144), .A(n11051), .ZN(n11053) );
  AOI22_X1 U11676 ( .A1(n11147), .A2(n11053), .B1(n7321), .B2(n11146), .ZN(
        P1_U3531) );
  AOI22_X1 U11677 ( .A1(n11150), .A2(n11053), .B1(n6073), .B2(n11148), .ZN(
        P1_U3480) );
  OAI21_X1 U11678 ( .B1(n5681), .B2(n11141), .A(n11054), .ZN(n11056) );
  AOI211_X1 U11679 ( .C1(n11144), .C2(n11057), .A(n11056), .B(n11055), .ZN(
        n11058) );
  AOI22_X1 U11680 ( .A1(n11147), .A2(n11058), .B1(n7368), .B2(n11146), .ZN(
        P1_U3532) );
  AOI22_X1 U11681 ( .A1(n11150), .A2(n11058), .B1(n6096), .B2(n11148), .ZN(
        P1_U3483) );
  AND2_X1 U11682 ( .A1(n11059), .A2(n11119), .ZN(n11063) );
  AND2_X1 U11683 ( .A1(n11060), .A2(n11121), .ZN(n11061) );
  NOR3_X1 U11684 ( .A1(n11063), .A2(n11062), .A3(n11061), .ZN(n11065) );
  AOI22_X1 U11685 ( .A1(n11127), .A2(n11065), .B1(n7838), .B2(n11126), .ZN(
        P2_U3469) );
  INV_X1 U11686 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U11687 ( .A1(n11131), .A2(n11065), .B1(n11064), .B2(n11128), .ZN(
        P2_U3420) );
  OAI21_X1 U11688 ( .B1(n11068), .B2(n11067), .A(n11066), .ZN(n11076) );
  OR3_X1 U11689 ( .A1(n11071), .A2(n11070), .A3(n11069), .ZN(n11073) );
  AOI21_X1 U11690 ( .B1(n11074), .B2(n11073), .A(n11072), .ZN(n11075) );
  AOI211_X1 U11691 ( .C1(n11085), .C2(n11077), .A(n11076), .B(n11075), .ZN(
        n11078) );
  OAI21_X1 U11692 ( .B1(n11080), .B2(n11079), .A(n11078), .ZN(P2_U3176) );
  AOI21_X1 U11693 ( .B1(n11083), .B2(n11082), .A(n11081), .ZN(n11084) );
  INV_X1 U11694 ( .A(n11084), .ZN(n11088) );
  AOI222_X1 U11695 ( .A1(n11111), .A2(n11088), .B1(n11087), .B2(n11086), .C1(
        n11085), .C2(n11106), .ZN(n11089) );
  OAI21_X1 U11696 ( .B1(n11111), .B2(n11090), .A(n11089), .ZN(P2_U3222) );
  INV_X1 U11697 ( .A(n11091), .ZN(n11096) );
  OAI21_X1 U11698 ( .B1(n11093), .B2(n11141), .A(n11092), .ZN(n11095) );
  AOI211_X1 U11699 ( .C1(n11097), .C2(n11096), .A(n11095), .B(n11094), .ZN(
        n11098) );
  AOI22_X1 U11700 ( .A1(n11147), .A2(n11098), .B1(n7481), .B2(n11146), .ZN(
        P1_U3533) );
  AOI22_X1 U11701 ( .A1(n11150), .A2(n11098), .B1(n6126), .B2(n11148), .ZN(
        P1_U3486) );
  INV_X1 U11702 ( .A(n11099), .ZN(n11103) );
  INV_X1 U11703 ( .A(n11100), .ZN(n11101) );
  OAI21_X1 U11704 ( .B1(n11103), .B2(n11102), .A(n11101), .ZN(n11108) );
  AOI222_X1 U11705 ( .A1(n11108), .A2(n11111), .B1(n11107), .B2(n11106), .C1(
        n11105), .C2(n11104), .ZN(n11109) );
  OAI21_X1 U11706 ( .B1(n11111), .B2(n11110), .A(n11109), .ZN(P2_U3221) );
  OAI211_X1 U11707 ( .C1(n11114), .C2(n11141), .A(n11113), .B(n11112), .ZN(
        n11115) );
  AOI21_X1 U11708 ( .B1(n11116), .B2(n11144), .A(n11115), .ZN(n11118) );
  AOI22_X1 U11709 ( .A1(n11147), .A2(n11118), .B1(n11117), .B2(n11146), .ZN(
        P1_U3535) );
  AOI22_X1 U11710 ( .A1(n11150), .A2(n11118), .B1(n6178), .B2(n11148), .ZN(
        P1_U3492) );
  AND2_X1 U11711 ( .A1(n11120), .A2(n11119), .ZN(n11125) );
  AND2_X1 U11712 ( .A1(n11122), .A2(n11121), .ZN(n11123) );
  NOR3_X1 U11713 ( .A1(n11125), .A2(n11124), .A3(n11123), .ZN(n11130) );
  AOI22_X1 U11714 ( .A1(n11127), .A2(n11130), .B1(n8305), .B2(n11126), .ZN(
        P2_U3472) );
  INV_X1 U11715 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U11716 ( .A1(n11131), .A2(n11130), .B1(n11129), .B2(n11128), .ZN(
        P2_U3429) );
  OAI211_X1 U11717 ( .C1(n11134), .C2(n11141), .A(n11133), .B(n11132), .ZN(
        n11135) );
  AOI21_X1 U11718 ( .B1(n11136), .B2(n11144), .A(n11135), .ZN(n11138) );
  INV_X1 U11719 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U11720 ( .A1(n11147), .A2(n11138), .B1(n11137), .B2(n11146), .ZN(
        P1_U3537) );
  AOI22_X1 U11721 ( .A1(n11150), .A2(n11138), .B1(n6234), .B2(n11148), .ZN(
        P1_U3498) );
  OAI211_X1 U11722 ( .C1(n11142), .C2(n11141), .A(n11140), .B(n11139), .ZN(
        n11143) );
  AOI21_X1 U11723 ( .B1(n11145), .B2(n11144), .A(n11143), .ZN(n11149) );
  AOI22_X1 U11724 ( .A1(n11147), .A2(n11149), .B1(n9934), .B2(n11146), .ZN(
        P1_U3539) );
  AOI22_X1 U11725 ( .A1(n11150), .A2(n11149), .B1(n6284), .B2(n11148), .ZN(
        P1_U3504) );
  XNOR2_X1 U11726 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X1 U5157 ( .A(n5913), .Z(n6548) );
  CLKBUF_X1 U5165 ( .A(n5099), .Z(n7035) );
  CLKBUF_X1 U5167 ( .A(n5992), .Z(n6561) );
  CLKBUF_X3 U5205 ( .A(n5090), .Z(n5101) );
  CLKBUF_X1 U5222 ( .A(n7037), .Z(n8884) );
  CLKBUF_X1 U5492 ( .A(n7231), .Z(n5103) );
  NAND3_X1 U6177 ( .A1(n5925), .A2(n5924), .A3(n5923), .ZN(n10968) );
endmodule

