

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7189, n7190, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233;

  INV_X1 U7290 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n15913) );
  OR2_X1 U7291 ( .A1(n11669), .A2(n11668), .ZN(n11898) );
  INV_X1 U7292 ( .A(n15094), .ZN(n15050) );
  CLKBUF_X2 U7293 ( .A(n11678), .Z(n14267) );
  AND2_X1 U7294 ( .A1(n8721), .A2(n8720), .ZN(n12295) );
  INV_X1 U7295 ( .A(n10024), .ZN(n10044) );
  INV_X1 U7296 ( .A(n10691), .ZN(n12835) );
  CLKBUF_X2 U7297 ( .A(n10756), .Z(n12966) );
  INV_X2 U7298 ( .A(n13051), .ZN(n13004) );
  NAND2_X1 U7299 ( .A1(n7726), .A2(n7723), .ZN(n13321) );
  INV_X1 U7300 ( .A(n15913), .ZN(n7189) );
  INV_X1 U7301 ( .A(n7189), .ZN(n7190) );
  INV_X1 U7302 ( .A(n7189), .ZN(P1_U3086) );
  AND2_X1 U7303 ( .A1(n8394), .A2(n8477), .ZN(n8393) );
  INV_X1 U7304 ( .A(n14352), .ZN(n14304) );
  NOR2_X2 U7305 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8643) );
  INV_X1 U7306 ( .A(n15062), .ZN(n15096) );
  NAND2_X1 U7307 ( .A1(n7486), .A2(n7485), .ZN(n11823) );
  BUF_X1 U7308 ( .A(n9405), .Z(n10431) );
  CLKBUF_X2 U7309 ( .A(n11099), .Z(n13405) );
  NAND2_X1 U7310 ( .A1(n7924), .A2(n7923), .ZN(n7922) );
  INV_X1 U7311 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7446) );
  NOR2_X1 U7312 ( .A1(n8415), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8414) );
  INV_X1 U7313 ( .A(n11714), .ZN(n7486) );
  INV_X1 U7314 ( .A(n8288), .ZN(n12742) );
  INV_X1 U7315 ( .A(n10410), .ZN(n16096) );
  XNOR2_X1 U7316 ( .A(n13809), .B(n7449), .ZN(n13790) );
  NAND2_X1 U7317 ( .A1(n14342), .A2(n14341), .ZN(n14340) );
  NAND2_X1 U7318 ( .A1(n11808), .A2(n11807), .ZN(n16152) );
  NAND2_X1 U7319 ( .A1(n10210), .A2(n10209), .ZN(n12733) );
  XOR2_X1 U7320 ( .A(n10211), .B(P1_IR_REG_31__SCAN_IN), .Z(n7192) );
  NAND2_X1 U7321 ( .A1(n8393), .A2(n8643), .ZN(n8675) );
  OR2_X2 U7322 ( .A1(n12302), .A2(n7926), .ZN(n7925) );
  AOI21_X2 U7323 ( .B1(n13928), .B2(n8046), .A(n7261), .ZN(n8045) );
  NOR2_X2 U7324 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8481) );
  MUX2_X2 U7325 ( .A(n14205), .B(n14204), .S(n16232), .Z(n14206) );
  MUX2_X2 U7326 ( .A(n14131), .B(n14204), .S(n16228), .Z(n14132) );
  XNOR2_X1 U7327 ( .A(n14482), .B(n9900), .ZN(n10994) );
  OAI211_X2 U7328 ( .C1(n10024), .C2(n10748), .A(n8660), .B(n8659), .ZN(n9900)
         );
  NAND2_X2 U7329 ( .A1(n10691), .A2(n9343), .ZN(n12987) );
  BUF_X2 U7330 ( .A(n11522), .Z(n7193) );
  OR2_X2 U7331 ( .A1(n10617), .A2(n10493), .ZN(n13755) );
  AND3_X1 U7332 ( .A1(n10116), .A2(n8503), .A3(n10832), .ZN(n10034) );
  XNOR2_X2 U7333 ( .A(n7386), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8503) );
  OAI222_X1 U7334 ( .A1(n10526), .A2(P3_U3151), .B1(n13319), .B2(n10174), .C1(
        n10173), .C2(n14252), .ZN(P3_U3294) );
  OAI21_X2 U7335 ( .B1(n10526), .B2(n10514), .A(n10515), .ZN(n10563) );
  XNOR2_X2 U7336 ( .A(n9358), .B(P3_IR_REG_30__SCAN_IN), .ZN(n9360) );
  NOR2_X2 U7337 ( .A1(n15946), .A2(n9188), .ZN(n15994) );
  AOI22_X1 U7338 ( .A1(n10004), .A2(n10003), .B1(n7384), .B2(n10002), .ZN(
        n10007) );
  OR2_X1 U7339 ( .A1(n12661), .A2(n12660), .ZN(n15366) );
  INV_X2 U7340 ( .A(n10057), .ZN(n10085) );
  NAND2_X1 U7341 ( .A1(n8680), .A2(n7728), .ZN(n11603) );
  INV_X1 U7343 ( .A(n12762), .ZN(n16070) );
  INV_X4 U7344 ( .A(n10055), .ZN(n7194) );
  INV_X1 U7345 ( .A(n15234), .ZN(n11239) );
  CLKBUF_X1 U7346 ( .A(n10725), .Z(n15109) );
  INV_X1 U7347 ( .A(n13521), .ZN(n7730) );
  XNOR2_X1 U7348 ( .A(n8139), .B(n8655), .ZN(n10748) );
  NAND2_X1 U7349 ( .A1(n9790), .A2(n7234), .ZN(n10956) );
  INV_X4 U7350 ( .A(n7251), .ZN(n15065) );
  INV_X4 U7351 ( .A(n15095), .ZN(n11123) );
  NAND2_X2 U7352 ( .A1(n10290), .A2(n15351), .ZN(n10691) );
  INV_X2 U7353 ( .A(n8610), .ZN(n12718) );
  NAND2_X1 U7354 ( .A1(n12264), .A2(n9342), .ZN(n9405) );
  MUX2_X1 U7355 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10208), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n10210) );
  OR2_X1 U7356 ( .A1(n10214), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n10378) );
  AND2_X1 U7357 ( .A1(n8057), .A2(n8058), .ZN(n11612) );
  AND2_X1 U7358 ( .A1(n7258), .A2(n8414), .ZN(n8412) );
  OAI21_X1 U7359 ( .B1(n9805), .B2(n16039), .A(n9804), .ZN(n13907) );
  OAI21_X1 U7360 ( .B1(n9247), .B2(n16206), .A(n8137), .ZN(n9246) );
  INV_X1 U7361 ( .A(n7784), .ZN(n7783) );
  OAI21_X1 U7362 ( .B1(n15647), .B2(n16116), .A(n15645), .ZN(n7784) );
  NOR2_X1 U7363 ( .A1(n15436), .A2(n7243), .ZN(n15647) );
  XNOR2_X1 U7364 ( .A(n8177), .B(n15412), .ZN(n15629) );
  OAI21_X1 U7365 ( .B1(n8069), .B2(n16180), .A(n8066), .ZN(n7706) );
  NOR2_X1 U7366 ( .A1(n9233), .A2(n10110), .ZN(n9235) );
  OR2_X1 U7367 ( .A1(n15628), .A2(n16074), .ZN(n8069) );
  AOI21_X1 U7368 ( .B1(n7693), .B2(n9112), .A(n7691), .ZN(n14821) );
  NOR2_X1 U7369 ( .A1(n15465), .A2(n15408), .ZN(n15454) );
  OR2_X1 U7370 ( .A1(n14440), .A2(n14439), .ZN(n14442) );
  OR2_X1 U7371 ( .A1(n7635), .A2(n7633), .ZN(n7625) );
  NOR2_X1 U7372 ( .A1(n9109), .A2(n8466), .ZN(n9111) );
  OR2_X1 U7373 ( .A1(n15466), .A2(n15469), .ZN(n8187) );
  NAND2_X1 U7374 ( .A1(n15168), .A2(n15170), .ZN(n15169) );
  NAND2_X1 U7375 ( .A1(n15480), .A2(n7545), .ZN(n15466) );
  NAND2_X1 U7376 ( .A1(n13993), .A2(n13194), .ZN(n13980) );
  NAND2_X1 U7377 ( .A1(n8108), .A2(n8110), .ZN(n15468) );
  AOI21_X1 U7378 ( .B1(n7847), .B2(n14399), .A(n14303), .ZN(n7850) );
  XNOR2_X1 U7379 ( .A(n14298), .B(n14296), .ZN(n14335) );
  AOI21_X1 U7380 ( .B1(n7221), .B2(n13838), .A(n7700), .ZN(n13875) );
  NAND2_X1 U7381 ( .A1(n14419), .A2(n14422), .ZN(n14421) );
  OR2_X1 U7382 ( .A1(n14035), .A2(n14034), .ZN(n14033) );
  OAI21_X1 U7383 ( .B1(n14340), .B2(n7869), .A(n7868), .ZN(n14294) );
  AOI21_X1 U7384 ( .B1(n13398), .B2(n7650), .A(n7648), .ZN(n7647) );
  NAND2_X1 U7385 ( .A1(n14730), .A2(n14731), .ZN(n14729) );
  AND2_X1 U7386 ( .A1(n14055), .A2(n9645), .ZN(n14048) );
  AND2_X1 U7387 ( .A1(n14743), .A2(n8861), .ZN(n14730) );
  NAND2_X1 U7388 ( .A1(n7796), .A2(n7266), .ZN(n8170) );
  NOR2_X1 U7389 ( .A1(n12709), .A2(n12710), .ZN(n14980) );
  NAND2_X1 U7390 ( .A1(n8404), .A2(n8402), .ZN(n14379) );
  NAND2_X1 U7391 ( .A1(n7469), .A2(n12895), .ZN(n15667) );
  AOI22_X1 U7392 ( .A1(n7838), .A2(n7254), .B1(n12587), .B2(n7832), .ZN(n12706) );
  NAND2_X1 U7393 ( .A1(n12568), .A2(n7214), .ZN(n7867) );
  OAI21_X1 U7394 ( .B1(n9719), .B2(n9718), .A(n9308), .ZN(n9310) );
  AND2_X1 U7395 ( .A1(n8919), .A2(n8918), .ZN(n14925) );
  NAND2_X1 U7396 ( .A1(n9702), .A2(n9701), .ZN(n9704) );
  NAND2_X1 U7397 ( .A1(n8026), .A2(n8025), .ZN(n12663) );
  NAND2_X1 U7398 ( .A1(n7846), .A2(n8401), .ZN(n12495) );
  NAND2_X1 U7399 ( .A1(n7403), .A2(n12358), .ZN(n12480) );
  NAND2_X1 U7400 ( .A1(n9688), .A2(n9687), .ZN(n9690) );
  NAND2_X1 U7401 ( .A1(n12141), .A2(n12140), .ZN(n12331) );
  OR2_X1 U7402 ( .A1(n12069), .A2(n12068), .ZN(n12072) );
  NAND2_X1 U7403 ( .A1(n12043), .A2(n12042), .ZN(n12044) );
  NAND2_X1 U7404 ( .A1(n12825), .A2(n12824), .ZN(n15711) );
  AOI21_X1 U7405 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12306), .A(n12300), .ZN(
        n12450) );
  NOR2_X1 U7406 ( .A1(n11975), .A2(n11974), .ZN(n11976) );
  NOR2_X1 U7407 ( .A1(n11961), .A2(n9534), .ZN(n11974) );
  NAND2_X1 U7408 ( .A1(n11622), .A2(n13259), .ZN(n11621) );
  INV_X1 U7409 ( .A(n7754), .ZN(n11973) );
  NAND2_X1 U7410 ( .A1(n11188), .A2(n8257), .ZN(n11314) );
  AND2_X1 U7411 ( .A1(n11936), .A2(n8742), .ZN(n11895) );
  OAI22_X1 U7412 ( .A1(n11113), .A2(n11112), .B1(n11086), .B2(n11085), .ZN(
        n11090) );
  NAND2_X1 U7413 ( .A1(n11468), .A2(n13260), .ZN(n11467) );
  NAND2_X2 U7414 ( .A1(n12077), .A2(n12076), .ZN(n12797) );
  INV_X1 U7415 ( .A(n11901), .ZN(n16133) );
  AND2_X1 U7416 ( .A1(n11357), .A2(n16095), .ZN(n11348) );
  AND2_X1 U7417 ( .A1(n8734), .A2(n8733), .ZN(n11901) );
  AND2_X1 U7418 ( .A1(n8008), .A2(n8007), .ZN(n9580) );
  OR2_X1 U7419 ( .A1(n9287), .A2(n7342), .ZN(n8008) );
  NAND2_X1 U7420 ( .A1(n7232), .A2(n7442), .ZN(n11018) );
  NOR2_X1 U7421 ( .A1(n10982), .A2(n10981), .ZN(n10984) );
  NAND2_X1 U7422 ( .A1(n7911), .A2(n7910), .ZN(n11594) );
  INV_X2 U7423 ( .A(n16180), .ZN(n16183) );
  NAND4_X2 U7424 ( .A1(n11138), .A2(n11137), .A3(n11136), .A4(n11135), .ZN(
        n15233) );
  NAND4_X1 U7425 ( .A1(n10765), .A2(n10764), .A3(n10763), .A4(n10762), .ZN(
        n15234) );
  NAND2_X1 U7426 ( .A1(n7430), .A2(n7428), .ZN(n9186) );
  OAI21_X1 U7427 ( .B1(n10748), .B2(n12987), .A(n7798), .ZN(n12757) );
  CLKBUF_X1 U7428 ( .A(n10980), .Z(n7718) );
  NAND2_X1 U7429 ( .A1(n8498), .A2(n8497), .ZN(n9094) );
  NAND4_X1 U7430 ( .A1(n9388), .A2(n9386), .A3(n9387), .A4(n9385), .ZN(n13740)
         );
  NAND4_X1 U7431 ( .A1(n9411), .A2(n9410), .A3(n9409), .A4(n9408), .ZN(n13522)
         );
  NAND4_X1 U7432 ( .A1(n9399), .A2(n9398), .A3(n9397), .A4(n9396), .ZN(n13523)
         );
  INV_X2 U7433 ( .A(n8699), .ZN(n9104) );
  AND4_X1 U7434 ( .A1(n10699), .A2(n10698), .A3(n10697), .A4(n10696), .ZN(
        n10864) );
  NAND4_X1 U7435 ( .A1(n8636), .A2(n8635), .A3(n8634), .A4(n8633), .ZN(n14483)
         );
  NAND4_X1 U7436 ( .A1(n8654), .A2(n8653), .A3(n8652), .A4(n8651), .ZN(n14482)
         );
  NAND2_X1 U7437 ( .A1(n11046), .A2(n10406), .ZN(n16151) );
  OAI211_X1 U7438 ( .C1(n10628), .C2(n10431), .A(n9417), .B(n9416), .ZN(n10737) );
  AND2_X1 U7439 ( .A1(n13078), .A2(n15764), .ZN(n10761) );
  AND2_X2 U7440 ( .A1(n8288), .A2(n8287), .ZN(n15062) );
  XNOR2_X1 U7441 ( .A(n8505), .B(n8504), .ZN(n10115) );
  AND2_X4 U7442 ( .A1(n12718), .A2(n8611), .ZN(n8650) );
  INV_X2 U7443 ( .A(n12987), .ZN(n12998) );
  AOI21_X1 U7444 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(n9134), .A(n9133), .ZN(
        n9184) );
  BUF_X2 U7445 ( .A(n10757), .Z(n12965) );
  NOR2_X1 U7446 ( .A1(n9179), .A2(n15938), .ZN(n9181) );
  MUX2_X1 U7447 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15780), .S(n10691), .Z(n10786)
         );
  NAND2_X1 U7448 ( .A1(n8493), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8505) );
  NAND2_X2 U7449 ( .A1(n9360), .A2(n12397), .ZN(n13246) );
  INV_X1 U7450 ( .A(n9360), .ZN(n13320) );
  NAND2_X1 U7451 ( .A1(n8607), .A2(n8608), .ZN(n8609) );
  AND2_X1 U7452 ( .A1(n10379), .A2(n10378), .ZN(n12731) );
  OR2_X1 U7453 ( .A1(n8500), .A2(n8810), .ZN(n7386) );
  MUX2_X1 U7454 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8606), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n8608) );
  NAND2_X1 U7455 ( .A1(n10368), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10219) );
  XNOR2_X1 U7456 ( .A(n10404), .B(P1_IR_REG_19__SCAN_IN), .ZN(n12730) );
  NAND2_X1 U7457 ( .A1(n7683), .A2(n7681), .ZN(n12264) );
  XNOR2_X1 U7458 ( .A(n8210), .B(n10220), .ZN(n15351) );
  INV_X1 U7459 ( .A(n7776), .ZN(n9129) );
  NAND2_X1 U7460 ( .A1(n7939), .A2(n7943), .ZN(n10522) );
  NAND2_X2 U7461 ( .A1(n9343), .A2(P1_U3086), .ZN(n15771) );
  INV_X4 U7462 ( .A(n9343), .ZN(n10689) );
  INV_X1 U7463 ( .A(n10239), .ZN(n8058) );
  CLKBUF_X1 U7464 ( .A(n9400), .Z(n10524) );
  NAND4_X1 U7465 ( .A1(n10190), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10239) );
  NAND2_X1 U7466 ( .A1(n9128), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7777) );
  AND2_X1 U7467 ( .A1(n9400), .A2(n7941), .ZN(n9412) );
  XOR2_X1 U7468 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), .Z(
        n9169) );
  INV_X1 U7469 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n9230) );
  NOR2_X1 U7470 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n10133) );
  NOR2_X1 U7471 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n10134) );
  NOR2_X1 U7472 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n10135) );
  INV_X1 U7473 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n11432) );
  INV_X1 U7474 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n11182) );
  INV_X1 U7475 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9424) );
  INV_X1 U7476 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9075) );
  CLKBUF_X2 U7477 ( .A(P3_IR_REG_0__SCAN_IN), .Z(n7731) );
  INV_X1 U7478 ( .A(P1_RD_REG_SCAN_IN), .ZN(n16000) );
  INV_X1 U7479 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n15348) );
  NOR2_X1 U7480 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8478) );
  INV_X4 U7481 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7482 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n10212) );
  NOR2_X1 U7483 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n9325) );
  XNOR2_X2 U7484 ( .A(n10219), .B(n10218), .ZN(n10290) );
  NOR2_X2 U7485 ( .A1(n15965), .A2(n15964), .ZN(n15963) );
  NOR2_X2 U7486 ( .A1(n7436), .A2(n15959), .ZN(n15965) );
  OAI21_X2 U7487 ( .B1(n9213), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n15970), .ZN(
        n15976) );
  INV_X1 U7488 ( .A(n9335), .ZN(n7421) );
  AND2_X1 U7489 ( .A1(n11118), .A2(n11119), .ZN(n11127) );
  NOR2_X1 U7490 ( .A1(n8282), .A2(n7840), .ZN(n7839) );
  NOR2_X1 U7491 ( .A1(n7841), .A2(n12019), .ZN(n7840) );
  NAND2_X1 U7492 ( .A1(n8205), .A2(n8207), .ZN(n8202) );
  NAND2_X1 U7493 ( .A1(n8201), .A2(n8207), .ZN(n8200) );
  NAND2_X1 U7494 ( .A1(n15667), .A2(n15406), .ZN(n8207) );
  NOR2_X1 U7495 ( .A1(n12602), .A2(n8106), .ZN(n8105) );
  INV_X1 U7496 ( .A(n12519), .ZN(n8106) );
  NAND2_X1 U7497 ( .A1(n7450), .A2(n7453), .ZN(n8943) );
  AOI21_X1 U7498 ( .B1(n7454), .B2(n8563), .A(n7354), .ZN(n7453) );
  OR2_X1 U7499 ( .A1(n8906), .A2(n7451), .ZN(n7450) );
  AOI21_X1 U7500 ( .B1(n7661), .B2(n7663), .A(n7659), .ZN(n7658) );
  INV_X1 U7501 ( .A(n12125), .ZN(n7659) );
  INV_X1 U7502 ( .A(n9605), .ZN(n9778) );
  INV_X1 U7503 ( .A(n7639), .ZN(n7638) );
  INV_X1 U7504 ( .A(n8885), .ZN(n10032) );
  AOI21_X1 U7505 ( .B1(n7578), .B2(n7576), .A(n7284), .ZN(n7575) );
  INV_X1 U7506 ( .A(n14613), .ZN(n7576) );
  NOR2_X1 U7507 ( .A1(n9050), .A2(n8125), .ZN(n8124) );
  INV_X1 U7508 ( .A(n9049), .ZN(n8125) );
  AND2_X1 U7509 ( .A1(n10101), .A2(n9045), .ZN(n7610) );
  AND2_X1 U7510 ( .A1(n11935), .A2(n9038), .ZN(n12141) );
  XNOR2_X1 U7511 ( .A(n11944), .B(n12038), .ZN(n11937) );
  NAND2_X1 U7512 ( .A1(n10980), .A2(n8631), .ZN(n9027) );
  NOR2_X1 U7513 ( .A1(n9094), .A2(n10115), .ZN(n11522) );
  NOR2_X1 U7514 ( .A1(n15586), .A2(n8209), .ZN(n8208) );
  INV_X1 U7515 ( .A(n15396), .ZN(n8209) );
  INV_X1 U7516 ( .A(n7373), .ZN(n9911) );
  NAND2_X1 U7517 ( .A1(n8244), .A2(n8243), .ZN(n8248) );
  INV_X1 U7518 ( .A(n7272), .ZN(n8243) );
  NAND2_X1 U7519 ( .A1(n9929), .A2(n9930), .ZN(n9928) );
  INV_X1 U7520 ( .A(n12810), .ZN(n8306) );
  INV_X1 U7521 ( .A(n9959), .ZN(n9962) );
  INV_X1 U7522 ( .A(n9981), .ZN(n8223) );
  NAND2_X1 U7523 ( .A1(n8216), .A2(n8215), .ZN(n8214) );
  INV_X1 U7524 ( .A(n8217), .ZN(n8215) );
  INV_X1 U7525 ( .A(n8219), .ZN(n8216) );
  NAND2_X1 U7526 ( .A1(n12884), .A2(n12887), .ZN(n7503) );
  OR2_X1 U7527 ( .A1(n9988), .A2(n9985), .ZN(n8465) );
  INV_X1 U7528 ( .A(n8053), .ZN(n8052) );
  OAI21_X1 U7529 ( .B1(n14093), .B2(n8054), .A(n14074), .ZN(n8053) );
  XNOR2_X1 U7530 ( .A(n12991), .B(n12730), .ZN(n12734) );
  INV_X1 U7531 ( .A(n15222), .ZN(n15410) );
  INV_X1 U7532 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U7533 ( .A1(n7560), .A2(n10690), .ZN(n7561) );
  NAND2_X1 U7534 ( .A1(n12547), .A2(n12548), .ZN(n8330) );
  NAND2_X1 U7535 ( .A1(n13467), .A2(n7646), .ZN(n13360) );
  INV_X1 U7536 ( .A(n7765), .ZN(n11099) );
  AND2_X1 U7537 ( .A1(n7261), .A2(n13295), .ZN(n8043) );
  NOR4_X1 U7538 ( .A1(n13094), .A2(n13938), .A3(n13961), .A4(n13093), .ZN(
        n13256) );
  NAND2_X1 U7539 ( .A1(n11018), .A2(n11017), .ZN(n7757) );
  NAND2_X1 U7540 ( .A1(n7699), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7796) );
  INV_X1 U7541 ( .A(n7632), .ZN(n7631) );
  OAI21_X1 U7542 ( .B1(n8030), .B2(n13938), .A(n13205), .ZN(n7632) );
  NAND2_X1 U7543 ( .A1(n13369), .A2(n13953), .ZN(n13204) );
  NAND2_X1 U7544 ( .A1(n14227), .A2(n14001), .ZN(n8441) );
  OR2_X1 U7545 ( .A1(n16223), .A2(n14089), .ZN(n13157) );
  NAND2_X1 U7546 ( .A1(n12480), .A2(n12551), .ZN(n9561) );
  OR2_X1 U7547 ( .A1(n13522), .A2(n10737), .ZN(n13107) );
  OAI21_X1 U7548 ( .B1(n9812), .B2(n14047), .A(n7616), .ZN(n14035) );
  INV_X1 U7549 ( .A(n7617), .ZN(n7616) );
  OAI21_X1 U7550 ( .B1(n14047), .B2(n13173), .A(n13175), .ZN(n7617) );
  NOR2_X1 U7551 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n8056) );
  XNOR2_X1 U7552 ( .A(n9341), .B(n9340), .ZN(n9342) );
  NOR2_X1 U7553 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n9333) );
  NOR2_X1 U7554 ( .A1(n9616), .A2(n9329), .ZN(n7420) );
  INV_X1 U7555 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9328) );
  AND2_X1 U7556 ( .A1(n9546), .A2(n9545), .ZN(n9549) );
  NAND2_X1 U7557 ( .A1(n7446), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7943) );
  OAI21_X1 U7558 ( .B1(n10524), .B2(n7942), .A(n7940), .ZN(n7939) );
  AND2_X1 U7559 ( .A1(n7941), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U7560 ( .A1(n10524), .A2(n7941), .ZN(n7940) );
  NAND2_X1 U7561 ( .A1(n8368), .A2(n8369), .ZN(n14576) );
  INV_X1 U7562 ( .A(n14929), .ZN(n9051) );
  NOR2_X1 U7563 ( .A1(n10110), .A2(n7207), .ZN(n7695) );
  NAND2_X1 U7564 ( .A1(n10109), .A2(n8370), .ZN(n8369) );
  INV_X1 U7565 ( .A(n8371), .ZN(n8370) );
  AOI21_X1 U7566 ( .B1(n8154), .B2(n14594), .A(n8372), .ZN(n8371) );
  INV_X1 U7567 ( .A(n14577), .ZN(n8372) );
  NAND2_X1 U7568 ( .A1(n14351), .A2(n7591), .ZN(n7590) );
  INV_X1 U7569 ( .A(n7714), .ZN(n7591) );
  NAND2_X1 U7570 ( .A1(n14778), .A2(n8834), .ZN(n14756) );
  INV_X1 U7571 ( .A(n8656), .ZN(n8699) );
  AND2_X1 U7572 ( .A1(n7615), .A2(n8414), .ZN(n7612) );
  NAND2_X1 U7573 ( .A1(n7727), .A2(n8486), .ZN(n7614) );
  NOR2_X1 U7574 ( .A1(n8585), .A2(n8484), .ZN(n8500) );
  AND2_X1 U7575 ( .A1(n15189), .A2(n8272), .ZN(n8271) );
  NAND2_X1 U7576 ( .A1(n15142), .A2(n8273), .ZN(n8272) );
  INV_X1 U7577 ( .A(n15054), .ZN(n8279) );
  NAND2_X1 U7578 ( .A1(n16096), .A2(n15062), .ZN(n15094) );
  NAND2_X1 U7579 ( .A1(n15481), .A2(n15487), .ZN(n15480) );
  INV_X1 U7580 ( .A(n12073), .ZN(n8072) );
  NOR2_X1 U7581 ( .A1(n8182), .A2(n12767), .ZN(n8178) );
  AND2_X1 U7582 ( .A1(n7198), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n8080) );
  OAI21_X1 U7583 ( .B1(n7198), .B2(n8082), .A(n8077), .ZN(n8076) );
  NAND2_X1 U7584 ( .A1(n8078), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n8077) );
  OAI21_X1 U7585 ( .B1(n8574), .B2(n7902), .A(n7900), .ZN(n9000) );
  INV_X1 U7586 ( .A(n7901), .ZN(n7900) );
  OAI21_X1 U7587 ( .B1(n7903), .B2(n7902), .A(n8580), .ZN(n7901) );
  INV_X1 U7588 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10140) );
  INV_X1 U7589 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U7590 ( .A1(n8570), .A2(n8569), .ZN(n8961) );
  NAND2_X1 U7591 ( .A1(n8943), .A2(n8566), .ZN(n8570) );
  NAND2_X1 U7592 ( .A1(n7889), .A2(n7886), .ZN(n8906) );
  AOI21_X1 U7593 ( .B1(n7888), .B2(n7887), .A(n7339), .ZN(n7886) );
  XNOR2_X1 U7594 ( .A(n8554), .B(n13659), .ZN(n8835) );
  NAND2_X1 U7595 ( .A1(n7876), .A2(n7462), .ZN(n7461) );
  INV_X1 U7596 ( .A(n8822), .ZN(n7462) );
  NAND2_X1 U7597 ( .A1(n8762), .A2(n8761), .ZN(n8764) );
  NAND2_X1 U7598 ( .A1(n8392), .A2(SI_3_), .ZN(n8523) );
  NAND2_X1 U7599 ( .A1(n7791), .A2(n7790), .ZN(n8356) );
  INV_X1 U7600 ( .A(n13359), .ZN(n7790) );
  INV_X1 U7601 ( .A(n13360), .ZN(n7791) );
  OAI21_X1 U7602 ( .B1(n13493), .B2(n7233), .A(n7667), .ZN(n13442) );
  INV_X1 U7603 ( .A(n7668), .ZN(n7667) );
  OAI21_X1 U7604 ( .B1(n7233), .B2(n13337), .A(n13340), .ZN(n7668) );
  AND2_X1 U7605 ( .A1(n13425), .A2(n13363), .ZN(n13450) );
  NAND2_X1 U7606 ( .A1(n13360), .A2(n13359), .ZN(n13449) );
  XNOR2_X1 U7607 ( .A(n10737), .B(n11099), .ZN(n11098) );
  NAND2_X1 U7608 ( .A1(n7306), .A2(n8338), .ZN(n7661) );
  NAND2_X1 U7609 ( .A1(n11927), .A2(n7666), .ZN(n7665) );
  AND2_X1 U7610 ( .A1(n8340), .A2(n8339), .ZN(n11928) );
  NAND2_X1 U7611 ( .A1(n11793), .A2(n13519), .ZN(n8339) );
  XNOR2_X1 U7612 ( .A(n16029), .B(n11099), .ZN(n10736) );
  NAND2_X1 U7613 ( .A1(n7669), .A2(n7708), .ZN(n7793) );
  INV_X1 U7614 ( .A(n10641), .ZN(n7708) );
  OR2_X1 U7615 ( .A1(n11653), .A2(n11654), .ZN(n8340) );
  INV_X1 U7616 ( .A(n13426), .ZN(n8337) );
  AOI21_X1 U7617 ( .B1(n13426), .B2(n8336), .A(n8335), .ZN(n8334) );
  INV_X1 U7618 ( .A(n13368), .ZN(n8335) );
  OR2_X1 U7619 ( .A1(n14249), .A2(n10132), .ZN(n10462) );
  NAND2_X1 U7620 ( .A1(n10956), .A2(n9851), .ZN(n13293) );
  NAND2_X2 U7621 ( .A1(n9361), .A2(n9360), .ZN(n9605) );
  AND2_X1 U7622 ( .A1(n10520), .A2(n10519), .ZN(n7745) );
  NOR2_X1 U7623 ( .A1(n11014), .A2(n16146), .ZN(n11559) );
  NAND2_X1 U7624 ( .A1(n8165), .A2(n8164), .ZN(n13792) );
  INV_X1 U7625 ( .A(n12455), .ZN(n8164) );
  NAND2_X1 U7626 ( .A1(n8170), .A2(n8169), .ZN(n8168) );
  INV_X1 U7627 ( .A(n13824), .ZN(n8169) );
  AOI21_X1 U7628 ( .B1(n13868), .B2(n7741), .A(n13867), .ZN(n13871) );
  NOR2_X1 U7629 ( .A1(n13871), .A2(n13870), .ZN(n7447) );
  NAND2_X1 U7630 ( .A1(n9814), .A2(n13218), .ZN(n13915) );
  AND2_X1 U7631 ( .A1(n8033), .A2(n13952), .ZN(n8031) );
  INV_X1 U7632 ( .A(n13974), .ZN(n13979) );
  NOR2_X1 U7633 ( .A1(n13999), .A2(n7637), .ZN(n7636) );
  INV_X1 U7634 ( .A(n13189), .ZN(n7637) );
  OR2_X1 U7635 ( .A1(n14227), .A2(n14029), .ZN(n13189) );
  INV_X1 U7636 ( .A(n14074), .ZN(n8458) );
  NAND2_X1 U7637 ( .A1(n11619), .A2(n13126), .ZN(n12101) );
  AND2_X1 U7638 ( .A1(n13096), .A2(n7643), .ZN(n16028) );
  NAND2_X1 U7639 ( .A1(n13098), .A2(n11648), .ZN(n7643) );
  OR2_X1 U7640 ( .A1(n13740), .A2(n11064), .ZN(n11648) );
  INV_X1 U7641 ( .A(n9705), .ZN(n13241) );
  INV_X1 U7642 ( .A(n9443), .ZN(n9668) );
  INV_X1 U7643 ( .A(n10431), .ZN(n9667) );
  INV_X1 U7644 ( .A(n10462), .ZN(n10466) );
  NAND2_X1 U7645 ( .A1(n10956), .A2(n9820), .ZN(n16222) );
  INV_X1 U7646 ( .A(n7986), .ZN(n7985) );
  OAI21_X1 U7647 ( .B1(n9661), .B2(n7987), .A(n9676), .ZN(n7986) );
  XNOR2_X1 U7648 ( .A(n9666), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13881) );
  INV_X1 U7649 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n9545) );
  OAI21_X1 U7650 ( .B1(n9274), .B2(n8004), .A(n8002), .ZN(n9491) );
  INV_X1 U7651 ( .A(n8003), .ZN(n8002) );
  OAI21_X1 U7652 ( .B1(n8005), .B2(n8004), .A(n9488), .ZN(n8003) );
  INV_X1 U7653 ( .A(n9276), .ZN(n8004) );
  AND4_X1 U7654 ( .A1(n9322), .A2(n9455), .A3(n9424), .A4(n9457), .ZN(n9323)
         );
  NOR2_X1 U7655 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n9322) );
  NAND2_X1 U7656 ( .A1(n9274), .A2(n8005), .ZN(n9474) );
  AOI21_X1 U7657 ( .B1(n7999), .B2(n8001), .A(n7997), .ZN(n7996) );
  INV_X1 U7658 ( .A(n9271), .ZN(n7997) );
  NAND2_X1 U7659 ( .A1(n9064), .A2(n13321), .ZN(n8629) );
  OR2_X1 U7660 ( .A1(n12496), .A2(n12498), .ZN(n12568) );
  AND3_X1 U7661 ( .A1(n8925), .A2(n8924), .A3(n8923), .ZN(n14289) );
  AND3_X1 U7662 ( .A1(n8913), .A2(n8912), .A3(n8911), .ZN(n14361) );
  NAND2_X1 U7663 ( .A1(n7574), .A2(n7573), .ZN(n14585) );
  AOI21_X1 U7664 ( .B1(n7575), .B2(n7577), .A(n10109), .ZN(n7573) );
  OR2_X1 U7665 ( .A1(n14618), .A2(n14601), .ZN(n14603) );
  NAND2_X1 U7666 ( .A1(n9053), .A2(n8972), .ZN(n14613) );
  NOR2_X1 U7667 ( .A1(n7270), .A2(n7598), .ZN(n7596) );
  NAND2_X1 U7668 ( .A1(n14728), .A2(n9048), .ZN(n9049) );
  NAND2_X1 U7669 ( .A1(n14729), .A2(n8874), .ZN(n14708) );
  AND2_X1 U7670 ( .A1(n14879), .A2(n14774), .ZN(n14763) );
  NAND2_X1 U7671 ( .A1(n14771), .A2(n9044), .ZN(n7611) );
  NAND2_X1 U7672 ( .A1(n12401), .A2(n16202), .ZN(n14801) );
  NAND2_X1 U7673 ( .A1(n12325), .A2(n8794), .ZN(n12406) );
  INV_X1 U7674 ( .A(n12329), .ZN(n12326) );
  NAND2_X1 U7675 ( .A1(n8760), .A2(n7269), .ZN(n8149) );
  NAND2_X1 U7676 ( .A1(n11934), .A2(n11937), .ZN(n8760) );
  NAND2_X1 U7677 ( .A1(n7694), .A2(n9037), .ZN(n11935) );
  AOI21_X1 U7678 ( .B1(n7236), .B2(n9036), .A(n8134), .ZN(n8133) );
  OAI21_X1 U7679 ( .B1(n7583), .B2(n10096), .A(n7581), .ZN(n11892) );
  AOI21_X1 U7680 ( .B1(n11661), .B2(n7582), .A(n7268), .ZN(n7581) );
  INV_X1 U7681 ( .A(n7767), .ZN(n7582) );
  OR2_X1 U7682 ( .A1(n11416), .A2(n8702), .ZN(n7584) );
  OAI211_X1 U7683 ( .C1(n8131), .C2(n11393), .A(n8130), .B(n11407), .ZN(n11406) );
  AND2_X1 U7684 ( .A1(n8629), .A2(n9343), .ZN(n8656) );
  INV_X1 U7685 ( .A(n14719), .ZN(n9112) );
  AND3_X1 U7686 ( .A1(n7609), .A2(n7607), .A3(n7606), .ZN(n9109) );
  INV_X1 U7687 ( .A(n14351), .ZN(n7606) );
  INV_X1 U7688 ( .A(n7590), .ZN(n7588) );
  OR2_X1 U7689 ( .A1(n11508), .A2(n14479), .ZN(n7767) );
  XNOR2_X1 U7690 ( .A(n8605), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U7691 ( .A1(n8607), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U7692 ( .A1(n8485), .A2(n8471), .ZN(n8489) );
  NOR2_X1 U7693 ( .A1(n8482), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7385) );
  XNOR2_X1 U7694 ( .A(n10843), .B(n15065), .ZN(n11118) );
  OAI21_X1 U7695 ( .B1(n7237), .B2(n15100), .A(n7824), .ZN(n7823) );
  NAND2_X1 U7696 ( .A1(n7237), .A2(n7825), .ZN(n7824) );
  OR2_X1 U7697 ( .A1(n15100), .A2(n15092), .ZN(n7825) );
  AOI21_X1 U7698 ( .B1(n8253), .B2(n8256), .A(n8251), .ZN(n8250) );
  INV_X1 U7699 ( .A(n15150), .ZN(n8251) );
  AOI21_X1 U7700 ( .B1(n7839), .B2(n7841), .A(n7837), .ZN(n7836) );
  AOI21_X1 U7701 ( .B1(n8283), .B2(n8281), .A(n7263), .ZN(n8280) );
  AND2_X1 U7702 ( .A1(n10371), .A2(n15764), .ZN(n10756) );
  AND2_X1 U7703 ( .A1(n10371), .A2(n10372), .ZN(n10757) );
  OR2_X1 U7704 ( .A1(n15451), .A2(n7477), .ZN(n8090) );
  AND2_X1 U7705 ( .A1(n15459), .A2(n15409), .ZN(n7477) );
  NAND2_X1 U7706 ( .A1(n12963), .A2(n12962), .ZN(n15634) );
  NAND2_X1 U7707 ( .A1(n15468), .A2(n8468), .ZN(n15451) );
  OR2_X1 U7708 ( .A1(n15470), .A2(n15378), .ZN(n8468) );
  NOR2_X1 U7709 ( .A1(n15662), .A2(n8118), .ZN(n8117) );
  NAND2_X1 U7710 ( .A1(n15499), .A2(n8113), .ZN(n8110) );
  NAND2_X1 U7711 ( .A1(n8116), .A2(n15509), .ZN(n8115) );
  INV_X1 U7712 ( .A(n15499), .ZN(n8116) );
  AOI21_X1 U7713 ( .B1(n15533), .B2(n15404), .A(n15403), .ZN(n15523) );
  NAND2_X1 U7714 ( .A1(n15534), .A2(n15375), .ZN(n15516) );
  OR2_X1 U7715 ( .A1(n15679), .A2(n15374), .ZN(n15375) );
  XNOR2_X1 U7716 ( .A(n15705), .B(n15369), .ZN(n15586) );
  AND2_X1 U7717 ( .A1(n15603), .A2(n15394), .ZN(n7549) );
  NAND2_X1 U7718 ( .A1(n15366), .A2(n15365), .ZN(n15604) );
  AOI21_X1 U7719 ( .B1(n8105), .B2(n13027), .A(n7259), .ZN(n8103) );
  NOR2_X1 U7720 ( .A1(n13028), .A2(n7548), .ZN(n7547) );
  INV_X1 U7721 ( .A(n12524), .ZN(n7548) );
  NAND2_X1 U7722 ( .A1(n10023), .A2(n10021), .ZN(n10040) );
  AOI21_X1 U7723 ( .B1(n10019), .B2(n10018), .A(n7230), .ZN(n10023) );
  NAND2_X1 U7724 ( .A1(n7246), .A2(n15943), .ZN(n7428) );
  NAND2_X1 U7725 ( .A1(n7966), .A2(n7235), .ZN(n7430) );
  AND4_X1 U7726 ( .A1(n9659), .A2(n9658), .A3(n9657), .A4(n9656), .ZN(n14028)
         );
  NAND2_X1 U7727 ( .A1(n8237), .A2(n10123), .ZN(n8236) );
  NAND2_X1 U7728 ( .A1(n10113), .A2(n10114), .ZN(n8237) );
  OR2_X1 U7729 ( .A1(n14567), .A2(n9058), .ZN(n8616) );
  NAND2_X1 U7730 ( .A1(n8138), .A2(n7704), .ZN(n7703) );
  INV_X1 U7731 ( .A(n9240), .ZN(n7704) );
  NAND2_X1 U7732 ( .A1(n15123), .A2(n8277), .ZN(n8275) );
  NAND2_X1 U7733 ( .A1(n10308), .A2(n10307), .ZN(n10312) );
  NOR2_X1 U7734 ( .A1(n15988), .A2(n15989), .ZN(n15987) );
  OR2_X1 U7735 ( .A1(n9882), .A2(n11399), .ZN(n9883) );
  NAND2_X1 U7736 ( .A1(n9891), .A2(n9890), .ZN(n9904) );
  AND2_X1 U7737 ( .A1(n12748), .A2(n8462), .ZN(n7762) );
  NAND2_X1 U7738 ( .A1(n9902), .A2(n9901), .ZN(n7373) );
  NAND2_X1 U7739 ( .A1(n12773), .A2(n12772), .ZN(n7498) );
  AOI21_X1 U7740 ( .B1(n7377), .B2(n9917), .A(n9916), .ZN(n9919) );
  NAND2_X1 U7741 ( .A1(n9923), .A2(n7272), .ZN(n8249) );
  INV_X1 U7742 ( .A(n9925), .ZN(n7366) );
  NOR2_X1 U7743 ( .A1(n12781), .A2(n12784), .ZN(n7509) );
  NAND2_X1 U7744 ( .A1(n12778), .A2(n8291), .ZN(n8290) );
  INV_X1 U7745 ( .A(n12779), .ZN(n8291) );
  NAND2_X1 U7746 ( .A1(n12784), .A2(n12781), .ZN(n7508) );
  NOR2_X1 U7747 ( .A1(n12812), .A2(n12810), .ZN(n8307) );
  INV_X1 U7748 ( .A(n8307), .ZN(n8305) );
  OAI22_X1 U7749 ( .A1(n12807), .A2(n7530), .B1(n7529), .B2(n12808), .ZN(n7528) );
  INV_X1 U7750 ( .A(n12806), .ZN(n7529) );
  NOR2_X1 U7751 ( .A1(n12809), .A2(n12806), .ZN(n7530) );
  AOI21_X1 U7752 ( .B1(n8303), .B2(n12814), .A(n8302), .ZN(n8301) );
  INV_X1 U7753 ( .A(n12813), .ZN(n8302) );
  NOR2_X1 U7754 ( .A1(n8303), .A2(n12814), .ZN(n8300) );
  NAND2_X1 U7755 ( .A1(n9954), .A2(n9953), .ZN(n7376) );
  NAND2_X1 U7756 ( .A1(n9952), .A2(n9951), .ZN(n7375) );
  NAND2_X1 U7757 ( .A1(n8240), .A2(n9955), .ZN(n8239) );
  INV_X1 U7758 ( .A(n9957), .ZN(n8240) );
  NAND2_X1 U7759 ( .A1(n12826), .A2(n12828), .ZN(n8293) );
  INV_X1 U7760 ( .A(n12874), .ZN(n8314) );
  AND2_X1 U7761 ( .A1(n8220), .A2(n9982), .ZN(n8219) );
  NAND2_X1 U7762 ( .A1(n8224), .A2(n8221), .ZN(n8220) );
  NOR2_X1 U7763 ( .A1(n8221), .A2(n8224), .ZN(n8217) );
  NAND2_X1 U7764 ( .A1(n8224), .A2(n7275), .ZN(n8222) );
  NAND2_X1 U7765 ( .A1(n8313), .A2(n12874), .ZN(n8312) );
  NAND2_X1 U7766 ( .A1(n7516), .A2(n7517), .ZN(n7760) );
  INV_X1 U7767 ( .A(n12873), .ZN(n8313) );
  INV_X1 U7768 ( .A(n12884), .ZN(n7504) );
  NAND2_X1 U7769 ( .A1(n12900), .A2(n12899), .ZN(n7535) );
  AOI21_X1 U7770 ( .B1(n8226), .B2(n9994), .A(n7369), .ZN(n7368) );
  INV_X1 U7771 ( .A(n9993), .ZN(n7369) );
  NAND2_X1 U7772 ( .A1(n12922), .A2(n12920), .ZN(n8310) );
  NAND2_X1 U7773 ( .A1(n7513), .A2(n12931), .ZN(n7512) );
  AND2_X1 U7774 ( .A1(n12933), .A2(n7515), .ZN(n7514) );
  INV_X1 U7775 ( .A(n12931), .ZN(n7515) );
  NAND2_X1 U7776 ( .A1(n7650), .A2(n7653), .ZN(n7649) );
  AND2_X1 U7777 ( .A1(n13354), .A2(n13351), .ZN(n8359) );
  NAND2_X1 U7778 ( .A1(n13214), .A2(n13229), .ZN(n7398) );
  OR2_X1 U7779 ( .A1(n13256), .A2(n8014), .ZN(n7396) );
  OR2_X1 U7780 ( .A1(n13213), .A2(n13229), .ZN(n8014) );
  AOI21_X1 U7781 ( .B1(n13256), .B2(n13215), .A(n13915), .ZN(n7397) );
  NAND2_X1 U7782 ( .A1(n7348), .A2(n8578), .ZN(n7902) );
  AND2_X1 U7783 ( .A1(n7463), .A2(n7344), .ZN(n7872) );
  OAI21_X1 U7784 ( .B1(n7875), .B2(n7460), .A(n7458), .ZN(n7463) );
  AOI21_X1 U7785 ( .B1(n7461), .B2(n8553), .A(n7459), .ZN(n7458) );
  OR2_X1 U7786 ( .A1(n7210), .A2(n8745), .ZN(n8377) );
  OR2_X1 U7787 ( .A1(n8539), .A2(n8381), .ZN(n8376) );
  INV_X1 U7788 ( .A(n8535), .ZN(n7471) );
  INV_X1 U7789 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9130) );
  INV_X1 U7790 ( .A(n12621), .ZN(n8329) );
  NOR2_X1 U7791 ( .A1(n13230), .A2(n8048), .ZN(n8047) );
  INV_X1 U7792 ( .A(n7943), .ZN(n7938) );
  NOR2_X2 U7793 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n9400) );
  NAND2_X1 U7794 ( .A1(n8158), .A2(n10544), .ZN(n8159) );
  AND2_X1 U7795 ( .A1(n10628), .A2(n10528), .ZN(n8158) );
  AND3_X1 U7796 ( .A1(n8162), .A2(n8161), .A3(n7265), .ZN(n10802) );
  NOR2_X1 U7797 ( .A1(n9552), .A2(n14190), .ZN(n7926) );
  NAND2_X1 U7798 ( .A1(n13792), .A2(n13791), .ZN(n7782) );
  NAND2_X1 U7799 ( .A1(n13844), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8167) );
  INV_X1 U7800 ( .A(n8453), .ZN(n13916) );
  AOI21_X1 U7801 ( .B1(n8447), .B2(n9754), .A(n7297), .ZN(n8445) );
  INV_X1 U7802 ( .A(n8447), .ZN(n8446) );
  INV_X1 U7803 ( .A(n8455), .ZN(n8451) );
  NAND2_X1 U7804 ( .A1(n13369), .A2(n13510), .ZN(n8454) );
  OR2_X1 U7805 ( .A1(n14155), .A2(n13469), .ZN(n13352) );
  OR2_X1 U7806 ( .A1(n14039), .A2(n13462), .ZN(n13184) );
  OR2_X1 U7807 ( .A1(n14169), .A2(n14028), .ZN(n13177) );
  INV_X1 U7808 ( .A(n16031), .ZN(n13270) );
  NOR2_X1 U7809 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n8460) );
  INV_X1 U7810 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n9785) );
  NOR2_X1 U7811 ( .A1(n9634), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n9786) );
  INV_X1 U7812 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U7813 ( .A1(n9544), .A2(n9286), .ZN(n9287) );
  INV_X1 U7814 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9486) );
  NOR2_X1 U7815 ( .A1(n9471), .A2(n8006), .ZN(n8005) );
  INV_X1 U7816 ( .A(n9273), .ZN(n8006) );
  INV_X1 U7817 ( .A(n14334), .ZN(n7849) );
  INV_X1 U7818 ( .A(n14413), .ZN(n14285) );
  NOR2_X1 U7819 ( .A1(n10112), .A2(n7909), .ZN(n7908) );
  AND2_X1 U7820 ( .A1(n10072), .A2(n10071), .ZN(n10082) );
  NAND2_X1 U7821 ( .A1(n9122), .A2(n7915), .ZN(n7914) );
  NOR2_X1 U7822 ( .A1(n14560), .A2(n14569), .ZN(n7915) );
  NOR2_X1 U7823 ( .A1(n8154), .A2(n7579), .ZN(n7578) );
  INV_X1 U7824 ( .A(n8973), .ZN(n7579) );
  AND2_X1 U7825 ( .A1(n10109), .A2(n8154), .ZN(n8362) );
  NOR2_X1 U7826 ( .A1(n10974), .A2(n8503), .ZN(n11230) );
  OR2_X1 U7827 ( .A1(n9067), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9079) );
  INV_X1 U7828 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8416) );
  INV_X1 U7829 ( .A(n7807), .ZN(n7815) );
  OAI21_X1 U7830 ( .B1(n11312), .B2(n11313), .A(n7249), .ZN(n7807) );
  INV_X1 U7831 ( .A(n15031), .ZN(n8255) );
  INV_X1 U7832 ( .A(n7816), .ZN(n7812) );
  INV_X1 U7833 ( .A(n15455), .ZN(n8192) );
  OAI22_X1 U7834 ( .A1(n15455), .A2(n15407), .B1(n15409), .B2(n15648), .ZN(
        n8191) );
  NOR2_X1 U7835 ( .A1(n15459), .A2(n8020), .ZN(n8019) );
  OR2_X1 U7836 ( .A1(n15654), .A2(n15662), .ZN(n8020) );
  NOR2_X1 U7837 ( .A1(n8114), .A2(n15487), .ZN(n8113) );
  INV_X1 U7838 ( .A(n8464), .ZN(n8114) );
  NOR2_X1 U7839 ( .A1(n15552), .A2(n15679), .ZN(n8027) );
  NOR2_X1 U7840 ( .A1(n8102), .A2(n12658), .ZN(n8101) );
  INV_X1 U7841 ( .A(n8103), .ZN(n8102) );
  INV_X1 U7842 ( .A(n12088), .ZN(n7544) );
  OAI21_X1 U7843 ( .B1(n8073), .B2(n8072), .A(n12182), .ZN(n8071) );
  AND2_X1 U7844 ( .A1(n13023), .A2(n12071), .ZN(n8073) );
  AOI21_X1 U7845 ( .B1(n8062), .B2(n8065), .A(n7282), .ZN(n8060) );
  OR2_X1 U7846 ( .A1(n9009), .A2(n9008), .ZN(n9103) );
  INV_X1 U7847 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10149) );
  INV_X1 U7848 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10148) );
  INV_X1 U7849 ( .A(SI_22_), .ZN(n13652) );
  NAND2_X1 U7850 ( .A1(n11612), .A2(n7523), .ZN(n10214) );
  NOR2_X1 U7851 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n7523) );
  OAI22_X1 U7852 ( .A1(n8863), .A2(n8862), .B1(SI_17_), .B2(n8557), .ZN(n8558)
         );
  NAND2_X1 U7853 ( .A1(n8851), .A2(n8556), .ZN(n8863) );
  XNOR2_X1 U7854 ( .A(n8557), .B(SI_17_), .ZN(n8862) );
  NAND2_X1 U7855 ( .A1(n7361), .A2(n13629), .ZN(n8373) );
  INV_X1 U7856 ( .A(n7872), .ZN(n7361) );
  INV_X1 U7857 ( .A(n8553), .ZN(n7460) );
  AND2_X1 U7858 ( .A1(n7363), .A2(n8550), .ZN(n7876) );
  NAND2_X1 U7859 ( .A1(n7877), .A2(n7883), .ZN(n7363) );
  AOI21_X1 U7860 ( .B1(n7884), .B2(n7882), .A(n7299), .ZN(n7881) );
  INV_X1 U7861 ( .A(n8546), .ZN(n7882) );
  AOI21_X1 U7862 ( .B1(n8780), .B2(n8546), .A(n7885), .ZN(n7884) );
  INV_X1 U7863 ( .A(n8795), .ZN(n7885) );
  NAND2_X1 U7864 ( .A1(n8764), .A2(n8543), .ZN(n8781) );
  NAND2_X1 U7865 ( .A1(n8730), .A2(n8538), .ZN(n8540) );
  NAND2_X1 U7866 ( .A1(n8360), .A2(n8532), .ZN(n7897) );
  OAI21_X1 U7867 ( .B1(n8690), .B2(n8361), .A(n8531), .ZN(n8360) );
  INV_X1 U7868 ( .A(n8510), .ZN(n8518) );
  INV_X1 U7869 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7845) );
  NOR2_X1 U7870 ( .A1(n9142), .A2(n9141), .ZN(n9196) );
  NOR2_X1 U7871 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9193), .ZN(n9141) );
  AOI22_X1 U7872 ( .A1(n9203), .A2(n9150), .B1(P1_ADDR_REG_11__SCAN_IN), .B2(
        n9149), .ZN(n9206) );
  NAND2_X1 U7873 ( .A1(n13407), .A2(n13403), .ZN(n8352) );
  NAND2_X1 U7874 ( .A1(n11926), .A2(n13518), .ZN(n7666) );
  INV_X1 U7875 ( .A(n12549), .ZN(n8326) );
  NAND2_X1 U7876 ( .A1(n11300), .A2(n11301), .ZN(n11652) );
  NAND2_X1 U7877 ( .A1(n7654), .A2(n7658), .ZN(n12241) );
  OR2_X1 U7878 ( .A1(n11928), .A2(n7660), .ZN(n7654) );
  INV_X1 U7879 ( .A(n13348), .ZN(n7653) );
  AND2_X1 U7880 ( .A1(n13459), .A2(n7651), .ZN(n7650) );
  NAND2_X1 U7881 ( .A1(n7652), .A2(n13348), .ZN(n7651) );
  INV_X1 U7882 ( .A(n13397), .ZN(n7652) );
  NAND2_X1 U7883 ( .A1(n8329), .A2(n8325), .ZN(n8321) );
  NAND2_X1 U7884 ( .A1(n8320), .A2(n8329), .ZN(n8319) );
  INV_X1 U7885 ( .A(n8323), .ZN(n8320) );
  AOI21_X1 U7886 ( .B1(n8325), .B2(n8328), .A(n8324), .ZN(n8323) );
  NAND2_X1 U7887 ( .A1(n13358), .A2(n13357), .ZN(n7646) );
  NAND2_X1 U7888 ( .A1(n11652), .A2(n7794), .ZN(n11653) );
  NAND2_X1 U7889 ( .A1(n11651), .A2(n7795), .ZN(n7794) );
  NAND2_X1 U7890 ( .A1(n7673), .A2(n13450), .ZN(n13424) );
  NAND2_X1 U7891 ( .A1(n8334), .A2(n8337), .ZN(n8332) );
  NAND2_X1 U7892 ( .A1(n13334), .A2(n13333), .ZN(n13493) );
  AND2_X1 U7893 ( .A1(n13251), .A2(n13250), .ZN(n13902) );
  AND4_X1 U7894 ( .A1(n9577), .A2(n9576), .A3(n9575), .A4(n9574), .ZN(n13384)
         );
  OAI21_X1 U7895 ( .B1(n10498), .B2(n7406), .A(n7404), .ZN(n10509) );
  INV_X1 U7896 ( .A(n7405), .ZN(n7404) );
  OAI21_X1 U7897 ( .B1(n10614), .B2(n7406), .A(n13742), .ZN(n7405) );
  OAI21_X1 U7898 ( .B1(n7435), .B2(n7434), .A(n7432), .ZN(n13772) );
  INV_X1 U7899 ( .A(n7433), .ZN(n7432) );
  OAI21_X1 U7900 ( .B1(n13746), .B2(n7434), .A(n10539), .ZN(n7433) );
  INV_X1 U7901 ( .A(n7780), .ZN(n7434) );
  AOI21_X1 U7902 ( .B1(n13780), .B2(n7949), .A(n7946), .ZN(n7945) );
  NAND2_X1 U7903 ( .A1(n7947), .A2(n7951), .ZN(n7946) );
  NAND2_X1 U7904 ( .A1(n10813), .A2(n10812), .ZN(n10815) );
  NAND2_X1 U7905 ( .A1(n13779), .A2(n7956), .ZN(n7955) );
  OR2_X1 U7906 ( .A1(n11559), .A2(n11560), .ZN(n7921) );
  NAND2_X1 U7907 ( .A1(n7921), .A2(n7920), .ZN(n11950) );
  INV_X1 U7908 ( .A(n11564), .ZN(n7920) );
  OAI21_X1 U7909 ( .B1(n11567), .B2(n11566), .A(n11568), .ZN(n11570) );
  OR2_X1 U7910 ( .A1(n11576), .A2(n11577), .ZN(n8173) );
  INV_X1 U7911 ( .A(n7757), .ZN(n11574) );
  NAND2_X1 U7912 ( .A1(n11950), .A2(n11949), .ZN(n7732) );
  XNOR2_X1 U7913 ( .A(n7754), .B(n11965), .ZN(n11961) );
  XNOR2_X1 U7914 ( .A(n7925), .B(n12311), .ZN(n12303) );
  NAND2_X1 U7915 ( .A1(n12310), .A2(n7411), .ZN(n12469) );
  AND2_X1 U7916 ( .A1(n7412), .A2(n12309), .ZN(n7411) );
  OR2_X1 U7917 ( .A1(n12462), .A2(n12461), .ZN(n13789) );
  XNOR2_X1 U7918 ( .A(n7782), .B(n7449), .ZN(n7699) );
  INV_X1 U7919 ( .A(n7796), .ZN(n13821) );
  NOR2_X1 U7920 ( .A1(n13836), .A2(n14063), .ZN(n13867) );
  NAND2_X1 U7921 ( .A1(n9814), .A2(n13207), .ZN(n8048) );
  NAND2_X1 U7922 ( .A1(n13406), .A2(n8050), .ZN(n8049) );
  INV_X1 U7923 ( .A(n7633), .ZN(n7629) );
  NAND2_X1 U7924 ( .A1(n8012), .A2(n8011), .ZN(n13207) );
  OR2_X1 U7925 ( .A1(n7631), .A2(n13094), .ZN(n7627) );
  INV_X1 U7926 ( .A(n13980), .ZN(n7635) );
  NOR2_X1 U7927 ( .A1(n8450), .A2(n13930), .ZN(n8447) );
  AOI21_X1 U7928 ( .B1(n8031), .B2(n8034), .A(n7220), .ZN(n8030) );
  NAND2_X1 U7929 ( .A1(n8036), .A2(n7288), .ZN(n8033) );
  NAND2_X1 U7930 ( .A1(n8036), .A2(n13200), .ZN(n8034) );
  NAND2_X1 U7931 ( .A1(n13944), .A2(n9778), .ZN(n7387) );
  AOI21_X1 U7932 ( .B1(n13975), .B2(n13974), .A(n7401), .ZN(n13963) );
  AND2_X1 U7933 ( .A1(n13988), .A2(n13392), .ZN(n7401) );
  OAI22_X1 U7934 ( .A1(n9717), .A2(n9716), .B1(n13977), .B2(n13475), .ZN(
        n13975) );
  NOR2_X1 U7935 ( .A1(n14151), .A2(n14002), .ZN(n9716) );
  NAND2_X1 U7936 ( .A1(n14004), .A2(n13355), .ZN(n13991) );
  NAND2_X1 U7937 ( .A1(n7402), .A2(n8431), .ZN(n9717) );
  AOI21_X1 U7938 ( .B1(n8434), .B2(n8436), .A(n8432), .ZN(n8431) );
  NAND2_X1 U7939 ( .A1(n14026), .A2(n8434), .ZN(n7402) );
  INV_X1 U7940 ( .A(n7334), .ZN(n8432) );
  OR2_X1 U7941 ( .A1(n8439), .A2(n8438), .ZN(n8437) );
  INV_X1 U7942 ( .A(n8441), .ZN(n8438) );
  AND2_X1 U7943 ( .A1(n13281), .A2(n8440), .ZN(n8439) );
  NAND2_X1 U7944 ( .A1(n7244), .A2(n9675), .ZN(n8440) );
  AND2_X1 U7945 ( .A1(n14056), .A2(n13171), .ZN(n8456) );
  AOI21_X1 U7946 ( .B1(n7622), .B2(n7624), .A(n7619), .ZN(n7618) );
  INV_X1 U7947 ( .A(n13157), .ZN(n7624) );
  AOI21_X1 U7948 ( .B1(n14105), .B2(n8425), .A(n8424), .ZN(n8423) );
  NAND2_X1 U7949 ( .A1(n9561), .A2(n8422), .ZN(n8421) );
  NAND2_X1 U7950 ( .A1(n7621), .A2(n13157), .ZN(n14094) );
  NAND2_X1 U7951 ( .A1(n14102), .A2(n8426), .ZN(n7621) );
  NAND2_X1 U7952 ( .A1(n14094), .A2(n14093), .ZN(n14092) );
  AND2_X1 U7953 ( .A1(n13156), .A2(n13331), .ZN(n13275) );
  AOI21_X1 U7954 ( .B1(n7195), .B2(n13271), .A(n12152), .ZN(n8039) );
  NAND2_X1 U7955 ( .A1(n8037), .A2(n7195), .ZN(n8038) );
  NAND2_X1 U7956 ( .A1(n12101), .A2(n13257), .ZN(n12100) );
  OR2_X1 U7957 ( .A1(n9478), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U7958 ( .A1(n11467), .A2(n9462), .ZN(n11622) );
  AND2_X1 U7959 ( .A1(n13114), .A2(n13115), .ZN(n13113) );
  NAND2_X1 U7960 ( .A1(n11633), .A2(n9418), .ZN(n11032) );
  INV_X1 U7961 ( .A(n13265), .ZN(n11031) );
  OR2_X1 U7962 ( .A1(n9705), .A2(n10158), .ZN(n9417) );
  NAND2_X1 U7963 ( .A1(n16030), .A2(n13270), .ZN(n8461) );
  OR2_X1 U7964 ( .A1(n9705), .A2(n10164), .ZN(n9404) );
  INV_X1 U7965 ( .A(n14108), .ZN(n16034) );
  NAND2_X1 U7966 ( .A1(n10601), .A2(n13229), .ZN(n16032) );
  AND2_X1 U7967 ( .A1(n9852), .A2(n13304), .ZN(n16039) );
  INV_X1 U7968 ( .A(n16039), .ZN(n14103) );
  AND3_X1 U7969 ( .A1(n9384), .A2(n9383), .A3(n9382), .ZN(n11640) );
  OR2_X1 U7970 ( .A1(n9443), .A2(n10173), .ZN(n9383) );
  OR2_X1 U7971 ( .A1(n9705), .A2(n10174), .ZN(n9384) );
  OR2_X1 U7972 ( .A1(n9443), .A2(n13643), .ZN(n9375) );
  NAND2_X1 U7973 ( .A1(n13980), .A2(n13979), .ZN(n14147) );
  NAND2_X1 U7974 ( .A1(n9620), .A2(n9619), .ZN(n14179) );
  OR2_X1 U7975 ( .A1(n10429), .A2(n9705), .ZN(n9620) );
  AND3_X1 U7976 ( .A1(n14250), .A2(n9850), .A3(n14248), .ZN(n10464) );
  INV_X1 U7977 ( .A(n16032), .ZN(n14107) );
  INV_X1 U7978 ( .A(n9845), .ZN(n10244) );
  NAND2_X1 U7979 ( .A1(n14255), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9358) );
  XNOR2_X1 U7980 ( .A(n9823), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9858) );
  XNOR2_X1 U7981 ( .A(n9310), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n9729) );
  INV_X1 U7982 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9332) );
  INV_X1 U7983 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9331) );
  INV_X1 U7984 ( .A(n9825), .ZN(n9827) );
  NAND2_X1 U7985 ( .A1(n9704), .A2(n9306), .ZN(n9719) );
  XNOR2_X1 U7986 ( .A(n9856), .B(n9855), .ZN(n10432) );
  INV_X1 U7987 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9855) );
  OAI21_X1 U7988 ( .B1(n7234), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9856) );
  INV_X1 U7989 ( .A(n9299), .ZN(n7987) );
  NAND2_X1 U7990 ( .A1(n9664), .A2(n9299), .ZN(n9677) );
  AND2_X1 U7991 ( .A1(n9301), .A2(n9300), .ZN(n9676) );
  NAND2_X1 U7992 ( .A1(n9662), .A2(n9661), .ZN(n9664) );
  NAND2_X1 U7993 ( .A1(n9649), .A2(n9297), .ZN(n9662) );
  NAND2_X1 U7994 ( .A1(n9647), .A2(n9646), .ZN(n9649) );
  INV_X1 U7995 ( .A(n7993), .ZN(n7992) );
  OAI21_X1 U7996 ( .B1(n9612), .B2(n7994), .A(n9628), .ZN(n7993) );
  INV_X1 U7997 ( .A(n9293), .ZN(n7994) );
  NAND2_X1 U7998 ( .A1(n9615), .A2(n9293), .ZN(n9629) );
  NAND2_X1 U7999 ( .A1(n9613), .A2(n9612), .ZN(n9615) );
  NAND2_X1 U8000 ( .A1(n9597), .A2(n9291), .ZN(n9613) );
  NAND2_X1 U8001 ( .A1(n9582), .A2(n9289), .ZN(n9595) );
  NAND2_X1 U8002 ( .A1(n9595), .A2(n9594), .ZN(n9597) );
  NAND2_X1 U8003 ( .A1(n9580), .A2(n9579), .ZN(n9582) );
  INV_X1 U8004 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9583) );
  AND2_X1 U8005 ( .A1(n9549), .A2(n9548), .ZN(n9567) );
  NAND2_X1 U8006 ( .A1(n9542), .A2(n9541), .ZN(n9544) );
  INV_X1 U8007 ( .A(n9282), .ZN(n7980) );
  NAND2_X1 U8008 ( .A1(n9521), .A2(n9282), .ZN(n9527) );
  AND2_X1 U8009 ( .A1(n9284), .A2(n9283), .ZN(n9526) );
  INV_X1 U8010 ( .A(n7979), .ZN(n7978) );
  OAI21_X1 U8011 ( .B1(n9518), .B2(n7980), .A(n9526), .ZN(n7979) );
  NAND2_X1 U8012 ( .A1(n9519), .A2(n9518), .ZN(n9521) );
  NAND2_X1 U8013 ( .A1(n9504), .A2(n9280), .ZN(n9519) );
  NAND2_X1 U8014 ( .A1(n9502), .A2(n9501), .ZN(n9504) );
  OR2_X1 U8015 ( .A1(n9506), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9617) );
  AND2_X1 U8016 ( .A1(n9278), .A2(n9277), .ZN(n9488) );
  AND2_X1 U8017 ( .A1(n9269), .A2(n9268), .ZN(n9429) );
  NAND2_X1 U8018 ( .A1(n9267), .A2(n9266), .ZN(n9430) );
  XNOR2_X1 U8019 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9259) );
  INV_X1 U8020 ( .A(n11682), .ZN(n7857) );
  NAND2_X1 U8021 ( .A1(n14421), .A2(n14295), .ZN(n14298) );
  XNOR2_X1 U8022 ( .A(n14304), .B(n11603), .ZN(n11088) );
  NAND2_X1 U8023 ( .A1(n12044), .A2(n12045), .ZN(n12228) );
  NAND2_X1 U8024 ( .A1(n8600), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8909) );
  OR2_X1 U8025 ( .A1(n8909), .A2(n14414), .ZN(n8921) );
  XNOR2_X1 U8026 ( .A(n14294), .B(n14292), .ZN(n14419) );
  INV_X1 U8027 ( .A(n14273), .ZN(n7866) );
  INV_X1 U8028 ( .A(n7865), .ZN(n7864) );
  OAI21_X1 U8029 ( .B1(n14378), .B2(n7866), .A(n14390), .ZN(n7865) );
  NAND2_X1 U8030 ( .A1(n8403), .A2(n14270), .ZN(n8402) );
  NAND2_X1 U8031 ( .A1(n7867), .A2(n7215), .ZN(n8404) );
  INV_X1 U8032 ( .A(n8405), .ZN(n8403) );
  AND4_X1 U8033 ( .A1(n8845), .A2(n8844), .A3(n8843), .A4(n8842), .ZN(n14381)
         );
  AND4_X1 U8034 ( .A1(n8728), .A2(n8727), .A3(n8726), .A4(n8725), .ZN(n11679)
         );
  AND3_X1 U8035 ( .A1(n8618), .A2(n7771), .A3(n8617), .ZN(n8631) );
  AOI22_X1 U8036 ( .A1(n8649), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n8885), .B2(
        P2_REG2_REG_1__SCAN_IN), .ZN(n7771) );
  OAI21_X1 U8037 ( .B1(n7590), .B2(n8366), .A(n9100), .ZN(n7586) );
  INV_X1 U8038 ( .A(n14465), .ZN(n14318) );
  OAI21_X1 U8039 ( .B1(n8365), .B2(n8363), .A(n10110), .ZN(n9238) );
  NAND2_X1 U8040 ( .A1(n8369), .A2(n8364), .ZN(n8363) );
  INV_X1 U8041 ( .A(n7578), .ZN(n7577) );
  AND2_X1 U8042 ( .A1(n8991), .A2(n8990), .ZN(n14582) );
  OAI21_X1 U8043 ( .B1(n14611), .B2(n14594), .A(n8154), .ZN(n14593) );
  OAI22_X1 U8044 ( .A1(n14667), .A2(n7602), .B1(n14648), .B2(n14925), .ZN(
        n7598) );
  NAND2_X1 U8045 ( .A1(n14682), .A2(n7600), .ZN(n7599) );
  NOR2_X1 U8046 ( .A1(n14667), .A2(n7601), .ZN(n7600) );
  INV_X1 U8047 ( .A(n14681), .ZN(n7601) );
  NOR2_X1 U8048 ( .A1(n8914), .A2(n8151), .ZN(n8150) );
  NAND2_X1 U8049 ( .A1(n8891), .A2(n8890), .ZN(n14692) );
  INV_X1 U8050 ( .A(n14688), .ZN(n14693) );
  NAND2_X1 U8051 ( .A1(n8882), .A2(n8881), .ZN(n14713) );
  OR2_X1 U8052 ( .A1(n12834), .A2(n10024), .ZN(n8882) );
  INV_X1 U8053 ( .A(n10104), .ZN(n14707) );
  NAND2_X1 U8054 ( .A1(n14872), .A2(n14470), .ZN(n7746) );
  NAND3_X1 U8055 ( .A1(n7556), .A2(n14779), .A3(n7554), .ZN(n14778) );
  INV_X1 U8056 ( .A(n7558), .ZN(n7555) );
  AND2_X1 U8057 ( .A1(n12326), .A2(n7256), .ZN(n8148) );
  AND2_X1 U8058 ( .A1(n9040), .A2(n8793), .ZN(n12329) );
  NAND2_X1 U8059 ( .A1(n11894), .A2(n8744), .ZN(n11934) );
  INV_X1 U8060 ( .A(n14600), .ZN(n14791) );
  NAND2_X1 U8061 ( .A1(n11420), .A2(n9033), .ZN(n7595) );
  NAND2_X1 U8062 ( .A1(n7604), .A2(n10994), .ZN(n7603) );
  NAND2_X1 U8063 ( .A1(n11412), .A2(n11413), .ZN(n11411) );
  XNOR2_X1 U8064 ( .A(n14483), .B(n11724), .ZN(n11407) );
  NAND2_X1 U8065 ( .A1(n9026), .A2(n11393), .ZN(n11392) );
  NAND2_X1 U8066 ( .A1(n10896), .A2(n9064), .ZN(n14600) );
  NAND2_X1 U8067 ( .A1(n10896), .A2(n9065), .ZN(n14794) );
  INV_X1 U8068 ( .A(n14584), .ZN(n14819) );
  AND2_X1 U8069 ( .A1(n14603), .A2(n14602), .ZN(n14824) );
  NAND2_X1 U8070 ( .A1(n8963), .A2(n8962), .ZN(n14830) );
  XNOR2_X1 U8071 ( .A(n14641), .B(n14646), .ZN(n14629) );
  NAND2_X1 U8072 ( .A1(n14756), .A2(n14757), .ZN(n8147) );
  NAND2_X1 U8073 ( .A1(n8147), .A2(n8145), .ZN(n14743) );
  NOR2_X1 U8074 ( .A1(n14740), .A2(n8146), .ZN(n8145) );
  INV_X1 U8075 ( .A(n8847), .ZN(n8146) );
  AND2_X1 U8076 ( .A1(n14786), .A2(n8806), .ZN(n8141) );
  AND2_X1 U8077 ( .A1(n8801), .A2(n8800), .ZN(n16202) );
  NAND2_X1 U8078 ( .A1(n8751), .A2(n8750), .ZN(n11944) );
  OR2_X1 U8079 ( .A1(n11805), .A2(n10024), .ZN(n8751) );
  NAND2_X1 U8080 ( .A1(n7247), .A2(n7584), .ZN(n7583) );
  NAND2_X1 U8081 ( .A1(n8715), .A2(n8714), .ZN(n11508) );
  NAND2_X1 U8082 ( .A1(n7747), .A2(n8682), .ZN(n11416) );
  XNOR2_X1 U8083 ( .A(n11603), .B(n14481), .ZN(n11597) );
  NAND2_X1 U8084 ( .A1(n11230), .A2(n10832), .ZN(n16201) );
  NAND2_X1 U8085 ( .A1(n8656), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7772) );
  OR2_X1 U8086 ( .A1(n14965), .A2(n9078), .ZN(n9097) );
  INV_X1 U8087 ( .A(n8588), .ZN(n7725) );
  INV_X1 U8088 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9069) );
  OAI21_X1 U8089 ( .B1(n9079), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9076) );
  INV_X1 U8090 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8477) );
  AOI21_X1 U8091 ( .B1(n8277), .B2(n8279), .A(n7298), .ZN(n8274) );
  INV_X1 U8092 ( .A(n7349), .ZN(n7841) );
  AOI21_X1 U8093 ( .B1(n8271), .B2(n8269), .A(n7283), .ZN(n8268) );
  INV_X1 U8094 ( .A(n8273), .ZN(n8269) );
  AND2_X1 U8095 ( .A1(n15200), .A2(n8278), .ZN(n8277) );
  OR2_X1 U8096 ( .A1(n15124), .A2(n8279), .ZN(n8278) );
  AND2_X1 U8097 ( .A1(n11772), .A2(n11773), .ZN(n7816) );
  NAND2_X1 U8098 ( .A1(n15161), .A2(n7271), .ZN(n15113) );
  NOR2_X1 U8099 ( .A1(n11127), .A2(n11126), .ZN(n8264) );
  AOI21_X1 U8100 ( .B1(n8263), .B2(n10860), .A(n8261), .ZN(n8260) );
  NAND2_X1 U8101 ( .A1(n10859), .A2(n8263), .ZN(n8262) );
  INV_X1 U8102 ( .A(n11126), .ZN(n8261) );
  NAND2_X1 U8103 ( .A1(n7805), .A2(n7804), .ZN(n11907) );
  AND2_X1 U8104 ( .A1(n7802), .A2(n7811), .ZN(n7804) );
  NAND2_X1 U8105 ( .A1(n11314), .A2(n7806), .ZN(n7805) );
  AND2_X1 U8106 ( .A1(n11783), .A2(n7812), .ZN(n7811) );
  NAND2_X1 U8107 ( .A1(n10384), .A2(n10383), .ZN(n10851) );
  OR2_X1 U8108 ( .A1(n12582), .A2(n7835), .ZN(n7834) );
  INV_X1 U8109 ( .A(n7842), .ZN(n7835) );
  INV_X1 U8110 ( .A(n8285), .ZN(n8284) );
  NAND2_X1 U8111 ( .A1(n13002), .A2(n13001), .ZN(n15354) );
  NAND2_X1 U8112 ( .A1(n7487), .A2(n15427), .ZN(n15423) );
  NOR2_X1 U8113 ( .A1(n8191), .A2(n15434), .ZN(n8189) );
  INV_X1 U8114 ( .A(n8191), .ZN(n8188) );
  NAND2_X1 U8115 ( .A1(n7546), .A2(n8118), .ZN(n7545) );
  INV_X1 U8116 ( .A(n8187), .ZN(n15465) );
  NOR2_X1 U8117 ( .A1(n15504), .A2(n15662), .ZN(n15491) );
  INV_X1 U8118 ( .A(n15377), .ZN(n15487) );
  OR2_X1 U8119 ( .A1(n15508), .A2(n15406), .ZN(n8464) );
  AND2_X1 U8120 ( .A1(n8115), .A2(n8113), .ZN(n15485) );
  NOR2_X1 U8121 ( .A1(n15509), .A2(n8204), .ZN(n8203) );
  INV_X1 U8122 ( .A(n15405), .ZN(n8204) );
  NAND2_X1 U8123 ( .A1(n8027), .A2(n15529), .ZN(n15524) );
  NAND2_X1 U8124 ( .A1(n7468), .A2(n7467), .ZN(n7464) );
  NAND2_X1 U8125 ( .A1(n7469), .A2(n7466), .ZN(n7465) );
  NOR2_X1 U8126 ( .A1(n7468), .A2(n7467), .ZN(n7466) );
  AND2_X1 U8127 ( .A1(n15672), .A2(n15376), .ZN(n7362) );
  NAND2_X1 U8128 ( .A1(n8205), .A2(n8206), .ZN(n15520) );
  AOI21_X1 U8129 ( .B1(n8096), .B2(n8094), .A(n7285), .ZN(n8093) );
  INV_X1 U8130 ( .A(n8096), .ZN(n8095) );
  NAND2_X1 U8131 ( .A1(n8197), .A2(n15401), .ZN(n8194) );
  NAND2_X1 U8132 ( .A1(n15568), .A2(n15550), .ZN(n15552) );
  NAND2_X1 U8133 ( .A1(n15562), .A2(n8094), .ZN(n15561) );
  NOR2_X1 U8134 ( .A1(n13029), .A2(n8199), .ZN(n8198) );
  NAND2_X1 U8135 ( .A1(n12655), .A2(n12660), .ZN(n15395) );
  INV_X1 U8136 ( .A(n8105), .ZN(n8104) );
  NAND2_X1 U8137 ( .A1(n12195), .A2(n12194), .ZN(n12805) );
  NAND2_X1 U8138 ( .A1(n12072), .A2(n8073), .ZN(n12173) );
  NAND2_X1 U8139 ( .A1(n12018), .A2(n12017), .ZN(n12793) );
  XNOR2_X1 U8140 ( .A(n12770), .B(n15233), .ZN(n12767) );
  INV_X1 U8141 ( .A(n12767), .ZN(n13014) );
  NOR2_X1 U8142 ( .A1(n16070), .A2(n11239), .ZN(n8182) );
  NAND2_X1 U8143 ( .A1(n16070), .A2(n11239), .ZN(n8183) );
  OAI21_X1 U8144 ( .B1(n10779), .B2(n13012), .A(n7540), .ZN(n10750) );
  AOI21_X1 U8145 ( .B1(n7539), .B2(n10705), .A(n7538), .ZN(n7540) );
  INV_X1 U8146 ( .A(n10695), .ZN(n7539) );
  INV_X1 U8147 ( .A(n10746), .ZN(n7538) );
  INV_X1 U8148 ( .A(n12754), .ZN(n13013) );
  OAI21_X1 U8149 ( .B1(n8023), .B2(n7490), .A(n10691), .ZN(n7491) );
  OR2_X1 U8150 ( .A1(n10691), .A2(n10693), .ZN(n8024) );
  NOR2_X1 U8151 ( .A1(n9343), .A2(n10690), .ZN(n7490) );
  NAND2_X1 U8152 ( .A1(n8089), .A2(n8087), .ZN(n15419) );
  NAND2_X1 U8153 ( .A1(n8090), .A2(n7241), .ZN(n8089) );
  NAND2_X1 U8154 ( .A1(n12943), .A2(n12942), .ZN(n15643) );
  OAI22_X1 U8155 ( .A1(n13000), .A2(n10749), .B1(n10691), .B2(n15270), .ZN(
        n7799) );
  NAND2_X1 U8156 ( .A1(n9103), .A2(n9102), .ZN(n10019) );
  INV_X1 U8157 ( .A(n8076), .ZN(n8075) );
  NAND2_X1 U8158 ( .A1(n8084), .A2(n8080), .ZN(n8079) );
  XNOR2_X1 U8159 ( .A(n10370), .B(P1_IR_REG_29__SCAN_IN), .ZN(n10372) );
  NAND2_X1 U8160 ( .A1(n7550), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10370) );
  AND4_X1 U8161 ( .A1(n8058), .A2(n8057), .A3(n10218), .A4(n8469), .ZN(n7551)
         );
  OR2_X1 U8162 ( .A1(n10150), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n7204) );
  XNOR2_X1 U8163 ( .A(n8984), .B(n7348), .ZN(n14963) );
  NAND2_X1 U8164 ( .A1(n7899), .A2(n8578), .ZN(n8984) );
  NAND2_X1 U8165 ( .A1(n8574), .A2(n7903), .ZN(n7899) );
  NAND2_X1 U8166 ( .A1(n8574), .A2(n8573), .ZN(n8975) );
  XNOR2_X1 U8167 ( .A(n10144), .B(P1_IR_REG_23__SCAN_IN), .ZN(n10421) );
  XNOR2_X1 U8168 ( .A(n8948), .B(n8947), .ZN(n14971) );
  XNOR2_X1 U8169 ( .A(n8943), .B(n13652), .ZN(n12882) );
  NAND2_X1 U8170 ( .A1(n10217), .A2(n7711), .ZN(n12991) );
  AND2_X1 U8171 ( .A1(n10216), .A2(n7712), .ZN(n7711) );
  OR2_X1 U8172 ( .A1(n10214), .A2(n10213), .ZN(n10217) );
  NAND2_X1 U8173 ( .A1(n7303), .A2(n7192), .ZN(n7712) );
  NAND2_X1 U8174 ( .A1(n7455), .A2(n8561), .ZN(n8917) );
  NAND2_X1 U8175 ( .A1(n10403), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10404) );
  NAND2_X1 U8176 ( .A1(n11612), .A2(n10146), .ZN(n10403) );
  XNOR2_X1 U8177 ( .A(n8893), .B(n8892), .ZN(n12727) );
  OAI21_X1 U8178 ( .B1(n8558), .B2(n7893), .A(n7892), .ZN(n8893) );
  NAND2_X1 U8179 ( .A1(n8384), .A2(n8383), .ZN(n8877) );
  NAND2_X1 U8180 ( .A1(n8374), .A2(SI_9_), .ZN(n8382) );
  NAND2_X1 U8181 ( .A1(n8540), .A2(n8539), .ZN(n8374) );
  NAND2_X1 U8182 ( .A1(n8524), .A2(n8523), .ZN(n8671) );
  OAI21_X1 U8183 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n9146), .A(n9145), .ZN(
        n9165) );
  INV_X1 U8184 ( .A(n15961), .ZN(n7438) );
  NAND2_X1 U8185 ( .A1(n9205), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7963) );
  AOI21_X1 U8186 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n12305), .A(n9152), .ZN(
        n9215) );
  AOI21_X1 U8187 ( .B1(n7658), .B2(n7660), .A(n7300), .ZN(n7655) );
  INV_X1 U8188 ( .A(n10739), .ZN(n8343) );
  NAND2_X1 U8189 ( .A1(n13476), .A2(n13345), .ZN(n13398) );
  NOR2_X1 U8190 ( .A1(n8348), .A2(n13440), .ZN(n8346) );
  NOR2_X1 U8191 ( .A1(n8349), .A2(n8351), .ZN(n8348) );
  NOR2_X1 U8192 ( .A1(n13407), .A2(n13403), .ZN(n8351) );
  INV_X1 U8193 ( .A(n8352), .ZN(n8349) );
  NAND2_X1 U8194 ( .A1(n8352), .A2(n8353), .ZN(n8350) );
  INV_X1 U8195 ( .A(n13407), .ZN(n8353) );
  NAND2_X1 U8196 ( .A1(n9763), .A2(n9762), .ZN(n13412) );
  OR2_X1 U8197 ( .A1(n9730), .A2(n13534), .ZN(n9762) );
  OR2_X1 U8198 ( .A1(n9705), .A2(n10167), .ZN(n9493) );
  OAI21_X1 U8199 ( .B1(n13102), .B2(n13888), .A(n10775), .ZN(n10596) );
  AND3_X1 U8200 ( .A1(n9686), .A2(n9685), .A3(n9684), .ZN(n14029) );
  NAND2_X1 U8201 ( .A1(n11102), .A2(n11101), .ZN(n11299) );
  AND2_X1 U8202 ( .A1(n9532), .A2(n9531), .ZN(n12366) );
  OR2_X1 U8203 ( .A1(n10640), .A2(n10639), .ZN(n7669) );
  XNOR2_X1 U8204 ( .A(n10736), .B(n13523), .ZN(n10641) );
  NAND2_X1 U8205 ( .A1(n7684), .A2(n7389), .ZN(n7388) );
  NAND2_X1 U8206 ( .A1(n13307), .A2(n13308), .ZN(n7684) );
  NAND2_X1 U8207 ( .A1(n13306), .A2(n13305), .ZN(n7389) );
  OAI22_X1 U8208 ( .A1(n13307), .A2(n13294), .B1(n13292), .B2(n13293), .ZN(
        n7390) );
  AND2_X1 U8209 ( .A1(n13251), .A2(n9783), .ZN(n13919) );
  NAND2_X1 U8210 ( .A1(n9700), .A2(n9699), .ZN(n14015) );
  INV_X1 U8211 ( .A(n14029), .ZN(n14001) );
  NAND2_X1 U8212 ( .A1(n7410), .A2(n10552), .ZN(n10562) );
  OR2_X1 U8213 ( .A1(n11983), .A2(n11982), .ZN(n12310) );
  OR2_X1 U8214 ( .A1(n12451), .A2(n12452), .ZN(n8165) );
  OR2_X1 U8215 ( .A1(n13814), .A2(n13813), .ZN(n7924) );
  INV_X1 U8216 ( .A(n8170), .ZN(n13825) );
  INV_X1 U8217 ( .A(n8168), .ZN(n13835) );
  NOR2_X1 U8218 ( .A1(n7416), .A2(n7257), .ZN(n7413) );
  OAI21_X1 U8219 ( .B1(n7932), .B2(n13882), .A(n13865), .ZN(n7416) );
  NAND2_X1 U8220 ( .A1(n13862), .A2(n7931), .ZN(n7930) );
  NOR2_X1 U8221 ( .A1(n13896), .A2(n8175), .ZN(n8174) );
  OR2_X1 U8222 ( .A1(n13864), .A2(n7929), .ZN(n7928) );
  XNOR2_X1 U8223 ( .A(n7756), .B(n7755), .ZN(n8176) );
  INV_X1 U8224 ( .A(n13892), .ZN(n7755) );
  NOR2_X1 U8225 ( .A1(n7447), .A2(n13891), .ZN(n7756) );
  INV_X1 U8226 ( .A(n14218), .ZN(n13968) );
  NAND2_X1 U8227 ( .A1(n10466), .A2(n10465), .ZN(n16128) );
  NAND2_X1 U8228 ( .A1(n9681), .A2(n9680), .ZN(n14227) );
  OR2_X1 U8229 ( .A1(n10777), .A2(n9705), .ZN(n9681) );
  NAND2_X1 U8230 ( .A1(n9637), .A2(n9636), .ZN(n14237) );
  OR2_X1 U8231 ( .A1(n9705), .A2(n10168), .ZN(n9476) );
  OR2_X1 U8232 ( .A1(n9705), .A2(n10161), .ZN(n9445) );
  OR2_X1 U8233 ( .A1(n9338), .A2(n9337), .ZN(n7683) );
  AOI21_X1 U8234 ( .B1(n9825), .B2(n7199), .A(n7682), .ZN(n7681) );
  OAI21_X1 U8235 ( .B1(n9339), .B2(P3_IR_REG_27__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9338) );
  XNOR2_X1 U8236 ( .A(n9787), .B(P3_IR_REG_22__SCAN_IN), .ZN(n13313) );
  AND2_X1 U8237 ( .A1(n8941), .A2(n8940), .ZN(n14362) );
  AND2_X1 U8238 ( .A1(n8772), .A2(n8771), .ZN(n16186) );
  INV_X1 U8239 ( .A(n14925), .ZN(n14368) );
  OAI22_X1 U8240 ( .A1(n12495), .A2(n12494), .B1(n12493), .B2(n12492), .ZN(
        n12496) );
  NAND2_X1 U8241 ( .A1(n8398), .A2(n11254), .ZN(n8395) );
  NAND2_X1 U8242 ( .A1(n8397), .A2(n8398), .ZN(n8396) );
  INV_X1 U8243 ( .A(n11258), .ZN(n8398) );
  OAI21_X1 U8244 ( .B1(n14379), .B2(n7866), .A(n7864), .ZN(n14388) );
  AND2_X1 U8245 ( .A1(n8957), .A2(n8956), .ZN(n14401) );
  AND4_X1 U8246 ( .A1(n8805), .A2(n8804), .A3(n8803), .A4(n8802), .ZN(n14795)
         );
  NAND2_X1 U8247 ( .A1(n8813), .A2(n8812), .ZN(n14800) );
  INV_X1 U8248 ( .A(n14654), .ZN(n14840) );
  AND4_X1 U8249 ( .A1(n8779), .A2(n8778), .A3(n8777), .A4(n8776), .ZN(n12335)
         );
  NOR2_X1 U8250 ( .A1(n8235), .A2(n10126), .ZN(n8233) );
  NOR2_X1 U8251 ( .A1(n10113), .A2(n10120), .ZN(n8235) );
  NAND2_X1 U8252 ( .A1(n8983), .A2(n8982), .ZN(n14614) );
  NAND2_X1 U8253 ( .A1(n8971), .A2(n8970), .ZN(n14633) );
  INV_X1 U8254 ( .A(n14401), .ZN(n14646) );
  INV_X1 U8255 ( .A(n14289), .ZN(n14648) );
  AND4_X1 U8256 ( .A1(n8873), .A2(n8872), .A3(n8871), .A4(n8870), .ZN(n14433)
         );
  INV_X1 U8257 ( .A(n12038), .ZN(n14476) );
  AND2_X1 U8258 ( .A1(n10929), .A2(n13321), .ZN(n15888) );
  INV_X1 U8259 ( .A(n14563), .ZN(n7749) );
  NAND2_X1 U8260 ( .A1(n7611), .A2(n9045), .ZN(n14758) );
  AND2_X1 U8261 ( .A1(n8839), .A2(n8838), .ZN(n14879) );
  OR2_X1 U8262 ( .A1(n16094), .A2(n11547), .ZN(n16062) );
  OR2_X1 U8263 ( .A1(n10838), .A2(n15818), .ZN(n14697) );
  NOR2_X1 U8264 ( .A1(n16208), .A2(n8391), .ZN(n8390) );
  INV_X1 U8265 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8391) );
  NOR2_X1 U8266 ( .A1(n9066), .A2(n14356), .ZN(n14557) );
  NAND2_X1 U8267 ( .A1(n7609), .A2(n7607), .ZN(n9057) );
  INV_X1 U8268 ( .A(n9025), .ZN(n14559) );
  NAND2_X1 U8269 ( .A1(n7589), .A2(n7588), .ZN(n9101) );
  NAND2_X1 U8270 ( .A1(n16208), .A2(n16204), .ZN(n8387) );
  OR2_X1 U8271 ( .A1(n14562), .A2(n16206), .ZN(n8389) );
  OR2_X1 U8272 ( .A1(n9235), .A2(n9234), .ZN(n9249) );
  INV_X1 U8273 ( .A(n12425), .ZN(n12422) );
  NAND2_X1 U8274 ( .A1(n16208), .A2(n16134), .ZN(n14896) );
  NAND2_X1 U8275 ( .A1(n10046), .A2(n10045), .ZN(n14902) );
  NAND2_X1 U8276 ( .A1(n10027), .A2(n10026), .ZN(n14905) );
  OAI211_X1 U8277 ( .C1(n14559), .C2(n16138), .A(n14557), .B(n8157), .ZN(n8156) );
  AND2_X1 U8278 ( .A1(n14562), .A2(n14948), .ZN(n8157) );
  NAND2_X1 U8279 ( .A1(n14575), .A2(n14571), .ZN(n9247) );
  AND2_X2 U8280 ( .A1(n9125), .A2(n15820), .ZN(n14948) );
  INV_X1 U8281 ( .A(n15821), .ZN(n15818) );
  XNOR2_X1 U8282 ( .A(n8502), .B(n8501), .ZN(n12683) );
  INV_X1 U8283 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10360) );
  NAND2_X1 U8284 ( .A1(n12523), .A2(n12522), .ZN(n15733) );
  NOR2_X1 U8285 ( .A1(n7820), .A2(n15205), .ZN(n7818) );
  AND2_X1 U8286 ( .A1(n7823), .A2(n7324), .ZN(n7820) );
  INV_X1 U8287 ( .A(n15100), .ZN(n7822) );
  NAND2_X1 U8288 ( .A1(n7823), .A2(n7826), .ZN(n7821) );
  NAND2_X1 U8289 ( .A1(n15100), .A2(n15092), .ZN(n7826) );
  INV_X1 U8290 ( .A(n15225), .ZN(n12584) );
  NAND2_X1 U8291 ( .A1(n15046), .A2(n15045), .ZN(n15123) );
  NAND2_X1 U8292 ( .A1(n12654), .A2(n12653), .ZN(n15719) );
  NAND2_X1 U8293 ( .A1(n12838), .A2(n12837), .ZN(n15705) );
  OR2_X1 U8294 ( .A1(n12834), .A2(n12987), .ZN(n12838) );
  INV_X1 U8295 ( .A(n15220), .ZN(n15196) );
  AND2_X1 U8296 ( .A1(n10861), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15216) );
  NAND2_X1 U8297 ( .A1(n15299), .A2(n7274), .ZN(n10308) );
  NOR2_X1 U8298 ( .A1(n10313), .A2(n10314), .ZN(n10346) );
  NAND2_X1 U8299 ( .A1(n15312), .A2(n7336), .ZN(n10579) );
  NAND2_X1 U8300 ( .A1(n12989), .A2(n12988), .ZN(n15361) );
  XNOR2_X1 U8301 ( .A(n15382), .B(n15412), .ZN(n15628) );
  OAI21_X1 U8302 ( .B1(n8090), .B2(n8088), .A(n8085), .ZN(n15382) );
  AOI21_X1 U8303 ( .B1(n8087), .B2(n8086), .A(n7276), .ZN(n8085) );
  AND2_X1 U8304 ( .A1(n7484), .A2(n7536), .ZN(n8068) );
  NOR2_X1 U8305 ( .A1(n15632), .A2(n7537), .ZN(n7536) );
  NAND2_X1 U8306 ( .A1(n15629), .A2(n16176), .ZN(n7484) );
  INV_X1 U8307 ( .A(n8022), .ZN(n7537) );
  INV_X1 U8308 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10359) );
  INV_X1 U8309 ( .A(n9182), .ZN(n7429) );
  XNOR2_X1 U8310 ( .A(n9186), .B(n9187), .ZN(n15948) );
  XNOR2_X1 U8311 ( .A(n9209), .B(n7962), .ZN(n15969) );
  INV_X1 U8312 ( .A(n9208), .ZN(n7962) );
  NAND2_X1 U8313 ( .A1(n15969), .A2(n15968), .ZN(n15967) );
  NAND2_X1 U8314 ( .A1(n7972), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7971) );
  OR2_X1 U8315 ( .A1(n15991), .A2(n15990), .ZN(n7970) );
  AND2_X1 U8316 ( .A1(n10976), .A2(n9243), .ZN(n9881) );
  AND2_X1 U8317 ( .A1(n9905), .A2(n9904), .ZN(n7372) );
  AND2_X1 U8318 ( .A1(n12754), .A2(n12753), .ZN(n12755) );
  NAND2_X1 U8319 ( .A1(n7495), .A2(n12779), .ZN(n7494) );
  OR2_X1 U8320 ( .A1(n8248), .A2(n8246), .ZN(n7364) );
  OAI21_X1 U8321 ( .B1(n12782), .B2(n7509), .A(n7508), .ZN(n12787) );
  NAND2_X1 U8322 ( .A1(n7507), .A2(n7505), .ZN(n12786) );
  AND2_X1 U8323 ( .A1(n12788), .A2(n7506), .ZN(n7505) );
  NAND2_X1 U8324 ( .A1(n7509), .A2(n7508), .ZN(n7506) );
  NAND2_X1 U8325 ( .A1(n7753), .A2(n7752), .ZN(n9940) );
  OR2_X1 U8326 ( .A1(n9936), .A2(n9935), .ZN(n7752) );
  INV_X1 U8327 ( .A(n12799), .ZN(n8296) );
  NAND2_X1 U8328 ( .A1(n8297), .A2(n12799), .ZN(n8294) );
  INV_X1 U8329 ( .A(n12794), .ZN(n7527) );
  NAND2_X1 U8330 ( .A1(n12794), .A2(n7526), .ZN(n7525) );
  OR2_X1 U8331 ( .A1(n8231), .A2(n9947), .ZN(n8230) );
  INV_X1 U8332 ( .A(n9946), .ZN(n8231) );
  AOI22_X1 U8333 ( .A1(n8300), .A2(n8307), .B1(n8301), .B2(n8304), .ZN(n8299)
         );
  NAND2_X1 U8334 ( .A1(n8305), .A2(n12814), .ZN(n8304) );
  NAND2_X1 U8335 ( .A1(n7374), .A2(n8238), .ZN(n9959) );
  NAND2_X1 U8336 ( .A1(n9956), .A2(n9957), .ZN(n8238) );
  OAI21_X1 U8337 ( .B1(n7522), .B2(n12840), .A(n7521), .ZN(n12845) );
  INV_X1 U8338 ( .A(n9970), .ZN(n8228) );
  NAND2_X1 U8339 ( .A1(n12845), .A2(n12846), .ZN(n12844) );
  INV_X1 U8340 ( .A(n12859), .ZN(n7520) );
  AND2_X1 U8341 ( .A1(n7327), .A2(n7518), .ZN(n7517) );
  NAND2_X1 U8342 ( .A1(n7519), .A2(n12859), .ZN(n7518) );
  NAND2_X1 U8343 ( .A1(n7378), .A2(n8213), .ZN(n9988) );
  AOI22_X1 U8344 ( .A1(n8219), .A2(n8222), .B1(n8217), .B2(n8218), .ZN(n8213)
         );
  INV_X1 U8345 ( .A(n7275), .ZN(n8218) );
  OR2_X1 U8346 ( .A1(n12885), .A2(n7196), .ZN(n7499) );
  NAND2_X1 U8347 ( .A1(n7502), .A2(n7500), .ZN(n12897) );
  AOI21_X1 U8348 ( .B1(n7196), .B2(n7503), .A(n7501), .ZN(n7500) );
  INV_X1 U8349 ( .A(n9990), .ZN(n8227) );
  INV_X1 U8350 ( .A(n12911), .ZN(n7713) );
  NAND2_X1 U8351 ( .A1(n12921), .A2(n8309), .ZN(n8308) );
  INV_X1 U8352 ( .A(n12920), .ZN(n8309) );
  NAND2_X1 U8353 ( .A1(n8241), .A2(n8242), .ZN(n10000) );
  NAND2_X1 U8354 ( .A1(n9998), .A2(n9999), .ZN(n8242) );
  INV_X1 U8355 ( .A(n10000), .ZN(n7384) );
  INV_X1 U8356 ( .A(n8835), .ZN(n7459) );
  NAND2_X1 U8357 ( .A1(n14611), .A2(n8362), .ZN(n8368) );
  INV_X1 U8358 ( .A(n8942), .ZN(n7571) );
  NAND2_X1 U8359 ( .A1(n7511), .A2(n7510), .ZN(n12956) );
  AOI21_X1 U8360 ( .B1(n7205), .B2(n7514), .A(n7293), .ZN(n7510) );
  NAND2_X1 U8361 ( .A1(n12932), .A2(n7205), .ZN(n7511) );
  INV_X1 U8362 ( .A(n8203), .ZN(n8201) );
  AND2_X1 U8363 ( .A1(n13019), .A2(n8063), .ZN(n8062) );
  NAND2_X1 U8364 ( .A1(n8064), .A2(n11700), .ZN(n8063) );
  INV_X1 U8365 ( .A(n11698), .ZN(n8064) );
  INV_X1 U8366 ( .A(n11700), .ZN(n8065) );
  NAND2_X1 U8367 ( .A1(n8083), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8082) );
  INV_X1 U8368 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8083) );
  NAND2_X1 U8369 ( .A1(n7452), .A2(n8563), .ZN(n7451) );
  INV_X1 U8370 ( .A(n8562), .ZN(n7452) );
  INV_X1 U8371 ( .A(n8561), .ZN(n7454) );
  NOR2_X1 U8372 ( .A1(n8892), .A2(n7891), .ZN(n7890) );
  INV_X1 U8373 ( .A(n7892), .ZN(n7891) );
  INV_X1 U8374 ( .A(n8892), .ZN(n7888) );
  AND2_X1 U8375 ( .A1(n7893), .A2(n7892), .ZN(n7887) );
  NAND2_X1 U8376 ( .A1(n7252), .A2(n7874), .ZN(n7873) );
  NAND2_X1 U8377 ( .A1(n10178), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7874) );
  INV_X1 U8378 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9128) );
  INV_X1 U8379 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9134) );
  INV_X1 U8380 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13705) );
  NOR2_X1 U8381 ( .A1(n9535), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7400) );
  NAND2_X1 U8382 ( .A1(n8359), .A2(n7649), .ZN(n7648) );
  INV_X1 U8383 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13709) );
  NOR2_X1 U8384 ( .A1(n7674), .A2(n13988), .ZN(n7672) );
  INV_X1 U8385 ( .A(n13450), .ZN(n7674) );
  NAND2_X1 U8386 ( .A1(n7395), .A2(n8013), .ZN(n13228) );
  NOR2_X1 U8387 ( .A1(n13286), .A2(n13216), .ZN(n8013) );
  INV_X1 U8388 ( .A(n13228), .ZN(n13227) );
  NAND2_X1 U8389 ( .A1(n7781), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U8390 ( .A1(n7949), .A2(n7957), .ZN(n7947) );
  INV_X1 U8391 ( .A(n7955), .ZN(n7952) );
  NOR2_X1 U8392 ( .A1(n7957), .A2(n7953), .ZN(n7948) );
  OR2_X1 U8393 ( .A1(n7634), .A2(n13938), .ZN(n7633) );
  INV_X1 U8394 ( .A(n8031), .ZN(n7634) );
  OR2_X1 U8395 ( .A1(n9747), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9749) );
  NOR2_X1 U8396 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(n9722), .ZN(n7399) );
  AOI21_X1 U8397 ( .B1(n8437), .B2(n8435), .A(n7312), .ZN(n8434) );
  INV_X1 U8398 ( .A(n7242), .ZN(n8435) );
  INV_X1 U8399 ( .A(n8437), .ZN(n8436) );
  NOR2_X1 U8400 ( .A1(n9653), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7394) );
  INV_X1 U8401 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n13586) );
  INV_X1 U8402 ( .A(n8051), .ZN(n7619) );
  AOI21_X1 U8403 ( .B1(n8052), .B2(n8054), .A(n7218), .ZN(n8051) );
  AND2_X1 U8404 ( .A1(n8052), .A2(n7623), .ZN(n7622) );
  NAND2_X1 U8405 ( .A1(n14105), .A2(n13157), .ZN(n7623) );
  NOR2_X1 U8406 ( .A1(n9588), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7392) );
  NOR2_X1 U8407 ( .A1(n8426), .A2(n8428), .ZN(n8422) );
  INV_X1 U8408 ( .A(n14086), .ZN(n8424) );
  INV_X1 U8409 ( .A(n13332), .ZN(n8425) );
  OR2_X1 U8410 ( .A1(n16217), .A2(n14109), .ZN(n13156) );
  INV_X1 U8411 ( .A(n14250), .ZN(n9865) );
  NAND2_X1 U8412 ( .A1(n9359), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7642) );
  OAI22_X1 U8413 ( .A1(n7199), .A2(n7642), .B1(n9359), .B2(
        P3_IR_REG_31__SCAN_IN), .ZN(n7639) );
  INV_X1 U8414 ( .A(n8000), .ZN(n7999) );
  OAI21_X1 U8415 ( .B1(n9429), .B2(n8001), .A(n9441), .ZN(n8000) );
  INV_X1 U8416 ( .A(n9269), .ZN(n8001) );
  INV_X1 U8417 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9260) );
  INV_X1 U8418 ( .A(n7870), .ZN(n7869) );
  AOI21_X1 U8419 ( .B1(n7870), .B2(n8409), .A(n7212), .ZN(n7868) );
  INV_X1 U8420 ( .A(n9236), .ZN(n8364) );
  INV_X1 U8421 ( .A(n8368), .ZN(n8365) );
  NAND2_X1 U8422 ( .A1(n7759), .A2(n7568), .ZN(n7567) );
  NOR2_X1 U8423 ( .A1(n7571), .A2(n7569), .ZN(n7568) );
  INV_X1 U8424 ( .A(n8926), .ZN(n7569) );
  INV_X1 U8425 ( .A(n8903), .ZN(n8151) );
  AOI21_X1 U8426 ( .B1(n8123), .B2(n8127), .A(n7197), .ZN(n8122) );
  INV_X1 U8427 ( .A(n8124), .ZN(n8123) );
  AND2_X1 U8428 ( .A1(n12146), .A2(n16186), .ZN(n12145) );
  INV_X1 U8429 ( .A(n11936), .ZN(n8134) );
  INV_X1 U8430 ( .A(n12683), .ZN(n10974) );
  INV_X1 U8431 ( .A(n9034), .ZN(n7593) );
  INV_X1 U8432 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U8433 ( .A1(n8491), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8880) );
  OR2_X1 U8434 ( .A1(n8731), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8749) );
  OR2_X1 U8435 ( .A1(n8718), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8731) );
  OR2_X1 U8436 ( .A1(n7808), .A2(n7329), .ZN(n7803) );
  AND2_X1 U8437 ( .A1(n7249), .A2(n11312), .ZN(n7808) );
  NOR2_X1 U8438 ( .A1(n11702), .A2(n11701), .ZN(n11811) );
  INV_X1 U8439 ( .A(n11127), .ZN(n8263) );
  AND2_X1 U8440 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n11131) );
  AND2_X1 U8441 ( .A1(n7815), .A2(n11774), .ZN(n7806) );
  INV_X1 U8442 ( .A(n12025), .ZN(n8281) );
  AND2_X1 U8443 ( .A1(n11811), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12028) );
  AND2_X1 U8444 ( .A1(n12604), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n12667) );
  NOR2_X1 U8445 ( .A1(n12211), .A2(n12711), .ZN(n12530) );
  NAND2_X1 U8446 ( .A1(n12732), .A2(n12731), .ZN(n12735) );
  NAND2_X1 U8447 ( .A1(n15447), .A2(n15410), .ZN(n8193) );
  NAND2_X1 U8448 ( .A1(n12888), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12902) );
  INV_X1 U8449 ( .A(n12913), .ZN(n12912) );
  INV_X1 U8450 ( .A(n12902), .ZN(n12901) );
  INV_X1 U8451 ( .A(n12895), .ZN(n7467) );
  NOR3_X2 U8452 ( .A1(n12663), .A2(n15711), .A3(n15719), .ZN(n15591) );
  INV_X1 U8453 ( .A(n12614), .ZN(n8199) );
  OR2_X1 U8454 ( .A1(n11450), .A2(n11449), .ZN(n11702) );
  INV_X1 U8455 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11201) );
  INV_X1 U8456 ( .A(n10788), .ZN(n7489) );
  NOR2_X1 U8457 ( .A1(n10692), .A2(n10689), .ZN(n8023) );
  INV_X1 U8458 ( .A(n8472), .ZN(n8091) );
  NAND2_X1 U8459 ( .A1(n15643), .A2(n15410), .ZN(n8092) );
  NAND2_X1 U8460 ( .A1(n11193), .A2(n11192), .ZN(n12770) );
  INV_X1 U8461 ( .A(n8082), .ZN(n8074) );
  AND2_X1 U8462 ( .A1(n7904), .A2(n8573), .ZN(n7903) );
  INV_X1 U8463 ( .A(n8974), .ZN(n7904) );
  NAND2_X1 U8464 ( .A1(n8875), .A2(SI_18_), .ZN(n7892) );
  NOR2_X1 U8465 ( .A1(n8875), .A2(SI_18_), .ZN(n7893) );
  OAI21_X1 U8466 ( .B1(n8536), .B2(n7472), .A(n7296), .ZN(n8762) );
  NAND2_X1 U8467 ( .A1(n7250), .A2(n8538), .ZN(n7472) );
  AND2_X1 U8468 ( .A1(n8377), .A2(n8376), .ZN(n8375) );
  NOR2_X1 U8469 ( .A1(n11426), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U8470 ( .A1(n8536), .A2(n8535), .ZN(n8730) );
  OAI21_X1 U8471 ( .B1(SI_6_), .B2(n7873), .A(n8532), .ZN(n8711) );
  NAND2_X1 U8472 ( .A1(n8508), .A2(n10173), .ZN(n8516) );
  NAND2_X1 U8473 ( .A1(n7561), .A2(n7742), .ZN(n8508) );
  AOI21_X1 U8474 ( .B1(n7697), .B2(n7973), .A(n7696), .ZN(n9176) );
  AND2_X1 U8475 ( .A1(n9127), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7696) );
  INV_X1 U8476 ( .A(n9169), .ZN(n7697) );
  NOR2_X1 U8477 ( .A1(n9131), .A2(n9132), .ZN(n9167) );
  OAI22_X1 U8478 ( .A1(n9138), .A2(n9190), .B1(P3_ADDR_REG_6__SCAN_IN), .B2(
        n9137), .ZN(n9139) );
  INV_X1 U8479 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9137) );
  OAI21_X1 U8480 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n9156), .A(n9155), .ZN(
        n9158) );
  NAND2_X1 U8481 ( .A1(n9352), .A2(n9351), .ZN(n9588) );
  INV_X1 U8482 ( .A(n9572), .ZN(n9352) );
  INV_X1 U8483 ( .A(n7661), .ZN(n7660) );
  XNOR2_X1 U8484 ( .A(n7765), .B(n11640), .ZN(n7670) );
  INV_X1 U8485 ( .A(n13246), .ZN(n9795) );
  NAND2_X1 U8486 ( .A1(n7400), .A2(n13705), .ZN(n9572) );
  INV_X1 U8487 ( .A(n7400), .ZN(n9555) );
  NAND2_X1 U8488 ( .A1(n9354), .A2(n13701), .ZN(n9747) );
  INV_X1 U8489 ( .A(n9735), .ZN(n9354) );
  INV_X1 U8490 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9346) );
  INV_X1 U8491 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11104) );
  NAND2_X1 U8492 ( .A1(n7680), .A2(n7679), .ZN(n7645) );
  INV_X1 U8493 ( .A(n13357), .ZN(n7679) );
  INV_X1 U8494 ( .A(n13358), .ZN(n7680) );
  OR2_X1 U8495 ( .A1(n13514), .A2(n16193), .ZN(n13144) );
  NAND2_X1 U8496 ( .A1(n7391), .A2(n13709), .ZN(n9653) );
  INV_X1 U8497 ( .A(n7394), .ZN(n9671) );
  INV_X1 U8498 ( .A(n7392), .ZN(n9603) );
  AND2_X1 U8499 ( .A1(n13496), .A2(n13492), .ZN(n13337) );
  OAI21_X1 U8500 ( .B1(n7294), .B2(n8043), .A(n7208), .ZN(n8042) );
  INV_X1 U8501 ( .A(n13244), .ZN(n9799) );
  INV_X1 U8502 ( .A(n9407), .ZN(n9796) );
  NAND2_X1 U8503 ( .A1(n13320), .A2(n12397), .ZN(n8420) );
  OR2_X1 U8504 ( .A1(n10567), .A2(n11647), .ZN(n10569) );
  NAND2_X1 U8505 ( .A1(n7935), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7934) );
  NOR2_X1 U8506 ( .A1(n7938), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U8507 ( .A1(n10530), .A2(n8159), .ZN(n10620) );
  NAND2_X1 U8508 ( .A1(n10485), .A2(n10573), .ZN(n10552) );
  OR2_X1 U8509 ( .A1(n10562), .A2(n10561), .ZN(n10551) );
  NAND2_X1 U8510 ( .A1(n10517), .A2(n10529), .ZN(n13753) );
  NAND2_X1 U8511 ( .A1(n7435), .A2(n13746), .ZN(n13749) );
  NAND2_X1 U8512 ( .A1(n10509), .A2(n10508), .ZN(n10511) );
  AND3_X1 U8513 ( .A1(n8163), .A2(n13772), .A3(P3_REG2_REG_5__SCAN_IN), .ZN(
        n13775) );
  OR2_X1 U8514 ( .A1(n13772), .A2(n10671), .ZN(n8162) );
  NOR2_X1 U8515 ( .A1(n10672), .A2(n10659), .ZN(n10804) );
  NAND2_X1 U8516 ( .A1(n10657), .A2(n13763), .ZN(n13766) );
  XNOR2_X1 U8517 ( .A(n11558), .B(n11575), .ZN(n11014) );
  XNOR2_X1 U8518 ( .A(n7757), .B(n11019), .ZN(n11020) );
  OR2_X1 U8519 ( .A1(n11570), .A2(n11571), .ZN(n11956) );
  NAND2_X1 U8520 ( .A1(n11960), .A2(n11959), .ZN(n7754) );
  INV_X1 U8521 ( .A(n7732), .ZN(n11985) );
  INV_X1 U8522 ( .A(n7925), .ZN(n12457) );
  AND2_X1 U8523 ( .A1(n12469), .A2(n12468), .ZN(n12472) );
  INV_X1 U8524 ( .A(n7782), .ZN(n13820) );
  NAND2_X1 U8525 ( .A1(n13844), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7923) );
  XNOR2_X1 U8526 ( .A(n7741), .B(n13868), .ZN(n13836) );
  AOI21_X1 U8527 ( .B1(n7744), .B2(n7933), .A(n7743), .ZN(n7932) );
  INV_X1 U8528 ( .A(n13879), .ZN(n7743) );
  INV_X1 U8529 ( .A(n13882), .ZN(n7931) );
  NAND2_X1 U8530 ( .A1(n13865), .A2(n7358), .ZN(n7929) );
  NAND2_X1 U8531 ( .A1(n13894), .A2(n13893), .ZN(n8175) );
  NAND2_X1 U8532 ( .A1(n7399), .A2(n13712), .ZN(n9735) );
  INV_X1 U8533 ( .A(n7399), .ZN(n9733) );
  OR2_X1 U8534 ( .A1(n9708), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U8535 ( .A1(n7393), .A2(n13419), .ZN(n9708) );
  NAND2_X1 U8536 ( .A1(n7394), .A2(n13586), .ZN(n9682) );
  NAND2_X1 U8537 ( .A1(n7392), .A2(n9353), .ZN(n9621) );
  INV_X1 U8538 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U8539 ( .A1(n8430), .A2(n13332), .ZN(n14104) );
  NAND2_X1 U8540 ( .A1(n9561), .A2(n8427), .ZN(n8430) );
  NAND2_X1 U8541 ( .A1(n9561), .A2(n12552), .ZN(n12637) );
  NOR2_X1 U8542 ( .A1(n8443), .A2(n12357), .ZN(n8442) );
  INV_X1 U8543 ( .A(n9525), .ZN(n8443) );
  AND2_X1 U8544 ( .A1(n13144), .A2(n13145), .ZN(n13273) );
  OR2_X1 U8545 ( .A1(n9512), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9535) );
  AND3_X1 U8546 ( .A1(n7307), .A2(n9509), .A3(n9508), .ZN(n12119) );
  NAND2_X1 U8547 ( .A1(n9350), .A2(n9349), .ZN(n9512) );
  INV_X1 U8548 ( .A(n9495), .ZN(n9350) );
  NAND2_X1 U8549 ( .A1(n9348), .A2(n9347), .ZN(n9478) );
  INV_X1 U8550 ( .A(n9463), .ZN(n9348) );
  OR2_X1 U8551 ( .A1(n9447), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U8552 ( .A1(n13696), .A2(n11104), .ZN(n9434) );
  NAND2_X1 U8553 ( .A1(n16028), .A2(n16031), .ZN(n16027) );
  CLKBUF_X1 U8554 ( .A(n16031), .Z(n7707) );
  NOR2_X1 U8555 ( .A1(n13902), .A2(n13901), .ZN(n14193) );
  OR2_X1 U8556 ( .A1(n9443), .A2(n13640), .ZN(n9745) );
  NAND2_X1 U8557 ( .A1(n9707), .A2(n9706), .ZN(n14151) );
  OR2_X1 U8558 ( .A1(n11042), .A2(n9705), .ZN(n9707) );
  NAND2_X1 U8559 ( .A1(n9692), .A2(n9691), .ZN(n14155) );
  OR2_X1 U8560 ( .A1(n10958), .A2(n9705), .ZN(n9692) );
  AND2_X1 U8561 ( .A1(n14017), .A2(n16163), .ZN(n14182) );
  NAND2_X1 U8562 ( .A1(n7421), .A2(n8460), .ZN(n8459) );
  NOR2_X1 U8563 ( .A1(n7419), .A2(n7677), .ZN(n7418) );
  INV_X1 U8564 ( .A(n8460), .ZN(n7419) );
  NOR2_X1 U8565 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7682) );
  NAND2_X1 U8566 ( .A1(n9759), .A2(n9758), .ZN(n9773) );
  NAND2_X1 U8567 ( .A1(n9316), .A2(n9315), .ZN(n9744) );
  NAND2_X1 U8568 ( .A1(n9374), .A2(n9314), .ZN(n9316) );
  NAND2_X1 U8569 ( .A1(n7984), .A2(n7982), .ZN(n9688) );
  AOI21_X1 U8570 ( .B1(n7985), .B2(n7987), .A(n7983), .ZN(n7982) );
  INV_X1 U8571 ( .A(n9301), .ZN(n7983) );
  XNOR2_X1 U8572 ( .A(n9794), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9851) );
  AND2_X1 U8573 ( .A1(n9299), .A2(n9298), .ZN(n9661) );
  NAND2_X1 U8574 ( .A1(n7991), .A2(n7989), .ZN(n9647) );
  AOI21_X1 U8575 ( .B1(n7992), .B2(n7994), .A(n7990), .ZN(n7989) );
  INV_X1 U8576 ( .A(n9295), .ZN(n7990) );
  AND2_X1 U8577 ( .A1(n9297), .A2(n9296), .ZN(n9646) );
  NAND2_X1 U8578 ( .A1(n7678), .A2(n9330), .ZN(n9634) );
  AND2_X1 U8579 ( .A1(n9293), .A2(n9292), .ZN(n9612) );
  AND2_X1 U8580 ( .A1(n9291), .A2(n9290), .ZN(n9594) );
  NAND2_X1 U8581 ( .A1(n10679), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8007) );
  AND2_X1 U8582 ( .A1(n9289), .A2(n9288), .ZN(n9579) );
  OR2_X1 U8583 ( .A1(n9287), .A2(n10685), .ZN(n8009) );
  NAND2_X1 U8584 ( .A1(n9287), .A2(n10685), .ZN(n8010) );
  NOR2_X1 U8585 ( .A1(n9549), .A2(n7446), .ZN(n7444) );
  NAND2_X1 U8586 ( .A1(n7977), .A2(n7975), .ZN(n9542) );
  AOI21_X1 U8587 ( .B1(n7978), .B2(n7980), .A(n7976), .ZN(n7975) );
  INV_X1 U8588 ( .A(n9284), .ZN(n7976) );
  AND2_X1 U8589 ( .A1(n9286), .A2(n9285), .ZN(n9541) );
  AND2_X1 U8590 ( .A1(n9282), .A2(n9281), .ZN(n9518) );
  NAND2_X1 U8591 ( .A1(n9491), .A2(n9278), .ZN(n9502) );
  OR2_X1 U8592 ( .A1(n9456), .A2(n7446), .ZN(n9440) );
  AND2_X1 U8593 ( .A1(n9266), .A2(n9265), .ZN(n9414) );
  NAND2_X1 U8594 ( .A1(n7859), .A2(n7203), .ZN(n7858) );
  INV_X1 U8595 ( .A(n11505), .ZN(n7859) );
  NAND2_X1 U8596 ( .A1(n11505), .A2(n7856), .ZN(n7852) );
  INV_X1 U8597 ( .A(n7854), .ZN(n7853) );
  XNOR2_X1 U8598 ( .A(n7718), .B(n14352), .ZN(n10981) );
  NOR2_X1 U8599 ( .A1(n14365), .A2(n7871), .ZN(n7870) );
  INV_X1 U8600 ( .A(n14288), .ZN(n7871) );
  NOR2_X1 U8601 ( .A1(n8399), .A2(n7849), .ZN(n7848) );
  INV_X1 U8602 ( .A(n8855), .ZN(n8598) );
  INV_X1 U8603 ( .A(n11089), .ZN(n8397) );
  NAND2_X1 U8604 ( .A1(n14379), .A2(n14378), .ZN(n14377) );
  INV_X1 U8605 ( .A(n14614), .ZN(n14405) );
  NAND2_X1 U8606 ( .A1(n14340), .A2(n8408), .ZN(n14410) );
  INV_X1 U8607 ( .A(n8921), .ZN(n8601) );
  OR2_X1 U8608 ( .A1(n8934), .A2(n8933), .ZN(n8951) );
  INV_X1 U8609 ( .A(n14277), .ZN(n8407) );
  NOR2_X1 U8610 ( .A1(n14450), .A2(n8406), .ZN(n8405) );
  INV_X1 U8611 ( .A(n14266), .ZN(n8406) );
  AND2_X1 U8612 ( .A1(n7905), .A2(n12564), .ZN(n10113) );
  XNOR2_X1 U8613 ( .A(n7906), .B(n9093), .ZN(n7905) );
  XNOR2_X1 U8614 ( .A(n14905), .B(n14463), .ZN(n7907) );
  INV_X1 U8615 ( .A(n10082), .ZN(n10075) );
  AND4_X1 U8616 ( .A1(n8741), .A2(n8740), .A3(n8739), .A4(n8738), .ZN(n11875)
         );
  AND2_X1 U8617 ( .A1(n11230), .A2(n8212), .ZN(n11678) );
  NOR2_X1 U8618 ( .A1(n14905), .A2(n7914), .ZN(n7912) );
  NAND2_X1 U8619 ( .A1(n14581), .A2(n7913), .ZN(n14551) );
  INV_X1 U8620 ( .A(n7914), .ZN(n7913) );
  NAND2_X1 U8621 ( .A1(n9106), .A2(n9105), .ZN(n13086) );
  AND2_X1 U8622 ( .A1(n14581), .A2(n9248), .ZN(n9241) );
  NAND2_X1 U8623 ( .A1(n8602), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8965) );
  INV_X1 U8624 ( .A(n8951), .ZN(n8602) );
  NAND2_X1 U8625 ( .A1(n8603), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8989) );
  INV_X1 U8626 ( .A(n8965), .ZN(n8603) );
  OR2_X1 U8627 ( .A1(n8840), .A2(n14456), .ZN(n8855) );
  NOR2_X1 U8628 ( .A1(n7290), .A2(n7559), .ZN(n7558) );
  INV_X1 U8629 ( .A(n8794), .ZN(n7559) );
  OR2_X1 U8630 ( .A1(n8141), .A2(n7216), .ZN(n8140) );
  NOR2_X2 U8631 ( .A1(n11943), .A2(n11944), .ZN(n12146) );
  NAND2_X1 U8632 ( .A1(n7690), .A2(n8743), .ZN(n11894) );
  OR2_X1 U8633 ( .A1(n11660), .A2(n9036), .ZN(n8135) );
  NAND2_X1 U8634 ( .A1(n8135), .A2(n7236), .ZN(n11938) );
  INV_X1 U8635 ( .A(n12295), .ZN(n11668) );
  NOR2_X1 U8636 ( .A1(n10980), .A2(n11399), .ZN(n11412) );
  NAND2_X1 U8637 ( .A1(n14611), .A2(n7278), .ZN(n7607) );
  INV_X1 U8638 ( .A(n7695), .ZN(n7608) );
  OR2_X1 U8639 ( .A1(n7318), .A2(n7695), .ZN(n7609) );
  NOR2_X1 U8640 ( .A1(n7207), .A2(n9236), .ZN(n8367) );
  AND2_X1 U8641 ( .A1(n9100), .A2(n9023), .ZN(n14351) );
  INV_X1 U8642 ( .A(n9235), .ZN(n7589) );
  AND2_X1 U8643 ( .A1(n14569), .A2(n14580), .ZN(n7714) );
  INV_X1 U8644 ( .A(n7729), .ZN(n7728) );
  OAI21_X1 U8645 ( .B1(n11122), .B2(n10024), .A(n8679), .ZN(n7729) );
  AND2_X1 U8646 ( .A1(n7193), .A2(n12683), .ZN(n16190) );
  INV_X1 U8647 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U8648 ( .A1(n8588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8587) );
  INV_X1 U8649 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U8650 ( .A1(n9068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U8651 ( .A1(n9076), .A2(n9075), .ZN(n9068) );
  NAND2_X1 U8652 ( .A1(n9072), .A2(n9071), .ZN(n9074) );
  INV_X1 U8653 ( .A(n8927), .ZN(n8928) );
  INV_X1 U8654 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8499) );
  OR2_X1 U8655 ( .A1(n7386), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U8656 ( .A1(n8496), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n8497) );
  INV_X1 U8657 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8504) );
  INV_X1 U8658 ( .A(n8415), .ZN(n8413) );
  INV_X1 U8659 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8810) );
  NOR2_X1 U8660 ( .A1(n8675), .A2(n8482), .ZN(n8485) );
  INV_X1 U8661 ( .A(n7803), .ZN(n7813) );
  NAND2_X1 U8662 ( .A1(n14971), .A2(n12998), .ZN(n7469) );
  INV_X1 U8663 ( .A(n8271), .ZN(n8270) );
  NAND2_X1 U8664 ( .A1(n15091), .A2(n15090), .ZN(n7829) );
  OR2_X1 U8665 ( .A1(n8274), .A2(n7828), .ZN(n7827) );
  MUX2_X1 U8666 ( .A(n7251), .B(n10851), .S(n10850), .Z(n10852) );
  AND2_X1 U8667 ( .A1(n8254), .A2(n15038), .ZN(n8253) );
  NAND2_X1 U8668 ( .A1(n15074), .A2(n8255), .ZN(n8254) );
  INV_X1 U8669 ( .A(n15074), .ZN(n8256) );
  OR2_X1 U8670 ( .A1(n10859), .A2(n10860), .ZN(n8265) );
  AOI21_X1 U8671 ( .B1(n8268), .B2(n8270), .A(n8267), .ZN(n8266) );
  INV_X1 U8672 ( .A(n15081), .ZN(n8267) );
  NAND2_X1 U8673 ( .A1(n15016), .A2(n15015), .ZN(n15161) );
  NAND2_X1 U8674 ( .A1(n12028), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n12198) );
  OR3_X1 U8675 ( .A1(n12198), .A2(n12197), .A3(n12196), .ZN(n12211) );
  NAND2_X1 U8676 ( .A1(n12861), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12877) );
  NAND2_X1 U8677 ( .A1(n12370), .A2(n8286), .ZN(n8285) );
  OR2_X1 U8678 ( .A1(n12829), .A2(n15190), .ZN(n12831) );
  NAND2_X1 U8679 ( .A1(n12667), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n12829) );
  OR2_X1 U8680 ( .A1(n15000), .A2(n14999), .ZN(n8273) );
  NAND2_X1 U8681 ( .A1(n12982), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n11135) );
  OR2_X1 U8682 ( .A1(n10199), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n10233) );
  NOR2_X1 U8683 ( .A1(n11288), .A2(n11287), .ZN(n7427) );
  XNOR2_X1 U8684 ( .A(n11736), .B(n11735), .ZN(n11288) );
  NOR2_X1 U8685 ( .A1(n7427), .A2(n7426), .ZN(n11996) );
  NOR2_X1 U8686 ( .A1(n11736), .A2(n11735), .ZN(n7426) );
  AND2_X1 U8687 ( .A1(n12696), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n15330) );
  INV_X1 U8688 ( .A(n7241), .ZN(n8086) );
  OAI21_X1 U8689 ( .B1(n8187), .B2(n8186), .A(n8184), .ZN(n15416) );
  NAND2_X1 U8690 ( .A1(n8192), .A2(n8193), .ZN(n8186) );
  OR2_X1 U8691 ( .A1(n8189), .A2(n8185), .ZN(n8184) );
  INV_X1 U8692 ( .A(n8193), .ZN(n8185) );
  NAND2_X1 U8693 ( .A1(n8019), .A2(n15447), .ZN(n8018) );
  INV_X1 U8694 ( .A(n8090), .ZN(n15379) );
  NOR2_X1 U8695 ( .A1(n15504), .A2(n8017), .ZN(n15457) );
  INV_X1 U8696 ( .A(n8019), .ZN(n8017) );
  NOR2_X1 U8697 ( .A1(n15504), .A2(n8020), .ZN(n15472) );
  NOR2_X1 U8698 ( .A1(n8111), .A2(n8109), .ZN(n8108) );
  INV_X1 U8699 ( .A(n15469), .ZN(n8109) );
  INV_X1 U8700 ( .A(n8027), .ZN(n15539) );
  AND2_X1 U8701 ( .A1(n15549), .A2(n15372), .ZN(n8096) );
  NAND2_X1 U8702 ( .A1(n15566), .A2(n15565), .ZN(n15564) );
  AOI21_X1 U8703 ( .B1(n15604), .B2(n15608), .A(n15368), .ZN(n15587) );
  NAND2_X1 U8704 ( .A1(n15587), .A2(n15586), .ZN(n15585) );
  AOI21_X1 U8705 ( .B1(n13029), .B2(n7253), .A(n8100), .ZN(n8099) );
  NOR2_X1 U8706 ( .A1(n15729), .A2(n12657), .ZN(n8100) );
  INV_X1 U8707 ( .A(n8026), .ZN(n12600) );
  OAI21_X1 U8708 ( .B1(n12163), .B2(n7267), .A(n7542), .ZN(n12345) );
  INV_X1 U8709 ( .A(n7543), .ZN(n7542) );
  OAI21_X1 U8710 ( .B1(n12204), .B2(n7281), .A(n12206), .ZN(n7543) );
  INV_X1 U8711 ( .A(n8071), .ZN(n8070) );
  NAND2_X1 U8712 ( .A1(n12166), .A2(n16172), .ZN(n12165) );
  NAND2_X1 U8713 ( .A1(n8061), .A2(n11700), .ZN(n11809) );
  NAND2_X1 U8714 ( .A1(n11699), .A2(n11698), .ZN(n8061) );
  NAND2_X1 U8715 ( .A1(n7489), .A2(n7488), .ZN(n11358) );
  AND2_X1 U8716 ( .A1(n8021), .A2(n12749), .ZN(n7488) );
  XNOR2_X1 U8717 ( .A(n15235), .B(n12757), .ZN(n12754) );
  INV_X1 U8718 ( .A(n15482), .ZN(n15583) );
  NAND2_X1 U8719 ( .A1(n7489), .A2(n12749), .ZN(n10768) );
  AND4_X1 U8720 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n12741) );
  NAND2_X1 U8721 ( .A1(n10778), .A2(n12746), .ZN(n10782) );
  NAND2_X1 U8722 ( .A1(n10710), .A2(n15343), .ZN(n16002) );
  AOI21_X1 U8723 ( .B1(n15634), .B2(n16151), .A(n15633), .ZN(n8022) );
  NAND2_X1 U8724 ( .A1(n12615), .A2(n12614), .ZN(n12648) );
  NAND2_X1 U8725 ( .A1(n12072), .A2(n12071), .ZN(n12172) );
  INV_X1 U8726 ( .A(n16151), .ZN(n16171) );
  INV_X1 U8728 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10369) );
  XNOR2_X1 U8729 ( .A(n10019), .B(n10018), .ZN(n14958) );
  NAND2_X1 U8730 ( .A1(n7209), .A2(n7552), .ZN(n10368) );
  INV_X1 U8731 ( .A(n10152), .ZN(n7552) );
  NAND2_X1 U8732 ( .A1(n9103), .A2(n9010), .ZN(n13080) );
  XNOR2_X1 U8733 ( .A(n9000), .B(n8581), .ZN(n12940) );
  XNOR2_X1 U8734 ( .A(n10151), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10229) );
  AND2_X1 U8735 ( .A1(n10154), .A2(n7238), .ZN(n10230) );
  NAND2_X1 U8736 ( .A1(n10143), .A2(n10142), .ZN(n10209) );
  INV_X1 U8737 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10142) );
  NAND2_X1 U8738 ( .A1(n8556), .A2(n8373), .ZN(n8849) );
  INV_X1 U8739 ( .A(n7456), .ZN(n8836) );
  AOI21_X1 U8740 ( .B1(n7875), .B2(n7457), .A(n7460), .ZN(n7456) );
  INV_X1 U8741 ( .A(n7461), .ZN(n7457) );
  NAND2_X1 U8742 ( .A1(n7879), .A2(n7881), .ZN(n8808) );
  NAND2_X1 U8743 ( .A1(n7880), .A2(n7884), .ZN(n7879) );
  INV_X1 U8744 ( .A(n8781), .ZN(n7880) );
  OAI21_X1 U8745 ( .B1(n8781), .B2(n8780), .A(n8546), .ZN(n8796) );
  AND2_X1 U8746 ( .A1(n7898), .A2(n7897), .ZN(n8717) );
  XNOR2_X1 U8747 ( .A(n8712), .B(n8711), .ZN(n11315) );
  NAND2_X1 U8748 ( .A1(n8693), .A2(n8530), .ZN(n8712) );
  OAI21_X1 U8749 ( .B1(n8671), .B2(n7564), .A(n7562), .ZN(n8693) );
  INV_X1 U8750 ( .A(n8527), .ZN(n7564) );
  AND2_X1 U8751 ( .A1(n7563), .A2(n8690), .ZN(n7562) );
  NAND2_X1 U8752 ( .A1(n8526), .A2(n8527), .ZN(n7563) );
  NAND2_X1 U8753 ( .A1(n8671), .A2(n8670), .ZN(n8673) );
  OR2_X1 U8754 ( .A1(n10202), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U8755 ( .A1(n8642), .A2(n8521), .ZN(n8139) );
  OAI21_X1 U8756 ( .B1(SI_3_), .B2(n8392), .A(n8523), .ZN(n8522) );
  INV_X1 U8757 ( .A(n7479), .ZN(n7478) );
  OAI21_X1 U8758 ( .B1(n8515), .B2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .ZN(
        n7479) );
  INV_X1 U8759 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9171) );
  NOR2_X1 U8760 ( .A1(n15996), .A2(n9174), .ZN(n9178) );
  AOI22_X1 U8761 ( .A1(n9184), .A2(n9136), .B1(P1_ADDR_REG_5__SCAN_IN), .B2(
        n9135), .ZN(n9190) );
  OR2_X1 U8762 ( .A1(n9135), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n9136) );
  INV_X1 U8763 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9135) );
  OAI21_X1 U8764 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n9144), .A(n9143), .ZN(
        n9202) );
  AOI21_X1 U8765 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n9148), .A(n9147), .ZN(
        n9203) );
  AOI21_X1 U8766 ( .B1(n15936), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n9151), .ZN(
        n9211) );
  AND2_X1 U8767 ( .A1(n9207), .A2(n9206), .ZN(n9151) );
  AND2_X1 U8768 ( .A1(n7960), .A2(n15974), .ZN(n9217) );
  INV_X1 U8769 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U8770 ( .A1(n13329), .A2(n13411), .ZN(n7778) );
  INV_X1 U8771 ( .A(n8355), .ZN(n8354) );
  NAND2_X1 U8772 ( .A1(n9721), .A2(n9720), .ZN(n13392) );
  OR2_X1 U8773 ( .A1(n9443), .A2(n13650), .ZN(n9720) );
  NAND2_X1 U8774 ( .A1(n13398), .A2(n13397), .ZN(n13396) );
  OR2_X1 U8775 ( .A1(n11928), .A2(n11927), .ZN(n7664) );
  OAI21_X1 U8776 ( .B1(n10431), .B2(n7710), .A(n7709), .ZN(n10597) );
  NAND2_X1 U8777 ( .A1(n9405), .A2(n14260), .ZN(n7709) );
  OAI21_X1 U8778 ( .B1(n7670), .B2(n16035), .A(n10638), .ZN(n10600) );
  NAND2_X1 U8779 ( .A1(n13458), .A2(n13351), .ZN(n13417) );
  NAND2_X1 U8780 ( .A1(n8322), .A2(n8325), .ZN(n12623) );
  NAND2_X1 U8781 ( .A1(n12356), .A2(n8327), .ZN(n8322) );
  INV_X1 U8782 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n13701) );
  NAND2_X1 U8783 ( .A1(n13424), .A2(n13425), .ZN(n8333) );
  NAND2_X1 U8784 ( .A1(n13494), .A2(n13339), .ZN(n13434) );
  NAND2_X1 U8785 ( .A1(n11098), .A2(n13522), .ZN(n8341) );
  NAND2_X1 U8786 ( .A1(n7657), .A2(n7661), .ZN(n12124) );
  NAND2_X1 U8787 ( .A1(n11928), .A2(n7662), .ZN(n7657) );
  OAI21_X1 U8788 ( .B1(n13398), .B2(n7653), .A(n7650), .ZN(n13458) );
  NAND2_X1 U8789 ( .A1(n13396), .A2(n13348), .ZN(n13460) );
  NOR2_X1 U8790 ( .A1(n8317), .A2(n7286), .ZN(n8316) );
  INV_X1 U8791 ( .A(n12624), .ZN(n8317) );
  NAND2_X1 U8792 ( .A1(n8315), .A2(n8319), .ZN(n12625) );
  OR2_X1 U8793 ( .A1(n12356), .A2(n8321), .ZN(n8315) );
  INV_X1 U8794 ( .A(n14015), .ZN(n13469) );
  NAND2_X1 U8795 ( .A1(n12356), .A2(n12355), .ZN(n12550) );
  INV_X1 U8796 ( .A(n8340), .ZN(n11792) );
  OAI21_X1 U8797 ( .B1(n13424), .B2(n8337), .A(n8334), .ZN(n13485) );
  NAND2_X1 U8798 ( .A1(n13493), .A2(n13337), .ZN(n13494) );
  INV_X1 U8799 ( .A(n13384), .ZN(n14109) );
  OR2_X1 U8800 ( .A1(n9605), .A2(n10470), .ZN(n9385) );
  OR2_X1 U8801 ( .A1(n13246), .A2(n10523), .ZN(n9388) );
  OR2_X1 U8802 ( .A1(n9412), .A2(n7446), .ZN(n9413) );
  AOI21_X1 U8803 ( .B1(n13778), .B2(n10668), .A(n13779), .ZN(n13783) );
  OAI21_X1 U8804 ( .B1(n10657), .B2(n7409), .A(n7407), .ZN(n10813) );
  INV_X1 U8805 ( .A(n7408), .ZN(n7407) );
  OAI21_X1 U8806 ( .B1(n13763), .B2(n7409), .A(n10663), .ZN(n7408) );
  INV_X1 U8807 ( .A(n10665), .ZN(n7409) );
  NAND2_X1 U8808 ( .A1(n7954), .A2(n7955), .ZN(n10795) );
  NAND2_X1 U8809 ( .A1(n11006), .A2(n11005), .ZN(n11567) );
  INV_X1 U8810 ( .A(n7921), .ZN(n11565) );
  NAND2_X1 U8811 ( .A1(n8173), .A2(n8172), .ZN(n11960) );
  INV_X1 U8812 ( .A(n11579), .ZN(n8172) );
  INV_X1 U8813 ( .A(n8173), .ZN(n11580) );
  NAND2_X1 U8814 ( .A1(n12310), .A2(n12309), .ZN(n12313) );
  INV_X1 U8815 ( .A(n7699), .ZN(n13793) );
  XNOR2_X1 U8816 ( .A(n7922), .B(n13868), .ZN(n13833) );
  NOR2_X1 U8817 ( .A1(n13833), .A2(n13834), .ZN(n13858) );
  AND2_X1 U8818 ( .A1(n13871), .A2(n13870), .ZN(n7797) );
  INV_X1 U8819 ( .A(n7701), .ZN(n7700) );
  AOI21_X1 U8820 ( .B1(n13874), .B2(n13884), .A(n7702), .ZN(n7701) );
  NAND2_X1 U8821 ( .A1(n13872), .A2(n13873), .ZN(n7702) );
  INV_X1 U8822 ( .A(n8048), .ZN(n8046) );
  NAND2_X1 U8823 ( .A1(n7628), .A2(n7626), .ZN(n13914) );
  AND2_X1 U8824 ( .A1(n7627), .A2(n13207), .ZN(n7626) );
  NAND2_X1 U8825 ( .A1(n13980), .A2(n7280), .ZN(n7628) );
  AOI22_X1 U8826 ( .A1(n13929), .A2(n13930), .B1(n8448), .B2(n8447), .ZN(
        n13931) );
  NAND2_X1 U8827 ( .A1(n8448), .A2(n8449), .ZN(n13929) );
  NAND2_X1 U8828 ( .A1(n13951), .A2(n8452), .ZN(n8448) );
  NAND2_X1 U8829 ( .A1(n7630), .A2(n8030), .ZN(n13939) );
  NAND2_X1 U8830 ( .A1(n13980), .A2(n8031), .ZN(n7630) );
  NAND2_X1 U8831 ( .A1(n8032), .A2(n8033), .ZN(n13949) );
  OR2_X1 U8832 ( .A1(n13980), .A2(n8034), .ZN(n8032) );
  NAND2_X1 U8833 ( .A1(n14147), .A2(n13200), .ZN(n13970) );
  AND2_X1 U8834 ( .A1(n14014), .A2(n13189), .ZN(n8463) );
  NAND2_X1 U8835 ( .A1(n8433), .A2(n8437), .ZN(n14000) );
  NAND2_X1 U8836 ( .A1(n14026), .A2(n7242), .ZN(n8433) );
  OAI21_X1 U8837 ( .B1(n14026), .B2(n7244), .A(n9675), .ZN(n14010) );
  NAND2_X1 U8838 ( .A1(n9670), .A2(n9669), .ZN(n14039) );
  OR2_X1 U8839 ( .A1(n10648), .A2(n9705), .ZN(n9670) );
  NAND2_X1 U8840 ( .A1(n9652), .A2(n9651), .ZN(n14169) );
  OR2_X1 U8841 ( .A1(n10609), .A2(n9705), .ZN(n9652) );
  NAND2_X1 U8842 ( .A1(n9812), .A2(n13173), .ZN(n14042) );
  AND2_X1 U8843 ( .A1(n8457), .A2(n13171), .ZN(n14057) );
  NAND2_X1 U8844 ( .A1(n14084), .A2(n9611), .ZN(n14073) );
  INV_X1 U8845 ( .A(n8457), .ZN(n14072) );
  NAND2_X1 U8846 ( .A1(n14092), .A2(n13164), .ZN(n14071) );
  NAND2_X1 U8847 ( .A1(n9586), .A2(n9585), .ZN(n16223) );
  OR2_X1 U8848 ( .A1(n10221), .A2(n9705), .ZN(n9554) );
  INV_X1 U8849 ( .A(n12366), .ZN(n16193) );
  NAND2_X1 U8850 ( .A1(n8038), .A2(n8039), .ZN(n12251) );
  INV_X1 U8851 ( .A(n12119), .ZN(n16142) );
  NAND2_X1 U8852 ( .A1(n12100), .A2(n9809), .ZN(n12153) );
  NAND2_X1 U8853 ( .A1(n11621), .A2(n9477), .ZN(n12104) );
  NAND2_X1 U8854 ( .A1(n11030), .A2(n9433), .ZN(n11481) );
  INV_X1 U8855 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n13696) );
  NAND2_X1 U8856 ( .A1(n8461), .A2(n9406), .ZN(n11631) );
  NAND2_X1 U8857 ( .A1(n11063), .A2(n11062), .ZN(n16126) );
  NAND2_X1 U8858 ( .A1(n13243), .A2(n13242), .ZN(n14119) );
  AND2_X1 U8859 ( .A1(n9732), .A2(n9731), .ZN(n14218) );
  INV_X1 U8860 ( .A(n13392), .ZN(n14222) );
  NAND2_X1 U8861 ( .A1(n9602), .A2(n9601), .ZN(n14242) );
  AND3_X1 U8862 ( .A1(n9461), .A2(n9460), .A3(n9459), .ZN(n11746) );
  INV_X1 U8863 ( .A(n10597), .ZN(n11064) );
  AND2_X1 U8864 ( .A1(n9833), .A2(n9832), .ZN(n14248) );
  NAND2_X1 U8865 ( .A1(n10432), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14249) );
  NAND3_X1 U8866 ( .A1(n7678), .A2(n7676), .A3(n7675), .ZN(n14255) );
  AND2_X1 U8867 ( .A1(n8056), .A2(n7326), .ZN(n7676) );
  INV_X1 U8868 ( .A(n8459), .ZN(n7675) );
  NAND2_X1 U8869 ( .A1(n9826), .A2(n9827), .ZN(n11731) );
  MUX2_X1 U8870 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9824), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9826) );
  MUX2_X1 U8871 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9789), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9790) );
  INV_X1 U8872 ( .A(n9851), .ZN(n10775) );
  NAND2_X1 U8873 ( .A1(n7981), .A2(n7985), .ZN(n9679) );
  OR2_X1 U8874 ( .A1(n9662), .A2(n7987), .ZN(n7981) );
  INV_X1 U8875 ( .A(n13881), .ZN(n13888) );
  NAND2_X1 U8876 ( .A1(n7988), .A2(n7992), .ZN(n9631) );
  OR2_X1 U8877 ( .A1(n9613), .A2(n7994), .ZN(n7988) );
  INV_X1 U8878 ( .A(n13823), .ZN(n13844) );
  INV_X1 U8879 ( .A(SI_15_), .ZN(n13659) );
  NOR2_X1 U8880 ( .A1(n9567), .A2(n7446), .ZN(n7445) );
  INV_X1 U8881 ( .A(SI_12_), .ZN(n10222) );
  INV_X1 U8882 ( .A(SI_11_), .ZN(n13666) );
  OR2_X1 U8883 ( .A1(n9546), .A2(n7446), .ZN(n9530) );
  NAND2_X1 U8884 ( .A1(n7974), .A2(n7978), .ZN(n9529) );
  OR2_X1 U8885 ( .A1(n9519), .A2(n7980), .ZN(n7974) );
  NAND2_X1 U8886 ( .A1(n9474), .A2(n9276), .ZN(n9489) );
  NOR2_X1 U8887 ( .A1(n9484), .A2(n7446), .ZN(n7443) );
  NAND2_X1 U8888 ( .A1(n9274), .A2(n9273), .ZN(n9472) );
  NAND2_X1 U8889 ( .A1(n7998), .A2(n9269), .ZN(n9442) );
  NAND2_X1 U8890 ( .A1(n9430), .A2(n9429), .ZN(n7998) );
  INV_X1 U8891 ( .A(n10522), .ZN(n10559) );
  INV_X1 U8892 ( .A(n9259), .ZN(n9377) );
  NAND2_X1 U8893 ( .A1(n7731), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9380) );
  NAND2_X1 U8894 ( .A1(n7858), .A2(n7856), .ZN(n11880) );
  AND2_X1 U8895 ( .A1(n8997), .A2(n8996), .ZN(n14599) );
  NOR2_X1 U8896 ( .A1(n14315), .A2(n8411), .ZN(n8410) );
  INV_X1 U8897 ( .A(n14311), .ZN(n8411) );
  NAND2_X1 U8898 ( .A1(n14442), .A2(n14311), .ZN(n14314) );
  NAND2_X1 U8899 ( .A1(n8827), .A2(n8826), .ZN(n14889) );
  NAND2_X1 U8900 ( .A1(n14335), .A2(n14334), .ZN(n14333) );
  NAND2_X1 U8901 ( .A1(n12229), .A2(n12230), .ZN(n12268) );
  NAND2_X1 U8902 ( .A1(n12228), .A2(n12227), .ZN(n12229) );
  AND4_X1 U8903 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n12038)
         );
  NAND2_X1 U8904 ( .A1(n14410), .A2(n14288), .ZN(n14364) );
  AND4_X1 U8905 ( .A1(n8792), .A2(n8791), .A3(n8790), .A4(n8789), .ZN(n12499)
         );
  NAND2_X1 U8906 ( .A1(n8977), .A2(n8976), .ZN(n14601) );
  NAND2_X1 U8907 ( .A1(n14377), .A2(n14273), .ZN(n14389) );
  NAND2_X1 U8908 ( .A1(n14333), .A2(n14299), .ZN(n14400) );
  NOR2_X1 U8909 ( .A1(n11090), .A2(n11089), .ZN(n11255) );
  NAND2_X1 U8910 ( .A1(n14340), .A2(n14284), .ZN(n14412) );
  NAND2_X1 U8911 ( .A1(n12568), .A2(n12567), .ZN(n14262) );
  AOI21_X1 U8912 ( .B1(n12230), .B2(n12226), .A(n12267), .ZN(n8401) );
  NAND2_X1 U8913 ( .A1(n12044), .A2(n8400), .ZN(n7846) );
  AND2_X1 U8914 ( .A1(n12045), .A2(n12230), .ZN(n8400) );
  OAI21_X2 U8915 ( .B1(n10839), .B2(n11550), .A(n14697), .ZN(n14423) );
  INV_X1 U8916 ( .A(n14713), .ZN(n14861) );
  NAND2_X1 U8917 ( .A1(n14388), .A2(n14277), .ZN(n14429) );
  NOR2_X1 U8918 ( .A1(n11505), .A2(n11504), .ZN(n11677) );
  NAND2_X1 U8919 ( .A1(n11091), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14403) );
  INV_X1 U8920 ( .A(n14449), .ZN(n14420) );
  NAND2_X1 U8921 ( .A1(n14324), .A2(n14266), .ZN(n14451) );
  INV_X1 U8922 ( .A(n14599), .ZN(n14466) );
  INV_X1 U8923 ( .A(n11679), .ZN(n14478) );
  NAND4_X1 U8924 ( .A1(n8669), .A2(n8668), .A3(n8667), .A4(n8666), .ZN(n14481)
         );
  NAND2_X1 U8925 ( .A1(n7587), .A2(n7585), .ZN(n9108) );
  INV_X1 U8926 ( .A(n7586), .ZN(n7585) );
  NAND2_X1 U8927 ( .A1(n9233), .A2(n7588), .ZN(n7587) );
  NAND2_X1 U8928 ( .A1(n7572), .A2(n7575), .ZN(n14586) );
  OR2_X1 U8929 ( .A1(n14610), .A2(n7577), .ZN(n7572) );
  AND2_X1 U8930 ( .A1(n8986), .A2(n8985), .ZN(n14584) );
  INV_X1 U8931 ( .A(n7692), .ZN(n7691) );
  NAND2_X1 U8932 ( .A1(n14579), .A2(n14578), .ZN(n7693) );
  AOI22_X1 U8933 ( .A1(n14580), .A2(n14791), .B1(n14647), .B2(n14614), .ZN(
        n7692) );
  NAND2_X1 U8934 ( .A1(n7580), .A2(n8973), .ZN(n14592) );
  NAND2_X1 U8935 ( .A1(n14610), .A2(n14613), .ZN(n7580) );
  NAND2_X1 U8936 ( .A1(n8385), .A2(n8949), .ZN(n14641) );
  NAND2_X1 U8937 ( .A1(n14971), .A2(n10044), .ZN(n8385) );
  AND2_X1 U8938 ( .A1(n8932), .A2(n8931), .ZN(n14654) );
  NAND2_X1 U8939 ( .A1(n7599), .A2(n7597), .ZN(n14645) );
  INV_X1 U8940 ( .A(n7598), .ZN(n7597) );
  AOI21_X1 U8941 ( .B1(n14682), .B2(n14681), .A(n9052), .ZN(n14668) );
  NAND2_X1 U8942 ( .A1(n8152), .A2(n8903), .ZN(n14675) );
  NAND2_X1 U8943 ( .A1(n8121), .A2(n8127), .ZN(n14689) );
  NAND2_X1 U8944 ( .A1(n14722), .A2(n8124), .ZN(n8121) );
  NAND2_X1 U8945 ( .A1(n14722), .A2(n9049), .ZN(n14704) );
  AND2_X1 U8946 ( .A1(n8866), .A2(n8865), .ZN(n14728) );
  AND2_X1 U8947 ( .A1(n8149), .A2(n7256), .ZN(n12327) );
  NAND2_X1 U8948 ( .A1(n8760), .A2(n8759), .ZN(n12139) );
  NAND2_X1 U8949 ( .A1(n7595), .A2(n9034), .ZN(n11495) );
  NAND2_X1 U8950 ( .A1(n11406), .A2(n9028), .ZN(n10995) );
  NAND2_X1 U8951 ( .A1(n9027), .A2(n11392), .ZN(n11408) );
  NAND2_X1 U8952 ( .A1(n8656), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8646) );
  INV_X1 U8953 ( .A(n16085), .ZN(n14747) );
  OR2_X1 U8954 ( .A1(n16094), .A2(n11550), .ZN(n16085) );
  NAND2_X1 U8955 ( .A1(n16206), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7721) );
  OR2_X1 U8956 ( .A1(n16208), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8137) );
  INV_X1 U8957 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U8958 ( .A1(n14811), .A2(n14813), .ZN(n14901) );
  INV_X1 U8959 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n7788) );
  INV_X1 U8960 ( .A(n14641), .ZN(n14914) );
  AND2_X1 U8961 ( .A1(n8908), .A2(n8907), .ZN(n14929) );
  NAND2_X1 U8962 ( .A1(n8147), .A2(n8847), .ZN(n14741) );
  OR3_X1 U8963 ( .A1(n14882), .A2(n14881), .A3(n14880), .ZN(n14883) );
  NAND2_X1 U8964 ( .A1(n8142), .A2(n8141), .ZN(n14785) );
  AND2_X1 U8965 ( .A1(n8142), .A2(n8806), .ZN(n14787) );
  NAND2_X1 U8966 ( .A1(n8144), .A2(n8143), .ZN(n8142) );
  AND2_X1 U8967 ( .A1(n8785), .A2(n8784), .ZN(n12425) );
  INV_X1 U8968 ( .A(n11944), .ZN(n12289) );
  NAND2_X1 U8969 ( .A1(n11662), .A2(n11661), .ZN(n11664) );
  NAND2_X1 U8970 ( .A1(n7583), .A2(n7767), .ZN(n11662) );
  AND2_X1 U8971 ( .A1(n10895), .A2(n9082), .ZN(n15821) );
  AND2_X1 U8972 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10827), .ZN(n9082) );
  OAI21_X1 U8973 ( .B1(n9097), .B2(P2_D_REG_0__SCAN_IN), .A(n9096), .ZN(n15820) );
  NAND2_X1 U8974 ( .A1(n7750), .A2(n7217), .ZN(n7726) );
  NOR2_X1 U8975 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n7724) );
  XNOR2_X1 U8976 ( .A(n9070), .B(n9069), .ZN(n14965) );
  NAND2_X1 U8977 ( .A1(n9074), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U8978 ( .A1(n9074), .A2(n9073), .ZN(n14967) );
  OR2_X1 U8979 ( .A1(n9072), .A2(n9071), .ZN(n9073) );
  XNOR2_X1 U8980 ( .A(n9076), .B(n9075), .ZN(n12688) );
  INV_X1 U8981 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10824) );
  INV_X1 U8982 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10635) );
  INV_X1 U8983 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10471) );
  INV_X1 U8984 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10367) );
  INV_X1 U8985 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10243) );
  INV_X1 U8986 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10237) );
  INV_X1 U8987 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10224) );
  INV_X1 U8988 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10183) );
  INV_X1 U8989 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10179) );
  INV_X1 U8990 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10157) );
  NAND2_X1 U8991 ( .A1(n7814), .A2(n7813), .ZN(n11775) );
  NAND2_X1 U8992 ( .A1(n15169), .A2(n15031), .ZN(n15073) );
  AOI21_X1 U8993 ( .B1(n12020), .B2(n12019), .A(n7841), .ZN(n12026) );
  NAND2_X1 U8994 ( .A1(n12026), .A2(n12025), .ZN(n12371) );
  INV_X1 U8995 ( .A(n8265), .ZN(n11128) );
  NAND2_X1 U8996 ( .A1(n7810), .A2(n7809), .ZN(n11784) );
  OR2_X1 U8997 ( .A1(n11774), .A2(n7816), .ZN(n7809) );
  NAND2_X1 U8998 ( .A1(n7814), .A2(n7353), .ZN(n7810) );
  NAND2_X1 U8999 ( .A1(n15161), .A2(n15020), .ZN(n15115) );
  NAND2_X1 U9000 ( .A1(n7838), .A2(n7836), .ZN(n12583) );
  AOI21_X1 U9001 ( .B1(n8264), .B2(n10860), .A(n11189), .ZN(n8258) );
  NAND2_X1 U9002 ( .A1(n10859), .A2(n8264), .ZN(n8259) );
  NAND2_X1 U9003 ( .A1(n12909), .A2(n12908), .ZN(n15662) );
  NAND2_X1 U9004 ( .A1(n12850), .A2(n12849), .ZN(n15688) );
  INV_X1 U9005 ( .A(n7834), .ZN(n7832) );
  AND2_X1 U9006 ( .A1(n12587), .A2(n7842), .ZN(n7833) );
  OAI21_X1 U9007 ( .B1(n7831), .B2(n7830), .A(n7834), .ZN(n12588) );
  NAND2_X1 U9008 ( .A1(n7836), .A2(n7842), .ZN(n7830) );
  INV_X1 U9009 ( .A(n7838), .ZN(n7831) );
  NAND2_X1 U9010 ( .A1(n12371), .A2(n8285), .ZN(n12373) );
  AOI21_X1 U9011 ( .B1(n11314), .B2(n11313), .A(n11312), .ZN(n11441) );
  NAND2_X1 U9012 ( .A1(n8276), .A2(n15054), .ZN(n15199) );
  NAND2_X1 U9013 ( .A1(n15123), .A2(n15124), .ZN(n8276) );
  AND2_X1 U9014 ( .A1(n10411), .A2(n15615), .ZN(n15220) );
  INV_X1 U9015 ( .A(n10864), .ZN(n15236) );
  NAND2_X1 U9016 ( .A1(n10761), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n10413) );
  OR2_X2 U9017 ( .A1(n10231), .A2(n8287), .ZN(n15237) );
  NAND2_X1 U9018 ( .A1(n15260), .A2(n15261), .ZN(n15259) );
  XNOR2_X1 U9019 ( .A(n15255), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n15261) );
  NAND2_X1 U9020 ( .A1(n10312), .A2(n7273), .ZN(n10313) );
  OAI21_X1 U9021 ( .B1(n15926), .B2(n15921), .A(n10941), .ZN(n15924) );
  NOR2_X1 U9022 ( .A1(n10579), .A2(n10580), .ZN(n15926) );
  NAND2_X1 U9023 ( .A1(n15924), .A2(n7422), .ZN(n10942) );
  OR2_X1 U9024 ( .A1(n15930), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7422) );
  INV_X1 U9025 ( .A(n7427), .ZN(n11734) );
  NOR2_X1 U9026 ( .A1(n15329), .A2(n7424), .ZN(n12696) );
  AND2_X1 U9027 ( .A1(n12694), .A2(n12699), .ZN(n7424) );
  XNOR2_X1 U9028 ( .A(n7423), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n15342) );
  NOR2_X1 U9029 ( .A1(n15330), .A2(n15329), .ZN(n7423) );
  AOI211_X1 U9030 ( .C1(n15423), .C2(n15634), .A(n16096), .B(n15383), .ZN(
        n15632) );
  NAND2_X1 U9031 ( .A1(n8190), .A2(n8188), .ZN(n15435) );
  INV_X1 U9032 ( .A(n15643), .ZN(n15447) );
  NAND2_X1 U9033 ( .A1(n8115), .A2(n8464), .ZN(n15486) );
  NAND2_X1 U9034 ( .A1(n15520), .A2(n15405), .ZN(n15510) );
  NAND2_X1 U9035 ( .A1(n12872), .A2(n12871), .ZN(n15679) );
  NAND2_X1 U9036 ( .A1(n15564), .A2(n8096), .ZN(n15692) );
  NAND2_X1 U9037 ( .A1(n15561), .A2(n8196), .ZN(n15546) );
  AND2_X1 U9038 ( .A1(n15561), .A2(n15399), .ZN(n15548) );
  NAND2_X1 U9039 ( .A1(n12729), .A2(n12728), .ZN(n15698) );
  NAND2_X1 U9040 ( .A1(n15605), .A2(n15396), .ZN(n15580) );
  INV_X1 U9041 ( .A(n15705), .ZN(n15597) );
  NAND2_X1 U9042 ( .A1(n15395), .A2(n15394), .ZN(n15607) );
  OR2_X1 U9043 ( .A1(n12518), .A2(n8104), .ZN(n8098) );
  NAND2_X1 U9044 ( .A1(n12525), .A2(n12524), .ZN(n12527) );
  NAND2_X1 U9045 ( .A1(n8107), .A2(n12519), .ZN(n12603) );
  NAND2_X1 U9046 ( .A1(n12518), .A2(n12517), .ZN(n8107) );
  NAND2_X1 U9047 ( .A1(n7541), .A2(n12088), .ZN(n12205) );
  NAND2_X1 U9048 ( .A1(n12163), .A2(n12171), .ZN(n7541) );
  AND2_X1 U9049 ( .A1(n8181), .A2(n8179), .ZN(n11336) );
  NAND2_X1 U9050 ( .A1(n11235), .A2(n11234), .ZN(n11356) );
  OR2_X1 U9051 ( .A1(n16022), .A2(n12168), .ZN(n15577) );
  OR2_X1 U9052 ( .A1(n10417), .A2(n10686), .ZN(n15615) );
  NAND2_X1 U9053 ( .A1(n10706), .A2(n10718), .ZN(n10747) );
  OR2_X1 U9054 ( .A1(n16022), .A2(n11046), .ZN(n16014) );
  NAND2_X1 U9055 ( .A1(n8069), .A2(n8068), .ZN(n7483) );
  INV_X1 U9056 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U9057 ( .A1(n15422), .A2(n7473), .ZN(n15743) );
  AND2_X1 U9058 ( .A1(n15642), .A2(n15421), .ZN(n7473) );
  INV_X1 U9059 ( .A(n10421), .ZN(n10145) );
  NAND2_X1 U9060 ( .A1(n8084), .A2(n7198), .ZN(n15759) );
  XNOR2_X1 U9061 ( .A(n10043), .B(n10042), .ZN(n15758) );
  NAND2_X1 U9062 ( .A1(n10040), .A2(n7894), .ZN(n13079) );
  INV_X1 U9063 ( .A(n7896), .ZN(n7895) );
  OAI21_X1 U9064 ( .B1(n10018), .B2(n7230), .A(n10022), .ZN(n7896) );
  INV_X1 U9065 ( .A(n10372), .ZN(n15764) );
  OAI21_X1 U9066 ( .B1(n10152), .B2(n7204), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8210) );
  XNOR2_X1 U9067 ( .A(n10155), .B(P1_IR_REG_24__SCAN_IN), .ZN(n12685) );
  XNOR2_X1 U9068 ( .A(n12883), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15778) );
  INV_X1 U9069 ( .A(n12731), .ZN(n12992) );
  NAND2_X1 U9070 ( .A1(n7245), .A2(n8384), .ZN(n8879) );
  INV_X1 U9071 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11435) );
  INV_X1 U9072 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11186) );
  INV_X1 U9073 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10822) );
  INV_X1 U9074 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10633) );
  INV_X1 U9075 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10476) );
  INV_X1 U9076 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10365) );
  NAND2_X1 U9077 ( .A1(n8378), .A2(n8382), .ZN(n8748) );
  AND2_X1 U9078 ( .A1(n8380), .A2(n8379), .ZN(n8378) );
  INV_X1 U9079 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10241) );
  INV_X1 U9080 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10235) );
  INV_X1 U9081 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10195) );
  NAND2_X1 U9082 ( .A1(n8673), .A2(n8672), .ZN(n11122) );
  OR2_X1 U9083 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  XNOR2_X1 U9084 ( .A(n7425), .B(n10197), .ZN(n15255) );
  NAND2_X1 U9085 ( .A1(n10196), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7425) );
  XNOR2_X1 U9086 ( .A(n9172), .B(n9173), .ZN(n15997) );
  NOR2_X1 U9087 ( .A1(n15997), .A2(n15998), .ZN(n15996) );
  INV_X1 U9088 ( .A(n7965), .ZN(n9198) );
  OAI21_X1 U9089 ( .B1(n7439), .B2(n7438), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n7437) );
  NAND2_X1 U9090 ( .A1(n15967), .A2(n9210), .ZN(n15972) );
  NOR2_X1 U9091 ( .A1(n15972), .A2(n15971), .ZN(n9213) );
  NAND2_X1 U9092 ( .A1(n15976), .A2(n15975), .ZN(n15974) );
  NOR2_X1 U9093 ( .A1(n9217), .A2(n9216), .ZN(n15979) );
  NAND2_X1 U9094 ( .A1(n15980), .A2(n15978), .ZN(n15985) );
  NAND2_X1 U9095 ( .A1(n15985), .A2(n15984), .ZN(n15983) );
  NAND2_X1 U9096 ( .A1(n7448), .A2(n15983), .ZN(n15988) );
  OAI21_X1 U9097 ( .B1(n15985), .B2(n15984), .A(n7959), .ZN(n7448) );
  INV_X1 U9098 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7959) );
  NOR2_X1 U9099 ( .A1(n14249), .A2(n10446), .ZN(P3_U3897) );
  NAND2_X1 U9100 ( .A1(n8350), .A2(n13495), .ZN(n8347) );
  INV_X1 U9101 ( .A(n7669), .ZN(n10642) );
  NOR2_X1 U9102 ( .A1(n7390), .A2(n7388), .ZN(n13316) );
  INV_X1 U9103 ( .A(n8165), .ZN(n12456) );
  INV_X1 U9104 ( .A(n7924), .ZN(n13832) );
  NAND2_X1 U9105 ( .A1(n8176), .A2(n13838), .ZN(n7740) );
  NOR2_X1 U9106 ( .A1(n7413), .A2(n7414), .ZN(n7415) );
  NAND2_X1 U9107 ( .A1(n7687), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7685) );
  OR2_X1 U9108 ( .A1(n16232), .A2(n9860), .ZN(n7688) );
  NAND2_X1 U9109 ( .A1(n8236), .A2(n14972), .ZN(n8234) );
  NAND2_X1 U9110 ( .A1(n10124), .A2(n8233), .ZN(n8232) );
  AOI21_X1 U9111 ( .B1(n14564), .B2(n14623), .A(n7748), .ZN(n14565) );
  OAI21_X1 U9112 ( .B1(n14559), .B2(n16062), .A(n7749), .ZN(n7748) );
  NAND2_X1 U9113 ( .A1(n7722), .A2(n7719), .ZN(P2_U3530) );
  INV_X1 U9114 ( .A(n7720), .ZN(n7719) );
  NAND2_X1 U9115 ( .A1(n14901), .A2(n16208), .ZN(n7722) );
  OAI21_X1 U9116 ( .B1(n14812), .B2(n14896), .A(n7721), .ZN(n7720) );
  OAI211_X1 U9117 ( .C1(n14557), .C2(n16206), .A(n8388), .B(n8386), .ZN(
        P2_U3527) );
  AND2_X1 U9118 ( .A1(n8389), .A2(n7341), .ZN(n8388) );
  OR2_X1 U9119 ( .A1(n14559), .A2(n8387), .ZN(n8386) );
  NAND2_X1 U9120 ( .A1(n7919), .A2(n7916), .ZN(P2_U3498) );
  AOI21_X1 U9121 ( .B1(n14902), .B2(n14906), .A(n7917), .ZN(n7916) );
  NAND2_X1 U9122 ( .A1(n14901), .A2(n14948), .ZN(n7919) );
  NOR2_X1 U9123 ( .A1(n14948), .A2(n7918), .ZN(n7917) );
  OR2_X1 U9124 ( .A1(n14948), .A2(n7769), .ZN(n7768) );
  INV_X1 U9125 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U9126 ( .A1(n8156), .A2(n8155), .ZN(n9252) );
  OR2_X1 U9127 ( .A1(n14948), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8155) );
  NOR2_X1 U9128 ( .A1(n9250), .A2(n7787), .ZN(n7786) );
  NOR2_X1 U9129 ( .A1(n14948), .A2(n7788), .ZN(n7787) );
  NAND2_X1 U9130 ( .A1(n7821), .A2(n15210), .ZN(n7819) );
  NAND2_X1 U9131 ( .A1(n7482), .A2(n7480), .ZN(P1_U3557) );
  OR2_X1 U9132 ( .A1(n16179), .A2(n7481), .ZN(n7480) );
  NAND2_X1 U9133 ( .A1(n7483), .A2(n16179), .ZN(n7482) );
  INV_X1 U9134 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7481) );
  OAI21_X1 U9135 ( .B1(n8068), .B2(n16180), .A(n7705), .ZN(P1_U3525) );
  INV_X1 U9136 ( .A(n7706), .ZN(n7705) );
  OR2_X1 U9137 ( .A1(n16183), .A2(n8067), .ZN(n8066) );
  NAND2_X1 U9138 ( .A1(n7476), .A2(n7474), .ZN(P1_U3524) );
  OR2_X1 U9139 ( .A1(n16183), .A2(n7475), .ZN(n7474) );
  NAND2_X1 U9140 ( .A1(n15743), .A2(n16183), .ZN(n7476) );
  INV_X1 U9141 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7475) );
  INV_X1 U9142 ( .A(n7966), .ZN(n7967) );
  NAND2_X1 U9143 ( .A1(n7970), .A2(n7775), .ZN(n7774) );
  XNOR2_X1 U9144 ( .A(n9232), .B(n7360), .ZN(n7968) );
  AND2_X1 U9145 ( .A1(n9809), .A2(n8040), .ZN(n7195) );
  INV_X1 U9146 ( .A(n15498), .ZN(n15509) );
  AND2_X1 U9147 ( .A1(n12886), .A2(n7504), .ZN(n7196) );
  AND2_X1 U9148 ( .A1(n8126), .A2(n14468), .ZN(n7197) );
  INV_X1 U9149 ( .A(n15565), .ZN(n8094) );
  AND2_X1 U9150 ( .A1(n10369), .A2(n10218), .ZN(n7198) );
  INV_X1 U9151 ( .A(n9994), .ZN(n7370) );
  AND2_X1 U9152 ( .A1(n8056), .A2(n7302), .ZN(n7199) );
  AND2_X1 U9153 ( .A1(n8354), .A2(n13449), .ZN(n7200) );
  INV_X1 U9154 ( .A(n10108), .ZN(n8154) );
  INV_X1 U9155 ( .A(n9983), .ZN(n8224) );
  NAND2_X1 U9156 ( .A1(n14581), .A2(n7915), .ZN(n7201) );
  OR2_X1 U9157 ( .A1(n13442), .A2(n13441), .ZN(n7202) );
  AND2_X1 U9158 ( .A1(n11676), .A2(n11503), .ZN(n7203) );
  AND2_X1 U9159 ( .A1(n7304), .A2(n7512), .ZN(n7205) );
  OR2_X1 U9160 ( .A1(n13369), .A2(n13953), .ZN(n13205) );
  AND2_X1 U9161 ( .A1(n8016), .A2(n8015), .ZN(n7206) );
  AND2_X1 U9162 ( .A1(n14569), .A2(n9054), .ZN(n7207) );
  NOR2_X1 U9163 ( .A1(n9094), .A2(n12564), .ZN(n10976) );
  NAND2_X1 U9164 ( .A1(n12121), .A2(n13517), .ZN(n8338) );
  NAND2_X1 U9165 ( .A1(n7873), .A2(SI_6_), .ZN(n8532) );
  AND2_X1 U9166 ( .A1(n13287), .A2(n13302), .ZN(n7208) );
  NOR2_X1 U9167 ( .A1(n7204), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U9168 ( .A1(n8895), .A2(n8894), .ZN(n14700) );
  INV_X1 U9169 ( .A(n14700), .ZN(n8126) );
  INV_X1 U9170 ( .A(n14399), .ZN(n8399) );
  AND2_X1 U9171 ( .A1(n8539), .A2(n8381), .ZN(n7210) );
  OR2_X1 U9172 ( .A1(n14179), .A2(n14088), .ZN(n13171) );
  INV_X1 U9173 ( .A(n9754), .ZN(n8452) );
  OAI211_X1 U9174 ( .C1(n7469), .C2(n15406), .A(n7465), .B(n7464), .ZN(n15498)
         );
  AND2_X1 U9175 ( .A1(n7727), .A2(n8586), .ZN(n7211) );
  AND2_X1 U9176 ( .A1(n7387), .A2(n9753), .ZN(n13953) );
  INV_X1 U9177 ( .A(n13953), .ZN(n13510) );
  AND2_X1 U9178 ( .A1(n14291), .A2(n14290), .ZN(n7212) );
  INV_X1 U9179 ( .A(n12898), .ZN(n7501) );
  INV_X1 U9180 ( .A(n14560), .ZN(n9251) );
  NAND2_X1 U9181 ( .A1(n9012), .A2(n9011), .ZN(n14560) );
  OR2_X1 U9182 ( .A1(n13077), .A2(n13076), .ZN(n7213) );
  AND2_X1 U9183 ( .A1(n7350), .A2(n12567), .ZN(n7214) );
  INV_X1 U9184 ( .A(n8328), .ZN(n8327) );
  NAND2_X1 U9185 ( .A1(n8330), .A2(n12355), .ZN(n8328) );
  NOR2_X1 U9186 ( .A1(n8306), .A2(n12811), .ZN(n8303) );
  AND2_X1 U9187 ( .A1(n7301), .A2(n14261), .ZN(n7215) );
  AND2_X1 U9188 ( .A1(n14800), .A2(n14472), .ZN(n7216) );
  AND2_X1 U9189 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7217) );
  AND2_X1 U9190 ( .A1(n14179), .A2(n13445), .ZN(n7218) );
  NAND2_X1 U9191 ( .A1(n9376), .A2(n9375), .ZN(n13364) );
  INV_X1 U9192 ( .A(n13364), .ZN(n14214) );
  OR2_X1 U9193 ( .A1(n13246), .A2(n11647), .ZN(n7219) );
  AND2_X1 U9194 ( .A1(n14214), .A2(n13511), .ZN(n7220) );
  INV_X1 U9195 ( .A(n13329), .ZN(n8012) );
  OR2_X1 U9196 ( .A1(n7797), .A2(n7447), .ZN(n7221) );
  AND2_X1 U9197 ( .A1(n9428), .A2(n9427), .ZN(n13752) );
  INV_X1 U9198 ( .A(n13752), .ZN(n7781) );
  INV_X1 U9199 ( .A(n14872), .ZN(n14748) );
  AND2_X1 U9200 ( .A1(n8854), .A2(n8853), .ZN(n14872) );
  AND4_X1 U9201 ( .A1(n8501), .A2(n9075), .A3(n9080), .A4(n9069), .ZN(n7222)
         );
  AND3_X1 U9202 ( .A1(n8532), .A2(n8527), .A3(n8530), .ZN(n7223) );
  NAND2_X1 U9203 ( .A1(n13210), .A2(n13207), .ZN(n13094) );
  INV_X1 U9204 ( .A(n13094), .ZN(n13930) );
  OR2_X1 U9205 ( .A1(n14428), .A2(n8407), .ZN(n7224) );
  AND2_X1 U9206 ( .A1(n8039), .A2(n8041), .ZN(n7225) );
  NOR2_X1 U9207 ( .A1(n8126), .A2(n14468), .ZN(n7226) );
  AND2_X1 U9208 ( .A1(n13774), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7227) );
  AND2_X1 U9209 ( .A1(n13271), .A2(n9477), .ZN(n7228) );
  AND2_X1 U9210 ( .A1(n8458), .A2(n9611), .ZN(n7229) );
  AND2_X1 U9211 ( .A1(n7881), .A2(n7878), .ZN(n7877) );
  INV_X1 U9212 ( .A(n14105), .ZN(n8426) );
  AND2_X1 U9213 ( .A1(n9051), .A2(n14361), .ZN(n9052) );
  INV_X1 U9214 ( .A(n15662), .ZN(n7546) );
  NAND2_X1 U9215 ( .A1(n9345), .A2(n9344), .ZN(n13329) );
  NAND2_X1 U9216 ( .A1(n9715), .A2(n9714), .ZN(n14002) );
  INV_X1 U9217 ( .A(n14002), .ZN(n13977) );
  NAND2_X1 U9218 ( .A1(n11314), .A2(n7815), .ZN(n7814) );
  INV_X1 U9219 ( .A(n13899), .ZN(n13865) );
  NOR2_X1 U9220 ( .A1(n10017), .A2(SI_29_), .ZN(n7230) );
  AND2_X1 U9221 ( .A1(n7858), .A2(n7861), .ZN(n7231) );
  OR2_X1 U9222 ( .A1(n10804), .A2(n10805), .ZN(n7232) );
  NAND2_X2 U9223 ( .A1(n13320), .A2(n9361), .ZN(n9407) );
  INV_X1 U9224 ( .A(n10755), .ZN(n12027) );
  INV_X2 U9225 ( .A(n12027), .ZN(n12875) );
  AND2_X1 U9226 ( .A1(n8357), .A2(n10596), .ZN(n7765) );
  OAI211_X1 U9227 ( .C1(n10024), .C2(n10701), .A(n8646), .B(n8645), .ZN(n11724) );
  INV_X1 U9228 ( .A(n10761), .ZN(n11704) );
  NAND2_X1 U9229 ( .A1(n8476), .A2(n13339), .ZN(n7233) );
  OR2_X1 U9230 ( .A1(n9788), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n7234) );
  AND2_X1 U9231 ( .A1(n9323), .A2(n9412), .ZN(n9484) );
  NAND2_X1 U9232 ( .A1(n9168), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7235) );
  INV_X1 U9233 ( .A(n8631), .ZN(n14484) );
  AND2_X1 U9234 ( .A1(n11895), .A2(n9035), .ZN(n7236) );
  NAND2_X1 U9235 ( .A1(n14718), .A2(n9047), .ZN(n14722) );
  AND2_X1 U9236 ( .A1(n7827), .A2(n7829), .ZN(n7237) );
  NAND2_X1 U9237 ( .A1(n16027), .A2(n9806), .ZN(n11635) );
  OAI211_X1 U9238 ( .C1(n10522), .C2(n10431), .A(n9404), .B(n9403), .ZN(n16029) );
  INV_X1 U9239 ( .A(n9926), .ZN(n8246) );
  OR2_X1 U9240 ( .A1(n10152), .A2(n10150), .ZN(n7238) );
  AND3_X1 U9241 ( .A1(n10229), .A2(n10230), .A3(n12685), .ZN(n10420) );
  NOR2_X1 U9242 ( .A1(n14662), .A2(n14661), .ZN(n7239) );
  NAND2_X1 U9243 ( .A1(n8168), .A2(n8167), .ZN(n7741) );
  NAND2_X1 U9244 ( .A1(n16070), .A2(n15234), .ZN(n7240) );
  XNOR2_X1 U9245 ( .A(n11508), .B(n14479), .ZN(n11494) );
  INV_X1 U9246 ( .A(n11494), .ZN(n7594) );
  AND2_X1 U9247 ( .A1(n15434), .A2(n8091), .ZN(n7241) );
  AND2_X1 U9248 ( .A1(n8441), .A2(n9675), .ZN(n7242) );
  AND2_X1 U9249 ( .A1(n8190), .A2(n8189), .ZN(n7243) );
  OR2_X1 U9250 ( .A1(n13412), .A2(n13932), .ZN(n9814) );
  XNOR2_X1 U9251 ( .A(n15529), .B(n15376), .ZN(n15522) );
  INV_X1 U9252 ( .A(n15522), .ZN(n8205) );
  NOR2_X1 U9253 ( .A1(n14039), .A2(n14050), .ZN(n7244) );
  INV_X1 U9254 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7727) );
  AND2_X1 U9255 ( .A1(n8383), .A2(n8875), .ZN(n7245) );
  AND2_X1 U9256 ( .A1(n7235), .A2(n15942), .ZN(n7246) );
  AND2_X1 U9257 ( .A1(n7594), .A2(n8703), .ZN(n7247) );
  AND2_X1 U9258 ( .A1(n8344), .A2(n8343), .ZN(n7248) );
  INV_X1 U9259 ( .A(n15092), .ZN(n7828) );
  INV_X1 U9260 ( .A(n10110), .ZN(n8366) );
  OR2_X1 U9261 ( .A1(n11437), .A2(n11438), .ZN(n7249) );
  INV_X1 U9262 ( .A(n16190), .ZN(n9243) );
  AND2_X1 U9263 ( .A1(n13205), .A2(n13204), .ZN(n13940) );
  INV_X1 U9264 ( .A(n13940), .ZN(n13938) );
  OAI211_X1 U9265 ( .C1(n10024), .C2(n10692), .A(n8623), .B(n7772), .ZN(n10980) );
  XNOR2_X1 U9266 ( .A(n9413), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10628) );
  OR2_X1 U9267 ( .A1(n8379), .A2(SI_9_), .ZN(n7250) );
  NOR2_X1 U9268 ( .A1(n12742), .A2(n10708), .ZN(n7251) );
  OR2_X1 U9269 ( .A1(n10178), .A2(n10227), .ZN(n7252) );
  INV_X1 U9270 ( .A(n12795), .ZN(n7526) );
  NAND2_X1 U9271 ( .A1(n8356), .A2(n13449), .ZN(n13389) );
  AND2_X1 U9272 ( .A1(n8103), .A2(n8104), .ZN(n7253) );
  NAND2_X1 U9273 ( .A1(n12947), .A2(n12946), .ZN(n15636) );
  INV_X1 U9274 ( .A(n15636), .ZN(n15427) );
  AND2_X1 U9275 ( .A1(n7836), .A2(n7833), .ZN(n7254) );
  INV_X1 U9276 ( .A(n10101), .ZN(n14757) );
  AND4_X1 U9277 ( .A1(n8584), .A2(n8583), .A3(n8582), .A4(n9071), .ZN(n7255)
         );
  INV_X1 U9278 ( .A(n12945), .ZN(n8311) );
  NAND2_X1 U9279 ( .A1(n16186), .A2(n12335), .ZN(n7256) );
  NAND2_X1 U9280 ( .A1(n15113), .A2(n15025), .ZN(n15168) );
  INV_X1 U9281 ( .A(n9900), .ZN(n7910) );
  NAND2_X1 U9282 ( .A1(n14400), .A2(n14399), .ZN(n14398) );
  AND2_X1 U9283 ( .A1(n7932), .A2(n7930), .ZN(n7257) );
  AND2_X1 U9284 ( .A1(n7255), .A2(n7222), .ZN(n7258) );
  AND2_X1 U9285 ( .A1(n15733), .A2(n12601), .ZN(n7259) );
  OR2_X1 U9286 ( .A1(n13092), .A2(n16138), .ZN(n7260) );
  NAND2_X1 U9287 ( .A1(n9171), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n9170) );
  INV_X1 U9288 ( .A(n9170), .ZN(n7973) );
  AND2_X1 U9289 ( .A1(n8049), .A2(n9814), .ZN(n7261) );
  NAND2_X1 U9290 ( .A1(n8643), .A2(n8394), .ZN(n8657) );
  AND2_X1 U9291 ( .A1(n8332), .A2(n13486), .ZN(n7262) );
  AND2_X1 U9292 ( .A1(n12510), .A2(n12511), .ZN(n7263) );
  INV_X1 U9293 ( .A(n7884), .ZN(n7883) );
  AND2_X1 U9294 ( .A1(n14410), .A2(n7870), .ZN(n7264) );
  INV_X1 U9295 ( .A(n7856), .ZN(n7855) );
  NOR2_X1 U9296 ( .A1(n7860), .A2(n7857), .ZN(n7856) );
  INV_X1 U9297 ( .A(n14569), .ZN(n9248) );
  NAND2_X1 U9298 ( .A1(n8590), .A2(n8589), .ZN(n14569) );
  INV_X1 U9299 ( .A(n13200), .ZN(n8035) );
  NAND2_X1 U9300 ( .A1(n13769), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7265) );
  NAND2_X1 U9301 ( .A1(n7670), .A2(n16035), .ZN(n10638) );
  OR2_X1 U9302 ( .A1(n7449), .A2(n13820), .ZN(n7266) );
  OR2_X1 U9303 ( .A1(n12204), .A2(n7544), .ZN(n7267) );
  INV_X1 U9304 ( .A(n8112), .ZN(n8111) );
  AOI21_X1 U9305 ( .B1(n15498), .B2(n8113), .A(n8117), .ZN(n8112) );
  AND2_X1 U9306 ( .A1(n12295), .A2(n11679), .ZN(n7268) );
  AND2_X1 U9307 ( .A1(n15778), .A2(n10691), .ZN(n15672) );
  INV_X1 U9308 ( .A(n15672), .ZN(n15529) );
  AND2_X1 U9309 ( .A1(n12138), .A2(n8759), .ZN(n7269) );
  AND2_X1 U9310 ( .A1(n14840), .A2(n14362), .ZN(n7270) );
  NOR2_X1 U9311 ( .A1(n8223), .A2(n9979), .ZN(n8221) );
  INV_X1 U9312 ( .A(n12860), .ZN(n7519) );
  INV_X1 U9313 ( .A(n7663), .ZN(n7662) );
  NAND2_X1 U9314 ( .A1(n8338), .A2(n7666), .ZN(n7663) );
  INV_X1 U9315 ( .A(n8409), .ZN(n8408) );
  NAND2_X1 U9316 ( .A1(n14285), .A2(n14284), .ZN(n8409) );
  AND2_X1 U9317 ( .A1(n15022), .A2(n15020), .ZN(n7271) );
  INV_X1 U9318 ( .A(n7487), .ZN(n15443) );
  NOR2_X1 U9319 ( .A1(n15504), .A2(n8018), .ZN(n7487) );
  AND2_X1 U9320 ( .A1(n9921), .A2(n9920), .ZN(n7272) );
  INV_X1 U9321 ( .A(n8450), .ZN(n8449) );
  OAI21_X1 U9322 ( .B1(n9754), .B2(n8451), .A(n8454), .ZN(n8450) );
  OR2_X1 U9323 ( .A1(n10317), .A2(n16118), .ZN(n7273) );
  OR2_X1 U9324 ( .A1(n15296), .A2(n10306), .ZN(n7274) );
  OR2_X1 U9325 ( .A1(n9981), .A2(n9980), .ZN(n7275) );
  INV_X1 U9326 ( .A(n8807), .ZN(n8143) );
  AND2_X1 U9327 ( .A1(n15427), .A2(n15438), .ZN(n7276) );
  NAND2_X1 U9328 ( .A1(n8326), .A2(n8330), .ZN(n8325) );
  OR2_X1 U9329 ( .A1(n13979), .A2(n8035), .ZN(n7277) );
  INV_X1 U9330 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n9340) );
  AND2_X1 U9331 ( .A1(n7608), .A2(n8362), .ZN(n7278) );
  AND2_X1 U9332 ( .A1(n14994), .A2(n14993), .ZN(n7279) );
  AND2_X1 U9333 ( .A1(n7629), .A2(n13930), .ZN(n7280) );
  OR2_X1 U9334 ( .A1(n12171), .A2(n7544), .ZN(n7281) );
  INV_X1 U9335 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9330) );
  NOR2_X1 U9336 ( .A1(n12780), .A2(n11916), .ZN(n7282) );
  NOR2_X1 U9337 ( .A1(n15002), .A2(n15001), .ZN(n7283) );
  NOR2_X1 U9338 ( .A1(n14601), .A2(n14614), .ZN(n7284) );
  NOR2_X1 U9339 ( .A1(n15688), .A2(n15373), .ZN(n7285) );
  AND2_X1 U9340 ( .A1(n8319), .A2(n8321), .ZN(n7286) );
  AND2_X1 U9341 ( .A1(n7371), .A2(n8225), .ZN(n7287) );
  INV_X1 U9342 ( .A(n8675), .ZN(n7615) );
  NAND2_X1 U9343 ( .A1(n9484), .A2(n7420), .ZN(n9632) );
  INV_X1 U9344 ( .A(n9632), .ZN(n7678) );
  NAND2_X1 U9345 ( .A1(n13283), .A2(n7277), .ZN(n7288) );
  AND2_X1 U9346 ( .A1(n8333), .A2(n13426), .ZN(n7289) );
  OR2_X1 U9347 ( .A1(n7216), .A2(n8807), .ZN(n7290) );
  INV_X1 U9348 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10146) );
  INV_X1 U9349 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U9350 ( .A1(n8160), .A2(n10529), .ZN(n10530) );
  INV_X1 U9351 ( .A(n9052), .ZN(n7602) );
  AND2_X1 U9352 ( .A1(n13749), .A2(n7780), .ZN(n7291) );
  AND2_X1 U9353 ( .A1(n7499), .A2(n7503), .ZN(n7292) );
  AND2_X1 U9354 ( .A1(n12944), .A2(n8311), .ZN(n7293) );
  OR2_X1 U9355 ( .A1(n13299), .A2(n13298), .ZN(n7294) );
  INV_X1 U9356 ( .A(n8428), .ZN(n8427) );
  OR2_X1 U9357 ( .A1(n9578), .A2(n8429), .ZN(n8428) );
  AND2_X1 U9358 ( .A1(n8295), .A2(n13025), .ZN(n7295) );
  AND2_X1 U9359 ( .A1(n8375), .A2(n7470), .ZN(n7296) );
  AND2_X1 U9360 ( .A1(n8012), .A2(n13943), .ZN(n7297) );
  XNOR2_X1 U9361 ( .A(n13364), .B(n13511), .ZN(n13952) );
  INV_X1 U9362 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10220) );
  INV_X1 U9363 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8486) );
  INV_X1 U9364 ( .A(n8088), .ZN(n8087) );
  NAND2_X1 U9365 ( .A1(n15420), .A2(n8092), .ZN(n8088) );
  INV_X1 U9366 ( .A(n8226), .ZN(n8225) );
  NOR2_X1 U9367 ( .A1(n8227), .A2(n9991), .ZN(n8226) );
  AND2_X1 U9368 ( .A1(n15061), .A2(n15060), .ZN(n7298) );
  AND2_X1 U9369 ( .A1(n8548), .A2(n10222), .ZN(n7299) );
  INV_X1 U9370 ( .A(n13369), .ZN(n14210) );
  NAND2_X1 U9371 ( .A1(n9746), .A2(n9745), .ZN(n13369) );
  NAND2_X1 U9372 ( .A1(n12242), .A2(n12240), .ZN(n7300) );
  AND2_X1 U9373 ( .A1(n14263), .A2(n14270), .ZN(n7301) );
  AND2_X1 U9374 ( .A1(n9337), .A2(n9340), .ZN(n7302) );
  NAND2_X1 U9375 ( .A1(n10212), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n7303) );
  OR2_X1 U9376 ( .A1(n8311), .A2(n12944), .ZN(n7304) );
  INV_X1 U9377 ( .A(n7391), .ZN(n9638) );
  NOR2_X1 U9378 ( .A1(n9621), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7391) );
  INV_X1 U9379 ( .A(n7393), .ZN(n9693) );
  NOR2_X1 U9380 ( .A1(n9682), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7393) );
  AND2_X1 U9381 ( .A1(n14654), .A2(n14632), .ZN(n7305) );
  INV_X1 U9382 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U9383 ( .A1(n7665), .A2(n12122), .ZN(n7306) );
  INV_X1 U9384 ( .A(n8197), .ZN(n8196) );
  NAND2_X1 U9385 ( .A1(n15547), .A2(n15399), .ZN(n8197) );
  INV_X1 U9386 ( .A(n12798), .ZN(n8297) );
  OR2_X1 U9387 ( .A1(n10180), .A2(n9705), .ZN(n7307) );
  OR2_X1 U9388 ( .A1(n9970), .A2(n9972), .ZN(n7308) );
  OR2_X1 U9389 ( .A1(n9990), .A2(n9992), .ZN(n7309) );
  OR2_X1 U9390 ( .A1(n9948), .A2(n9946), .ZN(n7310) );
  OR2_X1 U9391 ( .A1(n9998), .A2(n9999), .ZN(n7311) );
  AND2_X1 U9392 ( .A1(n14155), .A2(n14015), .ZN(n7312) );
  OR2_X1 U9393 ( .A1(n8228), .A2(n9971), .ZN(n7313) );
  INV_X1 U9394 ( .A(n15459), .ZN(n15648) );
  NAND2_X1 U9395 ( .A1(n12930), .A2(n12929), .ZN(n15459) );
  INV_X1 U9396 ( .A(n15654), .ZN(n15470) );
  NAND2_X1 U9397 ( .A1(n12919), .A2(n12918), .ZN(n15654) );
  AND2_X1 U9398 ( .A1(n9924), .A2(n11508), .ZN(n7314) );
  AND2_X1 U9399 ( .A1(n15520), .A2(n8203), .ZN(n7315) );
  OR2_X1 U9400 ( .A1(n8300), .A2(n8301), .ZN(n7316) );
  NOR2_X1 U9401 ( .A1(n13073), .A2(n13074), .ZN(n7317) );
  INV_X1 U9402 ( .A(n8530), .ZN(n8361) );
  AND2_X1 U9403 ( .A1(n8369), .A2(n8367), .ZN(n7318) );
  AND2_X1 U9404 ( .A1(n8094), .A2(n15401), .ZN(n7319) );
  INV_X1 U9405 ( .A(n8128), .ZN(n8127) );
  NOR2_X1 U9406 ( .A1(n14861), .A2(n14469), .ZN(n8128) );
  INV_X1 U9407 ( .A(n8745), .ZN(n8379) );
  AND2_X1 U9408 ( .A1(n7199), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n7320) );
  OR2_X1 U9409 ( .A1(n9335), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n7321) );
  INV_X1 U9410 ( .A(n12933), .ZN(n7513) );
  AND2_X1 U9411 ( .A1(n8110), .A2(n8112), .ZN(n7322) );
  OR2_X1 U9412 ( .A1(n12828), .A2(n12826), .ZN(n7323) );
  NAND2_X1 U9413 ( .A1(n7237), .A2(n7822), .ZN(n7324) );
  AND2_X1 U9414 ( .A1(n13769), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7957) );
  INV_X1 U9415 ( .A(n7957), .ZN(n7956) );
  AND2_X1 U9416 ( .A1(n7864), .A2(n7866), .ZN(n7325) );
  AND2_X1 U9417 ( .A1(n7302), .A2(n9359), .ZN(n7326) );
  NAND2_X1 U9418 ( .A1(n8314), .A2(n12873), .ZN(n7327) );
  INV_X1 U9419 ( .A(n8517), .ZN(n8520) );
  NAND3_X1 U9420 ( .A1(n7742), .A2(SI_1_), .A3(n7561), .ZN(n8517) );
  AND2_X1 U9421 ( .A1(n8089), .A2(n8092), .ZN(n7328) );
  NOR2_X1 U9422 ( .A1(n11440), .A2(n11439), .ZN(n7329) );
  NAND2_X1 U9423 ( .A1(n9935), .A2(n9936), .ZN(n7330) );
  NAND2_X1 U9424 ( .A1(n12860), .A2(n7520), .ZN(n7331) );
  NAND2_X1 U9425 ( .A1(n8549), .A2(SI_13_), .ZN(n8550) );
  INV_X1 U9426 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7941) );
  INV_X1 U9427 ( .A(n7950), .ZN(n7949) );
  NAND2_X1 U9428 ( .A1(n7955), .A2(n7953), .ZN(n7950) );
  AND2_X1 U9429 ( .A1(n12795), .A2(n7527), .ZN(n7332) );
  INV_X1 U9430 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10218) );
  INV_X1 U9431 ( .A(n13374), .ZN(n7739) );
  INV_X1 U9432 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10207) );
  INV_X1 U9433 ( .A(n15406), .ZN(n7468) );
  INV_X1 U9434 ( .A(n13268), .ZN(n8041) );
  NAND4_X1 U9435 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n9882)
         );
  INV_X1 U9436 ( .A(n11965), .ZN(n8171) );
  NAND2_X1 U9437 ( .A1(n15395), .A2(n7549), .ZN(n15605) );
  INV_X1 U9438 ( .A(n13990), .ZN(n8028) );
  NAND2_X1 U9439 ( .A1(n14104), .A2(n14105), .ZN(n14085) );
  INV_X1 U9440 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8078) );
  INV_X2 U9441 ( .A(n11704), .ZN(n12982) );
  AND2_X1 U9442 ( .A1(n9366), .A2(n9365), .ZN(n13943) );
  INV_X1 U9443 ( .A(n13943), .ZN(n8011) );
  AOI21_X1 U9444 ( .B1(n13923), .B2(n9778), .A(n9768), .ZN(n13932) );
  INV_X1 U9445 ( .A(n8809), .ZN(n7878) );
  INV_X1 U9446 ( .A(n13425), .ZN(n8336) );
  NAND2_X1 U9447 ( .A1(n8098), .A2(n8103), .ZN(n12659) );
  AND2_X1 U9448 ( .A1(n9728), .A2(n9727), .ZN(n13966) );
  INV_X1 U9449 ( .A(n13136), .ZN(n8040) );
  NAND2_X1 U9450 ( .A1(n7620), .A2(n7618), .ZN(n14067) );
  NAND2_X1 U9451 ( .A1(n8444), .A2(n9525), .ZN(n12429) );
  NAND2_X1 U9452 ( .A1(n12173), .A2(n12073), .ZN(n12183) );
  AND2_X1 U9453 ( .A1(n7867), .A2(n14261), .ZN(n7333) );
  INV_X1 U9454 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U9455 ( .A1(n9551), .A2(n9550), .ZN(n12306) );
  NAND2_X1 U9456 ( .A1(n8616), .A2(n8615), .ZN(n14580) );
  OR2_X1 U9457 ( .A1(n14155), .A2(n14015), .ZN(n7334) );
  NAND2_X1 U9458 ( .A1(n8457), .A2(n8456), .ZN(n14055) );
  OR2_X1 U9459 ( .A1(n12663), .A2(n15719), .ZN(n7335) );
  INV_X1 U9460 ( .A(n9807), .ZN(n13262) );
  NAND2_X1 U9461 ( .A1(n13107), .A2(n13108), .ZN(n9807) );
  OR2_X1 U9462 ( .A1(n14242), .A2(n14106), .ZN(n13164) );
  INV_X1 U9463 ( .A(n13164), .ZN(n8054) );
  NAND2_X1 U9464 ( .A1(n8798), .A2(n8483), .ZN(n8824) );
  INV_X1 U9465 ( .A(n13511), .ZN(n13965) );
  NAND2_X1 U9466 ( .A1(n9372), .A2(n9371), .ZN(n13511) );
  AND4_X1 U9467 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(n14453)
         );
  OR2_X1 U9468 ( .A1(n15316), .A2(n10578), .ZN(n7336) );
  NAND2_X1 U9469 ( .A1(n7333), .A2(n14263), .ZN(n14324) );
  NAND2_X1 U9470 ( .A1(n14324), .A2(n8405), .ZN(n7337) );
  INV_X1 U9471 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8495) );
  INV_X1 U9472 ( .A(n13966), .ZN(n13988) );
  NAND2_X1 U9473 ( .A1(n8798), .A2(n8413), .ZN(n7338) );
  AND2_X1 U9474 ( .A1(n8560), .A2(n10649), .ZN(n7339) );
  INV_X1 U9475 ( .A(n12552), .ZN(n8429) );
  INV_X1 U9476 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10679) );
  AND2_X1 U9477 ( .A1(n13377), .A2(n7778), .ZN(n7340) );
  NOR2_X1 U9478 ( .A1(n9099), .A2(n8390), .ZN(n7341) );
  AND2_X1 U9479 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n10685), .ZN(n7342) );
  AND2_X1 U9480 ( .A1(n15564), .A2(n15372), .ZN(n7343) );
  OR2_X1 U9481 ( .A1(n8554), .A2(SI_15_), .ZN(n7344) );
  AND2_X1 U9482 ( .A1(n9880), .A2(n7685), .ZN(n7345) );
  AND2_X1 U9483 ( .A1(n9863), .A2(n7688), .ZN(n7346) );
  AND2_X1 U9484 ( .A1(n7645), .A2(n7646), .ZN(n7347) );
  INV_X1 U9485 ( .A(SI_9_), .ZN(n8381) );
  AND3_X2 U9486 ( .A1(n11058), .A2(n9876), .A3(n9875), .ZN(n16228) );
  INV_X1 U9487 ( .A(n16228), .ZN(n7687) );
  INV_X2 U9488 ( .A(n15611), .ZN(n16022) );
  NAND2_X1 U9489 ( .A1(n10705), .A2(n10746), .ZN(n13012) );
  NAND2_X1 U9490 ( .A1(n12020), .A2(n7839), .ZN(n7838) );
  INV_X1 U9491 ( .A(n13801), .ZN(n7449) );
  INV_X1 U9492 ( .A(n15502), .ZN(n8118) );
  INV_X1 U9493 ( .A(n9342), .ZN(n10438) );
  NAND2_X1 U9494 ( .A1(n7656), .A2(n7655), .ZN(n12356) );
  NAND2_X1 U9495 ( .A1(n13313), .A2(n13102), .ZN(n13217) );
  INV_X1 U9496 ( .A(n13217), .ZN(n13229) );
  NAND2_X1 U9497 ( .A1(n12598), .A2(n12597), .ZN(n15729) );
  INV_X1 U9498 ( .A(n15729), .ZN(n8025) );
  INV_X1 U9499 ( .A(SI_18_), .ZN(n13630) );
  AND2_X1 U9500 ( .A1(n9848), .A2(n9847), .ZN(n14250) );
  INV_X1 U9501 ( .A(n16208), .ZN(n16206) );
  AND2_X2 U9502 ( .A1(n9125), .A2(n9098), .ZN(n16208) );
  NAND2_X1 U9503 ( .A1(n7664), .A2(n7666), .ZN(n12123) );
  XOR2_X1 U9504 ( .A(n8579), .B(SI_26_), .Z(n7348) );
  OR2_X1 U9505 ( .A1(n11914), .A2(n11913), .ZN(n7349) );
  OR2_X1 U9506 ( .A1(n12570), .A2(n12569), .ZN(n7350) );
  AND2_X1 U9507 ( .A1(n12371), .A2(n8283), .ZN(n7351) );
  NOR2_X1 U9508 ( .A1(n11255), .A2(n11254), .ZN(n7352) );
  INV_X1 U9509 ( .A(n8016), .ZN(n12349) );
  NOR2_X1 U9510 ( .A1(n12165), .A2(n12797), .ZN(n8016) );
  AND2_X1 U9511 ( .A1(n7813), .A2(n7812), .ZN(n7353) );
  AND2_X1 U9512 ( .A1(n8564), .A2(SI_21_), .ZN(n7354) );
  NAND2_X1 U9513 ( .A1(n8265), .A2(n8264), .ZN(n7355) );
  AND2_X1 U9514 ( .A1(n8135), .A2(n9035), .ZN(n7356) );
  INV_X1 U9515 ( .A(n15205), .ZN(n15210) );
  INV_X1 U9516 ( .A(n13520), .ZN(n7795) );
  XNOR2_X1 U9517 ( .A(n8587), .B(n8586), .ZN(n9064) );
  INV_X1 U9518 ( .A(n12780), .ZN(n7485) );
  AND2_X1 U9519 ( .A1(n10498), .A2(n10614), .ZN(n7357) );
  NAND2_X1 U9520 ( .A1(n12189), .A2(n12188), .ZN(n12801) );
  INV_X1 U9521 ( .A(n12801), .ZN(n8015) );
  AND2_X1 U9522 ( .A1(n10458), .A2(n10466), .ZN(n13495) );
  NAND2_X2 U9523 ( .A1(n8629), .A2(n10689), .ZN(n10024) );
  AND2_X1 U9524 ( .A1(n7933), .A2(n13882), .ZN(n7358) );
  INV_X1 U9525 ( .A(n13741), .ZN(n7406) );
  AND2_X1 U9526 ( .A1(n14876), .A2(n9243), .ZN(n16138) );
  INV_X1 U9527 ( .A(n12622), .ZN(n8324) );
  NAND2_X1 U9528 ( .A1(n7248), .A2(n7793), .ZN(n8342) );
  INV_X1 U9529 ( .A(n13862), .ZN(n7933) );
  INV_X1 U9530 ( .A(n7861), .ZN(n7860) );
  NAND2_X1 U9531 ( .A1(n11674), .A2(n11675), .ZN(n7861) );
  INV_X1 U9532 ( .A(n13868), .ZN(n8166) );
  INV_X1 U9533 ( .A(n10368), .ZN(n8084) );
  INV_X1 U9534 ( .A(n13779), .ZN(n7958) );
  INV_X1 U9535 ( .A(n10807), .ZN(n7442) );
  AND2_X1 U9536 ( .A1(n7967), .A2(n15941), .ZN(n7359) );
  XOR2_X1 U9537 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n7360) );
  INV_X1 U9538 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8419) );
  INV_X1 U9539 ( .A(n7731), .ZN(n7710) );
  INV_X1 U9540 ( .A(n10803), .ZN(n7953) );
  NAND2_X1 U9541 ( .A1(n7952), .A2(n10803), .ZN(n7951) );
  XNOR2_X1 U9542 ( .A(n10802), .B(n10803), .ZN(n10672) );
  NAND3_X1 U9543 ( .A1(n8556), .A2(n8555), .A3(n8373), .ZN(n8851) );
  NOR2_X2 U9544 ( .A1(n15515), .A2(n7362), .ZN(n15499) );
  OAI211_X1 U9546 ( .C1(n7367), .C2(n8247), .A(n7365), .B(n7364), .ZN(n9929)
         );
  OR2_X1 U9547 ( .A1(n8245), .A2(n7366), .ZN(n7365) );
  NOR2_X1 U9548 ( .A1(n9925), .A2(n9926), .ZN(n7367) );
  OAI21_X1 U9549 ( .B1(n7371), .B2(n7370), .A(n7368), .ZN(n9996) );
  NAND3_X1 U9550 ( .A1(n9989), .A2(n8465), .A3(n7309), .ZN(n7371) );
  AOI21_X1 U9551 ( .B1(n7373), .B2(n9909), .A(n7372), .ZN(n9906) );
  NAND3_X1 U9552 ( .A1(n7376), .A2(n7375), .A3(n8239), .ZN(n7374) );
  NOR2_X1 U9553 ( .A1(n7377), .A2(n9917), .ZN(n9918) );
  NAND2_X1 U9554 ( .A1(n9913), .A2(n9912), .ZN(n7377) );
  AND2_X4 U9555 ( .A1(n16190), .A2(n8503), .ZN(n10055) );
  NAND2_X1 U9556 ( .A1(n7379), .A2(n8214), .ZN(n7378) );
  NAND2_X1 U9557 ( .A1(n7381), .A2(n7380), .ZN(n7379) );
  NAND2_X1 U9558 ( .A1(n9978), .A2(n9977), .ZN(n7380) );
  NAND2_X1 U9559 ( .A1(n9974), .A2(n9973), .ZN(n7381) );
  NAND2_X1 U9560 ( .A1(n7382), .A2(n10091), .ZN(n10124) );
  NAND2_X1 U9561 ( .A1(n7383), .A2(n10076), .ZN(n7382) );
  NAND3_X1 U9562 ( .A1(n8211), .A2(n10015), .A3(n10011), .ZN(n7383) );
  AND2_X2 U9563 ( .A1(n7615), .A2(n7385), .ZN(n8798) );
  NAND4_X1 U9564 ( .A1(n8478), .A2(n8481), .A3(n8479), .A4(n8480), .ZN(n8482)
         );
  NAND3_X1 U9565 ( .A1(n13696), .A2(n11104), .A3(n9346), .ZN(n9447) );
  NAND3_X1 U9566 ( .A1(n7398), .A2(n7397), .A3(n7396), .ZN(n7395) );
  NAND2_X1 U9567 ( .A1(n8444), .A2(n8442), .ZN(n7403) );
  AND2_X2 U9568 ( .A1(n11479), .A2(n9446), .ZN(n11468) );
  NOR2_X2 U9569 ( .A1(n13950), .A2(n13952), .ZN(n13951) );
  NAND2_X1 U9570 ( .A1(n14048), .A2(n14047), .ZN(n14046) );
  NAND2_X1 U9571 ( .A1(n14084), .A2(n7229), .ZN(n8457) );
  NAND3_X1 U9572 ( .A1(n8461), .A2(n9406), .A3(n9807), .ZN(n11633) );
  NAND2_X1 U9573 ( .A1(n10551), .A2(n10552), .ZN(n10492) );
  NAND2_X1 U9574 ( .A1(n10486), .A2(n10526), .ZN(n7410) );
  NAND2_X1 U9575 ( .A1(n12472), .A2(n12471), .ZN(n13800) );
  INV_X1 U9576 ( .A(n12312), .ZN(n7412) );
  NAND3_X1 U9577 ( .A1(n7928), .A2(n7927), .A3(n8174), .ZN(n7414) );
  NAND3_X1 U9578 ( .A1(n7740), .A2(n7417), .A3(n7415), .ZN(P3_U3201) );
  NAND2_X1 U9579 ( .A1(n13898), .A2(n13897), .ZN(n7417) );
  NAND4_X1 U9580 ( .A1(n9484), .A2(n7418), .A3(n7421), .A4(n7420), .ZN(n9339)
         );
  NOR2_X2 U9581 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n10190) );
  XNOR2_X1 U9582 ( .A(n9181), .B(n7429), .ZN(n15943) );
  NAND2_X1 U9583 ( .A1(n9183), .A2(n7431), .ZN(n7966) );
  INV_X1 U9584 ( .A(n15945), .ZN(n7431) );
  INV_X1 U9585 ( .A(n10622), .ZN(n13747) );
  NAND2_X1 U9586 ( .A1(n10530), .A2(n10622), .ZN(n7435) );
  INV_X1 U9587 ( .A(n7439), .ZN(n15960) );
  AND2_X1 U9588 ( .A1(n7439), .A2(n7438), .ZN(n15959) );
  INV_X1 U9589 ( .A(n7437), .ZN(n7436) );
  OR2_X2 U9590 ( .A1(n7440), .A2(n15955), .ZN(n7439) );
  NOR2_X1 U9591 ( .A1(n15957), .A2(n15956), .ZN(n15955) );
  AOI21_X1 U9592 ( .B1(n15957), .B2(n15956), .A(n7441), .ZN(n7440) );
  INV_X1 U9593 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7441) );
  NOR2_X1 U9594 ( .A1(n11020), .A2(n11007), .ZN(n11576) );
  MUX2_X1 U9595 ( .A(n7446), .B(n7443), .S(P3_IR_REG_8__SCAN_IN), .Z(n9485) );
  MUX2_X1 U9596 ( .A(n7446), .B(n7444), .S(P3_IR_REG_12__SCAN_IN), .Z(n9547)
         );
  MUX2_X1 U9597 ( .A(n7446), .B(n7445), .S(P3_IR_REG_13__SCAN_IN), .Z(n9565)
         );
  NAND2_X1 U9598 ( .A1(n8162), .A2(n8161), .ZN(n13776) );
  OR2_X1 U9599 ( .A1(n8906), .A2(n8562), .ZN(n7455) );
  NAND2_X1 U9600 ( .A1(n7875), .A2(n7876), .ZN(n8823) );
  NAND2_X1 U9601 ( .A1(n7872), .A2(SI_16_), .ZN(n8556) );
  NAND3_X1 U9602 ( .A1(n7250), .A2(n8538), .A3(n7471), .ZN(n7470) );
  NAND2_X1 U9603 ( .A1(n15422), .A2(n15421), .ZN(n15635) );
  NAND2_X1 U9604 ( .A1(n8509), .A2(n7478), .ZN(n8510) );
  AND2_X2 U9605 ( .A1(n7844), .A2(n7843), .ZN(n8515) );
  NOR2_X2 U9606 ( .A1(n11823), .A2(n16152), .ZN(n12166) );
  NAND2_X1 U9607 ( .A1(n15597), .A2(n15591), .ZN(n15592) );
  NOR2_X2 U9608 ( .A1(n15423), .A2(n15634), .ZN(n15383) );
  NAND2_X2 U9609 ( .A1(n10691), .A2(n10689), .ZN(n13000) );
  NAND2_X1 U9610 ( .A1(n8024), .A2(n7491), .ZN(n10725) );
  NAND3_X1 U9611 ( .A1(n7496), .A2(n7494), .A3(n7492), .ZN(n8289) );
  NAND2_X1 U9612 ( .A1(n7493), .A2(n12777), .ZN(n7492) );
  INV_X1 U9613 ( .A(n7498), .ZN(n7493) );
  INV_X1 U9614 ( .A(n12778), .ZN(n7495) );
  NAND2_X1 U9615 ( .A1(n7497), .A2(n12775), .ZN(n7496) );
  NAND2_X1 U9616 ( .A1(n7498), .A2(n12776), .ZN(n7497) );
  NAND2_X1 U9617 ( .A1(n12885), .A2(n7503), .ZN(n7502) );
  NAND2_X1 U9618 ( .A1(n12782), .A2(n7508), .ZN(n7507) );
  NAND3_X1 U9619 ( .A1(n7736), .A2(n7733), .A3(n7331), .ZN(n7516) );
  NAND2_X1 U9620 ( .A1(n12839), .A2(n12842), .ZN(n7521) );
  NOR2_X1 U9621 ( .A1(n12842), .A2(n12839), .ZN(n7522) );
  NAND2_X1 U9622 ( .A1(n7524), .A2(n7295), .ZN(n12804) );
  OAI211_X1 U9623 ( .C1(n12796), .C2(n7332), .A(n7525), .B(n8294), .ZN(n7524)
         );
  NAND2_X1 U9624 ( .A1(n7528), .A2(n7316), .ZN(n8298) );
  NAND3_X1 U9625 ( .A1(n7533), .A2(n7531), .A3(n8308), .ZN(n7698) );
  NAND2_X1 U9626 ( .A1(n7532), .A2(n7713), .ZN(n7531) );
  INV_X1 U9627 ( .A(n7535), .ZN(n7532) );
  NAND2_X1 U9628 ( .A1(n7534), .A2(n12910), .ZN(n7533) );
  NAND2_X1 U9629 ( .A1(n7535), .A2(n12911), .ZN(n7534) );
  INV_X1 U9630 ( .A(n13012), .ZN(n10718) );
  NAND2_X1 U9631 ( .A1(n10779), .A2(n10695), .ZN(n10706) );
  NAND2_X1 U9632 ( .A1(n10717), .A2(n10694), .ZN(n10779) );
  INV_X1 U9633 ( .A(n12345), .ZN(n12208) );
  NAND2_X1 U9634 ( .A1(n12525), .A2(n7547), .ZN(n12615) );
  NAND2_X1 U9635 ( .A1(n12615), .A2(n8198), .ZN(n12650) );
  NAND2_X1 U9636 ( .A1(n7551), .A2(n7209), .ZN(n7550) );
  NAND3_X1 U9637 ( .A1(n8057), .A2(n8058), .A3(n8469), .ZN(n10152) );
  NAND2_X1 U9638 ( .A1(n8149), .A2(n8148), .ZN(n12325) );
  INV_X1 U9639 ( .A(n12325), .ZN(n7557) );
  NAND2_X1 U9640 ( .A1(n7553), .A2(n8140), .ZN(n14780) );
  NAND2_X1 U9641 ( .A1(n12325), .A2(n7558), .ZN(n7553) );
  NAND2_X1 U9642 ( .A1(n8140), .A2(n7555), .ZN(n7554) );
  NAND2_X1 U9643 ( .A1(n7557), .A2(n8140), .ZN(n7556) );
  INV_X1 U9644 ( .A(n8515), .ZN(n7560) );
  NAND2_X1 U9645 ( .A1(n8673), .A2(n8527), .ZN(n8691) );
  NAND2_X1 U9646 ( .A1(n7759), .A2(n8926), .ZN(n14656) );
  NAND2_X1 U9647 ( .A1(n7567), .A2(n7565), .ZN(n8959) );
  INV_X1 U9648 ( .A(n7566), .ZN(n7565) );
  OAI21_X1 U9649 ( .B1(n7571), .B2(n14655), .A(n14630), .ZN(n7566) );
  NAND2_X1 U9650 ( .A1(n7570), .A2(n8942), .ZN(n14628) );
  NAND2_X1 U9651 ( .A1(n14656), .A2(n14655), .ZN(n7570) );
  NAND2_X1 U9652 ( .A1(n14610), .A2(n7575), .ZN(n7574) );
  NAND2_X1 U9653 ( .A1(n7584), .A2(n8703), .ZN(n11493) );
  NOR2_X1 U9654 ( .A1(n9235), .A2(n7714), .ZN(n9024) );
  OAI21_X2 U9655 ( .B1(n7595), .B2(n7594), .A(n7592), .ZN(n11660) );
  AOI21_X1 U9656 ( .B1(n7593), .B2(n11494), .A(n7314), .ZN(n7592) );
  AOI21_X2 U9657 ( .B1(n7599), .B2(n7596), .A(n7305), .ZN(n14631) );
  OAI211_X1 U9658 ( .C1(n11406), .C2(n7605), .A(n9030), .B(n7603), .ZN(n11596)
         );
  INV_X1 U9659 ( .A(n10994), .ZN(n7605) );
  INV_X1 U9660 ( .A(n9028), .ZN(n7604) );
  NAND2_X1 U9661 ( .A1(n7611), .A2(n7610), .ZN(n14760) );
  NAND3_X1 U9662 ( .A1(n7613), .A2(n7258), .A3(n7612), .ZN(n8588) );
  NOR2_X1 U9663 ( .A1(n8482), .A2(n7614), .ZN(n7613) );
  NAND2_X1 U9664 ( .A1(n14102), .A2(n7622), .ZN(n7620) );
  AND2_X2 U9665 ( .A1(n7625), .A2(n7631), .ZN(n13928) );
  INV_X1 U9666 ( .A(n13991), .ZN(n8029) );
  NAND2_X1 U9667 ( .A1(n14014), .A2(n7636), .ZN(n14004) );
  NAND2_X1 U9668 ( .A1(n9825), .A2(n7320), .ZN(n7640) );
  OR2_X1 U9669 ( .A1(n9825), .A2(n7642), .ZN(n7641) );
  NAND3_X1 U9670 ( .A1(n7641), .A2(n7640), .A3(n7638), .ZN(n9361) );
  INV_X2 U9671 ( .A(n9361), .ZN(n12397) );
  INV_X2 U9672 ( .A(n13738), .ZN(n16035) );
  OAI211_X2 U9673 ( .C1(n9605), .C2(n10603), .A(n8417), .B(n7219), .ZN(n13738)
         );
  NAND2_X1 U9674 ( .A1(n13373), .A2(n13374), .ZN(n13404) );
  OAI211_X1 U9675 ( .C1(n13373), .C2(n7739), .A(n13495), .B(n7644), .ZN(n7779)
         );
  NAND2_X1 U9676 ( .A1(n13373), .A2(n7739), .ZN(n7644) );
  NAND3_X1 U9677 ( .A1(n7645), .A2(n13977), .A3(n7646), .ZN(n13467) );
  INV_X1 U9678 ( .A(n7647), .ZN(n13356) );
  NAND2_X1 U9679 ( .A1(n11928), .A2(n7658), .ZN(n7656) );
  NAND2_X1 U9680 ( .A1(n8356), .A2(n13966), .ZN(n8355) );
  OAI211_X1 U9681 ( .C1(n13449), .C2(n7674), .A(n7671), .B(n8334), .ZN(n8331)
         );
  NAND2_X1 U9682 ( .A1(n8356), .A2(n7672), .ZN(n7671) );
  NAND2_X1 U9683 ( .A1(n8355), .A2(n13449), .ZN(n7673) );
  INV_X1 U9684 ( .A(n8056), .ZN(n7677) );
  NOR2_X2 U9685 ( .A1(n9632), .A2(n8459), .ZN(n9825) );
  AOI21_X1 U9686 ( .B1(n11648), .B2(n10598), .A(n10600), .ZN(n10640) );
  NAND2_X1 U9687 ( .A1(n8044), .A2(n8042), .ZN(n13303) );
  NAND2_X1 U9688 ( .A1(n8029), .A2(n8028), .ZN(n13993) );
  NAND2_X1 U9689 ( .A1(n9810), .A2(n13140), .ZN(n12434) );
  AOI21_X1 U9690 ( .B1(n14126), .B2(n16226), .A(n14125), .ZN(n14200) );
  XNOR2_X1 U9691 ( .A(n13914), .B(n13915), .ZN(n14126) );
  NAND2_X1 U9692 ( .A1(n11028), .A2(n9808), .ZN(n11478) );
  NAND2_X1 U9693 ( .A1(n11465), .A2(n13121), .ZN(n11620) );
  NAND2_X1 U9694 ( .A1(n11636), .A2(n13107), .ZN(n11029) );
  NAND2_X1 U9695 ( .A1(n11635), .A2(n13262), .ZN(n11636) );
  NAND2_X1 U9696 ( .A1(n7686), .A2(n7345), .ZN(P3_U3488) );
  OR2_X1 U9697 ( .A1(n9877), .A2(n7687), .ZN(n7686) );
  NAND2_X1 U9698 ( .A1(n7689), .A2(n7346), .ZN(P3_U3456) );
  OR2_X1 U9699 ( .A1(n9877), .A2(n16229), .ZN(n7689) );
  INV_X1 U9700 ( .A(n11892), .ZN(n7690) );
  NOR2_X2 U9701 ( .A1(n14612), .A2(n14613), .ZN(n14611) );
  NAND2_X1 U9702 ( .A1(n14736), .A2(n7746), .ZN(n14718) );
  NAND2_X1 U9703 ( .A1(n12399), .A2(n12405), .ZN(n12398) );
  NAND2_X1 U9704 ( .A1(n11596), .A2(n11597), .ZN(n11595) );
  NAND2_X1 U9705 ( .A1(n14790), .A2(n14789), .ZN(n14788) );
  NAND2_X1 U9706 ( .A1(n12328), .A2(n9040), .ZN(n12399) );
  NAND2_X1 U9707 ( .A1(n9253), .A2(n16208), .ZN(n9256) );
  NAND2_X1 U9708 ( .A1(n9124), .A2(n7260), .ZN(n9253) );
  NAND2_X1 U9709 ( .A1(n8630), .A2(n14484), .ZN(n8624) );
  OAI22_X1 U9710 ( .A1(n14631), .A2(n14630), .B1(n14401), .B2(n14641), .ZN(
        n14612) );
  NAND2_X1 U9711 ( .A1(n8132), .A2(n8133), .ZN(n7694) );
  NOR2_X1 U9712 ( .A1(n13810), .A2(n13811), .ZN(n13814) );
  NOR2_X1 U9713 ( .A1(n12458), .A2(n12459), .ZN(n12462) );
  XNOR2_X2 U9714 ( .A(n9380), .B(n9381), .ZN(n10526) );
  OR2_X2 U9715 ( .A1(n13859), .A2(n8166), .ZN(n13863) );
  OR2_X2 U9716 ( .A1(n10801), .A2(n10800), .ZN(n11013) );
  NOR2_X1 U9717 ( .A1(n10796), .A2(n10797), .ZN(n10801) );
  NOR2_X2 U9718 ( .A1(n11986), .A2(n11987), .ZN(n11989) );
  NOR2_X2 U9719 ( .A1(n11951), .A2(n9533), .ZN(n11986) );
  XNOR2_X1 U9720 ( .A(n9194), .B(n9192), .ZN(n15950) );
  NAND2_X1 U9721 ( .A1(n15991), .A2(n15990), .ZN(n7972) );
  NAND2_X1 U9722 ( .A1(n7970), .A2(n7971), .ZN(n7969) );
  XNOR2_X1 U9723 ( .A(n7969), .B(n7968), .ZN(SUB_1596_U4) );
  NAND2_X1 U9724 ( .A1(n12792), .A2(n12791), .ZN(n12796) );
  NAND2_X1 U9725 ( .A1(n7698), .A2(n8310), .ZN(n12932) );
  NAND2_X1 U9726 ( .A1(n14760), .A2(n9046), .ZN(n14737) );
  NAND2_X1 U9727 ( .A1(n8382), .A2(n8380), .ZN(n8746) );
  NAND2_X1 U9728 ( .A1(n9247), .A2(n14948), .ZN(n7789) );
  AOI21_X1 U9729 ( .B1(n14573), .B2(n14884), .A(n7703), .ZN(n14575) );
  NAND2_X1 U9730 ( .A1(n11595), .A2(n9032), .ZN(n11420) );
  INV_X1 U9731 ( .A(n9239), .ZN(n8138) );
  MUX2_X1 U9732 ( .A(n10488), .B(P3_REG2_REG_2__SCAN_IN), .S(n10522), .Z(
        n10546) );
  NAND2_X1 U9733 ( .A1(n12804), .A2(n12803), .ZN(n12807) );
  NAND2_X1 U9734 ( .A1(n7789), .A2(n7786), .ZN(P2_U3494) );
  NAND2_X1 U9735 ( .A1(n15578), .A2(n15398), .ZN(n15562) );
  NAND2_X1 U9736 ( .A1(n11235), .A2(n8180), .ZN(n8181) );
  NAND2_X1 U9737 ( .A1(n8195), .A2(n8194), .ZN(n15533) );
  OAI21_X1 U9738 ( .B1(n15523), .B2(n8202), .A(n8200), .ZN(n15481) );
  NAND2_X1 U9739 ( .A1(n15605), .A2(n8208), .ZN(n15578) );
  OAI22_X2 U9740 ( .A1(n12155), .A2(n9510), .B1(n12238), .B2(n16142), .ZN(
        n12252) );
  NAND2_X1 U9741 ( .A1(n11031), .A2(n11032), .ZN(n11030) );
  NAND2_X1 U9742 ( .A1(n15141), .A2(n8268), .ZN(n7800) );
  AOI21_X1 U9743 ( .B1(n14982), .B2(n14981), .A(n14980), .ZN(n14988) );
  INV_X1 U9744 ( .A(n8283), .ZN(n8282) );
  NOR2_X1 U9745 ( .A1(n12374), .A2(n8284), .ZN(n8283) );
  AOI21_X2 U9746 ( .B1(n15132), .B2(n15133), .A(n7279), .ZN(n15141) );
  INV_X1 U9747 ( .A(n10738), .ZN(n8344) );
  INV_X1 U9748 ( .A(n7793), .ZN(n10740) );
  INV_X1 U9749 ( .A(n10956), .ZN(n13102) );
  NAND2_X1 U9750 ( .A1(n11299), .A2(n11298), .ZN(n11300) );
  NAND2_X1 U9751 ( .A1(n9822), .A2(n9829), .ZN(n11891) );
  NAND2_X1 U9752 ( .A1(n13478), .A2(n13477), .ZN(n13476) );
  NAND3_X1 U9753 ( .A1(n7764), .A2(n7213), .A3(n7317), .ZN(P1_U3242) );
  OR2_X1 U9754 ( .A1(n12749), .A2(n10864), .ZN(n10705) );
  AND2_X1 U9755 ( .A1(n12761), .A2(n13011), .ZN(n7737) );
  NAND2_X1 U9756 ( .A1(n7715), .A2(n8632), .ZN(n11405) );
  NAND2_X1 U9757 ( .A1(n13356), .A2(n13415), .ZN(n13358) );
  NAND2_X1 U9758 ( .A1(n7716), .A2(n7717), .ZN(n7715) );
  NOR2_X1 U9759 ( .A1(n7725), .A2(n7724), .ZN(n7723) );
  NAND2_X1 U9760 ( .A1(n8624), .A2(n9027), .ZN(n7716) );
  OR2_X1 U9761 ( .A1(n8699), .A2(n10207), .ZN(n8660) );
  INV_X1 U9762 ( .A(n11391), .ZN(n7717) );
  NAND2_X1 U9763 ( .A1(n14692), .A2(n14693), .ZN(n8152) );
  NAND2_X1 U9764 ( .A1(n8662), .A2(n8661), .ZN(n11598) );
  INV_X1 U9765 ( .A(n7716), .ZN(n9026) );
  AND2_X2 U9766 ( .A1(n14662), .A2(n14654), .ZN(n14651) );
  AND2_X2 U9767 ( .A1(n14676), .A2(n14925), .ZN(n14662) );
  NOR2_X4 U9768 ( .A1(n14603), .A2(n14819), .ZN(n14581) );
  INV_X1 U9769 ( .A(n10980), .ZN(n8630) );
  NAND2_X1 U9770 ( .A1(n8959), .A2(n8958), .ZN(n14610) );
  NAND2_X1 U9771 ( .A1(n11620), .A2(n13124), .ZN(n11619) );
  NAND2_X1 U9772 ( .A1(n11029), .A2(n13265), .ZN(n11028) );
  XNOR2_X1 U9773 ( .A(n13111), .B(n7730), .ZN(n13265) );
  NAND2_X1 U9774 ( .A1(n11477), .A2(n13114), .ZN(n11466) );
  NAND2_X1 U9775 ( .A1(n7735), .A2(n7734), .ZN(n7733) );
  OAI21_X1 U9776 ( .B1(n13004), .B2(n12736), .A(n15109), .ZN(n12740) );
  NAND2_X4 U9777 ( .A1(n12735), .A2(n13048), .ZN(n13051) );
  NAND2_X1 U9778 ( .A1(n8483), .A2(n8416), .ZN(n8415) );
  NOR2_X2 U9779 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8480) );
  NAND2_X1 U9780 ( .A1(n7939), .A2(n7943), .ZN(n7935) );
  NAND2_X1 U9781 ( .A1(n7934), .A2(n7936), .ZN(n10542) );
  NOR2_X1 U9782 ( .A1(n12303), .A2(n9571), .ZN(n12458) );
  NOR2_X1 U9783 ( .A1(n13790), .A2(n14185), .ZN(n13810) );
  INV_X1 U9784 ( .A(n13863), .ZN(n7744) );
  XNOR2_X2 U9785 ( .A(n7732), .B(n11965), .ZN(n11951) );
  NOR2_X1 U9786 ( .A1(n13913), .A2(n14182), .ZN(n9821) );
  INV_X1 U9787 ( .A(n9792), .ZN(n9791) );
  NAND2_X1 U9788 ( .A1(n9786), .A2(n9785), .ZN(n9792) );
  INV_X1 U9789 ( .A(n12846), .ZN(n7734) );
  INV_X1 U9790 ( .A(n12845), .ZN(n7735) );
  NAND2_X1 U9791 ( .A1(n12844), .A2(n12843), .ZN(n7736) );
  AND3_X2 U9792 ( .A1(n10703), .A2(n10704), .A3(n10702), .ZN(n12749) );
  NAND2_X1 U9793 ( .A1(n7738), .A2(n7737), .ZN(n12768) );
  NAND2_X1 U9794 ( .A1(n12756), .A2(n12755), .ZN(n7738) );
  INV_X1 U9795 ( .A(n14299), .ZN(n7847) );
  NOR2_X1 U9796 ( .A1(n7224), .A2(n7325), .ZN(n7863) );
  NAND2_X1 U9797 ( .A1(n7851), .A2(n7850), .ZN(n14372) );
  NAND2_X1 U9798 ( .A1(n8512), .A2(n8516), .ZN(n7766) );
  OAI21_X1 U9799 ( .B1(n9176), .B2(n9175), .A(n7777), .ZN(n7776) );
  AND2_X2 U9800 ( .A1(n8610), .A2(n8609), .ZN(n8885) );
  NAND2_X1 U9801 ( .A1(n7758), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8606) );
  OR2_X1 U9802 ( .A1(n10563), .A2(n10484), .ZN(n10564) );
  NAND2_X1 U9803 ( .A1(n10564), .A2(n10515), .ZN(n10541) );
  NAND2_X1 U9804 ( .A1(n11533), .A2(n11532), .ZN(n11699) );
  INV_X1 U9805 ( .A(n7922), .ZN(n13859) );
  NAND2_X1 U9806 ( .A1(n8515), .A2(n9260), .ZN(n7742) );
  OAI21_X1 U9807 ( .B1(n12072), .B2(n8072), .A(n8070), .ZN(n12186) );
  NAND2_X2 U9808 ( .A1(n12191), .A2(n12190), .ZN(n12518) );
  NAND2_X1 U9809 ( .A1(n15646), .A2(n7783), .ZN(n15744) );
  NAND2_X1 U9810 ( .A1(n8621), .A2(n8517), .ZN(n7773) );
  NAND2_X1 U9811 ( .A1(n7773), .A2(SI_2_), .ZN(n8521) );
  NAND2_X1 U9812 ( .A1(n15536), .A2(n15535), .ZN(n15534) );
  NAND2_X2 U9813 ( .A1(n10521), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n13778) );
  NOR2_X2 U9814 ( .A1(n13780), .A2(n7745), .ZN(n10521) );
  AND2_X2 U9815 ( .A1(n15442), .A2(n15723), .ZN(n7785) );
  NOR2_X1 U9816 ( .A1(n11989), .A2(n11988), .ZN(n12302) );
  NAND4_X2 U9817 ( .A1(n10413), .A2(n10414), .A3(n10415), .A4(n10412), .ZN(
        n12736) );
  NOR2_X1 U9818 ( .A1(n15379), .A2(n8472), .ZN(n15433) );
  NAND2_X1 U9819 ( .A1(n11598), .A2(n8681), .ZN(n7747) );
  NAND2_X1 U9820 ( .A1(n8358), .A2(n14250), .ZN(n8357) );
  NAND2_X1 U9821 ( .A1(n13484), .A2(n13372), .ZN(n13373) );
  NAND2_X1 U9822 ( .A1(n8637), .A2(n8638), .ZN(n8642) );
  NAND2_X1 U9823 ( .A1(n8120), .A2(n8119), .ZN(n14682) );
  NAND4_X1 U9824 ( .A1(n8798), .A2(n8412), .A3(n8136), .A4(n7211), .ZN(n8607)
         );
  INV_X1 U9825 ( .A(n8609), .ZN(n8611) );
  NAND2_X1 U9826 ( .A1(n8798), .A2(n8412), .ZN(n7750) );
  NAND2_X1 U9827 ( .A1(n7751), .A2(n7313), .ZN(n9975) );
  NAND3_X1 U9828 ( .A1(n9969), .A2(n9968), .A3(n7308), .ZN(n7751) );
  OAI21_X1 U9829 ( .B1(n9919), .B2(n9918), .A(n8249), .ZN(n8247) );
  NAND3_X1 U9830 ( .A1(n9934), .A2(n9933), .A3(n7330), .ZN(n7753) );
  AOI22_X1 U9831 ( .A1(n9964), .A2(n9963), .B1(n9961), .B2(n9962), .ZN(n9967)
         );
  NAND2_X1 U9832 ( .A1(n10244), .A2(n9846), .ZN(n9848) );
  NAND2_X1 U9833 ( .A1(n7792), .A2(n9858), .ZN(n9845) );
  NAND2_X1 U9834 ( .A1(n10546), .A2(n10545), .ZN(n10544) );
  XNOR2_X1 U9835 ( .A(n12450), .B(n12466), .ZN(n12301) );
  NAND3_X1 U9836 ( .A1(n8798), .A2(n7211), .A3(n8412), .ZN(n7758) );
  NAND2_X1 U9837 ( .A1(n9253), .A2(n14948), .ZN(n7770) );
  NAND2_X1 U9838 ( .A1(n14660), .A2(n14667), .ZN(n7759) );
  NAND2_X1 U9839 ( .A1(n8518), .A2(n8519), .ZN(n8621) );
  AND2_X1 U9840 ( .A1(n8183), .A2(n11234), .ZN(n8180) );
  OAI21_X2 U9841 ( .B1(n11122), .B2(n12987), .A(n11121), .ZN(n12762) );
  NAND2_X1 U9842 ( .A1(n7760), .A2(n8312), .ZN(n12885) );
  NAND3_X1 U9843 ( .A1(n12821), .A2(n7761), .A3(n7323), .ZN(n8292) );
  NAND2_X1 U9844 ( .A1(n12819), .A2(n12820), .ZN(n7761) );
  NAND2_X1 U9845 ( .A1(n7763), .A2(n7762), .ZN(n12756) );
  NAND2_X1 U9846 ( .A1(n12740), .A2(n12739), .ZN(n7763) );
  NAND2_X1 U9847 ( .A1(n13077), .A2(n13075), .ZN(n7764) );
  NAND2_X1 U9848 ( .A1(n9791), .A2(n9793), .ZN(n9788) );
  NAND2_X1 U9849 ( .A1(n9825), .A2(n9336), .ZN(n9822) );
  OAI21_X1 U9850 ( .B1(n9632), .B2(n7321), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9824) );
  AND3_X1 U9851 ( .A1(n7766), .A2(n8514), .A3(n8513), .ZN(n8637) );
  AOI21_X1 U9852 ( .B1(n8122), .B2(n8128), .A(n7226), .ZN(n8119) );
  NAND2_X1 U9853 ( .A1(n7770), .A2(n7768), .ZN(P2_U3496) );
  NOR2_X2 U9854 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n8479) );
  INV_X1 U9855 ( .A(n16029), .ZN(n8055) );
  NOR2_X1 U9856 ( .A1(n15950), .A2(n15951), .ZN(n15949) );
  NOR2_X1 U9857 ( .A1(n9821), .A2(n13907), .ZN(n9877) );
  INV_X1 U9858 ( .A(n8045), .ZN(n13296) );
  OAI21_X1 U9859 ( .B1(n15976), .B2(n15975), .A(n7961), .ZN(n7960) );
  XNOR2_X1 U9860 ( .A(n7774), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9861 ( .A1(n15991), .A2(n15990), .ZN(n7775) );
  INV_X1 U9862 ( .A(n15963), .ZN(n7964) );
  NAND2_X2 U9863 ( .A1(n9405), .A2(n9343), .ZN(n9705) );
  NOR2_X1 U9864 ( .A1(n12301), .A2(n12642), .ZN(n12451) );
  NAND2_X1 U9865 ( .A1(n7779), .A2(n7340), .ZN(P3_U3154) );
  NOR2_X2 U9866 ( .A1(n15441), .A2(n7785), .ZN(n15646) );
  INV_X1 U9867 ( .A(n8182), .ZN(n8179) );
  NAND2_X1 U9868 ( .A1(n14788), .A2(n9043), .ZN(n14771) );
  NAND2_X1 U9869 ( .A1(n8153), .A2(n8915), .ZN(n14660) );
  NAND2_X1 U9870 ( .A1(n9830), .A2(n11891), .ZN(n7792) );
  NAND2_X1 U9871 ( .A1(n7202), .A2(n13342), .ZN(n13478) );
  NAND2_X1 U9872 ( .A1(n8318), .A2(n8316), .ZN(n13334) );
  NAND3_X1 U9873 ( .A1(n8159), .A2(n10530), .A3(P3_REG2_REG_3__SCAN_IN), .ZN(
        n10622) );
  INV_X1 U9874 ( .A(n8624), .ZN(n8129) );
  NAND2_X1 U9875 ( .A1(n8129), .A2(n9027), .ZN(n8130) );
  INV_X1 U9876 ( .A(n7799), .ZN(n7798) );
  NAND2_X1 U9877 ( .A1(n7800), .A2(n8266), .ZN(n15010) );
  NAND2_X1 U9878 ( .A1(n15207), .A2(n7801), .ZN(n15132) );
  OR2_X1 U9879 ( .A1(n14988), .A2(n14987), .ZN(n7801) );
  NAND2_X1 U9880 ( .A1(n7803), .A2(n11774), .ZN(n7802) );
  NAND2_X1 U9881 ( .A1(n8275), .A2(n7818), .ZN(n7817) );
  OAI211_X1 U9882 ( .C1(n8275), .C2(n7819), .A(n15104), .B(n7817), .ZN(
        P1_U3220) );
  NAND2_X1 U9883 ( .A1(n8275), .A2(n8274), .ZN(n15093) );
  INV_X1 U9884 ( .A(n8280), .ZN(n7837) );
  NAND2_X1 U9885 ( .A1(n12580), .A2(n12581), .ZN(n7842) );
  NAND4_X1 U9886 ( .A1(n9230), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n16001), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7843) );
  NAND4_X1 U9887 ( .A1(n15348), .A2(n16000), .A3(n7845), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7844) );
  NAND2_X1 U9888 ( .A1(n8516), .A2(n8518), .ZN(n8511) );
  NAND2_X1 U9889 ( .A1(n14335), .A2(n7848), .ZN(n7851) );
  NAND2_X1 U9890 ( .A1(n14372), .A2(n14371), .ZN(n14370) );
  NAND2_X1 U9891 ( .A1(n7853), .A2(n7852), .ZN(n11881) );
  OAI21_X1 U9892 ( .B1(n7855), .B2(n7203), .A(n11879), .ZN(n7854) );
  NAND2_X1 U9893 ( .A1(n14379), .A2(n7864), .ZN(n7862) );
  NAND2_X1 U9894 ( .A1(n7863), .A2(n7862), .ZN(n14430) );
  INV_X1 U9895 ( .A(n7333), .ZN(n14323) );
  NAND2_X1 U9896 ( .A1(n8781), .A2(n7877), .ZN(n7875) );
  NAND2_X1 U9897 ( .A1(n8558), .A2(n7890), .ZN(n7889) );
  NAND2_X1 U9898 ( .A1(n8558), .A2(n13630), .ZN(n8383) );
  OR2_X1 U9899 ( .A1(n8558), .A2(n13630), .ZN(n8384) );
  OAI21_X1 U9900 ( .B1(n10019), .B2(n7230), .A(n7895), .ZN(n7894) );
  INV_X1 U9901 ( .A(n13079), .ZN(n10025) );
  NAND2_X1 U9902 ( .A1(n7223), .A2(n8673), .ZN(n7898) );
  NAND3_X1 U9903 ( .A1(n7898), .A2(n8534), .A3(n7897), .ZN(n8536) );
  NAND4_X1 U9904 ( .A1(n10092), .A2(n7908), .A3(n10111), .A4(n7907), .ZN(n7906) );
  NAND3_X1 U9905 ( .A1(n10110), .A2(n14629), .A3(n10109), .ZN(n7909) );
  NOR2_X2 U9906 ( .A1(n11594), .A2(n11603), .ZN(n11593) );
  INV_X1 U9907 ( .A(n11411), .ZN(n7911) );
  NAND2_X1 U9908 ( .A1(n7912), .A2(n14581), .ZN(n14552) );
  NOR2_X2 U9909 ( .A1(n14802), .A2(n14889), .ZN(n14774) );
  OR2_X2 U9910 ( .A1(n14801), .A2(n14800), .ZN(n14802) );
  AND2_X2 U9911 ( .A1(n12145), .A2(n12425), .ZN(n12401) );
  NOR2_X2 U9912 ( .A1(n14711), .A2(n14700), .ZN(n14696) );
  NAND2_X2 U9913 ( .A1(n14724), .A2(n14861), .ZN(n14711) );
  AND2_X2 U9914 ( .A1(n14745), .A2(n14728), .ZN(n14724) );
  AND2_X2 U9915 ( .A1(n14763), .A2(n14872), .ZN(n14745) );
  AND2_X2 U9916 ( .A1(n13789), .A2(n13788), .ZN(n13809) );
  NAND4_X1 U9917 ( .A1(n7932), .A2(n13864), .A3(n7931), .A4(n13865), .ZN(n7927) );
  AOI21_X1 U9918 ( .B1(n13864), .B2(n13863), .A(n13862), .ZN(n13880) );
  NAND2_X1 U9919 ( .A1(n10541), .A2(n10542), .ZN(n10540) );
  NAND2_X1 U9920 ( .A1(n7939), .A2(n7937), .ZN(n7936) );
  OAI211_X1 U9921 ( .C1(n13778), .C2(n7950), .A(n7944), .B(n7945), .ZN(n10669)
         );
  NAND3_X1 U9922 ( .A1(n10668), .A2(n7948), .A3(n13778), .ZN(n7944) );
  NOR2_X1 U9923 ( .A1(n10669), .A2(n10658), .ZN(n10796) );
  NAND3_X1 U9924 ( .A1(n10668), .A2(n13778), .A3(n7956), .ZN(n7954) );
  AND2_X2 U9925 ( .A1(n7964), .A2(n7963), .ZN(n9209) );
  XNOR2_X2 U9926 ( .A(n7965), .B(n9199), .ZN(n15954) );
  OR2_X2 U9927 ( .A1(n15949), .A2(n9195), .ZN(n7965) );
  NAND2_X1 U9928 ( .A1(n15943), .A2(n15942), .ZN(n15941) );
  NAND2_X1 U9929 ( .A1(n15941), .A2(n9183), .ZN(n15944) );
  XNOR2_X1 U9930 ( .A(n9169), .B(n7973), .ZN(n9172) );
  NAND2_X1 U9931 ( .A1(n9519), .A2(n7978), .ZN(n7977) );
  NAND2_X1 U9932 ( .A1(n9662), .A2(n7985), .ZN(n7984) );
  NAND2_X1 U9933 ( .A1(n9613), .A2(n7992), .ZN(n7991) );
  NAND2_X1 U9934 ( .A1(n9430), .A2(n7999), .ZN(n7995) );
  NAND2_X1 U9935 ( .A1(n7995), .A2(n7996), .ZN(n9454) );
  NAND3_X1 U9936 ( .A1(n8009), .A2(n8010), .A3(P1_DATAO_REG_13__SCAN_IN), .ZN(
        n9564) );
  NAND2_X1 U9937 ( .A1(n8009), .A2(n8010), .ZN(n9562) );
  AND2_X2 U9938 ( .A1(n11348), .A2(n11385), .ZN(n11538) );
  NOR2_X2 U9939 ( .A1(n11358), .A2(n12762), .ZN(n11357) );
  INV_X2 U9940 ( .A(n12757), .ZN(n8021) );
  NOR2_X2 U9941 ( .A1(n12528), .A2(n15733), .ZN(n8026) );
  NOR2_X2 U9942 ( .A1(n15592), .A2(n15698), .ZN(n15568) );
  INV_X1 U9943 ( .A(n13961), .ZN(n8036) );
  INV_X1 U9944 ( .A(n12101), .ZN(n8037) );
  NAND2_X1 U9945 ( .A1(n8038), .A2(n7225), .ZN(n9810) );
  NAND3_X1 U9946 ( .A1(n13928), .A2(n8047), .A3(n7208), .ZN(n8044) );
  NAND2_X1 U9947 ( .A1(n13094), .A2(n13207), .ZN(n8050) );
  XNOR2_X1 U9948 ( .A(n13523), .B(n8055), .ZN(n16031) );
  NOR2_X2 U9949 ( .A1(n11427), .A2(n10141), .ZN(n8057) );
  INV_X2 U9950 ( .A(n12736), .ZN(n10845) );
  NAND2_X1 U9951 ( .A1(n12744), .A2(n12745), .ZN(n10717) );
  NAND2_X1 U9952 ( .A1(n12737), .A2(n12736), .ZN(n12745) );
  NAND2_X1 U9953 ( .A1(n11699), .A2(n8062), .ZN(n8059) );
  NAND2_X1 U9954 ( .A1(n8059), .A2(n8060), .ZN(n12069) );
  NAND2_X1 U9955 ( .A1(n10368), .A2(n8074), .ZN(n8081) );
  NAND3_X1 U9956 ( .A1(n8081), .A2(n8079), .A3(n8075), .ZN(n10371) );
  OAI21_X1 U9957 ( .B1(n15566), .B2(n8095), .A(n8093), .ZN(n15536) );
  NAND2_X1 U9958 ( .A1(n12518), .A2(n8101), .ZN(n8097) );
  NAND2_X1 U9959 ( .A1(n8097), .A2(n8099), .ZN(n12661) );
  NAND2_X1 U9960 ( .A1(n10754), .A2(n10753), .ZN(n11238) );
  NOR2_X1 U9961 ( .A1(n8205), .A2(n15516), .ZN(n15515) );
  NAND2_X1 U9962 ( .A1(n11241), .A2(n12767), .ZN(n11342) );
  NAND2_X1 U9963 ( .A1(n11342), .A2(n11341), .ZN(n11343) );
  OAI21_X2 U9964 ( .B1(n11238), .B2(n11237), .A(n11236), .ZN(n11355) );
  AOI21_X2 U9965 ( .B1(n11240), .B2(n7240), .A(n8470), .ZN(n11241) );
  NAND2_X1 U9966 ( .A1(n13244), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U9967 ( .A1(n12433), .A2(n13144), .ZN(n12479) );
  NAND2_X1 U9968 ( .A1(n9378), .A2(n9261), .ZN(n9402) );
  NAND2_X1 U9969 ( .A1(n9320), .A2(n9319), .ZN(n9757) );
  INV_X1 U9970 ( .A(n11355), .ZN(n11240) );
  NAND2_X1 U9971 ( .A1(n14722), .A2(n8122), .ZN(n8120) );
  INV_X1 U9972 ( .A(n9027), .ZN(n8131) );
  NAND2_X1 U9973 ( .A1(n11660), .A2(n7236), .ZN(n8132) );
  AND2_X2 U9974 ( .A1(n8611), .A2(n8610), .ZN(n8649) );
  NAND2_X1 U9975 ( .A1(n8139), .A2(n8655), .ZN(n8524) );
  INV_X1 U9976 ( .A(n12406), .ZN(n8144) );
  NAND2_X1 U9977 ( .A1(n8152), .A2(n8150), .ZN(n8153) );
  NAND2_X1 U9978 ( .A1(n10544), .A2(n10528), .ZN(n8160) );
  NAND3_X1 U9979 ( .A1(n8163), .A2(n13772), .A3(n7227), .ZN(n8161) );
  NAND2_X1 U9980 ( .A1(n8163), .A2(n13772), .ZN(n10532) );
  NAND2_X1 U9981 ( .A1(n7291), .A2(n10519), .ZN(n8163) );
  NAND2_X1 U9982 ( .A1(n15418), .A2(n15411), .ZN(n8177) );
  NAND2_X1 U9983 ( .A1(n8181), .A2(n8178), .ZN(n11339) );
  NAND2_X1 U9984 ( .A1(n15465), .A2(n8192), .ZN(n8190) );
  NAND2_X1 U9985 ( .A1(n15562), .A2(n7319), .ZN(n8195) );
  INV_X1 U9986 ( .A(n15523), .ZN(n8206) );
  NAND3_X1 U9987 ( .A1(n10012), .A2(n10008), .A3(n10013), .ZN(n8211) );
  NAND2_X2 U9988 ( .A1(n10034), .A2(n8212), .ZN(n10050) );
  NAND2_X2 U9989 ( .A1(n10115), .A2(n8212), .ZN(n10832) );
  INV_X1 U9990 ( .A(n9094), .ZN(n8212) );
  NAND2_X1 U9991 ( .A1(n8229), .A2(n8230), .ZN(n9949) );
  NAND3_X1 U9992 ( .A1(n9945), .A2(n7310), .A3(n9944), .ZN(n8229) );
  OAI211_X1 U9993 ( .C1(n10124), .C2(n8234), .A(n10130), .B(n8232), .ZN(
        P2_U3328) );
  NAND2_X1 U9994 ( .A1(n9940), .A2(n9941), .ZN(n9939) );
  NAND3_X1 U9995 ( .A1(n9996), .A2(n9995), .A3(n7311), .ZN(n8241) );
  INV_X1 U9996 ( .A(n9923), .ZN(n8244) );
  AND2_X1 U9997 ( .A1(n8248), .A2(n8246), .ZN(n8245) );
  OAI21_X1 U9998 ( .B1(n15169), .B2(n8256), .A(n8253), .ZN(n15149) );
  NAND2_X1 U9999 ( .A1(n8252), .A2(n8250), .ZN(n15046) );
  NAND2_X1 U10000 ( .A1(n15169), .A2(n8253), .ZN(n8252) );
  NAND2_X1 U10001 ( .A1(n8259), .A2(n8258), .ZN(n8257) );
  NAND2_X1 U10002 ( .A1(n8262), .A2(n8260), .ZN(n11188) );
  OAI21_X1 U10003 ( .B1(n15141), .B2(n8270), .A(n8268), .ZN(n15082) );
  OAI21_X1 U10004 ( .B1(n15141), .B2(n15142), .A(n8273), .ZN(n15188) );
  INV_X1 U10005 ( .A(n12372), .ZN(n8286) );
  OR2_X2 U10006 ( .A1(n12733), .A2(n12731), .ZN(n8288) );
  INV_X1 U10007 ( .A(n10420), .ZN(n8287) );
  INV_X2 U10008 ( .A(n13000), .ZN(n12836) );
  NAND2_X1 U10009 ( .A1(n8289), .A2(n8290), .ZN(n12782) );
  NAND2_X1 U10010 ( .A1(n8292), .A2(n8293), .ZN(n12840) );
  NAND2_X1 U10011 ( .A1(n12798), .A2(n8296), .ZN(n8295) );
  NAND2_X1 U10012 ( .A1(n8298), .A2(n8299), .ZN(n12818) );
  NAND2_X1 U10013 ( .A1(n12356), .A2(n8319), .ZN(n8318) );
  NAND2_X1 U10014 ( .A1(n8331), .A2(n7262), .ZN(n13484) );
  AND2_X1 U10015 ( .A1(n8342), .A2(n8341), .ZN(n11102) );
  OAI211_X1 U10016 ( .C1(n13404), .C2(n8347), .A(n8345), .B(n13413), .ZN(
        P3_U3160) );
  NAND2_X1 U10017 ( .A1(n13404), .A2(n8346), .ZN(n8345) );
  INV_X1 U10018 ( .A(n13293), .ZN(n8358) );
  NAND2_X1 U10019 ( .A1(n8540), .A2(n7210), .ZN(n8380) );
  INV_X2 U10020 ( .A(n7560), .ZN(n10178) );
  MUX2_X1 U10021 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n9343), .Z(n8392) );
  INV_X1 U10022 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8394) );
  OAI21_X2 U10023 ( .B1(n8396), .B2(n11090), .A(n8395), .ZN(n11505) );
  NAND2_X1 U10024 ( .A1(n14442), .A2(n8410), .ZN(n14349) );
  NAND2_X1 U10025 ( .A1(n8798), .A2(n8414), .ZN(n8585) );
  INV_X2 U10026 ( .A(n8420), .ZN(n13244) );
  INV_X1 U10027 ( .A(n8418), .ZN(n8417) );
  OAI22_X1 U10028 ( .A1(n8420), .A2(n8419), .B1(n10484), .B2(n9407), .ZN(n8418) );
  NAND2_X1 U10029 ( .A1(n8421), .A2(n8423), .ZN(n9610) );
  INV_X1 U10030 ( .A(n9717), .ZN(n13987) );
  NAND2_X1 U10031 ( .A1(n12252), .A2(n13268), .ZN(n8444) );
  OAI21_X1 U10032 ( .B1(n13951), .B2(n8446), .A(n8445), .ZN(n8453) );
  NOR2_X1 U10033 ( .A1(n13951), .A2(n8455), .ZN(n13941) );
  AND2_X1 U10034 ( .A1(n13364), .A2(n13511), .ZN(n8455) );
  NAND2_X1 U10035 ( .A1(n11621), .A2(n7228), .ZN(n12102) );
  NAND3_X1 U10036 ( .A1(n11030), .A2(n9433), .A3(n13261), .ZN(n11479) );
  OAI21_X1 U10037 ( .B1(n15647), .B2(n16002), .A(n15440), .ZN(n15441) );
  INV_X1 U10038 ( .A(n15163), .ZN(n15016) );
  NAND2_X1 U10039 ( .A1(n15010), .A2(n15009), .ZN(n15163) );
  INV_X1 U10040 ( .A(n10378), .ZN(n10143) );
  OAI21_X1 U10041 ( .B1(n15640), .B2(n15732), .A(n15639), .ZN(n15641) );
  NAND2_X1 U10042 ( .A1(n15418), .A2(n15417), .ZN(n15640) );
  NAND2_X1 U10043 ( .A1(n12734), .A2(n12733), .ZN(n13048) );
  NAND2_X1 U10044 ( .A1(n12973), .A2(n12974), .ZN(n12978) );
  NAND2_X1 U10045 ( .A1(n11804), .A2(n11803), .ZN(n12085) );
  INV_X1 U10046 ( .A(n12991), .ZN(n15779) );
  INV_X1 U10047 ( .A(n12730), .ZN(n15343) );
  NAND2_X1 U10048 ( .A1(n15208), .A2(n15209), .ZN(n15207) );
  INV_X2 U10049 ( .A(n8515), .ZN(n9343) );
  AND2_X1 U10050 ( .A1(n14484), .A2(n14350), .ZN(n10982) );
  AOI211_X1 U10051 ( .C1(n16190), .C2(n16189), .A(n16188), .B(n16187), .ZN(
        n16192) );
  NAND2_X1 U10052 ( .A1(n14948), .A2(n16190), .ZN(n14953) );
  NAND2_X1 U10053 ( .A1(n16208), .A2(n16190), .ZN(n14897) );
  NAND2_X1 U10054 ( .A1(n13922), .A2(n13921), .ZN(n14125) );
  NAND2_X1 U10055 ( .A1(n14483), .A2(n10055), .ZN(n9891) );
  NAND2_X1 U10056 ( .A1(n10055), .A2(n11399), .ZN(n9884) );
  NAND2_X1 U10057 ( .A1(n10047), .A2(n10092), .ZN(n10070) );
  OR2_X1 U10058 ( .A1(n15416), .A2(n15415), .ZN(n15417) );
  OR2_X1 U10059 ( .A1(n16094), .A2(n9093), .ZN(n14751) );
  CLKBUF_X1 U10060 ( .A(n11641), .Z(n13258) );
  INV_X1 U10061 ( .A(n10115), .ZN(n9093) );
  NAND2_X1 U10062 ( .A1(n12102), .A2(n9494), .ZN(n12155) );
  AND2_X1 U10063 ( .A1(n10981), .A2(n10982), .ZN(n10983) );
  NAND2_X1 U10064 ( .A1(n9959), .A2(n9958), .ZN(n9964) );
  AND2_X1 U10065 ( .A1(n15435), .A2(n15434), .ZN(n15436) );
  NOR2_X1 U10066 ( .A1(n10983), .A2(n10984), .ZN(n11222) );
  INV_X1 U10067 ( .A(n13029), .ZN(n12658) );
  AND2_X1 U10068 ( .A1(n12747), .A2(n13012), .ZN(n8462) );
  INV_X2 U10069 ( .A(n16052), .ZN(n16131) );
  AND2_X2 U10070 ( .A1(n11061), .A2(n16128), .ZN(n16052) );
  INV_X1 U10071 ( .A(n14192), .ZN(n9879) );
  INV_X1 U10072 ( .A(n14948), .ZN(n16209) );
  AND2_X1 U10073 ( .A1(n10721), .A2(n10720), .ZN(n16074) );
  INV_X1 U10074 ( .A(n16074), .ZN(n15723) );
  INV_X1 U10075 ( .A(n13412), .ZN(n14203) );
  NAND2_X1 U10076 ( .A1(n16232), .A2(n16054), .ZN(n14246) );
  AND2_X1 U10077 ( .A1(n9251), .A2(n14465), .ZN(n8466) );
  OR2_X1 U10078 ( .A1(n9251), .A2(n14951), .ZN(n8467) );
  AND4_X1 U10079 ( .A1(n10212), .A2(n10147), .A3(n10146), .A4(n10211), .ZN(
        n8469) );
  AND2_X1 U10080 ( .A1(n11239), .A2(n12762), .ZN(n8470) );
  AND3_X1 U10081 ( .A1(n8488), .A2(n8487), .A3(n8486), .ZN(n8471) );
  INV_X1 U10082 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n14251) );
  INV_X1 U10083 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n14456) );
  AND2_X1 U10084 ( .A1(n15648), .A2(n15439), .ZN(n8472) );
  CLKBUF_X1 U10085 ( .A(n10650), .Z(n14252) );
  OR2_X1 U10086 ( .A1(n14218), .A2(n13978), .ZN(n8473) );
  INV_X1 U10087 ( .A(n13978), .ZN(n13512) );
  XNOR2_X1 U10088 ( .A(n13086), .B(n9107), .ZN(n10112) );
  NOR2_X1 U10089 ( .A1(n13943), .A2(n16034), .ZN(n8474) );
  INV_X1 U10090 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n13419) );
  AND2_X1 U10091 ( .A1(n10059), .A2(n10058), .ZN(n8475) );
  INV_X1 U10092 ( .A(n10371), .ZN(n13078) );
  OR2_X1 U10093 ( .A1(n13432), .A2(n13445), .ZN(n8476) );
  INV_X1 U10094 ( .A(n14728), .ZN(n14867) );
  OAI21_X1 U10095 ( .B1(n10007), .B2(n10006), .A(n10005), .ZN(n10012) );
  NAND2_X1 U10096 ( .A1(n11724), .A2(n10050), .ZN(n9890) );
  OAI22_X1 U10097 ( .A1(n12295), .A2(n7194), .B1(n11679), .B2(n10073), .ZN(
        n9927) );
  INV_X1 U10098 ( .A(n9941), .ZN(n9942) );
  NAND2_X1 U10099 ( .A1(n9943), .A2(n9942), .ZN(n9944) );
  OAI22_X1 U10100 ( .A1(n12425), .A2(n7194), .B1(n12499), .B2(n10073), .ZN(
        n9953) );
  INV_X1 U10101 ( .A(n12841), .ZN(n12842) );
  NAND2_X1 U10102 ( .A1(n7287), .A2(n7370), .ZN(n9995) );
  OAI22_X1 U10103 ( .A1(n14654), .A2(n7194), .B1(n14362), .B2(n10073), .ZN(
        n9997) );
  OAI22_X1 U10104 ( .A1(n14914), .A2(n10085), .B1(n14401), .B2(n7194), .ZN(
        n10001) );
  INV_X1 U10105 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9327) );
  INV_X1 U10106 ( .A(n13932), .ZN(n9769) );
  INV_X1 U10107 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U10108 ( .A1(n13301), .A2(n14119), .ZN(n13302) );
  NAND2_X1 U10109 ( .A1(n14218), .A2(n13978), .ZN(n9741) );
  NAND2_X1 U10110 ( .A1(n13412), .A2(n9769), .ZN(n9770) );
  NOR2_X1 U10111 ( .A1(n10075), .A2(n10074), .ZN(n10076) );
  INV_X1 U10112 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8586) );
  INV_X1 U10113 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9351) );
  INV_X1 U10114 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n9337) );
  INV_X1 U10115 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9336) );
  INV_X1 U10116 ( .A(n10112), .ZN(n9110) );
  INV_X1 U10117 ( .A(n14433), .ZN(n9048) );
  OR2_X1 U10118 ( .A1(n8753), .A2(n8752), .ZN(n8774) );
  INV_X1 U10119 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8492) );
  OR2_X1 U10120 ( .A1(n10845), .A2(n15094), .ZN(n10847) );
  INV_X1 U10121 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11701) );
  INV_X1 U10122 ( .A(n13025), .ZN(n12207) );
  NOR2_X1 U10123 ( .A1(n8510), .A2(n10166), .ZN(n8512) );
  AND2_X1 U10124 ( .A1(n13378), .A2(n13379), .ZN(n13333) );
  NAND2_X1 U10125 ( .A1(n9356), .A2(n9355), .ZN(n9764) );
  INV_X1 U10126 ( .A(n13999), .ZN(n9813) );
  OR2_X1 U10127 ( .A1(n9310), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9311) );
  AND2_X1 U10128 ( .A1(n9280), .A2(n9279), .ZN(n9501) );
  INV_X1 U10129 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U10130 ( .A1(n14271), .A2(n14272), .ZN(n14273) );
  NAND2_X1 U10131 ( .A1(n8601), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8934) );
  OR3_X1 U10132 ( .A1(n8989), .A2(n8987), .A3(n8988), .ZN(n8990) );
  INV_X1 U10133 ( .A(n10119), .ZN(n10120) );
  INV_X1 U10134 ( .A(n8897), .ZN(n8600) );
  OR2_X1 U10135 ( .A1(n8828), .A2(n10931), .ZN(n8840) );
  OAI22_X1 U10136 ( .A1(n14318), .A2(n14794), .B1(n14546), .B2(n10033), .ZN(
        n9118) );
  OR2_X1 U10137 ( .A1(n8787), .A2(n8786), .ZN(n8816) );
  INV_X1 U10138 ( .A(n8816), .ZN(n8597) );
  INV_X1 U10139 ( .A(n10109), .ZN(n14587) );
  AND2_X1 U10140 ( .A1(n10974), .A2(n8503), .ZN(n10896) );
  INV_X1 U10141 ( .A(n15164), .ZN(n15015) );
  INV_X1 U10142 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n12197) );
  AND2_X1 U10143 ( .A1(n12530), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12604) );
  NOR2_X1 U10144 ( .A1(n12831), .A2(n12721), .ZN(n12851) );
  INV_X1 U10145 ( .A(n15484), .ZN(n15582) );
  NOR2_X1 U10146 ( .A1(n10715), .A2(n12994), .ZN(n15437) );
  AND2_X1 U10147 ( .A1(n15638), .A2(n15637), .ZN(n15639) );
  INV_X1 U10148 ( .A(n12733), .ZN(n10719) );
  AND2_X1 U10149 ( .A1(n10716), .A2(n10416), .ZN(n10423) );
  INV_X1 U10150 ( .A(n8848), .ZN(n8555) );
  OR2_X1 U10151 ( .A1(n10631), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n11184) );
  INV_X1 U10152 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9127) );
  NOR2_X1 U10153 ( .A1(n9165), .A2(n9164), .ZN(n9147) );
  AND2_X1 U10154 ( .A1(n9212), .A2(n9211), .ZN(n9152) );
  INV_X1 U10155 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9347) );
  INV_X1 U10156 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n13712) );
  INV_X1 U10157 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U10158 ( .A1(n12354), .A2(n13515), .ZN(n12355) );
  OR2_X1 U10159 ( .A1(n10602), .A2(n10461), .ZN(n13470) );
  OR2_X1 U10160 ( .A1(n9764), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n13903) );
  NOR2_X1 U10161 ( .A1(n8474), .A2(n13920), .ZN(n13921) );
  INV_X1 U10162 ( .A(n13281), .ZN(n14011) );
  AND2_X1 U10163 ( .A1(n13148), .A2(n13149), .ZN(n13272) );
  AND2_X1 U10164 ( .A1(n10775), .A2(n13881), .ZN(n16045) );
  OR2_X1 U10165 ( .A1(n9443), .A2(n13632), .ZN(n9344) );
  NAND2_X1 U10166 ( .A1(n9312), .A2(n9311), .ZN(n9374) );
  NAND2_X1 U10167 ( .A1(n9690), .A2(n9303), .ZN(n9702) );
  AND2_X1 U10168 ( .A1(n9295), .A2(n9294), .ZN(n9628) );
  AND2_X1 U10169 ( .A1(n9271), .A2(n9270), .ZN(n9441) );
  AND2_X1 U10170 ( .A1(n9263), .A2(n9262), .ZN(n9401) );
  NAND2_X1 U10171 ( .A1(n8598), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8868) );
  OR2_X1 U10172 ( .A1(n8883), .A2(n14434), .ZN(n8897) );
  OR2_X1 U10173 ( .A1(n14621), .A2(n9058), .ZN(n8971) );
  INV_X1 U10174 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10931) );
  INV_X1 U10175 ( .A(n14633), .ZN(n14598) );
  INV_X1 U10176 ( .A(n14472), .ZN(n14327) );
  OR2_X1 U10177 ( .A1(n9243), .A2(n8503), .ZN(n10838) );
  NAND2_X1 U10178 ( .A1(n10025), .A2(n10044), .ZN(n10027) );
  AND2_X1 U10179 ( .A1(n9042), .A2(n9041), .ZN(n12405) );
  AND2_X1 U10180 ( .A1(n9056), .A2(n9055), .ZN(n14719) );
  INV_X1 U10181 ( .A(n15438), .ZN(n15381) );
  OR2_X1 U10182 ( .A1(n10857), .A2(n10856), .ZN(n10858) );
  NAND2_X1 U10183 ( .A1(n11907), .A2(n11906), .ZN(n12020) );
  INV_X1 U10184 ( .A(n12889), .ZN(n12888) );
  INV_X1 U10185 ( .A(n15216), .ZN(n15192) );
  OR2_X1 U10186 ( .A1(n10418), .A2(n10419), .ZN(n15213) );
  AND2_X1 U10187 ( .A1(n12851), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n12861) );
  INV_X1 U10188 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n12711) );
  INV_X1 U10189 ( .A(n12279), .ZN(n12652) );
  NOR2_X1 U10190 ( .A1(n16005), .A2(n12731), .ZN(n10410) );
  INV_X1 U10191 ( .A(n15380), .ZN(n15434) );
  INV_X1 U10192 ( .A(n13031), .ZN(n12660) );
  INV_X1 U10193 ( .A(n12770), .ZN(n16095) );
  NOR2_X1 U10194 ( .A1(n10417), .A2(n10423), .ZN(n13061) );
  OAI21_X1 U10195 ( .B1(n10209), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10144) );
  AND2_X1 U10196 ( .A1(n9858), .A2(n9857), .ZN(n10132) );
  AND2_X1 U10197 ( .A1(n9740), .A2(n9739), .ZN(n13978) );
  INV_X1 U10198 ( .A(n13889), .ZN(n13874) );
  AND2_X1 U10199 ( .A1(n10461), .A2(n13229), .ZN(n14108) );
  INV_X1 U10200 ( .A(n16126), .ZN(n14065) );
  INV_X1 U10201 ( .A(n14118), .ZN(n14099) );
  AND2_X1 U10202 ( .A1(n9867), .A2(n9866), .ZN(n11058) );
  INV_X1 U10203 ( .A(n14246), .ZN(n9862) );
  INV_X1 U10204 ( .A(n16222), .ZN(n16054) );
  INV_X1 U10205 ( .A(n14182), .ZN(n16226) );
  INV_X1 U10206 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9457) );
  NOR3_X1 U10207 ( .A1(n14965), .A2(n12688), .A3(n14967), .ZN(n10131) );
  INV_X1 U10208 ( .A(n14403), .ZN(n14459) );
  AND3_X1 U10209 ( .A1(n9117), .A2(n9116), .A3(n9115), .ZN(n10033) );
  INV_X1 U10210 ( .A(n8649), .ZN(n9058) );
  INV_X1 U10211 ( .A(n9882), .ZN(n11395) );
  AND2_X1 U10212 ( .A1(n10933), .A2(n10932), .ZN(n15892) );
  INV_X1 U10213 ( .A(n14697), .ZN(n16080) );
  INV_X1 U10214 ( .A(n14794), .ZN(n14647) );
  INV_X1 U10215 ( .A(n14751), .ZN(n16088) );
  INV_X1 U10216 ( .A(n16062), .ZN(n14753) );
  INV_X1 U10217 ( .A(n16094), .ZN(n14805) );
  INV_X1 U10218 ( .A(n14897), .ZN(n11947) );
  NOR2_X1 U10219 ( .A1(n15812), .A2(n9095), .ZN(n9125) );
  INV_X1 U10220 ( .A(n16138), .ZN(n16204) );
  INV_X1 U10221 ( .A(n14876), .ZN(n14884) );
  INV_X1 U10222 ( .A(n16201), .ZN(n16134) );
  XNOR2_X1 U10223 ( .A(n9081), .B(n9080), .ZN(n10895) );
  INV_X1 U10224 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8501) );
  AND2_X1 U10225 ( .A1(n8782), .A2(n8770), .ZN(n10924) );
  INV_X1 U10226 ( .A(n12749), .ZN(n15181) );
  INV_X1 U10227 ( .A(n12972), .ZN(n12977) );
  OR2_X1 U10228 ( .A1(n15917), .A2(n10715), .ZN(n15337) );
  INV_X1 U10229 ( .A(n12275), .ZN(n15927) );
  INV_X1 U10230 ( .A(n16014), .ZN(n15617) );
  INV_X1 U10231 ( .A(n15404), .ZN(n15535) );
  AND2_X1 U10232 ( .A1(n10716), .A2(n10715), .ZN(n15500) );
  INV_X1 U10233 ( .A(n15577), .ZN(n15620) );
  INV_X1 U10234 ( .A(n16002), .ZN(n15490) );
  NAND2_X1 U10235 ( .A1(n15387), .A2(n15615), .ZN(n15611) );
  INV_X1 U10236 ( .A(n15361), .ZN(n15627) );
  NAND2_X1 U10237 ( .A1(n12992), .A2(n10707), .ZN(n16116) );
  INV_X1 U10238 ( .A(n16176), .ZN(n15732) );
  NAND2_X1 U10239 ( .A1(n16002), .A2(n16116), .ZN(n16176) );
  INV_X1 U10240 ( .A(n11044), .ZN(n10688) );
  OR2_X1 U10241 ( .A1(n10229), .A2(n12685), .ZN(n10390) );
  NAND2_X1 U10242 ( .A1(n10145), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10231) );
  AND2_X1 U10243 ( .A1(n10683), .A2(n10820), .ZN(n12193) );
  INV_X1 U10244 ( .A(n10132), .ZN(n10446) );
  INV_X1 U10245 ( .A(n13495), .ZN(n13440) );
  INV_X1 U10246 ( .A(n13411), .ZN(n13507) );
  INV_X1 U10247 ( .A(n14028), .ZN(n14058) );
  NAND2_X1 U10248 ( .A1(n10437), .A2(n10436), .ZN(n13895) );
  INV_X1 U10249 ( .A(n13897), .ZN(n13877) );
  NAND2_X1 U10250 ( .A1(n16131), .A2(n16123), .ZN(n14118) );
  NAND2_X1 U10251 ( .A1(n9861), .A2(n9879), .ZN(n9880) );
  NAND2_X1 U10252 ( .A1(n16228), .A2(n16054), .ZN(n14192) );
  NAND2_X1 U10253 ( .A1(n9861), .A2(n9862), .ZN(n9863) );
  INV_X1 U10254 ( .A(n16232), .ZN(n16229) );
  AND2_X2 U10255 ( .A1(n9859), .A2(n10466), .ZN(n16232) );
  INV_X1 U10256 ( .A(SI_14_), .ZN(n13624) );
  INV_X1 U10257 ( .A(n10628), .ZN(n10529) );
  CLKBUF_X1 U10258 ( .A(n12396), .Z(n13319) );
  NAND2_X1 U10259 ( .A1(n10835), .A2(n10834), .ZN(n14449) );
  INV_X1 U10260 ( .A(n14423), .ZN(n14462) );
  NAND2_X1 U10261 ( .A1(n9022), .A2(n9021), .ZN(n14465) );
  INV_X1 U10262 ( .A(n14361), .ZN(n14467) );
  INV_X1 U10263 ( .A(n12335), .ZN(n14475) );
  OR2_X1 U10264 ( .A1(n10933), .A2(P2_U3088), .ZN(n15904) );
  INV_X1 U10265 ( .A(n15898), .ZN(n15859) );
  XNOR2_X1 U10266 ( .A(n9108), .B(n9110), .ZN(n13092) );
  INV_X1 U10267 ( .A(n14805), .ZN(n16082) );
  OR2_X1 U10268 ( .A1(n16094), .A2(n11546), .ZN(n14806) );
  AND2_X1 U10269 ( .A1(n11516), .A2(n14697), .ZN(n16094) );
  OR2_X1 U10270 ( .A1(n16208), .A2(n9254), .ZN(n9255) );
  INV_X1 U10271 ( .A(n14601), .ZN(n14912) );
  NAND2_X1 U10272 ( .A1(n14948), .A2(n16134), .ZN(n14951) );
  OR2_X1 U10273 ( .A1(n15818), .A2(n15815), .ZN(n15816) );
  INV_X1 U10274 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11425) );
  INV_X1 U10275 ( .A(n12793), .ZN(n16172) );
  INV_X1 U10276 ( .A(n12805), .ZN(n12594) );
  OR2_X1 U10277 ( .A1(n10419), .A2(n10408), .ZN(n15205) );
  OR2_X1 U10278 ( .A1(n15917), .A2(n15905), .ZN(n12275) );
  OR2_X1 U10279 ( .A1(n15917), .A2(n10291), .ZN(n15338) );
  OR2_X1 U10280 ( .A1(n16022), .A2(n12996), .ZN(n15598) );
  INV_X2 U10281 ( .A(n10228), .ZN(n15811) );
  INV_X1 U10282 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11925) );
  INV_X1 U10283 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10685) );
  AND2_X1 U10284 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10894), .ZN(P2_U3947) );
  NOR2_X2 U10285 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8583) );
  NOR2_X2 U10286 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8584) );
  NAND3_X1 U10287 ( .A1(n8583), .A2(n8584), .A3(n8495), .ZN(n8484) );
  NOR2_X1 U10288 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8488) );
  NOR2_X1 U10289 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n8487) );
  NAND2_X1 U10290 ( .A1(n8489), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8864) );
  INV_X1 U10291 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U10292 ( .A1(n8864), .A2(n8490), .ZN(n8491) );
  NAND2_X1 U10293 ( .A1(n8880), .A2(n8492), .ZN(n8493) );
  NAND2_X1 U10294 ( .A1(n8505), .A2(n8504), .ZN(n8494) );
  NAND2_X1 U10295 ( .A1(n8494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8496) );
  INV_X1 U10296 ( .A(n8503), .ZN(n12564) );
  NAND2_X1 U10297 ( .A1(n8500), .A2(n8499), .ZN(n9067) );
  NAND2_X1 U10298 ( .A1(n9067), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8502) );
  OR2_X1 U10299 ( .A1(n10976), .A2(n10974), .ZN(n8507) );
  NOR2_X1 U10300 ( .A1(n10896), .A2(n9093), .ZN(n8506) );
  NAND2_X1 U10301 ( .A1(n8507), .A2(n8506), .ZN(n14876) );
  INV_X1 U10302 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10690) );
  NAND2_X1 U10303 ( .A1(n8520), .A2(SI_2_), .ZN(n8514) );
  INV_X1 U10304 ( .A(SI_1_), .ZN(n10173) );
  INV_X1 U10305 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10381) );
  INV_X1 U10306 ( .A(SI_0_), .ZN(n10380) );
  INV_X1 U10307 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9257) );
  NAND2_X1 U10308 ( .A1(n8515), .A2(n9257), .ZN(n8509) );
  INV_X1 U10309 ( .A(SI_2_), .ZN(n10166) );
  NAND3_X1 U10310 ( .A1(n8511), .A2(n10166), .A3(n8517), .ZN(n8513) );
  MUX2_X1 U10311 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n10689), .Z(n8638) );
  NAND2_X1 U10312 ( .A1(n8517), .A2(n8516), .ZN(n8619) );
  INV_X1 U10313 ( .A(n8619), .ZN(n8519) );
  INV_X1 U10314 ( .A(n8522), .ZN(n8655) );
  MUX2_X1 U10315 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8515), .Z(n8525) );
  NAND2_X1 U10316 ( .A1(n8525), .A2(SI_4_), .ZN(n8527) );
  OAI21_X1 U10317 ( .B1(n8525), .B2(SI_4_), .A(n8527), .ZN(n8526) );
  INV_X1 U10318 ( .A(n8526), .ZN(n8670) );
  MUX2_X1 U10319 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10689), .Z(n8528) );
  NAND2_X1 U10320 ( .A1(n8528), .A2(SI_5_), .ZN(n8530) );
  OAI21_X1 U10321 ( .B1(n8528), .B2(SI_5_), .A(n8530), .ZN(n8529) );
  INV_X1 U10322 ( .A(n8529), .ZN(n8690) );
  INV_X1 U10323 ( .A(n8711), .ZN(n8531) );
  MUX2_X1 U10324 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10689), .Z(n8533) );
  NAND2_X1 U10325 ( .A1(n8533), .A2(SI_7_), .ZN(n8535) );
  OAI21_X1 U10326 ( .B1(SI_7_), .B2(n8533), .A(n8535), .ZN(n8716) );
  INV_X1 U10327 ( .A(n8716), .ZN(n8534) );
  MUX2_X1 U10328 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10689), .Z(n8537) );
  NAND2_X1 U10329 ( .A1(n8537), .A2(SI_8_), .ZN(n8539) );
  OAI21_X1 U10330 ( .B1(SI_8_), .B2(n8537), .A(n8539), .ZN(n8729) );
  INV_X1 U10331 ( .A(n8729), .ZN(n8538) );
  MUX2_X1 U10332 ( .A(n10359), .B(n10360), .S(n10178), .Z(n8745) );
  MUX2_X1 U10333 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10689), .Z(n8541) );
  NAND2_X1 U10334 ( .A1(n8541), .A2(SI_10_), .ZN(n8543) );
  OAI21_X1 U10335 ( .B1(SI_10_), .B2(n8541), .A(n8543), .ZN(n8542) );
  INV_X1 U10336 ( .A(n8542), .ZN(n8761) );
  MUX2_X1 U10337 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n10178), .Z(n8544) );
  XNOR2_X1 U10338 ( .A(n8544), .B(SI_11_), .ZN(n8780) );
  INV_X1 U10339 ( .A(n8544), .ZN(n8545) );
  NAND2_X1 U10340 ( .A1(n8545), .A2(n13666), .ZN(n8546) );
  MUX2_X1 U10341 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n10689), .Z(n8547) );
  XNOR2_X1 U10342 ( .A(n8547), .B(n10222), .ZN(n8795) );
  INV_X1 U10343 ( .A(n8547), .ZN(n8548) );
  MUX2_X1 U10344 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10689), .Z(n8549) );
  OAI21_X1 U10345 ( .B1(n8549), .B2(SI_13_), .A(n8550), .ZN(n8809) );
  MUX2_X1 U10346 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n10178), .Z(n8551) );
  XNOR2_X1 U10347 ( .A(n8551), .B(SI_14_), .ZN(n8822) );
  INV_X1 U10348 ( .A(n8551), .ZN(n8552) );
  NAND2_X1 U10349 ( .A1(n8552), .A2(n13624), .ZN(n8553) );
  MUX2_X1 U10350 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n10689), .Z(n8554) );
  MUX2_X1 U10351 ( .A(n11435), .B(n11425), .S(n10178), .Z(n8848) );
  MUX2_X1 U10352 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n10689), .Z(n8557) );
  MUX2_X1 U10353 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10178), .Z(n8875) );
  MUX2_X1 U10354 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10178), .Z(n8559) );
  XNOR2_X1 U10355 ( .A(n8559), .B(SI_19_), .ZN(n8892) );
  INV_X1 U10356 ( .A(n8559), .ZN(n8560) );
  INV_X1 U10357 ( .A(SI_19_), .ZN(n10649) );
  MUX2_X1 U10358 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n10178), .Z(n8904) );
  NOR2_X1 U10359 ( .A1(n8904), .A2(SI_20_), .ZN(n8562) );
  NAND2_X1 U10360 ( .A1(n8904), .A2(SI_20_), .ZN(n8561) );
  MUX2_X1 U10361 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10689), .Z(n8564) );
  XNOR2_X1 U10362 ( .A(n8564), .B(SI_21_), .ZN(n8916) );
  INV_X1 U10363 ( .A(n8916), .ZN(n8563) );
  MUX2_X1 U10364 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10178), .Z(n8927) );
  MUX2_X1 U10365 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10178), .Z(n8946) );
  INV_X1 U10366 ( .A(n8946), .ZN(n8565) );
  INV_X1 U10367 ( .A(SI_23_), .ZN(n13650) );
  AOI22_X1 U10368 ( .A1(n13652), .A2(n8928), .B1(n8565), .B2(n13650), .ZN(
        n8566) );
  OAI21_X1 U10369 ( .B1(n8928), .B2(n13652), .A(n13650), .ZN(n8568) );
  AND2_X1 U10370 ( .A1(SI_22_), .A2(SI_23_), .ZN(n8567) );
  AOI22_X1 U10371 ( .A1(n8568), .A2(n8946), .B1(n8927), .B2(n8567), .ZN(n8569)
         );
  MUX2_X1 U10372 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10178), .Z(n8572) );
  XNOR2_X1 U10373 ( .A(n8572), .B(SI_24_), .ZN(n8960) );
  INV_X1 U10374 ( .A(n8960), .ZN(n8571) );
  NAND2_X1 U10375 ( .A1(n8961), .A2(n8571), .ZN(n8574) );
  NAND2_X1 U10376 ( .A1(n8572), .A2(SI_24_), .ZN(n8573) );
  INV_X1 U10377 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15772) );
  INV_X1 U10378 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14969) );
  MUX2_X1 U10379 ( .A(n15772), .B(n14969), .S(n10689), .Z(n8575) );
  NAND2_X1 U10380 ( .A1(n8575), .A2(n13643), .ZN(n8578) );
  INV_X1 U10381 ( .A(n8575), .ZN(n8576) );
  NAND2_X1 U10382 ( .A1(n8576), .A2(SI_25_), .ZN(n8577) );
  NAND2_X1 U10383 ( .A1(n8578), .A2(n8577), .ZN(n8974) );
  MUX2_X1 U10384 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10178), .Z(n8579) );
  NAND2_X1 U10385 ( .A1(n8579), .A2(SI_26_), .ZN(n8580) );
  INV_X1 U10386 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12941) );
  INV_X1 U10387 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13323) );
  MUX2_X1 U10388 ( .A(n12941), .B(n13323), .S(n10178), .Z(n9001) );
  XNOR2_X1 U10389 ( .A(n9001), .B(SI_27_), .ZN(n8999) );
  INV_X1 U10390 ( .A(n8999), .ZN(n8581) );
  NOR2_X1 U10391 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8582) );
  NAND2_X1 U10392 ( .A1(n12940), .A2(n10044), .ZN(n8590) );
  NAND2_X1 U10393 ( .A1(n9104), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U10394 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8684) );
  INV_X1 U10395 ( .A(n8684), .ZN(n8591) );
  NAND2_X1 U10396 ( .A1(n8591), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8705) );
  INV_X1 U10397 ( .A(n8705), .ZN(n8592) );
  NAND2_X1 U10398 ( .A1(n8592), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8723) );
  INV_X1 U10399 ( .A(n8723), .ZN(n8593) );
  NAND2_X1 U10400 ( .A1(n8593), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8736) );
  INV_X1 U10401 ( .A(n8736), .ZN(n8594) );
  NAND2_X1 U10402 ( .A1(n8594), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8753) );
  INV_X1 U10403 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8752) );
  INV_X1 U10404 ( .A(n8774), .ZN(n8595) );
  NAND2_X1 U10405 ( .A1(n8595), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8787) );
  INV_X1 U10406 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8786) );
  AND2_X1 U10407 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .ZN(n8596) );
  NAND2_X1 U10408 ( .A1(n8597), .A2(n8596), .ZN(n8828) );
  INV_X1 U10409 ( .A(n8868), .ZN(n8599) );
  NAND2_X1 U10410 ( .A1(n8599), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8883) );
  INV_X1 U10411 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n14434) );
  INV_X1 U10412 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n14414) );
  INV_X1 U10413 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8933) );
  INV_X1 U10414 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8987) );
  INV_X1 U10415 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8988) );
  INV_X1 U10416 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n14317) );
  NOR2_X1 U10417 ( .A1(n8990), .A2(n14317), .ZN(n9013) );
  INV_X1 U10418 ( .A(n9013), .ZN(n9015) );
  NAND2_X1 U10419 ( .A1(n8990), .A2(n14317), .ZN(n8604) );
  NAND2_X1 U10420 ( .A1(n9015), .A2(n8604), .ZN(n14567) );
  INV_X1 U10421 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n14566) );
  NAND2_X1 U10422 ( .A1(n8650), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8613) );
  AND2_X2 U10423 ( .A1(n12718), .A2(n8609), .ZN(n8665) );
  NAND2_X1 U10424 ( .A1(n8665), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8612) );
  OAI211_X1 U10425 ( .C1(n14566), .C2(n10032), .A(n8613), .B(n8612), .ZN(n8614) );
  INV_X1 U10426 ( .A(n8614), .ZN(n8615) );
  NAND2_X1 U10427 ( .A1(n8665), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U10428 ( .A1(n8650), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U10429 ( .A1(n8619), .A2(n8510), .ZN(n8620) );
  NAND2_X1 U10430 ( .A1(n8621), .A2(n8620), .ZN(n10692) );
  INV_X2 U10431 ( .A(n8629), .ZN(n8674) );
  NAND2_X1 U10432 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8622) );
  XNOR2_X1 U10433 ( .A(n8622), .B(P2_IR_REG_1__SCAN_IN), .ZN(n14488) );
  NAND2_X1 U10434 ( .A1(n8674), .A2(n14488), .ZN(n8623) );
  NAND2_X1 U10435 ( .A1(n8665), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U10436 ( .A1(n8650), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U10437 ( .A1(n8649), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U10438 ( .A1(n8885), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U10439 ( .A1(n10689), .A2(SI_0_), .ZN(n9391) );
  XNOR2_X1 U10440 ( .A(n9391), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14976) );
  MUX2_X1 U10441 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14976), .S(n8629), .Z(n11399)
         );
  AND2_X1 U10442 ( .A1(n9882), .A2(n11399), .ZN(n11391) );
  NAND2_X1 U10443 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  NAND2_X1 U10444 ( .A1(n8665), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U10445 ( .A1(n8650), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U10446 ( .A1(n8649), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U10447 ( .A1(n8885), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8633) );
  INV_X1 U10448 ( .A(n8637), .ZN(n8640) );
  INV_X1 U10449 ( .A(n8638), .ZN(n8639) );
  NAND2_X1 U10450 ( .A1(n8640), .A2(n8639), .ZN(n8641) );
  NAND2_X1 U10451 ( .A1(n8642), .A2(n8641), .ZN(n10701) );
  OR2_X1 U10452 ( .A1(n8643), .A2(n8810), .ZN(n8644) );
  XNOR2_X1 U10453 ( .A(n8644), .B(P2_IR_REG_2__SCAN_IN), .ZN(n11271) );
  NAND2_X1 U10454 ( .A1(n8674), .A2(n11271), .ZN(n8645) );
  INV_X1 U10455 ( .A(n11407), .ZN(n11404) );
  NAND2_X1 U10456 ( .A1(n11405), .A2(n11404), .ZN(n8648) );
  INV_X1 U10457 ( .A(n14483), .ZN(n11394) );
  INV_X1 U10458 ( .A(n11724), .ZN(n11413) );
  NAND2_X1 U10459 ( .A1(n11394), .A2(n11413), .ZN(n8647) );
  NAND2_X1 U10460 ( .A1(n8648), .A2(n8647), .ZN(n10993) );
  INV_X1 U10461 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n16060) );
  NAND2_X1 U10462 ( .A1(n8649), .A2(n16060), .ZN(n8654) );
  NAND2_X1 U10463 ( .A1(n8650), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U10464 ( .A1(n8665), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U10465 ( .A1(n8885), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U10466 ( .A1(n8657), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8658) );
  XNOR2_X1 U10467 ( .A(n8658), .B(P2_IR_REG_3__SCAN_IN), .ZN(n14504) );
  NAND2_X1 U10468 ( .A1(n8674), .A2(n14504), .ZN(n8659) );
  NAND2_X1 U10469 ( .A1(n10993), .A2(n7605), .ZN(n8662) );
  INV_X1 U10470 ( .A(n14482), .ZN(n9029) );
  NAND2_X1 U10471 ( .A1(n9029), .A2(n7910), .ZN(n8661) );
  NAND2_X1 U10472 ( .A1(n8650), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8669) );
  INV_X1 U10473 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U10474 ( .A1(n16060), .A2(n8663), .ZN(n8664) );
  AND2_X1 U10475 ( .A1(n8664), .A2(n8684), .ZN(n16081) );
  NAND2_X1 U10476 ( .A1(n8649), .A2(n16081), .ZN(n8668) );
  NAND2_X1 U10477 ( .A1(n8665), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U10478 ( .A1(n8885), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U10479 ( .A1(n9104), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U10480 ( .A1(n8675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8676) );
  MUX2_X1 U10481 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8676), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8678) );
  INV_X1 U10482 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U10483 ( .A1(n7615), .A2(n8677), .ZN(n8695) );
  NAND2_X1 U10484 ( .A1(n8678), .A2(n8695), .ZN(n14521) );
  INV_X1 U10485 ( .A(n14521), .ZN(n14515) );
  NAND2_X1 U10486 ( .A1(n8674), .A2(n14515), .ZN(n8679) );
  INV_X1 U10487 ( .A(n11597), .ZN(n8681) );
  INV_X1 U10488 ( .A(n14481), .ZN(n9031) );
  INV_X1 U10489 ( .A(n11603), .ZN(n16084) );
  NAND2_X1 U10490 ( .A1(n9031), .A2(n16084), .ZN(n8682) );
  NAND2_X1 U10491 ( .A1(n8650), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8689) );
  INV_X1 U10492 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U10493 ( .A1(n8684), .A2(n8683), .ZN(n8685) );
  AND2_X1 U10494 ( .A1(n8705), .A2(n8685), .ZN(n11839) );
  NAND2_X1 U10495 ( .A1(n8649), .A2(n11839), .ZN(n8688) );
  NAND2_X1 U10496 ( .A1(n8665), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U10497 ( .A1(n8885), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8686) );
  NAND4_X1 U10498 ( .A1(n8689), .A2(n8688), .A3(n8687), .A4(n8686), .ZN(n14480) );
  OR2_X1 U10499 ( .A1(n8691), .A2(n8690), .ZN(n8692) );
  NAND2_X1 U10500 ( .A1(n8693), .A2(n8692), .ZN(n11190) );
  NOR2_X1 U10501 ( .A1(n11190), .A2(n10024), .ZN(n8701) );
  NAND2_X1 U10502 ( .A1(n8695), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8694) );
  MUX2_X1 U10503 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8694), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8698) );
  INV_X1 U10504 ( .A(n8695), .ZN(n8697) );
  INV_X1 U10505 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U10506 ( .A1(n8697), .A2(n8696), .ZN(n8718) );
  NAND2_X1 U10507 ( .A1(n8698), .A2(n8718), .ZN(n10911) );
  OAI22_X1 U10508 ( .A1(n8699), .A2(n10183), .B1(n8629), .B2(n10911), .ZN(
        n8700) );
  OR2_X2 U10509 ( .A1(n8701), .A2(n8700), .ZN(n11840) );
  NOR2_X1 U10510 ( .A1(n14480), .A2(n11840), .ZN(n8702) );
  NAND2_X1 U10511 ( .A1(n14480), .A2(n11840), .ZN(n8703) );
  NAND2_X1 U10512 ( .A1(n8650), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8710) );
  INV_X1 U10513 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U10514 ( .A1(n8705), .A2(n8704), .ZN(n8706) );
  AND2_X1 U10515 ( .A1(n8723), .A2(n8706), .ZN(n11506) );
  NAND2_X1 U10516 ( .A1(n8649), .A2(n11506), .ZN(n8709) );
  NAND2_X1 U10517 ( .A1(n8665), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U10518 ( .A1(n8885), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8707) );
  NAND4_X1 U10519 ( .A1(n8710), .A2(n8709), .A3(n8708), .A4(n8707), .ZN(n14479) );
  NAND2_X1 U10520 ( .A1(n11315), .A2(n10044), .ZN(n8715) );
  NAND2_X1 U10521 ( .A1(n8718), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8713) );
  XNOR2_X1 U10522 ( .A(n8713), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14539) );
  AOI22_X1 U10523 ( .A1(n9104), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8674), .B2(
        n14539), .ZN(n8714) );
  XNOR2_X1 U10524 ( .A(n8717), .B(n8716), .ZN(n11442) );
  NAND2_X1 U10525 ( .A1(n11442), .A2(n10044), .ZN(n8721) );
  NAND2_X1 U10526 ( .A1(n8731), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8719) );
  XNOR2_X1 U10527 ( .A(n8719), .B(P2_IR_REG_7__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U10528 ( .A1(n9104), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8674), .B2(
        n11166), .ZN(n8720) );
  INV_X1 U10529 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U10530 ( .A1(n8723), .A2(n8722), .ZN(n8724) );
  AND2_X1 U10531 ( .A1(n8736), .A2(n8724), .ZN(n11685) );
  NAND2_X1 U10532 ( .A1(n8649), .A2(n11685), .ZN(n8728) );
  NAND2_X1 U10533 ( .A1(n8650), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8727) );
  NAND2_X1 U10534 ( .A1(n8665), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U10535 ( .A1(n8885), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U10536 ( .A(n11668), .B(n14478), .ZN(n10096) );
  INV_X1 U10537 ( .A(n10096), .ZN(n11661) );
  XNOR2_X1 U10538 ( .A(n8730), .B(n8729), .ZN(n11694) );
  NAND2_X1 U10539 ( .A1(n11694), .A2(n10044), .ZN(n8734) );
  NAND2_X1 U10540 ( .A1(n8749), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8732) );
  XNOR2_X1 U10541 ( .A(n8732), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U10542 ( .A1(n9104), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8674), .B2(
        n10920), .ZN(n8733) );
  NAND2_X1 U10543 ( .A1(n8650), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8741) );
  INV_X1 U10544 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U10545 ( .A1(n8736), .A2(n8735), .ZN(n8737) );
  AND2_X1 U10546 ( .A1(n8753), .A2(n8737), .ZN(n11884) );
  NAND2_X1 U10547 ( .A1(n8649), .A2(n11884), .ZN(n8740) );
  NAND2_X1 U10548 ( .A1(n8665), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U10549 ( .A1(n8885), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U10550 ( .A1(n16133), .A2(n11875), .ZN(n11936) );
  OR2_X1 U10551 ( .A1(n16133), .A2(n11875), .ZN(n8742) );
  INV_X1 U10552 ( .A(n11895), .ZN(n8743) );
  OR2_X1 U10553 ( .A1(n11901), .A2(n11875), .ZN(n8744) );
  NAND2_X1 U10554 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  NAND2_X1 U10555 ( .A1(n8748), .A2(n8747), .ZN(n11805) );
  OAI21_X1 U10556 ( .B1(n8749), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8766) );
  XNOR2_X1 U10557 ( .A(n8766), .B(P2_IR_REG_9__SCAN_IN), .ZN(n15891) );
  AOI22_X1 U10558 ( .A1(n9104), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8674), .B2(
        n15891), .ZN(n8750) );
  NAND2_X1 U10559 ( .A1(n8650), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U10560 ( .A1(n8753), .A2(n8752), .ZN(n8754) );
  AND2_X1 U10561 ( .A1(n8774), .A2(n8754), .ZN(n12093) );
  NAND2_X1 U10562 ( .A1(n8649), .A2(n12093), .ZN(n8757) );
  NAND2_X1 U10563 ( .A1(n8665), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U10564 ( .A1(n8885), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U10565 ( .A1(n11944), .A2(n14476), .ZN(n8759) );
  OR2_X1 U10566 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  AND2_X1 U10567 ( .A1(n8764), .A2(n8763), .ZN(n12016) );
  NAND2_X1 U10568 ( .A1(n12016), .A2(n10044), .ZN(n8772) );
  INV_X1 U10569 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U10570 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  NAND2_X1 U10571 ( .A1(n8767), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8769) );
  INV_X1 U10572 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U10573 ( .A1(n8769), .A2(n8768), .ZN(n8782) );
  OR2_X1 U10574 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  AOI22_X1 U10575 ( .A1(n9104), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8674), 
        .B2(n10924), .ZN(n8771) );
  INV_X1 U10576 ( .A(n16186), .ZN(n12149) );
  NAND2_X1 U10577 ( .A1(n8650), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8779) );
  INV_X1 U10578 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U10579 ( .A1(n8774), .A2(n8773), .ZN(n8775) );
  AND2_X1 U10580 ( .A1(n8787), .A2(n8775), .ZN(n12144) );
  NAND2_X1 U10581 ( .A1(n8649), .A2(n12144), .ZN(n8778) );
  NAND2_X1 U10582 ( .A1(n8665), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U10583 ( .A1(n8885), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8776) );
  XNOR2_X1 U10584 ( .A(n12149), .B(n14475), .ZN(n12140) );
  XNOR2_X1 U10585 ( .A(n8781), .B(n8780), .ZN(n12074) );
  NAND2_X1 U10586 ( .A1(n12074), .A2(n10044), .ZN(n8785) );
  NAND2_X1 U10587 ( .A1(n8782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8783) );
  XNOR2_X1 U10588 ( .A(n8783), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U10589 ( .A1(n9104), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8674), 
        .B2(n10970), .ZN(n8784) );
  NAND2_X1 U10590 ( .A1(n8650), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U10591 ( .A1(n8787), .A2(n8786), .ZN(n8788) );
  AND2_X1 U10592 ( .A1(n8816), .A2(n8788), .ZN(n12337) );
  NAND2_X1 U10593 ( .A1(n8649), .A2(n12337), .ZN(n8791) );
  NAND2_X1 U10594 ( .A1(n8665), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U10595 ( .A1(n8885), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U10596 ( .A1(n12422), .A2(n12499), .ZN(n9040) );
  OR2_X1 U10597 ( .A1(n12422), .A2(n12499), .ZN(n8793) );
  OR2_X1 U10598 ( .A1(n12425), .A2(n12499), .ZN(n8794) );
  XNOR2_X1 U10599 ( .A(n8796), .B(n8795), .ZN(n12187) );
  NAND2_X1 U10600 ( .A1(n12187), .A2(n10044), .ZN(n8801) );
  NOR2_X1 U10601 ( .A1(n8485), .A2(n8810), .ZN(n8797) );
  MUX2_X1 U10602 ( .A(n8810), .B(n8797), .S(P2_IR_REG_12__SCAN_IN), .Z(n8799)
         );
  OR2_X1 U10603 ( .A1(n8799), .A2(n8798), .ZN(n10926) );
  INV_X1 U10604 ( .A(n10926), .ZN(n15882) );
  AOI22_X1 U10605 ( .A1(n9104), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8674), 
        .B2(n15882), .ZN(n8800) );
  NAND2_X1 U10606 ( .A1(n8650), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8805) );
  XNOR2_X1 U10607 ( .A(n8816), .B(P2_REG3_REG_12__SCAN_IN), .ZN(n12500) );
  NAND2_X1 U10608 ( .A1(n8649), .A2(n12500), .ZN(n8804) );
  NAND2_X1 U10609 ( .A1(n8665), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U10610 ( .A1(n8885), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8802) );
  NOR2_X1 U10611 ( .A1(n16202), .A2(n14795), .ZN(n8807) );
  NAND2_X1 U10612 ( .A1(n16202), .A2(n14795), .ZN(n8806) );
  XNOR2_X1 U10613 ( .A(n8808), .B(n7878), .ZN(n12192) );
  NAND2_X1 U10614 ( .A1(n12192), .A2(n10044), .ZN(n8813) );
  OR2_X1 U10615 ( .A1(n8798), .A2(n8810), .ZN(n8811) );
  XNOR2_X1 U10616 ( .A(n8811), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U10617 ( .A1(n9104), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8674), 
        .B2(n11367), .ZN(n8812) );
  NAND2_X1 U10618 ( .A1(n8650), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8821) );
  INV_X1 U10619 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8815) );
  INV_X1 U10620 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8814) );
  OAI21_X1 U10621 ( .B1(n8816), .B2(n8815), .A(n8814), .ZN(n8817) );
  AND2_X1 U10622 ( .A1(n8828), .A2(n8817), .ZN(n14799) );
  NAND2_X1 U10623 ( .A1(n8649), .A2(n14799), .ZN(n8820) );
  NAND2_X1 U10624 ( .A1(n8665), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U10625 ( .A1(n8885), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8818) );
  NAND4_X1 U10626 ( .A1(n8821), .A2(n8820), .A3(n8819), .A4(n8818), .ZN(n14472) );
  XNOR2_X1 U10627 ( .A(n14800), .B(n14327), .ZN(n14786) );
  XNOR2_X1 U10628 ( .A(n8823), .B(n8822), .ZN(n12520) );
  NAND2_X1 U10629 ( .A1(n12520), .A2(n10044), .ZN(n8827) );
  NAND2_X1 U10630 ( .A1(n8824), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8825) );
  XNOR2_X1 U10631 ( .A(n8825), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U10632 ( .A1(n9104), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8674), 
        .B2(n10901), .ZN(n8826) );
  NAND2_X1 U10633 ( .A1(n8650), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8833) );
  NAND2_X1 U10634 ( .A1(n8828), .A2(n10931), .ZN(n8829) );
  AND2_X1 U10635 ( .A1(n8840), .A2(n8829), .ZN(n14775) );
  NAND2_X1 U10636 ( .A1(n8649), .A2(n14775), .ZN(n8832) );
  NAND2_X1 U10637 ( .A1(n8665), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U10638 ( .A1(n8885), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8830) );
  NAND4_X1 U10639 ( .A1(n8833), .A2(n8832), .A3(n8831), .A4(n8830), .ZN(n14792) );
  XNOR2_X1 U10640 ( .A(n14889), .B(n14792), .ZN(n14770) );
  INV_X1 U10641 ( .A(n14770), .ZN(n14779) );
  OR2_X1 U10642 ( .A1(n14889), .A2(n14792), .ZN(n8834) );
  XNOR2_X1 U10643 ( .A(n8836), .B(n8835), .ZN(n12595) );
  NAND2_X1 U10644 ( .A1(n12595), .A2(n10044), .ZN(n8839) );
  NAND2_X1 U10645 ( .A1(n7338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8837) );
  XNOR2_X1 U10646 ( .A(n8837), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U10647 ( .A1(n9104), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8674), 
        .B2(n11864), .ZN(n8838) );
  INV_X1 U10648 ( .A(n14879), .ZN(n8846) );
  NAND2_X1 U10649 ( .A1(n8650), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U10650 ( .A1(n8840), .A2(n14456), .ZN(n8841) );
  AND2_X1 U10651 ( .A1(n8855), .A2(n8841), .ZN(n14765) );
  NAND2_X1 U10652 ( .A1(n8649), .A2(n14765), .ZN(n8844) );
  NAND2_X1 U10653 ( .A1(n8665), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U10654 ( .A1(n8885), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8842) );
  INV_X1 U10655 ( .A(n14381), .ZN(n14471) );
  XNOR2_X1 U10656 ( .A(n8846), .B(n14471), .ZN(n10101) );
  NAND2_X1 U10657 ( .A1(n14879), .A2(n14381), .ZN(n8847) );
  NAND2_X1 U10658 ( .A1(n8849), .A2(n8848), .ZN(n8850) );
  AND2_X1 U10659 ( .A1(n8851), .A2(n8850), .ZN(n12651) );
  NAND2_X1 U10660 ( .A1(n12651), .A2(n10044), .ZN(n8854) );
  NAND2_X1 U10661 ( .A1(n8585), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8852) );
  XNOR2_X1 U10662 ( .A(n8852), .B(P2_IR_REG_16__SCAN_IN), .ZN(n15849) );
  AOI22_X1 U10663 ( .A1(n9104), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8674), 
        .B2(n15849), .ZN(n8853) );
  NAND2_X1 U10664 ( .A1(n8650), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8860) );
  INV_X1 U10665 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n14384) );
  NAND2_X1 U10666 ( .A1(n8855), .A2(n14384), .ZN(n8856) );
  AND2_X1 U10667 ( .A1(n8868), .A2(n8856), .ZN(n14746) );
  NAND2_X1 U10668 ( .A1(n8649), .A2(n14746), .ZN(n8859) );
  NAND2_X1 U10669 ( .A1(n8665), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U10670 ( .A1(n8885), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8857) );
  INV_X1 U10671 ( .A(n14453), .ZN(n14470) );
  XNOR2_X1 U10672 ( .A(n14748), .B(n14470), .ZN(n14740) );
  NAND2_X1 U10673 ( .A1(n14748), .A2(n14470), .ZN(n8861) );
  XNOR2_X1 U10674 ( .A(n8863), .B(n8862), .ZN(n12822) );
  NAND2_X1 U10675 ( .A1(n12822), .A2(n10044), .ZN(n8866) );
  XNOR2_X1 U10676 ( .A(n8864), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15864) );
  AOI22_X1 U10677 ( .A1(n9104), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8674), 
        .B2(n15864), .ZN(n8865) );
  NAND2_X1 U10678 ( .A1(n8650), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8873) );
  INV_X1 U10679 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8867) );
  NAND2_X1 U10680 ( .A1(n8868), .A2(n8867), .ZN(n8869) );
  AND2_X1 U10681 ( .A1(n8883), .A2(n8869), .ZN(n14726) );
  NAND2_X1 U10682 ( .A1(n8649), .A2(n14726), .ZN(n8872) );
  NAND2_X1 U10683 ( .A1(n8665), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U10684 ( .A1(n8885), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8870) );
  XNOR2_X1 U10685 ( .A(n14867), .B(n14433), .ZN(n14731) );
  NAND2_X1 U10686 ( .A1(n14728), .A2(n14433), .ZN(n8874) );
  INV_X1 U10687 ( .A(n8875), .ZN(n8876) );
  NAND2_X1 U10688 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  NAND2_X1 U10689 ( .A1(n8879), .A2(n8878), .ZN(n12834) );
  XNOR2_X1 U10690 ( .A(n8880), .B(P2_IR_REG_18__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U10691 ( .A1(n9104), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8674), 
        .B2(n11870), .ZN(n8881) );
  NAND2_X1 U10692 ( .A1(n8883), .A2(n14434), .ZN(n8884) );
  AND2_X1 U10693 ( .A1(n8897), .A2(n8884), .ZN(n14712) );
  NAND2_X1 U10694 ( .A1(n8649), .A2(n14712), .ZN(n8889) );
  NAND2_X1 U10695 ( .A1(n8650), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U10696 ( .A1(n8665), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U10697 ( .A1(n8885), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8886) );
  NAND4_X1 U10698 ( .A1(n8889), .A2(n8888), .A3(n8887), .A4(n8886), .ZN(n14469) );
  XNOR2_X1 U10699 ( .A(n14713), .B(n14469), .ZN(n10104) );
  NAND2_X1 U10700 ( .A1(n14708), .A2(n14707), .ZN(n8891) );
  INV_X1 U10701 ( .A(n14469), .ZN(n14343) );
  NAND2_X1 U10702 ( .A1(n14861), .A2(n14343), .ZN(n8890) );
  NAND2_X1 U10703 ( .A1(n12727), .A2(n10044), .ZN(n8895) );
  AOI22_X1 U10704 ( .A1(n9104), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9093), 
        .B2(n8674), .ZN(n8894) );
  INV_X1 U10705 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U10706 ( .A1(n8897), .A2(n8896), .ZN(n8898) );
  NAND2_X1 U10707 ( .A1(n8909), .A2(n8898), .ZN(n14698) );
  NAND2_X1 U10708 ( .A1(n8650), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U10709 ( .A1(n8665), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8899) );
  AND2_X1 U10710 ( .A1(n8900), .A2(n8899), .ZN(n8902) );
  NAND2_X1 U10711 ( .A1(n8885), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8901) );
  OAI211_X1 U10712 ( .C1(n14698), .C2(n9058), .A(n8902), .B(n8901), .ZN(n14468) );
  XNOR2_X1 U10713 ( .A(n14700), .B(n14468), .ZN(n14688) );
  OR2_X1 U10714 ( .A1(n14700), .A2(n14468), .ZN(n8903) );
  INV_X1 U10715 ( .A(SI_20_), .ZN(n10776) );
  XNOR2_X1 U10716 ( .A(n8904), .B(n10776), .ZN(n8905) );
  XNOR2_X1 U10717 ( .A(n8906), .B(n8905), .ZN(n12847) );
  NAND2_X1 U10718 ( .A1(n12847), .A2(n10044), .ZN(n8908) );
  NAND2_X1 U10719 ( .A1(n9104), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U10720 ( .A1(n8909), .A2(n14414), .ZN(n8910) );
  AND2_X1 U10721 ( .A1(n8921), .A2(n8910), .ZN(n14678) );
  NAND2_X1 U10722 ( .A1(n14678), .A2(n8649), .ZN(n8913) );
  AOI22_X1 U10723 ( .A1(n8650), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n8665), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U10724 ( .A1(n8885), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8911) );
  AND2_X1 U10725 ( .A1(n14929), .A2(n14361), .ZN(n8914) );
  NAND2_X1 U10726 ( .A1(n9051), .A2(n14467), .ZN(n8915) );
  XNOR2_X1 U10727 ( .A(n8917), .B(n8916), .ZN(n12869) );
  NAND2_X1 U10728 ( .A1(n12869), .A2(n10044), .ZN(n8919) );
  NAND2_X1 U10729 ( .A1(n9104), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8918) );
  INV_X1 U10730 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U10731 ( .A1(n8921), .A2(n8920), .ZN(n8922) );
  NAND2_X1 U10732 ( .A1(n8934), .A2(n8922), .ZN(n14663) );
  OR2_X1 U10733 ( .A1(n14663), .A2(n9058), .ZN(n8925) );
  AOI22_X1 U10734 ( .A1(n8650), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n8665), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U10735 ( .A1(n8885), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8923) );
  XNOR2_X1 U10736 ( .A(n14368), .B(n14289), .ZN(n14667) );
  OR2_X1 U10737 ( .A1(n14925), .A2(n14289), .ZN(n8926) );
  NAND2_X1 U10738 ( .A1(n12882), .A2(n8927), .ZN(n8945) );
  INV_X1 U10739 ( .A(n12882), .ZN(n8929) );
  NAND2_X1 U10740 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  NAND2_X1 U10741 ( .A1(n8945), .A2(n8930), .ZN(n12682) );
  OR2_X1 U10742 ( .A1(n12682), .A2(n10024), .ZN(n8932) );
  NAND2_X1 U10743 ( .A1(n9104), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U10744 ( .A1(n8934), .A2(n8933), .ZN(n8935) );
  AND2_X1 U10745 ( .A1(n8951), .A2(n8935), .ZN(n14652) );
  NAND2_X1 U10746 ( .A1(n14652), .A2(n8649), .ZN(n8941) );
  INV_X1 U10747 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U10748 ( .A1(n8650), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U10749 ( .A1(n8665), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8936) );
  OAI211_X1 U10750 ( .C1(n8938), .C2(n10032), .A(n8937), .B(n8936), .ZN(n8939)
         );
  INV_X1 U10751 ( .A(n8939), .ZN(n8940) );
  XNOR2_X1 U10752 ( .A(n14840), .B(n14362), .ZN(n14655) );
  OR2_X1 U10753 ( .A1(n14654), .A2(n14362), .ZN(n8942) );
  NAND2_X1 U10754 ( .A1(n8943), .A2(SI_22_), .ZN(n8944) );
  NAND2_X1 U10755 ( .A1(n8945), .A2(n8944), .ZN(n8948) );
  XNOR2_X1 U10756 ( .A(n8946), .B(SI_23_), .ZN(n8947) );
  NAND2_X1 U10757 ( .A1(n9104), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8949) );
  INV_X1 U10758 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U10759 ( .A1(n8951), .A2(n8950), .ZN(n8952) );
  NAND2_X1 U10760 ( .A1(n8965), .A2(n8952), .ZN(n14638) );
  OR2_X1 U10761 ( .A1(n14638), .A2(n9058), .ZN(n8957) );
  INV_X1 U10762 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14639) );
  NAND2_X1 U10763 ( .A1(n8650), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U10764 ( .A1(n8665), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8953) );
  OAI211_X1 U10765 ( .C1(n10032), .C2(n14639), .A(n8954), .B(n8953), .ZN(n8955) );
  INV_X1 U10766 ( .A(n8955), .ZN(n8956) );
  INV_X1 U10767 ( .A(n14629), .ZN(n14630) );
  OR2_X1 U10768 ( .A1(n14914), .A2(n14401), .ZN(n8958) );
  XNOR2_X1 U10769 ( .A(n8961), .B(n8960), .ZN(n12907) );
  NAND2_X1 U10770 ( .A1(n12907), .A2(n10044), .ZN(n8963) );
  NAND2_X1 U10771 ( .A1(n9104), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8962) );
  INV_X1 U10772 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8964) );
  NAND2_X1 U10773 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  NAND2_X1 U10774 ( .A1(n8989), .A2(n8966), .ZN(n14621) );
  INV_X1 U10775 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14622) );
  NAND2_X1 U10776 ( .A1(n8650), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8968) );
  NAND2_X1 U10777 ( .A1(n8665), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8967) );
  OAI211_X1 U10778 ( .C1(n14622), .C2(n10032), .A(n8968), .B(n8967), .ZN(n8969) );
  INV_X1 U10779 ( .A(n8969), .ZN(n8970) );
  NAND2_X1 U10780 ( .A1(n14830), .A2(n14598), .ZN(n9053) );
  OR2_X1 U10781 ( .A1(n14830), .A2(n14598), .ZN(n8972) );
  NAND2_X1 U10782 ( .A1(n14830), .A2(n14633), .ZN(n8973) );
  XNOR2_X1 U10783 ( .A(n8975), .B(n8974), .ZN(n14966) );
  NAND2_X1 U10784 ( .A1(n14966), .A2(n10044), .ZN(n8977) );
  NAND2_X1 U10785 ( .A1(n9104), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8976) );
  XNOR2_X1 U10786 ( .A(n8989), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n14604) );
  NAND2_X1 U10787 ( .A1(n14604), .A2(n8649), .ZN(n8983) );
  INV_X1 U10788 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U10789 ( .A1(n8650), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U10790 ( .A1(n8665), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8978) );
  OAI211_X1 U10791 ( .C1(n8980), .C2(n10032), .A(n8979), .B(n8978), .ZN(n8981)
         );
  INV_X1 U10792 ( .A(n8981), .ZN(n8982) );
  XNOR2_X1 U10793 ( .A(n14601), .B(n14405), .ZN(n10108) );
  NAND2_X1 U10794 ( .A1(n14963), .A2(n10044), .ZN(n8986) );
  NAND2_X1 U10795 ( .A1(n9104), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8985) );
  OAI21_X1 U10796 ( .B1(n8989), .B2(n8988), .A(n8987), .ZN(n8991) );
  NAND2_X1 U10797 ( .A1(n14582), .A2(n8649), .ZN(n8997) );
  INV_X1 U10798 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U10799 ( .A1(n8650), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U10800 ( .A1(n8665), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8992) );
  OAI211_X1 U10801 ( .C1(n8994), .C2(n10032), .A(n8993), .B(n8992), .ZN(n8995)
         );
  INV_X1 U10802 ( .A(n8995), .ZN(n8996) );
  XNOR2_X1 U10803 ( .A(n14819), .B(n14466), .ZN(n10109) );
  NAND2_X1 U10804 ( .A1(n14584), .A2(n14599), .ZN(n8998) );
  NAND2_X1 U10805 ( .A1(n14585), .A2(n8998), .ZN(n9233) );
  XNOR2_X1 U10806 ( .A(n14569), .B(n14580), .ZN(n10110) );
  NAND2_X1 U10807 ( .A1(n9000), .A2(n8999), .ZN(n9004) );
  INV_X1 U10808 ( .A(n9001), .ZN(n9002) );
  NAND2_X1 U10809 ( .A1(n9002), .A2(SI_27_), .ZN(n9003) );
  NAND2_X1 U10810 ( .A1(n9004), .A2(n9003), .ZN(n9009) );
  INV_X1 U10811 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13081) );
  INV_X1 U10812 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9760) );
  MUX2_X1 U10813 ( .A(n13081), .B(n9760), .S(n10689), .Z(n9005) );
  NAND2_X1 U10814 ( .A1(n9005), .A2(n13534), .ZN(n9102) );
  INV_X1 U10815 ( .A(n9005), .ZN(n9006) );
  NAND2_X1 U10816 ( .A1(n9006), .A2(SI_28_), .ZN(n9007) );
  NAND2_X1 U10817 ( .A1(n9102), .A2(n9007), .ZN(n9008) );
  NAND2_X1 U10818 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  NAND2_X1 U10819 ( .A1(n13080), .A2(n10044), .ZN(n9012) );
  NAND2_X1 U10820 ( .A1(n9104), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9011) );
  NAND2_X1 U10821 ( .A1(n9013), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13084) );
  INV_X1 U10822 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U10823 ( .A1(n9015), .A2(n9014), .ZN(n9016) );
  NAND2_X1 U10824 ( .A1(n13084), .A2(n9016), .ZN(n14558) );
  OR2_X1 U10825 ( .A1(n14558), .A2(n9058), .ZN(n9022) );
  INV_X1 U10826 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U10827 ( .A1(n8650), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9018) );
  NAND2_X1 U10828 ( .A1(n8665), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9017) );
  OAI211_X1 U10829 ( .C1(n10032), .C2(n9019), .A(n9018), .B(n9017), .ZN(n9020)
         );
  INV_X1 U10830 ( .A(n9020), .ZN(n9021) );
  NAND2_X1 U10831 ( .A1(n9251), .A2(n14318), .ZN(n9100) );
  NAND2_X1 U10832 ( .A1(n14560), .A2(n14465), .ZN(n9023) );
  OAI21_X1 U10833 ( .B1(n9024), .B2(n14351), .A(n9101), .ZN(n9025) );
  INV_X1 U10834 ( .A(n14362), .ZN(n14632) );
  NAND2_X1 U10835 ( .A1(n11395), .A2(n11399), .ZN(n10093) );
  INV_X1 U10836 ( .A(n10093), .ZN(n11393) );
  NAND2_X1 U10837 ( .A1(n11394), .A2(n11724), .ZN(n9028) );
  NAND2_X1 U10838 ( .A1(n9029), .A2(n9900), .ZN(n9030) );
  NAND2_X1 U10839 ( .A1(n9031), .A2(n11603), .ZN(n9032) );
  INV_X2 U10840 ( .A(n11840), .ZN(n11418) );
  NAND2_X1 U10841 ( .A1(n14480), .A2(n11418), .ZN(n9033) );
  INV_X1 U10842 ( .A(n14480), .ZN(n9922) );
  NAND2_X1 U10843 ( .A1(n9922), .A2(n11840), .ZN(n9034) );
  INV_X1 U10844 ( .A(n14479), .ZN(n9924) );
  NOR2_X1 U10845 ( .A1(n12295), .A2(n14478), .ZN(n9036) );
  NAND2_X1 U10846 ( .A1(n12295), .A2(n14478), .ZN(n9035) );
  INV_X1 U10847 ( .A(n11937), .ZN(n9037) );
  NAND2_X1 U10848 ( .A1(n11944), .A2(n12038), .ZN(n9038) );
  INV_X1 U10849 ( .A(n12140), .ZN(n12138) );
  NAND2_X1 U10850 ( .A1(n16186), .A2(n14475), .ZN(n12330) );
  AND2_X1 U10851 ( .A1(n12329), .A2(n12330), .ZN(n9039) );
  NAND2_X1 U10852 ( .A1(n12331), .A2(n9039), .ZN(n12328) );
  INV_X1 U10853 ( .A(n16202), .ZN(n12504) );
  NAND2_X1 U10854 ( .A1(n12504), .A2(n14795), .ZN(n9042) );
  OR2_X1 U10855 ( .A1(n12504), .A2(n14795), .ZN(n9041) );
  NAND2_X1 U10856 ( .A1(n12398), .A2(n9042), .ZN(n14790) );
  INV_X1 U10857 ( .A(n14786), .ZN(n14789) );
  NAND2_X1 U10858 ( .A1(n14800), .A2(n14327), .ZN(n9043) );
  INV_X1 U10859 ( .A(n14792), .ZN(n12574) );
  OR2_X1 U10860 ( .A1(n14889), .A2(n12574), .ZN(n9044) );
  NAND2_X1 U10861 ( .A1(n14889), .A2(n12574), .ZN(n9045) );
  NAND2_X1 U10862 ( .A1(n14879), .A2(n14471), .ZN(n9046) );
  NAND2_X1 U10863 ( .A1(n14737), .A2(n14740), .ZN(n14736) );
  INV_X1 U10864 ( .A(n14731), .ZN(n9047) );
  NOR2_X1 U10865 ( .A1(n14713), .A2(n14343), .ZN(n9050) );
  XNOR2_X1 U10866 ( .A(n9051), .B(n14467), .ZN(n14681) );
  INV_X1 U10867 ( .A(n9053), .ZN(n14594) );
  NAND2_X1 U10868 ( .A1(n14601), .A2(n14405), .ZN(n14577) );
  NOR2_X1 U10869 ( .A1(n14584), .A2(n14466), .ZN(n9236) );
  INV_X1 U10870 ( .A(n14580), .ZN(n9054) );
  NAND2_X1 U10871 ( .A1(n9094), .A2(n8503), .ZN(n9056) );
  NAND2_X1 U10872 ( .A1(n10974), .A2(n9093), .ZN(n9055) );
  AOI211_X1 U10873 ( .C1(n14351), .C2(n9057), .A(n14719), .B(n9109), .ZN(n9066) );
  OR2_X1 U10874 ( .A1(n13084), .A2(n9058), .ZN(n9063) );
  INV_X1 U10875 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13083) );
  NAND2_X1 U10876 ( .A1(n8650), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9060) );
  NAND2_X1 U10877 ( .A1(n8665), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9059) );
  OAI211_X1 U10878 ( .C1(n13083), .C2(n10032), .A(n9060), .B(n9059), .ZN(n9061) );
  INV_X1 U10879 ( .A(n9061), .ZN(n9062) );
  NAND2_X1 U10880 ( .A1(n9063), .A2(n9062), .ZN(n14464) );
  INV_X1 U10881 ( .A(n14464), .ZN(n9107) );
  INV_X1 U10882 ( .A(n9064), .ZN(n9065) );
  OAI22_X1 U10883 ( .A1(n9107), .A2(n14600), .B1(n9054), .B2(n14794), .ZN(
        n14356) );
  AND2_X1 U10884 ( .A1(n11593), .A2(n11418), .ZN(n11417) );
  INV_X1 U10885 ( .A(n11508), .ZN(n12321) );
  NAND2_X1 U10886 ( .A1(n11417), .A2(n12321), .ZN(n11669) );
  OR2_X2 U10887 ( .A1(n11898), .A2(n16133), .ZN(n11943) );
  AND2_X2 U10888 ( .A1(n14929), .A2(n14696), .ZN(n14676) );
  NAND2_X1 U10889 ( .A1(n14914), .A2(n14651), .ZN(n14637) );
  OR2_X2 U10890 ( .A1(n14637), .A2(n14830), .ZN(n14618) );
  OAI211_X1 U10891 ( .C1(n9251), .C2(n9241), .A(n7201), .B(n14267), .ZN(n14562) );
  XNOR2_X1 U10892 ( .A(P2_B_REG_SCAN_IN), .B(n12688), .ZN(n9077) );
  AND2_X1 U10893 ( .A1(n14967), .A2(n9077), .ZN(n9078) );
  INV_X1 U10894 ( .A(n9097), .ZN(n15815) );
  INV_X1 U10895 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15814) );
  AOI22_X1 U10896 ( .A1(n15815), .A2(n15814), .B1(n14965), .B2(n14967), .ZN(
        n10826) );
  NAND2_X1 U10897 ( .A1(n9079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9081) );
  INV_X1 U10898 ( .A(n10131), .ZN(n10827) );
  OR2_X1 U10899 ( .A1(n10826), .A2(n15818), .ZN(n15812) );
  NOR4_X1 U10900 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9086) );
  NOR4_X1 U10901 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9085) );
  NOR4_X1 U10902 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9084) );
  NOR4_X1 U10903 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9083) );
  NAND4_X1 U10904 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(n9092)
         );
  NOR2_X1 U10905 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9090) );
  NOR4_X1 U10906 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9089) );
  NOR4_X1 U10907 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9088) );
  NOR4_X1 U10908 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9087) );
  NAND4_X1 U10909 ( .A1(n9090), .A2(n9089), .A3(n9088), .A4(n9087), .ZN(n9091)
         );
  OAI21_X1 U10910 ( .B1(n9092), .B2(n9091), .A(n15815), .ZN(n10825) );
  NAND2_X1 U10911 ( .A1(n10896), .A2(n10832), .ZN(n11514) );
  NAND3_X1 U10912 ( .A1(n10825), .A2(n10838), .A3(n11514), .ZN(n9095) );
  NAND2_X1 U10913 ( .A1(n14965), .A2(n12688), .ZN(n9096) );
  INV_X1 U10914 ( .A(n15820), .ZN(n9098) );
  NOR2_X1 U10915 ( .A1(n9251), .A2(n14896), .ZN(n9099) );
  INV_X1 U10916 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15765) );
  INV_X1 U10917 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14959) );
  MUX2_X1 U10918 ( .A(n15765), .B(n14959), .S(n10178), .Z(n10016) );
  XNOR2_X1 U10919 ( .A(n10016), .B(SI_29_), .ZN(n10018) );
  NAND2_X1 U10920 ( .A1(n14958), .A2(n10044), .ZN(n9106) );
  NAND2_X1 U10921 ( .A1(n9104), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9105) );
  XNOR2_X1 U10922 ( .A(n9111), .B(n9110), .ZN(n9113) );
  NAND2_X1 U10923 ( .A1(n9113), .A2(n9112), .ZN(n9120) );
  INV_X1 U10924 ( .A(n13321), .ZN(n10900) );
  NAND2_X1 U10925 ( .A1(n10900), .A2(P2_B_REG_SCAN_IN), .ZN(n9114) );
  NAND2_X1 U10926 ( .A1(n14791), .A2(n9114), .ZN(n14546) );
  NAND2_X1 U10927 ( .A1(n8650), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U10928 ( .A1(n8885), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U10929 ( .A1(n8665), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9115) );
  INV_X1 U10930 ( .A(n9118), .ZN(n9119) );
  NAND2_X1 U10931 ( .A1(n9120), .A2(n9119), .ZN(n13082) );
  INV_X1 U10932 ( .A(n13086), .ZN(n9122) );
  AOI21_X1 U10933 ( .B1(n7201), .B2(n13086), .A(n14300), .ZN(n9121) );
  NAND2_X1 U10934 ( .A1(n14551), .A2(n9121), .ZN(n13088) );
  OAI21_X1 U10935 ( .B1(n9122), .B2(n16201), .A(n13088), .ZN(n9123) );
  NOR2_X1 U10936 ( .A1(n13082), .A2(n9123), .ZN(n9124) );
  INV_X1 U10937 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n13843) );
  INV_X1 U10938 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n9156) );
  NOR2_X1 U10939 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n9156), .ZN(n9126) );
  AOI21_X1 U10940 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n9156), .A(n9126), .ZN(
        n9163) );
  INV_X1 U10941 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9154) );
  INV_X1 U10942 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n12305) );
  XNOR2_X1 U10943 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9212) );
  INV_X1 U10944 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15936) );
  XNOR2_X1 U10945 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9207) );
  INV_X1 U10946 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9148) );
  INV_X1 U10947 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9146) );
  XNOR2_X1 U10948 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9201) );
  INV_X1 U10949 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9144) );
  XNOR2_X1 U10950 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9197) );
  INV_X1 U10951 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n9140) );
  AND2_X1 U10952 ( .A1(n9137), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n9138) );
  XNOR2_X1 U10953 ( .A(n9128), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n9175) );
  NOR2_X1 U10954 ( .A1(n9129), .A2(n9130), .ZN(n9132) );
  XNOR2_X1 U10955 ( .A(n9130), .B(n9129), .ZN(n9180) );
  NOR2_X1 U10956 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n9180), .ZN(n9131) );
  XNOR2_X1 U10957 ( .A(n9134), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n9166) );
  NOR2_X1 U10958 ( .A1(n9167), .A2(n9166), .ZN(n9133) );
  NOR2_X1 U10959 ( .A1(n9140), .A2(n9139), .ZN(n9142) );
  XNOR2_X1 U10960 ( .A(n9140), .B(n9139), .ZN(n9193) );
  NAND2_X1 U10961 ( .A1(n9197), .A2(n9196), .ZN(n9143) );
  NAND2_X1 U10962 ( .A1(n9201), .A2(n9202), .ZN(n9145) );
  XOR2_X1 U10963 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n9164) );
  INV_X1 U10964 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n9149) );
  OR2_X1 U10965 ( .A1(n9149), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n9150) );
  XOR2_X1 U10966 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n9214) );
  NOR2_X1 U10967 ( .A1(n9215), .A2(n9214), .ZN(n9153) );
  AOI21_X1 U10968 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n9154), .A(n9153), .ZN(
        n9162) );
  NAND2_X1 U10969 ( .A1(n9163), .A2(n9162), .ZN(n9155) );
  INV_X1 U10970 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9157) );
  NOR2_X1 U10971 ( .A1(n9158), .A2(n9157), .ZN(n9160) );
  XOR2_X1 U10972 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n9158), .Z(n9218) );
  NOR2_X1 U10973 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n9218), .ZN(n9159) );
  NOR2_X1 U10974 ( .A1(n9160), .A2(n9159), .ZN(n9221) );
  XOR2_X1 U10975 ( .A(n9221), .B(P1_ADDR_REG_17__SCAN_IN), .Z(n9222) );
  XNOR2_X1 U10976 ( .A(n13843), .B(n9222), .ZN(n9161) );
  AND2_X1 U10977 ( .A1(n9161), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n9219) );
  XNOR2_X1 U10978 ( .A(n9161), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(n15989) );
  XNOR2_X1 U10979 ( .A(n9163), .B(n9162), .ZN(n9216) );
  XOR2_X1 U10980 ( .A(n9165), .B(n9164), .Z(n15961) );
  XNOR2_X1 U10981 ( .A(n9167), .B(n9166), .ZN(n9168) );
  XNOR2_X1 U10982 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n9168), .ZN(n15945) );
  INV_X1 U10983 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9173) );
  NOR2_X1 U10984 ( .A1(n9172), .A2(n9173), .ZN(n9174) );
  OAI21_X1 U10985 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9171), .A(n9170), .ZN(
        n15937) );
  NAND2_X1 U10986 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15937), .ZN(n15998) );
  XOR2_X1 U10987 ( .A(n9176), .B(n9175), .Z(n9177) );
  NOR2_X1 U10988 ( .A1(n9178), .A2(n9177), .ZN(n9179) );
  XNOR2_X1 U10989 ( .A(n9178), .B(n9177), .ZN(n15940) );
  INV_X1 U10990 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15939) );
  NOR2_X1 U10991 ( .A1(n15940), .A2(n15939), .ZN(n15938) );
  XOR2_X1 U10992 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n9180), .Z(n9182) );
  NAND2_X1 U10993 ( .A1(n9181), .A2(n9182), .ZN(n9183) );
  INV_X1 U10994 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15942) );
  XNOR2_X1 U10995 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n9185) );
  XNOR2_X1 U10996 ( .A(n9185), .B(n9184), .ZN(n9187) );
  NOR2_X1 U10997 ( .A1(n9186), .A2(n9187), .ZN(n9188) );
  INV_X1 U10998 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15947) );
  NOR2_X1 U10999 ( .A1(n15948), .A2(n15947), .ZN(n15946) );
  XOR2_X1 U11000 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), .Z(
        n9189) );
  XNOR2_X1 U11001 ( .A(n9190), .B(n9189), .ZN(n15993) );
  NAND2_X1 U11002 ( .A1(n15994), .A2(n15993), .ZN(n9191) );
  NOR2_X1 U11003 ( .A1(n15994), .A2(n15993), .ZN(n15992) );
  AOI21_X2 U11004 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(n9191), .A(n15992), .ZN(
        n9194) );
  INV_X1 U11005 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9192) );
  NOR2_X1 U11006 ( .A1(n9194), .A2(n9192), .ZN(n9195) );
  XOR2_X1 U11007 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9193), .Z(n15951) );
  XNOR2_X1 U11008 ( .A(n9197), .B(n9196), .ZN(n9199) );
  NAND2_X1 U11009 ( .A1(n9198), .A2(n9199), .ZN(n9200) );
  INV_X1 U11010 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15953) );
  NAND2_X1 U11011 ( .A1(n15954), .A2(n15953), .ZN(n15952) );
  NAND2_X1 U11012 ( .A1(n9200), .A2(n15952), .ZN(n15957) );
  XNOR2_X1 U11013 ( .A(n9202), .B(n9201), .ZN(n15956) );
  XNOR2_X1 U11014 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9204) );
  XNOR2_X1 U11015 ( .A(n9204), .B(n9203), .ZN(n15964) );
  NAND2_X1 U11016 ( .A1(n15965), .A2(n15964), .ZN(n9205) );
  XOR2_X1 U11017 ( .A(n9207), .B(n9206), .Z(n9208) );
  NAND2_X1 U11018 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  INV_X1 U11019 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15968) );
  XNOR2_X1 U11020 ( .A(n9212), .B(n9211), .ZN(n15971) );
  NAND2_X1 U11021 ( .A1(n15972), .A2(n15971), .ZN(n15970) );
  XNOR2_X1 U11022 ( .A(n9215), .B(n9214), .ZN(n15975) );
  INV_X1 U11023 ( .A(n15979), .ZN(n15980) );
  INV_X1 U11024 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15982) );
  NAND2_X1 U11025 ( .A1(n9217), .A2(n9216), .ZN(n15981) );
  NAND2_X1 U11026 ( .A1(n15982), .A2(n15981), .ZN(n15978) );
  XNOR2_X1 U11027 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n9218), .ZN(n15984) );
  NOR2_X2 U11028 ( .A1(n9219), .A2(n15987), .ZN(n15991) );
  INV_X1 U11029 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9220) );
  NOR2_X1 U11030 ( .A1(n9221), .A2(n9220), .ZN(n9224) );
  NOR2_X1 U11031 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n9222), .ZN(n9223) );
  NOR2_X1 U11032 ( .A1(n9224), .A2(n9223), .ZN(n9227) );
  INV_X1 U11033 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U11034 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9229), .ZN(n9225) );
  OAI21_X1 U11035 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9229), .A(n9225), .ZN(
        n9226) );
  XNOR2_X1 U11036 ( .A(n9227), .B(n9226), .ZN(n15990) );
  NOR2_X1 U11037 ( .A1(n9227), .A2(n9226), .ZN(n9228) );
  AOI21_X1 U11038 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9229), .A(n9228), .ZN(
        n9231) );
  XNOR2_X1 U11039 ( .A(n9231), .B(n9230), .ZN(n9232) );
  AND2_X1 U11040 ( .A1(n9233), .A2(n10110), .ZN(n9234) );
  INV_X1 U11041 ( .A(n9249), .ZN(n14573) );
  OAI22_X1 U11042 ( .A1(n14318), .A2(n14600), .B1(n14599), .B2(n14794), .ZN(
        n9240) );
  OR3_X1 U11043 ( .A1(n14576), .A2(n9236), .A3(n10110), .ZN(n9237) );
  AOI21_X1 U11044 ( .B1(n9238), .B2(n9237), .A(n14719), .ZN(n9239) );
  INV_X1 U11045 ( .A(n9241), .ZN(n9242) );
  OAI211_X1 U11046 ( .C1(n9248), .C2(n14581), .A(n9242), .B(n14267), .ZN(
        n14571) );
  OAI22_X1 U11047 ( .A1(n9249), .A2(n14897), .B1(n9248), .B2(n14896), .ZN(
        n9244) );
  INV_X1 U11048 ( .A(n9244), .ZN(n9245) );
  NAND2_X1 U11049 ( .A1(n9246), .A2(n9245), .ZN(P2_U3526) );
  OAI22_X1 U11050 ( .A1(n9249), .A2(n14953), .B1(n9248), .B2(n14951), .ZN(
        n9250) );
  NAND2_X1 U11051 ( .A1(n9252), .A2(n8467), .ZN(P2_U3495) );
  INV_X1 U11052 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U11053 ( .A1(n9256), .A2(n9255), .ZN(P2_U3528) );
  INV_X1 U11054 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U11055 ( .A1(n9257), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9390) );
  INV_X1 U11056 ( .A(n9390), .ZN(n9258) );
  NAND2_X1 U11057 ( .A1(n9259), .A2(n9258), .ZN(n9378) );
  NAND2_X1 U11058 ( .A1(n9260), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9261) );
  NAND2_X1 U11059 ( .A1(n10157), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9263) );
  INV_X1 U11060 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10700) );
  NAND2_X1 U11061 ( .A1(n10700), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9262) );
  NAND2_X1 U11062 ( .A1(n9402), .A2(n9401), .ZN(n9264) );
  NAND2_X1 U11063 ( .A1(n9264), .A2(n9263), .ZN(n9415) );
  NAND2_X1 U11064 ( .A1(n10207), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9266) );
  INV_X1 U11065 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10749) );
  NAND2_X1 U11066 ( .A1(n10749), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9265) );
  NAND2_X1 U11067 ( .A1(n9415), .A2(n9414), .ZN(n9267) );
  NAND2_X1 U11068 ( .A1(n10179), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9269) );
  INV_X1 U11069 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10201) );
  NAND2_X1 U11070 ( .A1(n10201), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U11071 ( .A1(n10183), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9271) );
  NAND2_X1 U11072 ( .A1(n10195), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11073 ( .A1(n10227), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n9272) );
  NAND2_X1 U11074 ( .A1(n9454), .A2(n9272), .ZN(n9274) );
  NAND2_X1 U11075 ( .A1(n10224), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U11076 ( .A1(n10235), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U11077 ( .A1(n10237), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11078 ( .A1(n9276), .A2(n9275), .ZN(n9471) );
  NAND2_X1 U11079 ( .A1(n10241), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11080 ( .A1(n10243), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11081 ( .A1(n10359), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11082 ( .A1(n10360), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U11083 ( .A1(n10365), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U11084 ( .A1(n10367), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U11085 ( .A1(n10476), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n9284) );
  NAND2_X1 U11086 ( .A1(n10471), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n9283) );
  NAND2_X1 U11087 ( .A1(n10633), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U11088 ( .A1(n10635), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U11089 ( .A1(n10822), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U11090 ( .A1(n10824), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U11091 ( .A1(n11186), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9291) );
  INV_X1 U11092 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11179) );
  NAND2_X1 U11093 ( .A1(n11179), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9290) );
  NAND2_X1 U11094 ( .A1(n11435), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11095 ( .A1(n11425), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9292) );
  INV_X1 U11096 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11615) );
  NAND2_X1 U11097 ( .A1(n11615), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n9295) );
  INV_X1 U11098 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11618) );
  NAND2_X1 U11099 ( .A1(n11618), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11100 ( .A1(n11925), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9297) );
  INV_X1 U11101 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11923) );
  NAND2_X1 U11102 ( .A1(n11923), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n9296) );
  INV_X1 U11103 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12132) );
  NAND2_X1 U11104 ( .A1(n12132), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9299) );
  INV_X1 U11105 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12720) );
  NAND2_X1 U11106 ( .A1(n12720), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9298) );
  INV_X1 U11107 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12848) );
  NAND2_X1 U11108 ( .A1(n12848), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9301) );
  INV_X1 U11109 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12441) );
  NAND2_X1 U11110 ( .A1(n12441), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9300) );
  INV_X1 U11111 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12870) );
  NAND2_X1 U11112 ( .A1(n12870), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9303) );
  INV_X1 U11113 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n12565) );
  NAND2_X1 U11114 ( .A1(n12565), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9302) );
  AND2_X1 U11115 ( .A1(n9303), .A2(n9302), .ZN(n9687) );
  INV_X1 U11116 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9304) );
  NAND2_X1 U11117 ( .A1(n9304), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9306) );
  INV_X1 U11118 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12684) );
  NAND2_X1 U11119 ( .A1(n12684), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9305) );
  AND2_X1 U11120 ( .A1(n9306), .A2(n9305), .ZN(n9701) );
  INV_X1 U11121 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9307) );
  XNOR2_X1 U11122 ( .A(n9307), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U11123 ( .A1(n9307), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9308) );
  INV_X1 U11124 ( .A(n9729), .ZN(n9309) );
  NAND2_X1 U11125 ( .A1(n9309), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U11126 ( .A1(n15772), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U11127 ( .A1(n14969), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U11128 ( .A1(n9315), .A2(n9313), .ZN(n9373) );
  INV_X1 U11129 ( .A(n9373), .ZN(n9314) );
  INV_X1 U11130 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15766) );
  NAND2_X1 U11131 ( .A1(n15766), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9319) );
  INV_X1 U11132 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14964) );
  NAND2_X1 U11133 ( .A1(n14964), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11134 ( .A1(n9319), .A2(n9317), .ZN(n9743) );
  INV_X1 U11135 ( .A(n9743), .ZN(n9318) );
  NAND2_X1 U11136 ( .A1(n9744), .A2(n9318), .ZN(n9320) );
  NAND2_X1 U11137 ( .A1(n12941), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U11138 ( .A1(n13323), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9321) );
  NAND2_X1 U11139 ( .A1(n9758), .A2(n9321), .ZN(n9755) );
  XNOR2_X1 U11140 ( .A(n9757), .B(n9755), .ZN(n12265) );
  NOR2_X1 U11141 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n9326) );
  NAND4_X1 U11142 ( .A1(n9326), .A2(n9325), .A3(n9324), .A4(n9583), .ZN(n9616)
         );
  NAND3_X1 U11143 ( .A1(n9486), .A2(n9328), .A3(n9327), .ZN(n9329) );
  NOR2_X1 U11144 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n9334) );
  NAND4_X1 U11145 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n9335)
         );
  NAND2_X1 U11146 ( .A1(n9339), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U11147 ( .A1(n12265), .A2(n13241), .ZN(n9345) );
  NAND2_X2 U11148 ( .A1(n9405), .A2(n10178), .ZN(n9443) );
  INV_X1 U11149 ( .A(SI_27_), .ZN(n13632) );
  INV_X1 U11150 ( .A(n9749), .ZN(n9356) );
  INV_X1 U11151 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9355) );
  NAND2_X1 U11152 ( .A1(n9749), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U11153 ( .A1(n9764), .A2(n9357), .ZN(n13933) );
  NAND2_X1 U11154 ( .A1(n13933), .A2(n9778), .ZN(n9366) );
  INV_X1 U11155 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n14205) );
  NAND2_X1 U11156 ( .A1(n9795), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U11157 ( .A1(n9796), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9362) );
  OAI211_X1 U11158 ( .C1(n9799), .C2(n14205), .A(n9363), .B(n9362), .ZN(n9364)
         );
  INV_X1 U11159 ( .A(n9364), .ZN(n9365) );
  NAND2_X1 U11160 ( .A1(n9735), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U11161 ( .A1(n9747), .A2(n9367), .ZN(n13956) );
  NAND2_X1 U11162 ( .A1(n13956), .A2(n9778), .ZN(n9372) );
  INV_X1 U11163 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n14212) );
  NAND2_X1 U11164 ( .A1(n9795), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U11165 ( .A1(n9796), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9368) );
  OAI211_X1 U11166 ( .C1(n9799), .C2(n14212), .A(n9369), .B(n9368), .ZN(n9370)
         );
  INV_X1 U11167 ( .A(n9370), .ZN(n9371) );
  XNOR2_X1 U11168 ( .A(n9374), .B(n9373), .ZN(n11889) );
  NAND2_X1 U11169 ( .A1(n11889), .A2(n13241), .ZN(n9376) );
  INV_X1 U11170 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10603) );
  INV_X1 U11171 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11647) );
  INV_X1 U11172 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10484) );
  NAND2_X1 U11173 ( .A1(n9377), .A2(n9390), .ZN(n9379) );
  AND2_X1 U11174 ( .A1(n9379), .A2(n9378), .ZN(n10174) );
  INV_X1 U11175 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9381) );
  OR2_X1 U11176 ( .A1(n9405), .A2(n10526), .ZN(n9382) );
  NAND2_X1 U11177 ( .A1(n16035), .A2(n9393), .ZN(n13098) );
  NAND2_X1 U11178 ( .A1(n13738), .A2(n11640), .ZN(n13096) );
  NAND2_X1 U11179 ( .A1(n13098), .A2(n13096), .ZN(n11641) );
  INV_X1 U11180 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10523) );
  INV_X1 U11181 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10513) );
  OR2_X1 U11182 ( .A1(n9407), .A2(n10513), .ZN(n9387) );
  NAND2_X1 U11183 ( .A1(n13244), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9386) );
  INV_X1 U11184 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U11185 ( .A1(n10381), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9389) );
  AND2_X1 U11186 ( .A1(n9390), .A2(n9389), .ZN(n9392) );
  OAI21_X1 U11187 ( .B1(n10689), .B2(n9392), .A(n9391), .ZN(n14260) );
  NAND2_X1 U11188 ( .A1(n13740), .A2(n10597), .ZN(n11642) );
  NAND2_X1 U11189 ( .A1(n11641), .A2(n11642), .ZN(n9395) );
  INV_X1 U11190 ( .A(n11640), .ZN(n9393) );
  OR2_X1 U11191 ( .A1(n13738), .A2(n9393), .ZN(n9394) );
  NAND2_X1 U11192 ( .A1(n9395), .A2(n9394), .ZN(n16030) );
  INV_X1 U11193 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10488) );
  OR2_X1 U11194 ( .A1(n13246), .A2(n10488), .ZN(n9399) );
  INV_X1 U11195 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10487) );
  OR2_X1 U11196 ( .A1(n9407), .A2(n10487), .ZN(n9398) );
  INV_X1 U11197 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n16044) );
  OR2_X1 U11198 ( .A1(n9605), .A2(n16044), .ZN(n9396) );
  XNOR2_X1 U11199 ( .A(n9402), .B(n9401), .ZN(n10164) );
  OR2_X1 U11200 ( .A1(n9443), .A2(SI_2_), .ZN(n9403) );
  OR2_X1 U11201 ( .A1(n13523), .A2(n8055), .ZN(n9406) );
  NAND2_X1 U11202 ( .A1(n13244), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9411) );
  INV_X1 U11203 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10493) );
  OR2_X1 U11204 ( .A1(n9407), .A2(n10493), .ZN(n9410) );
  INV_X1 U11205 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10494) );
  OR2_X1 U11206 ( .A1(n13246), .A2(n10494), .ZN(n9409) );
  OR2_X1 U11207 ( .A1(n9605), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9408) );
  XNOR2_X1 U11208 ( .A(n9415), .B(n9414), .ZN(n10158) );
  BUF_X1 U11209 ( .A(n9443), .Z(n9730) );
  OR2_X1 U11210 ( .A1(n9730), .A2(SI_3_), .ZN(n9416) );
  NAND2_X1 U11211 ( .A1(n13522), .A2(n10737), .ZN(n13108) );
  INV_X1 U11212 ( .A(n10737), .ZN(n16053) );
  NAND2_X1 U11213 ( .A1(n13522), .A2(n16053), .ZN(n9418) );
  NAND2_X1 U11214 ( .A1(n13244), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9423) );
  INV_X1 U11215 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10518) );
  OR2_X1 U11216 ( .A1(n9407), .A2(n10518), .ZN(n9422) );
  NAND2_X1 U11217 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9419) );
  AND2_X1 U11218 ( .A1(n9434), .A2(n9419), .ZN(n11587) );
  OR2_X1 U11219 ( .A1(n9605), .A2(n11587), .ZN(n9421) );
  INV_X1 U11220 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10531) );
  OR2_X1 U11221 ( .A1(n13246), .A2(n10531), .ZN(n9420) );
  NAND4_X1 U11222 ( .A1(n9423), .A2(n9422), .A3(n9421), .A4(n9420), .ZN(n13521) );
  NAND2_X1 U11223 ( .A1(n9412), .A2(n9424), .ZN(n9425) );
  NOR2_X1 U11224 ( .A1(n9425), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9456) );
  INV_X1 U11225 ( .A(n9456), .ZN(n9428) );
  NAND2_X1 U11226 ( .A1(n9425), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9426) );
  MUX2_X1 U11227 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9426), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9427) );
  XNOR2_X1 U11228 ( .A(n9430), .B(n9429), .ZN(n10170) );
  OR2_X1 U11229 ( .A1(n9705), .A2(n10170), .ZN(n9432) );
  OR2_X1 U11230 ( .A1(n9730), .A2(SI_4_), .ZN(n9431) );
  OAI211_X1 U11231 ( .C1(n13752), .C2(n10431), .A(n9432), .B(n9431), .ZN(
        n13111) );
  INV_X1 U11232 ( .A(n13111), .ZN(n11106) );
  NAND2_X1 U11233 ( .A1(n13521), .A2(n11106), .ZN(n9433) );
  NAND2_X1 U11234 ( .A1(n13244), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9439) );
  INV_X1 U11235 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10502) );
  OR2_X1 U11236 ( .A1(n9407), .A2(n10502), .ZN(n9438) );
  NAND2_X1 U11237 ( .A1(n9434), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9435) );
  AND2_X1 U11238 ( .A1(n9447), .A2(n9435), .ZN(n11762) );
  OR2_X1 U11239 ( .A1(n9605), .A2(n11762), .ZN(n9437) );
  INV_X1 U11240 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10503) );
  OR2_X1 U11241 ( .A1(n13246), .A2(n10503), .ZN(n9436) );
  NAND4_X1 U11242 ( .A1(n9439), .A2(n9438), .A3(n9437), .A4(n9436), .ZN(n13520) );
  XNOR2_X1 U11243 ( .A(n9440), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10519) );
  XNOR2_X1 U11244 ( .A(n9442), .B(n9441), .ZN(n10161) );
  OR2_X1 U11245 ( .A1(n9730), .A2(SI_5_), .ZN(n9444) );
  OAI211_X1 U11246 ( .C1(n10519), .C2(n10431), .A(n9445), .B(n9444), .ZN(
        n11763) );
  OR2_X1 U11247 ( .A1(n13520), .A2(n11763), .ZN(n13114) );
  NAND2_X1 U11248 ( .A1(n13520), .A2(n11763), .ZN(n13115) );
  INV_X1 U11249 ( .A(n11763), .ZN(n11305) );
  OR2_X1 U11250 ( .A1(n13520), .A2(n11305), .ZN(n9446) );
  NAND2_X1 U11251 ( .A1(n13244), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9452) );
  INV_X1 U11252 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10667) );
  OR2_X1 U11253 ( .A1(n9407), .A2(n10667), .ZN(n9451) );
  NAND2_X1 U11254 ( .A1(n9447), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9448) );
  AND2_X1 U11255 ( .A1(n9463), .A2(n9448), .ZN(n11745) );
  OR2_X1 U11256 ( .A1(n9605), .A2(n11745), .ZN(n9450) );
  INV_X1 U11257 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10652) );
  OR2_X1 U11258 ( .A1(n13246), .A2(n10652), .ZN(n9449) );
  NAND4_X1 U11259 ( .A1(n9452), .A2(n9451), .A3(n9450), .A4(n9449), .ZN(n13519) );
  INV_X1 U11260 ( .A(SI_6_), .ZN(n13566) );
  OR2_X1 U11261 ( .A1(n9443), .A2(n13566), .ZN(n9461) );
  XNOR2_X1 U11262 ( .A(n10224), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n9453) );
  XNOR2_X1 U11263 ( .A(n9454), .B(n9453), .ZN(n10175) );
  OR2_X1 U11264 ( .A1(n9705), .A2(n10175), .ZN(n9460) );
  NAND2_X1 U11265 ( .A1(n9456), .A2(n9455), .ZN(n9469) );
  NAND2_X1 U11266 ( .A1(n9469), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9458) );
  XNOR2_X1 U11267 ( .A(n9457), .B(n9458), .ZN(n13769) );
  OR2_X1 U11268 ( .A1(n10431), .A2(n13769), .ZN(n9459) );
  OR2_X1 U11269 ( .A1(n13519), .A2(n11746), .ZN(n13121) );
  NAND2_X1 U11270 ( .A1(n13519), .A2(n11746), .ZN(n13122) );
  NAND2_X1 U11271 ( .A1(n13121), .A2(n13122), .ZN(n13260) );
  INV_X1 U11272 ( .A(n11746), .ZN(n11657) );
  NAND2_X1 U11273 ( .A1(n13519), .A2(n11657), .ZN(n9462) );
  NAND2_X1 U11274 ( .A1(n13244), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9468) );
  INV_X1 U11275 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10658) );
  OR2_X1 U11276 ( .A1(n9407), .A2(n10658), .ZN(n9467) );
  NAND2_X1 U11277 ( .A1(n9463), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9464) );
  AND2_X1 U11278 ( .A1(n9478), .A2(n9464), .ZN(n16106) );
  OR2_X1 U11279 ( .A1(n9605), .A2(n16106), .ZN(n9466) );
  INV_X1 U11280 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10659) );
  OR2_X1 U11281 ( .A1(n13246), .A2(n10659), .ZN(n9465) );
  NAND4_X1 U11282 ( .A1(n9468), .A2(n9467), .A3(n9466), .A4(n9465), .ZN(n13518) );
  OAI21_X1 U11283 ( .B1(n9469), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9470) );
  XNOR2_X1 U11284 ( .A(n9470), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10803) );
  NAND2_X1 U11285 ( .A1(n9472), .A2(n9471), .ZN(n9473) );
  AND2_X1 U11286 ( .A1(n9474), .A2(n9473), .ZN(n10168) );
  OR2_X1 U11287 ( .A1(n9443), .A2(SI_7_), .ZN(n9475) );
  OAI211_X1 U11288 ( .C1(n10803), .C2(n10431), .A(n9476), .B(n9475), .ZN(
        n16108) );
  OR2_X1 U11289 ( .A1(n13518), .A2(n16108), .ZN(n13126) );
  NAND2_X1 U11290 ( .A1(n13518), .A2(n16108), .ZN(n13127) );
  NAND2_X1 U11291 ( .A1(n13126), .A2(n13127), .ZN(n13259) );
  INV_X1 U11292 ( .A(n16108), .ZN(n11798) );
  NAND2_X1 U11293 ( .A1(n13518), .A2(n11798), .ZN(n9477) );
  NAND2_X1 U11294 ( .A1(n13244), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9483) );
  INV_X1 U11295 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10798) );
  OR2_X1 U11296 ( .A1(n9407), .A2(n10798), .ZN(n9482) );
  NAND2_X1 U11297 ( .A1(n9478), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9479) );
  AND2_X1 U11298 ( .A1(n9495), .A2(n9479), .ZN(n16127) );
  OR2_X1 U11299 ( .A1(n9605), .A2(n16127), .ZN(n9481) );
  INV_X1 U11300 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10806) );
  OR2_X1 U11301 ( .A1(n13246), .A2(n10806), .ZN(n9480) );
  NAND4_X1 U11302 ( .A1(n9483), .A2(n9482), .A3(n9481), .A4(n9480), .ZN(n13517) );
  INV_X1 U11303 ( .A(n9485), .ZN(n9487) );
  NAND2_X1 U11304 ( .A1(n9484), .A2(n9486), .ZN(n9506) );
  NAND2_X1 U11305 ( .A1(n9487), .A2(n9506), .ZN(n11016) );
  OR2_X1 U11306 ( .A1(n9489), .A2(n9488), .ZN(n9490) );
  NAND2_X1 U11307 ( .A1(n9491), .A2(n9490), .ZN(n10167) );
  INV_X1 U11308 ( .A(SI_8_), .ZN(n13671) );
  OR2_X1 U11309 ( .A1(n9443), .A2(n13671), .ZN(n9492) );
  OAI211_X1 U11310 ( .C1(n10431), .C2(n11016), .A(n9493), .B(n9492), .ZN(
        n13130) );
  XNOR2_X1 U11311 ( .A(n13517), .B(n13130), .ZN(n13257) );
  OR2_X1 U11312 ( .A1(n13517), .A2(n13130), .ZN(n9494) );
  NAND2_X1 U11313 ( .A1(n13244), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9500) );
  OR2_X1 U11314 ( .A1(n9407), .A2(n16146), .ZN(n9499) );
  NAND2_X1 U11315 ( .A1(n9495), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9496) );
  AND2_X1 U11316 ( .A1(n9512), .A2(n9496), .ZN(n12159) );
  OR2_X1 U11317 ( .A1(n9605), .A2(n12159), .ZN(n9498) );
  INV_X1 U11318 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11007) );
  OR2_X1 U11319 ( .A1(n13246), .A2(n11007), .ZN(n9497) );
  NAND4_X1 U11320 ( .A1(n9500), .A2(n9499), .A3(n9498), .A4(n9497), .ZN(n13516) );
  OR2_X1 U11321 ( .A1(n9502), .A2(n9501), .ZN(n9503) );
  AND2_X1 U11322 ( .A1(n9504), .A2(n9503), .ZN(n10180) );
  OR2_X1 U11323 ( .A1(n9443), .A2(SI_9_), .ZN(n9509) );
  NAND2_X1 U11324 ( .A1(n9506), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9505) );
  MUX2_X1 U11325 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9505), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n9507) );
  NAND2_X1 U11326 ( .A1(n9507), .A2(n9617), .ZN(n11019) );
  INV_X1 U11327 ( .A(n11019), .ZN(n11575) );
  OR2_X1 U11328 ( .A1(n10431), .A2(n11575), .ZN(n9508) );
  NOR2_X1 U11329 ( .A1(n13516), .A2(n12119), .ZN(n9510) );
  INV_X1 U11330 ( .A(n13516), .ZN(n12238) );
  NAND2_X1 U11331 ( .A1(n9796), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9517) );
  INV_X1 U11332 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n9511) );
  OR2_X1 U11333 ( .A1(n9799), .A2(n9511), .ZN(n9516) );
  NAND2_X1 U11334 ( .A1(n9512), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9513) );
  AND2_X1 U11335 ( .A1(n9535), .A2(n9513), .ZN(n12256) );
  OR2_X1 U11336 ( .A1(n9605), .A2(n12256), .ZN(n9515) );
  INV_X1 U11337 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12257) );
  OR2_X1 U11338 ( .A1(n13246), .A2(n12257), .ZN(n9514) );
  NAND4_X1 U11339 ( .A1(n9517), .A2(n9516), .A3(n9515), .A4(n9514), .ZN(n13515) );
  OR2_X1 U11340 ( .A1(n9519), .A2(n9518), .ZN(n9520) );
  NAND2_X1 U11341 ( .A1(n9521), .A2(n9520), .ZN(n10182) );
  NAND2_X1 U11342 ( .A1(n10182), .A2(n13241), .ZN(n9524) );
  NAND2_X1 U11343 ( .A1(n9617), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9522) );
  XNOR2_X1 U11344 ( .A(n9522), .B(P3_IR_REG_10__SCAN_IN), .ZN(n11953) );
  OR2_X1 U11345 ( .A1(n10431), .A2(n11953), .ZN(n9523) );
  OAI211_X1 U11346 ( .C1(n9730), .C2(SI_10_), .A(n9524), .B(n9523), .ZN(n16162) );
  OR2_X1 U11347 ( .A1(n13515), .A2(n16162), .ZN(n13140) );
  NAND2_X1 U11348 ( .A1(n13515), .A2(n16162), .ZN(n13141) );
  NAND2_X1 U11349 ( .A1(n13140), .A2(n13141), .ZN(n13268) );
  INV_X1 U11350 ( .A(n16162), .ZN(n12259) );
  NAND2_X1 U11351 ( .A1(n13515), .A2(n12259), .ZN(n9525) );
  OR2_X1 U11352 ( .A1(n9527), .A2(n9526), .ZN(n9528) );
  NAND2_X1 U11353 ( .A1(n9529), .A2(n9528), .ZN(n10189) );
  NAND2_X1 U11354 ( .A1(n10189), .A2(n13241), .ZN(n9532) );
  NOR2_X1 U11355 ( .A1(n9617), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n9546) );
  XNOR2_X1 U11356 ( .A(n9530), .B(n9545), .ZN(n11965) );
  AOI22_X1 U11357 ( .A1(n9668), .A2(n13666), .B1(n9667), .B2(n11965), .ZN(
        n9531) );
  NAND2_X1 U11358 ( .A1(n13244), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9540) );
  INV_X1 U11359 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n9533) );
  OR2_X1 U11360 ( .A1(n9407), .A2(n9533), .ZN(n9539) );
  INV_X1 U11361 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n9534) );
  OR2_X1 U11362 ( .A1(n13246), .A2(n9534), .ZN(n9538) );
  NAND2_X1 U11363 ( .A1(n9535), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9536) );
  AND2_X1 U11364 ( .A1(n9555), .A2(n9536), .ZN(n12435) );
  OR2_X1 U11365 ( .A1(n9605), .A2(n12435), .ZN(n9537) );
  NAND4_X1 U11366 ( .A1(n9540), .A2(n9539), .A3(n9538), .A4(n9537), .ZN(n13514) );
  AND2_X1 U11367 ( .A1(n12366), .A2(n13514), .ZN(n12357) );
  OR2_X1 U11368 ( .A1(n12366), .A2(n13514), .ZN(n12358) );
  OR2_X1 U11369 ( .A1(n9542), .A2(n9541), .ZN(n9543) );
  NAND2_X1 U11370 ( .A1(n9544), .A2(n9543), .ZN(n10221) );
  INV_X1 U11371 ( .A(n9547), .ZN(n9551) );
  INV_X1 U11372 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9548) );
  INV_X1 U11373 ( .A(n9567), .ZN(n9550) );
  INV_X1 U11374 ( .A(n12306), .ZN(n9552) );
  AOI22_X1 U11375 ( .A1(n9668), .A2(SI_12_), .B1(n9667), .B2(n9552), .ZN(n9553) );
  NAND2_X1 U11376 ( .A1(n9554), .A2(n9553), .ZN(n14187) );
  NAND2_X1 U11377 ( .A1(n13244), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9560) );
  INV_X1 U11378 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14190) );
  OR2_X1 U11379 ( .A1(n9407), .A2(n14190), .ZN(n9559) );
  NAND2_X1 U11380 ( .A1(n9555), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9556) );
  AND2_X1 U11381 ( .A1(n9572), .A2(n9556), .ZN(n12560) );
  OR2_X1 U11382 ( .A1(n9605), .A2(n12560), .ZN(n9558) );
  INV_X1 U11383 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12484) );
  OR2_X1 U11384 ( .A1(n13246), .A2(n12484), .ZN(n9557) );
  NAND4_X1 U11385 ( .A1(n9560), .A2(n9559), .A3(n9558), .A4(n9557), .ZN(n13513) );
  NAND2_X1 U11386 ( .A1(n14187), .A2(n13513), .ZN(n12551) );
  OR2_X1 U11387 ( .A1(n14187), .A2(n13513), .ZN(n12552) );
  NAND2_X1 U11388 ( .A1(n9562), .A2(n10679), .ZN(n9563) );
  NAND2_X1 U11389 ( .A1(n9564), .A2(n9563), .ZN(n10341) );
  NAND2_X1 U11390 ( .A1(n10341), .A2(n13241), .ZN(n9570) );
  INV_X1 U11391 ( .A(SI_13_), .ZN(n10342) );
  INV_X1 U11392 ( .A(n9565), .ZN(n9568) );
  INV_X1 U11393 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U11394 ( .A1(n9567), .A2(n9566), .ZN(n9598) );
  NAND2_X1 U11395 ( .A1(n9568), .A2(n9598), .ZN(n12311) );
  AOI22_X1 U11396 ( .A1(n9668), .A2(n10342), .B1(n9667), .B2(n12311), .ZN(
        n9569) );
  NAND2_X1 U11397 ( .A1(n9570), .A2(n9569), .ZN(n16217) );
  NAND2_X1 U11398 ( .A1(n13244), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9577) );
  INV_X1 U11399 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n9571) );
  OR2_X1 U11400 ( .A1(n9407), .A2(n9571), .ZN(n9576) );
  NAND2_X1 U11401 ( .A1(n9572), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9573) );
  AND2_X1 U11402 ( .A1(n9588), .A2(n9573), .ZN(n12641) );
  OR2_X1 U11403 ( .A1(n9605), .A2(n12641), .ZN(n9575) );
  INV_X1 U11404 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12642) );
  OR2_X1 U11405 ( .A1(n13246), .A2(n12642), .ZN(n9574) );
  AND2_X1 U11406 ( .A1(n16217), .A2(n13384), .ZN(n9578) );
  OR2_X1 U11407 ( .A1(n16217), .A2(n13384), .ZN(n13332) );
  OR2_X1 U11408 ( .A1(n9580), .A2(n9579), .ZN(n9581) );
  NAND2_X1 U11409 ( .A1(n9582), .A2(n9581), .ZN(n10361) );
  NAND2_X1 U11410 ( .A1(n10361), .A2(n13241), .ZN(n9586) );
  NAND2_X1 U11411 ( .A1(n9598), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9584) );
  XNOR2_X1 U11412 ( .A(n9584), .B(n9583), .ZN(n13797) );
  AOI22_X1 U11413 ( .A1(n9668), .A2(n13624), .B1(n9667), .B2(n13797), .ZN(
        n9585) );
  NAND2_X1 U11414 ( .A1(n13244), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9593) );
  INV_X1 U11415 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n9587) );
  OR2_X1 U11416 ( .A1(n9407), .A2(n9587), .ZN(n9592) );
  NAND2_X1 U11417 ( .A1(n9588), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9589) );
  AND2_X1 U11418 ( .A1(n9603), .A2(n9589), .ZN(n14112) );
  OR2_X1 U11419 ( .A1(n9605), .A2(n14112), .ZN(n9591) );
  INV_X1 U11420 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n14113) );
  OR2_X1 U11421 ( .A1(n13246), .A2(n14113), .ZN(n9590) );
  NAND4_X1 U11422 ( .A1(n9593), .A2(n9592), .A3(n9591), .A4(n9590), .ZN(n14089) );
  NAND2_X1 U11423 ( .A1(n16223), .A2(n14089), .ZN(n13155) );
  NAND2_X1 U11424 ( .A1(n13157), .A2(n13155), .ZN(n14105) );
  INV_X1 U11425 ( .A(n14089), .ZN(n13501) );
  OR2_X1 U11426 ( .A1(n16223), .A2(n13501), .ZN(n14086) );
  OR2_X1 U11427 ( .A1(n9595), .A2(n9594), .ZN(n9596) );
  NAND2_X1 U11428 ( .A1(n9597), .A2(n9596), .ZN(n10362) );
  NAND2_X1 U11429 ( .A1(n10362), .A2(n13241), .ZN(n9602) );
  OAI21_X1 U11430 ( .B1(n9598), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9600) );
  INV_X1 U11431 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9599) );
  XNOR2_X1 U11432 ( .A(n9600), .B(n9599), .ZN(n13801) );
  AOI22_X1 U11433 ( .A1(n9668), .A2(n13659), .B1(n9667), .B2(n13801), .ZN(
        n9601) );
  NAND2_X1 U11434 ( .A1(n13244), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9609) );
  INV_X1 U11435 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14185) );
  OR2_X1 U11436 ( .A1(n9407), .A2(n14185), .ZN(n9608) );
  NAND2_X1 U11437 ( .A1(n9603), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9604) );
  AND2_X1 U11438 ( .A1(n9621), .A2(n9604), .ZN(n14095) );
  OR2_X1 U11439 ( .A1(n9605), .A2(n14095), .ZN(n9607) );
  INV_X1 U11440 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14096) );
  OR2_X1 U11441 ( .A1(n13246), .A2(n14096), .ZN(n9606) );
  NAND4_X1 U11442 ( .A1(n9609), .A2(n9608), .A3(n9607), .A4(n9606), .ZN(n14106) );
  NAND2_X1 U11443 ( .A1(n14242), .A2(n14106), .ZN(n13166) );
  NAND2_X1 U11444 ( .A1(n13164), .A2(n13166), .ZN(n13277) );
  NAND2_X1 U11445 ( .A1(n9610), .A2(n13277), .ZN(n14084) );
  INV_X1 U11446 ( .A(n14106), .ZN(n14076) );
  OR2_X1 U11447 ( .A1(n14242), .A2(n14076), .ZN(n9611) );
  OR2_X1 U11448 ( .A1(n9613), .A2(n9612), .ZN(n9614) );
  NAND2_X1 U11449 ( .A1(n9615), .A2(n9614), .ZN(n10429) );
  OAI21_X1 U11450 ( .B1(n9617), .B2(n9616), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n9618) );
  XNOR2_X1 U11451 ( .A(n9618), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13823) );
  AOI22_X1 U11452 ( .A1(n9668), .A2(SI_16_), .B1(n9667), .B2(n13823), .ZN(
        n9619) );
  NAND2_X1 U11453 ( .A1(n9621), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U11454 ( .A1(n9638), .A2(n9622), .ZN(n14078) );
  NAND2_X1 U11455 ( .A1(n9778), .A2(n14078), .ZN(n9627) );
  INV_X1 U11456 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n9623) );
  OR2_X1 U11457 ( .A1(n9799), .A2(n9623), .ZN(n9626) );
  INV_X1 U11458 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13812) );
  OR2_X1 U11459 ( .A1(n9407), .A2(n13812), .ZN(n9625) );
  INV_X1 U11460 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13822) );
  OR2_X1 U11461 ( .A1(n13246), .A2(n13822), .ZN(n9624) );
  NAND4_X1 U11462 ( .A1(n9627), .A2(n9626), .A3(n9625), .A4(n9624), .ZN(n14088) );
  NAND2_X1 U11463 ( .A1(n14179), .A2(n14088), .ZN(n13163) );
  NAND2_X1 U11464 ( .A1(n13171), .A2(n13163), .ZN(n14074) );
  OR2_X1 U11465 ( .A1(n9629), .A2(n9628), .ZN(n9630) );
  NAND2_X1 U11466 ( .A1(n9631), .A2(n9630), .ZN(n10483) );
  NAND2_X1 U11467 ( .A1(n10483), .A2(n13241), .ZN(n9637) );
  INV_X1 U11468 ( .A(SI_17_), .ZN(n13627) );
  NAND2_X1 U11469 ( .A1(n9632), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9633) );
  MUX2_X1 U11470 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9633), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9635) );
  NAND2_X1 U11471 ( .A1(n9635), .A2(n9634), .ZN(n13868) );
  AOI22_X1 U11472 ( .A1(n9668), .A2(n13627), .B1(n9667), .B2(n13868), .ZN(
        n9636) );
  NAND2_X1 U11473 ( .A1(n9638), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U11474 ( .A1(n9653), .A2(n9639), .ZN(n14061) );
  NAND2_X1 U11475 ( .A1(n9778), .A2(n14061), .ZN(n9644) );
  INV_X1 U11476 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13834) );
  OR2_X1 U11477 ( .A1(n9407), .A2(n13834), .ZN(n9643) );
  INV_X1 U11478 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14063) );
  OR2_X1 U11479 ( .A1(n13246), .A2(n14063), .ZN(n9642) );
  INV_X1 U11480 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n9640) );
  OR2_X1 U11481 ( .A1(n9799), .A2(n9640), .ZN(n9641) );
  NAND4_X1 U11482 ( .A1(n9644), .A2(n9643), .A3(n9642), .A4(n9641), .ZN(n14049) );
  XNOR2_X1 U11483 ( .A(n14237), .B(n14049), .ZN(n14056) );
  INV_X1 U11484 ( .A(n14049), .ZN(n14077) );
  OR2_X1 U11485 ( .A1(n14237), .A2(n14077), .ZN(n9645) );
  OR2_X1 U11486 ( .A1(n9647), .A2(n9646), .ZN(n9648) );
  NAND2_X1 U11487 ( .A1(n9649), .A2(n9648), .ZN(n10609) );
  NAND2_X1 U11488 ( .A1(n9634), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9650) );
  XNOR2_X1 U11489 ( .A(n9650), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U11490 ( .A1(n9668), .A2(SI_18_), .B1(n9667), .B2(n13884), .ZN(
        n9651) );
  NAND2_X1 U11491 ( .A1(n9653), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9654) );
  NAND2_X1 U11492 ( .A1(n9671), .A2(n9654), .ZN(n14043) );
  NAND2_X1 U11493 ( .A1(n14043), .A2(n9778), .ZN(n9659) );
  INV_X1 U11494 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13860) );
  OR2_X1 U11495 ( .A1(n9407), .A2(n13860), .ZN(n9658) );
  INV_X1 U11496 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n9655) );
  OR2_X1 U11497 ( .A1(n9799), .A2(n9655), .ZN(n9657) );
  INV_X1 U11498 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n14045) );
  OR2_X1 U11499 ( .A1(n13246), .A2(n14045), .ZN(n9656) );
  NAND2_X1 U11500 ( .A1(n14169), .A2(n14028), .ZN(n13175) );
  NAND2_X1 U11501 ( .A1(n13177), .A2(n13175), .ZN(n14047) );
  OR2_X1 U11502 ( .A1(n14169), .A2(n14058), .ZN(n9660) );
  NAND2_X1 U11503 ( .A1(n14046), .A2(n9660), .ZN(n14026) );
  OR2_X1 U11504 ( .A1(n9662), .A2(n9661), .ZN(n9663) );
  NAND2_X1 U11505 ( .A1(n9664), .A2(n9663), .ZN(n10648) );
  INV_X1 U11506 ( .A(n9786), .ZN(n9665) );
  NAND2_X1 U11507 ( .A1(n9665), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9666) );
  AOI22_X1 U11508 ( .A1(n9668), .A2(SI_19_), .B1(n13881), .B2(n9667), .ZN(
        n9669) );
  INV_X1 U11509 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n14031) );
  NAND2_X1 U11510 ( .A1(n9671), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U11511 ( .A1(n9682), .A2(n9672), .ZN(n14030) );
  NAND2_X1 U11512 ( .A1(n14030), .A2(n9778), .ZN(n9674) );
  AOI22_X1 U11513 ( .A1(n13244), .A2(P3_REG0_REG_19__SCAN_IN), .B1(n9796), 
        .B2(P3_REG1_REG_19__SCAN_IN), .ZN(n9673) );
  OAI211_X1 U11514 ( .C1(n13246), .C2(n14031), .A(n9674), .B(n9673), .ZN(
        n14050) );
  NAND2_X1 U11515 ( .A1(n14039), .A2(n14050), .ZN(n9675) );
  OR2_X1 U11516 ( .A1(n9677), .A2(n9676), .ZN(n9678) );
  NAND2_X1 U11517 ( .A1(n9679), .A2(n9678), .ZN(n10777) );
  OR2_X1 U11518 ( .A1(n9730), .A2(n10776), .ZN(n9680) );
  NAND2_X1 U11519 ( .A1(n9682), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U11520 ( .A1(n9693), .A2(n9683), .ZN(n14020) );
  NAND2_X1 U11521 ( .A1(n14020), .A2(n9778), .ZN(n9686) );
  AOI22_X1 U11522 ( .A1(n13244), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n9796), 
        .B2(P3_REG1_REG_20__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U11523 ( .A1(n9795), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U11524 ( .A1(n14227), .A2(n14029), .ZN(n13190) );
  NAND2_X1 U11525 ( .A1(n13189), .A2(n13190), .ZN(n13281) );
  OR2_X1 U11526 ( .A1(n9688), .A2(n9687), .ZN(n9689) );
  NAND2_X1 U11527 ( .A1(n9690), .A2(n9689), .ZN(n10958) );
  INV_X1 U11528 ( .A(SI_21_), .ZN(n10957) );
  OR2_X1 U11529 ( .A1(n9730), .A2(n10957), .ZN(n9691) );
  NAND2_X1 U11530 ( .A1(n9693), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U11531 ( .A1(n9708), .A2(n9694), .ZN(n14005) );
  NAND2_X1 U11532 ( .A1(n14005), .A2(n9778), .ZN(n9700) );
  INV_X1 U11533 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n9697) );
  NAND2_X1 U11534 ( .A1(n9796), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U11535 ( .A1(n9795), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9695) );
  OAI211_X1 U11536 ( .C1(n9697), .C2(n9799), .A(n9696), .B(n9695), .ZN(n9698)
         );
  INV_X1 U11537 ( .A(n9698), .ZN(n9699) );
  OR2_X1 U11538 ( .A1(n9702), .A2(n9701), .ZN(n9703) );
  NAND2_X1 U11539 ( .A1(n9704), .A2(n9703), .ZN(n11042) );
  OR2_X1 U11540 ( .A1(n9730), .A2(n13652), .ZN(n9706) );
  NAND2_X1 U11541 ( .A1(n9708), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U11542 ( .A1(n9722), .A2(n9709), .ZN(n13994) );
  NAND2_X1 U11543 ( .A1(n13994), .A2(n9778), .ZN(n9715) );
  INV_X1 U11544 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n9712) );
  NAND2_X1 U11545 ( .A1(n9796), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9711) );
  NAND2_X1 U11546 ( .A1(n9795), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9710) );
  OAI211_X1 U11547 ( .C1(n9712), .C2(n9799), .A(n9711), .B(n9710), .ZN(n9713)
         );
  INV_X1 U11548 ( .A(n9713), .ZN(n9714) );
  INV_X1 U11549 ( .A(n14151), .ZN(n13475) );
  XNOR2_X1 U11550 ( .A(n9719), .B(n9718), .ZN(n11295) );
  NAND2_X1 U11551 ( .A1(n11295), .A2(n13241), .ZN(n9721) );
  NAND2_X1 U11552 ( .A1(n9722), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U11553 ( .A1(n9733), .A2(n9723), .ZN(n13982) );
  NAND2_X1 U11554 ( .A1(n13982), .A2(n9778), .ZN(n9728) );
  INV_X1 U11555 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n14220) );
  NAND2_X1 U11556 ( .A1(n9796), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U11557 ( .A1(n9795), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9724) );
  OAI211_X1 U11558 ( .C1(n14220), .C2(n9799), .A(n9725), .B(n9724), .ZN(n9726)
         );
  INV_X1 U11559 ( .A(n9726), .ZN(n9727) );
  XNOR2_X1 U11560 ( .A(n13392), .B(n13966), .ZN(n13974) );
  XNOR2_X1 U11561 ( .A(n9729), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U11562 ( .A1(n11729), .A2(n13241), .ZN(n9732) );
  INV_X1 U11563 ( .A(SI_24_), .ZN(n13646) );
  OR2_X1 U11564 ( .A1(n9443), .A2(n13646), .ZN(n9731) );
  NAND2_X1 U11565 ( .A1(n9733), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9734) );
  NAND2_X1 U11566 ( .A1(n9735), .A2(n9734), .ZN(n13967) );
  NAND2_X1 U11567 ( .A1(n13967), .A2(n9778), .ZN(n9740) );
  INV_X1 U11568 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n14216) );
  NAND2_X1 U11569 ( .A1(n9795), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9737) );
  NAND2_X1 U11570 ( .A1(n9796), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9736) );
  OAI211_X1 U11571 ( .C1(n9799), .C2(n14216), .A(n9737), .B(n9736), .ZN(n9738)
         );
  INV_X1 U11572 ( .A(n9738), .ZN(n9739) );
  NAND2_X1 U11573 ( .A1(n13963), .A2(n8473), .ZN(n9742) );
  NAND2_X1 U11574 ( .A1(n9742), .A2(n9741), .ZN(n13950) );
  XNOR2_X1 U11575 ( .A(n9744), .B(n9743), .ZN(n11970) );
  NAND2_X1 U11576 ( .A1(n11970), .A2(n13241), .ZN(n9746) );
  INV_X1 U11577 ( .A(SI_26_), .ZN(n13640) );
  NAND2_X1 U11578 ( .A1(n9747), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U11579 ( .A1(n9749), .A2(n9748), .ZN(n13944) );
  INV_X1 U11580 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n14208) );
  NAND2_X1 U11581 ( .A1(n9795), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9751) );
  NAND2_X1 U11582 ( .A1(n9796), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9750) );
  OAI211_X1 U11583 ( .C1(n9799), .C2(n14208), .A(n9751), .B(n9750), .ZN(n9752)
         );
  INV_X1 U11584 ( .A(n9752), .ZN(n9753) );
  NOR2_X1 U11585 ( .A1(n13369), .A2(n13510), .ZN(n9754) );
  NAND2_X1 U11586 ( .A1(n13329), .A2(n13943), .ZN(n13210) );
  INV_X1 U11587 ( .A(n9755), .ZN(n9756) );
  NAND2_X1 U11588 ( .A1(n9757), .A2(n9756), .ZN(n9759) );
  NAND2_X1 U11589 ( .A1(n13081), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9774) );
  NAND2_X1 U11590 ( .A1(n9760), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U11591 ( .A1(n9774), .A2(n9761), .ZN(n9771) );
  XNOR2_X1 U11592 ( .A(n9773), .B(n9771), .ZN(n12262) );
  NAND2_X1 U11593 ( .A1(n12262), .A2(n13241), .ZN(n9763) );
  NAND2_X1 U11594 ( .A1(n9764), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9765) );
  NAND2_X1 U11595 ( .A1(n13903), .A2(n9765), .ZN(n13923) );
  INV_X1 U11596 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n14201) );
  NAND2_X1 U11597 ( .A1(n9795), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U11598 ( .A1(n9796), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9766) );
  OAI211_X1 U11599 ( .C1(n9799), .C2(n14201), .A(n9767), .B(n9766), .ZN(n9768)
         );
  NAND2_X1 U11600 ( .A1(n13412), .A2(n13932), .ZN(n13218) );
  NAND2_X1 U11601 ( .A1(n13916), .A2(n13915), .ZN(n13918) );
  NAND2_X1 U11602 ( .A1(n13918), .A2(n9770), .ZN(n9784) );
  INV_X1 U11603 ( .A(n9771), .ZN(n9772) );
  NAND2_X1 U11604 ( .A1(n9773), .A2(n9772), .ZN(n9775) );
  NAND2_X1 U11605 ( .A1(n9775), .A2(n9774), .ZN(n13221) );
  XNOR2_X1 U11606 ( .A(n14959), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n13219) );
  XNOR2_X1 U11607 ( .A(n13221), .B(n13219), .ZN(n12393) );
  NAND2_X1 U11608 ( .A1(n12393), .A2(n13241), .ZN(n9777) );
  INV_X1 U11609 ( .A(SI_29_), .ZN(n12394) );
  OR2_X1 U11610 ( .A1(n9730), .A2(n12394), .ZN(n9776) );
  NAND2_X1 U11611 ( .A1(n9777), .A2(n9776), .ZN(n9861) );
  INV_X1 U11612 ( .A(n13903), .ZN(n9779) );
  NAND2_X1 U11613 ( .A1(n9779), .A2(n9778), .ZN(n13251) );
  INV_X1 U11614 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U11615 ( .A1(n13244), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U11616 ( .A1(n9795), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9780) );
  OAI211_X1 U11617 ( .C1(n9878), .C2(n9407), .A(n9781), .B(n9780), .ZN(n9782)
         );
  INV_X1 U11618 ( .A(n9782), .ZN(n9783) );
  OR2_X1 U11619 ( .A1(n9861), .A2(n13919), .ZN(n13295) );
  NAND2_X1 U11620 ( .A1(n9861), .A2(n13919), .ZN(n13297) );
  NAND2_X1 U11621 ( .A1(n13295), .A2(n13297), .ZN(n13286) );
  XNOR2_X1 U11622 ( .A(n9784), .B(n13286), .ZN(n9805) );
  NAND2_X1 U11623 ( .A1(n7234), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U11624 ( .A1(n13313), .A2(n13881), .ZN(n9852) );
  NAND2_X1 U11625 ( .A1(n9788), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U11626 ( .A1(n9792), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U11627 ( .A1(n13102), .A2(n9851), .ZN(n13304) );
  INV_X1 U11628 ( .A(n12264), .ZN(n13310) );
  NAND2_X1 U11629 ( .A1(n13310), .A2(n10438), .ZN(n10435) );
  NAND2_X1 U11630 ( .A1(n10435), .A2(n10431), .ZN(n10601) );
  INV_X1 U11631 ( .A(n10601), .ZN(n10461) );
  INV_X1 U11632 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14199) );
  NAND2_X1 U11633 ( .A1(n9795), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U11634 ( .A1(n9796), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9797) );
  OAI211_X1 U11635 ( .C1(n9799), .C2(n14199), .A(n9798), .B(n9797), .ZN(n9800)
         );
  INV_X1 U11636 ( .A(n9800), .ZN(n9801) );
  NAND2_X1 U11637 ( .A1(n13251), .A2(n9801), .ZN(n13509) );
  INV_X1 U11638 ( .A(P3_B_REG_SCAN_IN), .ZN(n9802) );
  NOR2_X1 U11639 ( .A1(n12264), .A2(n9802), .ZN(n9803) );
  NOR2_X1 U11640 ( .A1(n16032), .A2(n9803), .ZN(n13900) );
  AOI22_X1 U11641 ( .A1(n14108), .A2(n9769), .B1(n13509), .B2(n13900), .ZN(
        n9804) );
  OR2_X1 U11642 ( .A1(n13523), .A2(n16029), .ZN(n9806) );
  OR2_X1 U11643 ( .A1(n13521), .A2(n13111), .ZN(n9808) );
  NAND2_X1 U11644 ( .A1(n11478), .A2(n13113), .ZN(n11477) );
  INV_X1 U11645 ( .A(n13260), .ZN(n13119) );
  NAND2_X1 U11646 ( .A1(n11466), .A2(n13119), .ZN(n11465) );
  INV_X1 U11647 ( .A(n13259), .ZN(n13124) );
  INV_X1 U11648 ( .A(n13130), .ZN(n16125) );
  OR2_X1 U11649 ( .A1(n13517), .A2(n16125), .ZN(n9809) );
  NOR2_X1 U11650 ( .A1(n13516), .A2(n16142), .ZN(n13136) );
  NAND2_X1 U11651 ( .A1(n13516), .A2(n16142), .ZN(n13137) );
  NAND2_X1 U11652 ( .A1(n13514), .A2(n16193), .ZN(n13145) );
  NAND2_X1 U11653 ( .A1(n12434), .A2(n13273), .ZN(n12433) );
  INV_X1 U11654 ( .A(n13513), .ZN(n12432) );
  OR2_X1 U11655 ( .A1(n14187), .A2(n12432), .ZN(n13148) );
  NAND2_X1 U11656 ( .A1(n14187), .A2(n12432), .ZN(n13149) );
  NAND2_X1 U11657 ( .A1(n12479), .A2(n13272), .ZN(n9811) );
  NAND2_X1 U11658 ( .A1(n9811), .A2(n13149), .ZN(n12633) );
  NAND2_X1 U11659 ( .A1(n16217), .A2(n14109), .ZN(n13331) );
  NAND2_X1 U11660 ( .A1(n12633), .A2(n13275), .ZN(n12635) );
  NAND2_X1 U11661 ( .A1(n12635), .A2(n13156), .ZN(n14102) );
  INV_X1 U11662 ( .A(n13277), .ZN(n14093) );
  INV_X1 U11663 ( .A(n14088), .ZN(n13445) );
  INV_X1 U11664 ( .A(n14056), .ZN(n14068) );
  NAND2_X1 U11665 ( .A1(n14067), .A2(n14068), .ZN(n9812) );
  OR2_X1 U11666 ( .A1(n14237), .A2(n14049), .ZN(n13173) );
  INV_X1 U11667 ( .A(n14047), .ZN(n13279) );
  INV_X1 U11668 ( .A(n14050), .ZN(n13462) );
  NAND2_X1 U11669 ( .A1(n14039), .A2(n13462), .ZN(n13183) );
  NAND2_X1 U11670 ( .A1(n13184), .A2(n13183), .ZN(n14034) );
  NAND2_X1 U11671 ( .A1(n14033), .A2(n13184), .ZN(n14012) );
  NAND2_X1 U11672 ( .A1(n14012), .A2(n14011), .ZN(n14014) );
  NAND2_X1 U11673 ( .A1(n14155), .A2(n13469), .ZN(n13355) );
  NAND2_X1 U11674 ( .A1(n13352), .A2(n13355), .ZN(n13999) );
  XNOR2_X1 U11675 ( .A(n14151), .B(n13977), .ZN(n13990) );
  NAND2_X1 U11676 ( .A1(n13475), .A2(n14002), .ZN(n13194) );
  NAND2_X1 U11677 ( .A1(n14222), .A2(n13988), .ZN(n13200) );
  NAND2_X1 U11678 ( .A1(n13968), .A2(n13978), .ZN(n13283) );
  NOR2_X1 U11679 ( .A1(n13968), .A2(n13978), .ZN(n13961) );
  INV_X1 U11680 ( .A(n13952), .ZN(n13093) );
  INV_X1 U11681 ( .A(n13915), .ZN(n13406) );
  XNOR2_X1 U11682 ( .A(n13296), .B(n13286), .ZN(n13913) );
  AND2_X1 U11683 ( .A1(n10956), .A2(n10775), .ZN(n9874) );
  INV_X1 U11684 ( .A(n9874), .ZN(n9815) );
  XNOR2_X1 U11685 ( .A(n13313), .B(n9815), .ZN(n9817) );
  NAND2_X1 U11686 ( .A1(n10956), .A2(n13888), .ZN(n9816) );
  NAND2_X1 U11687 ( .A1(n9817), .A2(n9816), .ZN(n10454) );
  INV_X1 U11688 ( .A(n13313), .ZN(n9820) );
  NAND2_X1 U11689 ( .A1(n10775), .A2(n13888), .ZN(n9869) );
  INV_X1 U11690 ( .A(n9869), .ZN(n13308) );
  AND2_X1 U11691 ( .A1(n16222), .A2(n13308), .ZN(n9818) );
  NAND2_X1 U11692 ( .A1(n10454), .A2(n9818), .ZN(n9819) );
  NAND2_X1 U11693 ( .A1(n9852), .A2(n9869), .ZN(n9871) );
  OR2_X1 U11694 ( .A1(n9871), .A2(n9820), .ZN(n9868) );
  AND2_X1 U11695 ( .A1(n9819), .A2(n9868), .ZN(n14017) );
  NAND2_X1 U11696 ( .A1(n9820), .A2(n16045), .ZN(n16163) );
  NAND2_X1 U11697 ( .A1(n9822), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9823) );
  XNOR2_X1 U11698 ( .A(n11731), .B(P3_B_REG_SCAN_IN), .ZN(n9830) );
  NAND2_X1 U11699 ( .A1(n9827), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9828) );
  MUX2_X1 U11700 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9828), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9829) );
  INV_X1 U11701 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9831) );
  NAND2_X1 U11702 ( .A1(n10244), .A2(n9831), .ZN(n9833) );
  INV_X1 U11703 ( .A(n9858), .ZN(n11972) );
  NAND2_X1 U11704 ( .A1(n11972), .A2(n11891), .ZN(n9832) );
  NOR2_X1 U11705 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9837) );
  NOR4_X1 U11706 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9836) );
  NOR4_X1 U11707 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9835) );
  NOR4_X1 U11708 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9834) );
  NAND4_X1 U11709 ( .A1(n9837), .A2(n9836), .A3(n9835), .A4(n9834), .ZN(n9843)
         );
  NOR4_X1 U11710 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9841) );
  NOR4_X1 U11711 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9840) );
  NOR4_X1 U11712 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9839) );
  NOR4_X1 U11713 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9838) );
  NAND4_X1 U11714 ( .A1(n9841), .A2(n9840), .A3(n9839), .A4(n9838), .ZN(n9842)
         );
  NOR2_X1 U11715 ( .A1(n9843), .A2(n9842), .ZN(n9844) );
  NOR2_X1 U11716 ( .A1(n9845), .A2(n9844), .ZN(n9864) );
  NOR2_X1 U11717 ( .A1(n14248), .A2(n9864), .ZN(n9849) );
  INV_X1 U11718 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9846) );
  NAND2_X1 U11719 ( .A1(n11972), .A2(n11731), .ZN(n9847) );
  NAND2_X1 U11720 ( .A1(n9849), .A2(n9865), .ZN(n10459) );
  INV_X1 U11721 ( .A(n10454), .ZN(n10450) );
  INV_X1 U11722 ( .A(n9864), .ZN(n9850) );
  OR2_X1 U11723 ( .A1(n13293), .A2(n9852), .ZN(n10455) );
  OR2_X1 U11724 ( .A1(n13217), .A2(n9869), .ZN(n10477) );
  NAND2_X1 U11725 ( .A1(n10455), .A2(n10477), .ZN(n9853) );
  NAND2_X1 U11726 ( .A1(n10464), .A2(n9853), .ZN(n9854) );
  OAI21_X1 U11727 ( .B1(n10459), .B2(n10450), .A(n9854), .ZN(n9859) );
  NOR2_X1 U11728 ( .A1(n11891), .A2(n11731), .ZN(n9857) );
  INV_X1 U11729 ( .A(n9861), .ZN(n13908) );
  NOR2_X1 U11730 ( .A1(n10462), .A2(n9864), .ZN(n9867) );
  XNOR2_X1 U11731 ( .A(n9865), .B(n14248), .ZN(n9866) );
  NAND2_X1 U11732 ( .A1(n9868), .A2(n13217), .ZN(n11059) );
  NAND2_X1 U11733 ( .A1(n13229), .A2(n9869), .ZN(n11055) );
  NAND2_X1 U11734 ( .A1(n11059), .A2(n11055), .ZN(n9870) );
  NAND2_X1 U11735 ( .A1(n9870), .A2(n14248), .ZN(n9876) );
  NAND2_X1 U11736 ( .A1(n9871), .A2(n10956), .ZN(n9873) );
  INV_X1 U11737 ( .A(n14248), .ZN(n9872) );
  OAI211_X1 U11738 ( .C1(n13313), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9875)
         );
  NAND2_X1 U11739 ( .A1(n7193), .A2(n10974), .ZN(n10116) );
  NAND2_X1 U11740 ( .A1(n9882), .A2(n10050), .ZN(n9885) );
  OAI21_X1 U11741 ( .B1(n9885), .B2(n11399), .A(n9881), .ZN(n9887) );
  NAND3_X1 U11742 ( .A1(n9885), .A2(n9884), .A3(n9883), .ZN(n9886) );
  NAND2_X1 U11743 ( .A1(n9887), .A2(n9886), .ZN(n9898) );
  NAND2_X1 U11744 ( .A1(n14484), .A2(n10055), .ZN(n9889) );
  NAND2_X1 U11745 ( .A1(n7718), .A2(n10050), .ZN(n9888) );
  NAND2_X1 U11746 ( .A1(n9889), .A2(n9888), .ZN(n9897) );
  INV_X1 U11747 ( .A(n9904), .ZN(n9894) );
  NAND2_X1 U11748 ( .A1(n14483), .A2(n10050), .ZN(n9893) );
  NAND2_X1 U11749 ( .A1(n11724), .A2(n10055), .ZN(n9892) );
  NAND2_X1 U11750 ( .A1(n9893), .A2(n9892), .ZN(n9903) );
  NAND2_X1 U11751 ( .A1(n9894), .A2(n9903), .ZN(n9895) );
  OAI21_X1 U11752 ( .B1(n9898), .B2(n9897), .A(n9895), .ZN(n9908) );
  AOI22_X1 U11753 ( .A1(n14484), .A2(n10050), .B1(n10055), .B2(n7718), .ZN(
        n9896) );
  AOI21_X1 U11754 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(n9907) );
  AND2_X1 U11755 ( .A1(n10055), .A2(n9900), .ZN(n9899) );
  AOI21_X1 U11756 ( .B1(n14482), .B2(n10057), .A(n9899), .ZN(n9909) );
  NAND2_X1 U11757 ( .A1(n14482), .A2(n10055), .ZN(n9902) );
  NAND2_X1 U11758 ( .A1(n10050), .A2(n9900), .ZN(n9901) );
  INV_X1 U11759 ( .A(n9903), .ZN(n9905) );
  OAI21_X1 U11760 ( .B1(n9908), .B2(n9907), .A(n9906), .ZN(n9913) );
  INV_X1 U11761 ( .A(n9909), .ZN(n9910) );
  NAND2_X1 U11762 ( .A1(n9911), .A2(n9910), .ZN(n9912) );
  NAND2_X1 U11763 ( .A1(n14481), .A2(n10050), .ZN(n9915) );
  NAND2_X1 U11764 ( .A1(n11603), .A2(n10055), .ZN(n9914) );
  NAND2_X1 U11765 ( .A1(n9915), .A2(n9914), .ZN(n9917) );
  BUF_X2 U11766 ( .A(n10050), .Z(n10057) );
  AOI22_X1 U11767 ( .A1(n14481), .A2(n10055), .B1(n11603), .B2(n10057), .ZN(
        n9916) );
  NAND2_X1 U11768 ( .A1(n14480), .A2(n10055), .ZN(n9921) );
  NAND2_X1 U11769 ( .A1(n10050), .A2(n11840), .ZN(n9920) );
  OAI22_X1 U11770 ( .A1(n9922), .A2(n10085), .B1(n11418), .B2(n7194), .ZN(
        n9923) );
  AOI22_X1 U11771 ( .A1(n10055), .A2(n11508), .B1(n14479), .B2(n10057), .ZN(
        n9926) );
  OAI22_X1 U11772 ( .A1(n9924), .A2(n7194), .B1(n12321), .B2(n10085), .ZN(
        n9925) );
  INV_X1 U11773 ( .A(n10057), .ZN(n10073) );
  OAI22_X1 U11774 ( .A1(n12295), .A2(n10073), .B1(n11679), .B2(n7194), .ZN(
        n9930) );
  NAND2_X1 U11775 ( .A1(n9928), .A2(n9927), .ZN(n9934) );
  INV_X1 U11776 ( .A(n9929), .ZN(n9932) );
  INV_X1 U11777 ( .A(n9930), .ZN(n9931) );
  NAND2_X1 U11778 ( .A1(n9932), .A2(n9931), .ZN(n9933) );
  OAI22_X1 U11779 ( .A1(n11901), .A2(n7194), .B1(n11875), .B2(n10073), .ZN(
        n9936) );
  INV_X1 U11780 ( .A(n11875), .ZN(n14477) );
  AOI22_X1 U11781 ( .A1(n16133), .A2(n10050), .B1(n10055), .B2(n14477), .ZN(
        n9935) );
  OAI22_X1 U11782 ( .A1(n12289), .A2(n10073), .B1(n12038), .B2(n7194), .ZN(
        n9941) );
  AOI22_X1 U11783 ( .A1(n11944), .A2(n10055), .B1(n14476), .B2(n10057), .ZN(
        n9937) );
  INV_X1 U11784 ( .A(n9937), .ZN(n9938) );
  NAND2_X1 U11785 ( .A1(n9939), .A2(n9938), .ZN(n9945) );
  INV_X1 U11786 ( .A(n9940), .ZN(n9943) );
  OAI22_X1 U11787 ( .A1(n16186), .A2(n7194), .B1(n12335), .B2(n10073), .ZN(
        n9947) );
  OAI22_X1 U11788 ( .A1(n16186), .A2(n10073), .B1(n12335), .B2(n7194), .ZN(
        n9946) );
  INV_X1 U11789 ( .A(n9947), .ZN(n9948) );
  OAI22_X1 U11790 ( .A1(n12425), .A2(n10073), .B1(n12499), .B2(n7194), .ZN(
        n9950) );
  NAND2_X1 U11791 ( .A1(n9949), .A2(n9950), .ZN(n9954) );
  INV_X1 U11792 ( .A(n9949), .ZN(n9952) );
  INV_X1 U11793 ( .A(n9950), .ZN(n9951) );
  OAI22_X1 U11794 ( .A1(n16202), .A2(n7194), .B1(n14795), .B2(n10073), .ZN(
        n9955) );
  OAI22_X1 U11795 ( .A1(n16202), .A2(n10073), .B1(n14795), .B2(n7194), .ZN(
        n9957) );
  INV_X1 U11796 ( .A(n9955), .ZN(n9956) );
  AOI22_X1 U11797 ( .A1(n14800), .A2(n10050), .B1(n10055), .B2(n14472), .ZN(
        n9961) );
  INV_X1 U11798 ( .A(n9961), .ZN(n9958) );
  INV_X1 U11799 ( .A(n14800), .ZN(n14952) );
  OAI22_X1 U11800 ( .A1(n14952), .A2(n7194), .B1(n14327), .B2(n10073), .ZN(
        n9963) );
  AOI22_X1 U11801 ( .A1(n14889), .A2(n10055), .B1(n14792), .B2(n10057), .ZN(
        n9966) );
  INV_X1 U11802 ( .A(n14889), .ZN(n14777) );
  OAI22_X1 U11803 ( .A1(n14777), .A2(n10085), .B1(n12574), .B2(n7194), .ZN(
        n9965) );
  OAI21_X1 U11804 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(n9969) );
  NAND2_X1 U11805 ( .A1(n9967), .A2(n9966), .ZN(n9968) );
  OAI22_X1 U11806 ( .A1(n14879), .A2(n10085), .B1(n14381), .B2(n7194), .ZN(
        n9971) );
  OAI22_X1 U11807 ( .A1(n14879), .A2(n7194), .B1(n14381), .B2(n10073), .ZN(
        n9970) );
  INV_X1 U11808 ( .A(n9971), .ZN(n9972) );
  OAI22_X1 U11809 ( .A1(n14872), .A2(n7194), .B1(n14453), .B2(n10073), .ZN(
        n9976) );
  NAND2_X1 U11810 ( .A1(n9975), .A2(n9976), .ZN(n9974) );
  OAI22_X1 U11811 ( .A1(n14872), .A2(n10085), .B1(n14453), .B2(n7194), .ZN(
        n9973) );
  INV_X1 U11812 ( .A(n9975), .ZN(n9978) );
  INV_X1 U11813 ( .A(n9976), .ZN(n9977) );
  OAI22_X1 U11814 ( .A1(n14728), .A2(n10085), .B1(n14433), .B2(n7194), .ZN(
        n9979) );
  OAI22_X1 U11815 ( .A1(n14728), .A2(n7194), .B1(n14433), .B2(n10073), .ZN(
        n9981) );
  INV_X1 U11816 ( .A(n9979), .ZN(n9980) );
  AOI22_X1 U11817 ( .A1(n14713), .A2(n10055), .B1(n14469), .B2(n10050), .ZN(
        n9983) );
  OAI22_X1 U11818 ( .A1(n14861), .A2(n10085), .B1(n14343), .B2(n7194), .ZN(
        n9982) );
  AOI22_X1 U11819 ( .A1(n14700), .A2(n10050), .B1(n10055), .B2(n14468), .ZN(
        n9987) );
  INV_X1 U11820 ( .A(n9987), .ZN(n9985) );
  AOI22_X1 U11821 ( .A1(n14700), .A2(n10055), .B1(n14468), .B2(n10050), .ZN(
        n9984) );
  AOI21_X1 U11822 ( .B1(n9988), .B2(n9985), .A(n9984), .ZN(n9986) );
  INV_X1 U11823 ( .A(n9986), .ZN(n9989) );
  OAI22_X1 U11824 ( .A1(n14929), .A2(n7194), .B1(n14361), .B2(n10073), .ZN(
        n9991) );
  OAI22_X1 U11825 ( .A1(n14929), .A2(n10085), .B1(n14361), .B2(n7194), .ZN(
        n9990) );
  INV_X1 U11826 ( .A(n9991), .ZN(n9992) );
  OAI22_X1 U11827 ( .A1(n14925), .A2(n10085), .B1(n14289), .B2(n7194), .ZN(
        n9994) );
  OAI22_X1 U11828 ( .A1(n14925), .A2(n7194), .B1(n14289), .B2(n10073), .ZN(
        n9993) );
  INV_X1 U11829 ( .A(n9997), .ZN(n9999) );
  OAI22_X1 U11830 ( .A1(n14654), .A2(n10073), .B1(n14362), .B2(n7194), .ZN(
        n9998) );
  NAND2_X1 U11831 ( .A1(n10000), .A2(n10001), .ZN(n10004) );
  OAI22_X1 U11832 ( .A1(n14914), .A2(n7194), .B1(n14401), .B2(n10073), .ZN(
        n10003) );
  INV_X1 U11833 ( .A(n10001), .ZN(n10002) );
  AOI22_X1 U11834 ( .A1(n14830), .A2(n10055), .B1(n14633), .B2(n10050), .ZN(
        n10006) );
  INV_X1 U11835 ( .A(n14830), .ZN(n14620) );
  OAI22_X1 U11836 ( .A1(n14620), .A2(n10085), .B1(n14598), .B2(n7194), .ZN(
        n10005) );
  NAND2_X1 U11837 ( .A1(n10007), .A2(n10006), .ZN(n10013) );
  OAI22_X1 U11838 ( .A1(n14912), .A2(n7194), .B1(n14405), .B2(n10073), .ZN(
        n10008) );
  INV_X1 U11839 ( .A(n10008), .ZN(n10010) );
  AOI22_X1 U11840 ( .A1(n14601), .A2(n10057), .B1(n10055), .B2(n14614), .ZN(
        n10014) );
  INV_X1 U11841 ( .A(n10014), .ZN(n10009) );
  OR2_X1 U11842 ( .A1(n10010), .A2(n10009), .ZN(n10011) );
  NAND3_X1 U11843 ( .A1(n10012), .A2(n10014), .A3(n10013), .ZN(n10015) );
  INV_X1 U11844 ( .A(n10016), .ZN(n10017) );
  MUX2_X1 U11845 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10178), .Z(n10020) );
  NAND2_X1 U11846 ( .A1(n10020), .A2(SI_30_), .ZN(n10039) );
  OAI21_X1 U11847 ( .B1(SI_30_), .B2(n10020), .A(n10039), .ZN(n10022) );
  INV_X1 U11848 ( .A(n10022), .ZN(n10021) );
  NAND2_X1 U11849 ( .A1(n9104), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10026) );
  NAND2_X1 U11850 ( .A1(n14905), .A2(n10057), .ZN(n10029) );
  INV_X1 U11851 ( .A(n10033), .ZN(n14463) );
  NAND2_X1 U11852 ( .A1(n14463), .A2(n10055), .ZN(n10028) );
  NAND2_X1 U11853 ( .A1(n10029), .A2(n10028), .ZN(n10067) );
  INV_X1 U11854 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n14545) );
  NAND2_X1 U11855 ( .A1(n8650), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U11856 ( .A1(n8665), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n10030) );
  OAI211_X1 U11857 ( .C1(n10032), .C2(n14545), .A(n10031), .B(n10030), .ZN(
        n14548) );
  NAND2_X1 U11858 ( .A1(n14548), .A2(n10057), .ZN(n10086) );
  AOI21_X1 U11859 ( .B1(n10034), .B2(n10086), .A(n10033), .ZN(n10035) );
  AOI21_X1 U11860 ( .B1(n14905), .B2(n10055), .A(n10035), .ZN(n10068) );
  AND2_X1 U11861 ( .A1(n14464), .A2(n10050), .ZN(n10036) );
  AOI21_X1 U11862 ( .B1(n13086), .B2(n10055), .A(n10036), .ZN(n10065) );
  NAND2_X1 U11863 ( .A1(n13086), .A2(n10057), .ZN(n10038) );
  NAND2_X1 U11864 ( .A1(n14464), .A2(n10055), .ZN(n10037) );
  NAND2_X1 U11865 ( .A1(n10038), .A2(n10037), .ZN(n10064) );
  OAI22_X1 U11866 ( .A1(n10067), .A2(n10068), .B1(n10065), .B2(n10064), .ZN(
        n10047) );
  NAND2_X1 U11867 ( .A1(n10040), .A2(n10039), .ZN(n10043) );
  MUX2_X1 U11868 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10178), .Z(n10041) );
  XNOR2_X1 U11869 ( .A(n10041), .B(SI_31_), .ZN(n10042) );
  NAND2_X1 U11870 ( .A1(n15758), .A2(n10044), .ZN(n10046) );
  NAND2_X1 U11871 ( .A1(n9104), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n10045) );
  XNOR2_X1 U11872 ( .A(n14902), .B(n14548), .ZN(n10092) );
  NAND2_X1 U11873 ( .A1(n14560), .A2(n10057), .ZN(n10049) );
  NAND2_X1 U11874 ( .A1(n14465), .A2(n10055), .ZN(n10048) );
  NAND2_X1 U11875 ( .A1(n10049), .A2(n10048), .ZN(n10062) );
  INV_X1 U11876 ( .A(n10062), .ZN(n10053) );
  AND2_X1 U11877 ( .A1(n14465), .A2(n10050), .ZN(n10051) );
  AOI21_X1 U11878 ( .B1(n14560), .B2(n10055), .A(n10051), .ZN(n10063) );
  INV_X1 U11879 ( .A(n10063), .ZN(n10052) );
  NAND2_X1 U11880 ( .A1(n10053), .A2(n10052), .ZN(n10054) );
  NAND2_X1 U11881 ( .A1(n10070), .A2(n10054), .ZN(n10084) );
  INV_X1 U11882 ( .A(n10084), .ZN(n10061) );
  AND2_X1 U11883 ( .A1(n14580), .A2(n10055), .ZN(n10056) );
  AOI21_X1 U11884 ( .B1(n14569), .B2(n10050), .A(n10056), .ZN(n10077) );
  INV_X1 U11885 ( .A(n10077), .ZN(n10060) );
  NAND2_X1 U11886 ( .A1(n14569), .A2(n10055), .ZN(n10059) );
  NAND2_X1 U11887 ( .A1(n14580), .A2(n10057), .ZN(n10058) );
  NAND3_X1 U11888 ( .A1(n10061), .A2(n10060), .A3(n8475), .ZN(n10072) );
  AOI22_X1 U11889 ( .A1(n10065), .A2(n10064), .B1(n10063), .B2(n10062), .ZN(
        n10066) );
  NAND2_X1 U11890 ( .A1(n10092), .A2(n10066), .ZN(n10069) );
  AOI22_X1 U11891 ( .A1(n10070), .A2(n10069), .B1(n10068), .B2(n10067), .ZN(
        n10071) );
  AOI22_X1 U11892 ( .A1(n14819), .A2(n10050), .B1(n10055), .B2(n14466), .ZN(
        n10079) );
  OAI22_X1 U11893 ( .A1(n14584), .A2(n7194), .B1(n14599), .B2(n10073), .ZN(
        n10078) );
  NOR2_X1 U11894 ( .A1(n10079), .A2(n10078), .ZN(n10074) );
  INV_X1 U11895 ( .A(n10078), .ZN(n10081) );
  INV_X1 U11896 ( .A(n10079), .ZN(n10080) );
  OAI22_X1 U11897 ( .A1(n8475), .A2(n10060), .B1(n10081), .B2(n10080), .ZN(
        n10083) );
  OAI21_X1 U11898 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(n10090) );
  NAND2_X1 U11899 ( .A1(n14548), .A2(n10085), .ZN(n10088) );
  NAND2_X1 U11900 ( .A1(n10086), .A2(n7194), .ZN(n10087) );
  MUX2_X1 U11901 ( .A(n10088), .B(n10087), .S(n14902), .Z(n10089) );
  AND2_X1 U11902 ( .A1(n10090), .A2(n10089), .ZN(n10091) );
  INV_X1 U11903 ( .A(n7193), .ZN(n10114) );
  INV_X1 U11904 ( .A(n11399), .ZN(n10979) );
  NAND2_X1 U11905 ( .A1(n9882), .A2(n10979), .ZN(n10836) );
  AND2_X1 U11906 ( .A1(n10093), .A2(n10836), .ZN(n11523) );
  NAND4_X1 U11907 ( .A1(n11523), .A2(n9026), .A3(n9094), .A4(n11597), .ZN(
        n10095) );
  XNOR2_X1 U11908 ( .A(n14480), .B(n11418), .ZN(n11419) );
  NAND2_X1 U11909 ( .A1(n10994), .A2(n11407), .ZN(n10094) );
  NOR3_X1 U11910 ( .A1(n10095), .A2(n11419), .A3(n10094), .ZN(n10097) );
  NAND4_X1 U11911 ( .A1(n10097), .A2(n11895), .A3(n11494), .A4(n10096), .ZN(
        n10098) );
  NOR2_X1 U11912 ( .A1(n11937), .A2(n10098), .ZN(n10099) );
  NAND4_X1 U11913 ( .A1(n12405), .A2(n12329), .A3(n10099), .A4(n12140), .ZN(
        n10100) );
  NOR2_X1 U11914 ( .A1(n14786), .A2(n10100), .ZN(n10102) );
  NAND4_X1 U11915 ( .A1(n14740), .A2(n10102), .A3(n10101), .A4(n14770), .ZN(
        n10103) );
  NOR2_X1 U11916 ( .A1(n14731), .A2(n10103), .ZN(n10105) );
  NAND4_X1 U11917 ( .A1(n14681), .A2(n10105), .A3(n14688), .A4(n10104), .ZN(
        n10106) );
  OR3_X1 U11918 ( .A1(n14613), .A2(n14667), .A3(n10106), .ZN(n10107) );
  NOR4_X1 U11919 ( .A1(n14351), .A2(n10108), .A3(n14655), .A4(n10107), .ZN(
        n10111) );
  NOR2_X1 U11920 ( .A1(n12564), .A2(n10115), .ZN(n10118) );
  INV_X1 U11921 ( .A(n10116), .ZN(n10117) );
  AOI21_X1 U11922 ( .B1(n10118), .B2(n9094), .A(n10117), .ZN(n10119) );
  NOR2_X1 U11923 ( .A1(n12564), .A2(n9093), .ZN(n10122) );
  INV_X1 U11924 ( .A(n10832), .ZN(n10121) );
  AOI211_X1 U11925 ( .C1(n10976), .C2(n12683), .A(n10122), .B(n10121), .ZN(
        n10123) );
  INV_X1 U11926 ( .A(n10895), .ZN(n10125) );
  NAND2_X1 U11927 ( .A1(n10125), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10126) );
  INV_X1 U11928 ( .A(n10126), .ZN(n14972) );
  INV_X1 U11929 ( .A(P2_B_REG_SCAN_IN), .ZN(n10128) );
  NOR4_X1 U11930 ( .A1(n15818), .A2(n14794), .A3(n13321), .A4(n10832), .ZN(
        n10127) );
  AOI211_X1 U11931 ( .C1(n14972), .C2(n12683), .A(n10128), .B(n10127), .ZN(
        n10129) );
  INV_X1 U11932 ( .A(n10129), .ZN(n10130) );
  AND2_X1 U11933 ( .A1(n10895), .A2(n10131), .ZN(n10894) );
  INV_X2 U11934 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U11935 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n10138) );
  NOR2_X2 U11936 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .ZN(n10137) );
  NOR2_X2 U11937 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .ZN(n10136) );
  NAND4_X1 U11938 ( .A1(n10138), .A2(n10137), .A3(n10136), .A4(n11182), .ZN(
        n11427) );
  NAND3_X1 U11939 ( .A1(n11432), .A2(n10140), .A3(n10139), .ZN(n10141) );
  NOR2_X1 U11940 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n10147) );
  NAND2_X1 U11941 ( .A1(n10149), .A2(n10148), .ZN(n10150) );
  NAND2_X1 U11942 ( .A1(n7238), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10151) );
  OAI21_X1 U11943 ( .B1(n10152), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10153) );
  MUX2_X1 U11944 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10153), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n10154) );
  NAND2_X1 U11945 ( .A1(n10152), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10155) );
  INV_X1 U11946 ( .A(n15237), .ZN(P1_U4016) );
  NAND2_X1 U11947 ( .A1(n10178), .A2(P2_U3088), .ZN(n14975) );
  NOR2_X1 U11948 ( .A1(n10178), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14973) );
  AOI22_X1 U11949 ( .A1(n14973), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n14488), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n10156) );
  OAI21_X1 U11950 ( .B1(n10692), .B2(n14975), .A(n10156), .ZN(P2_U3326) );
  INV_X2 U11951 ( .A(n14973), .ZN(n14970) );
  INV_X1 U11952 ( .A(n11271), .ZN(n11280) );
  OAI222_X1 U11953 ( .A1(n14975), .A2(n10701), .B1(n14970), .B2(n10157), .C1(
        P2_U3088), .C2(n11280), .ZN(P2_U3325) );
  NAND2_X1 U11954 ( .A1(n10689), .A2(P3_U3151), .ZN(n10650) );
  INV_X1 U11955 ( .A(SI_3_), .ZN(n10160) );
  NOR2_X1 U11956 ( .A1(n10689), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14257) );
  INV_X1 U11957 ( .A(n14257), .ZN(n12396) );
  INV_X1 U11958 ( .A(n10158), .ZN(n10159) );
  OAI222_X1 U11959 ( .A1(P3_U3151), .A2(n10529), .B1(n14252), .B2(n10160), 
        .C1(n13319), .C2(n10159), .ZN(P3_U3292) );
  INV_X1 U11960 ( .A(n10519), .ZN(n10539) );
  INV_X1 U11961 ( .A(SI_5_), .ZN(n10163) );
  INV_X1 U11962 ( .A(n10161), .ZN(n10162) );
  OAI222_X1 U11963 ( .A1(P3_U3151), .A2(n10539), .B1(n14252), .B2(n10163), 
        .C1(n13319), .C2(n10162), .ZN(P3_U3290) );
  INV_X1 U11964 ( .A(n10164), .ZN(n10165) );
  OAI222_X1 U11965 ( .A1(P3_U3151), .A2(n10559), .B1(n14252), .B2(n10166), 
        .C1(n13319), .C2(n10165), .ZN(P3_U3293) );
  OAI222_X1 U11966 ( .A1(P3_U3151), .A2(n11016), .B1(n14252), .B2(n13671), 
        .C1(n13319), .C2(n10167), .ZN(P3_U3287) );
  INV_X1 U11967 ( .A(SI_7_), .ZN(n13673) );
  INV_X1 U11968 ( .A(n10168), .ZN(n10169) );
  OAI222_X1 U11969 ( .A1(P3_U3151), .A2(n7953), .B1(n14252), .B2(n13673), .C1(
        n13319), .C2(n10169), .ZN(P3_U3288) );
  INV_X1 U11970 ( .A(SI_4_), .ZN(n10172) );
  INV_X1 U11971 ( .A(n10170), .ZN(n10171) );
  OAI222_X1 U11972 ( .A1(P3_U3151), .A2(n7781), .B1(n14252), .B2(n10172), .C1(
        n13319), .C2(n10171), .ZN(P3_U3291) );
  OAI222_X1 U11973 ( .A1(P3_U3151), .A2(n13769), .B1(n13319), .B2(n10175), 
        .C1(n13566), .C2(n14252), .ZN(P3_U3289) );
  NAND2_X1 U11974 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10176) );
  MUX2_X1 U11975 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10176), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n10177) );
  INV_X1 U11976 ( .A(n10190), .ZN(n10196) );
  NAND2_X1 U11977 ( .A1(n10177), .A2(n10196), .ZN(n10693) );
  AND2_X1 U11978 ( .A1(n10178), .A2(n7190), .ZN(n15774) );
  INV_X2 U11979 ( .A(n15774), .ZN(n15773) );
  OAI222_X1 U11980 ( .A1(P1_U3086), .A2(n10693), .B1(n15771), .B2(n10692), 
        .C1(n10690), .C2(n15773), .ZN(P1_U3354) );
  OAI222_X1 U11981 ( .A1(P2_U3088), .A2(n14521), .B1(n14975), .B2(n11122), 
        .C1(n10179), .C2(n14970), .ZN(P2_U3323) );
  INV_X1 U11982 ( .A(n10180), .ZN(n10181) );
  OAI222_X1 U11983 ( .A1(P3_U3151), .A2(n11019), .B1(n14252), .B2(n8381), .C1(
        n13319), .C2(n10181), .ZN(P3_U3286) );
  INV_X1 U11984 ( .A(n11953), .ZN(n11583) );
  INV_X1 U11985 ( .A(SI_10_), .ZN(n13669) );
  OAI222_X1 U11986 ( .A1(P3_U3151), .A2(n11583), .B1(n14252), .B2(n13669), 
        .C1(n12396), .C2(n10182), .ZN(P3_U3285) );
  OAI222_X1 U11987 ( .A1(n14970), .A2(n10183), .B1(n14975), .B2(n11190), .C1(
        n10911), .C2(P2_U3088), .ZN(P2_U3322) );
  INV_X1 U11988 ( .A(P1_B_REG_SCAN_IN), .ZN(n15350) );
  NOR2_X1 U11989 ( .A1(n10230), .A2(n15350), .ZN(n10184) );
  MUX2_X1 U11990 ( .A(n10184), .B(n15350), .S(n12685), .Z(n10185) );
  INV_X1 U11991 ( .A(n10185), .ZN(n10186) );
  NAND2_X1 U11992 ( .A1(n10186), .A2(n10229), .ZN(n10388) );
  INV_X1 U11993 ( .A(n10388), .ZN(n10402) );
  OR2_X1 U11994 ( .A1(n10231), .A2(n10420), .ZN(n10417) );
  OR2_X1 U11995 ( .A1(n10402), .A2(n10417), .ZN(n10228) );
  INV_X1 U11996 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10389) );
  INV_X1 U11997 ( .A(n10231), .ZN(n10188) );
  INV_X1 U11998 ( .A(n10390), .ZN(n10187) );
  AOI22_X1 U11999 ( .A1(n10228), .A2(n10389), .B1(n10188), .B2(n10187), .ZN(
        P1_U3445) );
  OAI222_X1 U12000 ( .A1(n11965), .A2(P3_U3151), .B1(n13319), .B2(n10189), 
        .C1(n10650), .C2(n13666), .ZN(P3_U3284) );
  INV_X1 U12001 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10197) );
  NAND2_X1 U12002 ( .A1(n10190), .A2(n10197), .ZN(n10202) );
  INV_X1 U12003 ( .A(n10204), .ZN(n10192) );
  INV_X1 U12004 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n10191) );
  NAND2_X1 U12005 ( .A1(n10192), .A2(n10191), .ZN(n10199) );
  NAND2_X1 U12006 ( .A1(n10199), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10193) );
  MUX2_X1 U12007 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10193), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n10194) );
  AND2_X1 U12008 ( .A1(n10194), .A2(n10233), .ZN(n11191) );
  INV_X1 U12009 ( .A(n11191), .ZN(n10331) );
  OAI222_X1 U12010 ( .A1(n15773), .A2(n10195), .B1(n15771), .B2(n11190), .C1(
        n10331), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U12011 ( .A1(n7190), .A2(n15255), .B1(n15771), .B2(n10701), .C1(
        n10700), .C2(n15773), .ZN(P1_U3353) );
  NAND2_X1 U12012 ( .A1(n10204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10198) );
  MUX2_X1 U12013 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10198), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n10200) );
  NAND2_X1 U12014 ( .A1(n10200), .A2(n10199), .ZN(n15286) );
  OAI222_X1 U12015 ( .A1(P1_U3086), .A2(n15286), .B1(n15771), .B2(n11122), 
        .C1(n10201), .C2(n15773), .ZN(P1_U3351) );
  NAND2_X1 U12016 ( .A1(n10202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10203) );
  MUX2_X1 U12017 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10203), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n10205) );
  NAND2_X1 U12018 ( .A1(n10205), .A2(n10204), .ZN(n15270) );
  OAI222_X1 U12019 ( .A1(n15773), .A2(n10749), .B1(n15771), .B2(n10748), .C1(
        P1_U3086), .C2(n15270), .ZN(P1_U3352) );
  INV_X1 U12020 ( .A(n14975), .ZN(n13325) );
  INV_X1 U12021 ( .A(n13325), .ZN(n14968) );
  INV_X1 U12022 ( .A(n14504), .ZN(n10206) );
  OAI222_X1 U12023 ( .A1(n14970), .A2(n10207), .B1(n14968), .B2(n10748), .C1(
        P2_U3088), .C2(n10206), .ZN(P2_U3324) );
  NAND2_X1 U12024 ( .A1(n10421), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15775) );
  NAND2_X1 U12025 ( .A1(n10417), .A2(n15775), .ZN(n10289) );
  NAND2_X1 U12026 ( .A1(n10378), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U12027 ( .A1(n10212), .A2(n10211), .ZN(n10213) );
  AND2_X1 U12028 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n10215) );
  NAND2_X1 U12029 ( .A1(n10214), .A2(n10215), .ZN(n10216) );
  NAND2_X1 U12030 ( .A1(n10719), .A2(n15779), .ZN(n12994) );
  OAI21_X1 U12031 ( .B1(n10421), .B2(n12994), .A(n10691), .ZN(n10287) );
  AND2_X1 U12032 ( .A1(n10289), .A2(n10287), .ZN(n15914) );
  NOR2_X1 U12033 ( .A1(n15914), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U12034 ( .A1(n10650), .A2(n10222), .B1(n13319), .B2(n10221), .C1(
        n12306), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12035 ( .A(n11315), .ZN(n10226) );
  INV_X1 U12036 ( .A(n14539), .ZN(n10223) );
  OAI222_X1 U12037 ( .A1(n14970), .A2(n10224), .B1(n14968), .B2(n10226), .C1(
        P2_U3088), .C2(n10223), .ZN(P2_U3321) );
  NAND2_X1 U12038 ( .A1(n10233), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10225) );
  XNOR2_X1 U12039 ( .A(n10225), .B(P1_IR_REG_6__SCAN_IN), .ZN(n15303) );
  INV_X1 U12040 ( .A(n15303), .ZN(n15296) );
  OAI222_X1 U12041 ( .A1(n15773), .A2(n10227), .B1(n15771), .B2(n10226), .C1(
        n7190), .C2(n15296), .ZN(P1_U3349) );
  INV_X1 U12042 ( .A(n10229), .ZN(n15768) );
  INV_X1 U12043 ( .A(n10230), .ZN(n15769) );
  NAND2_X1 U12044 ( .A1(n15768), .A2(n15769), .ZN(n10387) );
  OAI22_X1 U12045 ( .A1(n15811), .A2(P1_D_REG_1__SCAN_IN), .B1(n10231), .B2(
        n10387), .ZN(n10232) );
  INV_X1 U12046 ( .A(n10232), .ZN(P1_U3446) );
  INV_X1 U12047 ( .A(n11442), .ZN(n10236) );
  OAI21_X1 U12048 ( .B1(n10233), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10234) );
  XNOR2_X1 U12049 ( .A(n10234), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11443) );
  INV_X1 U12050 ( .A(n11443), .ZN(n10317) );
  OAI222_X1 U12051 ( .A1(n15773), .A2(n10235), .B1(n15771), .B2(n10236), .C1(
        P1_U3086), .C2(n10317), .ZN(P1_U3348) );
  INV_X1 U12052 ( .A(n11166), .ZN(n11178) );
  OAI222_X1 U12053 ( .A1(n14970), .A2(n10237), .B1(n14968), .B2(n10236), .C1(
        P2_U3088), .C2(n11178), .ZN(P2_U3320) );
  INV_X1 U12054 ( .A(n11694), .ZN(n10242) );
  NAND2_X1 U12055 ( .A1(n10239), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10238) );
  MUX2_X1 U12056 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10238), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n10240) );
  OR2_X1 U12057 ( .A1(n10239), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n11426) );
  AND2_X1 U12058 ( .A1(n10240), .A2(n11426), .ZN(n11695) );
  INV_X1 U12059 ( .A(n11695), .ZN(n10347) );
  OAI222_X1 U12060 ( .A1(n15773), .A2(n10241), .B1(n15771), .B2(n10242), .C1(
        n7190), .C2(n10347), .ZN(P1_U3347) );
  INV_X1 U12061 ( .A(n10920), .ZN(n11153) );
  OAI222_X1 U12062 ( .A1(n14970), .A2(n10243), .B1(n14968), .B2(n10242), .C1(
        P2_U3088), .C2(n11153), .ZN(P2_U3319) );
  NOR2_X1 U12063 ( .A1(n14249), .A2(n10244), .ZN(n10246) );
  INV_X1 U12064 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10245) );
  NOR2_X1 U12065 ( .A1(n10276), .A2(n10245), .ZN(P3_U3240) );
  CLKBUF_X1 U12066 ( .A(n10246), .Z(n10276) );
  INV_X1 U12067 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10247) );
  NOR2_X1 U12068 ( .A1(n10276), .A2(n10247), .ZN(P3_U3247) );
  INV_X1 U12069 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10248) );
  NOR2_X1 U12070 ( .A1(n10276), .A2(n10248), .ZN(P3_U3250) );
  INV_X1 U12071 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10249) );
  NOR2_X1 U12072 ( .A1(n10276), .A2(n10249), .ZN(P3_U3248) );
  INV_X1 U12073 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10250) );
  NOR2_X1 U12074 ( .A1(n10276), .A2(n10250), .ZN(P3_U3249) );
  INV_X1 U12075 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10251) );
  NOR2_X1 U12076 ( .A1(n10246), .A2(n10251), .ZN(P3_U3244) );
  INV_X1 U12077 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10252) );
  NOR2_X1 U12078 ( .A1(n10246), .A2(n10252), .ZN(P3_U3245) );
  INV_X1 U12079 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10253) );
  NOR2_X1 U12080 ( .A1(n10246), .A2(n10253), .ZN(P3_U3236) );
  INV_X1 U12081 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10254) );
  NOR2_X1 U12082 ( .A1(n10246), .A2(n10254), .ZN(P3_U3237) );
  INV_X1 U12083 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10255) );
  NOR2_X1 U12084 ( .A1(n10246), .A2(n10255), .ZN(P3_U3238) );
  INV_X1 U12085 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10256) );
  NOR2_X1 U12086 ( .A1(n10246), .A2(n10256), .ZN(P3_U3239) );
  INV_X1 U12087 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10257) );
  NOR2_X1 U12088 ( .A1(n10276), .A2(n10257), .ZN(P3_U3257) );
  INV_X1 U12089 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10258) );
  NOR2_X1 U12090 ( .A1(n10246), .A2(n10258), .ZN(P3_U3241) );
  INV_X1 U12091 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10259) );
  NOR2_X1 U12092 ( .A1(n10246), .A2(n10259), .ZN(P3_U3242) );
  INV_X1 U12093 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10260) );
  NOR2_X1 U12094 ( .A1(n10246), .A2(n10260), .ZN(P3_U3243) );
  INV_X1 U12095 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10261) );
  NOR2_X1 U12096 ( .A1(n10246), .A2(n10261), .ZN(P3_U3258) );
  INV_X1 U12097 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10262) );
  NOR2_X1 U12098 ( .A1(n10276), .A2(n10262), .ZN(P3_U3259) );
  INV_X1 U12099 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10263) );
  NOR2_X1 U12100 ( .A1(n10246), .A2(n10263), .ZN(P3_U3260) );
  INV_X1 U12101 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10264) );
  NOR2_X1 U12102 ( .A1(n10276), .A2(n10264), .ZN(P3_U3261) );
  INV_X1 U12103 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10265) );
  NOR2_X1 U12104 ( .A1(n10276), .A2(n10265), .ZN(P3_U3262) );
  INV_X1 U12105 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10266) );
  NOR2_X1 U12106 ( .A1(n10276), .A2(n10266), .ZN(P3_U3263) );
  INV_X1 U12107 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10267) );
  NOR2_X1 U12108 ( .A1(n10276), .A2(n10267), .ZN(P3_U3251) );
  INV_X1 U12109 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10268) );
  NOR2_X1 U12110 ( .A1(n10276), .A2(n10268), .ZN(P3_U3252) );
  INV_X1 U12111 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10269) );
  NOR2_X1 U12112 ( .A1(n10276), .A2(n10269), .ZN(P3_U3253) );
  INV_X1 U12113 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10270) );
  NOR2_X1 U12114 ( .A1(n10276), .A2(n10270), .ZN(P3_U3254) );
  INV_X1 U12115 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10271) );
  NOR2_X1 U12116 ( .A1(n10276), .A2(n10271), .ZN(P3_U3255) );
  INV_X1 U12117 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10272) );
  NOR2_X1 U12118 ( .A1(n10276), .A2(n10272), .ZN(P3_U3256) );
  INV_X1 U12119 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10273) );
  NOR2_X1 U12120 ( .A1(n10276), .A2(n10273), .ZN(P3_U3235) );
  INV_X1 U12121 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U12122 ( .A1(n10276), .A2(n10274), .ZN(P3_U3234) );
  INV_X1 U12123 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10275) );
  NOR2_X1 U12124 ( .A1(n10276), .A2(n10275), .ZN(P3_U3246) );
  INV_X1 U12125 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10277) );
  MUX2_X1 U12126 ( .A(n10277), .B(P1_REG2_REG_4__SCAN_IN), .S(n15286), .Z(
        n10284) );
  XNOR2_X1 U12127 ( .A(n10693), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n15243) );
  AND2_X1 U12128 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10278) );
  NAND2_X1 U12129 ( .A1(n15243), .A2(n10278), .ZN(n15242) );
  INV_X1 U12130 ( .A(n10693), .ZN(n15244) );
  NAND2_X1 U12131 ( .A1(n15244), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U12132 ( .A1(n15242), .A2(n10279), .ZN(n15257) );
  INV_X1 U12133 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10280) );
  MUX2_X1 U12134 ( .A(n10280), .B(P1_REG2_REG_2__SCAN_IN), .S(n15255), .Z(
        n15258) );
  NAND2_X1 U12135 ( .A1(n15257), .A2(n15258), .ZN(n15272) );
  OR2_X1 U12136 ( .A1(n15255), .A2(n10280), .ZN(n15271) );
  NAND2_X1 U12137 ( .A1(n15272), .A2(n15271), .ZN(n10282) );
  INV_X1 U12138 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11068) );
  MUX2_X1 U12139 ( .A(n11068), .B(P1_REG2_REG_3__SCAN_IN), .S(n15270), .Z(
        n10281) );
  NAND2_X1 U12140 ( .A1(n10282), .A2(n10281), .ZN(n15281) );
  OR2_X1 U12141 ( .A1(n15270), .A2(n11068), .ZN(n15280) );
  NAND2_X1 U12142 ( .A1(n15281), .A2(n15280), .ZN(n10283) );
  NAND2_X1 U12143 ( .A1(n10284), .A2(n10283), .ZN(n15284) );
  INV_X1 U12144 ( .A(n15286), .ZN(n11120) );
  NAND2_X1 U12145 ( .A1(n11120), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10334) );
  INV_X1 U12146 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10285) );
  MUX2_X1 U12147 ( .A(n10285), .B(P1_REG2_REG_5__SCAN_IN), .S(n11191), .Z(
        n10335) );
  AOI21_X1 U12148 ( .B1(n15284), .B2(n10334), .A(n10335), .ZN(n15308) );
  NOR2_X1 U12149 ( .A1(n10331), .A2(n10285), .ZN(n15302) );
  INV_X1 U12150 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11381) );
  MUX2_X1 U12151 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11381), .S(n15303), .Z(
        n10286) );
  OAI21_X1 U12152 ( .B1(n15308), .B2(n15302), .A(n10286), .ZN(n15306) );
  NAND2_X1 U12153 ( .A1(n15303), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10293) );
  INV_X1 U12154 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10316) );
  MUX2_X1 U12155 ( .A(n10316), .B(P1_REG2_REG_7__SCAN_IN), .S(n11443), .Z(
        n10292) );
  AOI21_X1 U12156 ( .B1(n15306), .B2(n10293), .A(n10292), .ZN(n10324) );
  INV_X1 U12157 ( .A(n10287), .ZN(n10288) );
  NAND2_X1 U12158 ( .A1(n10289), .A2(n10288), .ZN(n15917) );
  OR2_X1 U12159 ( .A1(n10290), .A2(n15351), .ZN(n10291) );
  INV_X1 U12160 ( .A(n15338), .ZN(n15931) );
  NAND3_X1 U12161 ( .A1(n15306), .A2(n10293), .A3(n10292), .ZN(n10294) );
  NAND2_X1 U12162 ( .A1(n15931), .A2(n10294), .ZN(n10311) );
  INV_X1 U12163 ( .A(n10290), .ZN(n10715) );
  INV_X1 U12164 ( .A(n15337), .ZN(n15929) );
  INV_X1 U12165 ( .A(n15914), .ZN(n15935) );
  INV_X1 U12166 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10295) );
  NAND2_X1 U12167 ( .A1(n7190), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11456) );
  OAI21_X1 U12168 ( .B1(n15935), .B2(n10295), .A(n11456), .ZN(n10296) );
  AOI21_X1 U12169 ( .B1(n11443), .B2(n15929), .A(n10296), .ZN(n10310) );
  INV_X1 U12170 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10306) );
  INV_X1 U12171 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10305) );
  INV_X1 U12172 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10791) );
  MUX2_X1 U12173 ( .A(n10791), .B(P1_REG1_REG_1__SCAN_IN), .S(n10693), .Z(
        n15241) );
  AND2_X1 U12174 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n15240) );
  NAND2_X1 U12175 ( .A1(n15241), .A2(n15240), .ZN(n15239) );
  NAND2_X1 U12176 ( .A1(n15244), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10297) );
  NAND2_X1 U12177 ( .A1(n15239), .A2(n10297), .ZN(n15260) );
  INV_X1 U12178 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10298) );
  OR2_X1 U12179 ( .A1(n15255), .A2(n10298), .ZN(n10299) );
  NAND2_X1 U12180 ( .A1(n15259), .A2(n10299), .ZN(n15268) );
  INV_X1 U12181 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10771) );
  MUX2_X1 U12182 ( .A(n10771), .B(P1_REG1_REG_3__SCAN_IN), .S(n15270), .Z(
        n15269) );
  NAND2_X1 U12183 ( .A1(n15268), .A2(n15269), .ZN(n15267) );
  INV_X1 U12184 ( .A(n15270), .ZN(n10300) );
  NAND2_X1 U12185 ( .A1(n10300), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U12186 ( .A1(n15267), .A2(n10301), .ZN(n15289) );
  NAND2_X1 U12187 ( .A1(n11120), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10304) );
  INV_X1 U12188 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U12189 ( .A1(n15286), .A2(n10302), .ZN(n10303) );
  AND2_X1 U12190 ( .A1(n10304), .A2(n10303), .ZN(n15290) );
  NAND2_X1 U12191 ( .A1(n15289), .A2(n15290), .ZN(n15288) );
  NAND2_X1 U12192 ( .A1(n15288), .A2(n10304), .ZN(n10329) );
  MUX2_X1 U12193 ( .A(n10305), .B(P1_REG1_REG_5__SCAN_IN), .S(n11191), .Z(
        n10330) );
  NOR2_X1 U12194 ( .A1(n10329), .A2(n10330), .ZN(n10328) );
  AOI21_X1 U12195 ( .B1(n10305), .B2(n10331), .A(n10328), .ZN(n15300) );
  MUX2_X1 U12196 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10306), .S(n15303), .Z(
        n15301) );
  NAND2_X1 U12197 ( .A1(n15300), .A2(n15301), .ZN(n15299) );
  INV_X1 U12198 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n16118) );
  MUX2_X1 U12199 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n16118), .S(n11443), .Z(
        n10307) );
  INV_X1 U12200 ( .A(n15351), .ZN(n15905) );
  OAI211_X1 U12201 ( .C1(n10308), .C2(n10307), .A(n10312), .B(n15927), .ZN(
        n10309) );
  OAI211_X1 U12202 ( .C1(n10324), .C2(n10311), .A(n10310), .B(n10309), .ZN(
        P1_U3250) );
  INV_X1 U12203 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n11760) );
  MUX2_X1 U12204 ( .A(n11760), .B(P1_REG1_REG_8__SCAN_IN), .S(n11695), .Z(
        n10314) );
  AOI21_X1 U12205 ( .B1(n10314), .B2(n10313), .A(n10346), .ZN(n10327) );
  AND2_X1 U12206 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(n7190), .ZN(n11789) );
  NOR2_X1 U12207 ( .A1(n15337), .A2(n10347), .ZN(n10315) );
  AOI211_X1 U12208 ( .C1(n15914), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11789), .B(
        n10315), .ZN(n10326) );
  NOR2_X1 U12209 ( .A1(n10317), .A2(n10316), .ZN(n10322) );
  INV_X1 U12210 ( .A(n10322), .ZN(n10320) );
  INV_X1 U12211 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10318) );
  MUX2_X1 U12212 ( .A(n10318), .B(P1_REG2_REG_8__SCAN_IN), .S(n11695), .Z(
        n10319) );
  NAND2_X1 U12213 ( .A1(n10320), .A2(n10319), .ZN(n10323) );
  MUX2_X1 U12214 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10318), .S(n11695), .Z(
        n10321) );
  OAI21_X1 U12215 ( .B1(n10324), .B2(n10322), .A(n10321), .ZN(n10353) );
  OAI211_X1 U12216 ( .C1(n10324), .C2(n10323), .A(n10353), .B(n15931), .ZN(
        n10325) );
  OAI211_X1 U12217 ( .C1(n10327), .C2(n12275), .A(n10326), .B(n10325), .ZN(
        P1_U3251) );
  AOI21_X1 U12218 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(n10340) );
  NAND2_X1 U12219 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n11208) );
  INV_X1 U12220 ( .A(n11208), .ZN(n10333) );
  NOR2_X1 U12221 ( .A1(n15337), .A2(n10331), .ZN(n10332) );
  AOI211_X1 U12222 ( .C1(n15914), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n10333), .B(
        n10332), .ZN(n10339) );
  INV_X1 U12223 ( .A(n15308), .ZN(n10337) );
  NAND3_X1 U12224 ( .A1(n10335), .A2(n15284), .A3(n10334), .ZN(n10336) );
  NAND3_X1 U12225 ( .A1(n15931), .A2(n10337), .A3(n10336), .ZN(n10338) );
  OAI211_X1 U12226 ( .C1(n10340), .C2(n12275), .A(n10339), .B(n10338), .ZN(
        P1_U3248) );
  OAI222_X1 U12227 ( .A1(P3_U3151), .A2(n12311), .B1(n10650), .B2(n10342), 
        .C1(n12396), .C2(n10341), .ZN(P3_U3282) );
  INV_X1 U12228 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n16159) );
  NAND2_X1 U12229 ( .A1(n11426), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10343) );
  MUX2_X1 U12230 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10343), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n10344) );
  INV_X1 U12231 ( .A(n10344), .ZN(n10345) );
  NOR2_X1 U12232 ( .A1(n10345), .A2(n10473), .ZN(n11806) );
  MUX2_X1 U12233 ( .A(n16159), .B(P1_REG1_REG_9__SCAN_IN), .S(n11806), .Z(
        n10349) );
  AOI21_X1 U12234 ( .B1(n10347), .B2(n11760), .A(n10346), .ZN(n10348) );
  NOR2_X1 U12235 ( .A1(n10348), .A2(n10349), .ZN(n10577) );
  AOI21_X1 U12236 ( .B1(n10349), .B2(n10348), .A(n10577), .ZN(n10358) );
  AND2_X1 U12237 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11919) );
  INV_X1 U12238 ( .A(n11806), .ZN(n10585) );
  NOR2_X1 U12239 ( .A1(n15337), .A2(n10585), .ZN(n10350) );
  AOI211_X1 U12240 ( .C1(n15914), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n11919), .B(
        n10350), .ZN(n10357) );
  NAND2_X1 U12241 ( .A1(n11695), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10352) );
  INV_X1 U12242 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10584) );
  MUX2_X1 U12243 ( .A(n10584), .B(P1_REG2_REG_9__SCAN_IN), .S(n11806), .Z(
        n10351) );
  AOI21_X1 U12244 ( .B1(n10353), .B2(n10352), .A(n10351), .ZN(n15325) );
  INV_X1 U12245 ( .A(n15325), .ZN(n10355) );
  NAND3_X1 U12246 ( .A1(n10353), .A2(n10352), .A3(n10351), .ZN(n10354) );
  NAND3_X1 U12247 ( .A1(n10355), .A2(n15931), .A3(n10354), .ZN(n10356) );
  OAI211_X1 U12248 ( .C1(n10358), .C2(n12275), .A(n10357), .B(n10356), .ZN(
        P1_U3252) );
  OAI222_X1 U12249 ( .A1(n15773), .A2(n10359), .B1(n15771), .B2(n11805), .C1(
        n10585), .C2(n7190), .ZN(P1_U3346) );
  INV_X1 U12250 ( .A(n15891), .ZN(n10922) );
  OAI222_X1 U12251 ( .A1(n14970), .A2(n10360), .B1(n14975), .B2(n11805), .C1(
        n10922), .C2(P2_U3088), .ZN(P2_U3318) );
  OAI222_X1 U12252 ( .A1(n13797), .A2(P3_U3151), .B1(n13319), .B2(n10361), 
        .C1(n10650), .C2(n13624), .ZN(P3_U3281) );
  OAI222_X1 U12253 ( .A1(n13801), .A2(P3_U3151), .B1(n13319), .B2(n10362), 
        .C1(n14252), .C2(n13659), .ZN(P3_U3280) );
  INV_X1 U12254 ( .A(n10473), .ZN(n10363) );
  NAND2_X1 U12255 ( .A1(n10363), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10364) );
  XNOR2_X1 U12256 ( .A(n10364), .B(P1_IR_REG_10__SCAN_IN), .ZN(n15320) );
  INV_X1 U12257 ( .A(n15320), .ZN(n15316) );
  INV_X1 U12258 ( .A(n12016), .ZN(n10366) );
  OAI222_X1 U12259 ( .A1(n7190), .A2(n15316), .B1(n15771), .B2(n10366), .C1(
        n10365), .C2(n15773), .ZN(P1_U3345) );
  INV_X1 U12260 ( .A(n10924), .ZN(n11165) );
  OAI222_X1 U12261 ( .A1(n14970), .A2(n10367), .B1(n14968), .B2(n10366), .C1(
        n11165), .C2(P2_U3088), .ZN(P2_U3317) );
  NAND2_X1 U12262 ( .A1(n10756), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10376) );
  NAND2_X1 U12263 ( .A1(n10757), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10375) );
  NAND2_X1 U12264 ( .A1(n10761), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n10374) );
  AND2_X2 U12265 ( .A1(n13078), .A2(n10372), .ZN(n10755) );
  NAND2_X1 U12266 ( .A1(n10755), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10373) );
  NAND2_X1 U12267 ( .A1(n10214), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10377) );
  MUX2_X1 U12268 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10377), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n10379) );
  NAND2_X1 U12269 ( .A1(n12733), .A2(n12991), .ZN(n16005) );
  OR2_X1 U12270 ( .A1(n12741), .A2(n15094), .ZN(n10384) );
  NOR2_X1 U12271 ( .A1(n10689), .A2(n10380), .ZN(n10382) );
  XNOR2_X1 U12272 ( .A(n10382), .B(n10381), .ZN(n15780) );
  NAND2_X2 U12273 ( .A1(n12742), .A2(n8287), .ZN(n15095) );
  AOI22_X1 U12274 ( .A1(n10786), .A2(n11123), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n10420), .ZN(n10383) );
  OR2_X1 U12275 ( .A1(n12741), .A2(n15095), .ZN(n10386) );
  AOI22_X1 U12276 ( .A1(n10786), .A2(n15062), .B1(P1_REG1_REG_0__SCAN_IN), 
        .B2(n10420), .ZN(n10385) );
  NAND2_X1 U12277 ( .A1(n10386), .A2(n10385), .ZN(n10850) );
  XOR2_X1 U12278 ( .A(n10851), .B(n10850), .Z(n15250) );
  INV_X1 U12279 ( .A(n15250), .ZN(n10428) );
  OAI21_X1 U12280 ( .B1(n10388), .B2(P1_D_REG_1__SCAN_IN), .A(n10387), .ZN(
        n10687) );
  INV_X1 U12281 ( .A(n10687), .ZN(n11045) );
  NAND2_X1 U12282 ( .A1(n10402), .A2(n10389), .ZN(n10391) );
  NAND2_X1 U12283 ( .A1(n10391), .A2(n10390), .ZN(n11044) );
  NOR4_X1 U12284 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10400) );
  NOR4_X1 U12285 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10399) );
  INV_X1 U12286 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15810) );
  INV_X1 U12287 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15809) );
  INV_X1 U12288 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15808) );
  INV_X1 U12289 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15807) );
  NAND4_X1 U12290 ( .A1(n15810), .A2(n15809), .A3(n15808), .A4(n15807), .ZN(
        n10397) );
  NOR4_X1 U12291 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10395) );
  NOR4_X1 U12292 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10394) );
  NOR4_X1 U12293 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10393) );
  NOR4_X1 U12294 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10392) );
  NAND4_X1 U12295 ( .A1(n10395), .A2(n10394), .A3(n10393), .A4(n10392), .ZN(
        n10396) );
  NOR4_X1 U12296 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n10397), .A4(n10396), .ZN(n10398) );
  NAND3_X1 U12297 ( .A1(n10400), .A2(n10399), .A3(n10398), .ZN(n10401) );
  NAND2_X1 U12298 ( .A1(n10402), .A2(n10401), .ZN(n11043) );
  NAND3_X1 U12299 ( .A1(n11045), .A2(n10688), .A3(n11043), .ZN(n10419) );
  INV_X1 U12300 ( .A(n10417), .ZN(n10407) );
  NAND2_X1 U12301 ( .A1(n12733), .A2(n12731), .ZN(n13044) );
  INV_X1 U12302 ( .A(n13044), .ZN(n13041) );
  NAND2_X1 U12303 ( .A1(n13041), .A2(n12991), .ZN(n11046) );
  INV_X1 U12304 ( .A(n16005), .ZN(n10405) );
  NAND2_X1 U12305 ( .A1(n10405), .A2(n12730), .ZN(n10406) );
  NAND3_X1 U12306 ( .A1(n10407), .A2(n16171), .A3(n12994), .ZN(n10408) );
  OR2_X1 U12307 ( .A1(n10417), .A2(n11046), .ZN(n10409) );
  OR2_X1 U12308 ( .A1(n10409), .A2(n10419), .ZN(n10411) );
  NAND2_X1 U12309 ( .A1(n16153), .A2(n12730), .ZN(n10686) );
  NAND2_X1 U12310 ( .A1(n10756), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10415) );
  NAND2_X1 U12311 ( .A1(n10755), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10414) );
  NAND2_X1 U12312 ( .A1(n10757), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10412) );
  INV_X1 U12313 ( .A(n15437), .ZN(n15482) );
  NOR2_X1 U12314 ( .A1(n10845), .A2(n15482), .ZN(n16003) );
  INV_X1 U12315 ( .A(n12994), .ZN(n10716) );
  NAND2_X1 U12316 ( .A1(n12992), .A2(n15343), .ZN(n10416) );
  INV_X1 U12317 ( .A(n13061), .ZN(n10418) );
  INV_X1 U12318 ( .A(n15213), .ZN(n15159) );
  AOI22_X1 U12319 ( .A1(n15196), .A2(n10786), .B1(n16003), .B2(n15159), .ZN(
        n10427) );
  NAND2_X1 U12320 ( .A1(n10419), .A2(n10686), .ZN(n10425) );
  OR2_X1 U12321 ( .A1(n10421), .A2(n10420), .ZN(n10422) );
  NOR2_X1 U12322 ( .A1(n10423), .A2(n10422), .ZN(n10424) );
  NAND2_X1 U12323 ( .A1(n10425), .A2(n10424), .ZN(n10861) );
  OR2_X1 U12324 ( .A1(n10861), .A2(n7190), .ZN(n15183) );
  NAND2_X1 U12325 ( .A1(n15183), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10426) );
  OAI211_X1 U12326 ( .C1(n10428), .C2(n15205), .A(n10427), .B(n10426), .ZN(
        P1_U3232) );
  INV_X1 U12327 ( .A(SI_16_), .ZN(n13629) );
  OAI222_X1 U12328 ( .A1(P3_U3151), .A2(n13844), .B1(n14252), .B2(n13629), 
        .C1(n12396), .C2(n10429), .ZN(P3_U3279) );
  NAND2_X1 U12329 ( .A1(n13229), .A2(n10432), .ZN(n10430) );
  NAND2_X1 U12330 ( .A1(n10431), .A2(n10430), .ZN(n10442) );
  INV_X1 U12331 ( .A(n10442), .ZN(n10433) );
  OR2_X1 U12332 ( .A1(n10432), .A2(P3_U3151), .ZN(n13315) );
  NAND2_X1 U12333 ( .A1(n10462), .A2(n13315), .ZN(n10443) );
  NAND2_X1 U12334 ( .A1(n10433), .A2(n10443), .ZN(n10434) );
  INV_X2 U12335 ( .A(P3_U3897), .ZN(n13739) );
  MUX2_X1 U12336 ( .A(n10434), .B(n13739), .S(n13310), .Z(n13889) );
  INV_X1 U12337 ( .A(n10434), .ZN(n10437) );
  NAND2_X1 U12338 ( .A1(n10437), .A2(n13309), .ZN(n13899) );
  INV_X1 U12339 ( .A(n10435), .ZN(n10436) );
  AND2_X1 U12340 ( .A1(P3_U3897), .A2(n12264), .ZN(n13897) );
  NAND3_X1 U12341 ( .A1(n13899), .A2(n13895), .A3(n13877), .ZN(n10441) );
  INV_X2 U12342 ( .A(n10438), .ZN(n13309) );
  MUX2_X1 U12343 ( .A(n10523), .B(n10513), .S(n13309), .Z(n10439) );
  NAND2_X1 U12344 ( .A1(n10439), .A2(n7731), .ZN(n10561) );
  OAI21_X1 U12345 ( .B1(n7731), .B2(n10439), .A(n10561), .ZN(n10440) );
  NAND2_X1 U12346 ( .A1(n10441), .A2(n10440), .ZN(n10445) );
  AND2_X1 U12347 ( .A1(n10443), .A2(n10442), .ZN(n15817) );
  AOI22_X1 U12348 ( .A1(n15817), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10444) );
  OAI211_X1 U12349 ( .C1(n13889), .C2(n7710), .A(n10445), .B(n10444), .ZN(
        P3_U3182) );
  AND2_X1 U12350 ( .A1(n11055), .A2(n10446), .ZN(n10449) );
  INV_X1 U12351 ( .A(n10455), .ZN(n10447) );
  NAND2_X1 U12352 ( .A1(n10459), .A2(n10447), .ZN(n10448) );
  OAI211_X1 U12353 ( .C1(n10464), .C2(n10450), .A(n10449), .B(n10448), .ZN(
        n10451) );
  NAND2_X1 U12354 ( .A1(n10451), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10453) );
  NOR2_X1 U12355 ( .A1(n10462), .A2(n10477), .ZN(n13311) );
  NAND2_X1 U12356 ( .A1(n13311), .A2(n10459), .ZN(n10452) );
  NAND2_X1 U12357 ( .A1(n10453), .A2(n10452), .ZN(n10735) );
  NOR2_X1 U12358 ( .A1(n10735), .A2(n14249), .ZN(n10643) );
  NAND3_X1 U12359 ( .A1(n10464), .A2(n10454), .A3(n16222), .ZN(n10457) );
  OR2_X1 U12360 ( .A1(n10459), .A2(n10455), .ZN(n10456) );
  NAND2_X1 U12361 ( .A1(n10457), .A2(n10456), .ZN(n10458) );
  NAND2_X1 U12362 ( .A1(n13740), .A2(n11064), .ZN(n13095) );
  NAND2_X1 U12363 ( .A1(n11648), .A2(n13095), .ZN(n13263) );
  INV_X1 U12364 ( .A(n10459), .ZN(n10460) );
  NAND2_X1 U12365 ( .A1(n10460), .A2(n13311), .ZN(n10602) );
  NOR2_X1 U12366 ( .A1(n10462), .A2(n16222), .ZN(n10463) );
  NAND2_X1 U12367 ( .A1(n10464), .A2(n10463), .ZN(n10467) );
  INV_X1 U12368 ( .A(n16045), .ZN(n13294) );
  NOR2_X1 U12369 ( .A1(n16222), .A2(n13294), .ZN(n10465) );
  NAND2_X1 U12370 ( .A1(n10467), .A2(n16128), .ZN(n13411) );
  OAI22_X1 U12371 ( .A1(n16035), .A2(n13470), .B1(n11064), .B2(n13507), .ZN(
        n10468) );
  AOI21_X1 U12372 ( .B1(n13495), .B2(n13263), .A(n10468), .ZN(n10469) );
  OAI21_X1 U12373 ( .B1(n10643), .B2(n10470), .A(n10469), .ZN(P3_U3172) );
  INV_X1 U12374 ( .A(n12074), .ZN(n10475) );
  INV_X1 U12375 ( .A(n10970), .ZN(n10887) );
  OAI222_X1 U12376 ( .A1(n14970), .A2(n10471), .B1(n14968), .B2(n10475), .C1(
        P2_U3088), .C2(n10887), .ZN(P2_U3316) );
  INV_X1 U12377 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10472) );
  NAND2_X1 U12378 ( .A1(n10473), .A2(n10472), .ZN(n10631) );
  NAND2_X1 U12379 ( .A1(n10631), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10474) );
  XNOR2_X1 U12380 ( .A(n10474), .B(P1_IR_REG_11__SCAN_IN), .ZN(n12075) );
  INV_X1 U12381 ( .A(n12075), .ZN(n10581) );
  OAI222_X1 U12382 ( .A1(n15773), .A2(n10476), .B1(n15771), .B2(n10475), .C1(
        P1_U3086), .C2(n10581), .ZN(P1_U3344) );
  NAND3_X1 U12383 ( .A1(n13263), .A2(n16222), .A3(n10477), .ZN(n10479) );
  NAND2_X1 U12384 ( .A1(n13738), .A2(n14107), .ZN(n10478) );
  NAND2_X1 U12385 ( .A1(n10479), .A2(n10478), .ZN(n11060) );
  INV_X1 U12386 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10480) );
  OAI22_X1 U12387 ( .A1(n14246), .A2(n11064), .B1(n16232), .B2(n10480), .ZN(
        n10481) );
  AOI21_X1 U12388 ( .B1(n11060), .B2(n16232), .A(n10481), .ZN(n10482) );
  INV_X1 U12389 ( .A(n10482), .ZN(P3_U3390) );
  OAI222_X1 U12390 ( .A1(n13868), .A2(P3_U3151), .B1(n13319), .B2(n10483), 
        .C1(n14252), .C2(n13627), .ZN(P3_U3278) );
  MUX2_X1 U12391 ( .A(n11647), .B(n10484), .S(n13309), .Z(n10485) );
  INV_X1 U12392 ( .A(n10526), .ZN(n10573) );
  INV_X1 U12393 ( .A(n10485), .ZN(n10486) );
  MUX2_X1 U12394 ( .A(n10488), .B(n10487), .S(n13309), .Z(n10489) );
  NAND2_X1 U12395 ( .A1(n10489), .A2(n10522), .ZN(n10612) );
  INV_X1 U12396 ( .A(n10489), .ZN(n10490) );
  NAND2_X1 U12397 ( .A1(n10490), .A2(n10559), .ZN(n10491) );
  AND2_X1 U12398 ( .A1(n10612), .A2(n10491), .ZN(n10553) );
  NAND2_X1 U12399 ( .A1(n10492), .A2(n10553), .ZN(n10615) );
  NAND2_X1 U12400 ( .A1(n10615), .A2(n10612), .ZN(n10498) );
  MUX2_X1 U12401 ( .A(n10494), .B(n10493), .S(n13309), .Z(n10495) );
  NAND2_X1 U12402 ( .A1(n10495), .A2(n10628), .ZN(n13741) );
  INV_X1 U12403 ( .A(n10495), .ZN(n10496) );
  NAND2_X1 U12404 ( .A1(n10496), .A2(n10529), .ZN(n10497) );
  AND2_X1 U12405 ( .A1(n13741), .A2(n10497), .ZN(n10614) );
  MUX2_X1 U12406 ( .A(n10531), .B(n10518), .S(n13309), .Z(n10499) );
  NAND2_X1 U12407 ( .A1(n10499), .A2(n13752), .ZN(n10508) );
  INV_X1 U12408 ( .A(n10499), .ZN(n10500) );
  NAND2_X1 U12409 ( .A1(n10500), .A2(n7781), .ZN(n10501) );
  AND2_X1 U12410 ( .A1(n10508), .A2(n10501), .ZN(n13742) );
  INV_X1 U12411 ( .A(n10509), .ZN(n13743) );
  INV_X1 U12412 ( .A(n10508), .ZN(n10507) );
  MUX2_X1 U12413 ( .A(n10503), .B(n10502), .S(n13309), .Z(n10504) );
  NAND2_X1 U12414 ( .A1(n10504), .A2(n10519), .ZN(n13762) );
  INV_X1 U12415 ( .A(n10504), .ZN(n10505) );
  NAND2_X1 U12416 ( .A1(n10505), .A2(n10539), .ZN(n10506) );
  AND2_X1 U12417 ( .A1(n13762), .A2(n10506), .ZN(n10510) );
  NOR3_X1 U12418 ( .A1(n13743), .A2(n10507), .A3(n10510), .ZN(n10512) );
  NAND2_X1 U12419 ( .A1(n10511), .A2(n10510), .ZN(n10651) );
  INV_X1 U12420 ( .A(n10651), .ZN(n13765) );
  OAI21_X1 U12421 ( .B1(n10512), .B2(n13765), .A(n13897), .ZN(n10538) );
  NOR2_X1 U12422 ( .A1(n10513), .A2(n7731), .ZN(n10514) );
  NAND2_X1 U12423 ( .A1(n10524), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10515) );
  NAND2_X1 U12424 ( .A1(n10559), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10516) );
  NAND2_X1 U12425 ( .A1(n10540), .A2(n10516), .ZN(n10517) );
  OAI21_X1 U12426 ( .B1(n10517), .B2(n10529), .A(n13753), .ZN(n10617) );
  MUX2_X1 U12427 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10518), .S(n13752), .Z(
        n13754) );
  AOI21_X1 U12428 ( .B1(n13755), .B2(n13753), .A(n13754), .ZN(n13757) );
  AOI21_X1 U12429 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n7781), .A(n13757), .ZN(
        n10520) );
  NOR2_X1 U12430 ( .A1(n10520), .A2(n10519), .ZN(n13780) );
  OAI21_X1 U12431 ( .B1(n10521), .B2(P3_REG1_REG_5__SCAN_IN), .A(n13778), .ZN(
        n10536) );
  NOR2_X1 U12432 ( .A1(n10523), .A2(n7731), .ZN(n10525) );
  NAND2_X1 U12433 ( .A1(n10524), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10527) );
  OAI21_X1 U12434 ( .B1(n10526), .B2(n10525), .A(n10527), .ZN(n10567) );
  NAND2_X1 U12435 ( .A1(n10569), .A2(n10527), .ZN(n10545) );
  NAND2_X1 U12436 ( .A1(n10559), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10528) );
  INV_X1 U12437 ( .A(n10530), .ZN(n13745) );
  MUX2_X1 U12438 ( .A(n10531), .B(P3_REG2_REG_4__SCAN_IN), .S(n13752), .Z(
        n13746) );
  AOI21_X1 U12439 ( .B1(n10503), .B2(n10532), .A(n13775), .ZN(n10534) );
  NOR2_X1 U12440 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9346), .ZN(n11304) );
  AOI21_X1 U12441 ( .B1(n15817), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11304), .ZN(
        n10533) );
  OAI21_X1 U12442 ( .B1(n10534), .B2(n13895), .A(n10533), .ZN(n10535) );
  AOI21_X1 U12443 ( .B1(n13865), .B2(n10536), .A(n10535), .ZN(n10537) );
  OAI211_X1 U12444 ( .C1(n13889), .C2(n10539), .A(n10538), .B(n10537), .ZN(
        P3_U3187) );
  OAI21_X1 U12445 ( .B1(n10542), .B2(n10541), .A(n10540), .ZN(n10550) );
  INV_X1 U12446 ( .A(n15817), .ZN(n13842) );
  INV_X1 U12447 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10543) );
  OAI22_X1 U12448 ( .A1(n13842), .A2(n10543), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n16044), .ZN(n10549) );
  INV_X1 U12449 ( .A(n13895), .ZN(n13838) );
  OAI21_X1 U12450 ( .B1(n10546), .B2(n10545), .A(n10544), .ZN(n10547) );
  AND2_X1 U12451 ( .A1(n13838), .A2(n10547), .ZN(n10548) );
  AOI211_X1 U12452 ( .C1(n13865), .C2(n10550), .A(n10549), .B(n10548), .ZN(
        n10558) );
  INV_X1 U12453 ( .A(n10551), .ZN(n10560) );
  INV_X1 U12454 ( .A(n10552), .ZN(n10554) );
  NOR3_X1 U12455 ( .A1(n10560), .A2(n10554), .A3(n10553), .ZN(n10556) );
  INV_X1 U12456 ( .A(n10615), .ZN(n10555) );
  OAI21_X1 U12457 ( .B1(n10556), .B2(n10555), .A(n13897), .ZN(n10557) );
  OAI211_X1 U12458 ( .C1(n13889), .C2(n10559), .A(n10558), .B(n10557), .ZN(
        P3_U3184) );
  AOI21_X1 U12459 ( .B1(n10562), .B2(n10561), .A(n10560), .ZN(n10576) );
  INV_X1 U12460 ( .A(n10563), .ZN(n10565) );
  OAI21_X1 U12461 ( .B1(n10565), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10564), .ZN(
        n10572) );
  INV_X1 U12462 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n10566) );
  OAI22_X1 U12463 ( .A1(n13842), .A2(n10566), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10603), .ZN(n10571) );
  NAND2_X1 U12464 ( .A1(n10567), .A2(n11647), .ZN(n10568) );
  AOI21_X1 U12465 ( .B1(n10569), .B2(n10568), .A(n13895), .ZN(n10570) );
  AOI211_X1 U12466 ( .C1(n13865), .C2(n10572), .A(n10571), .B(n10570), .ZN(
        n10575) );
  NAND2_X1 U12467 ( .A1(n13874), .A2(n10573), .ZN(n10574) );
  OAI211_X1 U12468 ( .C1(n10576), .C2(n13877), .A(n10575), .B(n10574), .ZN(
        P3_U3183) );
  INV_X1 U12469 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n12392) );
  MUX2_X1 U12470 ( .A(n12392), .B(P1_REG1_REG_11__SCAN_IN), .S(n12075), .Z(
        n10580) );
  INV_X1 U12471 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10578) );
  AOI21_X1 U12472 ( .B1(n16159), .B2(n10585), .A(n10577), .ZN(n15314) );
  MUX2_X1 U12473 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10578), .S(n15320), .Z(
        n15313) );
  NAND2_X1 U12474 ( .A1(n15314), .A2(n15313), .ZN(n15312) );
  AOI21_X1 U12475 ( .B1(n10580), .B2(n10579), .A(n15926), .ZN(n10595) );
  INV_X1 U12476 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n12375) );
  NOR2_X1 U12477 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12375), .ZN(n10583) );
  NOR2_X1 U12478 ( .A1(n15337), .A2(n10581), .ZN(n10582) );
  AOI211_X1 U12479 ( .C1(n15914), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10583), 
        .B(n10582), .ZN(n10594) );
  NOR2_X1 U12480 ( .A1(n10585), .A2(n10584), .ZN(n15319) );
  INV_X1 U12481 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10586) );
  MUX2_X1 U12482 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10586), .S(n15320), .Z(
        n10587) );
  OAI21_X1 U12483 ( .B1(n15325), .B2(n15319), .A(n10587), .ZN(n15323) );
  NAND2_X1 U12484 ( .A1(n15320), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10590) );
  INV_X1 U12485 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10588) );
  MUX2_X1 U12486 ( .A(n10588), .B(P1_REG2_REG_11__SCAN_IN), .S(n12075), .Z(
        n10589) );
  AOI21_X1 U12487 ( .B1(n15323), .B2(n10590), .A(n10589), .ZN(n10944) );
  INV_X1 U12488 ( .A(n10944), .ZN(n10592) );
  NAND3_X1 U12489 ( .A1(n15323), .A2(n10590), .A3(n10589), .ZN(n10591) );
  NAND3_X1 U12490 ( .A1(n10592), .A2(n15931), .A3(n10591), .ZN(n10593) );
  OAI211_X1 U12491 ( .C1(n10595), .C2(n12275), .A(n10594), .B(n10593), .ZN(
        P1_U3254) );
  OAI21_X1 U12492 ( .B1(n7765), .B2(n10597), .A(n11642), .ZN(n10599) );
  NAND2_X1 U12493 ( .A1(n11064), .A2(n7765), .ZN(n10598) );
  AOI21_X1 U12494 ( .B1(n10600), .B2(n10599), .A(n10640), .ZN(n10607) );
  OR2_X1 U12495 ( .A1(n10602), .A2(n10601), .ZN(n13500) );
  INV_X1 U12496 ( .A(n13500), .ZN(n12630) );
  INV_X1 U12497 ( .A(n13523), .ZN(n13100) );
  OAI22_X1 U12498 ( .A1(n13100), .A2(n13470), .B1(n11640), .B2(n13507), .ZN(
        n10605) );
  NOR2_X1 U12499 ( .A1(n10643), .A2(n10603), .ZN(n10604) );
  AOI211_X1 U12500 ( .C1(n12630), .C2(n13740), .A(n10605), .B(n10604), .ZN(
        n10606) );
  OAI21_X1 U12501 ( .B1(n10607), .B2(n13440), .A(n10606), .ZN(P3_U3162) );
  INV_X2 U12502 ( .A(P2_U3947), .ZN(n14485) );
  NAND2_X1 U12503 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n14485), .ZN(n10608) );
  OAI21_X1 U12504 ( .B1(n14433), .B2(n14485), .A(n10608), .ZN(P2_U3548) );
  INV_X1 U12505 ( .A(n13884), .ZN(n10610) );
  OAI222_X1 U12506 ( .A1(P3_U3151), .A2(n10610), .B1(n10650), .B2(n13630), 
        .C1(n12396), .C2(n10609), .ZN(P3_U3277) );
  INV_X1 U12507 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12686) );
  NAND2_X1 U12508 ( .A1(n14633), .A2(P2_U3947), .ZN(n10611) );
  OAI21_X1 U12509 ( .B1(n12686), .B2(P2_U3947), .A(n10611), .ZN(P2_U3555) );
  INV_X1 U12510 ( .A(n10612), .ZN(n10613) );
  NOR2_X1 U12511 ( .A1(n10614), .A2(n10613), .ZN(n10616) );
  AOI21_X1 U12512 ( .B1(n10616), .B2(n10615), .A(n7357), .ZN(n10630) );
  NAND2_X1 U12513 ( .A1(n10617), .A2(n10493), .ZN(n10618) );
  NAND2_X1 U12514 ( .A1(n13755), .A2(n10618), .ZN(n10619) );
  NAND2_X1 U12515 ( .A1(n13865), .A2(n10619), .ZN(n10626) );
  NAND2_X1 U12516 ( .A1(n10620), .A2(n10494), .ZN(n10621) );
  NAND2_X1 U12517 ( .A1(n10622), .A2(n10621), .ZN(n10623) );
  NAND2_X1 U12518 ( .A1(n13838), .A2(n10623), .ZN(n10625) );
  NOR2_X1 U12519 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13696), .ZN(n10743) );
  AOI21_X1 U12520 ( .B1(n15817), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10743), .ZN(
        n10624) );
  NAND3_X1 U12521 ( .A1(n10626), .A2(n10625), .A3(n10624), .ZN(n10627) );
  AOI21_X1 U12522 ( .B1(n10628), .B2(n13874), .A(n10627), .ZN(n10629) );
  OAI21_X1 U12523 ( .B1(n10630), .B2(n13877), .A(n10629), .ZN(P3_U3185) );
  INV_X1 U12524 ( .A(n12187), .ZN(n10634) );
  NAND2_X1 U12525 ( .A1(n11184), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10680) );
  XNOR2_X1 U12526 ( .A(n10680), .B(P1_IR_REG_12__SCAN_IN), .ZN(n15930) );
  INV_X1 U12527 ( .A(n15930), .ZN(n10632) );
  OAI222_X1 U12528 ( .A1(n15773), .A2(n10633), .B1(n15771), .B2(n10634), .C1(
        n10632), .C2(P1_U3086), .ZN(P1_U3343) );
  OAI222_X1 U12529 ( .A1(n14970), .A2(n10635), .B1(n14968), .B2(n10634), .C1(
        n10926), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI22_X1 U12530 ( .A1(n14192), .A2(n11064), .B1(n16228), .B2(n10513), .ZN(
        n10636) );
  AOI21_X1 U12531 ( .B1(n11060), .B2(n16228), .A(n10636), .ZN(n10637) );
  INV_X1 U12532 ( .A(n10637), .ZN(P3_U3459) );
  INV_X1 U12533 ( .A(n10638), .ZN(n10639) );
  AOI21_X1 U12534 ( .B1(n10642), .B2(n10641), .A(n10740), .ZN(n10647) );
  INV_X1 U12535 ( .A(n13522), .ZN(n16033) );
  OAI22_X1 U12536 ( .A1(n16033), .A2(n13470), .B1(n13507), .B2(n16029), .ZN(
        n10645) );
  NOR2_X1 U12537 ( .A1(n10643), .A2(n16044), .ZN(n10644) );
  AOI211_X1 U12538 ( .C1(n12630), .C2(n13738), .A(n10645), .B(n10644), .ZN(
        n10646) );
  OAI21_X1 U12539 ( .B1(n10647), .B2(n13440), .A(n10646), .ZN(P3_U3177) );
  OAI222_X1 U12540 ( .A1(n10650), .A2(n10649), .B1(P3_U3151), .B2(n13888), 
        .C1(n12396), .C2(n10648), .ZN(P3_U3276) );
  NAND2_X1 U12541 ( .A1(n10651), .A2(n13762), .ZN(n10657) );
  MUX2_X1 U12542 ( .A(n10652), .B(n10667), .S(n13309), .Z(n10654) );
  INV_X1 U12543 ( .A(n13769), .ZN(n10653) );
  NAND2_X1 U12544 ( .A1(n10654), .A2(n10653), .ZN(n10665) );
  INV_X1 U12545 ( .A(n10654), .ZN(n10655) );
  NAND2_X1 U12546 ( .A1(n10655), .A2(n13769), .ZN(n10656) );
  AND2_X1 U12547 ( .A1(n10665), .A2(n10656), .ZN(n13763) );
  MUX2_X1 U12548 ( .A(n10659), .B(n10658), .S(n13309), .Z(n10660) );
  NAND2_X1 U12549 ( .A1(n10660), .A2(n10803), .ZN(n10812) );
  INV_X1 U12550 ( .A(n10660), .ZN(n10661) );
  NAND2_X1 U12551 ( .A1(n10661), .A2(n7953), .ZN(n10662) );
  AND2_X1 U12552 ( .A1(n10812), .A2(n10662), .ZN(n10663) );
  INV_X1 U12553 ( .A(n10663), .ZN(n10664) );
  NAND3_X1 U12554 ( .A1(n13766), .A2(n10665), .A3(n10664), .ZN(n10666) );
  AOI21_X1 U12555 ( .B1(n10813), .B2(n10666), .A(n13877), .ZN(n10678) );
  INV_X1 U12556 ( .A(n13780), .ZN(n10668) );
  MUX2_X1 U12557 ( .A(n10667), .B(P3_REG1_REG_6__SCAN_IN), .S(n13769), .Z(
        n13779) );
  AOI21_X1 U12558 ( .B1(n10658), .B2(n10669), .A(n10796), .ZN(n10670) );
  NOR2_X1 U12559 ( .A1(n10670), .A2(n13899), .ZN(n10677) );
  MUX2_X1 U12560 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n10652), .S(n13769), .Z(
        n13774) );
  INV_X1 U12561 ( .A(n13774), .ZN(n10671) );
  AOI21_X1 U12562 ( .B1(n10659), .B2(n10672), .A(n10804), .ZN(n10675) );
  AND2_X1 U12563 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11797) );
  NOR2_X1 U12564 ( .A1(n13889), .A2(n7953), .ZN(n10673) );
  AOI211_X1 U12565 ( .C1(n15817), .C2(P3_ADDR_REG_7__SCAN_IN), .A(n11797), .B(
        n10673), .ZN(n10674) );
  OAI21_X1 U12566 ( .B1(n10675), .B2(n13895), .A(n10674), .ZN(n10676) );
  OR3_X1 U12567 ( .A1(n10678), .A2(n10677), .A3(n10676), .ZN(P3_U3189) );
  INV_X1 U12568 ( .A(n11367), .ZN(n11380) );
  INV_X1 U12569 ( .A(n12192), .ZN(n10684) );
  OAI222_X1 U12570 ( .A1(P2_U3088), .A2(n11380), .B1(n14968), .B2(n10684), 
        .C1(n10679), .C2(n14970), .ZN(P2_U3314) );
  INV_X1 U12571 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n11181) );
  AOI21_X1 U12572 ( .B1(n10680), .B2(n11181), .A(n8078), .ZN(n10681) );
  NAND2_X1 U12573 ( .A1(n10681), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n10683) );
  INV_X1 U12574 ( .A(n10681), .ZN(n10682) );
  NAND2_X1 U12575 ( .A1(n10682), .A2(n11182), .ZN(n10820) );
  INV_X1 U12576 ( .A(n12193), .ZN(n10952) );
  OAI222_X1 U12577 ( .A1(n15773), .A2(n10685), .B1(n15771), .B2(n10684), .C1(
        n10952), .C2(n7190), .ZN(P1_U3342) );
  NAND4_X1 U12578 ( .A1(n13061), .A2(n10687), .A3(n11043), .A4(n10686), .ZN(
        n10731) );
  OR2_X1 U12579 ( .A1(n10731), .A2(n10688), .ZN(n16180) );
  INV_X1 U12580 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10730) );
  INV_X1 U12581 ( .A(n10725), .ZN(n12737) );
  NAND2_X1 U12582 ( .A1(n10845), .A2(n10725), .ZN(n12744) );
  INV_X1 U12583 ( .A(n10786), .ZN(n16013) );
  NOR2_X1 U12584 ( .A1(n12741), .A2(n16013), .ZN(n10781) );
  INV_X1 U12585 ( .A(n10781), .ZN(n10694) );
  NAND2_X1 U12586 ( .A1(n10845), .A2(n12737), .ZN(n10695) );
  NAND2_X1 U12587 ( .A1(n10756), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10699) );
  NAND2_X1 U12588 ( .A1(n10757), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n10698) );
  NAND2_X1 U12589 ( .A1(n10761), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n10697) );
  NAND2_X1 U12590 ( .A1(n10755), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10696) );
  OR2_X1 U12591 ( .A1(n13000), .A2(n10700), .ZN(n10704) );
  OR2_X1 U12592 ( .A1(n12987), .A2(n10701), .ZN(n10703) );
  OR2_X1 U12593 ( .A1(n10691), .A2(n15255), .ZN(n10702) );
  NAND2_X1 U12594 ( .A1(n10864), .A2(n12749), .ZN(n10746) );
  OAI21_X1 U12595 ( .B1(n10706), .B2(n10718), .A(n10747), .ZN(n11052) );
  INV_X1 U12596 ( .A(n11052), .ZN(n10728) );
  AND2_X1 U12597 ( .A1(n12991), .A2(n12730), .ZN(n10707) );
  NOR2_X1 U12598 ( .A1(n12991), .A2(n12730), .ZN(n10708) );
  NAND2_X1 U12599 ( .A1(n12742), .A2(n15779), .ZN(n10709) );
  NAND2_X1 U12600 ( .A1(n15065), .A2(n10709), .ZN(n12168) );
  INV_X1 U12601 ( .A(n12168), .ZN(n10710) );
  INV_X1 U12602 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10758) );
  NAND2_X1 U12603 ( .A1(n10757), .A2(n10758), .ZN(n10714) );
  NAND2_X1 U12604 ( .A1(n10755), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10713) );
  NAND2_X1 U12605 ( .A1(n10761), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n10712) );
  NAND2_X1 U12606 ( .A1(n10756), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10711) );
  NAND4_X1 U12607 ( .A1(n10714), .A2(n10713), .A3(n10712), .A4(n10711), .ZN(
        n15235) );
  INV_X1 U12608 ( .A(n15235), .ZN(n11233) );
  INV_X1 U12609 ( .A(n15500), .ZN(n15484) );
  OAI22_X1 U12610 ( .A1(n11233), .A2(n15482), .B1(n10845), .B2(n15484), .ZN(
        n10724) );
  INV_X1 U12611 ( .A(n10717), .ZN(n10778) );
  NAND2_X1 U12612 ( .A1(n12741), .A2(n10786), .ZN(n13010) );
  INV_X1 U12613 ( .A(n13010), .ZN(n12746) );
  NAND2_X1 U12614 ( .A1(n10782), .A2(n12744), .ZN(n10752) );
  XNOR2_X1 U12615 ( .A(n10752), .B(n10718), .ZN(n10722) );
  NAND2_X1 U12616 ( .A1(n10719), .A2(n12731), .ZN(n10721) );
  NAND2_X1 U12617 ( .A1(n15779), .A2(n12730), .ZN(n10720) );
  NOR2_X1 U12618 ( .A1(n10722), .A2(n16074), .ZN(n10723) );
  AOI211_X1 U12619 ( .C1(n15490), .C2(n11052), .A(n10724), .B(n10723), .ZN(
        n11054) );
  OR2_X1 U12620 ( .A1(n15109), .A2(n10786), .ZN(n10788) );
  NAND2_X1 U12621 ( .A1(n15181), .A2(n10788), .ZN(n10726) );
  AND2_X1 U12622 ( .A1(n10768), .A2(n10726), .ZN(n11049) );
  AOI22_X1 U12623 ( .A1(n11049), .A2(n16153), .B1(n15181), .B2(n16151), .ZN(
        n10727) );
  OAI211_X1 U12624 ( .C1(n10728), .C2(n16116), .A(n11054), .B(n10727), .ZN(
        n10732) );
  NAND2_X1 U12625 ( .A1(n10732), .A2(n16183), .ZN(n10729) );
  OAI21_X1 U12626 ( .B1(n16183), .B2(n10730), .A(n10729), .ZN(P1_U3465) );
  OR2_X1 U12627 ( .A1(n10731), .A2(n11044), .ZN(n16178) );
  INV_X2 U12628 ( .A(n16178), .ZN(n16179) );
  NAND2_X1 U12629 ( .A1(n10732), .A2(n16179), .ZN(n10733) );
  OAI21_X1 U12630 ( .B1(n16179), .B2(n10298), .A(n10733), .ZN(P1_U3530) );
  INV_X1 U12631 ( .A(n13315), .ZN(n10734) );
  OR2_X1 U12632 ( .A1(n10735), .A2(n10734), .ZN(n13503) );
  INV_X1 U12633 ( .A(n13503), .ZN(n12627) );
  NOR2_X1 U12634 ( .A1(n10736), .A2(n13523), .ZN(n10739) );
  XNOR2_X1 U12635 ( .A(n11098), .B(n13522), .ZN(n10738) );
  OAI21_X1 U12636 ( .B1(n10740), .B2(n10739), .A(n10738), .ZN(n10741) );
  NAND3_X1 U12637 ( .A1(n8342), .A2(n13495), .A3(n10741), .ZN(n10745) );
  OAI22_X1 U12638 ( .A1(n13100), .A2(n13500), .B1(n7730), .B2(n13470), .ZN(
        n10742) );
  AOI211_X1 U12639 ( .C1(n16053), .C2(n13411), .A(n10743), .B(n10742), .ZN(
        n10744) );
  OAI211_X1 U12640 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12627), .A(n10745), .B(
        n10744), .ZN(P3_U3158) );
  NAND2_X1 U12641 ( .A1(n10750), .A2(n13013), .ZN(n11235) );
  OAI21_X1 U12642 ( .B1(n10750), .B2(n13013), .A(n11235), .ZN(n10751) );
  INV_X1 U12643 ( .A(n10751), .ZN(n11073) );
  NAND2_X1 U12644 ( .A1(n10752), .A2(n13012), .ZN(n10754) );
  NAND2_X1 U12645 ( .A1(n10864), .A2(n15181), .ZN(n10753) );
  XNOR2_X1 U12646 ( .A(n11238), .B(n12754), .ZN(n10766) );
  NAND2_X1 U12647 ( .A1(n12875), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10765) );
  NAND2_X1 U12648 ( .A1(n12966), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10764) );
  INV_X1 U12649 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U12650 ( .A1(n10759), .A2(n10758), .ZN(n10760) );
  INV_X1 U12651 ( .A(n11131), .ZN(n11133) );
  AND2_X1 U12652 ( .A1(n10760), .A2(n11133), .ZN(n11359) );
  NAND2_X1 U12653 ( .A1(n12965), .A2(n11359), .ZN(n10763) );
  NAND2_X1 U12654 ( .A1(n10761), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10762) );
  AOI222_X1 U12655 ( .A1(n15723), .A2(n10766), .B1(n15234), .B2(n15583), .C1(
        n15236), .C2(n15500), .ZN(n11067) );
  INV_X1 U12656 ( .A(n11358), .ZN(n10767) );
  AOI21_X1 U12657 ( .B1(n12757), .B2(n10768), .A(n10767), .ZN(n11070) );
  AOI22_X1 U12658 ( .A1(n11070), .A2(n16153), .B1(n12757), .B2(n16151), .ZN(
        n10769) );
  OAI211_X1 U12659 ( .C1(n15732), .C2(n11073), .A(n11067), .B(n10769), .ZN(
        n10772) );
  NAND2_X1 U12660 ( .A1(n10772), .A2(n16179), .ZN(n10770) );
  OAI21_X1 U12661 ( .B1(n16179), .B2(n10771), .A(n10770), .ZN(P1_U3531) );
  INV_X1 U12662 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U12663 ( .A1(n10772), .A2(n16183), .ZN(n10773) );
  OAI21_X1 U12664 ( .B1(n16183), .B2(n10774), .A(n10773), .ZN(P1_U3468) );
  OAI222_X1 U12665 ( .A1(n12396), .A2(n10777), .B1(n10650), .B2(n10776), .C1(
        P3_U3151), .C2(n10775), .ZN(P3_U3275) );
  INV_X1 U12666 ( .A(n10779), .ZN(n10780) );
  AOI21_X1 U12667 ( .B1(n10781), .B2(n10778), .A(n10780), .ZN(n11074) );
  OAI21_X1 U12668 ( .B1(n10778), .B2(n12746), .A(n10782), .ZN(n10785) );
  OAI22_X1 U12669 ( .A1(n12741), .A2(n15484), .B1(n10864), .B2(n15482), .ZN(
        n10784) );
  NOR2_X1 U12670 ( .A1(n11074), .A2(n16002), .ZN(n10783) );
  AOI211_X1 U12671 ( .C1(n15723), .C2(n10785), .A(n10784), .B(n10783), .ZN(
        n11081) );
  NAND2_X1 U12672 ( .A1(n15109), .A2(n10786), .ZN(n10787) );
  AND3_X1 U12673 ( .A1(n10788), .A2(n16153), .A3(n10787), .ZN(n11075) );
  AOI21_X1 U12674 ( .B1(n15109), .B2(n16151), .A(n11075), .ZN(n10789) );
  OAI211_X1 U12675 ( .C1(n11074), .C2(n16116), .A(n11081), .B(n10789), .ZN(
        n10792) );
  NAND2_X1 U12676 ( .A1(n10792), .A2(n16179), .ZN(n10790) );
  OAI21_X1 U12677 ( .B1(n16179), .B2(n10791), .A(n10790), .ZN(P1_U3529) );
  INV_X1 U12678 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10794) );
  NAND2_X1 U12679 ( .A1(n10792), .A2(n16183), .ZN(n10793) );
  OAI21_X1 U12680 ( .B1(n16183), .B2(n10794), .A(n10793), .ZN(P1_U3462) );
  NOR2_X1 U12681 ( .A1(n10803), .A2(n10795), .ZN(n10797) );
  MUX2_X1 U12682 ( .A(n10798), .B(P3_REG1_REG_8__SCAN_IN), .S(n11016), .Z(
        n10800) );
  INV_X1 U12683 ( .A(n11013), .ZN(n10799) );
  AOI21_X1 U12684 ( .B1(n10801), .B2(n10800), .A(n10799), .ZN(n10819) );
  NOR2_X1 U12685 ( .A1(n10803), .A2(n10802), .ZN(n10805) );
  MUX2_X1 U12686 ( .A(n10806), .B(P3_REG2_REG_8__SCAN_IN), .S(n11016), .Z(
        n10807) );
  OAI21_X1 U12687 ( .B1(n7232), .B2(n7442), .A(n11018), .ZN(n10811) );
  INV_X1 U12688 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10808) );
  NOR2_X1 U12689 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10808), .ZN(n11931) );
  AOI21_X1 U12690 ( .B1(n15817), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11931), .ZN(
        n10809) );
  OAI21_X1 U12691 ( .B1(n13889), .B2(n11016), .A(n10809), .ZN(n10810) );
  AOI21_X1 U12692 ( .B1(n10811), .B2(n13838), .A(n10810), .ZN(n10818) );
  MUX2_X1 U12693 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13309), .Z(n11002) );
  INV_X1 U12694 ( .A(n11016), .ZN(n11003) );
  XNOR2_X1 U12695 ( .A(n11002), .B(n11003), .ZN(n10814) );
  NAND2_X1 U12696 ( .A1(n10815), .A2(n10814), .ZN(n11006) );
  OAI21_X1 U12697 ( .B1(n10815), .B2(n10814), .A(n11006), .ZN(n10816) );
  NAND2_X1 U12698 ( .A1(n10816), .A2(n13897), .ZN(n10817) );
  OAI211_X1 U12699 ( .C1(n10819), .C2(n13899), .A(n10818), .B(n10817), .ZN(
        P3_U3190) );
  INV_X1 U12700 ( .A(n12520), .ZN(n10823) );
  NAND2_X1 U12701 ( .A1(n10820), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10821) );
  XNOR2_X1 U12702 ( .A(n10821), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12521) );
  INV_X1 U12703 ( .A(n12521), .ZN(n11735) );
  OAI222_X1 U12704 ( .A1(n15773), .A2(n10822), .B1(n15771), .B2(n10823), .C1(
        n7190), .C2(n11735), .ZN(P1_U3341) );
  INV_X1 U12705 ( .A(n10901), .ZN(n11861) );
  OAI222_X1 U12706 ( .A1(n14970), .A2(n10824), .B1(n14968), .B2(n10823), .C1(
        P2_U3088), .C2(n11861), .ZN(P2_U3313) );
  NAND2_X1 U12707 ( .A1(n10826), .A2(n10825), .ZN(n10830) );
  OAI21_X1 U12708 ( .B1(n15820), .B2(n10830), .A(n10838), .ZN(n10829) );
  AND3_X1 U12709 ( .A1(n11514), .A2(n10895), .A3(n10827), .ZN(n10828) );
  NAND2_X1 U12710 ( .A1(n10829), .A2(n10828), .ZN(n11091) );
  NOR2_X1 U12711 ( .A1(n11091), .A2(P2_U3088), .ZN(n11227) );
  INV_X1 U12712 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11519) );
  AND2_X1 U12713 ( .A1(n14484), .A2(n14791), .ZN(n11228) );
  INV_X1 U12714 ( .A(n10830), .ZN(n11515) );
  NAND2_X1 U12715 ( .A1(n15821), .A2(n11515), .ZN(n10831) );
  OR2_X1 U12716 ( .A1(n15820), .A2(n10831), .ZN(n10839) );
  NOR2_X2 U12717 ( .A1(n10839), .A2(n10832), .ZN(n14392) );
  INV_X1 U12718 ( .A(n10839), .ZN(n10835) );
  INV_X1 U12719 ( .A(n10896), .ZN(n10833) );
  AND2_X1 U12720 ( .A1(n16201), .A2(n10833), .ZN(n10834) );
  NOR3_X1 U12721 ( .A1(n14449), .A2(n14267), .A3(n10836), .ZN(n10837) );
  AOI21_X1 U12722 ( .B1(n11228), .B2(n14392), .A(n10837), .ZN(n10842) );
  AOI21_X1 U12723 ( .B1(n14300), .B2(n9882), .A(n14449), .ZN(n10840) );
  NAND2_X1 U12724 ( .A1(n11230), .A2(n9094), .ZN(n11550) );
  OAI21_X1 U12725 ( .B1(n10840), .B2(n14423), .A(n11399), .ZN(n10841) );
  OAI211_X1 U12726 ( .C1(n11227), .C2(n11519), .A(n10842), .B(n10841), .ZN(
        P2_U3204) );
  OAI22_X1 U12727 ( .A1(n11233), .A2(n15095), .B1(n8021), .B2(n15096), .ZN(
        n10843) );
  OAI22_X1 U12728 ( .A1(n11233), .A2(n15094), .B1(n8021), .B2(n15095), .ZN(
        n11119) );
  XNOR2_X1 U12729 ( .A(n11118), .B(n11119), .ZN(n10860) );
  OAI22_X1 U12730 ( .A1(n10845), .A2(n15095), .B1(n12737), .B2(n15096), .ZN(
        n10844) );
  XNOR2_X1 U12731 ( .A(n10844), .B(n15065), .ZN(n10849) );
  NAND2_X1 U12732 ( .A1(n15109), .A2(n11123), .ZN(n10846) );
  NAND2_X1 U12733 ( .A1(n10847), .A2(n10846), .ZN(n10848) );
  NOR2_X1 U12734 ( .A1(n10849), .A2(n10848), .ZN(n10853) );
  AOI21_X1 U12735 ( .B1(n10849), .B2(n10848), .A(n10853), .ZN(n15106) );
  INV_X1 U12736 ( .A(n10852), .ZN(n15107) );
  NAND2_X1 U12737 ( .A1(n15106), .A2(n15107), .ZN(n15105) );
  INV_X1 U12738 ( .A(n10853), .ZN(n10854) );
  NAND2_X1 U12739 ( .A1(n15105), .A2(n10854), .ZN(n15178) );
  OAI22_X1 U12740 ( .A1(n10864), .A2(n15094), .B1(n12749), .B2(n15095), .ZN(
        n10857) );
  OAI22_X1 U12741 ( .A1(n10864), .A2(n15095), .B1(n12749), .B2(n15096), .ZN(
        n10855) );
  XNOR2_X1 U12742 ( .A(n10855), .B(n15065), .ZN(n10856) );
  XOR2_X1 U12743 ( .A(n10857), .B(n10856), .Z(n15179) );
  NAND2_X1 U12744 ( .A1(n15178), .A2(n15179), .ZN(n15177) );
  NAND2_X1 U12745 ( .A1(n15177), .A2(n10858), .ZN(n10859) );
  AOI211_X1 U12746 ( .C1(n10860), .C2(n10859), .A(n15205), .B(n11128), .ZN(
        n10866) );
  NAND2_X1 U12747 ( .A1(n15159), .A2(n15500), .ZN(n15191) );
  NAND2_X1 U12748 ( .A1(n15159), .A2(n15437), .ZN(n15193) );
  INV_X1 U12749 ( .A(n15193), .ZN(n15182) );
  AOI22_X1 U12750 ( .A1(n15182), .A2(n15234), .B1(n15196), .B2(n12757), .ZN(
        n10863) );
  MUX2_X1 U12751 ( .A(n15192), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n10862) );
  OAI211_X1 U12752 ( .C1(n10864), .C2(n15191), .A(n10863), .B(n10862), .ZN(
        n10865) );
  OR2_X1 U12753 ( .A1(n10866), .A2(n10865), .ZN(P1_U3218) );
  INV_X1 U12754 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n14804) );
  INV_X1 U12755 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10888) );
  INV_X1 U12756 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10884) );
  INV_X1 U12757 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10867) );
  MUX2_X1 U12758 ( .A(n10867), .B(P2_REG2_REG_4__SCAN_IN), .S(n14521), .Z(
        n10874) );
  INV_X1 U12759 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11721) );
  XNOR2_X1 U12760 ( .A(n11271), .B(n11721), .ZN(n11268) );
  AND2_X1 U12761 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10868) );
  NAND2_X1 U12762 ( .A1(n14488), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10869) );
  OAI211_X1 U12763 ( .C1(n14488), .C2(P2_REG2_REG_1__SCAN_IN), .A(n10868), .B(
        n10869), .ZN(n14493) );
  NAND2_X1 U12764 ( .A1(n14493), .A2(n10869), .ZN(n11269) );
  NAND2_X1 U12765 ( .A1(n11268), .A2(n11269), .ZN(n10871) );
  NAND2_X1 U12766 ( .A1(n11271), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10870) );
  NAND2_X1 U12767 ( .A1(n10871), .A2(n10870), .ZN(n14502) );
  INV_X1 U12768 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10872) );
  MUX2_X1 U12769 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10872), .S(n14504), .Z(
        n14503) );
  NAND2_X1 U12770 ( .A1(n14502), .A2(n14503), .ZN(n14517) );
  NAND2_X1 U12771 ( .A1(n14504), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n14516) );
  NAND2_X1 U12772 ( .A1(n14517), .A2(n14516), .ZN(n10873) );
  NAND2_X1 U12773 ( .A1(n10874), .A2(n10873), .ZN(n14520) );
  NAND2_X1 U12774 ( .A1(n14515), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10875) );
  NAND2_X1 U12775 ( .A1(n14520), .A2(n10875), .ZN(n15832) );
  INV_X1 U12776 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10876) );
  MUX2_X1 U12777 ( .A(n10876), .B(P2_REG2_REG_5__SCAN_IN), .S(n10911), .Z(
        n15831) );
  NAND2_X1 U12778 ( .A1(n15832), .A2(n15831), .ZN(n15830) );
  INV_X1 U12779 ( .A(n10911), .ZN(n15822) );
  NAND2_X1 U12780 ( .A1(n15822), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n14531) );
  NAND2_X1 U12781 ( .A1(n15830), .A2(n14531), .ZN(n10878) );
  INV_X1 U12782 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11549) );
  MUX2_X1 U12783 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11549), .S(n14539), .Z(
        n10877) );
  NAND2_X1 U12784 ( .A1(n10878), .A2(n10877), .ZN(n14533) );
  NAND2_X1 U12785 ( .A1(n14539), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n11168) );
  NAND2_X1 U12786 ( .A1(n14533), .A2(n11168), .ZN(n10881) );
  INV_X1 U12787 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10879) );
  MUX2_X1 U12788 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10879), .S(n11166), .Z(
        n10880) );
  NAND2_X1 U12789 ( .A1(n10881), .A2(n10880), .ZN(n11170) );
  NAND2_X1 U12790 ( .A1(n11166), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U12791 ( .A1(n11170), .A2(n10882), .ZN(n11148) );
  INV_X1 U12792 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11897) );
  MUX2_X1 U12793 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11897), .S(n10920), .Z(
        n11147) );
  NAND2_X1 U12794 ( .A1(n11148), .A2(n11147), .ZN(n11146) );
  NAND2_X1 U12795 ( .A1(n10920), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U12796 ( .A1(n11146), .A2(n10883), .ZN(n15894) );
  MUX2_X1 U12797 ( .A(n10884), .B(P2_REG2_REG_9__SCAN_IN), .S(n15891), .Z(
        n15893) );
  OR2_X1 U12798 ( .A1(n15894), .A2(n15893), .ZN(n15896) );
  OAI21_X1 U12799 ( .B1(n15891), .B2(P2_REG2_REG_9__SCAN_IN), .A(n15896), .ZN(
        n11156) );
  INV_X1 U12800 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10885) );
  MUX2_X1 U12801 ( .A(n10885), .B(P2_REG2_REG_10__SCAN_IN), .S(n10924), .Z(
        n11155) );
  NOR2_X1 U12802 ( .A1(n11156), .A2(n11155), .ZN(n11154) );
  AOI21_X1 U12803 ( .B1(n10924), .B2(P2_REG2_REG_10__SCAN_IN), .A(n11154), 
        .ZN(n10963) );
  INV_X1 U12804 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10886) );
  MUX2_X1 U12805 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10886), .S(n10970), .Z(
        n10964) );
  NAND2_X1 U12806 ( .A1(n10963), .A2(n10964), .ZN(n15878) );
  NAND2_X1 U12807 ( .A1(n10887), .A2(n10886), .ZN(n15876) );
  MUX2_X1 U12808 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10888), .S(n10926), .Z(
        n15877) );
  AOI21_X1 U12809 ( .B1(n15878), .B2(n15876), .A(n15877), .ZN(n15875) );
  AOI21_X1 U12810 ( .B1(n10888), .B2(n10926), .A(n15875), .ZN(n11370) );
  NAND2_X1 U12811 ( .A1(n11380), .A2(n14804), .ZN(n10889) );
  OAI211_X1 U12812 ( .C1(n14804), .C2(n11380), .A(n11370), .B(n10889), .ZN(
        n11368) );
  OAI21_X1 U12813 ( .B1(n14804), .B2(n11380), .A(n11368), .ZN(n10893) );
  INV_X1 U12814 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10891) );
  NOR2_X1 U12815 ( .A1(n10901), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11850) );
  INV_X1 U12816 ( .A(n11850), .ZN(n10890) );
  OAI21_X1 U12817 ( .B1(n10891), .B2(n11861), .A(n10890), .ZN(n10892) );
  NOR2_X1 U12818 ( .A1(n10892), .A2(n10893), .ZN(n11849) );
  AOI21_X1 U12819 ( .B1(n10893), .B2(n10892), .A(n11849), .ZN(n10938) );
  INV_X1 U12820 ( .A(n10894), .ZN(n10899) );
  NAND2_X1 U12821 ( .A1(n10896), .A2(n10895), .ZN(n10897) );
  NAND2_X1 U12822 ( .A1(n10897), .A2(n8629), .ZN(n10898) );
  NAND2_X1 U12823 ( .A1(n10899), .A2(n10898), .ZN(n10933) );
  NOR2_X1 U12824 ( .A1(n9064), .A2(P2_U3088), .ZN(n14960) );
  AND2_X1 U12825 ( .A1(n10933), .A2(n14960), .ZN(n10929) );
  AND2_X1 U12826 ( .A1(n10929), .A2(n10900), .ZN(n15898) );
  XNOR2_X1 U12827 ( .A(n10901), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11862) );
  INV_X1 U12828 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11945) );
  INV_X1 U12829 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10902) );
  MUX2_X1 U12830 ( .A(n10902), .B(P2_REG1_REG_4__SCAN_IN), .S(n14521), .Z(
        n10909) );
  INV_X1 U12831 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n11272) );
  MUX2_X1 U12832 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n11272), .S(n11271), .Z(
        n10904) );
  INV_X1 U12833 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n11400) );
  XNOR2_X1 U12834 ( .A(n14488), .B(n11400), .ZN(n14496) );
  AND2_X1 U12835 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14495) );
  NAND2_X1 U12836 ( .A1(n14496), .A2(n14495), .ZN(n14494) );
  NAND2_X1 U12837 ( .A1(n14488), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U12838 ( .A1(n14494), .A2(n10903), .ZN(n11270) );
  NAND2_X1 U12839 ( .A1(n10904), .A2(n11270), .ZN(n14507) );
  NAND2_X1 U12840 ( .A1(n11271), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n14505) );
  NAND2_X1 U12841 ( .A1(n14507), .A2(n14505), .ZN(n10907) );
  INV_X1 U12842 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10905) );
  MUX2_X1 U12843 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10905), .S(n14504), .Z(
        n10906) );
  NAND2_X1 U12844 ( .A1(n10907), .A2(n10906), .ZN(n14523) );
  NAND2_X1 U12845 ( .A1(n14504), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n14522) );
  NAND2_X1 U12846 ( .A1(n14523), .A2(n14522), .ZN(n10908) );
  NAND2_X1 U12847 ( .A1(n10909), .A2(n10908), .ZN(n14526) );
  NAND2_X1 U12848 ( .A1(n14515), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10910) );
  NAND2_X1 U12849 ( .A1(n14526), .A2(n10910), .ZN(n15828) );
  INV_X1 U12850 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10912) );
  MUX2_X1 U12851 ( .A(n10912), .B(P2_REG1_REG_5__SCAN_IN), .S(n10911), .Z(
        n15829) );
  NAND2_X1 U12852 ( .A1(n15828), .A2(n15829), .ZN(n15827) );
  NAND2_X1 U12853 ( .A1(n15822), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n14535) );
  NAND2_X1 U12854 ( .A1(n15827), .A2(n14535), .ZN(n10915) );
  INV_X1 U12855 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10913) );
  MUX2_X1 U12856 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10913), .S(n14539), .Z(
        n10914) );
  NAND2_X1 U12857 ( .A1(n10915), .A2(n10914), .ZN(n14537) );
  NAND2_X1 U12858 ( .A1(n14539), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10916) );
  NAND2_X1 U12859 ( .A1(n14537), .A2(n10916), .ZN(n11172) );
  INV_X1 U12860 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10917) );
  MUX2_X1 U12861 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10917), .S(n11166), .Z(
        n11173) );
  NAND2_X1 U12862 ( .A1(n11172), .A2(n11173), .ZN(n11171) );
  NAND2_X1 U12863 ( .A1(n11166), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10918) );
  NAND2_X1 U12864 ( .A1(n11171), .A2(n10918), .ZN(n11144) );
  INV_X1 U12865 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10919) );
  MUX2_X1 U12866 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10919), .S(n10920), .Z(
        n11145) );
  NAND2_X1 U12867 ( .A1(n11144), .A2(n11145), .ZN(n11143) );
  NAND2_X1 U12868 ( .A1(n10920), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10921) );
  NAND2_X1 U12869 ( .A1(n11143), .A2(n10921), .ZN(n15887) );
  MUX2_X1 U12870 ( .A(n11945), .B(P2_REG1_REG_9__SCAN_IN), .S(n15891), .Z(
        n15886) );
  NOR2_X1 U12871 ( .A1(n15887), .A2(n15886), .ZN(n15890) );
  AOI21_X1 U12872 ( .B1(n11945), .B2(n10922), .A(n15890), .ZN(n11160) );
  INV_X1 U12873 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10923) );
  MUX2_X1 U12874 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10923), .S(n10924), .Z(
        n11159) );
  NAND2_X1 U12875 ( .A1(n11160), .A2(n11159), .ZN(n11158) );
  NAND2_X1 U12876 ( .A1(n10924), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10960) );
  INV_X1 U12877 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10925) );
  MUX2_X1 U12878 ( .A(n10925), .B(P2_REG1_REG_11__SCAN_IN), .S(n10970), .Z(
        n10959) );
  AOI21_X1 U12879 ( .B1(n11158), .B2(n10960), .A(n10959), .ZN(n10973) );
  AOI21_X1 U12880 ( .B1(n10970), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10973), 
        .ZN(n15874) );
  INV_X1 U12881 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n16207) );
  MUX2_X1 U12882 ( .A(n16207), .B(P2_REG1_REG_12__SCAN_IN), .S(n10926), .Z(
        n15873) );
  NAND2_X1 U12883 ( .A1(n15874), .A2(n15873), .ZN(n15872) );
  OAI21_X1 U12884 ( .B1(n15882), .B2(P2_REG1_REG_12__SCAN_IN), .A(n15872), 
        .ZN(n11373) );
  OR2_X1 U12885 ( .A1(n11367), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10928) );
  NAND2_X1 U12886 ( .A1(n11367), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10927) );
  NAND2_X1 U12887 ( .A1(n10928), .A2(n10927), .ZN(n11374) );
  NOR2_X1 U12888 ( .A1(n11373), .A2(n11374), .ZN(n11372) );
  AOI21_X1 U12889 ( .B1(n11367), .B2(P2_REG1_REG_13__SCAN_IN), .A(n11372), 
        .ZN(n11863) );
  XOR2_X1 U12890 ( .A(n11862), .B(n11863), .Z(n10930) );
  NAND2_X1 U12891 ( .A1(n10930), .A2(n15888), .ZN(n10937) );
  INV_X1 U12892 ( .A(n15904), .ZN(n15858) );
  NOR2_X1 U12893 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10931), .ZN(n10935) );
  AND2_X1 U12894 ( .A1(n9064), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10932) );
  INV_X1 U12895 ( .A(n15892), .ZN(n15837) );
  NOR2_X1 U12896 ( .A1(n15837), .A2(n11861), .ZN(n10934) );
  AOI211_X1 U12897 ( .C1(n15858), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n10935), 
        .B(n10934), .ZN(n10936) );
  OAI211_X1 U12898 ( .C1(n10938), .C2(n15859), .A(n10937), .B(n10936), .ZN(
        P2_U3228) );
  INV_X1 U12899 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10939) );
  MUX2_X1 U12900 ( .A(n10939), .B(P1_REG1_REG_13__SCAN_IN), .S(n12193), .Z(
        n10943) );
  NOR2_X1 U12901 ( .A1(n12075), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n15921) );
  INV_X1 U12902 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10940) );
  MUX2_X1 U12903 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10940), .S(n15930), .Z(
        n10941) );
  NOR2_X1 U12904 ( .A1(n10942), .A2(n10943), .ZN(n11286) );
  AOI211_X1 U12905 ( .C1(n10943), .C2(n10942), .A(n12275), .B(n11286), .ZN(
        n10955) );
  AOI21_X1 U12906 ( .B1(n12075), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10944), 
        .ZN(n15919) );
  INV_X1 U12907 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10945) );
  MUX2_X1 U12908 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10945), .S(n15930), .Z(
        n15920) );
  NAND2_X1 U12909 ( .A1(n15919), .A2(n15920), .ZN(n15918) );
  OAI21_X1 U12910 ( .B1(n15930), .B2(P1_REG2_REG_12__SCAN_IN), .A(n15918), 
        .ZN(n10949) );
  INV_X1 U12911 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10946) );
  MUX2_X1 U12912 ( .A(n10946), .B(P1_REG2_REG_13__SCAN_IN), .S(n12193), .Z(
        n10948) );
  OR2_X1 U12913 ( .A1(n10949), .A2(n10948), .ZN(n11284) );
  INV_X1 U12914 ( .A(n11284), .ZN(n10947) );
  AOI211_X1 U12915 ( .C1(n10949), .C2(n10948), .A(n15338), .B(n10947), .ZN(
        n10954) );
  NOR2_X1 U12916 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12197), .ZN(n10950) );
  AOI21_X1 U12917 ( .B1(n15914), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10950), 
        .ZN(n10951) );
  OAI21_X1 U12918 ( .B1(n15337), .B2(n10952), .A(n10951), .ZN(n10953) );
  OR3_X1 U12919 ( .A1(n10955), .A2(n10954), .A3(n10953), .ZN(P1_U3256) );
  OAI222_X1 U12920 ( .A1(n12396), .A2(n10958), .B1(n14252), .B2(n10957), .C1(
        P3_U3151), .C2(n10956), .ZN(P3_U3274) );
  NAND3_X1 U12921 ( .A1(n11158), .A2(n10960), .A3(n10959), .ZN(n10961) );
  NAND2_X1 U12922 ( .A1(n10961), .A2(n15888), .ZN(n10972) );
  INV_X1 U12923 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U12924 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12269)
         );
  OAI21_X1 U12925 ( .B1(n15904), .B2(n10962), .A(n12269), .ZN(n10969) );
  INV_X1 U12926 ( .A(n10963), .ZN(n10966) );
  INV_X1 U12927 ( .A(n10964), .ZN(n10965) );
  NAND2_X1 U12928 ( .A1(n10966), .A2(n10965), .ZN(n10967) );
  AOI21_X1 U12929 ( .B1(n10967), .B2(n15878), .A(n15859), .ZN(n10968) );
  AOI211_X1 U12930 ( .C1(n15892), .C2(n10970), .A(n10969), .B(n10968), .ZN(
        n10971) );
  OAI21_X1 U12931 ( .B1(n10973), .B2(n10972), .A(n10971), .ZN(P2_U3225) );
  INV_X1 U12932 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11720) );
  INV_X1 U12933 ( .A(n11678), .ZN(n14350) );
  AND2_X1 U12934 ( .A1(n14483), .A2(n14350), .ZN(n10978) );
  AND2_X1 U12935 ( .A1(n10974), .A2(n10115), .ZN(n10975) );
  OR2_X4 U12936 ( .A1(n10976), .A2(n10975), .ZN(n14352) );
  XNOR2_X1 U12937 ( .A(n11724), .B(n14352), .ZN(n10977) );
  NOR2_X1 U12938 ( .A1(n10978), .A2(n10977), .ZN(n11082) );
  AOI21_X1 U12939 ( .B1(n10978), .B2(n10977), .A(n11082), .ZN(n10987) );
  AOI22_X1 U12940 ( .A1(n11391), .A2(n14350), .B1(n14304), .B2(n10979), .ZN(
        n11223) );
  NAND2_X1 U12941 ( .A1(n11223), .A2(n11222), .ZN(n11221) );
  INV_X1 U12942 ( .A(n10984), .ZN(n10985) );
  NAND2_X1 U12943 ( .A1(n11221), .A2(n10985), .ZN(n10986) );
  NAND2_X1 U12944 ( .A1(n10986), .A2(n10987), .ZN(n11084) );
  OAI21_X1 U12945 ( .B1(n10987), .B2(n10986), .A(n11084), .ZN(n10988) );
  NAND2_X1 U12946 ( .A1(n10988), .A2(n14420), .ZN(n10992) );
  NAND2_X1 U12947 ( .A1(n14482), .A2(n14791), .ZN(n10990) );
  NAND2_X1 U12948 ( .A1(n14484), .A2(n14647), .ZN(n10989) );
  NAND2_X1 U12949 ( .A1(n10990), .A2(n10989), .ZN(n11409) );
  AOI22_X1 U12950 ( .A1(n11724), .A2(n14423), .B1(n14392), .B2(n11409), .ZN(
        n10991) );
  OAI211_X1 U12951 ( .C1(n11227), .C2(n11720), .A(n10992), .B(n10991), .ZN(
        P2_U3209) );
  XNOR2_X1 U12952 ( .A(n10993), .B(n10994), .ZN(n16063) );
  XNOR2_X1 U12953 ( .A(n10995), .B(n10994), .ZN(n10998) );
  NAND2_X1 U12954 ( .A1(n14481), .A2(n14791), .ZN(n10997) );
  NAND2_X1 U12955 ( .A1(n14483), .A2(n14647), .ZN(n10996) );
  NAND2_X1 U12956 ( .A1(n10997), .A2(n10996), .ZN(n11109) );
  AOI21_X1 U12957 ( .B1(n10998), .B2(n9112), .A(n11109), .ZN(n16068) );
  INV_X1 U12958 ( .A(n11594), .ZN(n10999) );
  AOI211_X1 U12959 ( .C1(n9900), .C2(n11411), .A(n14300), .B(n10999), .ZN(
        n16066) );
  AOI21_X1 U12960 ( .B1(n16134), .B2(n9900), .A(n16066), .ZN(n11000) );
  OAI211_X1 U12961 ( .C1(n16138), .C2(n16063), .A(n16068), .B(n11000), .ZN(
        n11769) );
  NAND2_X1 U12962 ( .A1(n11769), .A2(n16208), .ZN(n11001) );
  OAI21_X1 U12963 ( .B1(n16208), .B2(n10905), .A(n11001), .ZN(P2_U3502) );
  INV_X1 U12964 ( .A(n11002), .ZN(n11004) );
  NAND2_X1 U12965 ( .A1(n11004), .A2(n11003), .ZN(n11005) );
  MUX2_X1 U12966 ( .A(n11007), .B(n16146), .S(n13309), .Z(n11009) );
  INV_X1 U12967 ( .A(n11009), .ZN(n11008) );
  NAND2_X1 U12968 ( .A1(n11008), .A2(n11019), .ZN(n11568) );
  INV_X1 U12969 ( .A(n11568), .ZN(n11010) );
  AND2_X1 U12970 ( .A1(n11009), .A2(n11575), .ZN(n11566) );
  NOR2_X1 U12971 ( .A1(n11010), .A2(n11566), .ZN(n11011) );
  XNOR2_X1 U12972 ( .A(n11567), .B(n11011), .ZN(n11026) );
  INV_X1 U12973 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n16146) );
  NAND2_X1 U12974 ( .A1(n11016), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11012) );
  AND2_X2 U12975 ( .A1(n11013), .A2(n11012), .ZN(n11558) );
  AOI21_X1 U12976 ( .B1(n16146), .B2(n11014), .A(n11559), .ZN(n11015) );
  NOR2_X1 U12977 ( .A1(n11015), .A2(n13899), .ZN(n11025) );
  NAND2_X1 U12978 ( .A1(n11016), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11017) );
  AOI21_X1 U12979 ( .B1(n11007), .B2(n11020), .A(n11576), .ZN(n11023) );
  NOR2_X1 U12980 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9349), .ZN(n12129) );
  AOI21_X1 U12981 ( .B1(n15817), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12129), .ZN(
        n11022) );
  NAND2_X1 U12982 ( .A1(n13874), .A2(n11575), .ZN(n11021) );
  OAI211_X1 U12983 ( .C1(n11023), .C2(n13895), .A(n11022), .B(n11021), .ZN(
        n11024) );
  AOI211_X1 U12984 ( .C1(n11026), .C2(n13897), .A(n11025), .B(n11024), .ZN(
        n11027) );
  INV_X1 U12985 ( .A(n11027), .ZN(P3_U3191) );
  OAI21_X1 U12986 ( .B1(n11029), .B2(n13265), .A(n11028), .ZN(n11591) );
  OAI211_X1 U12987 ( .C1(n11032), .C2(n11031), .A(n11030), .B(n14103), .ZN(
        n11034) );
  AOI22_X1 U12988 ( .A1(n14108), .A2(n13522), .B1(n13520), .B2(n14107), .ZN(
        n11033) );
  NAND2_X1 U12989 ( .A1(n11034), .A2(n11033), .ZN(n11588) );
  AOI21_X1 U12990 ( .B1(n16226), .B2(n11591), .A(n11588), .ZN(n11040) );
  INV_X1 U12991 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n11035) );
  OAI22_X1 U12992 ( .A1(n14246), .A2(n13111), .B1(n16232), .B2(n11035), .ZN(
        n11036) );
  INV_X1 U12993 ( .A(n11036), .ZN(n11037) );
  OAI21_X1 U12994 ( .B1(n11040), .B2(n16229), .A(n11037), .ZN(P3_U3402) );
  OAI22_X1 U12995 ( .A1(n14192), .A2(n13111), .B1(n16228), .B2(n10518), .ZN(
        n11038) );
  INV_X1 U12996 ( .A(n11038), .ZN(n11039) );
  OAI21_X1 U12997 ( .B1(n11040), .B2(n7687), .A(n11039), .ZN(P3_U3463) );
  OAI22_X1 U12998 ( .A1(n13313), .A2(P3_U3151), .B1(SI_22_), .B2(n14252), .ZN(
        n11041) );
  AOI21_X1 U12999 ( .B1(n11042), .B2(n14257), .A(n11041), .ZN(P3_U3273) );
  NAND4_X1 U13000 ( .A1(n13061), .A2(n11045), .A3(n11044), .A4(n11043), .ZN(
        n15387) );
  NAND2_X1 U13001 ( .A1(n12742), .A2(n12730), .ZN(n12996) );
  INV_X1 U13002 ( .A(n15598), .ZN(n16018) );
  OR2_X1 U13003 ( .A1(n15387), .A2(n12730), .ZN(n15363) );
  NOR2_X2 U13004 ( .A1(n15363), .A2(n16096), .ZN(n15601) );
  INV_X1 U13005 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11047) );
  OAI22_X1 U13006 ( .A1(n15611), .A2(n10280), .B1(n11047), .B2(n15615), .ZN(
        n11048) );
  AOI21_X1 U13007 ( .B1(n15601), .B2(n11049), .A(n11048), .ZN(n11050) );
  OAI21_X1 U13008 ( .B1(n12749), .B2(n16014), .A(n11050), .ZN(n11051) );
  AOI21_X1 U13009 ( .B1(n16018), .B2(n11052), .A(n11051), .ZN(n11053) );
  OAI21_X1 U13010 ( .B1(n11054), .B2(n16022), .A(n11053), .ZN(P1_U3291) );
  INV_X1 U13011 ( .A(n11055), .ZN(n11056) );
  OAI21_X1 U13012 ( .B1(n11056), .B2(n14248), .A(n11059), .ZN(n11057) );
  OAI211_X1 U13013 ( .C1(n14248), .C2(n11059), .A(n11058), .B(n11057), .ZN(
        n11061) );
  MUX2_X1 U13014 ( .A(n11060), .B(P3_REG2_REG_0__SCAN_IN), .S(n16052), .Z(
        n11066) );
  INV_X1 U13015 ( .A(n11061), .ZN(n11063) );
  NOR2_X1 U13016 ( .A1(n16222), .A2(n16045), .ZN(n11062) );
  OAI22_X1 U13017 ( .A1(n16126), .A2(n11064), .B1(n10470), .B2(n16128), .ZN(
        n11065) );
  OR2_X1 U13018 ( .A1(n11066), .A2(n11065), .ZN(P3_U3233) );
  MUX2_X1 U13019 ( .A(n11068), .B(n11067), .S(n15611), .Z(n11072) );
  OAI22_X1 U13020 ( .A1(n16014), .A2(n8021), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n15615), .ZN(n11069) );
  AOI21_X1 U13021 ( .B1(n11070), .B2(n15601), .A(n11069), .ZN(n11071) );
  OAI211_X1 U13022 ( .C1(n11073), .C2(n15577), .A(n11072), .B(n11071), .ZN(
        P1_U3290) );
  INV_X1 U13023 ( .A(n11074), .ZN(n11079) );
  INV_X1 U13024 ( .A(n15363), .ZN(n15429) );
  INV_X1 U13025 ( .A(n15615), .ZN(n16011) );
  AOI22_X1 U13026 ( .A1(n15429), .A2(n11075), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n16011), .ZN(n11077) );
  NAND2_X1 U13027 ( .A1(n16022), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n11076) );
  OAI211_X1 U13028 ( .C1(n12737), .C2(n16014), .A(n11077), .B(n11076), .ZN(
        n11078) );
  AOI21_X1 U13029 ( .B1(n11079), .B2(n16018), .A(n11078), .ZN(n11080) );
  OAI21_X1 U13030 ( .B1(n11081), .B2(n16022), .A(n11080), .ZN(P1_U3292) );
  INV_X1 U13031 ( .A(n11082), .ZN(n11083) );
  NAND2_X1 U13032 ( .A1(n11084), .A2(n11083), .ZN(n11113) );
  XOR2_X1 U13033 ( .A(n14352), .B(n9900), .Z(n11086) );
  INV_X2 U13034 ( .A(n11678), .ZN(n14300) );
  NAND2_X1 U13035 ( .A1(n14482), .A2(n14300), .ZN(n11085) );
  XNOR2_X1 U13036 ( .A(n11086), .B(n11085), .ZN(n11112) );
  NAND2_X1 U13037 ( .A1(n14481), .A2(n14300), .ZN(n11087) );
  NAND2_X1 U13038 ( .A1(n11088), .A2(n11087), .ZN(n11253) );
  OAI21_X1 U13039 ( .B1(n11088), .B2(n11087), .A(n11253), .ZN(n11089) );
  AOI21_X1 U13040 ( .B1(n11090), .B2(n11089), .A(n11255), .ZN(n11097) );
  NAND2_X1 U13041 ( .A1(n14480), .A2(n14791), .ZN(n11093) );
  NAND2_X1 U13042 ( .A1(n14482), .A2(n14647), .ZN(n11092) );
  NAND2_X1 U13043 ( .A1(n11093), .A2(n11092), .ZN(n11600) );
  NAND2_X1 U13044 ( .A1(n14392), .A2(n11600), .ZN(n11094) );
  NAND2_X1 U13045 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n14512) );
  OAI211_X1 U13046 ( .C1(n14462), .C2(n16084), .A(n11094), .B(n14512), .ZN(
        n11095) );
  AOI21_X1 U13047 ( .B1(n16081), .B2(n14459), .A(n11095), .ZN(n11096) );
  OAI21_X1 U13048 ( .B1(n11097), .B2(n14449), .A(n11096), .ZN(P2_U3202) );
  XNOR2_X1 U13049 ( .A(n13111), .B(n11099), .ZN(n11100) );
  NOR2_X1 U13050 ( .A1(n11100), .A2(n13521), .ZN(n11297) );
  AOI21_X1 U13051 ( .B1(n13521), .B2(n11100), .A(n11297), .ZN(n11101) );
  OAI21_X1 U13052 ( .B1(n11102), .B2(n11101), .A(n11299), .ZN(n11103) );
  NAND2_X1 U13053 ( .A1(n11103), .A2(n13495), .ZN(n11108) );
  NOR2_X1 U13054 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11104), .ZN(n13751) );
  OAI22_X1 U13055 ( .A1(n16033), .A2(n13500), .B1(n7795), .B2(n13470), .ZN(
        n11105) );
  AOI211_X1 U13056 ( .C1(n11106), .C2(n13411), .A(n13751), .B(n11105), .ZN(
        n11107) );
  OAI211_X1 U13057 ( .C1(n11587), .C2(n12627), .A(n11108), .B(n11107), .ZN(
        P3_U3170) );
  NAND2_X1 U13058 ( .A1(n14423), .A2(n9900), .ZN(n11111) );
  NAND2_X1 U13059 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n14500) );
  NAND2_X1 U13060 ( .A1(n14392), .A2(n11109), .ZN(n11110) );
  NAND3_X1 U13061 ( .A1(n11111), .A2(n14500), .A3(n11110), .ZN(n11116) );
  XNOR2_X1 U13062 ( .A(n11113), .B(n11112), .ZN(n11114) );
  NOR2_X1 U13063 ( .A1(n11114), .A2(n14449), .ZN(n11115) );
  AOI211_X1 U13064 ( .C1(n14459), .C2(n16060), .A(n11116), .B(n11115), .ZN(
        n11117) );
  INV_X1 U13065 ( .A(n11117), .ZN(P2_U3190) );
  NAND2_X1 U13066 ( .A1(n15234), .A2(n15050), .ZN(n11125) );
  AOI22_X1 U13067 ( .A1(n12836), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n12835), 
        .B2(n11120), .ZN(n11121) );
  NAND2_X1 U13068 ( .A1(n12762), .A2(n11123), .ZN(n11124) );
  NAND2_X1 U13069 ( .A1(n11125), .A2(n11124), .ZN(n11126) );
  NAND2_X1 U13070 ( .A1(n7355), .A2(n11188), .ZN(n11130) );
  OAI22_X1 U13071 ( .A1(n11239), .A2(n15095), .B1(n16070), .B2(n15096), .ZN(
        n11129) );
  XOR2_X1 U13072 ( .A(n15065), .B(n11129), .Z(n11189) );
  XNOR2_X1 U13073 ( .A(n11130), .B(n11189), .ZN(n11142) );
  NAND2_X1 U13074 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(n7190), .ZN(n15278) );
  OAI21_X1 U13075 ( .B1(n15220), .B2(n16070), .A(n15278), .ZN(n11140) );
  NAND2_X1 U13076 ( .A1(n12875), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n11138) );
  NAND2_X1 U13077 ( .A1(n12966), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n11137) );
  NAND2_X1 U13078 ( .A1(n11131), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n11202) );
  INV_X1 U13079 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U13080 ( .A1(n11133), .A2(n11132), .ZN(n11134) );
  AND2_X1 U13081 ( .A1(n11202), .A2(n11134), .ZN(n11246) );
  NAND2_X1 U13082 ( .A1(n12965), .A2(n11246), .ZN(n11136) );
  INV_X1 U13083 ( .A(n15233), .ZN(n11337) );
  OAI22_X1 U13084 ( .A1(n11233), .A2(n15191), .B1(n15193), .B2(n11337), .ZN(
        n11139) );
  AOI211_X1 U13085 ( .C1(n11359), .C2(n15216), .A(n11140), .B(n11139), .ZN(
        n11141) );
  OAI21_X1 U13086 ( .B1(n11142), .B2(n15205), .A(n11141), .ZN(P1_U3230) );
  OAI211_X1 U13087 ( .C1(n11145), .C2(n11144), .A(n15888), .B(n11143), .ZN(
        n11150) );
  OAI211_X1 U13088 ( .C1(n11148), .C2(n11147), .A(n15898), .B(n11146), .ZN(
        n11149) );
  NAND2_X1 U13089 ( .A1(n11150), .A2(n11149), .ZN(n11151) );
  AND2_X1 U13090 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11886) );
  AOI211_X1 U13091 ( .C1(n15858), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n11151), .B(
        n11886), .ZN(n11152) );
  OAI21_X1 U13092 ( .B1(n11153), .B2(n15837), .A(n11152), .ZN(P2_U3222) );
  AOI211_X1 U13093 ( .C1(n11156), .C2(n11155), .A(n11154), .B(n15859), .ZN(
        n11157) );
  INV_X1 U13094 ( .A(n11157), .ZN(n11164) );
  NAND2_X1 U13095 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n12232)
         );
  OAI211_X1 U13096 ( .C1(n11160), .C2(n11159), .A(n15888), .B(n11158), .ZN(
        n11161) );
  NAND2_X1 U13097 ( .A1(n12232), .A2(n11161), .ZN(n11162) );
  AOI21_X1 U13098 ( .B1(n15858), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n11162), 
        .ZN(n11163) );
  OAI211_X1 U13099 ( .C1(n15837), .C2(n11165), .A(n11164), .B(n11163), .ZN(
        P2_U3224) );
  MUX2_X1 U13100 ( .A(n10879), .B(P2_REG2_REG_7__SCAN_IN), .S(n11166), .Z(
        n11167) );
  NAND3_X1 U13101 ( .A1(n14533), .A2(n11168), .A3(n11167), .ZN(n11169) );
  NAND3_X1 U13102 ( .A1(n15898), .A2(n11170), .A3(n11169), .ZN(n11177) );
  NAND2_X1 U13103 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11684) );
  OAI211_X1 U13104 ( .C1(n11173), .C2(n11172), .A(n15888), .B(n11171), .ZN(
        n11174) );
  NAND2_X1 U13105 ( .A1(n11684), .A2(n11174), .ZN(n11175) );
  AOI21_X1 U13106 ( .B1(n15858), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n11175), .ZN(
        n11176) );
  OAI211_X1 U13107 ( .C1(n15837), .C2(n11178), .A(n11177), .B(n11176), .ZN(
        P2_U3221) );
  INV_X1 U13108 ( .A(n11864), .ZN(n15836) );
  INV_X1 U13109 ( .A(n12595), .ZN(n11187) );
  OAI222_X1 U13110 ( .A1(P2_U3088), .A2(n15836), .B1(n14968), .B2(n11187), 
        .C1(n11179), .C2(n14970), .ZN(P2_U3312) );
  INV_X1 U13111 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n11180) );
  NAND3_X1 U13112 ( .A1(n11182), .A2(n11181), .A3(n11180), .ZN(n11183) );
  OAI21_X1 U13113 ( .B1(n11184), .B2(n11183), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n11185) );
  XNOR2_X1 U13114 ( .A(n11185), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12596) );
  INV_X1 U13115 ( .A(n12596), .ZN(n12001) );
  OAI222_X1 U13116 ( .A1(P1_U3086), .A2(n12001), .B1(n15771), .B2(n11187), 
        .C1(n11186), .C2(n15773), .ZN(P1_U3340) );
  OR2_X1 U13117 ( .A1(n11190), .A2(n12987), .ZN(n11193) );
  AOI22_X1 U13118 ( .A1(n12836), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n12835), 
        .B2(n11191), .ZN(n11192) );
  NAND2_X1 U13119 ( .A1(n12770), .A2(n15062), .ZN(n11195) );
  NAND2_X1 U13120 ( .A1(n15233), .A2(n11123), .ZN(n11194) );
  NAND2_X1 U13121 ( .A1(n11195), .A2(n11194), .ZN(n11196) );
  XNOR2_X1 U13122 ( .A(n11196), .B(n7251), .ZN(n11198) );
  AOI22_X1 U13123 ( .A1(n12770), .A2(n11123), .B1(n15050), .B2(n15233), .ZN(
        n11197) );
  NOR2_X1 U13124 ( .A1(n11198), .A2(n11197), .ZN(n11312) );
  NAND2_X1 U13125 ( .A1(n11198), .A2(n11197), .ZN(n11313) );
  INV_X1 U13126 ( .A(n11313), .ZN(n11199) );
  NOR2_X1 U13127 ( .A1(n11312), .A2(n11199), .ZN(n11200) );
  XNOR2_X1 U13128 ( .A(n11314), .B(n11200), .ZN(n11212) );
  NAND2_X1 U13129 ( .A1(n12875), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n11207) );
  NAND2_X1 U13130 ( .A1(n12966), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n11206) );
  NOR2_X1 U13131 ( .A1(n11202), .A2(n11201), .ZN(n11324) );
  INV_X1 U13132 ( .A(n11324), .ZN(n11326) );
  NAND2_X1 U13133 ( .A1(n11202), .A2(n11201), .ZN(n11203) );
  AND2_X1 U13134 ( .A1(n11326), .A2(n11203), .ZN(n11383) );
  NAND2_X1 U13135 ( .A1(n12965), .A2(n11383), .ZN(n11205) );
  NAND2_X1 U13136 ( .A1(n12982), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n11204) );
  NAND4_X1 U13137 ( .A1(n11207), .A2(n11206), .A3(n11205), .A4(n11204), .ZN(
        n15232) );
  INV_X1 U13138 ( .A(n15232), .ZN(n11531) );
  OAI21_X1 U13139 ( .B1(n15193), .B2(n11531), .A(n11208), .ZN(n11210) );
  OAI22_X1 U13140 ( .A1(n15191), .A2(n11239), .B1(n15220), .B2(n16095), .ZN(
        n11209) );
  AOI211_X1 U13141 ( .C1(n11246), .C2(n15216), .A(n11210), .B(n11209), .ZN(
        n11211) );
  OAI21_X1 U13142 ( .B1(n11212), .B2(n15205), .A(n11211), .ZN(P1_U3227) );
  AOI22_X1 U13143 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n15898), .B1(n15888), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n11218) );
  INV_X1 U13144 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n11213) );
  NAND2_X1 U13145 ( .A1(n15898), .A2(n11213), .ZN(n11216) );
  INV_X1 U13146 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n11214) );
  NAND2_X1 U13147 ( .A1(n15888), .A2(n11214), .ZN(n11215) );
  AND3_X1 U13148 ( .A1(n11216), .A2(n11215), .A3(n15837), .ZN(n11217) );
  MUX2_X1 U13149 ( .A(n11218), .B(n11217), .S(P2_IR_REG_0__SCAN_IN), .Z(n11220) );
  AOI22_X1 U13150 ( .A1(n15858), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n11219) );
  NAND2_X1 U13151 ( .A1(n11220), .A2(n11219), .ZN(P2_U3214) );
  INV_X1 U13152 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n14486) );
  OAI21_X1 U13153 ( .B1(n11223), .B2(n11222), .A(n11221), .ZN(n11224) );
  NAND2_X1 U13154 ( .A1(n14392), .A2(n14791), .ZN(n14404) );
  INV_X1 U13155 ( .A(n14404), .ZN(n14444) );
  AOI22_X1 U13156 ( .A1(n11224), .A2(n14420), .B1(n14444), .B2(n14483), .ZN(
        n11226) );
  NAND2_X1 U13157 ( .A1(n14392), .A2(n14647), .ZN(n14402) );
  INV_X1 U13158 ( .A(n14402), .ZN(n14443) );
  AOI22_X1 U13159 ( .A1(n14443), .A2(n9882), .B1(n7718), .B2(n14423), .ZN(
        n11225) );
  OAI211_X1 U13160 ( .C1(n11227), .C2(n14486), .A(n11226), .B(n11225), .ZN(
        P2_U3194) );
  AOI21_X1 U13161 ( .B1(n14719), .B2(n14876), .A(n11523), .ZN(n11229) );
  NOR2_X1 U13162 ( .A1(n11229), .A2(n11228), .ZN(n11517) );
  NAND2_X1 U13163 ( .A1(n11399), .A2(n11230), .ZN(n11518) );
  NAND2_X1 U13164 ( .A1(n11517), .A2(n11518), .ZN(n11310) );
  NOR2_X1 U13165 ( .A1(n16208), .A2(n11214), .ZN(n11231) );
  AOI21_X1 U13166 ( .B1(n16208), .B2(n11310), .A(n11231), .ZN(n11232) );
  OAI21_X1 U13167 ( .B1(n11523), .B2(n14897), .A(n11232), .ZN(P2_U3499) );
  NAND2_X1 U13168 ( .A1(n11233), .A2(n8021), .ZN(n11234) );
  XNOR2_X1 U13169 ( .A(n11336), .B(n13014), .ZN(n16101) );
  INV_X1 U13170 ( .A(n16101), .ZN(n11252) );
  NOR2_X1 U13171 ( .A1(n15235), .A2(n8021), .ZN(n11237) );
  NAND2_X1 U13172 ( .A1(n15235), .A2(n8021), .ZN(n11236) );
  OAI211_X1 U13173 ( .C1(n11241), .C2(n12767), .A(n11342), .B(n15723), .ZN(
        n11243) );
  AOI22_X1 U13174 ( .A1(n15582), .A2(n15234), .B1(n15232), .B2(n15583), .ZN(
        n11242) );
  NAND2_X1 U13175 ( .A1(n11243), .A2(n11242), .ZN(n11244) );
  AOI21_X1 U13176 ( .B1(n16101), .B2(n15490), .A(n11244), .ZN(n16098) );
  MUX2_X1 U13177 ( .A(n10285), .B(n16098), .S(n15611), .Z(n11251) );
  NOR2_X1 U13178 ( .A1(n11357), .A2(n16095), .ZN(n11245) );
  OR2_X1 U13179 ( .A1(n11348), .A2(n11245), .ZN(n16097) );
  INV_X1 U13180 ( .A(n16097), .ZN(n11249) );
  INV_X1 U13181 ( .A(n11246), .ZN(n11247) );
  OAI22_X1 U13182 ( .A1(n16014), .A2(n16095), .B1(n11247), .B2(n15615), .ZN(
        n11248) );
  AOI21_X1 U13183 ( .B1(n11249), .B2(n15601), .A(n11248), .ZN(n11250) );
  OAI211_X1 U13184 ( .C1(n11252), .C2(n15598), .A(n11251), .B(n11250), .ZN(
        P1_U3288) );
  INV_X1 U13185 ( .A(n11253), .ZN(n11254) );
  NAND2_X1 U13186 ( .A1(n14480), .A2(n14300), .ZN(n11257) );
  XNOR2_X1 U13187 ( .A(n11840), .B(n14304), .ZN(n11256) );
  NAND2_X1 U13188 ( .A1(n11257), .A2(n11256), .ZN(n11503) );
  OAI21_X1 U13189 ( .B1(n11257), .B2(n11256), .A(n11503), .ZN(n11258) );
  AOI21_X1 U13190 ( .B1(n7352), .B2(n11258), .A(n11505), .ZN(n11267) );
  INV_X1 U13191 ( .A(n11839), .ZN(n11264) );
  NAND2_X1 U13192 ( .A1(n14479), .A2(n14791), .ZN(n11260) );
  NAND2_X1 U13193 ( .A1(n14481), .A2(n14647), .ZN(n11259) );
  AND2_X1 U13194 ( .A1(n11260), .A2(n11259), .ZN(n11421) );
  INV_X1 U13195 ( .A(n11421), .ZN(n11261) );
  AND2_X1 U13196 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n15823) );
  AOI21_X1 U13197 ( .B1(n14392), .B2(n11261), .A(n15823), .ZN(n11263) );
  NAND2_X1 U13198 ( .A1(n14423), .A2(n11840), .ZN(n11262) );
  OAI211_X1 U13199 ( .C1(n14403), .C2(n11264), .A(n11263), .B(n11262), .ZN(
        n11265) );
  INV_X1 U13200 ( .A(n11265), .ZN(n11266) );
  OAI21_X1 U13201 ( .B1(n11267), .B2(n14449), .A(n11266), .ZN(P2_U3199) );
  XOR2_X1 U13202 ( .A(n11269), .B(n11268), .Z(n11277) );
  INV_X1 U13203 ( .A(n11270), .ZN(n11275) );
  MUX2_X1 U13204 ( .A(n11272), .B(P2_REG1_REG_2__SCAN_IN), .S(n11271), .Z(
        n11274) );
  INV_X1 U13205 ( .A(n14507), .ZN(n11273) );
  INV_X1 U13206 ( .A(n15888), .ZN(n11371) );
  AOI211_X1 U13207 ( .C1(n11275), .C2(n11274), .A(n11273), .B(n11371), .ZN(
        n11276) );
  AOI21_X1 U13208 ( .B1(n15898), .B2(n11277), .A(n11276), .ZN(n11279) );
  AOI22_X1 U13209 ( .A1(n15858), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n11278) );
  OAI211_X1 U13210 ( .C1(n11280), .C2(n15837), .A(n11279), .B(n11278), .ZN(
        P2_U3216) );
  NAND2_X1 U13211 ( .A1(n12193), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11283) );
  INV_X1 U13212 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11281) );
  MUX2_X1 U13213 ( .A(n11281), .B(P1_REG2_REG_14__SCAN_IN), .S(n12521), .Z(
        n11282) );
  AOI21_X1 U13214 ( .B1(n11284), .B2(n11283), .A(n11282), .ZN(n11732) );
  NAND3_X1 U13215 ( .A1(n11284), .A2(n11283), .A3(n11282), .ZN(n11285) );
  NAND2_X1 U13216 ( .A1(n11285), .A2(n15931), .ZN(n11294) );
  AOI21_X1 U13217 ( .B1(n12193), .B2(P1_REG1_REG_13__SCAN_IN), .A(n11286), 
        .ZN(n11736) );
  INV_X1 U13218 ( .A(n11288), .ZN(n11289) );
  INV_X1 U13219 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11287) );
  OAI211_X1 U13220 ( .C1(n11289), .C2(P1_REG1_REG_14__SCAN_IN), .A(n11734), 
        .B(n15927), .ZN(n11293) );
  NOR2_X1 U13221 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12711), .ZN(n11291) );
  NOR2_X1 U13222 ( .A1(n15337), .A2(n11735), .ZN(n11290) );
  AOI211_X1 U13223 ( .C1(n15914), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n11291), 
        .B(n11290), .ZN(n11292) );
  OAI211_X1 U13224 ( .C1(n11732), .C2(n11294), .A(n11293), .B(n11292), .ZN(
        P1_U3257) );
  NAND2_X1 U13225 ( .A1(n11295), .A2(n14257), .ZN(n11296) );
  OAI211_X1 U13226 ( .C1(n13650), .C2(n14252), .A(n11296), .B(n13315), .ZN(
        P3_U3272) );
  XNOR2_X1 U13227 ( .A(n11305), .B(n13405), .ZN(n11651) );
  XNOR2_X1 U13228 ( .A(n11651), .B(n13520), .ZN(n11301) );
  INV_X1 U13229 ( .A(n11297), .ZN(n11298) );
  OAI21_X1 U13230 ( .B1(n11301), .B2(n11300), .A(n11652), .ZN(n11302) );
  NAND2_X1 U13231 ( .A1(n11302), .A2(n13495), .ZN(n11307) );
  INV_X1 U13232 ( .A(n13519), .ZN(n11795) );
  OAI22_X1 U13233 ( .A1(n7730), .A2(n13500), .B1(n11795), .B2(n13470), .ZN(
        n11303) );
  AOI211_X1 U13234 ( .C1(n11305), .C2(n13411), .A(n11304), .B(n11303), .ZN(
        n11306) );
  OAI211_X1 U13235 ( .C1(n11762), .C2(n12627), .A(n11307), .B(n11306), .ZN(
        P3_U3167) );
  INV_X1 U13236 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n11308) );
  NOR2_X1 U13237 ( .A1(n14948), .A2(n11308), .ZN(n11309) );
  AOI21_X1 U13238 ( .B1(n14948), .B2(n11310), .A(n11309), .ZN(n11311) );
  OAI21_X1 U13239 ( .B1(n11523), .B2(n14953), .A(n11311), .ZN(P2_U3430) );
  NAND2_X1 U13240 ( .A1(n11315), .A2(n12998), .ZN(n11317) );
  AOI22_X1 U13241 ( .A1(n12836), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12835), 
        .B2(n15303), .ZN(n11316) );
  NAND2_X1 U13242 ( .A1(n11317), .A2(n11316), .ZN(n12774) );
  NAND2_X1 U13243 ( .A1(n12774), .A2(n15062), .ZN(n11319) );
  NAND2_X1 U13244 ( .A1(n15232), .A2(n11123), .ZN(n11318) );
  NAND2_X1 U13245 ( .A1(n11319), .A2(n11318), .ZN(n11320) );
  XNOR2_X1 U13246 ( .A(n11320), .B(n15065), .ZN(n11437) );
  NAND2_X1 U13247 ( .A1(n12774), .A2(n11123), .ZN(n11322) );
  NAND2_X1 U13248 ( .A1(n15232), .A2(n15050), .ZN(n11321) );
  NAND2_X1 U13249 ( .A1(n11322), .A2(n11321), .ZN(n11438) );
  XNOR2_X1 U13250 ( .A(n11437), .B(n11438), .ZN(n11323) );
  XNOR2_X1 U13251 ( .A(n11441), .B(n11323), .ZN(n11335) );
  NAND2_X1 U13252 ( .A1(n12966), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U13253 ( .A1(n12982), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U13254 ( .A1(n11324), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11450) );
  INV_X1 U13255 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n11325) );
  NAND2_X1 U13256 ( .A1(n11326), .A2(n11325), .ZN(n11327) );
  AND2_X1 U13257 ( .A1(n11450), .A2(n11327), .ZN(n11540) );
  NAND2_X1 U13258 ( .A1(n12965), .A2(n11540), .ZN(n11329) );
  NAND2_X1 U13259 ( .A1(n12875), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11328) );
  NAND4_X1 U13260 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n15231) );
  INV_X1 U13261 ( .A(n15231), .ZN(n11786) );
  INV_X1 U13262 ( .A(n15191), .ZN(n15184) );
  AOI22_X1 U13263 ( .A1(n15184), .A2(n15233), .B1(n15216), .B2(n11383), .ZN(
        n11332) );
  NAND2_X1 U13264 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n15295) );
  OAI211_X1 U13265 ( .C1(n11786), .C2(n15193), .A(n11332), .B(n15295), .ZN(
        n11333) );
  AOI21_X1 U13266 ( .B1(n12774), .B2(n15196), .A(n11333), .ZN(n11334) );
  OAI21_X1 U13267 ( .B1(n11335), .B2(n15205), .A(n11334), .ZN(P1_U3239) );
  INV_X1 U13268 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11352) );
  NAND2_X1 U13269 ( .A1(n16095), .A2(n11337), .ZN(n11338) );
  NAND2_X1 U13270 ( .A1(n11339), .A2(n11338), .ZN(n11528) );
  XNOR2_X1 U13271 ( .A(n12774), .B(n15232), .ZN(n13016) );
  INV_X1 U13272 ( .A(n13016), .ZN(n11527) );
  XNOR2_X1 U13273 ( .A(n11528), .B(n11527), .ZN(n11340) );
  INV_X1 U13274 ( .A(n11340), .ZN(n11390) );
  NAND2_X1 U13275 ( .A1(n11340), .A2(n15490), .ZN(n11347) );
  NAND2_X1 U13276 ( .A1(n16095), .A2(n15233), .ZN(n11341) );
  NAND2_X1 U13277 ( .A1(n11343), .A2(n13016), .ZN(n11533) );
  OAI211_X1 U13278 ( .C1(n11343), .C2(n13016), .A(n11533), .B(n15723), .ZN(
        n11345) );
  AOI22_X1 U13279 ( .A1(n15582), .A2(n15233), .B1(n15231), .B2(n15583), .ZN(
        n11344) );
  AND2_X1 U13280 ( .A1(n11345), .A2(n11344), .ZN(n11346) );
  AND2_X1 U13281 ( .A1(n11347), .A2(n11346), .ZN(n11382) );
  INV_X1 U13282 ( .A(n11348), .ZN(n11349) );
  INV_X1 U13283 ( .A(n12774), .ZN(n11385) );
  AOI21_X1 U13284 ( .B1(n12774), .B2(n11349), .A(n11538), .ZN(n11387) );
  AOI22_X1 U13285 ( .A1(n11387), .A2(n16153), .B1(n12774), .B2(n16151), .ZN(
        n11350) );
  OAI211_X1 U13286 ( .C1(n16116), .C2(n11390), .A(n11382), .B(n11350), .ZN(
        n11353) );
  NAND2_X1 U13287 ( .A1(n11353), .A2(n16183), .ZN(n11351) );
  OAI21_X1 U13288 ( .B1(n16183), .B2(n11352), .A(n11351), .ZN(P1_U3477) );
  NAND2_X1 U13289 ( .A1(n11353), .A2(n16179), .ZN(n11354) );
  OAI21_X1 U13290 ( .B1(n16179), .B2(n10306), .A(n11354), .ZN(P1_U3534) );
  XNOR2_X1 U13291 ( .A(n15234), .B(n12762), .ZN(n13011) );
  XNOR2_X1 U13292 ( .A(n13011), .B(n11355), .ZN(n16075) );
  OR2_X1 U13293 ( .A1(n16022), .A2(n16074), .ZN(n15622) );
  XOR2_X1 U13294 ( .A(n13011), .B(n11356), .Z(n16077) );
  NAND2_X1 U13295 ( .A1(n16077), .A2(n15620), .ZN(n11365) );
  AOI21_X1 U13296 ( .B1(n12762), .B2(n11358), .A(n11357), .ZN(n16072) );
  AOI22_X1 U13297 ( .A1(n15500), .A2(n15235), .B1(n15233), .B2(n15437), .ZN(
        n16069) );
  INV_X1 U13298 ( .A(n16069), .ZN(n11360) );
  AOI22_X1 U13299 ( .A1(n11360), .A2(n15611), .B1(n11359), .B2(n16011), .ZN(
        n11362) );
  NAND2_X1 U13300 ( .A1(n15617), .A2(n12762), .ZN(n11361) );
  OAI211_X1 U13301 ( .C1(n10277), .C2(n15611), .A(n11362), .B(n11361), .ZN(
        n11363) );
  AOI21_X1 U13302 ( .B1(n15601), .B2(n16072), .A(n11363), .ZN(n11364) );
  OAI211_X1 U13303 ( .C1(n16075), .C2(n15622), .A(n11365), .B(n11364), .ZN(
        P1_U3289) );
  NAND2_X1 U13304 ( .A1(n11367), .A2(n14804), .ZN(n11366) );
  OAI21_X1 U13305 ( .B1(n11367), .B2(n14804), .A(n11366), .ZN(n11369) );
  OAI211_X1 U13306 ( .C1(n11370), .C2(n11369), .A(n11368), .B(n15898), .ZN(
        n11379) );
  NAND2_X1 U13307 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n12572)
         );
  AOI211_X1 U13308 ( .C1(n11374), .C2(n11373), .A(n11372), .B(n11371), .ZN(
        n11375) );
  INV_X1 U13309 ( .A(n11375), .ZN(n11376) );
  NAND2_X1 U13310 ( .A1(n12572), .A2(n11376), .ZN(n11377) );
  AOI21_X1 U13311 ( .B1(n15858), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n11377), 
        .ZN(n11378) );
  OAI211_X1 U13312 ( .C1(n15837), .C2(n11380), .A(n11379), .B(n11378), .ZN(
        P2_U3227) );
  MUX2_X1 U13313 ( .A(n11382), .B(n11381), .S(n16022), .Z(n11389) );
  INV_X1 U13314 ( .A(n11383), .ZN(n11384) );
  OAI22_X1 U13315 ( .A1(n11385), .A2(n16014), .B1(n15615), .B2(n11384), .ZN(
        n11386) );
  AOI21_X1 U13316 ( .B1(n11387), .B2(n15601), .A(n11386), .ZN(n11388) );
  OAI211_X1 U13317 ( .C1(n11390), .C2(n15598), .A(n11389), .B(n11388), .ZN(
        P1_U3287) );
  XNOR2_X1 U13318 ( .A(n9026), .B(n7717), .ZN(n11401) );
  OAI21_X1 U13319 ( .B1(n9026), .B2(n11393), .A(n11392), .ZN(n11397) );
  OAI22_X1 U13320 ( .A1(n11395), .A2(n14794), .B1(n11394), .B2(n14600), .ZN(
        n11396) );
  AOI21_X1 U13321 ( .B1(n11397), .B2(n9112), .A(n11396), .ZN(n11398) );
  OAI21_X1 U13322 ( .B1(n11401), .B2(n14876), .A(n11398), .ZN(n12117) );
  AOI211_X1 U13323 ( .C1(n11399), .C2(n7718), .A(n14300), .B(n11412), .ZN(
        n12113) );
  NOR2_X1 U13324 ( .A1(n12117), .A2(n12113), .ZN(n12133) );
  MUX2_X1 U13325 ( .A(n11400), .B(n12133), .S(n16208), .Z(n11403) );
  INV_X1 U13326 ( .A(n11401), .ZN(n12135) );
  NAND2_X1 U13327 ( .A1(n11947), .A2(n12135), .ZN(n11402) );
  OAI211_X1 U13328 ( .C1(n8630), .C2(n14896), .A(n11403), .B(n11402), .ZN(
        P2_U3500) );
  XNOR2_X1 U13329 ( .A(n11405), .B(n11404), .ZN(n11725) );
  OAI21_X1 U13330 ( .B1(n11408), .B2(n11407), .A(n11406), .ZN(n11410) );
  AOI21_X1 U13331 ( .B1(n11410), .B2(n9112), .A(n11409), .ZN(n11728) );
  OAI211_X1 U13332 ( .C1(n11413), .C2(n11412), .A(n11411), .B(n14267), .ZN(
        n11719) );
  OAI211_X1 U13333 ( .C1(n11413), .C2(n16201), .A(n11728), .B(n11719), .ZN(
        n11414) );
  AOI21_X1 U13334 ( .B1(n14884), .B2(n11725), .A(n11414), .ZN(n11464) );
  AOI22_X1 U13335 ( .A1(n11947), .A2(n11725), .B1(n16206), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n11415) );
  OAI21_X1 U13336 ( .B1(n11464), .B2(n16206), .A(n11415), .ZN(P2_U3501) );
  XNOR2_X1 U13337 ( .A(n11416), .B(n11419), .ZN(n11846) );
  INV_X1 U13338 ( .A(n11417), .ZN(n11499) );
  OAI211_X1 U13339 ( .C1(n11418), .C2(n11593), .A(n11499), .B(n14267), .ZN(
        n11842) );
  OAI21_X1 U13340 ( .B1(n11418), .B2(n16201), .A(n11842), .ZN(n11423) );
  XNOR2_X1 U13341 ( .A(n11420), .B(n11419), .ZN(n11422) );
  OAI21_X1 U13342 ( .B1(n11422), .B2(n14719), .A(n11421), .ZN(n11843) );
  AOI211_X1 U13343 ( .C1(n14884), .C2(n11846), .A(n11423), .B(n11843), .ZN(
        n11492) );
  AOI22_X1 U13344 ( .A1(n11846), .A2(n11947), .B1(n16206), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n11424) );
  OAI21_X1 U13345 ( .B1(n11492), .B2(n16206), .A(n11424), .ZN(P2_U3504) );
  INV_X1 U13346 ( .A(n12651), .ZN(n11436) );
  INV_X1 U13347 ( .A(n15849), .ZN(n11868) );
  OAI222_X1 U13348 ( .A1(n14970), .A2(n11425), .B1(n14968), .B2(n11436), .C1(
        n11868), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13349 ( .A(n11426), .ZN(n11429) );
  INV_X1 U13350 ( .A(n11427), .ZN(n11428) );
  NAND2_X1 U13351 ( .A1(n11429), .A2(n11428), .ZN(n11431) );
  NAND2_X1 U13352 ( .A1(n11431), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11430) );
  MUX2_X1 U13353 ( .A(P1_IR_REG_31__SCAN_IN), .B(n11430), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n11434) );
  INV_X1 U13354 ( .A(n11431), .ZN(n11433) );
  NAND2_X1 U13355 ( .A1(n11433), .A2(n11432), .ZN(n11610) );
  NAND2_X1 U13356 ( .A1(n11434), .A2(n11610), .ZN(n12279) );
  OAI222_X1 U13357 ( .A1(n7190), .A2(n12279), .B1(n15771), .B2(n11436), .C1(
        n11435), .C2(n15773), .ZN(P1_U3339) );
  INV_X1 U13358 ( .A(n11437), .ZN(n11440) );
  INV_X1 U13359 ( .A(n11438), .ZN(n11439) );
  NAND2_X1 U13360 ( .A1(n11442), .A2(n12998), .ZN(n11445) );
  AOI22_X1 U13361 ( .A1(n12836), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12835), 
        .B2(n11443), .ZN(n11444) );
  NAND2_X1 U13362 ( .A1(n11445), .A2(n11444), .ZN(n16111) );
  INV_X1 U13363 ( .A(n16111), .ZN(n11542) );
  OAI22_X1 U13364 ( .A1(n11542), .A2(n15095), .B1(n11786), .B2(n15094), .ZN(
        n11773) );
  NAND2_X1 U13365 ( .A1(n16111), .A2(n15062), .ZN(n11447) );
  NAND2_X1 U13366 ( .A1(n15231), .A2(n11123), .ZN(n11446) );
  NAND2_X1 U13367 ( .A1(n11447), .A2(n11446), .ZN(n11448) );
  XNOR2_X1 U13368 ( .A(n11448), .B(n15065), .ZN(n11772) );
  XOR2_X1 U13369 ( .A(n11773), .B(n11772), .Z(n11774) );
  XNOR2_X1 U13370 ( .A(n11775), .B(n11774), .ZN(n11460) );
  NAND2_X1 U13371 ( .A1(n10755), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n11455) );
  NAND2_X1 U13372 ( .A1(n12966), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n11454) );
  INV_X1 U13373 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n11449) );
  NAND2_X1 U13374 ( .A1(n11450), .A2(n11449), .ZN(n11451) );
  AND2_X1 U13375 ( .A1(n11702), .A2(n11451), .ZN(n11715) );
  NAND2_X1 U13376 ( .A1(n12965), .A2(n11715), .ZN(n11453) );
  NAND2_X1 U13377 ( .A1(n12982), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11452) );
  NAND4_X1 U13378 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n15230) );
  AOI22_X1 U13379 ( .A1(n15500), .A2(n15232), .B1(n15230), .B2(n15437), .ZN(
        n11534) );
  NAND2_X1 U13380 ( .A1(n15216), .A2(n11540), .ZN(n11457) );
  OAI211_X1 U13381 ( .C1(n11534), .C2(n15213), .A(n11457), .B(n11456), .ZN(
        n11458) );
  AOI21_X1 U13382 ( .B1(n16111), .B2(n15196), .A(n11458), .ZN(n11459) );
  OAI21_X1 U13383 ( .B1(n11460), .B2(n15205), .A(n11459), .ZN(P1_U3213) );
  INV_X1 U13384 ( .A(n14953), .ZN(n14919) );
  INV_X1 U13385 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11461) );
  NOR2_X1 U13386 ( .A1(n14948), .A2(n11461), .ZN(n11462) );
  AOI21_X1 U13387 ( .B1(n14919), .B2(n11725), .A(n11462), .ZN(n11463) );
  OAI21_X1 U13388 ( .B1(n11464), .B2(n16209), .A(n11463), .ZN(P2_U3436) );
  OAI21_X1 U13389 ( .B1(n11466), .B2(n13119), .A(n11465), .ZN(n11750) );
  OAI211_X1 U13390 ( .C1(n11468), .C2(n13260), .A(n11467), .B(n14103), .ZN(
        n11470) );
  AOI22_X1 U13391 ( .A1(n14108), .A2(n13520), .B1(n13518), .B2(n14107), .ZN(
        n11469) );
  NAND2_X1 U13392 ( .A1(n11470), .A2(n11469), .ZN(n11747) );
  AOI21_X1 U13393 ( .B1(n16226), .B2(n11750), .A(n11747), .ZN(n11476) );
  OAI22_X1 U13394 ( .A1(n14192), .A2(n11746), .B1(n16228), .B2(n10667), .ZN(
        n11471) );
  INV_X1 U13395 ( .A(n11471), .ZN(n11472) );
  OAI21_X1 U13396 ( .B1(n11476), .B2(n7687), .A(n11472), .ZN(P3_U3465) );
  INV_X1 U13397 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n11473) );
  OAI22_X1 U13398 ( .A1(n14246), .A2(n11746), .B1(n16232), .B2(n11473), .ZN(
        n11474) );
  INV_X1 U13399 ( .A(n11474), .ZN(n11475) );
  OAI21_X1 U13400 ( .B1(n11476), .B2(n16229), .A(n11475), .ZN(P3_U3408) );
  OAI21_X1 U13401 ( .B1(n11478), .B2(n13113), .A(n11477), .ZN(n11766) );
  INV_X1 U13402 ( .A(n11479), .ZN(n11480) );
  AOI21_X1 U13403 ( .B1(n13113), .B2(n11481), .A(n11480), .ZN(n11482) );
  OAI222_X1 U13404 ( .A1(n16032), .A2(n11795), .B1(n16034), .B2(n7730), .C1(
        n16039), .C2(n11482), .ZN(n11761) );
  AOI21_X1 U13405 ( .B1(n16226), .B2(n11766), .A(n11761), .ZN(n11488) );
  INV_X1 U13406 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n11483) );
  OAI22_X1 U13407 ( .A1(n14246), .A2(n11763), .B1(n16232), .B2(n11483), .ZN(
        n11484) );
  INV_X1 U13408 ( .A(n11484), .ZN(n11485) );
  OAI21_X1 U13409 ( .B1(n11488), .B2(n16229), .A(n11485), .ZN(P3_U3405) );
  OAI22_X1 U13410 ( .A1(n14192), .A2(n11763), .B1(n16228), .B2(n10502), .ZN(
        n11486) );
  INV_X1 U13411 ( .A(n11486), .ZN(n11487) );
  OAI21_X1 U13412 ( .B1(n11488), .B2(n7687), .A(n11487), .ZN(P3_U3464) );
  INV_X1 U13413 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11489) );
  NOR2_X1 U13414 ( .A1(n14948), .A2(n11489), .ZN(n11490) );
  AOI21_X1 U13415 ( .B1(n11846), .B2(n14919), .A(n11490), .ZN(n11491) );
  OAI21_X1 U13416 ( .B1(n11492), .B2(n16209), .A(n11491), .ZN(P2_U3445) );
  XOR2_X1 U13417 ( .A(n11493), .B(n11494), .Z(n11556) );
  XNOR2_X1 U13418 ( .A(n11495), .B(n11494), .ZN(n11497) );
  NAND2_X1 U13419 ( .A1(n14480), .A2(n14647), .ZN(n11496) );
  OAI21_X1 U13420 ( .B1(n11679), .B2(n14600), .A(n11496), .ZN(n11507) );
  AOI21_X1 U13421 ( .B1(n11497), .B2(n9112), .A(n11507), .ZN(n11548) );
  INV_X1 U13422 ( .A(n11669), .ZN(n11498) );
  AOI211_X1 U13423 ( .C1(n11508), .C2(n11499), .A(n14300), .B(n11498), .ZN(
        n11553) );
  INV_X1 U13424 ( .A(n11553), .ZN(n11500) );
  OAI211_X1 U13425 ( .C1(n11556), .C2(n16138), .A(n11548), .B(n11500), .ZN(
        n12323) );
  OAI22_X1 U13426 ( .A1(n14896), .A2(n12321), .B1(n16208), .B2(n10913), .ZN(
        n11501) );
  AOI21_X1 U13427 ( .B1(n12323), .B2(n16208), .A(n11501), .ZN(n11502) );
  INV_X1 U13428 ( .A(n11502), .ZN(P2_U3505) );
  INV_X1 U13429 ( .A(n11503), .ZN(n11504) );
  XNOR2_X1 U13430 ( .A(n11508), .B(n14352), .ZN(n11674) );
  NAND2_X1 U13431 ( .A1(n14479), .A2(n14300), .ZN(n11673) );
  XNOR2_X1 U13432 ( .A(n11674), .B(n11673), .ZN(n11676) );
  XOR2_X1 U13433 ( .A(n11677), .B(n11676), .Z(n11512) );
  INV_X1 U13434 ( .A(n11506), .ZN(n11551) );
  AND2_X1 U13435 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n14538) );
  AOI21_X1 U13436 ( .B1(n14392), .B2(n11507), .A(n14538), .ZN(n11510) );
  NAND2_X1 U13437 ( .A1(n14423), .A2(n11508), .ZN(n11509) );
  OAI211_X1 U13438 ( .C1(n14403), .C2(n11551), .A(n11510), .B(n11509), .ZN(
        n11511) );
  AOI21_X1 U13439 ( .B1(n11512), .B2(n14420), .A(n11511), .ZN(n11513) );
  INV_X1 U13440 ( .A(n11513), .ZN(P2_U3211) );
  NAND4_X1 U13441 ( .A1(n15820), .A2(n15821), .A3(n11515), .A4(n11514), .ZN(
        n11516) );
  INV_X1 U13442 ( .A(n16094), .ZN(n14623) );
  INV_X1 U13443 ( .A(n11517), .ZN(n11521) );
  OAI22_X1 U13444 ( .A1(n11519), .A2(n14697), .B1(n11518), .B2(n7193), .ZN(
        n11520) );
  OAI21_X1 U13445 ( .B1(n11521), .B2(n11520), .A(n14805), .ZN(n11526) );
  NAND2_X1 U13446 ( .A1(n7193), .A2(n8503), .ZN(n11546) );
  INV_X1 U13447 ( .A(n14806), .ZN(n16089) );
  INV_X1 U13448 ( .A(n11523), .ZN(n11524) );
  NAND2_X1 U13449 ( .A1(n16089), .A2(n11524), .ZN(n11525) );
  OAI211_X1 U13450 ( .C1(n11213), .C2(n14623), .A(n11526), .B(n11525), .ZN(
        P2_U3265) );
  NAND2_X1 U13451 ( .A1(n11528), .A2(n11527), .ZN(n11530) );
  OR2_X1 U13452 ( .A1(n12774), .A2(n15232), .ZN(n11529) );
  NAND2_X1 U13453 ( .A1(n11530), .A2(n11529), .ZN(n11691) );
  XNOR2_X1 U13454 ( .A(n16111), .B(n15231), .ZN(n13017) );
  INV_X1 U13455 ( .A(n13017), .ZN(n11690) );
  XNOR2_X1 U13456 ( .A(n11691), .B(n11690), .ZN(n11537) );
  INV_X1 U13457 ( .A(n11537), .ZN(n16115) );
  OR2_X1 U13458 ( .A1(n12774), .A2(n11531), .ZN(n11532) );
  XNOR2_X1 U13459 ( .A(n11699), .B(n13017), .ZN(n11535) );
  OAI21_X1 U13460 ( .B1(n11535), .B2(n16074), .A(n11534), .ZN(n11536) );
  AOI21_X1 U13461 ( .B1(n15490), .B2(n11537), .A(n11536), .ZN(n16114) );
  MUX2_X1 U13462 ( .A(n10316), .B(n16114), .S(n15611), .Z(n11545) );
  INV_X1 U13463 ( .A(n11538), .ZN(n11539) );
  NAND2_X1 U13464 ( .A1(n11538), .A2(n11542), .ZN(n11714) );
  AOI21_X1 U13465 ( .B1(n16111), .B2(n11539), .A(n7486), .ZN(n16112) );
  INV_X1 U13466 ( .A(n11540), .ZN(n11541) );
  OAI22_X1 U13467 ( .A1(n11542), .A2(n16014), .B1(n11541), .B2(n15615), .ZN(
        n11543) );
  AOI21_X1 U13468 ( .B1(n16112), .B2(n15601), .A(n11543), .ZN(n11544) );
  OAI211_X1 U13469 ( .C1(n16115), .C2(n15598), .A(n11545), .B(n11544), .ZN(
        P1_U3286) );
  AND2_X1 U13470 ( .A1(n14876), .A2(n11546), .ZN(n11547) );
  MUX2_X1 U13471 ( .A(n11549), .B(n11548), .S(n14623), .Z(n11555) );
  OAI22_X1 U13472 ( .A1(n16085), .A2(n12321), .B1(n14697), .B2(n11551), .ZN(
        n11552) );
  AOI21_X1 U13473 ( .B1(n11553), .B2(n16088), .A(n11552), .ZN(n11554) );
  OAI211_X1 U13474 ( .C1(n11556), .C2(n16062), .A(n11555), .B(n11554), .ZN(
        P2_U3259) );
  NAND2_X1 U13475 ( .A1(n13739), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11557) );
  OAI21_X1 U13476 ( .B1(n13919), .B2(n13739), .A(n11557), .ZN(P3_U3520) );
  NOR2_X1 U13477 ( .A1(n11575), .A2(n11558), .ZN(n11560) );
  INV_X1 U13478 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11561) );
  OR2_X1 U13479 ( .A1(n11953), .A2(n11561), .ZN(n11949) );
  NAND2_X1 U13480 ( .A1(n11953), .A2(n11561), .ZN(n11562) );
  NAND2_X1 U13481 ( .A1(n11949), .A2(n11562), .ZN(n11564) );
  INV_X1 U13482 ( .A(n11950), .ZN(n11563) );
  AOI21_X1 U13483 ( .B1(n11565), .B2(n11564), .A(n11563), .ZN(n11573) );
  MUX2_X1 U13484 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13309), .Z(n11952) );
  XNOR2_X1 U13485 ( .A(n11952), .B(n11583), .ZN(n11571) );
  INV_X1 U13486 ( .A(n11956), .ZN(n11569) );
  AOI21_X1 U13487 ( .B1(n11571), .B2(n11570), .A(n11569), .ZN(n11572) );
  OAI22_X1 U13488 ( .A1(n11573), .A2(n13899), .B1(n11572), .B2(n13877), .ZN(
        n11586) );
  NOR2_X1 U13489 ( .A1(n11575), .A2(n11574), .ZN(n11577) );
  OR2_X1 U13490 ( .A1(n11953), .A2(n12257), .ZN(n11959) );
  NAND2_X1 U13491 ( .A1(n11953), .A2(n12257), .ZN(n11578) );
  NAND2_X1 U13492 ( .A1(n11959), .A2(n11578), .ZN(n11579) );
  NAND2_X1 U13493 ( .A1(n11580), .A2(n11579), .ZN(n11581) );
  AOI21_X1 U13494 ( .B1(n11960), .B2(n11581), .A(n13895), .ZN(n11585) );
  INV_X1 U13495 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n13621) );
  NOR2_X1 U13496 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13621), .ZN(n12244) );
  AOI21_X1 U13497 ( .B1(n15817), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12244), 
        .ZN(n11582) );
  OAI21_X1 U13498 ( .B1(n13889), .B2(n11583), .A(n11582), .ZN(n11584) );
  OR3_X1 U13499 ( .A1(n11586), .A2(n11585), .A3(n11584), .ZN(P3_U3192) );
  NAND2_X1 U13500 ( .A1(n13102), .A2(n16045), .ZN(n12154) );
  NAND2_X1 U13501 ( .A1(n14017), .A2(n12154), .ZN(n16123) );
  OAI22_X1 U13502 ( .A1(n16126), .A2(n13111), .B1(n11587), .B2(n16128), .ZN(
        n11590) );
  MUX2_X1 U13503 ( .A(n11588), .B(P3_REG2_REG_4__SCAN_IN), .S(n16052), .Z(
        n11589) );
  AOI211_X1 U13504 ( .C1(n14099), .C2(n11591), .A(n11590), .B(n11589), .ZN(
        n11592) );
  INV_X1 U13505 ( .A(n11592), .ZN(P3_U3229) );
  AOI211_X1 U13506 ( .C1(n11603), .C2(n11594), .A(n14300), .B(n11593), .ZN(
        n16087) );
  OAI21_X1 U13507 ( .B1(n11596), .B2(n11597), .A(n11595), .ZN(n11601) );
  XNOR2_X1 U13508 ( .A(n11598), .B(n11597), .ZN(n11607) );
  NOR2_X1 U13509 ( .A1(n11607), .A2(n14876), .ZN(n11599) );
  AOI211_X1 U13510 ( .C1(n9112), .C2(n11601), .A(n11600), .B(n11599), .ZN(
        n16093) );
  INV_X1 U13511 ( .A(n16093), .ZN(n11602) );
  AOI211_X1 U13512 ( .C1(n16134), .C2(n11603), .A(n16087), .B(n11602), .ZN(
        n11609) );
  INV_X1 U13513 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11604) );
  OAI22_X1 U13514 ( .A1(n11607), .A2(n14953), .B1(n14948), .B2(n11604), .ZN(
        n11605) );
  INV_X1 U13515 ( .A(n11605), .ZN(n11606) );
  OAI21_X1 U13516 ( .B1(n11609), .B2(n16209), .A(n11606), .ZN(P2_U3442) );
  INV_X1 U13517 ( .A(n11607), .ZN(n16090) );
  AOI22_X1 U13518 ( .A1(n16090), .A2(n11947), .B1(n16206), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n11608) );
  OAI21_X1 U13519 ( .B1(n11609), .B2(n16206), .A(n11608), .ZN(P2_U3503) );
  INV_X1 U13520 ( .A(n12822), .ZN(n11617) );
  NAND2_X1 U13521 ( .A1(n11610), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11611) );
  MUX2_X1 U13522 ( .A(P1_IR_REG_31__SCAN_IN), .B(n11611), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n11614) );
  INV_X1 U13523 ( .A(n11612), .ZN(n11613) );
  AND2_X1 U13524 ( .A1(n11614), .A2(n11613), .ZN(n12823) );
  INV_X1 U13525 ( .A(n12823), .ZN(n12285) );
  OAI222_X1 U13526 ( .A1(n15773), .A2(n11615), .B1(n15771), .B2(n11617), .C1(
        P1_U3086), .C2(n12285), .ZN(P1_U3338) );
  INV_X1 U13527 ( .A(n15864), .ZN(n11616) );
  OAI222_X1 U13528 ( .A1(n14970), .A2(n11618), .B1(n14968), .B2(n11617), .C1(
        P2_U3088), .C2(n11616), .ZN(P2_U3310) );
  OAI21_X1 U13529 ( .B1(n11620), .B2(n13124), .A(n11619), .ZN(n16105) );
  OAI211_X1 U13530 ( .C1(n11622), .C2(n13259), .A(n11621), .B(n14103), .ZN(
        n11624) );
  AOI22_X1 U13531 ( .A1(n14107), .A2(n13517), .B1(n13519), .B2(n14108), .ZN(
        n11623) );
  NAND2_X1 U13532 ( .A1(n11624), .A2(n11623), .ZN(n16104) );
  AOI21_X1 U13533 ( .B1(n16226), .B2(n16105), .A(n16104), .ZN(n11630) );
  INV_X1 U13534 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11625) );
  OAI22_X1 U13535 ( .A1(n14246), .A2(n16108), .B1(n16232), .B2(n11625), .ZN(
        n11626) );
  INV_X1 U13536 ( .A(n11626), .ZN(n11627) );
  OAI21_X1 U13537 ( .B1(n11630), .B2(n16229), .A(n11627), .ZN(P3_U3411) );
  OAI22_X1 U13538 ( .A1(n14192), .A2(n16108), .B1(n16228), .B2(n10658), .ZN(
        n11628) );
  INV_X1 U13539 ( .A(n11628), .ZN(n11629) );
  OAI21_X1 U13540 ( .B1(n11630), .B2(n7687), .A(n11629), .ZN(P3_U3466) );
  AOI21_X1 U13541 ( .B1(n11631), .B2(n13262), .A(n16039), .ZN(n11634) );
  OAI22_X1 U13542 ( .A1(n13100), .A2(n16034), .B1(n7730), .B2(n16032), .ZN(
        n11632) );
  AOI21_X1 U13543 ( .B1(n11634), .B2(n11633), .A(n11632), .ZN(n16056) );
  OAI21_X1 U13544 ( .B1(n11635), .B2(n13262), .A(n11636), .ZN(n16055) );
  INV_X1 U13545 ( .A(n16128), .ZN(n14079) );
  AOI22_X1 U13546 ( .A1(n14065), .A2(n16053), .B1(n14079), .B2(n13696), .ZN(
        n11637) );
  OAI21_X1 U13547 ( .B1(n10494), .B2(n16131), .A(n11637), .ZN(n11638) );
  AOI21_X1 U13548 ( .B1(n16055), .B2(n14099), .A(n11638), .ZN(n11639) );
  OAI21_X1 U13549 ( .B1(n16056), .B2(n16052), .A(n11639), .ZN(P3_U3230) );
  NOR2_X1 U13550 ( .A1(n11640), .A2(n16222), .ZN(n16024) );
  XNOR2_X1 U13551 ( .A(n11642), .B(n13258), .ZN(n11643) );
  NAND2_X1 U13552 ( .A1(n11643), .A2(n14103), .ZN(n11645) );
  AOI22_X1 U13553 ( .A1(n14108), .A2(n13740), .B1(n13523), .B2(n14107), .ZN(
        n11644) );
  NAND2_X1 U13554 ( .A1(n11645), .A2(n11644), .ZN(n16023) );
  AOI21_X1 U13555 ( .B1(n16024), .B2(n13294), .A(n16023), .ZN(n11646) );
  MUX2_X1 U13556 ( .A(n11647), .B(n11646), .S(n16131), .Z(n11650) );
  XNOR2_X1 U13557 ( .A(n11648), .B(n13258), .ZN(n16025) );
  AOI22_X1 U13558 ( .A1(n16025), .A2(n14099), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n14079), .ZN(n11649) );
  NAND2_X1 U13559 ( .A1(n11650), .A2(n11649), .ZN(P3_U3232) );
  XNOR2_X1 U13560 ( .A(n11746), .B(n13405), .ZN(n11793) );
  XNOR2_X1 U13561 ( .A(n11793), .B(n13519), .ZN(n11654) );
  AOI211_X1 U13562 ( .C1(n11654), .C2(n11653), .A(n13440), .B(n11792), .ZN(
        n11655) );
  INV_X1 U13563 ( .A(n11655), .ZN(n11659) );
  INV_X1 U13564 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n13614) );
  NOR2_X1 U13565 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13614), .ZN(n13771) );
  INV_X1 U13566 ( .A(n13518), .ZN(n12106) );
  OAI22_X1 U13567 ( .A1(n7795), .A2(n13500), .B1(n12106), .B2(n13470), .ZN(
        n11656) );
  AOI211_X1 U13568 ( .C1(n11657), .C2(n13411), .A(n13771), .B(n11656), .ZN(
        n11658) );
  OAI211_X1 U13569 ( .C1(n11745), .C2(n12627), .A(n11659), .B(n11658), .ZN(
        P3_U3179) );
  XNOR2_X1 U13570 ( .A(n11660), .B(n11661), .ZN(n11667) );
  OR2_X1 U13571 ( .A1(n11662), .A2(n11661), .ZN(n11663) );
  NAND2_X1 U13572 ( .A1(n11664), .A2(n11663), .ZN(n12297) );
  NAND2_X1 U13573 ( .A1(n12297), .A2(n14884), .ZN(n11666) );
  AOI22_X1 U13574 ( .A1(n14477), .A2(n14791), .B1(n14647), .B2(n14479), .ZN(
        n11665) );
  OAI211_X1 U13575 ( .C1(n11667), .C2(n14719), .A(n11666), .B(n11665), .ZN(
        n11831) );
  AOI21_X1 U13576 ( .B1(n11669), .B2(n11668), .A(n14300), .ZN(n11670) );
  AND2_X1 U13577 ( .A1(n11670), .A2(n11898), .ZN(n11835) );
  NOR2_X1 U13578 ( .A1(n11831), .A2(n11835), .ZN(n12299) );
  OAI22_X1 U13579 ( .A1(n14896), .A2(n12295), .B1(n16208), .B2(n10917), .ZN(
        n11671) );
  AOI21_X1 U13580 ( .B1(n12297), .B2(n11947), .A(n11671), .ZN(n11672) );
  OAI21_X1 U13581 ( .B1(n12299), .B2(n16206), .A(n11672), .ZN(P2_U3506) );
  INV_X1 U13582 ( .A(n11673), .ZN(n11675) );
  NOR2_X1 U13583 ( .A1(n11679), .A2(n14267), .ZN(n11681) );
  XNOR2_X1 U13584 ( .A(n12295), .B(n14304), .ZN(n11680) );
  NOR2_X1 U13585 ( .A1(n11680), .A2(n11681), .ZN(n11878) );
  AOI21_X1 U13586 ( .B1(n11681), .B2(n11680), .A(n11878), .ZN(n11682) );
  OAI21_X1 U13587 ( .B1(n7231), .B2(n11682), .A(n11880), .ZN(n11683) );
  NAND2_X1 U13588 ( .A1(n11683), .A2(n14420), .ZN(n11689) );
  INV_X1 U13589 ( .A(n11684), .ZN(n11687) );
  INV_X1 U13590 ( .A(n11685), .ZN(n11833) );
  OAI22_X1 U13591 ( .A1(n14404), .A2(n11875), .B1(n14403), .B2(n11833), .ZN(
        n11686) );
  AOI211_X1 U13592 ( .C1(n14443), .C2(n14479), .A(n11687), .B(n11686), .ZN(
        n11688) );
  OAI211_X1 U13593 ( .C1(n12295), .C2(n14462), .A(n11689), .B(n11688), .ZN(
        P2_U3185) );
  NAND2_X1 U13594 ( .A1(n11691), .A2(n11690), .ZN(n11693) );
  OR2_X1 U13595 ( .A1(n16111), .A2(n15231), .ZN(n11692) );
  NAND2_X1 U13596 ( .A1(n11693), .A2(n11692), .ZN(n11802) );
  NAND2_X1 U13597 ( .A1(n11694), .A2(n12998), .ZN(n11697) );
  AOI22_X1 U13598 ( .A1(n12836), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12835), 
        .B2(n11695), .ZN(n11696) );
  NAND2_X1 U13599 ( .A1(n11697), .A2(n11696), .ZN(n12780) );
  XNOR2_X1 U13600 ( .A(n12780), .B(n15230), .ZN(n13019) );
  INV_X1 U13601 ( .A(n13019), .ZN(n11801) );
  XNOR2_X1 U13602 ( .A(n11802), .B(n11801), .ZN(n11712) );
  INV_X1 U13603 ( .A(n11712), .ZN(n11755) );
  NAND2_X1 U13604 ( .A1(n16111), .A2(n11786), .ZN(n11698) );
  OR2_X1 U13605 ( .A1(n16111), .A2(n11786), .ZN(n11700) );
  XNOR2_X1 U13606 ( .A(n11809), .B(n13019), .ZN(n11710) );
  NAND2_X1 U13607 ( .A1(n12966), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11708) );
  NAND2_X1 U13608 ( .A1(n10755), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11707) );
  INV_X1 U13609 ( .A(n11811), .ZN(n11813) );
  NAND2_X1 U13610 ( .A1(n11702), .A2(n11701), .ZN(n11703) );
  AND2_X1 U13611 ( .A1(n11813), .A2(n11703), .ZN(n11825) );
  NAND2_X1 U13612 ( .A1(n12965), .A2(n11825), .ZN(n11706) );
  NAND2_X1 U13613 ( .A1(n12982), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11705) );
  NAND4_X1 U13614 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n15229) );
  AOI22_X1 U13615 ( .A1(n15582), .A2(n15231), .B1(n15229), .B2(n15437), .ZN(
        n11709) );
  OAI21_X1 U13616 ( .B1(n11710), .B2(n16074), .A(n11709), .ZN(n11711) );
  AOI21_X1 U13617 ( .B1(n15490), .B2(n11712), .A(n11711), .ZN(n11754) );
  MUX2_X1 U13618 ( .A(n10318), .B(n11754), .S(n15611), .Z(n11718) );
  INV_X1 U13619 ( .A(n11823), .ZN(n11713) );
  AOI21_X1 U13620 ( .B1(n12780), .B2(n11714), .A(n11713), .ZN(n11752) );
  INV_X1 U13621 ( .A(n11715), .ZN(n11787) );
  OAI22_X1 U13622 ( .A1(n7485), .A2(n16014), .B1(n15615), .B2(n11787), .ZN(
        n11716) );
  AOI21_X1 U13623 ( .B1(n11752), .B2(n15601), .A(n11716), .ZN(n11717) );
  OAI211_X1 U13624 ( .C1(n11755), .C2(n15598), .A(n11718), .B(n11717), .ZN(
        P1_U3285) );
  NOR2_X1 U13625 ( .A1(n14751), .A2(n11719), .ZN(n11723) );
  OAI22_X1 U13626 ( .A1(n14805), .A2(n11721), .B1(n11720), .B2(n14697), .ZN(
        n11722) );
  AOI211_X1 U13627 ( .C1(n14747), .C2(n11724), .A(n11723), .B(n11722), .ZN(
        n11727) );
  NAND2_X1 U13628 ( .A1(n11725), .A2(n14753), .ZN(n11726) );
  OAI211_X1 U13629 ( .C1(n16094), .C2(n11728), .A(n11727), .B(n11726), .ZN(
        P2_U3263) );
  INV_X1 U13630 ( .A(n11729), .ZN(n11730) );
  OAI222_X1 U13631 ( .A1(n11731), .A2(P3_U3151), .B1(n13319), .B2(n11730), 
        .C1(n13646), .C2(n14252), .ZN(P3_U3271) );
  AOI21_X1 U13632 ( .B1(n12521), .B2(P1_REG2_REG_14__SCAN_IN), .A(n11732), 
        .ZN(n12002) );
  XNOR2_X1 U13633 ( .A(n12002), .B(n12001), .ZN(n11733) );
  NOR2_X1 U13634 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11733), .ZN(n12006) );
  AOI21_X1 U13635 ( .B1(n11733), .B2(P1_REG2_REG_15__SCAN_IN), .A(n12006), 
        .ZN(n11744) );
  XNOR2_X1 U13636 ( .A(n12596), .B(n11996), .ZN(n11738) );
  INV_X1 U13637 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11737) );
  NAND2_X1 U13638 ( .A1(n11738), .A2(n11737), .ZN(n11997) );
  OAI21_X1 U13639 ( .B1(n11738), .B2(n11737), .A(n11997), .ZN(n11739) );
  NAND2_X1 U13640 ( .A1(n11739), .A2(n15927), .ZN(n11743) );
  INV_X1 U13641 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n11740) );
  NAND2_X1 U13642 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15212)
         );
  OAI21_X1 U13643 ( .B1(n15935), .B2(n11740), .A(n15212), .ZN(n11741) );
  AOI21_X1 U13644 ( .B1(n12596), .B2(n15929), .A(n11741), .ZN(n11742) );
  OAI211_X1 U13645 ( .C1(n11744), .C2(n15338), .A(n11743), .B(n11742), .ZN(
        P1_U3258) );
  OAI22_X1 U13646 ( .A1(n16126), .A2(n11746), .B1(n11745), .B2(n16128), .ZN(
        n11749) );
  MUX2_X1 U13647 ( .A(n11747), .B(P3_REG2_REG_6__SCAN_IN), .S(n16052), .Z(
        n11748) );
  AOI211_X1 U13648 ( .C1(n14099), .C2(n11750), .A(n11749), .B(n11748), .ZN(
        n11751) );
  INV_X1 U13649 ( .A(n11751), .ZN(P3_U3227) );
  INV_X1 U13650 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U13651 ( .A1(n11752), .A2(n16153), .B1(n12780), .B2(n16151), .ZN(
        n11753) );
  OAI211_X1 U13652 ( .C1(n16116), .C2(n11755), .A(n11754), .B(n11753), .ZN(
        n11758) );
  NAND2_X1 U13653 ( .A1(n11758), .A2(n16183), .ZN(n11756) );
  OAI21_X1 U13654 ( .B1(n16183), .B2(n11757), .A(n11756), .ZN(P1_U3483) );
  NAND2_X1 U13655 ( .A1(n11758), .A2(n16179), .ZN(n11759) );
  OAI21_X1 U13656 ( .B1(n16179), .B2(n11760), .A(n11759), .ZN(P1_U3536) );
  INV_X1 U13657 ( .A(n11761), .ZN(n11768) );
  NOR2_X1 U13658 ( .A1(n16131), .A2(n10503), .ZN(n11765) );
  OAI22_X1 U13659 ( .A1(n16126), .A2(n11763), .B1(n11762), .B2(n16128), .ZN(
        n11764) );
  AOI211_X1 U13660 ( .C1(n11766), .C2(n14099), .A(n11765), .B(n11764), .ZN(
        n11767) );
  OAI21_X1 U13661 ( .B1(n11768), .B2(n16052), .A(n11767), .ZN(P3_U3228) );
  INV_X1 U13662 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11771) );
  NAND2_X1 U13663 ( .A1(n11769), .A2(n14948), .ZN(n11770) );
  OAI21_X1 U13664 ( .B1(n14948), .B2(n11771), .A(n11770), .ZN(P2_U3439) );
  NAND2_X1 U13665 ( .A1(n12780), .A2(n15062), .ZN(n11777) );
  NAND2_X1 U13666 ( .A1(n15230), .A2(n11123), .ZN(n11776) );
  NAND2_X1 U13667 ( .A1(n11777), .A2(n11776), .ZN(n11778) );
  XNOR2_X1 U13668 ( .A(n11778), .B(n15065), .ZN(n11782) );
  NAND2_X1 U13669 ( .A1(n12780), .A2(n11123), .ZN(n11780) );
  NAND2_X1 U13670 ( .A1(n15230), .A2(n15050), .ZN(n11779) );
  NAND2_X1 U13671 ( .A1(n11780), .A2(n11779), .ZN(n11781) );
  NOR2_X1 U13672 ( .A1(n11782), .A2(n11781), .ZN(n11905) );
  AOI21_X1 U13673 ( .B1(n11782), .B2(n11781), .A(n11905), .ZN(n11783) );
  OAI21_X1 U13674 ( .B1(n11784), .B2(n11783), .A(n11907), .ZN(n11785) );
  NAND2_X1 U13675 ( .A1(n11785), .A2(n15210), .ZN(n11791) );
  OAI22_X1 U13676 ( .A1(n15192), .A2(n11787), .B1(n11786), .B2(n15191), .ZN(
        n11788) );
  AOI211_X1 U13677 ( .C1(n15182), .C2(n15229), .A(n11789), .B(n11788), .ZN(
        n11790) );
  OAI211_X1 U13678 ( .C1(n7485), .C2(n15220), .A(n11791), .B(n11790), .ZN(
        P1_U3221) );
  XNOR2_X1 U13679 ( .A(n16108), .B(n13405), .ZN(n11926) );
  XNOR2_X1 U13680 ( .A(n11926), .B(n13518), .ZN(n11927) );
  XOR2_X1 U13681 ( .A(n11928), .B(n11927), .Z(n11794) );
  NAND2_X1 U13682 ( .A1(n11794), .A2(n13495), .ZN(n11800) );
  INV_X1 U13683 ( .A(n13517), .ZN(n12127) );
  OAI22_X1 U13684 ( .A1(n12127), .A2(n13470), .B1(n11795), .B2(n13500), .ZN(
        n11796) );
  AOI211_X1 U13685 ( .C1(n11798), .C2(n13411), .A(n11797), .B(n11796), .ZN(
        n11799) );
  OAI211_X1 U13686 ( .C1(n16106), .C2(n12627), .A(n11800), .B(n11799), .ZN(
        P3_U3153) );
  NAND2_X1 U13687 ( .A1(n11802), .A2(n11801), .ZN(n11804) );
  OR2_X1 U13688 ( .A1(n12780), .A2(n15230), .ZN(n11803) );
  OR2_X1 U13689 ( .A1(n11805), .A2(n12987), .ZN(n11808) );
  AOI22_X1 U13690 ( .A1(n12836), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n12835), 
        .B2(n11806), .ZN(n11807) );
  INV_X1 U13691 ( .A(n15229), .ZN(n12070) );
  XNOR2_X1 U13692 ( .A(n16152), .B(n12070), .ZN(n13021) );
  XNOR2_X1 U13693 ( .A(n12085), .B(n13021), .ZN(n16150) );
  INV_X1 U13694 ( .A(n16150), .ZN(n11830) );
  INV_X1 U13695 ( .A(n15230), .ZN(n11916) );
  INV_X1 U13696 ( .A(n13021), .ZN(n11810) );
  XNOR2_X1 U13697 ( .A(n12069), .B(n11810), .ZN(n11821) );
  NAND2_X1 U13698 ( .A1(n16150), .A2(n15490), .ZN(n11820) );
  NAND2_X1 U13699 ( .A1(n12875), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11818) );
  NAND2_X1 U13700 ( .A1(n12966), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11817) );
  INV_X1 U13701 ( .A(n12028), .ZN(n12029) );
  INV_X1 U13702 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11812) );
  NAND2_X1 U13703 ( .A1(n11813), .A2(n11812), .ZN(n11814) );
  AND2_X1 U13704 ( .A1(n12029), .A2(n11814), .ZN(n12169) );
  NAND2_X1 U13705 ( .A1(n12965), .A2(n12169), .ZN(n11816) );
  NAND2_X1 U13706 ( .A1(n12982), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n11815) );
  NAND4_X1 U13707 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n15228) );
  AOI22_X1 U13708 ( .A1(n15500), .A2(n15230), .B1(n15228), .B2(n15583), .ZN(
        n11819) );
  OAI211_X1 U13709 ( .C1(n16074), .C2(n11821), .A(n11820), .B(n11819), .ZN(
        n16158) );
  MUX2_X1 U13710 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n16158), .S(n15611), .Z(
        n11822) );
  INV_X1 U13711 ( .A(n11822), .ZN(n11829) );
  AND2_X1 U13712 ( .A1(n16152), .A2(n11823), .ZN(n11824) );
  NOR2_X1 U13713 ( .A1(n12166), .A2(n11824), .ZN(n16154) );
  INV_X1 U13714 ( .A(n16152), .ZN(n11826) );
  INV_X1 U13715 ( .A(n11825), .ZN(n11917) );
  OAI22_X1 U13716 ( .A1(n11826), .A2(n16014), .B1(n11917), .B2(n15615), .ZN(
        n11827) );
  AOI21_X1 U13717 ( .B1(n16154), .B2(n15601), .A(n11827), .ZN(n11828) );
  OAI211_X1 U13718 ( .C1(n11830), .C2(n15598), .A(n11829), .B(n11828), .ZN(
        P1_U3284) );
  INV_X1 U13719 ( .A(n12297), .ZN(n11838) );
  MUX2_X1 U13720 ( .A(n11831), .B(P2_REG2_REG_7__SCAN_IN), .S(n16094), .Z(
        n11832) );
  INV_X1 U13721 ( .A(n11832), .ZN(n11837) );
  OAI22_X1 U13722 ( .A1(n16085), .A2(n12295), .B1(n14697), .B2(n11833), .ZN(
        n11834) );
  AOI21_X1 U13723 ( .B1(n11835), .B2(n16088), .A(n11834), .ZN(n11836) );
  OAI211_X1 U13724 ( .C1(n11838), .C2(n14806), .A(n11837), .B(n11836), .ZN(
        P2_U3258) );
  AOI22_X1 U13725 ( .A1(n14747), .A2(n11840), .B1(n16080), .B2(n11839), .ZN(
        n11841) );
  OAI21_X1 U13726 ( .B1(n14751), .B2(n11842), .A(n11841), .ZN(n11845) );
  MUX2_X1 U13727 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11843), .S(n14805), .Z(
        n11844) );
  AOI211_X1 U13728 ( .C1(n11846), .C2(n14753), .A(n11845), .B(n11844), .ZN(
        n11847) );
  INV_X1 U13729 ( .A(n11847), .ZN(P2_U3260) );
  INV_X1 U13730 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11853) );
  NOR2_X1 U13731 ( .A1(n11868), .A2(n11853), .ZN(n11848) );
  AOI21_X1 U13732 ( .B1(n11853), .B2(n11868), .A(n11848), .ZN(n15847) );
  NOR2_X1 U13733 ( .A1(n11850), .A2(n11849), .ZN(n11851) );
  NAND2_X1 U13734 ( .A1(n11864), .A2(n11851), .ZN(n11852) );
  XNOR2_X1 U13735 ( .A(n15836), .B(n11851), .ZN(n15840) );
  NAND2_X1 U13736 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15840), .ZN(n15839) );
  NAND2_X1 U13737 ( .A1(n11852), .A2(n15839), .ZN(n15848) );
  NAND2_X1 U13738 ( .A1(n15847), .A2(n15848), .ZN(n15846) );
  OAI21_X1 U13739 ( .B1(n11868), .B2(n11853), .A(n15846), .ZN(n11854) );
  INV_X1 U13740 ( .A(n11854), .ZN(n15862) );
  INV_X1 U13741 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11855) );
  MUX2_X1 U13742 ( .A(n11855), .B(P2_REG2_REG_17__SCAN_IN), .S(n15864), .Z(
        n15861) );
  NOR2_X1 U13743 ( .A1(n15862), .A2(n15861), .ZN(n15860) );
  AOI21_X1 U13744 ( .B1(n15864), .B2(P2_REG2_REG_17__SCAN_IN), .A(n15860), 
        .ZN(n11856) );
  INV_X1 U13745 ( .A(n11870), .ZN(n12059) );
  NAND2_X1 U13746 ( .A1(n11856), .A2(n12059), .ZN(n12055) );
  OAI21_X1 U13747 ( .B1(n11856), .B2(n12059), .A(n12055), .ZN(n11857) );
  NOR2_X1 U13748 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11857), .ZN(n12053) );
  AOI21_X1 U13749 ( .B1(n11857), .B2(P2_REG2_REG_18__SCAN_IN), .A(n12053), 
        .ZN(n11874) );
  NAND2_X1 U13750 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n11858)
         );
  OAI21_X1 U13751 ( .B1(n15837), .B2(n12059), .A(n11858), .ZN(n11859) );
  AOI21_X1 U13752 ( .B1(n15858), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n11859), 
        .ZN(n11873) );
  INV_X1 U13753 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11867) );
  XNOR2_X1 U13754 ( .A(n11868), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15851) );
  INV_X1 U13755 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11860) );
  OAI22_X1 U13756 ( .A1(n11863), .A2(n11862), .B1(n11861), .B2(n11860), .ZN(
        n11865) );
  NAND2_X1 U13757 ( .A1(n11864), .A2(n11865), .ZN(n11866) );
  XNOR2_X1 U13758 ( .A(n11865), .B(n15836), .ZN(n15842) );
  NAND2_X1 U13759 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15842), .ZN(n15841) );
  NAND2_X1 U13760 ( .A1(n11866), .A2(n15841), .ZN(n15852) );
  NAND2_X1 U13761 ( .A1(n15851), .A2(n15852), .ZN(n15850) );
  OAI21_X1 U13762 ( .B1(n11868), .B2(n11867), .A(n15850), .ZN(n15865) );
  INV_X1 U13763 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11869) );
  XNOR2_X1 U13764 ( .A(n15864), .B(n11869), .ZN(n15866) );
  AOI22_X1 U13765 ( .A1(n15865), .A2(n15866), .B1(n15864), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n12060) );
  XNOR2_X1 U13766 ( .A(n12060), .B(n11870), .ZN(n11871) );
  NAND2_X1 U13767 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11871), .ZN(n12058) );
  OAI211_X1 U13768 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n11871), .A(n15888), 
        .B(n12058), .ZN(n11872) );
  OAI211_X1 U13769 ( .C1(n11874), .C2(n15859), .A(n11873), .B(n11872), .ZN(
        P2_U3232) );
  NOR2_X1 U13770 ( .A1(n11875), .A2(n14267), .ZN(n11877) );
  XNOR2_X1 U13771 ( .A(n11901), .B(n14304), .ZN(n11876) );
  NOR2_X1 U13772 ( .A1(n11876), .A2(n11877), .ZN(n12041) );
  AOI21_X1 U13773 ( .B1(n11877), .B2(n11876), .A(n12041), .ZN(n11882) );
  INV_X1 U13774 ( .A(n11878), .ZN(n11879) );
  NAND2_X1 U13775 ( .A1(n11881), .A2(n11882), .ZN(n12043) );
  OAI21_X1 U13776 ( .B1(n11882), .B2(n11881), .A(n12043), .ZN(n11883) );
  NAND2_X1 U13777 ( .A1(n11883), .A2(n14420), .ZN(n11888) );
  INV_X1 U13778 ( .A(n11884), .ZN(n11900) );
  OAI22_X1 U13779 ( .A1(n14404), .A2(n12038), .B1(n14403), .B2(n11900), .ZN(
        n11885) );
  AOI211_X1 U13780 ( .C1(n14443), .C2(n14478), .A(n11886), .B(n11885), .ZN(
        n11887) );
  OAI211_X1 U13781 ( .C1(n11901), .C2(n14462), .A(n11888), .B(n11887), .ZN(
        P2_U3193) );
  INV_X1 U13782 ( .A(n11889), .ZN(n11890) );
  OAI222_X1 U13783 ( .A1(n11891), .A2(P3_U3151), .B1(n13319), .B2(n11890), 
        .C1(n13643), .C2(n14252), .ZN(P3_U3270) );
  NAND2_X1 U13784 ( .A1(n11892), .A2(n11895), .ZN(n11893) );
  NAND2_X1 U13785 ( .A1(n11894), .A2(n11893), .ZN(n16137) );
  OAI21_X1 U13786 ( .B1(n7356), .B2(n11895), .A(n11938), .ZN(n11896) );
  AOI222_X1 U13787 ( .A1(n9112), .A2(n11896), .B1(n14476), .B2(n14791), .C1(
        n14478), .C2(n14647), .ZN(n16136) );
  MUX2_X1 U13788 ( .A(n11897), .B(n16136), .S(n14805), .Z(n11904) );
  AOI21_X1 U13789 ( .B1(n11898), .B2(n16133), .A(n14300), .ZN(n11899) );
  AND2_X1 U13790 ( .A1(n11943), .A2(n11899), .ZN(n16132) );
  OAI22_X1 U13791 ( .A1(n16085), .A2(n11901), .B1(n14697), .B2(n11900), .ZN(
        n11902) );
  AOI21_X1 U13792 ( .B1(n16132), .B2(n16088), .A(n11902), .ZN(n11903) );
  OAI211_X1 U13793 ( .C1(n16062), .C2(n16137), .A(n11904), .B(n11903), .ZN(
        P2_U3257) );
  INV_X1 U13794 ( .A(n11905), .ZN(n11906) );
  NAND2_X1 U13795 ( .A1(n16152), .A2(n15062), .ZN(n11909) );
  NAND2_X1 U13796 ( .A1(n15229), .A2(n11123), .ZN(n11908) );
  NAND2_X1 U13797 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  XNOR2_X1 U13798 ( .A(n11910), .B(n15065), .ZN(n11914) );
  NAND2_X1 U13799 ( .A1(n16152), .A2(n11123), .ZN(n11912) );
  NAND2_X1 U13800 ( .A1(n15229), .A2(n15050), .ZN(n11911) );
  NAND2_X1 U13801 ( .A1(n11912), .A2(n11911), .ZN(n11913) );
  NAND2_X1 U13802 ( .A1(n11914), .A2(n11913), .ZN(n12019) );
  NAND2_X1 U13803 ( .A1(n7349), .A2(n12019), .ZN(n11915) );
  XNOR2_X1 U13804 ( .A(n12020), .B(n11915), .ZN(n11922) );
  OAI22_X1 U13805 ( .A1(n15192), .A2(n11917), .B1(n11916), .B2(n15191), .ZN(
        n11918) );
  AOI211_X1 U13806 ( .C1(n15182), .C2(n15228), .A(n11919), .B(n11918), .ZN(
        n11921) );
  NAND2_X1 U13807 ( .A1(n16152), .A2(n15196), .ZN(n11920) );
  OAI211_X1 U13808 ( .C1(n11922), .C2(n15205), .A(n11921), .B(n11920), .ZN(
        P1_U3231) );
  OAI222_X1 U13809 ( .A1(P2_U3088), .A2(n12059), .B1(n14968), .B2(n12834), 
        .C1(n11923), .C2(n14970), .ZN(P2_U3309) );
  NAND2_X1 U13810 ( .A1(n11613), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11924) );
  XNOR2_X1 U13811 ( .A(n11924), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15331) );
  INV_X1 U13812 ( .A(n15331), .ZN(n12699) );
  OAI222_X1 U13813 ( .A1(n15773), .A2(n11925), .B1(n15771), .B2(n12834), .C1(
        n12699), .C2(P1_U3086), .ZN(P1_U3337) );
  XNOR2_X1 U13814 ( .A(n13130), .B(n13405), .ZN(n12120) );
  XNOR2_X1 U13815 ( .A(n12120), .B(n13517), .ZN(n12122) );
  XOR2_X1 U13816 ( .A(n12123), .B(n12122), .Z(n11929) );
  NAND2_X1 U13817 ( .A1(n11929), .A2(n13495), .ZN(n11933) );
  OAI22_X1 U13818 ( .A1(n12106), .A2(n13500), .B1(n12238), .B2(n13470), .ZN(
        n11930) );
  AOI211_X1 U13819 ( .C1(n13130), .C2(n13411), .A(n11931), .B(n11930), .ZN(
        n11932) );
  OAI211_X1 U13820 ( .C1(n16127), .C2(n12627), .A(n11933), .B(n11932), .ZN(
        P3_U3161) );
  XNOR2_X1 U13821 ( .A(n11934), .B(n11937), .ZN(n12099) );
  AOI22_X1 U13822 ( .A1(n14647), .A2(n14477), .B1(n14475), .B2(n14791), .ZN(
        n11942) );
  INV_X1 U13823 ( .A(n11935), .ZN(n11940) );
  AND3_X1 U13824 ( .A1(n11938), .A2(n11937), .A3(n11936), .ZN(n11939) );
  OAI21_X1 U13825 ( .B1(n11940), .B2(n11939), .A(n9112), .ZN(n11941) );
  OAI211_X1 U13826 ( .C1(n12099), .C2(n14876), .A(n11942), .B(n11941), .ZN(
        n12092) );
  AOI211_X1 U13827 ( .C1(n11944), .C2(n11943), .A(n14300), .B(n12146), .ZN(
        n12096) );
  NOR2_X1 U13828 ( .A1(n12092), .A2(n12096), .ZN(n12293) );
  INV_X1 U13829 ( .A(n12099), .ZN(n12291) );
  OAI22_X1 U13830 ( .A1(n14896), .A2(n12289), .B1(n16208), .B2(n11945), .ZN(
        n11946) );
  AOI21_X1 U13831 ( .B1(n12291), .B2(n11947), .A(n11946), .ZN(n11948) );
  OAI21_X1 U13832 ( .B1(n12293), .B2(n16206), .A(n11948), .ZN(P2_U3508) );
  AOI21_X1 U13833 ( .B1(n9533), .B2(n11951), .A(n11986), .ZN(n11969) );
  INV_X1 U13834 ( .A(n11952), .ZN(n11954) );
  NAND2_X1 U13835 ( .A1(n11954), .A2(n11953), .ZN(n11955) );
  NAND2_X1 U13836 ( .A1(n11956), .A2(n11955), .ZN(n11958) );
  MUX2_X1 U13837 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13309), .Z(n11977) );
  XNOR2_X1 U13838 ( .A(n11977), .B(n8171), .ZN(n11957) );
  NAND2_X1 U13839 ( .A1(n11958), .A2(n11957), .ZN(n11980) );
  OAI21_X1 U13840 ( .B1(n11958), .B2(n11957), .A(n11980), .ZN(n11967) );
  INV_X1 U13841 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n13722) );
  NOR2_X1 U13842 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13722), .ZN(n12361) );
  AOI21_X1 U13843 ( .B1(n9534), .B2(n11961), .A(n11974), .ZN(n11962) );
  NOR2_X1 U13844 ( .A1(n13895), .A2(n11962), .ZN(n11963) );
  AOI211_X1 U13845 ( .C1(n15817), .C2(P3_ADDR_REG_11__SCAN_IN), .A(n12361), 
        .B(n11963), .ZN(n11964) );
  OAI21_X1 U13846 ( .B1(n11965), .B2(n13889), .A(n11964), .ZN(n11966) );
  AOI21_X1 U13847 ( .B1(n11967), .B2(n13897), .A(n11966), .ZN(n11968) );
  OAI21_X1 U13848 ( .B1(n11969), .B2(n13899), .A(n11968), .ZN(P3_U3193) );
  INV_X1 U13849 ( .A(n11970), .ZN(n11971) );
  OAI222_X1 U13850 ( .A1(n11972), .A2(P3_U3151), .B1(n13319), .B2(n11971), 
        .C1(n13640), .C2(n10650), .ZN(P3_U3269) );
  NOR2_X1 U13851 ( .A1(n8171), .A2(n11973), .ZN(n11975) );
  NAND2_X1 U13852 ( .A1(n12306), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12308) );
  OAI21_X1 U13853 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12306), .A(n12308), 
        .ZN(n11981) );
  NOR2_X1 U13854 ( .A1(n11976), .A2(n11981), .ZN(n12300) );
  AOI21_X1 U13855 ( .B1(n11976), .B2(n11981), .A(n12300), .ZN(n11995) );
  INV_X1 U13856 ( .A(n11977), .ZN(n11978) );
  NAND2_X1 U13857 ( .A1(n11978), .A2(n8171), .ZN(n11979) );
  NAND2_X1 U13858 ( .A1(n11980), .A2(n11979), .ZN(n11983) );
  XNOR2_X1 U13859 ( .A(n12306), .B(P3_REG1_REG_12__SCAN_IN), .ZN(n11988) );
  MUX2_X1 U13860 ( .A(n11981), .B(n11988), .S(n13309), .Z(n11982) );
  AOI21_X1 U13861 ( .B1(n11983), .B2(n11982), .A(n13877), .ZN(n11993) );
  NAND2_X1 U13862 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n12556)
         );
  NAND2_X1 U13863 ( .A1(n15817), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n11984) );
  OAI211_X1 U13864 ( .C1(n13889), .C2(n12306), .A(n12556), .B(n11984), .ZN(
        n11992) );
  NOR2_X1 U13865 ( .A1(n8171), .A2(n11985), .ZN(n11987) );
  AOI21_X1 U13866 ( .B1(n11989), .B2(n11988), .A(n12302), .ZN(n11990) );
  NOR2_X1 U13867 ( .A1(n11990), .A2(n13899), .ZN(n11991) );
  AOI211_X1 U13868 ( .C1(n11993), .C2(n12310), .A(n11992), .B(n11991), .ZN(
        n11994) );
  OAI21_X1 U13869 ( .B1(n11995), .B2(n13895), .A(n11994), .ZN(P3_U3194) );
  NAND2_X1 U13870 ( .A1(n11996), .A2(n12001), .ZN(n11998) );
  NAND2_X1 U13871 ( .A1(n11998), .A2(n11997), .ZN(n12000) );
  XNOR2_X1 U13872 ( .A(n12652), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11999) );
  NOR2_X1 U13873 ( .A1(n12000), .A2(n11999), .ZN(n12274) );
  AOI211_X1 U13874 ( .C1(n12000), .C2(n11999), .A(n12275), .B(n12274), .ZN(
        n12015) );
  INV_X1 U13875 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12007) );
  NAND2_X1 U13876 ( .A1(n12002), .A2(n12001), .ZN(n12009) );
  INV_X1 U13877 ( .A(n12006), .ZN(n12003) );
  NAND2_X1 U13878 ( .A1(n12009), .A2(n12003), .ZN(n12005) );
  NAND2_X1 U13879 ( .A1(n12652), .A2(n12007), .ZN(n12004) );
  OAI211_X1 U13880 ( .C1(n12652), .C2(n12007), .A(n12005), .B(n12004), .ZN(
        n12010) );
  AOI21_X1 U13881 ( .B1(n12279), .B2(n12007), .A(n12006), .ZN(n12008) );
  OAI211_X1 U13882 ( .C1(n12007), .C2(n12279), .A(n12009), .B(n12008), .ZN(
        n12278) );
  NAND3_X1 U13883 ( .A1(n12010), .A2(n15931), .A3(n12278), .ZN(n12013) );
  INV_X1 U13884 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n15134) );
  NOR2_X1 U13885 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15134), .ZN(n12011) );
  AOI21_X1 U13886 ( .B1(n15914), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n12011), 
        .ZN(n12012) );
  OAI211_X1 U13887 ( .C1(n15337), .C2(n12279), .A(n12013), .B(n12012), .ZN(
        n12014) );
  OR2_X1 U13888 ( .A1(n12015), .A2(n12014), .ZN(P1_U3259) );
  NAND2_X1 U13889 ( .A1(n12016), .A2(n12998), .ZN(n12018) );
  AOI22_X1 U13890 ( .A1(n12836), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n12835), 
        .B2(n15320), .ZN(n12017) );
  NAND2_X1 U13891 ( .A1(n12793), .A2(n15062), .ZN(n12022) );
  NAND2_X1 U13892 ( .A1(n15228), .A2(n11123), .ZN(n12021) );
  NAND2_X1 U13893 ( .A1(n12022), .A2(n12021), .ZN(n12023) );
  XNOR2_X1 U13894 ( .A(n12023), .B(n15065), .ZN(n12370) );
  AND2_X1 U13895 ( .A1(n15228), .A2(n15050), .ZN(n12024) );
  AOI21_X1 U13896 ( .B1(n12793), .B2(n11123), .A(n12024), .ZN(n12372) );
  XNOR2_X1 U13897 ( .A(n12370), .B(n12372), .ZN(n12025) );
  OAI211_X1 U13898 ( .C1(n12026), .C2(n12025), .A(n12371), .B(n15210), .ZN(
        n12037) );
  NAND2_X1 U13899 ( .A1(n12966), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n12034) );
  NAND2_X1 U13900 ( .A1(n12875), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U13901 ( .A1(n12029), .A2(n12375), .ZN(n12030) );
  AND2_X1 U13902 ( .A1(n12198), .A2(n12030), .ZN(n12377) );
  NAND2_X1 U13903 ( .A1(n12965), .A2(n12377), .ZN(n12032) );
  NAND2_X1 U13904 ( .A1(n12982), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n12031) );
  NAND4_X1 U13905 ( .A1(n12034), .A2(n12033), .A3(n12032), .A4(n12031), .ZN(
        n15227) );
  INV_X1 U13906 ( .A(n15227), .ZN(n12184) );
  NOR2_X1 U13907 ( .A1(n12184), .A2(n15482), .ZN(n12164) );
  AND2_X1 U13908 ( .A1(n15229), .A2(n15582), .ZN(n12175) );
  NOR2_X1 U13909 ( .A1(n12164), .A2(n12175), .ZN(n16169) );
  NAND2_X1 U13910 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(n7190), .ZN(n15315) );
  OAI21_X1 U13911 ( .B1(n16169), .B2(n15213), .A(n15315), .ZN(n12035) );
  AOI21_X1 U13912 ( .B1(n12169), .B2(n15216), .A(n12035), .ZN(n12036) );
  OAI211_X1 U13913 ( .C1(n16172), .C2(n15220), .A(n12037), .B(n12036), .ZN(
        P1_U3217) );
  NOR2_X1 U13914 ( .A1(n12038), .A2(n14267), .ZN(n12040) );
  XNOR2_X1 U13915 ( .A(n12289), .B(n14304), .ZN(n12039) );
  NOR2_X1 U13916 ( .A1(n12039), .A2(n12040), .ZN(n12226) );
  AOI21_X1 U13917 ( .B1(n12040), .B2(n12039), .A(n12226), .ZN(n12045) );
  INV_X1 U13918 ( .A(n12041), .ZN(n12042) );
  OAI21_X1 U13919 ( .B1(n12045), .B2(n12044), .A(n12228), .ZN(n12046) );
  NAND2_X1 U13920 ( .A1(n12046), .A2(n14420), .ZN(n12051) );
  NAND2_X1 U13921 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n15902) );
  INV_X1 U13922 ( .A(n15902), .ZN(n12049) );
  INV_X1 U13923 ( .A(n12093), .ZN(n12047) );
  OAI22_X1 U13924 ( .A1(n14404), .A2(n12335), .B1(n14403), .B2(n12047), .ZN(
        n12048) );
  AOI211_X1 U13925 ( .C1(n14443), .C2(n14477), .A(n12049), .B(n12048), .ZN(
        n12050) );
  OAI211_X1 U13926 ( .C1(n12289), .C2(n14462), .A(n12051), .B(n12050), .ZN(
        P2_U3203) );
  INV_X1 U13927 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n12052) );
  MUX2_X1 U13928 ( .A(n12052), .B(P2_REG2_REG_19__SCAN_IN), .S(n10115), .Z(
        n12057) );
  INV_X1 U13929 ( .A(n12053), .ZN(n12054) );
  NAND2_X1 U13930 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  XOR2_X1 U13931 ( .A(n12057), .B(n12056), .Z(n12067) );
  OAI21_X1 U13932 ( .B1(n12060), .B2(n12059), .A(n12058), .ZN(n12062) );
  INV_X1 U13933 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14857) );
  XNOR2_X1 U13934 ( .A(n10115), .B(n14857), .ZN(n12061) );
  XNOR2_X1 U13935 ( .A(n12062), .B(n12061), .ZN(n12065) );
  AND2_X1 U13936 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14345) );
  AOI21_X1 U13937 ( .B1(n15858), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n14345), 
        .ZN(n12063) );
  OAI21_X1 U13938 ( .B1(n10115), .B2(n15837), .A(n12063), .ZN(n12064) );
  AOI21_X1 U13939 ( .B1(n15888), .B2(n12065), .A(n12064), .ZN(n12066) );
  OAI21_X1 U13940 ( .B1(n12067), .B2(n15859), .A(n12066), .ZN(P2_U3233) );
  NOR2_X1 U13941 ( .A1(n16152), .A2(n12070), .ZN(n12068) );
  NAND2_X1 U13942 ( .A1(n16152), .A2(n12070), .ZN(n12071) );
  XNOR2_X1 U13943 ( .A(n12793), .B(n15228), .ZN(n13023) );
  INV_X1 U13944 ( .A(n13023), .ZN(n12171) );
  INV_X1 U13945 ( .A(n15228), .ZN(n12378) );
  OR2_X1 U13946 ( .A1(n12793), .A2(n12378), .ZN(n12073) );
  NAND2_X1 U13947 ( .A1(n12074), .A2(n12998), .ZN(n12077) );
  AOI22_X1 U13948 ( .A1(n12836), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n12835), 
        .B2(n12075), .ZN(n12076) );
  XNOR2_X1 U13949 ( .A(n12797), .B(n15227), .ZN(n13022) );
  XOR2_X1 U13950 ( .A(n12183), .B(n13022), .Z(n12082) );
  NAND2_X1 U13951 ( .A1(n12966), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U13952 ( .A1(n12982), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n12080) );
  XNOR2_X1 U13953 ( .A(n12198), .B(P1_REG3_REG_12__SCAN_IN), .ZN(n12512) );
  NAND2_X1 U13954 ( .A1(n12965), .A2(n12512), .ZN(n12079) );
  NAND2_X1 U13955 ( .A1(n10755), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n12078) );
  NAND4_X1 U13956 ( .A1(n12081), .A2(n12080), .A3(n12079), .A4(n12078), .ZN(
        n15226) );
  AOI222_X1 U13957 ( .A1(n15723), .A2(n12082), .B1(n15226), .B2(n15583), .C1(
        n15228), .C2(n15500), .ZN(n12386) );
  AOI21_X1 U13958 ( .B1(n12797), .B2(n12165), .A(n8016), .ZN(n12384) );
  INV_X1 U13959 ( .A(n12797), .ZN(n12084) );
  AOI22_X1 U13960 ( .A1(n16022), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12377), 
        .B2(n16011), .ZN(n12083) );
  OAI21_X1 U13961 ( .B1(n12084), .B2(n16014), .A(n12083), .ZN(n12090) );
  NAND2_X1 U13962 ( .A1(n12085), .A2(n13021), .ZN(n12087) );
  OR2_X1 U13963 ( .A1(n16152), .A2(n15229), .ZN(n12086) );
  NAND2_X1 U13964 ( .A1(n12087), .A2(n12086), .ZN(n12163) );
  OR2_X1 U13965 ( .A1(n12793), .A2(n15228), .ZN(n12088) );
  XNOR2_X1 U13966 ( .A(n12205), .B(n13022), .ZN(n12387) );
  NOR2_X1 U13967 ( .A1(n12387), .A2(n15577), .ZN(n12089) );
  AOI211_X1 U13968 ( .C1(n12384), .C2(n15601), .A(n12090), .B(n12089), .ZN(
        n12091) );
  OAI21_X1 U13969 ( .B1(n12386), .B2(n16022), .A(n12091), .ZN(P1_U3282) );
  NAND2_X1 U13970 ( .A1(n12092), .A2(n14623), .ZN(n12098) );
  AOI22_X1 U13971 ( .A1(n16082), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n12093), 
        .B2(n16080), .ZN(n12094) );
  OAI21_X1 U13972 ( .B1(n12289), .B2(n16085), .A(n12094), .ZN(n12095) );
  AOI21_X1 U13973 ( .B1(n12096), .B2(n16088), .A(n12095), .ZN(n12097) );
  OAI211_X1 U13974 ( .C1(n12099), .C2(n14806), .A(n12098), .B(n12097), .ZN(
        P2_U3256) );
  OAI21_X1 U13975 ( .B1(n12101), .B2(n13257), .A(n12100), .ZN(n16122) );
  INV_X1 U13976 ( .A(n12102), .ZN(n12103) );
  AOI21_X1 U13977 ( .B1(n13257), .B2(n12104), .A(n12103), .ZN(n12105) );
  OAI222_X1 U13978 ( .A1(n16032), .A2(n12238), .B1(n16034), .B2(n12106), .C1(
        n16039), .C2(n12105), .ZN(n16121) );
  AOI21_X1 U13979 ( .B1(n16226), .B2(n16122), .A(n16121), .ZN(n12112) );
  INV_X1 U13980 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n12107) );
  OAI22_X1 U13981 ( .A1(n14246), .A2(n16125), .B1(n16232), .B2(n12107), .ZN(
        n12108) );
  INV_X1 U13982 ( .A(n12108), .ZN(n12109) );
  OAI21_X1 U13983 ( .B1(n12112), .B2(n16229), .A(n12109), .ZN(P3_U3414) );
  OAI22_X1 U13984 ( .A1(n14192), .A2(n16125), .B1(n16228), .B2(n10798), .ZN(
        n12110) );
  INV_X1 U13985 ( .A(n12110), .ZN(n12111) );
  OAI21_X1 U13986 ( .B1(n12112), .B2(n7687), .A(n12111), .ZN(P3_U3467) );
  AOI22_X1 U13987 ( .A1(n16088), .A2(n12113), .B1(n16089), .B2(n12135), .ZN(
        n12115) );
  AOI22_X1 U13988 ( .A1(n16082), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n16080), .ZN(n12114) );
  OAI211_X1 U13989 ( .C1(n8630), .C2(n16085), .A(n12115), .B(n12114), .ZN(
        n12116) );
  AOI21_X1 U13990 ( .B1(n14623), .B2(n12117), .A(n12116), .ZN(n12118) );
  INV_X1 U13991 ( .A(n12118), .ZN(P2_U3264) );
  XNOR2_X1 U13992 ( .A(n12119), .B(n13405), .ZN(n12239) );
  XNOR2_X1 U13993 ( .A(n12239), .B(n13516), .ZN(n12125) );
  INV_X1 U13994 ( .A(n12120), .ZN(n12121) );
  OAI21_X1 U13995 ( .B1(n12125), .B2(n12124), .A(n12241), .ZN(n12126) );
  NAND2_X1 U13996 ( .A1(n12126), .A2(n13495), .ZN(n12131) );
  INV_X1 U13997 ( .A(n13470), .ZN(n13498) );
  OAI22_X1 U13998 ( .A1(n12127), .A2(n13500), .B1(n13507), .B2(n16142), .ZN(
        n12128) );
  AOI211_X1 U13999 ( .C1(n13498), .C2(n13515), .A(n12129), .B(n12128), .ZN(
        n12130) );
  OAI211_X1 U14000 ( .C1(n12159), .C2(n12627), .A(n12131), .B(n12130), .ZN(
        P3_U3171) );
  INV_X1 U14001 ( .A(n12727), .ZN(n12719) );
  OAI222_X1 U14002 ( .A1(n15773), .A2(n12132), .B1(n15771), .B2(n12719), .C1(
        P1_U3086), .C2(n15343), .ZN(P1_U3336) );
  INV_X1 U14003 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n12134) );
  MUX2_X1 U14004 ( .A(n12134), .B(n12133), .S(n14948), .Z(n12137) );
  NAND2_X1 U14005 ( .A1(n14919), .A2(n12135), .ZN(n12136) );
  OAI211_X1 U14006 ( .C1(n8630), .C2(n14951), .A(n12137), .B(n12136), .ZN(
        P2_U3433) );
  XNOR2_X1 U14007 ( .A(n12139), .B(n12138), .ZN(n16184) );
  INV_X1 U14008 ( .A(n12499), .ZN(n14474) );
  AOI22_X1 U14009 ( .A1(n14647), .A2(n14476), .B1(n14474), .B2(n14791), .ZN(
        n12143) );
  OAI211_X1 U14010 ( .C1(n12141), .C2(n12140), .A(n9112), .B(n12331), .ZN(
        n12142) );
  OAI211_X1 U14011 ( .C1(n16184), .C2(n14876), .A(n12143), .B(n12142), .ZN(
        n16187) );
  NAND2_X1 U14012 ( .A1(n16187), .A2(n14805), .ZN(n12151) );
  INV_X1 U14013 ( .A(n12144), .ZN(n12233) );
  OAI22_X1 U14014 ( .A1(n14805), .A2(n10885), .B1(n12233), .B2(n14697), .ZN(
        n12148) );
  INV_X1 U14015 ( .A(n12145), .ZN(n12336) );
  OAI211_X1 U14016 ( .C1(n16186), .C2(n12146), .A(n12336), .B(n14267), .ZN(
        n16185) );
  NOR2_X1 U14017 ( .A1(n16185), .A2(n14751), .ZN(n12147) );
  AOI211_X1 U14018 ( .C1(n14747), .C2(n12149), .A(n12148), .B(n12147), .ZN(
        n12150) );
  OAI211_X1 U14019 ( .C1(n16184), .C2(n14806), .A(n12151), .B(n12150), .ZN(
        P2_U3255) );
  INV_X1 U14020 ( .A(n13137), .ZN(n12152) );
  OR2_X1 U14021 ( .A1(n13136), .A2(n12152), .ZN(n13264) );
  XNOR2_X1 U14022 ( .A(n12153), .B(n13264), .ZN(n16143) );
  INV_X1 U14023 ( .A(n12154), .ZN(n16050) );
  NAND2_X1 U14024 ( .A1(n16131), .A2(n16050), .ZN(n14023) );
  XNOR2_X1 U14025 ( .A(n12155), .B(n13264), .ZN(n12156) );
  NAND2_X1 U14026 ( .A1(n12156), .A2(n14103), .ZN(n12158) );
  AOI22_X1 U14027 ( .A1(n14108), .A2(n13517), .B1(n13515), .B2(n14107), .ZN(
        n12157) );
  OAI211_X1 U14028 ( .C1(n16143), .C2(n14017), .A(n12158), .B(n12157), .ZN(
        n16145) );
  NAND2_X1 U14029 ( .A1(n16145), .A2(n16131), .ZN(n12162) );
  OAI22_X1 U14030 ( .A1(n16126), .A2(n16142), .B1(n12159), .B2(n16128), .ZN(
        n12160) );
  AOI21_X1 U14031 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n16052), .A(n12160), .ZN(
        n12161) );
  OAI211_X1 U14032 ( .C1(n16143), .C2(n14023), .A(n12162), .B(n12161), .ZN(
        P3_U3224) );
  XNOR2_X1 U14033 ( .A(n12163), .B(n13023), .ZN(n16168) );
  INV_X1 U14034 ( .A(n12164), .ZN(n12167) );
  OAI211_X1 U14035 ( .C1(n16172), .C2(n12166), .A(n16153), .B(n12165), .ZN(
        n16170) );
  OAI211_X1 U14036 ( .C1(n16168), .C2(n12168), .A(n12167), .B(n16170), .ZN(
        n12180) );
  AOI22_X1 U14037 ( .A1(n12793), .A2(n15617), .B1(n16011), .B2(n12169), .ZN(
        n12170) );
  OAI21_X1 U14038 ( .B1(n16168), .B2(n15598), .A(n12170), .ZN(n12179) );
  AOI21_X1 U14039 ( .B1(n12172), .B2(n12171), .A(n16074), .ZN(n12174) );
  NAND2_X1 U14040 ( .A1(n12174), .A2(n12173), .ZN(n16173) );
  INV_X1 U14041 ( .A(n12175), .ZN(n12176) );
  NAND2_X1 U14042 ( .A1(n16173), .A2(n12176), .ZN(n12177) );
  MUX2_X1 U14043 ( .A(n12177), .B(P1_REG2_REG_10__SCAN_IN), .S(n16022), .Z(
        n12178) );
  AOI211_X1 U14044 ( .C1(n15429), .C2(n12180), .A(n12179), .B(n12178), .ZN(
        n12181) );
  INV_X1 U14045 ( .A(n12181), .ZN(P1_U3283) );
  NAND2_X1 U14046 ( .A1(n12797), .A2(n12184), .ZN(n12182) );
  OR2_X1 U14047 ( .A1(n12797), .A2(n12184), .ZN(n12185) );
  NAND2_X1 U14048 ( .A1(n12186), .A2(n12185), .ZN(n12342) );
  NAND2_X1 U14049 ( .A1(n12187), .A2(n12998), .ZN(n12189) );
  AOI22_X1 U14050 ( .A1(n12836), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n12835), 
        .B2(n15930), .ZN(n12188) );
  XNOR2_X1 U14051 ( .A(n12801), .B(n15226), .ZN(n13025) );
  NAND2_X1 U14052 ( .A1(n12342), .A2(n13025), .ZN(n12191) );
  INV_X1 U14053 ( .A(n15226), .ZN(n12376) );
  OR2_X1 U14054 ( .A1(n12801), .A2(n12376), .ZN(n12190) );
  NAND2_X1 U14055 ( .A1(n12192), .A2(n12998), .ZN(n12195) );
  AOI22_X1 U14056 ( .A1(n12836), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n12835), 
        .B2(n12193), .ZN(n12194) );
  NAND2_X1 U14057 ( .A1(n12875), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n12203) );
  NAND2_X1 U14058 ( .A1(n12966), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n12202) );
  INV_X1 U14059 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n12196) );
  OAI21_X1 U14060 ( .B1(n12198), .B2(n12196), .A(n12197), .ZN(n12199) );
  AND2_X1 U14061 ( .A1(n12199), .A2(n12211), .ZN(n12591) );
  NAND2_X1 U14062 ( .A1(n12965), .A2(n12591), .ZN(n12201) );
  NAND2_X1 U14063 ( .A1(n12982), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U14064 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n15225) );
  XNOR2_X1 U14065 ( .A(n12805), .B(n12584), .ZN(n13027) );
  INV_X1 U14066 ( .A(n13027), .ZN(n12517) );
  XNOR2_X1 U14067 ( .A(n12518), .B(n12517), .ZN(n12413) );
  NOR2_X1 U14068 ( .A1(n12797), .A2(n15227), .ZN(n12204) );
  NAND2_X1 U14069 ( .A1(n12797), .A2(n15227), .ZN(n12206) );
  NAND2_X1 U14070 ( .A1(n12208), .A2(n12207), .ZN(n12343) );
  OR2_X1 U14071 ( .A1(n12801), .A2(n15226), .ZN(n12209) );
  NAND2_X1 U14072 ( .A1(n12343), .A2(n12209), .ZN(n12210) );
  NAND2_X1 U14073 ( .A1(n12210), .A2(n13027), .ZN(n12525) );
  OAI21_X1 U14074 ( .B1(n12210), .B2(n13027), .A(n12525), .ZN(n12411) );
  NAND2_X1 U14075 ( .A1(n12411), .A2(n15620), .ZN(n12223) );
  NAND2_X1 U14076 ( .A1(n12594), .A2(n7206), .ZN(n12528) );
  OAI211_X1 U14077 ( .C1(n12594), .C2(n7206), .A(n16153), .B(n12528), .ZN(
        n12409) );
  NAND2_X1 U14078 ( .A1(n15226), .A2(n15500), .ZN(n12218) );
  NAND2_X1 U14079 ( .A1(n12875), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n12216) );
  NAND2_X1 U14080 ( .A1(n12966), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12215) );
  INV_X1 U14081 ( .A(n12530), .ZN(n12532) );
  NAND2_X1 U14082 ( .A1(n12211), .A2(n12711), .ZN(n12212) );
  AND2_X1 U14083 ( .A1(n12532), .A2(n12212), .ZN(n12713) );
  NAND2_X1 U14084 ( .A1(n12965), .A2(n12713), .ZN(n12214) );
  NAND2_X1 U14085 ( .A1(n12982), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n12213) );
  NAND4_X1 U14086 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n15224) );
  NAND2_X1 U14087 ( .A1(n15224), .A2(n15583), .ZN(n12217) );
  AND2_X1 U14088 ( .A1(n12218), .A2(n12217), .ZN(n12589) );
  NAND2_X1 U14089 ( .A1(n16011), .A2(n12591), .ZN(n12219) );
  OAI211_X1 U14090 ( .C1(n12409), .C2(n12730), .A(n12589), .B(n12219), .ZN(
        n12221) );
  OAI22_X1 U14091 ( .A1(n12594), .A2(n16014), .B1(n10946), .B2(n15611), .ZN(
        n12220) );
  AOI21_X1 U14092 ( .B1(n12221), .B2(n15611), .A(n12220), .ZN(n12222) );
  OAI211_X1 U14093 ( .C1(n12413), .C2(n15622), .A(n12223), .B(n12222), .ZN(
        P1_U3280) );
  NOR2_X1 U14094 ( .A1(n12335), .A2(n14267), .ZN(n12225) );
  XNOR2_X1 U14095 ( .A(n16186), .B(n14304), .ZN(n12224) );
  NOR2_X1 U14096 ( .A1(n12224), .A2(n12225), .ZN(n12267) );
  AOI21_X1 U14097 ( .B1(n12225), .B2(n12224), .A(n12267), .ZN(n12230) );
  INV_X1 U14098 ( .A(n12226), .ZN(n12227) );
  OAI21_X1 U14099 ( .B1(n12230), .B2(n12229), .A(n12268), .ZN(n12231) );
  NAND2_X1 U14100 ( .A1(n12231), .A2(n14420), .ZN(n12237) );
  INV_X1 U14101 ( .A(n12232), .ZN(n12235) );
  OAI22_X1 U14102 ( .A1(n14404), .A2(n12499), .B1(n14403), .B2(n12233), .ZN(
        n12234) );
  AOI211_X1 U14103 ( .C1(n14443), .C2(n14476), .A(n12235), .B(n12234), .ZN(
        n12236) );
  OAI211_X1 U14104 ( .C1(n16186), .C2(n14462), .A(n12237), .B(n12236), .ZN(
        P2_U3189) );
  NAND2_X1 U14105 ( .A1(n12239), .A2(n12238), .ZN(n12240) );
  AND2_X1 U14106 ( .A1(n12241), .A2(n12240), .ZN(n12243) );
  XNOR2_X1 U14107 ( .A(n16162), .B(n13405), .ZN(n12354) );
  XOR2_X1 U14108 ( .A(n13515), .B(n12354), .Z(n12242) );
  OAI211_X1 U14109 ( .C1(n12243), .C2(n12242), .A(n13495), .B(n12356), .ZN(
        n12250) );
  NAND2_X1 U14110 ( .A1(n12630), .A2(n13516), .ZN(n12248) );
  NAND2_X1 U14111 ( .A1(n13498), .A2(n13514), .ZN(n12247) );
  NAND2_X1 U14112 ( .A1(n12259), .A2(n13411), .ZN(n12246) );
  INV_X1 U14113 ( .A(n12244), .ZN(n12245) );
  AND4_X1 U14114 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n12245), .ZN(
        n12249) );
  OAI211_X1 U14115 ( .C1(n12256), .C2(n12627), .A(n12250), .B(n12249), .ZN(
        P3_U3157) );
  XNOR2_X1 U14116 ( .A(n12251), .B(n8041), .ZN(n16164) );
  XNOR2_X1 U14117 ( .A(n12252), .B(n8041), .ZN(n12253) );
  NAND2_X1 U14118 ( .A1(n12253), .A2(n14103), .ZN(n12255) );
  AOI22_X1 U14119 ( .A1(n14108), .A2(n13516), .B1(n13514), .B2(n14107), .ZN(
        n12254) );
  OAI211_X1 U14120 ( .C1(n14017), .C2(n16164), .A(n12255), .B(n12254), .ZN(
        n16166) );
  NAND2_X1 U14121 ( .A1(n16166), .A2(n16131), .ZN(n12261) );
  OAI22_X1 U14122 ( .A1(n16131), .A2(n12257), .B1(n12256), .B2(n16128), .ZN(
        n12258) );
  AOI21_X1 U14123 ( .B1(n12259), .B2(n14065), .A(n12258), .ZN(n12260) );
  OAI211_X1 U14124 ( .C1(n16164), .C2(n14023), .A(n12261), .B(n12260), .ZN(
        P3_U3223) );
  INV_X1 U14125 ( .A(n12262), .ZN(n12263) );
  OAI222_X1 U14126 ( .A1(P3_U3151), .A2(n12264), .B1(n13319), .B2(n12263), 
        .C1(n13534), .C2(n10650), .ZN(P3_U3267) );
  INV_X1 U14127 ( .A(n12265), .ZN(n12266) );
  OAI222_X1 U14128 ( .A1(P3_U3151), .A2(n13309), .B1(n13319), .B2(n12266), 
        .C1(n13632), .C2(n10650), .ZN(P3_U3268) );
  NOR2_X1 U14129 ( .A1(n12499), .A2(n14267), .ZN(n12491) );
  XNOR2_X1 U14130 ( .A(n12425), .B(n14352), .ZN(n12493) );
  XOR2_X1 U14131 ( .A(n12491), .B(n12493), .Z(n12494) );
  XNOR2_X1 U14132 ( .A(n12495), .B(n12494), .ZN(n12273) );
  INV_X1 U14133 ( .A(n14795), .ZN(n14473) );
  AOI22_X1 U14134 ( .A1(n14444), .A2(n14473), .B1(n14459), .B2(n12337), .ZN(
        n12270) );
  OAI211_X1 U14135 ( .C1(n12335), .C2(n14402), .A(n12270), .B(n12269), .ZN(
        n12271) );
  AOI21_X1 U14136 ( .B1(n12422), .B2(n14423), .A(n12271), .ZN(n12272) );
  OAI21_X1 U14137 ( .B1(n12273), .B2(n14449), .A(n12272), .ZN(P2_U3208) );
  AOI21_X1 U14138 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n12652), .A(n12274), 
        .ZN(n12277) );
  XNOR2_X1 U14139 ( .A(n12823), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n12276) );
  NOR2_X1 U14140 ( .A1(n12277), .A2(n12276), .ZN(n12693) );
  AOI211_X1 U14141 ( .C1(n12277), .C2(n12276), .A(n12275), .B(n12693), .ZN(
        n12287) );
  OAI21_X1 U14142 ( .B1(n12007), .B2(n12279), .A(n12278), .ZN(n12281) );
  XOR2_X1 U14143 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n12823), .Z(n12280) );
  NAND2_X1 U14144 ( .A1(n12280), .A2(n12281), .ZN(n12691) );
  OAI211_X1 U14145 ( .C1(n12281), .C2(n12280), .A(n12691), .B(n15931), .ZN(
        n12284) );
  AND2_X1 U14146 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n12282) );
  AOI21_X1 U14147 ( .B1(n15914), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n12282), 
        .ZN(n12283) );
  OAI211_X1 U14148 ( .C1(n15337), .C2(n12285), .A(n12284), .B(n12283), .ZN(
        n12286) );
  OR2_X1 U14149 ( .A1(n12287), .A2(n12286), .ZN(P1_U3260) );
  INV_X1 U14150 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n12288) );
  OAI22_X1 U14151 ( .A1(n14951), .A2(n12289), .B1(n14948), .B2(n12288), .ZN(
        n12290) );
  AOI21_X1 U14152 ( .B1(n12291), .B2(n14919), .A(n12290), .ZN(n12292) );
  OAI21_X1 U14153 ( .B1(n12293), .B2(n16209), .A(n12292), .ZN(P2_U3457) );
  INV_X1 U14154 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n12294) );
  OAI22_X1 U14155 ( .A1(n14951), .A2(n12295), .B1(n14948), .B2(n12294), .ZN(
        n12296) );
  AOI21_X1 U14156 ( .B1(n12297), .B2(n14919), .A(n12296), .ZN(n12298) );
  OAI21_X1 U14157 ( .B1(n12299), .B2(n16209), .A(n12298), .ZN(P2_U3451) );
  AOI21_X1 U14158 ( .B1(n12301), .B2(n12642), .A(n12451), .ZN(n12319) );
  AOI21_X1 U14159 ( .B1(n9571), .B2(n12303), .A(n12458), .ZN(n12304) );
  OR2_X1 U14160 ( .A1(n12304), .A2(n13899), .ZN(n12318) );
  INV_X1 U14161 ( .A(n12311), .ZN(n12466) );
  OR2_X1 U14162 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9351), .ZN(n12626) );
  OAI21_X1 U14163 ( .B1(n13842), .B2(n12305), .A(n12626), .ZN(n12316) );
  NAND2_X1 U14164 ( .A1(n12306), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12307) );
  MUX2_X1 U14165 ( .A(n12308), .B(n12307), .S(n13309), .Z(n12309) );
  MUX2_X1 U14166 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13309), .Z(n12465) );
  XNOR2_X1 U14167 ( .A(n12465), .B(n12311), .ZN(n12312) );
  NAND2_X1 U14168 ( .A1(n12313), .A2(n12312), .ZN(n12314) );
  AOI21_X1 U14169 ( .B1(n12469), .B2(n12314), .A(n13877), .ZN(n12315) );
  AOI211_X1 U14170 ( .C1(n13874), .C2(n12466), .A(n12316), .B(n12315), .ZN(
        n12317) );
  OAI211_X1 U14171 ( .C1(n12319), .C2(n13895), .A(n12318), .B(n12317), .ZN(
        P3_U3195) );
  INV_X1 U14172 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n12320) );
  OAI22_X1 U14173 ( .A1(n14951), .A2(n12321), .B1(n14948), .B2(n12320), .ZN(
        n12322) );
  AOI21_X1 U14174 ( .B1(n12323), .B2(n14948), .A(n12322), .ZN(n12324) );
  INV_X1 U14175 ( .A(n12324), .ZN(P2_U3448) );
  OAI21_X1 U14176 ( .B1(n12327), .B2(n12326), .A(n12325), .ZN(n12418) );
  INV_X1 U14177 ( .A(n12328), .ZN(n12333) );
  AOI21_X1 U14178 ( .B1(n12331), .B2(n12330), .A(n12329), .ZN(n12332) );
  NOR2_X1 U14179 ( .A1(n12333), .A2(n12332), .ZN(n12334) );
  OAI222_X1 U14180 ( .A1(n14600), .A2(n14795), .B1(n14794), .B2(n12335), .C1(
        n14719), .C2(n12334), .ZN(n12419) );
  NAND2_X1 U14181 ( .A1(n12419), .A2(n14805), .ZN(n12341) );
  AOI211_X1 U14182 ( .C1(n12422), .C2(n12336), .A(n14300), .B(n12401), .ZN(
        n12420) );
  AOI22_X1 U14183 ( .A1(n16082), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n12337), 
        .B2(n16080), .ZN(n12338) );
  OAI21_X1 U14184 ( .B1(n12425), .B2(n16085), .A(n12338), .ZN(n12339) );
  AOI21_X1 U14185 ( .B1(n12420), .B2(n16088), .A(n12339), .ZN(n12340) );
  OAI211_X1 U14186 ( .C1(n12418), .C2(n16062), .A(n12341), .B(n12340), .ZN(
        P2_U3254) );
  XOR2_X1 U14187 ( .A(n12342), .B(n13025), .Z(n12348) );
  INV_X1 U14188 ( .A(n12343), .ZN(n12344) );
  AOI21_X1 U14189 ( .B1(n13025), .B2(n12345), .A(n12344), .ZN(n12445) );
  AOI22_X1 U14190 ( .A1(n15582), .A2(n15227), .B1(n15225), .B2(n15437), .ZN(
        n12346) );
  OAI21_X1 U14191 ( .B1(n12445), .B2(n16002), .A(n12346), .ZN(n12347) );
  AOI21_X1 U14192 ( .B1(n12348), .B2(n15723), .A(n12347), .ZN(n12444) );
  AOI21_X1 U14193 ( .B1(n12801), .B2(n12349), .A(n7206), .ZN(n12442) );
  AOI22_X1 U14194 ( .A1(n16022), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12512), 
        .B2(n16011), .ZN(n12350) );
  OAI21_X1 U14195 ( .B1(n8015), .B2(n16014), .A(n12350), .ZN(n12352) );
  NOR2_X1 U14196 ( .A1(n12445), .A2(n15598), .ZN(n12351) );
  AOI211_X1 U14197 ( .C1(n12442), .C2(n15601), .A(n12352), .B(n12351), .ZN(
        n12353) );
  OAI21_X1 U14198 ( .B1(n16022), .B2(n12444), .A(n12353), .ZN(P1_U3281) );
  INV_X1 U14199 ( .A(n13515), .ZN(n12431) );
  OR2_X1 U14200 ( .A1(n12357), .A2(n13405), .ZN(n12547) );
  INV_X1 U14201 ( .A(n12358), .ZN(n12360) );
  INV_X1 U14202 ( .A(n13144), .ZN(n12359) );
  NAND2_X1 U14203 ( .A1(n13145), .A2(n13405), .ZN(n12548) );
  OAI22_X1 U14204 ( .A1(n12547), .A2(n12360), .B1(n12359), .B2(n12548), .ZN(
        n12549) );
  XNOR2_X1 U14205 ( .A(n12550), .B(n12549), .ZN(n12368) );
  AOI21_X1 U14206 ( .B1(n13498), .B2(n13513), .A(n12361), .ZN(n12364) );
  INV_X1 U14207 ( .A(n12435), .ZN(n12362) );
  NAND2_X1 U14208 ( .A1(n13503), .A2(n12362), .ZN(n12363) );
  OAI211_X1 U14209 ( .C1(n12431), .C2(n13500), .A(n12364), .B(n12363), .ZN(
        n12365) );
  AOI21_X1 U14210 ( .B1(n12366), .B2(n13411), .A(n12365), .ZN(n12367) );
  OAI21_X1 U14211 ( .B1(n12368), .B2(n13440), .A(n12367), .ZN(P3_U3176) );
  AOI22_X1 U14212 ( .A1(n12797), .A2(n15062), .B1(n11123), .B2(n15227), .ZN(
        n12369) );
  XNOR2_X1 U14213 ( .A(n12369), .B(n15065), .ZN(n12510) );
  AOI22_X1 U14214 ( .A1(n12797), .A2(n11123), .B1(n15050), .B2(n15227), .ZN(
        n12511) );
  XNOR2_X1 U14215 ( .A(n12510), .B(n12511), .ZN(n12374) );
  AOI21_X1 U14216 ( .B1(n12374), .B2(n12373), .A(n7351), .ZN(n12383) );
  OAI22_X1 U14217 ( .A1(n15193), .A2(n12376), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12375), .ZN(n12381) );
  INV_X1 U14218 ( .A(n12377), .ZN(n12379) );
  OAI22_X1 U14219 ( .A1(n15192), .A2(n12379), .B1(n12378), .B2(n15191), .ZN(
        n12380) );
  AOI211_X1 U14220 ( .C1(n12797), .C2(n15196), .A(n12381), .B(n12380), .ZN(
        n12382) );
  OAI21_X1 U14221 ( .B1(n12383), .B2(n15205), .A(n12382), .ZN(P1_U3236) );
  INV_X1 U14222 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U14223 ( .A1(n12384), .A2(n16153), .B1(n12797), .B2(n16151), .ZN(
        n12385) );
  OAI211_X1 U14224 ( .C1(n15732), .C2(n12387), .A(n12386), .B(n12385), .ZN(
        n12390) );
  NAND2_X1 U14225 ( .A1(n12390), .A2(n16183), .ZN(n12388) );
  OAI21_X1 U14226 ( .B1(n16183), .B2(n12389), .A(n12388), .ZN(P1_U3492) );
  NAND2_X1 U14227 ( .A1(n12390), .A2(n16179), .ZN(n12391) );
  OAI21_X1 U14228 ( .B1(n16179), .B2(n12392), .A(n12391), .ZN(P1_U3539) );
  INV_X1 U14229 ( .A(n12393), .ZN(n12395) );
  OAI222_X1 U14230 ( .A1(P3_U3151), .A2(n12397), .B1(n12396), .B2(n12395), 
        .C1(n12394), .C2(n10650), .ZN(P3_U3266) );
  OAI21_X1 U14231 ( .B1(n12405), .B2(n12399), .A(n12398), .ZN(n12400) );
  AOI222_X1 U14232 ( .A1(n9112), .A2(n12400), .B1(n14472), .B2(n14791), .C1(
        n14474), .C2(n14647), .ZN(n16200) );
  OAI211_X1 U14233 ( .C1(n12401), .C2(n16202), .A(n14267), .B(n14801), .ZN(
        n16199) );
  INV_X1 U14234 ( .A(n16199), .ZN(n12404) );
  AOI22_X1 U14235 ( .A1(n16082), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12500), 
        .B2(n16080), .ZN(n12402) );
  OAI21_X1 U14236 ( .B1(n16202), .B2(n16085), .A(n12402), .ZN(n12403) );
  AOI21_X1 U14237 ( .B1(n12404), .B2(n16088), .A(n12403), .ZN(n12408) );
  XNOR2_X1 U14238 ( .A(n12406), .B(n12405), .ZN(n16205) );
  NAND2_X1 U14239 ( .A1(n16205), .A2(n14753), .ZN(n12407) );
  OAI211_X1 U14240 ( .C1(n16200), .C2(n16082), .A(n12408), .B(n12407), .ZN(
        P2_U3253) );
  OAI211_X1 U14241 ( .C1(n12594), .C2(n16171), .A(n12409), .B(n12589), .ZN(
        n12410) );
  AOI21_X1 U14242 ( .B1(n12411), .B2(n16176), .A(n12410), .ZN(n12412) );
  OAI21_X1 U14243 ( .B1(n16074), .B2(n12413), .A(n12412), .ZN(n12415) );
  NAND2_X1 U14244 ( .A1(n12415), .A2(n16179), .ZN(n12414) );
  OAI21_X1 U14245 ( .B1(n16179), .B2(n10939), .A(n12414), .ZN(P1_U3541) );
  INV_X1 U14246 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U14247 ( .A1(n12415), .A2(n16183), .ZN(n12416) );
  OAI21_X1 U14248 ( .B1(n16183), .B2(n12417), .A(n12416), .ZN(P1_U3498) );
  INV_X1 U14249 ( .A(n12418), .ZN(n12421) );
  AOI211_X1 U14250 ( .C1(n12421), .C2(n16204), .A(n12420), .B(n12419), .ZN(
        n12428) );
  INV_X1 U14251 ( .A(n14896), .ZN(n14816) );
  AOI22_X1 U14252 ( .A1(n12422), .A2(n14816), .B1(n16206), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n12423) );
  OAI21_X1 U14253 ( .B1(n12428), .B2(n16206), .A(n12423), .ZN(P2_U3510) );
  INV_X1 U14254 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n12424) );
  OAI22_X1 U14255 ( .A1(n12425), .A2(n14951), .B1(n14948), .B2(n12424), .ZN(
        n12426) );
  INV_X1 U14256 ( .A(n12426), .ZN(n12427) );
  OAI21_X1 U14257 ( .B1(n12428), .B2(n16209), .A(n12427), .ZN(P2_U3463) );
  XOR2_X1 U14258 ( .A(n12429), .B(n13273), .Z(n12430) );
  OAI222_X1 U14259 ( .A1(n16032), .A2(n12432), .B1(n16034), .B2(n12431), .C1(
        n12430), .C2(n16039), .ZN(n16194) );
  INV_X1 U14260 ( .A(n16194), .ZN(n12439) );
  OAI21_X1 U14261 ( .B1(n12434), .B2(n13273), .A(n12433), .ZN(n16196) );
  NOR2_X1 U14262 ( .A1(n16193), .A2(n16126), .ZN(n12437) );
  OAI22_X1 U14263 ( .A1(n16131), .A2(n9534), .B1(n12435), .B2(n16128), .ZN(
        n12436) );
  AOI211_X1 U14264 ( .C1(n16196), .C2(n14099), .A(n12437), .B(n12436), .ZN(
        n12438) );
  OAI21_X1 U14265 ( .B1(n12439), .B2(n16052), .A(n12438), .ZN(P3_U3222) );
  INV_X1 U14266 ( .A(n12847), .ZN(n12440) );
  OAI222_X1 U14267 ( .A1(n15773), .A2(n12848), .B1(n15771), .B2(n12440), .C1(
        n12992), .C2(n7190), .ZN(P1_U3335) );
  OAI222_X1 U14268 ( .A1(n14970), .A2(n12441), .B1(P2_U3088), .B2(n8212), .C1(
        n14968), .C2(n12440), .ZN(P2_U3307) );
  INV_X1 U14269 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U14270 ( .A1(n12442), .A2(n16153), .B1(n12801), .B2(n16151), .ZN(
        n12443) );
  OAI211_X1 U14271 ( .C1(n12445), .C2(n16116), .A(n12444), .B(n12443), .ZN(
        n12448) );
  NAND2_X1 U14272 ( .A1(n12448), .A2(n16183), .ZN(n12446) );
  OAI21_X1 U14273 ( .B1(n16183), .B2(n12447), .A(n12446), .ZN(P1_U3495) );
  NAND2_X1 U14274 ( .A1(n12448), .A2(n16179), .ZN(n12449) );
  OAI21_X1 U14275 ( .B1(n16179), .B2(n10940), .A(n12449), .ZN(P1_U3540) );
  NOR2_X1 U14276 ( .A1(n12466), .A2(n12450), .ZN(n12452) );
  NAND2_X1 U14277 ( .A1(n13797), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13791) );
  OR2_X1 U14278 ( .A1(n13797), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12453) );
  NAND2_X1 U14279 ( .A1(n13791), .A2(n12453), .ZN(n12455) );
  INV_X1 U14280 ( .A(n13792), .ZN(n12454) );
  AOI21_X1 U14281 ( .B1(n12456), .B2(n12455), .A(n12454), .ZN(n12478) );
  NOR2_X1 U14282 ( .A1(n12466), .A2(n12457), .ZN(n12459) );
  INV_X1 U14283 ( .A(n12462), .ZN(n12464) );
  NAND2_X1 U14284 ( .A1(n13797), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13788) );
  OR2_X1 U14285 ( .A1(n13797), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12460) );
  NAND2_X1 U14286 ( .A1(n13788), .A2(n12460), .ZN(n12461) );
  INV_X1 U14287 ( .A(n12461), .ZN(n12463) );
  OAI21_X1 U14288 ( .B1(n12464), .B2(n12463), .A(n13789), .ZN(n12476) );
  INV_X1 U14289 ( .A(n12465), .ZN(n12467) );
  NAND2_X1 U14290 ( .A1(n12467), .A2(n12466), .ZN(n12468) );
  MUX2_X1 U14291 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13309), .Z(n13798) );
  INV_X1 U14292 ( .A(n13797), .ZN(n12470) );
  XNOR2_X1 U14293 ( .A(n13798), .B(n12470), .ZN(n12471) );
  OAI211_X1 U14294 ( .C1(n12472), .C2(n12471), .A(n13800), .B(n13897), .ZN(
        n12474) );
  INV_X1 U14295 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13576) );
  NOR2_X1 U14296 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13576), .ZN(n13382) );
  AOI21_X1 U14297 ( .B1(n15817), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13382), 
        .ZN(n12473) );
  OAI211_X1 U14298 ( .C1(n13889), .C2(n13797), .A(n12474), .B(n12473), .ZN(
        n12475) );
  AOI21_X1 U14299 ( .B1(n12476), .B2(n13865), .A(n12475), .ZN(n12477) );
  OAI21_X1 U14300 ( .B1(n12478), .B2(n13895), .A(n12477), .ZN(P3_U3196) );
  XNOR2_X1 U14301 ( .A(n12479), .B(n13272), .ZN(n14189) );
  INV_X1 U14302 ( .A(n14189), .ZN(n12488) );
  XNOR2_X1 U14303 ( .A(n12480), .B(n13272), .ZN(n12483) );
  AOI22_X1 U14304 ( .A1(n14109), .A2(n14107), .B1(n14108), .B2(n13514), .ZN(
        n12482) );
  INV_X1 U14305 ( .A(n14017), .ZN(n16212) );
  NAND2_X1 U14306 ( .A1(n14189), .A2(n16212), .ZN(n12481) );
  OAI211_X1 U14307 ( .C1(n12483), .C2(n16039), .A(n12482), .B(n12481), .ZN(
        n14188) );
  NAND2_X1 U14308 ( .A1(n14188), .A2(n16131), .ZN(n12487) );
  OAI22_X1 U14309 ( .A1(n16131), .A2(n12484), .B1(n12560), .B2(n16128), .ZN(
        n12485) );
  AOI21_X1 U14310 ( .B1(n14065), .B2(n14187), .A(n12485), .ZN(n12486) );
  OAI211_X1 U14311 ( .C1(n12488), .C2(n14023), .A(n12487), .B(n12486), .ZN(
        P3_U3221) );
  XNOR2_X1 U14312 ( .A(n16202), .B(n14352), .ZN(n12490) );
  OR2_X1 U14313 ( .A1(n14795), .A2(n14267), .ZN(n12489) );
  NAND2_X1 U14314 ( .A1(n12490), .A2(n12489), .ZN(n12567) );
  OAI21_X1 U14315 ( .B1(n12490), .B2(n12489), .A(n12567), .ZN(n12498) );
  INV_X1 U14316 ( .A(n12491), .ZN(n12492) );
  INV_X1 U14317 ( .A(n12568), .ZN(n12497) );
  AOI21_X1 U14318 ( .B1(n12498), .B2(n12496), .A(n12497), .ZN(n12506) );
  NAND2_X1 U14319 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n15884)
         );
  OAI21_X1 U14320 ( .B1(n14402), .B2(n12499), .A(n15884), .ZN(n12503) );
  INV_X1 U14321 ( .A(n12500), .ZN(n12501) );
  OAI22_X1 U14322 ( .A1(n14404), .A2(n14327), .B1(n14403), .B2(n12501), .ZN(
        n12502) );
  AOI211_X1 U14323 ( .C1(n12504), .C2(n14423), .A(n12503), .B(n12502), .ZN(
        n12505) );
  OAI21_X1 U14324 ( .B1(n12506), .B2(n14449), .A(n12505), .ZN(P2_U3196) );
  NAND2_X1 U14325 ( .A1(n12801), .A2(n15062), .ZN(n12508) );
  NAND2_X1 U14326 ( .A1(n15226), .A2(n11123), .ZN(n12507) );
  NAND2_X1 U14327 ( .A1(n12508), .A2(n12507), .ZN(n12509) );
  XNOR2_X1 U14328 ( .A(n12509), .B(n15065), .ZN(n12579) );
  AOI22_X1 U14329 ( .A1(n12801), .A2(n11123), .B1(n15050), .B2(n15226), .ZN(
        n12581) );
  XNOR2_X1 U14330 ( .A(n12579), .B(n12581), .ZN(n12582) );
  XOR2_X1 U14331 ( .A(n12582), .B(n12583), .Z(n12516) );
  AOI22_X1 U14332 ( .A1(n15184), .A2(n15227), .B1(n15216), .B2(n12512), .ZN(
        n12513) );
  NAND2_X1 U14333 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n15933)
         );
  OAI211_X1 U14334 ( .C1(n12584), .C2(n15193), .A(n12513), .B(n15933), .ZN(
        n12514) );
  AOI21_X1 U14335 ( .B1(n12801), .B2(n15196), .A(n12514), .ZN(n12515) );
  OAI21_X1 U14336 ( .B1(n12516), .B2(n15205), .A(n12515), .ZN(P1_U3224) );
  OR2_X1 U14337 ( .A1(n12805), .A2(n12584), .ZN(n12519) );
  NAND2_X1 U14338 ( .A1(n12520), .A2(n12998), .ZN(n12523) );
  AOI22_X1 U14339 ( .A1(n12836), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n12835), 
        .B2(n12521), .ZN(n12522) );
  XNOR2_X1 U14340 ( .A(n15733), .B(n15224), .ZN(n13028) );
  XNOR2_X1 U14341 ( .A(n12603), .B(n13028), .ZN(n15740) );
  OR2_X1 U14342 ( .A1(n12805), .A2(n15225), .ZN(n12524) );
  INV_X1 U14343 ( .A(n12615), .ZN(n12526) );
  AOI21_X1 U14344 ( .B1(n13028), .B2(n12527), .A(n12526), .ZN(n15738) );
  INV_X1 U14345 ( .A(n15601), .ZN(n16015) );
  INV_X1 U14346 ( .A(n12528), .ZN(n12529) );
  INV_X1 U14347 ( .A(n15733), .ZN(n12541) );
  OAI21_X1 U14348 ( .B1(n12529), .B2(n12541), .A(n12600), .ZN(n15736) );
  NAND2_X1 U14349 ( .A1(n15225), .A2(n15500), .ZN(n12539) );
  NAND2_X1 U14350 ( .A1(n12875), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n12537) );
  NAND2_X1 U14351 ( .A1(n12966), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n12536) );
  INV_X1 U14352 ( .A(n12604), .ZN(n12605) );
  INV_X1 U14353 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U14354 ( .A1(n12532), .A2(n12531), .ZN(n12533) );
  AND2_X1 U14355 ( .A1(n12605), .A2(n12533), .ZN(n15217) );
  NAND2_X1 U14356 ( .A1(n12965), .A2(n15217), .ZN(n12535) );
  NAND2_X1 U14357 ( .A1(n12982), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n12534) );
  NAND4_X1 U14358 ( .A1(n12537), .A2(n12536), .A3(n12535), .A4(n12534), .ZN(
        n15223) );
  NAND2_X1 U14359 ( .A1(n15223), .A2(n15583), .ZN(n12538) );
  AND2_X1 U14360 ( .A1(n12539), .A2(n12538), .ZN(n15735) );
  INV_X1 U14361 ( .A(n12713), .ZN(n12540) );
  OAI22_X1 U14362 ( .A1(n15735), .A2(n16022), .B1(n12540), .B2(n15615), .ZN(
        n12543) );
  NOR2_X1 U14363 ( .A1(n12541), .A2(n16014), .ZN(n12542) );
  AOI211_X1 U14364 ( .C1(n16022), .C2(P1_REG2_REG_14__SCAN_IN), .A(n12543), 
        .B(n12542), .ZN(n12544) );
  OAI21_X1 U14365 ( .B1(n16015), .B2(n15736), .A(n12544), .ZN(n12545) );
  AOI21_X1 U14366 ( .B1(n15738), .B2(n15620), .A(n12545), .ZN(n12546) );
  OAI21_X1 U14367 ( .B1(n15622), .B2(n15740), .A(n12546), .ZN(P1_U3279) );
  MUX2_X1 U14368 ( .A(n12551), .B(n13148), .S(n13405), .Z(n12622) );
  INV_X1 U14369 ( .A(n13149), .ZN(n12553) );
  MUX2_X1 U14370 ( .A(n8429), .B(n12553), .S(n13405), .Z(n12621) );
  NOR2_X1 U14371 ( .A1(n8324), .A2(n12621), .ZN(n12554) );
  XNOR2_X1 U14372 ( .A(n12623), .B(n12554), .ZN(n12562) );
  NAND2_X1 U14373 ( .A1(n12630), .A2(n13514), .ZN(n12555) );
  OAI211_X1 U14374 ( .C1(n13384), .C2(n13470), .A(n12556), .B(n12555), .ZN(
        n12557) );
  INV_X1 U14375 ( .A(n12557), .ZN(n12559) );
  NAND2_X1 U14376 ( .A1(n14187), .A2(n13411), .ZN(n12558) );
  OAI211_X1 U14377 ( .C1(n12627), .C2(n12560), .A(n12559), .B(n12558), .ZN(
        n12561) );
  AOI21_X1 U14378 ( .B1(n12562), .B2(n13495), .A(n12561), .ZN(n12563) );
  INV_X1 U14379 ( .A(n12563), .ZN(P3_U3164) );
  INV_X1 U14380 ( .A(n12869), .ZN(n12566) );
  OAI222_X1 U14381 ( .A1(n14970), .A2(n12565), .B1(n14968), .B2(n12566), .C1(
        n12564), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U14382 ( .A1(n15773), .A2(n12870), .B1(n15771), .B2(n12566), .C1(
        n7190), .C2(n12733), .ZN(P1_U3334) );
  XNOR2_X1 U14383 ( .A(n14800), .B(n14352), .ZN(n12570) );
  AND2_X1 U14384 ( .A1(n14472), .A2(n14350), .ZN(n12569) );
  NAND2_X1 U14385 ( .A1(n12570), .A2(n12569), .ZN(n14261) );
  NAND2_X1 U14386 ( .A1(n7350), .A2(n14261), .ZN(n12571) );
  XNOR2_X1 U14387 ( .A(n14262), .B(n12571), .ZN(n12578) );
  OAI21_X1 U14388 ( .B1(n14402), .B2(n14795), .A(n12572), .ZN(n12576) );
  INV_X1 U14389 ( .A(n14799), .ZN(n12573) );
  OAI22_X1 U14390 ( .A1(n14404), .A2(n12574), .B1(n14403), .B2(n12573), .ZN(
        n12575) );
  AOI211_X1 U14391 ( .C1(n14800), .C2(n14423), .A(n12576), .B(n12575), .ZN(
        n12577) );
  OAI21_X1 U14392 ( .B1(n12578), .B2(n14449), .A(n12577), .ZN(P2_U3206) );
  INV_X1 U14393 ( .A(n12579), .ZN(n12580) );
  OAI22_X1 U14394 ( .A1(n12594), .A2(n15096), .B1(n12584), .B2(n15095), .ZN(
        n12585) );
  XNOR2_X1 U14395 ( .A(n12585), .B(n15065), .ZN(n12705) );
  AND2_X1 U14396 ( .A1(n15225), .A2(n15050), .ZN(n12586) );
  AOI21_X1 U14397 ( .B1(n12805), .B2(n11123), .A(n12586), .ZN(n12708) );
  XNOR2_X1 U14398 ( .A(n12705), .B(n12708), .ZN(n12587) );
  OAI211_X1 U14399 ( .C1(n12588), .C2(n12587), .A(n12706), .B(n15210), .ZN(
        n12593) );
  OAI22_X1 U14400 ( .A1(n12589), .A2(n15213), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12197), .ZN(n12590) );
  AOI21_X1 U14401 ( .B1(n12591), .B2(n15216), .A(n12590), .ZN(n12592) );
  OAI211_X1 U14402 ( .C1(n12594), .C2(n15220), .A(n12593), .B(n12592), .ZN(
        P1_U3234) );
  NAND2_X1 U14403 ( .A1(n12595), .A2(n12998), .ZN(n12598) );
  AOI22_X1 U14404 ( .A1(n12836), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n12835), 
        .B2(n12596), .ZN(n12597) );
  INV_X1 U14405 ( .A(n12663), .ZN(n12599) );
  AOI211_X1 U14406 ( .C1(n15729), .C2(n12600), .A(n12599), .B(n16096), .ZN(
        n15728) );
  INV_X1 U14407 ( .A(n15224), .ZN(n12601) );
  NOR2_X1 U14408 ( .A1(n15733), .A2(n12601), .ZN(n12602) );
  XNOR2_X1 U14409 ( .A(n15729), .B(n15223), .ZN(n13029) );
  XNOR2_X1 U14410 ( .A(n12659), .B(n12658), .ZN(n12613) );
  NAND2_X1 U14411 ( .A1(n15224), .A2(n15500), .ZN(n12612) );
  NAND2_X1 U14412 ( .A1(n10755), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n12610) );
  NAND2_X1 U14413 ( .A1(n12966), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12609) );
  INV_X1 U14414 ( .A(n12667), .ZN(n12669) );
  NAND2_X1 U14415 ( .A1(n12605), .A2(n15134), .ZN(n12606) );
  AND2_X1 U14416 ( .A1(n12669), .A2(n12606), .ZN(n15137) );
  NAND2_X1 U14417 ( .A1(n12965), .A2(n15137), .ZN(n12608) );
  NAND2_X1 U14418 ( .A1(n12982), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n12607) );
  NAND4_X1 U14419 ( .A1(n12610), .A2(n12609), .A3(n12608), .A4(n12607), .ZN(
        n15393) );
  NAND2_X1 U14420 ( .A1(n15393), .A2(n15437), .ZN(n12611) );
  AND2_X1 U14421 ( .A1(n12612), .A2(n12611), .ZN(n15214) );
  OAI21_X1 U14422 ( .B1(n12613), .B2(n16074), .A(n15214), .ZN(n15727) );
  AOI21_X1 U14423 ( .B1(n15728), .B2(n15343), .A(n15727), .ZN(n12620) );
  NAND2_X1 U14424 ( .A1(n15733), .A2(n15224), .ZN(n12614) );
  XNOR2_X1 U14425 ( .A(n12648), .B(n12658), .ZN(n15731) );
  INV_X1 U14426 ( .A(n15731), .ZN(n12618) );
  AOI22_X1 U14427 ( .A1(n16022), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n15217), 
        .B2(n16011), .ZN(n12616) );
  OAI21_X1 U14428 ( .B1(n8025), .B2(n16014), .A(n12616), .ZN(n12617) );
  AOI21_X1 U14429 ( .B1(n12618), .B2(n15620), .A(n12617), .ZN(n12619) );
  OAI21_X1 U14430 ( .B1(n12620), .B2(n16022), .A(n12619), .ZN(P1_U3278) );
  INV_X1 U14431 ( .A(n13275), .ZN(n12636) );
  MUX2_X1 U14432 ( .A(n12636), .B(n13275), .S(n13405), .Z(n12624) );
  OAI211_X1 U14433 ( .C1(n12625), .C2(n12624), .A(n13334), .B(n13495), .ZN(
        n12632) );
  OAI21_X1 U14434 ( .B1(n13501), .B2(n13470), .A(n12626), .ZN(n12629) );
  NOR2_X1 U14435 ( .A1(n12627), .A2(n12641), .ZN(n12628) );
  AOI211_X1 U14436 ( .C1(n12630), .C2(n13513), .A(n12629), .B(n12628), .ZN(
        n12631) );
  OAI211_X1 U14437 ( .C1(n13507), .C2(n16217), .A(n12632), .B(n12631), .ZN(
        P3_U3174) );
  OR2_X1 U14438 ( .A1(n12633), .A2(n13275), .ZN(n12634) );
  NAND2_X1 U14439 ( .A1(n12635), .A2(n12634), .ZN(n16214) );
  INV_X1 U14440 ( .A(n16214), .ZN(n12647) );
  XNOR2_X1 U14441 ( .A(n12637), .B(n12636), .ZN(n12638) );
  NAND2_X1 U14442 ( .A1(n12638), .A2(n14103), .ZN(n12640) );
  AOI22_X1 U14443 ( .A1(n14108), .A2(n13513), .B1(n14089), .B2(n14107), .ZN(
        n12639) );
  NAND2_X1 U14444 ( .A1(n12640), .A2(n12639), .ZN(n16219) );
  NAND2_X1 U14445 ( .A1(n16219), .A2(n16131), .ZN(n12646) );
  INV_X1 U14446 ( .A(n16217), .ZN(n12644) );
  OAI22_X1 U14447 ( .A1(n16131), .A2(n12642), .B1(n12641), .B2(n16128), .ZN(
        n12643) );
  AOI21_X1 U14448 ( .B1(n12644), .B2(n14065), .A(n12643), .ZN(n12645) );
  OAI211_X1 U14449 ( .C1(n14118), .C2(n12647), .A(n12646), .B(n12645), .ZN(
        P3_U3220) );
  OR2_X1 U14450 ( .A1(n15729), .A2(n15223), .ZN(n12649) );
  NAND2_X1 U14451 ( .A1(n12650), .A2(n12649), .ZN(n12655) );
  NAND2_X1 U14452 ( .A1(n12651), .A2(n12998), .ZN(n12654) );
  AOI22_X1 U14453 ( .A1(n12836), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12835), 
        .B2(n12652), .ZN(n12653) );
  XNOR2_X1 U14454 ( .A(n15719), .B(n15393), .ZN(n13031) );
  OAI21_X1 U14455 ( .B1(n12655), .B2(n12660), .A(n15395), .ZN(n12656) );
  INV_X1 U14456 ( .A(n12656), .ZN(n15726) );
  INV_X1 U14457 ( .A(n15223), .ZN(n12657) );
  INV_X1 U14458 ( .A(n12661), .ZN(n12662) );
  OAI21_X1 U14459 ( .B1(n12662), .B2(n13031), .A(n15366), .ZN(n15724) );
  INV_X1 U14460 ( .A(n15622), .ZN(n15575) );
  NAND2_X1 U14461 ( .A1(n15719), .A2(n12663), .ZN(n12664) );
  NAND2_X1 U14462 ( .A1(n7335), .A2(n12664), .ZN(n15721) );
  NOR2_X1 U14463 ( .A1(n15721), .A2(n16015), .ZN(n12680) );
  INV_X1 U14464 ( .A(n15719), .ZN(n12678) );
  INV_X1 U14465 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n12673) );
  NAND2_X1 U14466 ( .A1(n12875), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n12666) );
  NAND2_X1 U14467 ( .A1(n12966), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n12665) );
  AND2_X1 U14468 ( .A1(n12666), .A2(n12665), .ZN(n12672) );
  INV_X1 U14469 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U14470 ( .A1(n12669), .A2(n12668), .ZN(n12670) );
  NAND2_X1 U14471 ( .A1(n12829), .A2(n12670), .ZN(n15614) );
  INV_X1 U14472 ( .A(n12965), .ZN(n12858) );
  OR2_X1 U14473 ( .A1(n15614), .A2(n12858), .ZN(n12671) );
  OAI211_X1 U14474 ( .C1(n11704), .C2(n12673), .A(n12672), .B(n12671), .ZN(
        n15581) );
  NAND2_X1 U14475 ( .A1(n15581), .A2(n15583), .ZN(n12675) );
  NAND2_X1 U14476 ( .A1(n15223), .A2(n15582), .ZN(n12674) );
  AND2_X1 U14477 ( .A1(n12675), .A2(n12674), .ZN(n15135) );
  INV_X1 U14478 ( .A(n15135), .ZN(n15718) );
  AOI22_X1 U14479 ( .A1(n15718), .A2(n15611), .B1(n15137), .B2(n16011), .ZN(
        n12677) );
  NAND2_X1 U14480 ( .A1(n16022), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12676) );
  OAI211_X1 U14481 ( .C1(n12678), .C2(n16014), .A(n12677), .B(n12676), .ZN(
        n12679) );
  AOI211_X1 U14482 ( .C1(n15724), .C2(n15575), .A(n12680), .B(n12679), .ZN(
        n12681) );
  OAI21_X1 U14483 ( .B1(n15726), .B2(n15577), .A(n12681), .ZN(P1_U3277) );
  OAI222_X1 U14484 ( .A1(n14970), .A2(n12684), .B1(P2_U3088), .B2(n12683), 
        .C1(n14968), .C2(n12682), .ZN(P2_U3305) );
  INV_X1 U14485 ( .A(n12685), .ZN(n12687) );
  INV_X1 U14486 ( .A(n12907), .ZN(n12689) );
  OAI222_X1 U14487 ( .A1(P1_U3086), .A2(n12687), .B1(n15771), .B2(n12689), 
        .C1(n15773), .C2(n12686), .ZN(P1_U3331) );
  INV_X1 U14488 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12690) );
  OAI222_X1 U14489 ( .A1(n14970), .A2(n12690), .B1(n14968), .B2(n12689), .C1(
        P2_U3088), .C2(n12688), .ZN(P2_U3303) );
  NAND2_X1 U14490 ( .A1(n12823), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n12692) );
  NAND2_X1 U14491 ( .A1(n12692), .A2(n12691), .ZN(n15332) );
  XNOR2_X1 U14492 ( .A(n15332), .B(n12699), .ZN(n15333) );
  XNOR2_X1 U14493 ( .A(n15333), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n12703) );
  AOI21_X1 U14494 ( .B1(n12823), .B2(P1_REG1_REG_17__SCAN_IN), .A(n12693), 
        .ZN(n12694) );
  NOR2_X1 U14495 ( .A1(n12694), .A2(n12699), .ZN(n15329) );
  INV_X1 U14496 ( .A(n15330), .ZN(n12695) );
  OAI211_X1 U14497 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n12696), .A(n12695), 
        .B(n15927), .ZN(n12702) );
  INV_X1 U14498 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n15190) );
  NOR2_X1 U14499 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15190), .ZN(n12697) );
  AOI21_X1 U14500 ( .B1(n15914), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n12697), 
        .ZN(n12698) );
  OAI21_X1 U14501 ( .B1(n15337), .B2(n12699), .A(n12698), .ZN(n12700) );
  INV_X1 U14502 ( .A(n12700), .ZN(n12701) );
  OAI211_X1 U14503 ( .C1(n12703), .C2(n15338), .A(n12702), .B(n12701), .ZN(
        P1_U3261) );
  AOI22_X1 U14504 ( .A1(n15733), .A2(n15062), .B1(n11123), .B2(n15224), .ZN(
        n12704) );
  XNOR2_X1 U14505 ( .A(n12704), .B(n15065), .ZN(n14981) );
  AOI22_X1 U14506 ( .A1(n15733), .A2(n11123), .B1(n15050), .B2(n15224), .ZN(
        n14982) );
  XNOR2_X1 U14507 ( .A(n14981), .B(n14982), .ZN(n12710) );
  INV_X1 U14508 ( .A(n12705), .ZN(n12707) );
  OAI21_X1 U14509 ( .B1(n12708), .B2(n12707), .A(n12706), .ZN(n12709) );
  AOI21_X1 U14510 ( .B1(n12710), .B2(n12709), .A(n14980), .ZN(n12716) );
  OAI22_X1 U14511 ( .A1(n15735), .A2(n15213), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12711), .ZN(n12712) );
  AOI21_X1 U14512 ( .B1(n12713), .B2(n15216), .A(n12712), .ZN(n12715) );
  NAND2_X1 U14513 ( .A1(n15733), .A2(n15196), .ZN(n12714) );
  OAI211_X1 U14514 ( .C1(n12716), .C2(n15205), .A(n12715), .B(n12714), .ZN(
        P1_U3215) );
  INV_X1 U14515 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12717) );
  OAI222_X1 U14516 ( .A1(n14975), .A2(n13079), .B1(P2_U3088), .B2(n12718), 
        .C1(n12717), .C2(n14970), .ZN(P2_U3297) );
  INV_X1 U14517 ( .A(n12940), .ZN(n13322) );
  OAI222_X1 U14518 ( .A1(n15773), .A2(n12941), .B1(n15771), .B2(n13322), .C1(
        n7190), .C2(n15351), .ZN(P1_U3328) );
  OAI222_X1 U14519 ( .A1(n14970), .A2(n12720), .B1(n14968), .B2(n12719), .C1(
        n10115), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U14520 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n12726) );
  INV_X1 U14521 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n12721) );
  INV_X1 U14522 ( .A(n12851), .ZN(n12723) );
  NAND2_X1 U14523 ( .A1(n12831), .A2(n12721), .ZN(n12722) );
  NAND2_X1 U14524 ( .A1(n12723), .A2(n12722), .ZN(n15569) );
  OR2_X1 U14525 ( .A1(n15569), .A2(n12858), .ZN(n12725) );
  AOI22_X1 U14526 ( .A1(n12966), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n12875), 
        .B2(P1_REG1_REG_19__SCAN_IN), .ZN(n12724) );
  OAI211_X1 U14527 ( .C1(n11704), .C2(n12726), .A(n12725), .B(n12724), .ZN(
        n15584) );
  NAND2_X1 U14528 ( .A1(n12727), .A2(n12998), .ZN(n12729) );
  AOI22_X1 U14529 ( .A1(n12836), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n12730), 
        .B2(n12835), .ZN(n12728) );
  INV_X1 U14530 ( .A(n12734), .ZN(n12732) );
  MUX2_X1 U14531 ( .A(n15584), .B(n15698), .S(n13004), .Z(n12846) );
  MUX2_X1 U14532 ( .A(n15729), .B(n15223), .S(n13051), .Z(n12814) );
  NAND2_X1 U14533 ( .A1(n12736), .A2(n13004), .ZN(n12738) );
  NAND2_X1 U14534 ( .A1(n12738), .A2(n12737), .ZN(n12739) );
  INV_X1 U14535 ( .A(n12741), .ZN(n15238) );
  NAND2_X1 U14536 ( .A1(n15238), .A2(n16013), .ZN(n13009) );
  NAND2_X1 U14537 ( .A1(n13009), .A2(n12742), .ZN(n12743) );
  NAND4_X1 U14538 ( .A1(n13010), .A2(n12744), .A3(n13004), .A4(n12743), .ZN(
        n12748) );
  NAND3_X1 U14539 ( .A1(n12746), .A2(n12745), .A3(n13051), .ZN(n12747) );
  OAI21_X1 U14540 ( .B1(n15236), .B2(n13051), .A(n15181), .ZN(n12752) );
  NAND2_X1 U14541 ( .A1(n15236), .A2(n13051), .ZN(n12750) );
  NAND2_X1 U14542 ( .A1(n12750), .A2(n12749), .ZN(n12751) );
  NAND2_X1 U14543 ( .A1(n12752), .A2(n12751), .ZN(n12753) );
  OAI21_X1 U14544 ( .B1(n15235), .B2(n13004), .A(n12757), .ZN(n12760) );
  NAND2_X1 U14545 ( .A1(n15235), .A2(n13004), .ZN(n12758) );
  NAND2_X1 U14546 ( .A1(n12758), .A2(n8021), .ZN(n12759) );
  NAND2_X1 U14547 ( .A1(n12760), .A2(n12759), .ZN(n12761) );
  OAI21_X1 U14548 ( .B1(n15234), .B2(n13051), .A(n12762), .ZN(n12765) );
  NAND2_X1 U14549 ( .A1(n15234), .A2(n13051), .ZN(n12763) );
  NAND2_X1 U14550 ( .A1(n12763), .A2(n16070), .ZN(n12764) );
  NAND2_X1 U14551 ( .A1(n12765), .A2(n12764), .ZN(n12766) );
  NAND3_X1 U14552 ( .A1(n12768), .A2(n12767), .A3(n12766), .ZN(n12773) );
  AND2_X1 U14553 ( .A1(n15233), .A2(n13004), .ZN(n12771) );
  OAI21_X1 U14554 ( .B1(n13004), .B2(n15233), .A(n12770), .ZN(n12769) );
  OAI21_X1 U14555 ( .B1(n12771), .B2(n12770), .A(n12769), .ZN(n12772) );
  MUX2_X1 U14556 ( .A(n15232), .B(n12774), .S(n13051), .Z(n12776) );
  MUX2_X1 U14557 ( .A(n15232), .B(n12774), .S(n13004), .Z(n12775) );
  INV_X1 U14558 ( .A(n12776), .ZN(n12777) );
  MUX2_X1 U14559 ( .A(n15231), .B(n16111), .S(n13004), .Z(n12779) );
  MUX2_X1 U14560 ( .A(n15231), .B(n16111), .S(n13051), .Z(n12778) );
  MUX2_X1 U14561 ( .A(n15230), .B(n12780), .S(n13051), .Z(n12783) );
  MUX2_X1 U14562 ( .A(n15230), .B(n12780), .S(n13004), .Z(n12781) );
  INV_X1 U14563 ( .A(n12783), .ZN(n12784) );
  MUX2_X1 U14564 ( .A(n16152), .B(n15229), .S(n13051), .Z(n12788) );
  MUX2_X1 U14565 ( .A(n16152), .B(n15229), .S(n13004), .Z(n12785) );
  NAND2_X1 U14566 ( .A1(n12786), .A2(n12785), .ZN(n12792) );
  INV_X1 U14567 ( .A(n12787), .ZN(n12790) );
  INV_X1 U14568 ( .A(n12788), .ZN(n12789) );
  NAND2_X1 U14569 ( .A1(n12790), .A2(n12789), .ZN(n12791) );
  MUX2_X1 U14570 ( .A(n15228), .B(n12793), .S(n13051), .Z(n12795) );
  MUX2_X1 U14571 ( .A(n12793), .B(n15228), .S(n13051), .Z(n12794) );
  MUX2_X1 U14572 ( .A(n15227), .B(n12797), .S(n13004), .Z(n12799) );
  MUX2_X1 U14573 ( .A(n15227), .B(n12797), .S(n13051), .Z(n12798) );
  AND2_X1 U14574 ( .A1(n15226), .A2(n13051), .ZN(n12802) );
  OAI21_X1 U14575 ( .B1(n15226), .B2(n13051), .A(n12801), .ZN(n12800) );
  OAI21_X1 U14576 ( .B1(n12802), .B2(n12801), .A(n12800), .ZN(n12803) );
  MUX2_X1 U14577 ( .A(n15225), .B(n12805), .S(n13004), .Z(n12808) );
  MUX2_X1 U14578 ( .A(n15225), .B(n12805), .S(n13051), .Z(n12806) );
  INV_X1 U14579 ( .A(n12808), .ZN(n12809) );
  MUX2_X1 U14580 ( .A(n15224), .B(n15733), .S(n13051), .Z(n12811) );
  MUX2_X1 U14581 ( .A(n15224), .B(n15733), .S(n13004), .Z(n12810) );
  INV_X1 U14582 ( .A(n12811), .ZN(n12812) );
  MUX2_X1 U14583 ( .A(n15729), .B(n15223), .S(n13004), .Z(n12813) );
  MUX2_X1 U14584 ( .A(n15719), .B(n15393), .S(n13004), .Z(n12817) );
  NAND2_X1 U14585 ( .A1(n12818), .A2(n12817), .ZN(n12816) );
  MUX2_X1 U14586 ( .A(n15719), .B(n15393), .S(n13051), .Z(n12815) );
  NAND2_X1 U14587 ( .A1(n12816), .A2(n12815), .ZN(n12821) );
  INV_X1 U14588 ( .A(n12817), .ZN(n12820) );
  INV_X1 U14589 ( .A(n12818), .ZN(n12819) );
  NAND2_X1 U14590 ( .A1(n12822), .A2(n12998), .ZN(n12825) );
  AOI22_X1 U14591 ( .A1(n12836), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12835), 
        .B2(n12823), .ZN(n12824) );
  MUX2_X1 U14592 ( .A(n15581), .B(n15711), .S(n13004), .Z(n12827) );
  MUX2_X1 U14593 ( .A(n15581), .B(n15711), .S(n13051), .Z(n12826) );
  INV_X1 U14594 ( .A(n12827), .ZN(n12828) );
  NAND2_X1 U14595 ( .A1(n12829), .A2(n15190), .ZN(n12830) );
  NAND2_X1 U14596 ( .A1(n12831), .A2(n12830), .ZN(n15594) );
  AOI22_X1 U14597 ( .A1(n12966), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n12982), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n12833) );
  NAND2_X1 U14598 ( .A1(n12875), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n12832) );
  OAI211_X1 U14599 ( .C1(n15594), .C2(n12858), .A(n12833), .B(n12832), .ZN(
        n15369) );
  AOI22_X1 U14600 ( .A1(n12836), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n12835), 
        .B2(n15331), .ZN(n12837) );
  MUX2_X1 U14601 ( .A(n15369), .B(n15705), .S(n13051), .Z(n12841) );
  MUX2_X1 U14602 ( .A(n15705), .B(n15369), .S(n13051), .Z(n12839) );
  MUX2_X1 U14603 ( .A(n15584), .B(n15698), .S(n13051), .Z(n12843) );
  NAND2_X1 U14604 ( .A1(n12847), .A2(n12998), .ZN(n12850) );
  OR2_X1 U14605 ( .A1(n13000), .A2(n12848), .ZN(n12849) );
  NOR2_X1 U14606 ( .A1(n12851), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n12852) );
  OR2_X1 U14607 ( .A1(n12861), .A2(n12852), .ZN(n15555) );
  INV_X1 U14608 ( .A(n12966), .ZN(n12985) );
  INV_X1 U14609 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n12855) );
  NAND2_X1 U14610 ( .A1(n12875), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n12854) );
  NAND2_X1 U14611 ( .A1(n12982), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n12853) );
  OAI211_X1 U14612 ( .C1(n12985), .C2(n12855), .A(n12854), .B(n12853), .ZN(
        n12856) );
  INV_X1 U14613 ( .A(n12856), .ZN(n12857) );
  OAI21_X1 U14614 ( .B1(n15555), .B2(n12858), .A(n12857), .ZN(n15400) );
  MUX2_X1 U14615 ( .A(n15688), .B(n15400), .S(n13004), .Z(n12860) );
  MUX2_X1 U14616 ( .A(n15688), .B(n15400), .S(n13051), .Z(n12859) );
  OR2_X1 U14617 ( .A1(n12861), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12862) );
  AND2_X1 U14618 ( .A1(n12862), .A2(n12877), .ZN(n15540) );
  NAND2_X1 U14619 ( .A1(n15540), .A2(n12965), .ZN(n12868) );
  INV_X1 U14620 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n12865) );
  NAND2_X1 U14621 ( .A1(n12875), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n12864) );
  NAND2_X1 U14622 ( .A1(n12982), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n12863) );
  OAI211_X1 U14623 ( .C1(n12985), .C2(n12865), .A(n12864), .B(n12863), .ZN(
        n12866) );
  INV_X1 U14624 ( .A(n12866), .ZN(n12867) );
  NAND2_X1 U14625 ( .A1(n12868), .A2(n12867), .ZN(n15402) );
  NAND2_X1 U14626 ( .A1(n12869), .A2(n12998), .ZN(n12872) );
  OR2_X1 U14627 ( .A1(n13000), .A2(n12870), .ZN(n12871) );
  MUX2_X1 U14628 ( .A(n15402), .B(n15679), .S(n13004), .Z(n12873) );
  MUX2_X1 U14629 ( .A(n15402), .B(n15679), .S(n13051), .Z(n12874) );
  NAND2_X1 U14630 ( .A1(n12875), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12881) );
  NAND2_X1 U14631 ( .A1(n12966), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n12880) );
  INV_X1 U14632 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15173) );
  INV_X1 U14633 ( .A(n12877), .ZN(n12876) );
  NAND2_X1 U14634 ( .A1(n12876), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12889) );
  AOI21_X1 U14635 ( .B1(n15173), .B2(n12877), .A(n12888), .ZN(n15526) );
  NAND2_X1 U14636 ( .A1(n12965), .A2(n15526), .ZN(n12879) );
  NAND2_X1 U14637 ( .A1(n12982), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n12878) );
  NAND4_X1 U14638 ( .A1(n12881), .A2(n12880), .A3(n12879), .A4(n12878), .ZN(
        n15501) );
  NAND2_X1 U14639 ( .A1(n12882), .A2(n7560), .ZN(n12883) );
  MUX2_X1 U14640 ( .A(n15501), .B(n15672), .S(n13051), .Z(n12886) );
  MUX2_X1 U14641 ( .A(n15501), .B(n15672), .S(n13004), .Z(n12884) );
  INV_X1 U14642 ( .A(n12886), .ZN(n12887) );
  NAND2_X1 U14643 ( .A1(n10755), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U14644 ( .A1(n12966), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n12892) );
  INV_X1 U14645 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n15075) );
  AOI21_X1 U14646 ( .B1(n15075), .B2(n12889), .A(n12901), .ZN(n15506) );
  NAND2_X1 U14647 ( .A1(n12965), .A2(n15506), .ZN(n12891) );
  NAND2_X1 U14648 ( .A1(n12982), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n12890) );
  NAND4_X1 U14649 ( .A1(n12893), .A2(n12892), .A3(n12891), .A4(n12890), .ZN(
        n15406) );
  INV_X1 U14650 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12894) );
  OR2_X1 U14651 ( .A1(n13000), .A2(n12894), .ZN(n12895) );
  MUX2_X1 U14652 ( .A(n15406), .B(n15667), .S(n13004), .Z(n12898) );
  MUX2_X1 U14653 ( .A(n15406), .B(n15667), .S(n13051), .Z(n12896) );
  NAND2_X1 U14654 ( .A1(n12897), .A2(n12896), .ZN(n12900) );
  NAND2_X1 U14655 ( .A1(n7292), .A2(n7501), .ZN(n12899) );
  NAND2_X1 U14656 ( .A1(n12875), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12906) );
  NAND2_X1 U14657 ( .A1(n12966), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12905) );
  INV_X1 U14658 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n15151) );
  NAND2_X1 U14659 ( .A1(n12901), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12913) );
  AOI21_X1 U14660 ( .B1(n15151), .B2(n12902), .A(n12912), .ZN(n15492) );
  NAND2_X1 U14661 ( .A1(n12965), .A2(n15492), .ZN(n12904) );
  NAND2_X1 U14662 ( .A1(n12982), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n12903) );
  NAND4_X1 U14663 ( .A1(n12906), .A2(n12905), .A3(n12904), .A4(n12903), .ZN(
        n15502) );
  NAND2_X1 U14664 ( .A1(n12907), .A2(n12998), .ZN(n12909) );
  OR2_X1 U14665 ( .A1(n13000), .A2(n12686), .ZN(n12908) );
  MUX2_X1 U14666 ( .A(n15502), .B(n15662), .S(n13051), .Z(n12911) );
  MUX2_X1 U14667 ( .A(n15502), .B(n15662), .S(n13004), .Z(n12910) );
  NAND2_X1 U14668 ( .A1(n12875), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12917) );
  NAND2_X1 U14669 ( .A1(n12966), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12916) );
  INV_X1 U14670 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n15127) );
  NAND2_X1 U14671 ( .A1(n12912), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n12924) );
  INV_X1 U14672 ( .A(n12924), .ZN(n12923) );
  AOI21_X1 U14673 ( .B1(n15127), .B2(n12913), .A(n12923), .ZN(n15473) );
  NAND2_X1 U14674 ( .A1(n12965), .A2(n15473), .ZN(n12915) );
  NAND2_X1 U14675 ( .A1(n12982), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n12914) );
  NAND4_X1 U14676 ( .A1(n12917), .A2(n12916), .A3(n12915), .A4(n12914), .ZN(
        n15378) );
  NAND2_X1 U14677 ( .A1(n14966), .A2(n12998), .ZN(n12919) );
  OR2_X1 U14678 ( .A1(n13000), .A2(n15772), .ZN(n12918) );
  MUX2_X1 U14679 ( .A(n15378), .B(n15654), .S(n13004), .Z(n12921) );
  MUX2_X1 U14680 ( .A(n15378), .B(n15654), .S(n13051), .Z(n12920) );
  INV_X1 U14681 ( .A(n12921), .ZN(n12922) );
  NAND2_X1 U14682 ( .A1(n12875), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12928) );
  NAND2_X1 U14683 ( .A1(n12966), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n12927) );
  INV_X1 U14684 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n15201) );
  NAND2_X1 U14685 ( .A1(n12923), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12935) );
  INV_X1 U14686 ( .A(n12935), .ZN(n12934) );
  AOI21_X1 U14687 ( .B1(n15201), .B2(n12924), .A(n12934), .ZN(n15458) );
  NAND2_X1 U14688 ( .A1(n12965), .A2(n15458), .ZN(n12926) );
  NAND2_X1 U14689 ( .A1(n12982), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n12925) );
  NAND4_X1 U14690 ( .A1(n12928), .A2(n12927), .A3(n12926), .A4(n12925), .ZN(
        n15439) );
  NAND2_X1 U14691 ( .A1(n14963), .A2(n12998), .ZN(n12930) );
  OR2_X1 U14692 ( .A1(n13000), .A2(n15766), .ZN(n12929) );
  MUX2_X1 U14693 ( .A(n15439), .B(n15459), .S(n13051), .Z(n12933) );
  MUX2_X1 U14694 ( .A(n15439), .B(n15459), .S(n13004), .Z(n12931) );
  NAND2_X1 U14695 ( .A1(n12966), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n12939) );
  NAND2_X1 U14696 ( .A1(n12875), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n12938) );
  INV_X1 U14697 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n15068) );
  NAND2_X1 U14698 ( .A1(n12934), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n12949) );
  INV_X1 U14699 ( .A(n12949), .ZN(n12948) );
  AOI21_X1 U14700 ( .B1(n15068), .B2(n12935), .A(n12948), .ZN(n15445) );
  NAND2_X1 U14701 ( .A1(n12965), .A2(n15445), .ZN(n12937) );
  NAND2_X1 U14702 ( .A1(n12982), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n12936) );
  NAND4_X1 U14703 ( .A1(n12939), .A2(n12938), .A3(n12937), .A4(n12936), .ZN(
        n15222) );
  NAND2_X1 U14704 ( .A1(n12940), .A2(n12998), .ZN(n12943) );
  OR2_X1 U14705 ( .A1(n13000), .A2(n12941), .ZN(n12942) );
  MUX2_X1 U14706 ( .A(n15222), .B(n15643), .S(n13004), .Z(n12945) );
  MUX2_X1 U14707 ( .A(n15222), .B(n15643), .S(n13051), .Z(n12944) );
  NAND2_X1 U14708 ( .A1(n13080), .A2(n12998), .ZN(n12947) );
  OR2_X1 U14709 ( .A1(n13000), .A2(n13081), .ZN(n12946) );
  NAND2_X1 U14710 ( .A1(n10755), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12953) );
  NAND2_X1 U14711 ( .A1(n12966), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12952) );
  INV_X1 U14712 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n15101) );
  NAND2_X1 U14713 ( .A1(n12948), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n15386) );
  INV_X1 U14714 ( .A(n15386), .ZN(n12964) );
  AOI21_X1 U14715 ( .B1(n15101), .B2(n12949), .A(n12964), .ZN(n15425) );
  NAND2_X1 U14716 ( .A1(n12965), .A2(n15425), .ZN(n12951) );
  NAND2_X1 U14717 ( .A1(n12982), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n12950) );
  NAND4_X1 U14718 ( .A1(n12953), .A2(n12952), .A3(n12951), .A4(n12950), .ZN(
        n15438) );
  MUX2_X1 U14719 ( .A(n15636), .B(n15438), .S(n13004), .Z(n12957) );
  NAND2_X1 U14720 ( .A1(n12956), .A2(n12957), .ZN(n12955) );
  MUX2_X1 U14721 ( .A(n15636), .B(n15438), .S(n13051), .Z(n12954) );
  NAND2_X1 U14722 ( .A1(n12955), .A2(n12954), .ZN(n12961) );
  INV_X1 U14723 ( .A(n12956), .ZN(n12959) );
  INV_X1 U14724 ( .A(n12957), .ZN(n12958) );
  NAND2_X1 U14725 ( .A1(n12959), .A2(n12958), .ZN(n12960) );
  NAND2_X1 U14726 ( .A1(n12961), .A2(n12960), .ZN(n12973) );
  NAND2_X1 U14727 ( .A1(n14958), .A2(n12998), .ZN(n12963) );
  OR2_X1 U14728 ( .A1(n13000), .A2(n15765), .ZN(n12962) );
  NAND2_X1 U14729 ( .A1(n12965), .A2(n12964), .ZN(n12970) );
  NAND2_X1 U14730 ( .A1(n12966), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12969) );
  NAND2_X1 U14731 ( .A1(n12982), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12968) );
  NAND2_X1 U14732 ( .A1(n12875), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12967) );
  NAND4_X1 U14733 ( .A1(n12970), .A2(n12969), .A3(n12968), .A4(n12967), .ZN(
        n15221) );
  MUX2_X1 U14734 ( .A(n15634), .B(n15221), .S(n13051), .Z(n12974) );
  INV_X1 U14735 ( .A(n15221), .ZN(n12971) );
  INV_X1 U14736 ( .A(n15634), .ZN(n15391) );
  MUX2_X1 U14737 ( .A(n12971), .B(n15391), .S(n13051), .Z(n12972) );
  INV_X1 U14738 ( .A(n12973), .ZN(n12976) );
  INV_X1 U14739 ( .A(n12974), .ZN(n12975) );
  AOI22_X1 U14740 ( .A1(n12978), .A2(n12977), .B1(n12976), .B2(n12975), .ZN(
        n13077) );
  INV_X1 U14741 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n12981) );
  NAND2_X1 U14742 ( .A1(n10755), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12980) );
  NAND2_X1 U14743 ( .A1(n12982), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12979) );
  OAI211_X1 U14744 ( .C1(n12985), .C2(n12981), .A(n12980), .B(n12979), .ZN(
        n15353) );
  INV_X1 U14745 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n15358) );
  NAND2_X1 U14746 ( .A1(n12875), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12984) );
  NAND2_X1 U14747 ( .A1(n12982), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12983) );
  OAI211_X1 U14748 ( .C1(n12985), .C2(n15358), .A(n12984), .B(n12983), .ZN(
        n15385) );
  OAI21_X1 U14749 ( .B1(n15353), .B2(n12992), .A(n15385), .ZN(n12986) );
  INV_X1 U14750 ( .A(n12986), .ZN(n12990) );
  OR2_X1 U14751 ( .A1(n13079), .A2(n12987), .ZN(n12989) );
  INV_X1 U14752 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13235) );
  OR2_X1 U14753 ( .A1(n13000), .A2(n13235), .ZN(n12988) );
  MUX2_X1 U14754 ( .A(n12990), .B(n15361), .S(n13051), .Z(n13057) );
  INV_X1 U14755 ( .A(n13057), .ZN(n13065) );
  NAND2_X1 U14756 ( .A1(n12992), .A2(n12991), .ZN(n12993) );
  NAND2_X1 U14757 ( .A1(n12994), .A2(n12993), .ZN(n12995) );
  AND2_X1 U14758 ( .A1(n12996), .A2(n12995), .ZN(n13043) );
  INV_X1 U14759 ( .A(n13043), .ZN(n13054) );
  AND2_X1 U14760 ( .A1(n13054), .A2(n13044), .ZN(n13072) );
  INV_X1 U14761 ( .A(n13072), .ZN(n12997) );
  NOR3_X1 U14762 ( .A1(n13065), .A2(n15775), .A3(n12997), .ZN(n13059) );
  NAND2_X1 U14763 ( .A1(n15758), .A2(n12998), .ZN(n13002) );
  INV_X1 U14764 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12999) );
  OR2_X1 U14765 ( .A1(n13000), .A2(n12999), .ZN(n13001) );
  INV_X1 U14766 ( .A(n15353), .ZN(n13003) );
  NAND2_X1 U14767 ( .A1(n15354), .A2(n13003), .ZN(n13006) );
  OR2_X1 U14768 ( .A1(n15354), .A2(n13003), .ZN(n13005) );
  MUX2_X1 U14769 ( .A(n13006), .B(n13005), .S(n13004), .Z(n13060) );
  XNOR2_X1 U14770 ( .A(n15354), .B(n15353), .ZN(n13071) );
  NAND2_X1 U14771 ( .A1(n15427), .A2(n15381), .ZN(n13007) );
  NAND2_X1 U14772 ( .A1(n15636), .A2(n15438), .ZN(n15411) );
  NAND2_X1 U14773 ( .A1(n13007), .A2(n15411), .ZN(n15420) );
  NAND2_X1 U14774 ( .A1(n15654), .A2(n15378), .ZN(n15407) );
  OR2_X1 U14775 ( .A1(n15654), .A2(n15378), .ZN(n13008) );
  NAND2_X1 U14776 ( .A1(n15407), .A2(n13008), .ZN(n15469) );
  INV_X1 U14777 ( .A(n15501), .ZN(n15376) );
  INV_X1 U14778 ( .A(n15402), .ZN(n15374) );
  XNOR2_X1 U14779 ( .A(n15679), .B(n15374), .ZN(n15404) );
  XNOR2_X1 U14780 ( .A(n15688), .B(n15400), .ZN(n15549) );
  INV_X1 U14781 ( .A(n15581), .ZN(n15367) );
  XNOR2_X1 U14782 ( .A(n15711), .B(n15367), .ZN(n15603) );
  AND2_X1 U14783 ( .A1(n13010), .A2(n13009), .ZN(n16012) );
  NAND4_X1 U14784 ( .A1(n16012), .A2(n10778), .A3(n13012), .A4(n13011), .ZN(
        n13015) );
  NOR3_X1 U14785 ( .A1(n13015), .A2(n13014), .A3(n13013), .ZN(n13018) );
  NAND4_X1 U14786 ( .A1(n13019), .A2(n13018), .A3(n13017), .A4(n13016), .ZN(
        n13020) );
  NOR2_X1 U14787 ( .A1(n13021), .A2(n13020), .ZN(n13024) );
  NAND4_X1 U14788 ( .A1(n13025), .A2(n13024), .A3(n13023), .A4(n13022), .ZN(
        n13026) );
  NOR2_X1 U14789 ( .A1(n13027), .A2(n13026), .ZN(n13030) );
  NAND4_X1 U14790 ( .A1(n13031), .A2(n13030), .A3(n13029), .A4(n13028), .ZN(
        n13032) );
  NOR2_X1 U14791 ( .A1(n15603), .A2(n13032), .ZN(n13033) );
  XNOR2_X1 U14792 ( .A(n15698), .B(n15584), .ZN(n15565) );
  NAND4_X1 U14793 ( .A1(n15549), .A2(n13033), .A3(n15565), .A4(n15586), .ZN(
        n13034) );
  NOR2_X1 U14794 ( .A1(n15404), .A2(n13034), .ZN(n13035) );
  XNOR2_X1 U14795 ( .A(n15662), .B(n15502), .ZN(n15377) );
  AND4_X1 U14796 ( .A1(n15469), .A2(n15522), .A3(n13035), .A4(n15377), .ZN(
        n13036) );
  XNOR2_X1 U14797 ( .A(n15459), .B(n15439), .ZN(n15455) );
  NAND4_X1 U14798 ( .A1(n15420), .A2(n13036), .A3(n15455), .A4(n15509), .ZN(
        n13037) );
  XNOR2_X1 U14799 ( .A(n15643), .B(n15410), .ZN(n15380) );
  NOR2_X1 U14800 ( .A1(n13037), .A2(n15380), .ZN(n13039) );
  XNOR2_X1 U14801 ( .A(n15634), .B(n15221), .ZN(n15412) );
  XNOR2_X1 U14802 ( .A(n15361), .B(n15385), .ZN(n13038) );
  NAND4_X1 U14803 ( .A1(n13071), .A2(n13039), .A3(n15412), .A4(n13038), .ZN(
        n13040) );
  XNOR2_X1 U14804 ( .A(n13040), .B(n15343), .ZN(n13042) );
  NAND2_X1 U14805 ( .A1(n13042), .A2(n13041), .ZN(n13047) );
  XNOR2_X1 U14806 ( .A(n13060), .B(n13043), .ZN(n13045) );
  NAND2_X1 U14807 ( .A1(n13045), .A2(n13044), .ZN(n13046) );
  NAND2_X1 U14808 ( .A1(n13047), .A2(n13046), .ZN(n13070) );
  INV_X1 U14809 ( .A(n13048), .ZN(n13049) );
  OAI21_X1 U14810 ( .B1(n15353), .B2(n13049), .A(n15385), .ZN(n13050) );
  INV_X1 U14811 ( .A(n13050), .ZN(n13052) );
  MUX2_X1 U14812 ( .A(n15361), .B(n13052), .S(n13051), .Z(n13064) );
  NOR3_X1 U14813 ( .A1(n13070), .A2(n13064), .A3(n15775), .ZN(n13053) );
  AOI21_X1 U14814 ( .B1(n13059), .B2(n13060), .A(n13053), .ZN(n13076) );
  INV_X1 U14815 ( .A(n13064), .ZN(n13058) );
  NOR2_X1 U14816 ( .A1(n13054), .A2(n15775), .ZN(n13063) );
  INV_X1 U14817 ( .A(n13063), .ZN(n13056) );
  INV_X1 U14818 ( .A(n13071), .ZN(n13055) );
  AOI211_X1 U14819 ( .C1(n13057), .C2(n13058), .A(n13056), .B(n13055), .ZN(
        n13075) );
  NAND2_X1 U14820 ( .A1(n13059), .A2(n13058), .ZN(n13069) );
  INV_X1 U14821 ( .A(n13060), .ZN(n13068) );
  NAND3_X1 U14822 ( .A1(n13061), .A2(n15905), .A3(n15582), .ZN(n13062) );
  OAI211_X1 U14823 ( .C1(n15779), .C2(n15775), .A(n13062), .B(P1_B_REG_SCAN_IN), .ZN(n13067) );
  NAND4_X1 U14824 ( .A1(n13071), .A2(n13065), .A3(n13064), .A4(n13063), .ZN(
        n13066) );
  OAI211_X1 U14825 ( .C1(n13069), .C2(n13068), .A(n13067), .B(n13066), .ZN(
        n13074) );
  AOI211_X1 U14826 ( .C1(n13072), .C2(n13071), .A(n15775), .B(n13070), .ZN(
        n13073) );
  OAI222_X1 U14827 ( .A1(n15771), .A2(n13079), .B1(P1_U3086), .B2(n13078), 
        .C1(n13235), .C2(n15773), .ZN(P1_U3325) );
  INV_X1 U14828 ( .A(n13080), .ZN(n14962) );
  OAI222_X1 U14829 ( .A1(n15773), .A2(n13081), .B1(n15771), .B2(n14962), .C1(
        P1_U3086), .C2(n10290), .ZN(P1_U3327) );
  NAND2_X1 U14830 ( .A1(n13082), .A2(n14805), .ZN(n13091) );
  OAI22_X1 U14831 ( .A1(n13084), .A2(n14697), .B1(n13083), .B2(n14805), .ZN(
        n13085) );
  AOI21_X1 U14832 ( .B1(n13086), .B2(n14747), .A(n13085), .ZN(n13087) );
  OAI21_X1 U14833 ( .B1(n13088), .B2(n14751), .A(n13087), .ZN(n13089) );
  INV_X1 U14834 ( .A(n13089), .ZN(n13090) );
  OAI211_X1 U14835 ( .C1(n13092), .C2(n16062), .A(n13091), .B(n13090), .ZN(
        P2_U3236) );
  MUX2_X1 U14836 ( .A(n14088), .B(n14179), .S(n13217), .Z(n13169) );
  AND2_X1 U14837 ( .A1(n13096), .A2(n13095), .ZN(n13101) );
  INV_X1 U14838 ( .A(n13101), .ZN(n13097) );
  NAND3_X1 U14839 ( .A1(n7707), .A2(n13098), .A3(n13097), .ZN(n13099) );
  OAI211_X1 U14840 ( .C1(n13100), .C2(n8055), .A(n13099), .B(n13108), .ZN(
        n13106) );
  INV_X1 U14841 ( .A(n11635), .ZN(n13104) );
  NAND3_X1 U14842 ( .A1(n7707), .A2(n13102), .A3(n13101), .ZN(n13103) );
  NAND3_X1 U14843 ( .A1(n13104), .A2(n13107), .A3(n13103), .ZN(n13105) );
  MUX2_X1 U14844 ( .A(n13106), .B(n13105), .S(n13217), .Z(n13110) );
  MUX2_X1 U14845 ( .A(n13108), .B(n13107), .S(n13229), .Z(n13109) );
  NAND4_X1 U14846 ( .A1(n13265), .A2(n13113), .A3(n13110), .A4(n13109), .ZN(
        n13120) );
  MUX2_X1 U14847 ( .A(n13521), .B(n13217), .S(n13111), .Z(n13112) );
  AOI21_X1 U14848 ( .B1(n13229), .B2(n7730), .A(n13112), .ZN(n13117) );
  INV_X1 U14849 ( .A(n13113), .ZN(n13261) );
  MUX2_X1 U14850 ( .A(n13115), .B(n13114), .S(n13229), .Z(n13116) );
  OAI21_X1 U14851 ( .B1(n13117), .B2(n13261), .A(n13116), .ZN(n13118) );
  NAND3_X1 U14852 ( .A1(n13120), .A2(n13119), .A3(n13118), .ZN(n13125) );
  MUX2_X1 U14853 ( .A(n13122), .B(n13121), .S(n13229), .Z(n13123) );
  NAND3_X1 U14854 ( .A1(n13125), .A2(n13124), .A3(n13123), .ZN(n13129) );
  MUX2_X1 U14855 ( .A(n13127), .B(n13126), .S(n13217), .Z(n13128) );
  NAND3_X1 U14856 ( .A1(n13129), .A2(n13257), .A3(n13128), .ZN(n13135) );
  INV_X1 U14857 ( .A(n13264), .ZN(n13134) );
  NAND2_X1 U14858 ( .A1(n13130), .A2(n13229), .ZN(n13132) );
  NAND2_X1 U14859 ( .A1(n16125), .A2(n13217), .ZN(n13131) );
  MUX2_X1 U14860 ( .A(n13132), .B(n13131), .S(n13517), .Z(n13133) );
  NAND3_X1 U14861 ( .A1(n13135), .A2(n13134), .A3(n13133), .ZN(n13139) );
  MUX2_X1 U14862 ( .A(n13137), .B(n8040), .S(n13217), .Z(n13138) );
  NAND3_X1 U14863 ( .A1(n13139), .A2(n8041), .A3(n13138), .ZN(n13143) );
  MUX2_X1 U14864 ( .A(n13141), .B(n13140), .S(n13229), .Z(n13142) );
  AND3_X1 U14865 ( .A1(n13143), .A2(n13273), .A3(n13142), .ZN(n13152) );
  NAND2_X1 U14866 ( .A1(n13149), .A2(n13144), .ZN(n13147) );
  NAND2_X1 U14867 ( .A1(n13148), .A2(n13145), .ZN(n13146) );
  MUX2_X1 U14868 ( .A(n13147), .B(n13146), .S(n13229), .Z(n13151) );
  MUX2_X1 U14869 ( .A(n13149), .B(n13148), .S(n13217), .Z(n13150) );
  OAI21_X1 U14870 ( .B1(n13152), .B2(n13151), .A(n13150), .ZN(n13153) );
  NAND2_X1 U14871 ( .A1(n13153), .A2(n13275), .ZN(n13154) );
  OAI21_X1 U14872 ( .B1(n13229), .B2(n13331), .A(n13154), .ZN(n13161) );
  INV_X1 U14873 ( .A(n13155), .ZN(n13159) );
  AOI21_X1 U14874 ( .B1(n13157), .B2(n13156), .A(n13159), .ZN(n13158) );
  MUX2_X1 U14875 ( .A(n13159), .B(n13158), .S(n13229), .Z(n13160) );
  AOI211_X1 U14876 ( .C1(n13161), .C2(n8426), .A(n13160), .B(n13277), .ZN(
        n13162) );
  AOI21_X1 U14877 ( .B1(n13163), .B2(n13169), .A(n13162), .ZN(n13168) );
  INV_X1 U14878 ( .A(n13177), .ZN(n13174) );
  NAND2_X1 U14879 ( .A1(n13177), .A2(n8054), .ZN(n13165) );
  MUX2_X1 U14880 ( .A(n13166), .B(n13165), .S(n13217), .Z(n13167) );
  OAI21_X1 U14881 ( .B1(n13168), .B2(n13174), .A(n13167), .ZN(n13182) );
  INV_X1 U14882 ( .A(n13169), .ZN(n13172) );
  INV_X1 U14883 ( .A(n13175), .ZN(n13170) );
  AOI211_X1 U14884 ( .C1(n13172), .C2(n13171), .A(n14056), .B(n13170), .ZN(
        n13181) );
  OAI211_X1 U14885 ( .C1(n13174), .C2(n13173), .A(n13183), .B(n13175), .ZN(
        n13179) );
  NAND3_X1 U14886 ( .A1(n13175), .A2(n14049), .A3(n14237), .ZN(n13176) );
  NAND3_X1 U14887 ( .A1(n13184), .A2(n13177), .A3(n13176), .ZN(n13178) );
  MUX2_X1 U14888 ( .A(n13179), .B(n13178), .S(n13229), .Z(n13180) );
  AOI21_X1 U14889 ( .B1(n13182), .B2(n13181), .A(n13180), .ZN(n13188) );
  INV_X1 U14890 ( .A(n13183), .ZN(n13186) );
  INV_X1 U14891 ( .A(n13184), .ZN(n13185) );
  MUX2_X1 U14892 ( .A(n13186), .B(n13185), .S(n13217), .Z(n13187) );
  OAI21_X1 U14893 ( .B1(n13188), .B2(n13187), .A(n14011), .ZN(n13192) );
  MUX2_X1 U14894 ( .A(n13190), .B(n13189), .S(n13217), .Z(n13191) );
  NAND3_X1 U14895 ( .A1(n13192), .A2(n9813), .A3(n13191), .ZN(n13199) );
  MUX2_X1 U14896 ( .A(n13355), .B(n13352), .S(n13229), .Z(n13193) );
  INV_X1 U14897 ( .A(n13193), .ZN(n13197) );
  NAND2_X1 U14898 ( .A1(n14151), .A2(n13977), .ZN(n13195) );
  MUX2_X1 U14899 ( .A(n13195), .B(n13194), .S(n13217), .Z(n13196) );
  OAI21_X1 U14900 ( .B1(n13990), .B2(n13197), .A(n13196), .ZN(n13198) );
  OAI211_X1 U14901 ( .C1(n13199), .C2(n13990), .A(n13198), .B(n13979), .ZN(
        n13203) );
  NAND2_X1 U14902 ( .A1(n13392), .A2(n13966), .ZN(n13201) );
  MUX2_X1 U14903 ( .A(n13201), .B(n13200), .S(n13217), .Z(n13202) );
  INV_X1 U14904 ( .A(n13283), .ZN(n13962) );
  AOI21_X1 U14905 ( .B1(n13203), .B2(n13202), .A(n13962), .ZN(n13215) );
  OAI21_X1 U14906 ( .B1(n14214), .B2(n13511), .A(n13204), .ZN(n13206) );
  NAND2_X1 U14907 ( .A1(n13206), .A2(n13205), .ZN(n13209) );
  INV_X1 U14908 ( .A(n13207), .ZN(n13208) );
  AOI21_X1 U14909 ( .B1(n13210), .B2(n13209), .A(n13208), .ZN(n13213) );
  INV_X1 U14910 ( .A(n13213), .ZN(n13212) );
  NAND4_X1 U14911 ( .A1(n13930), .A2(n13962), .A3(n13940), .A4(n13952), .ZN(
        n13211) );
  NAND2_X1 U14912 ( .A1(n13212), .A2(n13211), .ZN(n13214) );
  NOR3_X1 U14913 ( .A1(n13412), .A2(n13932), .A3(n13217), .ZN(n13216) );
  NAND3_X1 U14914 ( .A1(n13227), .A2(n13218), .A3(n13217), .ZN(n13232) );
  INV_X1 U14915 ( .A(n13219), .ZN(n13220) );
  NAND2_X1 U14916 ( .A1(n13221), .A2(n13220), .ZN(n13223) );
  NAND2_X1 U14917 ( .A1(n15765), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13222) );
  NAND2_X1 U14918 ( .A1(n13223), .A2(n13222), .ZN(n13234) );
  XNOR2_X1 U14919 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n13233) );
  INV_X1 U14920 ( .A(n13233), .ZN(n13224) );
  XNOR2_X1 U14921 ( .A(n13234), .B(n13224), .ZN(n13317) );
  NAND2_X1 U14922 ( .A1(n13317), .A2(n13241), .ZN(n13226) );
  INV_X1 U14923 ( .A(SI_30_), .ZN(n13634) );
  OR2_X1 U14924 ( .A1(n9730), .A2(n13634), .ZN(n13225) );
  NAND2_X1 U14925 ( .A1(n13226), .A2(n13225), .ZN(n14196) );
  INV_X1 U14926 ( .A(n13509), .ZN(n13252) );
  NOR2_X1 U14927 ( .A1(n14196), .A2(n13252), .ZN(n13301) );
  INV_X1 U14928 ( .A(n13301), .ZN(n13288) );
  INV_X1 U14929 ( .A(n13295), .ZN(n13230) );
  OAI211_X1 U14930 ( .C1(n13230), .C2(n13229), .A(n13228), .B(n13297), .ZN(
        n13231) );
  NAND3_X1 U14931 ( .A1(n13232), .A2(n13288), .A3(n13231), .ZN(n13255) );
  NAND2_X1 U14932 ( .A1(n13234), .A2(n13233), .ZN(n13237) );
  NAND2_X1 U14933 ( .A1(n13235), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U14934 ( .A1(n13237), .A2(n13236), .ZN(n13240) );
  INV_X1 U14935 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13238) );
  XNOR2_X1 U14936 ( .A(n13238), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n13239) );
  XNOR2_X1 U14937 ( .A(n13240), .B(n13239), .ZN(n14258) );
  NAND2_X1 U14938 ( .A1(n14258), .A2(n13241), .ZN(n13243) );
  INV_X1 U14939 ( .A(SI_31_), .ZN(n14253) );
  OR2_X1 U14940 ( .A1(n9730), .A2(n14253), .ZN(n13242) );
  INV_X1 U14941 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14121) );
  NAND2_X1 U14942 ( .A1(n13244), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13248) );
  INV_X1 U14943 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13245) );
  OR2_X1 U14944 ( .A1(n13246), .A2(n13245), .ZN(n13247) );
  OAI211_X1 U14945 ( .C1(n9407), .C2(n14121), .A(n13248), .B(n13247), .ZN(
        n13249) );
  INV_X1 U14946 ( .A(n13249), .ZN(n13250) );
  OR2_X1 U14947 ( .A1(n14119), .A2(n13902), .ZN(n13254) );
  NAND2_X1 U14948 ( .A1(n14196), .A2(n13252), .ZN(n13253) );
  NAND2_X1 U14949 ( .A1(n13254), .A2(n13253), .ZN(n13299) );
  INV_X1 U14950 ( .A(n13299), .ZN(n13290) );
  AND2_X1 U14951 ( .A1(n14119), .A2(n13902), .ZN(n13300) );
  AOI21_X1 U14952 ( .B1(n13255), .B2(n13290), .A(n13300), .ZN(n13307) );
  INV_X1 U14953 ( .A(n13256), .ZN(n13285) );
  INV_X1 U14954 ( .A(n13257), .ZN(n13271) );
  NOR4_X1 U14955 ( .A1(n13261), .A2(n13260), .A3(n13259), .A4(n13258), .ZN(
        n13267) );
  NOR3_X1 U14956 ( .A1(n9807), .A2(n13264), .A3(n13263), .ZN(n13266) );
  NAND3_X1 U14957 ( .A1(n13267), .A2(n13266), .A3(n13265), .ZN(n13269) );
  NOR4_X1 U14958 ( .A1(n13271), .A2(n13270), .A3(n13269), .A4(n13268), .ZN(
        n13274) );
  NAND4_X1 U14959 ( .A1(n13275), .A2(n13274), .A3(n13273), .A4(n13272), .ZN(
        n13276) );
  NOR3_X1 U14960 ( .A1(n13277), .A2(n14105), .A3(n13276), .ZN(n13278) );
  NAND4_X1 U14961 ( .A1(n13279), .A2(n14068), .A3(n13278), .A4(n14074), .ZN(
        n13280) );
  NOR4_X1 U14962 ( .A1(n13999), .A2(n13281), .A3(n14034), .A4(n13280), .ZN(
        n13282) );
  NAND4_X1 U14963 ( .A1(n13283), .A2(n13282), .A3(n8028), .A4(n13979), .ZN(
        n13284) );
  NOR4_X1 U14964 ( .A1(n13286), .A2(n13285), .A3(n13915), .A4(n13284), .ZN(
        n13289) );
  INV_X1 U14965 ( .A(n13300), .ZN(n13287) );
  NAND4_X1 U14966 ( .A1(n13290), .A2(n13289), .A3(n13288), .A4(n13287), .ZN(
        n13291) );
  XNOR2_X1 U14967 ( .A(n13291), .B(n13888), .ZN(n13292) );
  INV_X1 U14968 ( .A(n14196), .ZN(n14124) );
  INV_X1 U14969 ( .A(n13902), .ZN(n13508) );
  OAI21_X1 U14970 ( .B1(n14124), .B2(n13508), .A(n13297), .ZN(n13298) );
  XNOR2_X1 U14971 ( .A(n13303), .B(n13888), .ZN(n13306) );
  INV_X1 U14972 ( .A(n13304), .ZN(n13305) );
  NAND3_X1 U14973 ( .A1(n13311), .A2(n13310), .A3(n13309), .ZN(n13312) );
  OAI211_X1 U14974 ( .C1(n13313), .C2(n13315), .A(n13312), .B(P3_B_REG_SCAN_IN), .ZN(n13314) );
  OAI21_X1 U14975 ( .B1(n13316), .B2(n13315), .A(n13314), .ZN(P3_U3296) );
  INV_X1 U14976 ( .A(n13317), .ZN(n13318) );
  OAI222_X1 U14977 ( .A1(n13320), .A2(P3_U3151), .B1(n14252), .B2(n13634), 
        .C1(n13319), .C2(n13318), .ZN(P3_U3265) );
  OAI222_X1 U14978 ( .A1(n14970), .A2(n13323), .B1(n14968), .B2(n13322), .C1(
        P2_U3088), .C2(n13321), .ZN(P2_U3300) );
  INV_X1 U14979 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13324) );
  NAND3_X1 U14980 ( .A1(n13324), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13328) );
  NAND2_X1 U14981 ( .A1(n15758), .A2(n13325), .ZN(n13327) );
  NAND2_X1 U14982 ( .A1(n14973), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13326) );
  OAI211_X1 U14983 ( .C1(n8607), .C2(n13328), .A(n13327), .B(n13326), .ZN(
        P2_U3296) );
  XNOR2_X1 U14984 ( .A(n13329), .B(n7765), .ZN(n13330) );
  NOR2_X1 U14985 ( .A1(n13330), .A2(n8011), .ZN(n13403) );
  AOI21_X1 U14986 ( .B1(n13330), .B2(n8011), .A(n13403), .ZN(n13374) );
  XNOR2_X1 U14987 ( .A(n16223), .B(n13405), .ZN(n13335) );
  XNOR2_X1 U14988 ( .A(n13335), .B(n13501), .ZN(n13378) );
  MUX2_X1 U14989 ( .A(n13332), .B(n13331), .S(n13405), .Z(n13379) );
  XNOR2_X1 U14990 ( .A(n14242), .B(n13405), .ZN(n13338) );
  XNOR2_X1 U14991 ( .A(n13338), .B(n14076), .ZN(n13496) );
  INV_X1 U14992 ( .A(n13335), .ZN(n13336) );
  NAND2_X1 U14993 ( .A1(n13336), .A2(n13501), .ZN(n13492) );
  NAND2_X1 U14994 ( .A1(n13338), .A2(n14106), .ZN(n13339) );
  XNOR2_X1 U14995 ( .A(n14179), .B(n13405), .ZN(n13432) );
  NAND2_X1 U14996 ( .A1(n13432), .A2(n13445), .ZN(n13340) );
  XNOR2_X1 U14997 ( .A(n14237), .B(n13405), .ZN(n13341) );
  XNOR2_X1 U14998 ( .A(n13341), .B(n14049), .ZN(n13441) );
  NAND2_X1 U14999 ( .A1(n13341), .A2(n14049), .ZN(n13342) );
  XNOR2_X1 U15000 ( .A(n14169), .B(n13405), .ZN(n13343) );
  XNOR2_X1 U15001 ( .A(n13343), .B(n14058), .ZN(n13477) );
  INV_X1 U15002 ( .A(n13343), .ZN(n13344) );
  NAND2_X1 U15003 ( .A1(n13344), .A2(n14058), .ZN(n13345) );
  XNOR2_X1 U15004 ( .A(n14039), .B(n13405), .ZN(n13346) );
  XNOR2_X1 U15005 ( .A(n13346), .B(n14050), .ZN(n13397) );
  INV_X1 U15006 ( .A(n13346), .ZN(n13347) );
  NAND2_X1 U15007 ( .A1(n13347), .A2(n14050), .ZN(n13348) );
  XNOR2_X1 U15008 ( .A(n14227), .B(n13405), .ZN(n13349) );
  XNOR2_X1 U15009 ( .A(n13349), .B(n14001), .ZN(n13459) );
  INV_X1 U15010 ( .A(n13349), .ZN(n13350) );
  NAND2_X1 U15011 ( .A1(n13350), .A2(n14001), .ZN(n13351) );
  INV_X1 U15012 ( .A(n13352), .ZN(n13353) );
  MUX2_X1 U15013 ( .A(n7312), .B(n13353), .S(n13405), .Z(n13414) );
  INV_X1 U15014 ( .A(n13414), .ZN(n13354) );
  MUX2_X1 U15015 ( .A(n13355), .B(n7334), .S(n7765), .Z(n13415) );
  XNOR2_X1 U15016 ( .A(n14151), .B(n13405), .ZN(n13357) );
  XNOR2_X1 U15017 ( .A(n13392), .B(n13405), .ZN(n13359) );
  XNOR2_X1 U15018 ( .A(n14218), .B(n7765), .ZN(n13361) );
  NAND2_X1 U15019 ( .A1(n13361), .A2(n13978), .ZN(n13425) );
  INV_X1 U15020 ( .A(n13361), .ZN(n13362) );
  NAND2_X1 U15021 ( .A1(n13362), .A2(n13512), .ZN(n13363) );
  XNOR2_X1 U15022 ( .A(n13364), .B(n13405), .ZN(n13365) );
  NAND2_X1 U15023 ( .A1(n13365), .A2(n13965), .ZN(n13368) );
  INV_X1 U15024 ( .A(n13365), .ZN(n13366) );
  NAND2_X1 U15025 ( .A1(n13366), .A2(n13511), .ZN(n13367) );
  AND2_X1 U15026 ( .A1(n13368), .A2(n13367), .ZN(n13426) );
  XNOR2_X1 U15027 ( .A(n13369), .B(n7765), .ZN(n13370) );
  NOR2_X1 U15028 ( .A1(n13370), .A2(n13510), .ZN(n13371) );
  AOI21_X1 U15029 ( .B1(n13370), .B2(n13510), .A(n13371), .ZN(n13486) );
  INV_X1 U15030 ( .A(n13371), .ZN(n13372) );
  AOI22_X1 U15031 ( .A1(n13933), .A2(n13503), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13375) );
  OAI21_X1 U15032 ( .B1(n13953), .B2(n13500), .A(n13375), .ZN(n13376) );
  AOI21_X1 U15033 ( .B1(n9769), .B2(n13498), .A(n13376), .ZN(n13377) );
  INV_X1 U15034 ( .A(n13493), .ZN(n13381) );
  AOI21_X1 U15035 ( .B1(n13334), .B2(n13379), .A(n13378), .ZN(n13380) );
  OAI21_X1 U15036 ( .B1(n13381), .B2(n13380), .A(n13495), .ZN(n13388) );
  INV_X1 U15037 ( .A(n14112), .ZN(n13386) );
  AOI21_X1 U15038 ( .B1(n13498), .B2(n14106), .A(n13382), .ZN(n13383) );
  OAI21_X1 U15039 ( .B1(n13384), .B2(n13500), .A(n13383), .ZN(n13385) );
  AOI21_X1 U15040 ( .B1(n13386), .B2(n13503), .A(n13385), .ZN(n13387) );
  OAI211_X1 U15041 ( .C1(n13507), .C2(n16223), .A(n13388), .B(n13387), .ZN(
        P3_U3155) );
  AOI21_X1 U15042 ( .B1(n13988), .B2(n13389), .A(n7200), .ZN(n13395) );
  INV_X1 U15043 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n13684) );
  OAI22_X1 U15044 ( .A1(n13977), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13684), .ZN(n13391) );
  NOR2_X1 U15045 ( .A1(n13978), .A2(n13470), .ZN(n13390) );
  AOI211_X1 U15046 ( .C1(n13982), .C2(n13503), .A(n13391), .B(n13390), .ZN(
        n13394) );
  NAND2_X1 U15047 ( .A1(n13392), .A2(n13411), .ZN(n13393) );
  OAI211_X1 U15048 ( .C1(n13395), .C2(n13440), .A(n13394), .B(n13393), .ZN(
        P3_U3156) );
  INV_X1 U15049 ( .A(n14039), .ZN(n14232) );
  OAI211_X1 U15050 ( .C1(n13398), .C2(n13397), .A(n13396), .B(n13495), .ZN(
        n13402) );
  NAND2_X1 U15051 ( .A1(n14001), .A2(n13498), .ZN(n13399) );
  NAND2_X1 U15052 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13893)
         );
  OAI211_X1 U15053 ( .C1(n14028), .C2(n13500), .A(n13399), .B(n13893), .ZN(
        n13400) );
  AOI21_X1 U15054 ( .B1(n14030), .B2(n13503), .A(n13400), .ZN(n13401) );
  OAI211_X1 U15055 ( .C1(n14232), .C2(n13507), .A(n13402), .B(n13401), .ZN(
        P3_U3159) );
  XNOR2_X1 U15056 ( .A(n13406), .B(n13405), .ZN(n13407) );
  NOR2_X1 U15057 ( .A1(n13919), .A2(n13470), .ZN(n13410) );
  AOI22_X1 U15058 ( .A1(n13923), .A2(n13503), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13408) );
  OAI21_X1 U15059 ( .B1(n13943), .B2(n13500), .A(n13408), .ZN(n13409) );
  AOI211_X1 U15060 ( .C1(n13412), .C2(n13411), .A(n13410), .B(n13409), .ZN(
        n13413) );
  INV_X1 U15061 ( .A(n14155), .ZN(n14007) );
  NAND2_X1 U15062 ( .A1(n13354), .A2(n13415), .ZN(n13416) );
  XNOR2_X1 U15063 ( .A(n13417), .B(n13416), .ZN(n13418) );
  NAND2_X1 U15064 ( .A1(n13418), .A2(n13495), .ZN(n13423) );
  OAI22_X1 U15065 ( .A1(n14029), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13419), .ZN(n13421) );
  NOR2_X1 U15066 ( .A1(n13977), .A2(n13470), .ZN(n13420) );
  AOI211_X1 U15067 ( .C1(n14005), .C2(n13503), .A(n13421), .B(n13420), .ZN(
        n13422) );
  OAI211_X1 U15068 ( .C1(n14007), .C2(n13507), .A(n13423), .B(n13422), .ZN(
        P3_U3163) );
  INV_X1 U15069 ( .A(n13424), .ZN(n13452) );
  NOR3_X1 U15070 ( .A1(n13452), .A2(n8336), .A3(n13426), .ZN(n13427) );
  OAI21_X1 U15071 ( .B1(n13427), .B2(n7289), .A(n13495), .ZN(n13431) );
  OAI22_X1 U15072 ( .A1(n13978), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13701), .ZN(n13429) );
  NOR2_X1 U15073 ( .A1(n13953), .A2(n13470), .ZN(n13428) );
  AOI211_X1 U15074 ( .C1(n13956), .C2(n13503), .A(n13429), .B(n13428), .ZN(
        n13430) );
  OAI211_X1 U15075 ( .C1(n14214), .C2(n13507), .A(n13431), .B(n13430), .ZN(
        P3_U3165) );
  XNOR2_X1 U15076 ( .A(n13432), .B(n14088), .ZN(n13433) );
  XNOR2_X1 U15077 ( .A(n13434), .B(n13433), .ZN(n13439) );
  NAND2_X1 U15078 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n13819)
         );
  NAND2_X1 U15079 ( .A1(n13498), .A2(n14049), .ZN(n13435) );
  OAI211_X1 U15080 ( .C1(n14076), .C2(n13500), .A(n13819), .B(n13435), .ZN(
        n13437) );
  INV_X1 U15081 ( .A(n14179), .ZN(n14081) );
  NOR2_X1 U15082 ( .A1(n14081), .A2(n13507), .ZN(n13436) );
  AOI211_X1 U15083 ( .C1(n14078), .C2(n13503), .A(n13437), .B(n13436), .ZN(
        n13438) );
  OAI21_X1 U15084 ( .B1(n13439), .B2(n13440), .A(n13438), .ZN(P3_U3166) );
  AOI21_X1 U15085 ( .B1(n13442), .B2(n13441), .A(n13440), .ZN(n13443) );
  NAND2_X1 U15086 ( .A1(n13443), .A2(n7202), .ZN(n13448) );
  NAND2_X1 U15087 ( .A1(n14058), .A2(n13498), .ZN(n13444) );
  NAND2_X1 U15088 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13840)
         );
  OAI211_X1 U15089 ( .C1(n13445), .C2(n13500), .A(n13444), .B(n13840), .ZN(
        n13446) );
  AOI21_X1 U15090 ( .B1(n14061), .B2(n13503), .A(n13446), .ZN(n13447) );
  OAI211_X1 U15091 ( .C1(n13507), .C2(n14237), .A(n13448), .B(n13447), .ZN(
        P3_U3168) );
  INV_X1 U15092 ( .A(n13449), .ZN(n13451) );
  NOR3_X1 U15093 ( .A1(n7200), .A2(n13451), .A3(n13450), .ZN(n13453) );
  OAI21_X1 U15094 ( .B1(n13453), .B2(n13452), .A(n13495), .ZN(n13457) );
  OAI22_X1 U15095 ( .A1(n13966), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13712), .ZN(n13455) );
  NOR2_X1 U15096 ( .A1(n13965), .A2(n13470), .ZN(n13454) );
  AOI211_X1 U15097 ( .C1(n13967), .C2(n13503), .A(n13455), .B(n13454), .ZN(
        n13456) );
  OAI211_X1 U15098 ( .C1(n14218), .C2(n13507), .A(n13457), .B(n13456), .ZN(
        P3_U3169) );
  INV_X1 U15099 ( .A(n14227), .ZN(n13466) );
  OAI211_X1 U15100 ( .C1(n13460), .C2(n13459), .A(n13458), .B(n13495), .ZN(
        n13465) );
  AOI22_X1 U15101 ( .A1(n14015), .A2(n13498), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13461) );
  OAI21_X1 U15102 ( .B1(n13462), .B2(n13500), .A(n13461), .ZN(n13463) );
  AOI21_X1 U15103 ( .B1(n14020), .B2(n13503), .A(n13463), .ZN(n13464) );
  OAI211_X1 U15104 ( .C1(n13466), .C2(n13507), .A(n13465), .B(n13464), .ZN(
        P3_U3173) );
  OAI21_X1 U15105 ( .B1(n7347), .B2(n13977), .A(n13467), .ZN(n13468) );
  NAND2_X1 U15106 ( .A1(n13468), .A2(n13495), .ZN(n13474) );
  INV_X1 U15107 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13720) );
  OAI22_X1 U15108 ( .A1(n13469), .A2(n13500), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13720), .ZN(n13472) );
  NOR2_X1 U15109 ( .A1(n13966), .A2(n13470), .ZN(n13471) );
  AOI211_X1 U15110 ( .C1(n13994), .C2(n13503), .A(n13472), .B(n13471), .ZN(
        n13473) );
  OAI211_X1 U15111 ( .C1(n13475), .C2(n13507), .A(n13474), .B(n13473), .ZN(
        P3_U3175) );
  INV_X1 U15112 ( .A(n14169), .ZN(n13483) );
  OAI211_X1 U15113 ( .C1(n13478), .C2(n13477), .A(n13476), .B(n13495), .ZN(
        n13482) );
  NAND2_X1 U15114 ( .A1(n14050), .A2(n13498), .ZN(n13479) );
  NAND2_X1 U15115 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13873)
         );
  OAI211_X1 U15116 ( .C1(n14077), .C2(n13500), .A(n13479), .B(n13873), .ZN(
        n13480) );
  AOI21_X1 U15117 ( .B1(n14043), .B2(n13503), .A(n13480), .ZN(n13481) );
  OAI211_X1 U15118 ( .C1(n13483), .C2(n13507), .A(n13482), .B(n13481), .ZN(
        P3_U3178) );
  OAI21_X1 U15119 ( .B1(n13486), .B2(n13485), .A(n13484), .ZN(n13487) );
  NAND2_X1 U15120 ( .A1(n13487), .A2(n13495), .ZN(n13491) );
  AOI22_X1 U15121 ( .A1(n13944), .A2(n13503), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13488) );
  OAI21_X1 U15122 ( .B1(n13965), .B2(n13500), .A(n13488), .ZN(n13489) );
  AOI21_X1 U15123 ( .B1(n8011), .B2(n13498), .A(n13489), .ZN(n13490) );
  OAI211_X1 U15124 ( .C1(n14210), .C2(n13507), .A(n13491), .B(n13490), .ZN(
        P3_U3180) );
  AND2_X1 U15125 ( .A1(n13493), .A2(n13492), .ZN(n13497) );
  OAI211_X1 U15126 ( .C1(n13497), .C2(n13496), .A(n13495), .B(n13494), .ZN(
        n13506) );
  INV_X1 U15127 ( .A(n14095), .ZN(n13504) );
  AND2_X1 U15128 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13794) );
  AOI21_X1 U15129 ( .B1(n13498), .B2(n14088), .A(n13794), .ZN(n13499) );
  OAI21_X1 U15130 ( .B1(n13501), .B2(n13500), .A(n13499), .ZN(n13502) );
  AOI21_X1 U15131 ( .B1(n13504), .B2(n13503), .A(n13502), .ZN(n13505) );
  OAI211_X1 U15132 ( .C1(n13507), .C2(n14242), .A(n13506), .B(n13505), .ZN(
        P3_U3181) );
  MUX2_X1 U15133 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13508), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15134 ( .A(n13509), .B(P3_DATAO_REG_30__SCAN_IN), .S(n13739), .Z(
        P3_U3521) );
  MUX2_X1 U15135 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n9769), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15136 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n8011), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15137 ( .A(n13510), .B(P3_DATAO_REG_26__SCAN_IN), .S(n13739), .Z(
        P3_U3517) );
  MUX2_X1 U15138 ( .A(n13511), .B(P3_DATAO_REG_25__SCAN_IN), .S(n13739), .Z(
        P3_U3516) );
  MUX2_X1 U15139 ( .A(n13512), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13739), .Z(
        P3_U3515) );
  MUX2_X1 U15140 ( .A(n13988), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13739), .Z(
        P3_U3514) );
  MUX2_X1 U15141 ( .A(n14002), .B(P3_DATAO_REG_22__SCAN_IN), .S(n13739), .Z(
        P3_U3513) );
  MUX2_X1 U15142 ( .A(n14015), .B(P3_DATAO_REG_21__SCAN_IN), .S(n13739), .Z(
        P3_U3512) );
  MUX2_X1 U15143 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n14001), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15144 ( .A(n14050), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13739), .Z(
        P3_U3510) );
  MUX2_X1 U15145 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n14058), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15146 ( .A(n14049), .B(P3_DATAO_REG_17__SCAN_IN), .S(n13739), .Z(
        P3_U3508) );
  MUX2_X1 U15147 ( .A(n14088), .B(P3_DATAO_REG_16__SCAN_IN), .S(n13739), .Z(
        P3_U3507) );
  MUX2_X1 U15148 ( .A(n14106), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13739), .Z(
        P3_U3506) );
  MUX2_X1 U15149 ( .A(n14089), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13739), .Z(
        P3_U3505) );
  MUX2_X1 U15150 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n14109), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15151 ( .A(n13513), .B(P3_DATAO_REG_12__SCAN_IN), .S(n13739), .Z(
        P3_U3503) );
  MUX2_X1 U15152 ( .A(n13514), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13739), .Z(
        P3_U3502) );
  MUX2_X1 U15153 ( .A(n13515), .B(P3_DATAO_REG_10__SCAN_IN), .S(n13739), .Z(
        P3_U3501) );
  MUX2_X1 U15154 ( .A(n13516), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13739), .Z(
        P3_U3500) );
  MUX2_X1 U15155 ( .A(n13517), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13739), .Z(
        P3_U3499) );
  MUX2_X1 U15156 ( .A(n13518), .B(P3_DATAO_REG_7__SCAN_IN), .S(n13739), .Z(
        P3_U3498) );
  MUX2_X1 U15157 ( .A(n13519), .B(P3_DATAO_REG_6__SCAN_IN), .S(n13739), .Z(
        P3_U3497) );
  MUX2_X1 U15158 ( .A(n13520), .B(P3_DATAO_REG_5__SCAN_IN), .S(n13739), .Z(
        P3_U3496) );
  MUX2_X1 U15159 ( .A(n13521), .B(P3_DATAO_REG_4__SCAN_IN), .S(n13739), .Z(
        P3_U3495) );
  MUX2_X1 U15160 ( .A(n13522), .B(P3_DATAO_REG_3__SCAN_IN), .S(n13739), .Z(
        P3_U3494) );
  MUX2_X1 U15161 ( .A(n13523), .B(P3_DATAO_REG_2__SCAN_IN), .S(n13739), .Z(
        n13737) );
  OAI22_X1 U15162 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_60), .B1(
        keyinput_61), .B2(P3_REG3_REG_6__SCAN_IN), .ZN(n13524) );
  AOI221_X1 U15163 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .C1(
        P3_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n13524), .ZN(n13612) );
  INV_X1 U15164 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n13717) );
  INV_X1 U15165 ( .A(keyinput_55), .ZN(n13605) );
  OAI22_X1 U15166 ( .A1(n9349), .A2(keyinput_53), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_52), .ZN(n13525) );
  AOI221_X1 U15167 ( .B1(n9349), .B2(keyinput_53), .C1(keyinput_52), .C2(
        P3_REG3_REG_4__SCAN_IN), .A(n13525), .ZN(n13602) );
  INV_X1 U15168 ( .A(keyinput_51), .ZN(n13600) );
  INV_X1 U15169 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13617) );
  AOI22_X1 U15170 ( .A1(n9346), .A2(keyinput_49), .B1(n13617), .B2(keyinput_48), .ZN(n13526) );
  OAI221_X1 U15171 ( .B1(n9346), .B2(keyinput_49), .C1(n13617), .C2(
        keyinput_48), .A(n13526), .ZN(n13598) );
  OAI22_X1 U15172 ( .A1(n13701), .A2(keyinput_47), .B1(n13419), .B2(
        keyinput_45), .ZN(n13527) );
  AOI221_X1 U15173 ( .B1(n13701), .B2(keyinput_47), .C1(keyinput_45), .C2(
        n13419), .A(n13527), .ZN(n13594) );
  OAI22_X1 U15174 ( .A1(P3_REG3_REG_28__SCAN_IN), .A2(keyinput_42), .B1(
        P3_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .ZN(n13528) );
  AOI221_X1 U15175 ( .B1(P3_REG3_REG_28__SCAN_IN), .B2(keyinput_42), .C1(
        keyinput_43), .C2(P3_REG3_REG_8__SCAN_IN), .A(n13528), .ZN(n13591) );
  AOI22_X1 U15176 ( .A1(SI_4_), .A2(keyinput_28), .B1(SI_5_), .B2(keyinput_27), 
        .ZN(n13529) );
  OAI221_X1 U15177 ( .B1(SI_4_), .B2(keyinput_28), .C1(SI_5_), .C2(keyinput_27), .A(n13529), .ZN(n13571) );
  OAI22_X1 U15178 ( .A1(SI_9_), .A2(keyinput_23), .B1(keyinput_24), .B2(SI_8_), 
        .ZN(n13530) );
  AOI221_X1 U15179 ( .B1(SI_9_), .B2(keyinput_23), .C1(SI_8_), .C2(keyinput_24), .A(n13530), .ZN(n13569) );
  INV_X1 U15180 ( .A(keyinput_22), .ZN(n13564) );
  INV_X1 U15181 ( .A(keyinput_21), .ZN(n13562) );
  INV_X1 U15182 ( .A(keyinput_17), .ZN(n13556) );
  INV_X1 U15183 ( .A(keyinput_10), .ZN(n13547) );
  INV_X1 U15184 ( .A(keyinput_9), .ZN(n13545) );
  INV_X1 U15185 ( .A(keyinput_8), .ZN(n13543) );
  INV_X1 U15186 ( .A(keyinput_7), .ZN(n13541) );
  INV_X1 U15187 ( .A(SI_25_), .ZN(n13643) );
  INV_X1 U15188 ( .A(keyinput_6), .ZN(n13539) );
  OAI22_X1 U15189 ( .A1(SI_31_), .A2(keyinput_1), .B1(P3_WR_REG_SCAN_IN), .B2(
        keyinput_0), .ZN(n13531) );
  AOI221_X1 U15190 ( .B1(SI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P3_WR_REG_SCAN_IN), .A(n13531), .ZN(n13537) );
  AOI22_X1 U15191 ( .A1(n12394), .A2(keyinput_3), .B1(keyinput_5), .B2(n13632), 
        .ZN(n13532) );
  OAI221_X1 U15192 ( .B1(n12394), .B2(keyinput_3), .C1(n13632), .C2(keyinput_5), .A(n13532), .ZN(n13536) );
  INV_X1 U15193 ( .A(SI_28_), .ZN(n13534) );
  AOI22_X1 U15194 ( .A1(SI_30_), .A2(keyinput_2), .B1(n13534), .B2(keyinput_4), 
        .ZN(n13533) );
  OAI221_X1 U15195 ( .B1(SI_30_), .B2(keyinput_2), .C1(n13534), .C2(keyinput_4), .A(n13533), .ZN(n13535) );
  NOR3_X1 U15196 ( .A1(n13537), .A2(n13536), .A3(n13535), .ZN(n13538) );
  AOI221_X1 U15197 ( .B1(SI_26_), .B2(keyinput_6), .C1(n13640), .C2(n13539), 
        .A(n13538), .ZN(n13540) );
  AOI221_X1 U15198 ( .B1(SI_25_), .B2(n13541), .C1(n13643), .C2(keyinput_7), 
        .A(n13540), .ZN(n13542) );
  AOI221_X1 U15199 ( .B1(SI_24_), .B2(keyinput_8), .C1(n13646), .C2(n13543), 
        .A(n13542), .ZN(n13544) );
  AOI221_X1 U15200 ( .B1(SI_23_), .B2(n13545), .C1(n13650), .C2(keyinput_9), 
        .A(n13544), .ZN(n13546) );
  AOI221_X1 U15201 ( .B1(SI_22_), .B2(keyinput_10), .C1(n13652), .C2(n13547), 
        .A(n13546), .ZN(n13554) );
  AOI22_X1 U15202 ( .A1(SI_19_), .A2(keyinput_13), .B1(SI_21_), .B2(
        keyinput_11), .ZN(n13548) );
  OAI221_X1 U15203 ( .B1(SI_19_), .B2(keyinput_13), .C1(SI_21_), .C2(
        keyinput_11), .A(n13548), .ZN(n13553) );
  AOI22_X1 U15204 ( .A1(SI_20_), .A2(keyinput_12), .B1(n13627), .B2(
        keyinput_15), .ZN(n13549) );
  OAI221_X1 U15205 ( .B1(SI_20_), .B2(keyinput_12), .C1(n13627), .C2(
        keyinput_15), .A(n13549), .ZN(n13552) );
  AOI22_X1 U15206 ( .A1(n13629), .A2(keyinput_16), .B1(n13630), .B2(
        keyinput_14), .ZN(n13550) );
  OAI221_X1 U15207 ( .B1(n13629), .B2(keyinput_16), .C1(n13630), .C2(
        keyinput_14), .A(n13550), .ZN(n13551) );
  NOR4_X1 U15208 ( .A1(n13554), .A2(n13553), .A3(n13552), .A4(n13551), .ZN(
        n13555) );
  AOI221_X1 U15209 ( .B1(SI_15_), .B2(n13556), .C1(n13659), .C2(keyinput_17), 
        .A(n13555), .ZN(n13559) );
  AOI22_X1 U15210 ( .A1(SI_12_), .A2(keyinput_20), .B1(SI_13_), .B2(
        keyinput_19), .ZN(n13557) );
  OAI221_X1 U15211 ( .B1(SI_12_), .B2(keyinput_20), .C1(SI_13_), .C2(
        keyinput_19), .A(n13557), .ZN(n13558) );
  AOI211_X1 U15212 ( .C1(SI_14_), .C2(keyinput_18), .A(n13559), .B(n13558), 
        .ZN(n13560) );
  OAI21_X1 U15213 ( .B1(SI_14_), .B2(keyinput_18), .A(n13560), .ZN(n13561) );
  OAI221_X1 U15214 ( .B1(SI_11_), .B2(n13562), .C1(n13666), .C2(keyinput_21), 
        .A(n13561), .ZN(n13563) );
  OAI221_X1 U15215 ( .B1(SI_10_), .B2(keyinput_22), .C1(n13669), .C2(n13564), 
        .A(n13563), .ZN(n13568) );
  AOI22_X1 U15216 ( .A1(n13566), .A2(keyinput_26), .B1(n13673), .B2(
        keyinput_25), .ZN(n13565) );
  OAI221_X1 U15217 ( .B1(n13566), .B2(keyinput_26), .C1(n13673), .C2(
        keyinput_25), .A(n13565), .ZN(n13567) );
  AOI21_X1 U15218 ( .B1(n13569), .B2(n13568), .A(n13567), .ZN(n13570) );
  OAI22_X1 U15219 ( .A1(n13571), .A2(n13570), .B1(SI_1_), .B2(keyinput_31), 
        .ZN(n13572) );
  AOI21_X1 U15220 ( .B1(SI_1_), .B2(keyinput_31), .A(n13572), .ZN(n13584) );
  OAI22_X1 U15221 ( .A1(SI_3_), .A2(keyinput_29), .B1(SI_2_), .B2(keyinput_30), 
        .ZN(n13573) );
  AOI221_X1 U15222 ( .B1(SI_3_), .B2(keyinput_29), .C1(keyinput_30), .C2(SI_2_), .A(n13573), .ZN(n13583) );
  AOI22_X1 U15223 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_36), .B1(n13684), .B2(keyinput_38), .ZN(n13574) );
  OAI221_X1 U15224 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .C1(
        n13684), .C2(keyinput_38), .A(n13574), .ZN(n13582) );
  AOI22_X1 U15225 ( .A1(n13576), .A2(keyinput_37), .B1(P3_U3151), .B2(
        keyinput_34), .ZN(n13575) );
  OAI221_X1 U15226 ( .B1(n13576), .B2(keyinput_37), .C1(P3_U3151), .C2(
        keyinput_34), .A(n13575), .ZN(n13579) );
  INV_X1 U15227 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15999) );
  AOI22_X1 U15228 ( .A1(n15999), .A2(keyinput_33), .B1(n10380), .B2(
        keyinput_32), .ZN(n13577) );
  OAI221_X1 U15229 ( .B1(n15999), .B2(keyinput_33), .C1(n10380), .C2(
        keyinput_32), .A(n13577), .ZN(n13578) );
  AOI211_X1 U15230 ( .C1(keyinput_35), .C2(P3_REG3_REG_7__SCAN_IN), .A(n13579), 
        .B(n13578), .ZN(n13580) );
  OAI21_X1 U15231 ( .B1(keyinput_35), .B2(P3_REG3_REG_7__SCAN_IN), .A(n13580), 
        .ZN(n13581) );
  AOI211_X1 U15232 ( .C1(n13584), .C2(n13583), .A(n13582), .B(n13581), .ZN(
        n13588) );
  AOI22_X1 U15233 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_39), .B1(n13586), .B2(keyinput_41), .ZN(n13585) );
  OAI221_X1 U15234 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .C1(
        n13586), .C2(keyinput_41), .A(n13585), .ZN(n13587) );
  AOI211_X1 U15235 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(keyinput_40), .A(n13588), 
        .B(n13587), .ZN(n13589) );
  OAI21_X1 U15236 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .A(n13589), 
        .ZN(n13590) );
  AOI22_X1 U15237 ( .A1(n13591), .A2(n13590), .B1(keyinput_44), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n13592) );
  OAI21_X1 U15238 ( .B1(keyinput_44), .B2(P3_REG3_REG_1__SCAN_IN), .A(n13592), 
        .ZN(n13593) );
  OAI211_X1 U15239 ( .C1(n13705), .C2(keyinput_46), .A(n13594), .B(n13593), 
        .ZN(n13595) );
  AOI21_X1 U15240 ( .B1(n13705), .B2(keyinput_46), .A(n13595), .ZN(n13597) );
  NAND2_X1 U15241 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_50), .ZN(n13596) );
  OAI221_X1 U15242 ( .B1(n13598), .B2(n13597), .C1(P3_REG3_REG_17__SCAN_IN), 
        .C2(keyinput_50), .A(n13596), .ZN(n13599) );
  OAI221_X1 U15243 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(n13600), .C1(n13712), 
        .C2(keyinput_51), .A(n13599), .ZN(n13601) );
  OAI211_X1 U15244 ( .C1(P3_REG3_REG_0__SCAN_IN), .C2(keyinput_54), .A(n13602), 
        .B(n13601), .ZN(n13603) );
  AOI21_X1 U15245 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .A(n13603), 
        .ZN(n13604) );
  AOI221_X1 U15246 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_55), .C1(
        n13717), .C2(n13605), .A(n13604), .ZN(n13610) );
  AOI22_X1 U15247 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(keyinput_56), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .ZN(n13606) );
  OAI221_X1 U15248 ( .B1(P3_REG3_REG_13__SCAN_IN), .B2(keyinput_56), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_57), .A(n13606), .ZN(n13609) );
  OAI22_X1 U15249 ( .A1(n16044), .A2(keyinput_59), .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .ZN(n13607) );
  AOI221_X1 U15250 ( .B1(n16044), .B2(keyinput_59), .C1(keyinput_58), .C2(
        P3_REG3_REG_11__SCAN_IN), .A(n13607), .ZN(n13608) );
  OAI21_X1 U15251 ( .B1(n13610), .B2(n13609), .A(n13608), .ZN(n13611) );
  INV_X1 U15252 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n13734) );
  AOI22_X1 U15253 ( .A1(n13612), .A2(n13611), .B1(keyinput_62), .B2(n13734), 
        .ZN(n13735) );
  OAI22_X1 U15254 ( .A1(n13614), .A2(keyinput_125), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .ZN(n13613) );
  AOI221_X1 U15255 ( .B1(n13614), .B2(keyinput_125), .C1(keyinput_124), .C2(
        P3_REG3_REG_18__SCAN_IN), .A(n13613), .ZN(n13727) );
  INV_X1 U15256 ( .A(keyinput_119), .ZN(n13718) );
  OAI22_X1 U15257 ( .A1(n9349), .A2(keyinput_117), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_116), .ZN(n13615) );
  AOI221_X1 U15258 ( .B1(n9349), .B2(keyinput_117), .C1(keyinput_116), .C2(
        P3_REG3_REG_4__SCAN_IN), .A(n13615), .ZN(n13714) );
  INV_X1 U15259 ( .A(keyinput_115), .ZN(n13711) );
  OAI22_X1 U15260 ( .A1(n13617), .A2(keyinput_112), .B1(keyinput_113), .B2(
        P3_REG3_REG_5__SCAN_IN), .ZN(n13616) );
  AOI221_X1 U15261 ( .B1(n13617), .B2(keyinput_112), .C1(
        P3_REG3_REG_5__SCAN_IN), .C2(keyinput_113), .A(n13616), .ZN(n13707) );
  INV_X1 U15262 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13619) );
  AOI22_X1 U15263 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(n13619), .B2(keyinput_106), .ZN(n13618) );
  OAI221_X1 U15264 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        n13619), .C2(keyinput_106), .A(n13618), .ZN(n13698) );
  OAI22_X1 U15265 ( .A1(n13621), .A2(keyinput_103), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_105), .ZN(n13620) );
  AOI221_X1 U15266 ( .B1(n13621), .B2(keyinput_103), .C1(keyinput_105), .C2(
        P3_REG3_REG_19__SCAN_IN), .A(n13620), .ZN(n13694) );
  OAI22_X1 U15267 ( .A1(SI_5_), .A2(keyinput_91), .B1(SI_4_), .B2(keyinput_92), 
        .ZN(n13622) );
  AOI221_X1 U15268 ( .B1(SI_5_), .B2(keyinput_91), .C1(keyinput_92), .C2(SI_4_), .A(n13622), .ZN(n13678) );
  INV_X1 U15269 ( .A(keyinput_86), .ZN(n13668) );
  INV_X1 U15270 ( .A(keyinput_85), .ZN(n13665) );
  OAI22_X1 U15271 ( .A1(n13624), .A2(keyinput_82), .B1(SI_13_), .B2(
        keyinput_83), .ZN(n13623) );
  AOI221_X1 U15272 ( .B1(n13624), .B2(keyinput_82), .C1(keyinput_83), .C2(
        SI_13_), .A(n13623), .ZN(n13662) );
  INV_X1 U15273 ( .A(keyinput_81), .ZN(n13660) );
  OAI22_X1 U15274 ( .A1(SI_21_), .A2(keyinput_75), .B1(keyinput_76), .B2(
        SI_20_), .ZN(n13625) );
  AOI221_X1 U15275 ( .B1(SI_21_), .B2(keyinput_75), .C1(SI_20_), .C2(
        keyinput_76), .A(n13625), .ZN(n13657) );
  OAI22_X1 U15276 ( .A1(n13627), .A2(keyinput_79), .B1(keyinput_77), .B2(
        SI_19_), .ZN(n13626) );
  AOI221_X1 U15277 ( .B1(n13627), .B2(keyinput_79), .C1(SI_19_), .C2(
        keyinput_77), .A(n13626), .ZN(n13656) );
  OAI22_X1 U15278 ( .A1(n13630), .A2(keyinput_78), .B1(n13629), .B2(
        keyinput_80), .ZN(n13628) );
  AOI221_X1 U15279 ( .B1(n13630), .B2(keyinput_78), .C1(keyinput_80), .C2(
        n13629), .A(n13628), .ZN(n13655) );
  INV_X1 U15280 ( .A(keyinput_74), .ZN(n13653) );
  INV_X1 U15281 ( .A(keyinput_73), .ZN(n13649) );
  INV_X1 U15282 ( .A(keyinput_72), .ZN(n13647) );
  INV_X1 U15283 ( .A(keyinput_71), .ZN(n13644) );
  INV_X1 U15284 ( .A(keyinput_70), .ZN(n13641) );
  OAI22_X1 U15285 ( .A1(n12394), .A2(keyinput_67), .B1(n13632), .B2(
        keyinput_69), .ZN(n13631) );
  AOI221_X1 U15286 ( .B1(n12394), .B2(keyinput_67), .C1(keyinput_69), .C2(
        n13632), .A(n13631), .ZN(n13638) );
  OAI22_X1 U15287 ( .A1(n13634), .A2(keyinput_66), .B1(SI_28_), .B2(
        keyinput_68), .ZN(n13633) );
  AOI221_X1 U15288 ( .B1(n13634), .B2(keyinput_66), .C1(keyinput_68), .C2(
        SI_28_), .A(n13633), .ZN(n13637) );
  AOI22_X1 U15289 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n13635) );
  OAI221_X1 U15290 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n13635), .ZN(n13636) );
  NAND3_X1 U15291 ( .A1(n13638), .A2(n13637), .A3(n13636), .ZN(n13639) );
  OAI221_X1 U15292 ( .B1(SI_26_), .B2(n13641), .C1(n13640), .C2(keyinput_70), 
        .A(n13639), .ZN(n13642) );
  OAI221_X1 U15293 ( .B1(SI_25_), .B2(n13644), .C1(n13643), .C2(keyinput_71), 
        .A(n13642), .ZN(n13645) );
  OAI221_X1 U15294 ( .B1(SI_24_), .B2(n13647), .C1(n13646), .C2(keyinput_72), 
        .A(n13645), .ZN(n13648) );
  OAI221_X1 U15295 ( .B1(SI_23_), .B2(keyinput_73), .C1(n13650), .C2(n13649), 
        .A(n13648), .ZN(n13651) );
  OAI221_X1 U15296 ( .B1(SI_22_), .B2(n13653), .C1(n13652), .C2(keyinput_74), 
        .A(n13651), .ZN(n13654) );
  NAND4_X1 U15297 ( .A1(n13657), .A2(n13656), .A3(n13655), .A4(n13654), .ZN(
        n13658) );
  OAI221_X1 U15298 ( .B1(SI_15_), .B2(n13660), .C1(n13659), .C2(keyinput_81), 
        .A(n13658), .ZN(n13661) );
  OAI211_X1 U15299 ( .C1(SI_12_), .C2(keyinput_84), .A(n13662), .B(n13661), 
        .ZN(n13663) );
  AOI21_X1 U15300 ( .B1(SI_12_), .B2(keyinput_84), .A(n13663), .ZN(n13664) );
  AOI221_X1 U15301 ( .B1(SI_11_), .B2(keyinput_85), .C1(n13666), .C2(n13665), 
        .A(n13664), .ZN(n13667) );
  AOI221_X1 U15302 ( .B1(SI_10_), .B2(keyinput_86), .C1(n13669), .C2(n13668), 
        .A(n13667), .ZN(n13676) );
  AOI22_X1 U15303 ( .A1(SI_9_), .A2(keyinput_87), .B1(n13671), .B2(keyinput_88), .ZN(n13670) );
  OAI221_X1 U15304 ( .B1(SI_9_), .B2(keyinput_87), .C1(n13671), .C2(
        keyinput_88), .A(n13670), .ZN(n13675) );
  OAI22_X1 U15305 ( .A1(n13673), .A2(keyinput_89), .B1(keyinput_90), .B2(SI_6_), .ZN(n13672) );
  AOI221_X1 U15306 ( .B1(n13673), .B2(keyinput_89), .C1(SI_6_), .C2(
        keyinput_90), .A(n13672), .ZN(n13674) );
  OAI21_X1 U15307 ( .B1(n13676), .B2(n13675), .A(n13674), .ZN(n13677) );
  AOI22_X1 U15308 ( .A1(n13678), .A2(n13677), .B1(SI_3_), .B2(keyinput_93), 
        .ZN(n13679) );
  OAI21_X1 U15309 ( .B1(SI_3_), .B2(keyinput_93), .A(n13679), .ZN(n13692) );
  XOR2_X1 U15310 ( .A(n10173), .B(keyinput_95), .Z(n13681) );
  XNOR2_X1 U15311 ( .A(SI_2_), .B(keyinput_94), .ZN(n13680) );
  NAND2_X1 U15312 ( .A1(n13681), .A2(n13680), .ZN(n13691) );
  OAI22_X1 U15313 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_100), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .ZN(n13682) );
  AOI221_X1 U15314 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .C1(
        keyinput_101), .C2(P3_REG3_REG_14__SCAN_IN), .A(n13682), .ZN(n13686)
         );
  OAI22_X1 U15315 ( .A1(n13684), .A2(keyinput_102), .B1(n10380), .B2(
        keyinput_96), .ZN(n13683) );
  AOI221_X1 U15316 ( .B1(n13684), .B2(keyinput_102), .C1(keyinput_96), .C2(
        n10380), .A(n13683), .ZN(n13685) );
  OAI211_X1 U15317 ( .C1(P3_U3151), .C2(keyinput_98), .A(n13686), .B(n13685), 
        .ZN(n13687) );
  AOI21_X1 U15318 ( .B1(P3_U3151), .B2(keyinput_98), .A(n13687), .ZN(n13690)
         );
  OAI22_X1 U15319 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(keyinput_99), .B1(
        keyinput_97), .B2(P3_RD_REG_SCAN_IN), .ZN(n13688) );
  AOI221_X1 U15320 ( .B1(P3_REG3_REG_7__SCAN_IN), .B2(keyinput_99), .C1(
        P3_RD_REG_SCAN_IN), .C2(keyinput_97), .A(n13688), .ZN(n13689) );
  OAI211_X1 U15321 ( .C1(n13692), .C2(n13691), .A(n13690), .B(n13689), .ZN(
        n13693) );
  OAI211_X1 U15322 ( .C1(n13696), .C2(keyinput_104), .A(n13694), .B(n13693), 
        .ZN(n13695) );
  AOI21_X1 U15323 ( .B1(n13696), .B2(keyinput_104), .A(n13695), .ZN(n13697) );
  OAI22_X1 U15324 ( .A1(keyinput_108), .A2(n10603), .B1(n13698), .B2(n13697), 
        .ZN(n13699) );
  AOI21_X1 U15325 ( .B1(keyinput_108), .B2(n10603), .A(n13699), .ZN(n13703) );
  AOI22_X1 U15326 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_109), .B1(
        n13701), .B2(keyinput_111), .ZN(n13700) );
  OAI221_X1 U15327 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .C1(
        n13701), .C2(keyinput_111), .A(n13700), .ZN(n13702) );
  AOI211_X1 U15328 ( .C1(n13705), .C2(keyinput_110), .A(n13703), .B(n13702), 
        .ZN(n13704) );
  OAI21_X1 U15329 ( .B1(n13705), .B2(keyinput_110), .A(n13704), .ZN(n13706) );
  AOI22_X1 U15330 ( .A1(keyinput_114), .A2(n13709), .B1(n13707), .B2(n13706), 
        .ZN(n13708) );
  OAI21_X1 U15331 ( .B1(n13709), .B2(keyinput_114), .A(n13708), .ZN(n13710) );
  OAI221_X1 U15332 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .C1(
        n13712), .C2(n13711), .A(n13710), .ZN(n13713) );
  OAI211_X1 U15333 ( .C1(P3_REG3_REG_0__SCAN_IN), .C2(keyinput_118), .A(n13714), .B(n13713), .ZN(n13715) );
  AOI21_X1 U15334 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .A(n13715), 
        .ZN(n13716) );
  AOI221_X1 U15335 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(n13718), .C1(n13717), 
        .C2(keyinput_119), .A(n13716), .ZN(n13725) );
  AOI22_X1 U15336 ( .A1(n9351), .A2(keyinput_120), .B1(n13720), .B2(
        keyinput_121), .ZN(n13719) );
  OAI221_X1 U15337 ( .B1(n9351), .B2(keyinput_120), .C1(n13720), .C2(
        keyinput_121), .A(n13719), .ZN(n13724) );
  OAI22_X1 U15338 ( .A1(n13722), .A2(keyinput_122), .B1(n16044), .B2(
        keyinput_123), .ZN(n13721) );
  AOI221_X1 U15339 ( .B1(n13722), .B2(keyinput_122), .C1(keyinput_123), .C2(
        n16044), .A(n13721), .ZN(n13723) );
  OAI21_X1 U15340 ( .B1(n13725), .B2(n13724), .A(n13723), .ZN(n13726) );
  AOI22_X1 U15341 ( .A1(n13727), .A2(n13726), .B1(keyinput_126), .B2(
        P3_REG3_REG_26__SCAN_IN), .ZN(n13728) );
  OAI21_X1 U15342 ( .B1(keyinput_126), .B2(P3_REG3_REG_26__SCAN_IN), .A(n13728), .ZN(n13730) );
  AOI21_X1 U15343 ( .B1(keyinput_127), .B2(n13730), .A(keyinput_63), .ZN(
        n13732) );
  INV_X1 U15344 ( .A(keyinput_127), .ZN(n13729) );
  AOI21_X1 U15345 ( .B1(n13730), .B2(n13729), .A(P3_REG3_REG_15__SCAN_IN), 
        .ZN(n13731) );
  AOI22_X1 U15346 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(n13732), .B1(keyinput_63), .B2(n13731), .ZN(n13733) );
  AOI221_X1 U15347 ( .B1(keyinput_62), .B2(n13735), .C1(n13734), .C2(n13735), 
        .A(n13733), .ZN(n13736) );
  XOR2_X1 U15348 ( .A(n13737), .B(n13736), .Z(P3_U3493) );
  MUX2_X1 U15349 ( .A(n13738), .B(P3_DATAO_REG_1__SCAN_IN), .S(n13739), .Z(
        P3_U3492) );
  MUX2_X1 U15350 ( .A(n13740), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13739), .Z(
        P3_U3491) );
  NOR3_X1 U15351 ( .A1(n7357), .A2(n7406), .A3(n13742), .ZN(n13744) );
  OAI21_X1 U15352 ( .B1(n13744), .B2(n13743), .A(n13897), .ZN(n13761) );
  OR3_X1 U15353 ( .A1(n13747), .A2(n13746), .A3(n13745), .ZN(n13748) );
  AOI21_X1 U15354 ( .B1(n13749), .B2(n13748), .A(n13895), .ZN(n13750) );
  AOI211_X1 U15355 ( .C1(n15817), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n13751), .B(
        n13750), .ZN(n13760) );
  NAND2_X1 U15356 ( .A1(n13874), .A2(n13752), .ZN(n13759) );
  AND3_X1 U15357 ( .A1(n13755), .A2(n13754), .A3(n13753), .ZN(n13756) );
  OAI21_X1 U15358 ( .B1(n13757), .B2(n13756), .A(n13865), .ZN(n13758) );
  NAND4_X1 U15359 ( .A1(n13761), .A2(n13760), .A3(n13759), .A4(n13758), .ZN(
        P3_U3186) );
  INV_X1 U15360 ( .A(n13762), .ZN(n13764) );
  NOR3_X1 U15361 ( .A1(n13765), .A2(n13764), .A3(n13763), .ZN(n13768) );
  INV_X1 U15362 ( .A(n13766), .ZN(n13767) );
  OAI21_X1 U15363 ( .B1(n13768), .B2(n13767), .A(n13897), .ZN(n13787) );
  NOR2_X1 U15364 ( .A1(n13889), .A2(n13769), .ZN(n13770) );
  AOI211_X1 U15365 ( .C1(n15817), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n13771), .B(
        n13770), .ZN(n13786) );
  INV_X1 U15366 ( .A(n13772), .ZN(n13773) );
  NOR3_X1 U15367 ( .A1(n13775), .A2(n13774), .A3(n13773), .ZN(n13777) );
  OAI21_X1 U15368 ( .B1(n13777), .B2(n13776), .A(n13838), .ZN(n13785) );
  INV_X1 U15369 ( .A(n13778), .ZN(n13781) );
  NOR3_X1 U15370 ( .A1(n13781), .A2(n7958), .A3(n13780), .ZN(n13782) );
  OAI21_X1 U15371 ( .B1(n13783), .B2(n13782), .A(n13865), .ZN(n13784) );
  NAND4_X1 U15372 ( .A1(n13787), .A2(n13786), .A3(n13785), .A4(n13784), .ZN(
        P3_U3188) );
  AOI21_X1 U15373 ( .B1(n14185), .B2(n13790), .A(n13810), .ZN(n13808) );
  AOI21_X1 U15374 ( .B1(n14096), .B2(n13793), .A(n13821), .ZN(n13796) );
  AOI21_X1 U15375 ( .B1(n15817), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13794), 
        .ZN(n13795) );
  OAI21_X1 U15376 ( .B1(n13895), .B2(n13796), .A(n13795), .ZN(n13806) );
  MUX2_X1 U15377 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13309), .Z(n13803) );
  NAND2_X1 U15378 ( .A1(n13798), .A2(n13797), .ZN(n13799) );
  NAND2_X1 U15379 ( .A1(n13800), .A2(n13799), .ZN(n13815) );
  XNOR2_X1 U15380 ( .A(n13815), .B(n13801), .ZN(n13802) );
  NOR2_X1 U15381 ( .A1(n13802), .A2(n13803), .ZN(n13816) );
  AOI21_X1 U15382 ( .B1(n13803), .B2(n13802), .A(n13816), .ZN(n13804) );
  NOR2_X1 U15383 ( .A1(n13804), .A2(n13877), .ZN(n13805) );
  AOI211_X1 U15384 ( .C1(n13874), .C2(n7449), .A(n13806), .B(n13805), .ZN(
        n13807) );
  OAI21_X1 U15385 ( .B1(n13808), .B2(n13899), .A(n13807), .ZN(P3_U3197) );
  NOR2_X1 U15386 ( .A1(n7449), .A2(n13809), .ZN(n13811) );
  AOI22_X1 U15387 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13823), .B1(n13844), 
        .B2(n13812), .ZN(n13813) );
  AOI21_X1 U15388 ( .B1(n13814), .B2(n13813), .A(n13832), .ZN(n13831) );
  INV_X1 U15389 ( .A(n13815), .ZN(n13817) );
  AOI21_X1 U15390 ( .B1(n13817), .B2(n7449), .A(n13816), .ZN(n13847) );
  MUX2_X1 U15391 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13309), .Z(n13845) );
  XNOR2_X1 U15392 ( .A(n13845), .B(n13844), .ZN(n13846) );
  XNOR2_X1 U15393 ( .A(n13847), .B(n13846), .ZN(n13829) );
  NAND2_X1 U15394 ( .A1(n15817), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n13818) );
  OAI211_X1 U15395 ( .C1(n13889), .C2(n13844), .A(n13819), .B(n13818), .ZN(
        n13828) );
  AOI22_X1 U15396 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13823), .B1(n13844), 
        .B2(n13822), .ZN(n13824) );
  AOI21_X1 U15397 ( .B1(n13825), .B2(n13824), .A(n13835), .ZN(n13826) );
  NOR2_X1 U15398 ( .A1(n13826), .A2(n13895), .ZN(n13827) );
  AOI211_X1 U15399 ( .C1(n13897), .C2(n13829), .A(n13828), .B(n13827), .ZN(
        n13830) );
  OAI21_X1 U15400 ( .B1(n13831), .B2(n13899), .A(n13830), .ZN(P3_U3198) );
  AOI21_X1 U15401 ( .B1(n13834), .B2(n13833), .A(n13858), .ZN(n13853) );
  INV_X1 U15402 ( .A(n13836), .ZN(n13837) );
  NOR2_X1 U15403 ( .A1(P3_REG2_REG_17__SCAN_IN), .A2(n13837), .ZN(n13839) );
  OAI21_X1 U15404 ( .B1(n13867), .B2(n13839), .A(n13838), .ZN(n13841) );
  OAI211_X1 U15405 ( .C1(n13843), .C2(n13842), .A(n13841), .B(n13840), .ZN(
        n13851) );
  MUX2_X1 U15406 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13309), .Z(n13855) );
  XNOR2_X1 U15407 ( .A(n13855), .B(n13868), .ZN(n13849) );
  OAI22_X1 U15408 ( .A1(n13847), .A2(n13846), .B1(n13845), .B2(n13844), .ZN(
        n13848) );
  NOR2_X1 U15409 ( .A1(n13848), .A2(n13849), .ZN(n13854) );
  AOI211_X1 U15410 ( .C1(n13849), .C2(n13848), .A(n13877), .B(n13854), .ZN(
        n13850) );
  AOI211_X1 U15411 ( .C1(n13874), .C2(n8166), .A(n13851), .B(n13850), .ZN(
        n13852) );
  OAI21_X1 U15412 ( .B1(n13853), .B2(n13899), .A(n13852), .ZN(P3_U3199) );
  MUX2_X1 U15413 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13309), .Z(n13857) );
  AOI21_X1 U15414 ( .B1(n13855), .B2(n13868), .A(n13854), .ZN(n13885) );
  XNOR2_X1 U15415 ( .A(n13885), .B(n13884), .ZN(n13856) );
  NOR2_X1 U15416 ( .A1(n13856), .A2(n13857), .ZN(n13883) );
  AOI21_X1 U15417 ( .B1(n13857), .B2(n13856), .A(n13883), .ZN(n13878) );
  INV_X1 U15418 ( .A(n13858), .ZN(n13864) );
  OR2_X1 U15419 ( .A1(n13884), .A2(n13860), .ZN(n13879) );
  NAND2_X1 U15420 ( .A1(n13884), .A2(n13860), .ZN(n13861) );
  NAND2_X1 U15421 ( .A1(n13879), .A2(n13861), .ZN(n13862) );
  AND3_X1 U15422 ( .A1(n13864), .A2(n13863), .A3(n13862), .ZN(n13866) );
  OAI21_X1 U15423 ( .B1(n13880), .B2(n13866), .A(n13865), .ZN(n13876) );
  OR2_X1 U15424 ( .A1(n13884), .A2(n14045), .ZN(n13890) );
  NAND2_X1 U15425 ( .A1(n13884), .A2(n14045), .ZN(n13869) );
  NAND2_X1 U15426 ( .A1(n13890), .A2(n13869), .ZN(n13870) );
  NAND2_X1 U15427 ( .A1(n15817), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13872) );
  OAI211_X1 U15428 ( .C1(n13878), .C2(n13877), .A(n13876), .B(n13875), .ZN(
        P3_U3200) );
  XNOR2_X1 U15429 ( .A(n13881), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13882) );
  XNOR2_X1 U15430 ( .A(n13881), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13892) );
  MUX2_X1 U15431 ( .A(n13892), .B(n13882), .S(n13309), .Z(n13887) );
  AOI21_X1 U15432 ( .B1(n13885), .B2(n13884), .A(n13883), .ZN(n13886) );
  XOR2_X1 U15433 ( .A(n13887), .B(n13886), .Z(n13898) );
  NOR2_X1 U15434 ( .A1(n13889), .A2(n13888), .ZN(n13896) );
  INV_X1 U15435 ( .A(n13890), .ZN(n13891) );
  NAND2_X1 U15436 ( .A1(n15817), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13894) );
  INV_X1 U15437 ( .A(n14119), .ZN(n14195) );
  INV_X1 U15438 ( .A(n13900), .ZN(n13901) );
  NOR2_X1 U15439 ( .A1(n13903), .A2(n16128), .ZN(n13910) );
  NOR3_X1 U15440 ( .A1(n14193), .A2(n16052), .A3(n13910), .ZN(n13906) );
  NOR2_X1 U15441 ( .A1(n16131), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13904) );
  OAI22_X1 U15442 ( .A1(n14195), .A2(n16126), .B1(n13906), .B2(n13904), .ZN(
        P3_U3202) );
  NOR2_X1 U15443 ( .A1(n16131), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13905) );
  OAI22_X1 U15444 ( .A1(n14124), .A2(n16126), .B1(n13906), .B2(n13905), .ZN(
        P3_U3203) );
  NAND2_X1 U15445 ( .A1(n13907), .A2(n16131), .ZN(n13912) );
  NOR2_X1 U15446 ( .A1(n13908), .A2(n16126), .ZN(n13909) );
  AOI211_X1 U15447 ( .C1(n16052), .C2(P3_REG2_REG_29__SCAN_IN), .A(n13910), 
        .B(n13909), .ZN(n13911) );
  OAI211_X1 U15448 ( .C1(n13913), .C2(n14118), .A(n13912), .B(n13911), .ZN(
        P3_U3204) );
  INV_X1 U15449 ( .A(n14126), .ZN(n13927) );
  OR2_X1 U15450 ( .A1(n13916), .A2(n13915), .ZN(n13917) );
  NAND3_X1 U15451 ( .A1(n13918), .A2(n14103), .A3(n13917), .ZN(n13922) );
  NOR2_X1 U15452 ( .A1(n13919), .A2(n16032), .ZN(n13920) );
  AOI22_X1 U15453 ( .A1(n13923), .A2(n14079), .B1(n16052), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13924) );
  OAI21_X1 U15454 ( .B1(n14203), .B2(n16126), .A(n13924), .ZN(n13925) );
  AOI21_X1 U15455 ( .B1(n14125), .B2(n16131), .A(n13925), .ZN(n13926) );
  OAI21_X1 U15456 ( .B1(n13927), .B2(n14118), .A(n13926), .ZN(P3_U3205) );
  XNOR2_X1 U15457 ( .A(n13928), .B(n13930), .ZN(n14130) );
  INV_X1 U15458 ( .A(n14130), .ZN(n13937) );
  OAI222_X1 U15459 ( .A1(n16032), .A2(n13932), .B1(n16034), .B2(n13953), .C1(
        n16039), .C2(n13931), .ZN(n14129) );
  AOI22_X1 U15460 ( .A1(n13933), .A2(n14079), .B1(n16052), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13934) );
  OAI21_X1 U15461 ( .B1(n8012), .B2(n16126), .A(n13934), .ZN(n13935) );
  AOI21_X1 U15462 ( .B1(n14129), .B2(n16131), .A(n13935), .ZN(n13936) );
  OAI21_X1 U15463 ( .B1(n13937), .B2(n14118), .A(n13936), .ZN(P3_U3206) );
  XNOR2_X1 U15464 ( .A(n13939), .B(n13938), .ZN(n14134) );
  INV_X1 U15465 ( .A(n14134), .ZN(n13948) );
  XNOR2_X1 U15466 ( .A(n13941), .B(n13940), .ZN(n13942) );
  OAI222_X1 U15467 ( .A1(n16032), .A2(n13943), .B1(n16034), .B2(n13965), .C1(
        n13942), .C2(n16039), .ZN(n14133) );
  AOI22_X1 U15468 ( .A1(n13944), .A2(n14079), .B1(n16052), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13945) );
  OAI21_X1 U15469 ( .B1(n14210), .B2(n16126), .A(n13945), .ZN(n13946) );
  AOI21_X1 U15470 ( .B1(n14133), .B2(n16131), .A(n13946), .ZN(n13947) );
  OAI21_X1 U15471 ( .B1(n13948), .B2(n14118), .A(n13947), .ZN(P3_U3207) );
  XNOR2_X1 U15472 ( .A(n13949), .B(n13952), .ZN(n14138) );
  INV_X1 U15473 ( .A(n14138), .ZN(n13960) );
  AOI211_X1 U15474 ( .C1(n13952), .C2(n13950), .A(n16039), .B(n13951), .ZN(
        n13955) );
  OAI22_X1 U15475 ( .A1(n13953), .A2(n16032), .B1(n13978), .B2(n16034), .ZN(
        n13954) );
  OR2_X1 U15476 ( .A1(n13955), .A2(n13954), .ZN(n14137) );
  AOI22_X1 U15477 ( .A1(n13956), .A2(n14079), .B1(n16052), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13957) );
  OAI21_X1 U15478 ( .B1(n14214), .B2(n16126), .A(n13957), .ZN(n13958) );
  AOI21_X1 U15479 ( .B1(n14137), .B2(n16131), .A(n13958), .ZN(n13959) );
  OAI21_X1 U15480 ( .B1(n14118), .B2(n13960), .A(n13959), .ZN(P3_U3208) );
  OR2_X1 U15481 ( .A1(n13962), .A2(n13961), .ZN(n13969) );
  XOR2_X1 U15482 ( .A(n13969), .B(n13963), .Z(n13964) );
  OAI222_X1 U15483 ( .A1(n16034), .A2(n13966), .B1(n16032), .B2(n13965), .C1(
        n13964), .C2(n16039), .ZN(n14141) );
  AOI21_X1 U15484 ( .B1(n14079), .B2(n13967), .A(n14141), .ZN(n13973) );
  AOI22_X1 U15485 ( .A1(n13968), .A2(n14065), .B1(P3_REG2_REG_24__SCAN_IN), 
        .B2(n16052), .ZN(n13972) );
  XNOR2_X1 U15486 ( .A(n13970), .B(n13969), .ZN(n14142) );
  NAND2_X1 U15487 ( .A1(n14142), .A2(n14099), .ZN(n13971) );
  OAI211_X1 U15488 ( .C1(n13973), .C2(n16052), .A(n13972), .B(n13971), .ZN(
        P3_U3209) );
  XNOR2_X1 U15489 ( .A(n13975), .B(n13974), .ZN(n13976) );
  OAI222_X1 U15490 ( .A1(n16032), .A2(n13978), .B1(n16034), .B2(n13977), .C1(
        n16039), .C2(n13976), .ZN(n14146) );
  NOR2_X1 U15491 ( .A1(n13980), .A2(n13979), .ZN(n14145) );
  INV_X1 U15492 ( .A(n14147), .ZN(n13981) );
  NOR3_X1 U15493 ( .A1(n14145), .A2(n13981), .A3(n14118), .ZN(n13985) );
  AOI22_X1 U15494 ( .A1(n13982), .A2(n14079), .B1(n16052), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13983) );
  OAI21_X1 U15495 ( .B1(n14222), .B2(n16126), .A(n13983), .ZN(n13984) );
  AOI211_X1 U15496 ( .C1(n14146), .C2(n16131), .A(n13985), .B(n13984), .ZN(
        n13986) );
  INV_X1 U15497 ( .A(n13986), .ZN(P3_U3210) );
  XNOR2_X1 U15498 ( .A(n13987), .B(n8028), .ZN(n13989) );
  AOI222_X1 U15499 ( .A1(n14103), .A2(n13989), .B1(n14015), .B2(n14108), .C1(
        n13988), .C2(n14107), .ZN(n14153) );
  NAND2_X1 U15500 ( .A1(n13991), .A2(n13990), .ZN(n13992) );
  NAND2_X1 U15501 ( .A1(n13993), .A2(n13992), .ZN(n14154) );
  AOI22_X1 U15502 ( .A1(n13994), .A2(n14079), .B1(n16052), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n13996) );
  NAND2_X1 U15503 ( .A1(n14151), .A2(n14065), .ZN(n13995) );
  OAI211_X1 U15504 ( .C1(n14154), .C2(n14118), .A(n13996), .B(n13995), .ZN(
        n13997) );
  INV_X1 U15505 ( .A(n13997), .ZN(n13998) );
  OAI21_X1 U15506 ( .B1(n14153), .B2(n16052), .A(n13998), .ZN(P3_U3211) );
  XNOR2_X1 U15507 ( .A(n14000), .B(n13999), .ZN(n14003) );
  AOI222_X1 U15508 ( .A1(n14103), .A2(n14003), .B1(n14002), .B2(n14107), .C1(
        n14001), .C2(n14108), .ZN(n14158) );
  OAI21_X1 U15509 ( .B1(n8463), .B2(n9813), .A(n14004), .ZN(n14156) );
  AOI22_X1 U15510 ( .A1(n14005), .A2(n14079), .B1(n16052), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n14006) );
  OAI21_X1 U15511 ( .B1(n14007), .B2(n16126), .A(n14006), .ZN(n14008) );
  AOI21_X1 U15512 ( .B1(n14156), .B2(n14099), .A(n14008), .ZN(n14009) );
  OAI21_X1 U15513 ( .B1(n14158), .B2(n16052), .A(n14009), .ZN(P3_U3212) );
  XNOR2_X1 U15514 ( .A(n14010), .B(n14011), .ZN(n14019) );
  OR2_X1 U15515 ( .A1(n14012), .A2(n14011), .ZN(n14013) );
  NAND2_X1 U15516 ( .A1(n14014), .A2(n14013), .ZN(n14159) );
  AOI22_X1 U15517 ( .A1(n14015), .A2(n14107), .B1(n14108), .B2(n14050), .ZN(
        n14016) );
  OAI21_X1 U15518 ( .B1(n14159), .B2(n14017), .A(n14016), .ZN(n14018) );
  AOI21_X1 U15519 ( .B1(n14019), .B2(n14103), .A(n14018), .ZN(n14161) );
  AOI22_X1 U15520 ( .A1(n16052), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n14020), 
        .B2(n14079), .ZN(n14022) );
  NAND2_X1 U15521 ( .A1(n14227), .A2(n14065), .ZN(n14021) );
  OAI211_X1 U15522 ( .C1(n14159), .C2(n14023), .A(n14022), .B(n14021), .ZN(
        n14024) );
  INV_X1 U15523 ( .A(n14024), .ZN(n14025) );
  OAI21_X1 U15524 ( .B1(n14161), .B2(n16052), .A(n14025), .ZN(P3_U3213) );
  XOR2_X1 U15525 ( .A(n14034), .B(n14026), .Z(n14027) );
  OAI222_X1 U15526 ( .A1(n16032), .A2(n14029), .B1(n16034), .B2(n14028), .C1(
        n16039), .C2(n14027), .ZN(n14165) );
  INV_X1 U15527 ( .A(n14165), .ZN(n14041) );
  INV_X1 U15528 ( .A(n14030), .ZN(n14032) );
  OAI22_X1 U15529 ( .A1(n14032), .A2(n16128), .B1(n16131), .B2(n14031), .ZN(
        n14038) );
  INV_X1 U15530 ( .A(n14033), .ZN(n14036) );
  AND2_X1 U15531 ( .A1(n14035), .A2(n14034), .ZN(n14164) );
  NOR3_X1 U15532 ( .A1(n14036), .A2(n14164), .A3(n14118), .ZN(n14037) );
  AOI211_X1 U15533 ( .C1(n14065), .C2(n14039), .A(n14038), .B(n14037), .ZN(
        n14040) );
  OAI21_X1 U15534 ( .B1(n14041), .B2(n16052), .A(n14040), .ZN(P3_U3214) );
  XNOR2_X1 U15535 ( .A(n14042), .B(n14047), .ZN(n14172) );
  INV_X1 U15536 ( .A(n14043), .ZN(n14044) );
  OAI22_X1 U15537 ( .A1(n16131), .A2(n14045), .B1(n14044), .B2(n16128), .ZN(
        n14053) );
  OAI21_X1 U15538 ( .B1(n14048), .B2(n14047), .A(n14046), .ZN(n14051) );
  AOI222_X1 U15539 ( .A1(n14103), .A2(n14051), .B1(n14050), .B2(n14107), .C1(
        n14049), .C2(n14108), .ZN(n14171) );
  NOR2_X1 U15540 ( .A1(n14171), .A2(n16052), .ZN(n14052) );
  AOI211_X1 U15541 ( .C1(n14065), .C2(n14169), .A(n14053), .B(n14052), .ZN(
        n14054) );
  OAI21_X1 U15542 ( .B1(n14118), .B2(n14172), .A(n14054), .ZN(P3_U3215) );
  OAI211_X1 U15543 ( .C1(n14057), .C2(n14056), .A(n14055), .B(n14103), .ZN(
        n14060) );
  AOI22_X1 U15544 ( .A1(n14058), .A2(n14107), .B1(n14108), .B2(n14088), .ZN(
        n14059) );
  AND2_X1 U15545 ( .A1(n14060), .A2(n14059), .ZN(n14175) );
  INV_X1 U15546 ( .A(n14237), .ZN(n14066) );
  INV_X1 U15547 ( .A(n14061), .ZN(n14062) );
  OAI22_X1 U15548 ( .A1(n16131), .A2(n14063), .B1(n14062), .B2(n16128), .ZN(
        n14064) );
  AOI21_X1 U15549 ( .B1(n14066), .B2(n14065), .A(n14064), .ZN(n14070) );
  XNOR2_X1 U15550 ( .A(n14067), .B(n14068), .ZN(n14173) );
  NAND2_X1 U15551 ( .A1(n14173), .A2(n14099), .ZN(n14069) );
  OAI211_X1 U15552 ( .C1(n14175), .C2(n16052), .A(n14070), .B(n14069), .ZN(
        P3_U3216) );
  XOR2_X1 U15553 ( .A(n14074), .B(n14071), .Z(n14181) );
  AOI21_X1 U15554 ( .B1(n14074), .B2(n14073), .A(n14072), .ZN(n14075) );
  OAI222_X1 U15555 ( .A1(n16032), .A2(n14077), .B1(n16034), .B2(n14076), .C1(
        n16039), .C2(n14075), .ZN(n14178) );
  AOI22_X1 U15556 ( .A1(n16052), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n14079), 
        .B2(n14078), .ZN(n14080) );
  OAI21_X1 U15557 ( .B1(n14081), .B2(n16126), .A(n14080), .ZN(n14082) );
  AOI21_X1 U15558 ( .B1(n14178), .B2(n16131), .A(n14082), .ZN(n14083) );
  OAI21_X1 U15559 ( .B1(n14181), .B2(n14118), .A(n14083), .ZN(P3_U3217) );
  NAND3_X1 U15560 ( .A1(n14085), .A2(n14093), .A3(n14086), .ZN(n14087) );
  NAND3_X1 U15561 ( .A1(n14084), .A2(n14103), .A3(n14087), .ZN(n14091) );
  AOI22_X1 U15562 ( .A1(n14108), .A2(n14089), .B1(n14088), .B2(n14107), .ZN(
        n14090) );
  NAND2_X1 U15563 ( .A1(n14091), .A2(n14090), .ZN(n14183) );
  INV_X1 U15564 ( .A(n14183), .ZN(n14101) );
  OAI21_X1 U15565 ( .B1(n14094), .B2(n14093), .A(n14092), .ZN(n14184) );
  NOR2_X1 U15566 ( .A1(n14242), .A2(n16126), .ZN(n14098) );
  OAI22_X1 U15567 ( .A1(n16131), .A2(n14096), .B1(n14095), .B2(n16128), .ZN(
        n14097) );
  AOI211_X1 U15568 ( .C1(n14184), .C2(n14099), .A(n14098), .B(n14097), .ZN(
        n14100) );
  OAI21_X1 U15569 ( .B1(n14101), .B2(n16052), .A(n14100), .ZN(P3_U3218) );
  XNOR2_X1 U15570 ( .A(n14102), .B(n8426), .ZN(n16227) );
  INV_X1 U15571 ( .A(n16227), .ZN(n14117) );
  OAI211_X1 U15572 ( .C1(n14105), .C2(n14104), .A(n14085), .B(n14103), .ZN(
        n14111) );
  AOI22_X1 U15573 ( .A1(n14109), .A2(n14108), .B1(n14107), .B2(n14106), .ZN(
        n14110) );
  NAND2_X1 U15574 ( .A1(n14111), .A2(n14110), .ZN(n16224) );
  NOR2_X1 U15575 ( .A1(n16223), .A2(n16126), .ZN(n14115) );
  OAI22_X1 U15576 ( .A1(n16131), .A2(n14113), .B1(n14112), .B2(n16128), .ZN(
        n14114) );
  AOI211_X1 U15577 ( .C1(n16224), .C2(n16131), .A(n14115), .B(n14114), .ZN(
        n14116) );
  OAI21_X1 U15578 ( .B1(n14118), .B2(n14117), .A(n14116), .ZN(P3_U3219) );
  NAND2_X1 U15579 ( .A1(n14119), .A2(n9879), .ZN(n14120) );
  NAND2_X1 U15580 ( .A1(n14193), .A2(n16228), .ZN(n14123) );
  OAI211_X1 U15581 ( .C1(n16228), .C2(n14121), .A(n14120), .B(n14123), .ZN(
        P3_U3490) );
  NAND2_X1 U15582 ( .A1(n7687), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n14122) );
  OAI211_X1 U15583 ( .C1(n14124), .C2(n14192), .A(n14123), .B(n14122), .ZN(
        P3_U3489) );
  INV_X1 U15584 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n14127) );
  MUX2_X1 U15585 ( .A(n14127), .B(n14200), .S(n16228), .Z(n14128) );
  OAI21_X1 U15586 ( .B1(n14203), .B2(n14192), .A(n14128), .ZN(P3_U3487) );
  INV_X1 U15587 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n14131) );
  AOI21_X1 U15588 ( .B1(n16226), .B2(n14130), .A(n14129), .ZN(n14204) );
  OAI21_X1 U15589 ( .B1(n8012), .B2(n14192), .A(n14132), .ZN(P3_U3486) );
  INV_X1 U15590 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n14135) );
  AOI21_X1 U15591 ( .B1(n16226), .B2(n14134), .A(n14133), .ZN(n14207) );
  MUX2_X1 U15592 ( .A(n14135), .B(n14207), .S(n16228), .Z(n14136) );
  OAI21_X1 U15593 ( .B1(n14210), .B2(n14192), .A(n14136), .ZN(P3_U3485) );
  INV_X1 U15594 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n14139) );
  AOI21_X1 U15595 ( .B1(n14138), .B2(n16226), .A(n14137), .ZN(n14211) );
  MUX2_X1 U15596 ( .A(n14139), .B(n14211), .S(n16228), .Z(n14140) );
  OAI21_X1 U15597 ( .B1(n14214), .B2(n14192), .A(n14140), .ZN(P3_U3484) );
  INV_X1 U15598 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n14143) );
  AOI21_X1 U15599 ( .B1(n16226), .B2(n14142), .A(n14141), .ZN(n14215) );
  MUX2_X1 U15600 ( .A(n14143), .B(n14215), .S(n16228), .Z(n14144) );
  OAI21_X1 U15601 ( .B1(n14218), .B2(n14192), .A(n14144), .ZN(P3_U3483) );
  INV_X1 U15602 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n14149) );
  NOR2_X1 U15603 ( .A1(n14145), .A2(n14182), .ZN(n14148) );
  AOI21_X1 U15604 ( .B1(n14148), .B2(n14147), .A(n14146), .ZN(n14219) );
  MUX2_X1 U15605 ( .A(n14149), .B(n14219), .S(n16228), .Z(n14150) );
  OAI21_X1 U15606 ( .B1(n14222), .B2(n14192), .A(n14150), .ZN(P3_U3482) );
  NAND2_X1 U15607 ( .A1(n14151), .A2(n16054), .ZN(n14152) );
  OAI211_X1 U15608 ( .C1(n14182), .C2(n14154), .A(n14153), .B(n14152), .ZN(
        n14223) );
  MUX2_X1 U15609 ( .A(P3_REG1_REG_22__SCAN_IN), .B(n14223), .S(n16228), .Z(
        P3_U3481) );
  AOI22_X1 U15610 ( .A1(n14156), .A2(n16226), .B1(n16054), .B2(n14155), .ZN(
        n14157) );
  NAND2_X1 U15611 ( .A1(n14158), .A2(n14157), .ZN(n14224) );
  MUX2_X1 U15612 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n14224), .S(n16228), .Z(
        P3_U3480) );
  OR2_X1 U15613 ( .A1(n14159), .A2(n16163), .ZN(n14160) );
  NAND2_X1 U15614 ( .A1(n14161), .A2(n14160), .ZN(n14225) );
  MUX2_X1 U15615 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n14225), .S(n16228), .Z(
        n14162) );
  AOI21_X1 U15616 ( .B1(n9879), .B2(n14227), .A(n14162), .ZN(n14163) );
  INV_X1 U15617 ( .A(n14163), .ZN(P3_U3479) );
  INV_X1 U15618 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n14167) );
  NOR2_X1 U15619 ( .A1(n14164), .A2(n14182), .ZN(n14166) );
  AOI21_X1 U15620 ( .B1(n14166), .B2(n14033), .A(n14165), .ZN(n14229) );
  MUX2_X1 U15621 ( .A(n14167), .B(n14229), .S(n16228), .Z(n14168) );
  OAI21_X1 U15622 ( .B1(n14232), .B2(n14192), .A(n14168), .ZN(P3_U3478) );
  NAND2_X1 U15623 ( .A1(n14169), .A2(n16054), .ZN(n14170) );
  OAI211_X1 U15624 ( .C1(n14182), .C2(n14172), .A(n14171), .B(n14170), .ZN(
        n14233) );
  MUX2_X1 U15625 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n14233), .S(n16228), .Z(
        P3_U3477) );
  NAND2_X1 U15626 ( .A1(n14173), .A2(n16226), .ZN(n14174) );
  NAND2_X1 U15627 ( .A1(n14175), .A2(n14174), .ZN(n14234) );
  MUX2_X1 U15628 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n14234), .S(n16228), .Z(
        n14176) );
  INV_X1 U15629 ( .A(n14176), .ZN(n14177) );
  OAI21_X1 U15630 ( .B1(n14192), .B2(n14237), .A(n14177), .ZN(P3_U3476) );
  AOI21_X1 U15631 ( .B1(n16054), .B2(n14179), .A(n14178), .ZN(n14180) );
  OAI21_X1 U15632 ( .B1(n14182), .B2(n14181), .A(n14180), .ZN(n14238) );
  MUX2_X1 U15633 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n14238), .S(n16228), .Z(
        P3_U3475) );
  AOI21_X1 U15634 ( .B1(n16226), .B2(n14184), .A(n14183), .ZN(n14239) );
  MUX2_X1 U15635 ( .A(n14185), .B(n14239), .S(n16228), .Z(n14186) );
  OAI21_X1 U15636 ( .B1(n14192), .B2(n14242), .A(n14186), .ZN(P3_U3474) );
  INV_X1 U15637 ( .A(n14187), .ZN(n14247) );
  INV_X1 U15638 ( .A(n16163), .ZN(n16213) );
  AOI21_X1 U15639 ( .B1(n16213), .B2(n14189), .A(n14188), .ZN(n14243) );
  MUX2_X1 U15640 ( .A(n14190), .B(n14243), .S(n16228), .Z(n14191) );
  OAI21_X1 U15641 ( .B1(n14247), .B2(n14192), .A(n14191), .ZN(P3_U3471) );
  NAND2_X1 U15642 ( .A1(n16229), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n14194) );
  NAND2_X1 U15643 ( .A1(n14193), .A2(n16232), .ZN(n14197) );
  OAI211_X1 U15644 ( .C1(n14195), .C2(n14246), .A(n14194), .B(n14197), .ZN(
        P3_U3458) );
  NAND2_X1 U15645 ( .A1(n14196), .A2(n9862), .ZN(n14198) );
  OAI211_X1 U15646 ( .C1(n16232), .C2(n14199), .A(n14198), .B(n14197), .ZN(
        P3_U3457) );
  MUX2_X1 U15647 ( .A(n14201), .B(n14200), .S(n16232), .Z(n14202) );
  OAI21_X1 U15648 ( .B1(n14203), .B2(n14246), .A(n14202), .ZN(P3_U3455) );
  OAI21_X1 U15649 ( .B1(n8012), .B2(n14246), .A(n14206), .ZN(P3_U3454) );
  MUX2_X1 U15650 ( .A(n14208), .B(n14207), .S(n16232), .Z(n14209) );
  OAI21_X1 U15651 ( .B1(n14210), .B2(n14246), .A(n14209), .ZN(P3_U3453) );
  MUX2_X1 U15652 ( .A(n14212), .B(n14211), .S(n16232), .Z(n14213) );
  OAI21_X1 U15653 ( .B1(n14214), .B2(n14246), .A(n14213), .ZN(P3_U3452) );
  MUX2_X1 U15654 ( .A(n14216), .B(n14215), .S(n16232), .Z(n14217) );
  OAI21_X1 U15655 ( .B1(n14218), .B2(n14246), .A(n14217), .ZN(P3_U3451) );
  MUX2_X1 U15656 ( .A(n14220), .B(n14219), .S(n16232), .Z(n14221) );
  OAI21_X1 U15657 ( .B1(n14222), .B2(n14246), .A(n14221), .ZN(P3_U3450) );
  MUX2_X1 U15658 ( .A(P3_REG0_REG_22__SCAN_IN), .B(n14223), .S(n16232), .Z(
        P3_U3449) );
  MUX2_X1 U15659 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n14224), .S(n16232), .Z(
        P3_U3448) );
  MUX2_X1 U15660 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n14225), .S(n16232), .Z(
        n14226) );
  AOI21_X1 U15661 ( .B1(n9862), .B2(n14227), .A(n14226), .ZN(n14228) );
  INV_X1 U15662 ( .A(n14228), .ZN(P3_U3447) );
  INV_X1 U15663 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n14230) );
  MUX2_X1 U15664 ( .A(n14230), .B(n14229), .S(n16232), .Z(n14231) );
  OAI21_X1 U15665 ( .B1(n14232), .B2(n14246), .A(n14231), .ZN(P3_U3446) );
  MUX2_X1 U15666 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n14233), .S(n16232), .Z(
        P3_U3444) );
  MUX2_X1 U15667 ( .A(n14234), .B(P3_REG0_REG_17__SCAN_IN), .S(n16229), .Z(
        n14235) );
  INV_X1 U15668 ( .A(n14235), .ZN(n14236) );
  OAI21_X1 U15669 ( .B1(n14246), .B2(n14237), .A(n14236), .ZN(P3_U3441) );
  MUX2_X1 U15670 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n14238), .S(n16232), .Z(
        P3_U3438) );
  INV_X1 U15671 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14240) );
  MUX2_X1 U15672 ( .A(n14240), .B(n14239), .S(n16232), .Z(n14241) );
  OAI21_X1 U15673 ( .B1(n14246), .B2(n14242), .A(n14241), .ZN(P3_U3435) );
  INV_X1 U15674 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14244) );
  MUX2_X1 U15675 ( .A(n14244), .B(n14243), .S(n16232), .Z(n14245) );
  OAI21_X1 U15676 ( .B1(n14247), .B2(n14246), .A(n14245), .ZN(P3_U3426) );
  MUX2_X1 U15677 ( .A(n14248), .B(P3_D_REG_1__SCAN_IN), .S(n14249), .Z(
        P3_U3377) );
  MUX2_X1 U15678 ( .A(n14250), .B(P3_D_REG_0__SCAN_IN), .S(n14249), .Z(
        P3_U3376) );
  NAND3_X1 U15679 ( .A1(n14251), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n14254) );
  OAI22_X1 U15680 ( .A1(n14255), .A2(n14254), .B1(n14253), .B2(n14252), .ZN(
        n14256) );
  AOI21_X1 U15681 ( .B1(n14258), .B2(n14257), .A(n14256), .ZN(n14259) );
  INV_X1 U15682 ( .A(n14259), .ZN(P3_U3264) );
  MUX2_X1 U15683 ( .A(n14260), .B(n7731), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3295) );
  XNOR2_X1 U15684 ( .A(n14777), .B(n14352), .ZN(n14264) );
  NAND2_X1 U15685 ( .A1(n14792), .A2(n14300), .ZN(n14265) );
  XNOR2_X1 U15686 ( .A(n14264), .B(n14265), .ZN(n14326) );
  INV_X1 U15687 ( .A(n14326), .ZN(n14263) );
  NAND2_X1 U15688 ( .A1(n14264), .A2(n14265), .ZN(n14266) );
  XNOR2_X1 U15689 ( .A(n14879), .B(n14304), .ZN(n14269) );
  NOR2_X1 U15690 ( .A1(n14381), .A2(n14267), .ZN(n14268) );
  NAND2_X1 U15691 ( .A1(n14269), .A2(n14268), .ZN(n14270) );
  OAI21_X1 U15692 ( .B1(n14269), .B2(n14268), .A(n14270), .ZN(n14450) );
  NAND2_X1 U15693 ( .A1(n14470), .A2(n14300), .ZN(n14272) );
  XNOR2_X1 U15694 ( .A(n14872), .B(n14352), .ZN(n14271) );
  XOR2_X1 U15695 ( .A(n14272), .B(n14271), .Z(n14378) );
  XNOR2_X1 U15696 ( .A(n14728), .B(n14352), .ZN(n14276) );
  NOR2_X1 U15697 ( .A1(n14433), .A2(n14267), .ZN(n14274) );
  XNOR2_X1 U15698 ( .A(n14276), .B(n14274), .ZN(n14390) );
  INV_X1 U15699 ( .A(n14274), .ZN(n14275) );
  NAND2_X1 U15700 ( .A1(n14276), .A2(n14275), .ZN(n14277) );
  XNOR2_X1 U15701 ( .A(n14713), .B(n14352), .ZN(n14279) );
  AND2_X1 U15702 ( .A1(n14469), .A2(n14350), .ZN(n14278) );
  NAND2_X1 U15703 ( .A1(n14279), .A2(n14278), .ZN(n14280) );
  OAI21_X1 U15704 ( .B1(n14279), .B2(n14278), .A(n14280), .ZN(n14428) );
  NAND2_X1 U15705 ( .A1(n14430), .A2(n14280), .ZN(n14342) );
  XNOR2_X1 U15706 ( .A(n14700), .B(n14304), .ZN(n14282) );
  NAND2_X1 U15707 ( .A1(n14468), .A2(n14300), .ZN(n14281) );
  NOR2_X1 U15708 ( .A1(n14282), .A2(n14281), .ZN(n14283) );
  AOI21_X1 U15709 ( .B1(n14282), .B2(n14281), .A(n14283), .ZN(n14341) );
  INV_X1 U15710 ( .A(n14283), .ZN(n14284) );
  XNOR2_X1 U15711 ( .A(n14929), .B(n14352), .ZN(n14286) );
  NAND2_X1 U15712 ( .A1(n14467), .A2(n14300), .ZN(n14287) );
  XNOR2_X1 U15713 ( .A(n14286), .B(n14287), .ZN(n14413) );
  NAND2_X1 U15714 ( .A1(n14286), .A2(n14287), .ZN(n14288) );
  XNOR2_X1 U15715 ( .A(n14368), .B(n14352), .ZN(n14291) );
  NOR2_X1 U15716 ( .A1(n14289), .A2(n14267), .ZN(n14290) );
  XNOR2_X1 U15717 ( .A(n14291), .B(n14290), .ZN(n14365) );
  XNOR2_X1 U15718 ( .A(n14654), .B(n14352), .ZN(n14292) );
  NOR2_X1 U15719 ( .A1(n14362), .A2(n14267), .ZN(n14422) );
  INV_X1 U15720 ( .A(n14292), .ZN(n14293) );
  NAND2_X1 U15721 ( .A1(n14294), .A2(n14293), .ZN(n14295) );
  XNOR2_X1 U15722 ( .A(n14914), .B(n14352), .ZN(n14296) );
  NOR2_X1 U15723 ( .A1(n14401), .A2(n14267), .ZN(n14334) );
  INV_X1 U15724 ( .A(n14296), .ZN(n14297) );
  NAND2_X1 U15725 ( .A1(n14298), .A2(n14297), .ZN(n14299) );
  XNOR2_X1 U15726 ( .A(n14830), .B(n14304), .ZN(n14302) );
  NAND2_X1 U15727 ( .A1(n14633), .A2(n14300), .ZN(n14301) );
  NOR2_X1 U15728 ( .A1(n14302), .A2(n14301), .ZN(n14303) );
  AOI21_X1 U15729 ( .B1(n14302), .B2(n14301), .A(n14303), .ZN(n14399) );
  XNOR2_X1 U15730 ( .A(n14601), .B(n14304), .ZN(n14306) );
  NAND2_X1 U15731 ( .A1(n14614), .A2(n14300), .ZN(n14305) );
  NOR2_X1 U15732 ( .A1(n14306), .A2(n14305), .ZN(n14307) );
  AOI21_X1 U15733 ( .B1(n14306), .B2(n14305), .A(n14307), .ZN(n14371) );
  INV_X1 U15734 ( .A(n14307), .ZN(n14308) );
  NAND2_X1 U15735 ( .A1(n14370), .A2(n14308), .ZN(n14440) );
  XNOR2_X1 U15736 ( .A(n14584), .B(n14352), .ZN(n14310) );
  NAND2_X1 U15737 ( .A1(n14466), .A2(n14300), .ZN(n14309) );
  XNOR2_X1 U15738 ( .A(n14310), .B(n14309), .ZN(n14439) );
  NAND2_X1 U15739 ( .A1(n14310), .A2(n14309), .ZN(n14311) );
  XNOR2_X1 U15740 ( .A(n14569), .B(n14352), .ZN(n14313) );
  AND2_X1 U15741 ( .A1(n14580), .A2(n14350), .ZN(n14312) );
  NAND2_X1 U15742 ( .A1(n14313), .A2(n14312), .ZN(n14348) );
  OAI21_X1 U15743 ( .B1(n14313), .B2(n14312), .A(n14348), .ZN(n14315) );
  AOI21_X1 U15744 ( .B1(n14314), .B2(n14315), .A(n14449), .ZN(n14316) );
  NAND2_X1 U15745 ( .A1(n14316), .A2(n14349), .ZN(n14322) );
  OAI22_X1 U15746 ( .A1(n14599), .A2(n14402), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14317), .ZN(n14320) );
  OAI22_X1 U15747 ( .A1(n14318), .A2(n14404), .B1(n14567), .B2(n14403), .ZN(
        n14319) );
  AOI211_X1 U15748 ( .C1(n14569), .C2(n14423), .A(n14320), .B(n14319), .ZN(
        n14321) );
  NAND2_X1 U15749 ( .A1(n14322), .A2(n14321), .ZN(P2_U3186) );
  INV_X1 U15750 ( .A(n14324), .ZN(n14325) );
  AOI21_X1 U15751 ( .B1(n14326), .B2(n14323), .A(n14325), .ZN(n14332) );
  INV_X1 U15752 ( .A(n14775), .ZN(n14329) );
  OAI22_X1 U15753 ( .A1(n14327), .A2(n14794), .B1(n14381), .B2(n14600), .ZN(
        n14772) );
  AOI22_X1 U15754 ( .A1(n14392), .A2(n14772), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14328) );
  OAI21_X1 U15755 ( .B1(n14329), .B2(n14403), .A(n14328), .ZN(n14330) );
  AOI21_X1 U15756 ( .B1(n14889), .B2(n14423), .A(n14330), .ZN(n14331) );
  OAI21_X1 U15757 ( .B1(n14332), .B2(n14449), .A(n14331), .ZN(P2_U3187) );
  OAI211_X1 U15758 ( .C1(n14335), .C2(n14334), .A(n14333), .B(n14420), .ZN(
        n14339) );
  NOR2_X1 U15759 ( .A1(n14402), .A2(n14362), .ZN(n14337) );
  OAI22_X1 U15760 ( .A1(n14598), .A2(n14404), .B1(n14403), .B2(n14638), .ZN(
        n14336) );
  AOI211_X1 U15761 ( .C1(P2_REG3_REG_23__SCAN_IN), .C2(P2_U3088), .A(n14337), 
        .B(n14336), .ZN(n14338) );
  OAI211_X1 U15762 ( .C1(n14914), .C2(n14462), .A(n14339), .B(n14338), .ZN(
        P2_U3188) );
  OAI211_X1 U15763 ( .C1(n14342), .C2(n14341), .A(n14340), .B(n14420), .ZN(
        n14347) );
  OAI22_X1 U15764 ( .A1(n14361), .A2(n14600), .B1(n14343), .B2(n14794), .ZN(
        n14690) );
  NOR2_X1 U15765 ( .A1(n14403), .A2(n14698), .ZN(n14344) );
  AOI211_X1 U15766 ( .C1(n14392), .C2(n14690), .A(n14345), .B(n14344), .ZN(
        n14346) );
  OAI211_X1 U15767 ( .C1(n8126), .C2(n14462), .A(n14347), .B(n14346), .ZN(
        P2_U3191) );
  NAND2_X1 U15768 ( .A1(n14349), .A2(n14348), .ZN(n14355) );
  MUX2_X1 U15769 ( .A(n14560), .B(n14351), .S(n14350), .Z(n14353) );
  XNOR2_X1 U15770 ( .A(n14353), .B(n14352), .ZN(n14354) );
  XNOR2_X1 U15771 ( .A(n14355), .B(n14354), .ZN(n14360) );
  AOI22_X1 U15772 ( .A1(n14356), .A2(n14392), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14357) );
  OAI21_X1 U15773 ( .B1(n14558), .B2(n14403), .A(n14357), .ZN(n14358) );
  AOI21_X1 U15774 ( .B1(n14560), .B2(n14423), .A(n14358), .ZN(n14359) );
  OAI21_X1 U15775 ( .B1(n14360), .B2(n14449), .A(n14359), .ZN(P2_U3192) );
  OAI22_X1 U15776 ( .A1(n14362), .A2(n14600), .B1(n14361), .B2(n14794), .ZN(
        n14669) );
  AOI22_X1 U15777 ( .A1(n14669), .A2(n14392), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14363) );
  OAI21_X1 U15778 ( .B1(n14663), .B2(n14403), .A(n14363), .ZN(n14367) );
  AOI211_X1 U15779 ( .C1(n14365), .C2(n14364), .A(n14449), .B(n7264), .ZN(
        n14366) );
  AOI211_X1 U15780 ( .C1(n14368), .C2(n14423), .A(n14367), .B(n14366), .ZN(
        n14369) );
  INV_X1 U15781 ( .A(n14369), .ZN(P2_U3195) );
  OAI211_X1 U15782 ( .C1(n14372), .C2(n14371), .A(n14370), .B(n14420), .ZN(
        n14376) );
  AOI22_X1 U15783 ( .A1(n14443), .A2(n14633), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14375) );
  AOI22_X1 U15784 ( .A1(n14466), .A2(n14444), .B1(n14459), .B2(n14604), .ZN(
        n14374) );
  NAND2_X1 U15785 ( .A1(n14601), .A2(n14423), .ZN(n14373) );
  NAND4_X1 U15786 ( .A1(n14376), .A2(n14375), .A3(n14374), .A4(n14373), .ZN(
        P2_U3197) );
  OAI21_X1 U15787 ( .B1(n14379), .B2(n14378), .A(n14377), .ZN(n14380) );
  NAND2_X1 U15788 ( .A1(n14380), .A2(n14420), .ZN(n14387) );
  INV_X1 U15789 ( .A(n14392), .ZN(n14457) );
  OR2_X1 U15790 ( .A1(n14381), .A2(n14794), .ZN(n14383) );
  OR2_X1 U15791 ( .A1(n14433), .A2(n14600), .ZN(n14382) );
  AND2_X1 U15792 ( .A1(n14383), .A2(n14382), .ZN(n14738) );
  OAI22_X1 U15793 ( .A1(n14457), .A2(n14738), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14384), .ZN(n14385) );
  AOI21_X1 U15794 ( .B1(n14746), .B2(n14459), .A(n14385), .ZN(n14386) );
  OAI211_X1 U15795 ( .C1(n14872), .C2(n14462), .A(n14387), .B(n14386), .ZN(
        P2_U3198) );
  OAI21_X1 U15796 ( .B1(n14390), .B2(n14389), .A(n14388), .ZN(n14396) );
  NAND2_X1 U15797 ( .A1(n14469), .A2(n14791), .ZN(n14391) );
  OAI21_X1 U15798 ( .B1(n14453), .B2(n14794), .A(n14391), .ZN(n14721) );
  AOI22_X1 U15799 ( .A1(n14392), .A2(n14721), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14394) );
  NAND2_X1 U15800 ( .A1(n14459), .A2(n14726), .ZN(n14393) );
  OAI211_X1 U15801 ( .C1(n14728), .C2(n14462), .A(n14394), .B(n14393), .ZN(
        n14395) );
  AOI21_X1 U15802 ( .B1(n14396), .B2(n14420), .A(n14395), .ZN(n14397) );
  INV_X1 U15803 ( .A(n14397), .ZN(P2_U3200) );
  OAI211_X1 U15804 ( .C1(n14400), .C2(n14399), .A(n14398), .B(n14420), .ZN(
        n14409) );
  NOR2_X1 U15805 ( .A1(n14402), .A2(n14401), .ZN(n14407) );
  OAI22_X1 U15806 ( .A1(n14405), .A2(n14404), .B1(n14403), .B2(n14621), .ZN(
        n14406) );
  AOI211_X1 U15807 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3088), .A(n14407), 
        .B(n14406), .ZN(n14408) );
  OAI211_X1 U15808 ( .C1(n14620), .C2(n14462), .A(n14409), .B(n14408), .ZN(
        P2_U3201) );
  INV_X1 U15809 ( .A(n14410), .ZN(n14411) );
  AOI21_X1 U15810 ( .B1(n14413), .B2(n14412), .A(n14411), .ZN(n14418) );
  AOI22_X1 U15811 ( .A1(n14648), .A2(n14791), .B1(n14647), .B2(n14468), .ZN(
        n14683) );
  OAI22_X1 U15812 ( .A1(n14457), .A2(n14683), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14414), .ZN(n14416) );
  NOR2_X1 U15813 ( .A1(n14929), .A2(n14462), .ZN(n14415) );
  AOI211_X1 U15814 ( .C1(n14459), .C2(n14678), .A(n14416), .B(n14415), .ZN(
        n14417) );
  OAI21_X1 U15815 ( .B1(n14418), .B2(n14449), .A(n14417), .ZN(P2_U3205) );
  OAI211_X1 U15816 ( .C1(n14419), .C2(n14422), .A(n14421), .B(n14420), .ZN(
        n14427) );
  AOI22_X1 U15817 ( .A1(n14443), .A2(n14648), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14426) );
  AOI22_X1 U15818 ( .A1(n14444), .A2(n14646), .B1(n14459), .B2(n14652), .ZN(
        n14425) );
  NAND2_X1 U15819 ( .A1(n14840), .A2(n14423), .ZN(n14424) );
  NAND4_X1 U15820 ( .A1(n14427), .A2(n14426), .A3(n14425), .A4(n14424), .ZN(
        P2_U3207) );
  AOI21_X1 U15821 ( .B1(n14429), .B2(n14428), .A(n14449), .ZN(n14431) );
  NAND2_X1 U15822 ( .A1(n14431), .A2(n14430), .ZN(n14438) );
  NAND2_X1 U15823 ( .A1(n14468), .A2(n14791), .ZN(n14432) );
  OAI21_X1 U15824 ( .B1(n14433), .B2(n14794), .A(n14432), .ZN(n14705) );
  INV_X1 U15825 ( .A(n14705), .ZN(n14435) );
  OAI22_X1 U15826 ( .A1(n14457), .A2(n14435), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14434), .ZN(n14436) );
  AOI21_X1 U15827 ( .B1(n14712), .B2(n14459), .A(n14436), .ZN(n14437) );
  OAI211_X1 U15828 ( .C1(n14861), .C2(n14462), .A(n14438), .B(n14437), .ZN(
        P2_U3210) );
  NAND2_X1 U15829 ( .A1(n14440), .A2(n14439), .ZN(n14441) );
  AOI21_X1 U15830 ( .B1(n14442), .B2(n14441), .A(n14449), .ZN(n14448) );
  AOI22_X1 U15831 ( .A1(n14443), .A2(n14614), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14446) );
  AOI22_X1 U15832 ( .A1(n14580), .A2(n14444), .B1(n14459), .B2(n14582), .ZN(
        n14445) );
  OAI211_X1 U15833 ( .C1(n14584), .C2(n14462), .A(n14446), .B(n14445), .ZN(
        n14447) );
  OR2_X1 U15834 ( .A1(n14448), .A2(n14447), .ZN(P2_U3212) );
  AOI21_X1 U15835 ( .B1(n14451), .B2(n14450), .A(n14449), .ZN(n14452) );
  NAND2_X1 U15836 ( .A1(n14452), .A2(n7337), .ZN(n14461) );
  OR2_X1 U15837 ( .A1(n14453), .A2(n14600), .ZN(n14455) );
  NAND2_X1 U15838 ( .A1(n14792), .A2(n14647), .ZN(n14454) );
  AND2_X1 U15839 ( .A1(n14455), .A2(n14454), .ZN(n14761) );
  OAI22_X1 U15840 ( .A1(n14457), .A2(n14761), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14456), .ZN(n14458) );
  AOI21_X1 U15841 ( .B1(n14765), .B2(n14459), .A(n14458), .ZN(n14460) );
  OAI211_X1 U15842 ( .C1(n14879), .C2(n14462), .A(n14461), .B(n14460), .ZN(
        P2_U3213) );
  MUX2_X1 U15843 ( .A(n14548), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14485), .Z(
        P2_U3562) );
  MUX2_X1 U15844 ( .A(n14463), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14485), .Z(
        P2_U3561) );
  MUX2_X1 U15845 ( .A(n14464), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14485), .Z(
        P2_U3560) );
  MUX2_X1 U15846 ( .A(n14465), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14485), .Z(
        P2_U3559) );
  MUX2_X1 U15847 ( .A(n14580), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14485), .Z(
        P2_U3558) );
  MUX2_X1 U15848 ( .A(n14466), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14485), .Z(
        P2_U3557) );
  MUX2_X1 U15849 ( .A(n14614), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14485), .Z(
        P2_U3556) );
  MUX2_X1 U15850 ( .A(n14646), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14485), .Z(
        P2_U3554) );
  MUX2_X1 U15851 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14632), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15852 ( .A(n14648), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14485), .Z(
        P2_U3552) );
  MUX2_X1 U15853 ( .A(n14467), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14485), .Z(
        P2_U3551) );
  MUX2_X1 U15854 ( .A(n14468), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14485), .Z(
        P2_U3550) );
  MUX2_X1 U15855 ( .A(n14469), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14485), .Z(
        P2_U3549) );
  MUX2_X1 U15856 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n14470), .S(P2_U3947), .Z(
        P2_U3547) );
  MUX2_X1 U15857 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n14471), .S(P2_U3947), .Z(
        P2_U3546) );
  MUX2_X1 U15858 ( .A(n14792), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14485), .Z(
        P2_U3545) );
  MUX2_X1 U15859 ( .A(n14472), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14485), .Z(
        P2_U3544) );
  MUX2_X1 U15860 ( .A(n14473), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14485), .Z(
        P2_U3543) );
  MUX2_X1 U15861 ( .A(n14474), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14485), .Z(
        P2_U3542) );
  MUX2_X1 U15862 ( .A(n14475), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14485), .Z(
        P2_U3541) );
  MUX2_X1 U15863 ( .A(n14476), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14485), .Z(
        P2_U3540) );
  MUX2_X1 U15864 ( .A(n14477), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14485), .Z(
        P2_U3539) );
  MUX2_X1 U15865 ( .A(n14478), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14485), .Z(
        P2_U3538) );
  MUX2_X1 U15866 ( .A(n14479), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14485), .Z(
        P2_U3537) );
  MUX2_X1 U15867 ( .A(n14480), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14485), .Z(
        P2_U3536) );
  MUX2_X1 U15868 ( .A(n14481), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14485), .Z(
        P2_U3535) );
  MUX2_X1 U15869 ( .A(n14482), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14485), .Z(
        P2_U3534) );
  MUX2_X1 U15870 ( .A(n14483), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14485), .Z(
        P2_U3533) );
  MUX2_X1 U15871 ( .A(n14484), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14485), .Z(
        P2_U3532) );
  MUX2_X1 U15872 ( .A(n9882), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14485), .Z(
        P2_U3531) );
  OAI22_X1 U15873 ( .A1(n15904), .A2(n9173), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14486), .ZN(n14487) );
  AOI21_X1 U15874 ( .B1(n14488), .B2(n15892), .A(n14487), .ZN(n14499) );
  INV_X1 U15875 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n14491) );
  INV_X1 U15876 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n14489) );
  MUX2_X1 U15877 ( .A(n14489), .B(P2_REG2_REG_1__SCAN_IN), .S(n14488), .Z(
        n14490) );
  OAI21_X1 U15878 ( .B1(n11213), .B2(n14491), .A(n14490), .ZN(n14492) );
  NAND3_X1 U15879 ( .A1(n15898), .A2(n14493), .A3(n14492), .ZN(n14498) );
  OAI211_X1 U15880 ( .C1(n14496), .C2(n14495), .A(n15888), .B(n14494), .ZN(
        n14497) );
  NAND3_X1 U15881 ( .A1(n14499), .A2(n14498), .A3(n14497), .ZN(P2_U3215) );
  OAI21_X1 U15882 ( .B1(n15904), .B2(n15942), .A(n14500), .ZN(n14501) );
  AOI21_X1 U15883 ( .B1(n14504), .B2(n15892), .A(n14501), .ZN(n14511) );
  OAI211_X1 U15884 ( .C1(n14503), .C2(n14502), .A(n15898), .B(n14517), .ZN(
        n14510) );
  MUX2_X1 U15885 ( .A(n10905), .B(P2_REG1_REG_3__SCAN_IN), .S(n14504), .Z(
        n14506) );
  NAND3_X1 U15886 ( .A1(n14507), .A2(n14506), .A3(n14505), .ZN(n14508) );
  NAND3_X1 U15887 ( .A1(n15888), .A2(n14523), .A3(n14508), .ZN(n14509) );
  NAND3_X1 U15888 ( .A1(n14511), .A2(n14510), .A3(n14509), .ZN(P2_U3217) );
  INV_X1 U15889 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14513) );
  OAI21_X1 U15890 ( .B1(n15904), .B2(n14513), .A(n14512), .ZN(n14514) );
  AOI21_X1 U15891 ( .B1(n14515), .B2(n15892), .A(n14514), .ZN(n14529) );
  MUX2_X1 U15892 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10867), .S(n14521), .Z(
        n14518) );
  NAND3_X1 U15893 ( .A1(n14518), .A2(n14517), .A3(n14516), .ZN(n14519) );
  NAND3_X1 U15894 ( .A1(n15898), .A2(n14520), .A3(n14519), .ZN(n14528) );
  MUX2_X1 U15895 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10902), .S(n14521), .Z(
        n14524) );
  NAND3_X1 U15896 ( .A1(n14524), .A2(n14523), .A3(n14522), .ZN(n14525) );
  NAND3_X1 U15897 ( .A1(n15888), .A2(n14526), .A3(n14525), .ZN(n14527) );
  NAND3_X1 U15898 ( .A1(n14529), .A2(n14528), .A3(n14527), .ZN(P2_U3218) );
  MUX2_X1 U15899 ( .A(n11549), .B(P2_REG2_REG_6__SCAN_IN), .S(n14539), .Z(
        n14530) );
  NAND3_X1 U15900 ( .A1(n15830), .A2(n14531), .A3(n14530), .ZN(n14532) );
  NAND3_X1 U15901 ( .A1(n15898), .A2(n14533), .A3(n14532), .ZN(n14543) );
  MUX2_X1 U15902 ( .A(n10913), .B(P2_REG1_REG_6__SCAN_IN), .S(n14539), .Z(
        n14534) );
  NAND3_X1 U15903 ( .A1(n15827), .A2(n14535), .A3(n14534), .ZN(n14536) );
  NAND3_X1 U15904 ( .A1(n15888), .A2(n14537), .A3(n14536), .ZN(n14542) );
  AOI21_X1 U15905 ( .B1(n15858), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n14538), .ZN(
        n14541) );
  NAND2_X1 U15906 ( .A1(n15892), .A2(n14539), .ZN(n14540) );
  NAND4_X1 U15907 ( .A1(n14543), .A2(n14542), .A3(n14541), .A4(n14540), .ZN(
        P2_U3220) );
  INV_X1 U15908 ( .A(n14902), .ZN(n14812) );
  XNOR2_X1 U15909 ( .A(n14812), .B(n14552), .ZN(n14544) );
  NAND2_X1 U15910 ( .A1(n14544), .A2(n11678), .ZN(n14811) );
  NOR2_X1 U15911 ( .A1(n14805), .A2(n14545), .ZN(n14549) );
  INV_X1 U15912 ( .A(n14546), .ZN(n14547) );
  NAND2_X1 U15913 ( .A1(n14548), .A2(n14547), .ZN(n14813) );
  NOR2_X1 U15914 ( .A1(n16082), .A2(n14813), .ZN(n14554) );
  AOI211_X1 U15915 ( .C1(n14902), .C2(n14747), .A(n14549), .B(n14554), .ZN(
        n14550) );
  OAI21_X1 U15916 ( .B1(n14811), .B2(n14751), .A(n14550), .ZN(P2_U3234) );
  AOI21_X1 U15917 ( .B1(n14551), .B2(n14905), .A(n14300), .ZN(n14553) );
  NAND2_X1 U15918 ( .A1(n14553), .A2(n14552), .ZN(n14814) );
  AOI21_X1 U15919 ( .B1(n16094), .B2(P2_REG2_REG_30__SCAN_IN), .A(n14554), 
        .ZN(n14556) );
  NAND2_X1 U15920 ( .A1(n14905), .A2(n14747), .ZN(n14555) );
  OAI211_X1 U15921 ( .C1(n14814), .C2(n14751), .A(n14556), .B(n14555), .ZN(
        P2_U3235) );
  OAI21_X1 U15922 ( .B1(n14558), .B2(n14697), .A(n14557), .ZN(n14564) );
  AOI22_X1 U15923 ( .A1(n14560), .A2(n14747), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n16082), .ZN(n14561) );
  OAI21_X1 U15924 ( .B1(n14562), .B2(n14751), .A(n14561), .ZN(n14563) );
  INV_X1 U15925 ( .A(n14565), .ZN(P2_U3237) );
  OAI22_X1 U15926 ( .A1(n14567), .A2(n14697), .B1(n14566), .B2(n14805), .ZN(
        n14568) );
  AOI21_X1 U15927 ( .B1(n14569), .B2(n14747), .A(n14568), .ZN(n14570) );
  OAI21_X1 U15928 ( .B1(n14571), .B2(n14751), .A(n14570), .ZN(n14572) );
  AOI21_X1 U15929 ( .B1(n14573), .B2(n16089), .A(n14572), .ZN(n14574) );
  OAI21_X1 U15930 ( .B1(n14575), .B2(n16082), .A(n14574), .ZN(P2_U3238) );
  INV_X1 U15931 ( .A(n14576), .ZN(n14579) );
  NAND3_X1 U15932 ( .A1(n14593), .A2(n14587), .A3(n14577), .ZN(n14578) );
  AOI211_X1 U15933 ( .C1(n14819), .C2(n14603), .A(n14300), .B(n14581), .ZN(
        n14818) );
  AOI22_X1 U15934 ( .A1(n14582), .A2(n16080), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n16082), .ZN(n14583) );
  OAI21_X1 U15935 ( .B1(n14584), .B2(n16085), .A(n14583), .ZN(n14590) );
  OAI21_X1 U15936 ( .B1(n14587), .B2(n14586), .A(n14585), .ZN(n14588) );
  INV_X1 U15937 ( .A(n14588), .ZN(n14822) );
  NOR2_X1 U15938 ( .A1(n14822), .A2(n16062), .ZN(n14589) );
  AOI211_X1 U15939 ( .C1(n14818), .C2(n16088), .A(n14590), .B(n14589), .ZN(
        n14591) );
  OAI21_X1 U15940 ( .B1(n14821), .B2(n16082), .A(n14591), .ZN(P2_U3239) );
  XNOR2_X1 U15941 ( .A(n14592), .B(n8154), .ZN(n14825) );
  INV_X1 U15942 ( .A(n14825), .ZN(n14609) );
  INV_X1 U15943 ( .A(n14593), .ZN(n14596) );
  NOR3_X1 U15944 ( .A1(n14611), .A2(n14594), .A3(n8154), .ZN(n14595) );
  NOR2_X1 U15945 ( .A1(n14596), .A2(n14595), .ZN(n14597) );
  OAI222_X1 U15946 ( .A1(n14600), .A2(n14599), .B1(n14794), .B2(n14598), .C1(
        n14719), .C2(n14597), .ZN(n14823) );
  AOI21_X1 U15947 ( .B1(n14618), .B2(n14601), .A(n14300), .ZN(n14602) );
  NAND2_X1 U15948 ( .A1(n14824), .A2(n16088), .ZN(n14606) );
  AOI22_X1 U15949 ( .A1(n14604), .A2(n16080), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n16082), .ZN(n14605) );
  OAI211_X1 U15950 ( .C1(n14912), .C2(n16085), .A(n14606), .B(n14605), .ZN(
        n14607) );
  AOI21_X1 U15951 ( .B1(n14823), .B2(n14805), .A(n14607), .ZN(n14608) );
  OAI21_X1 U15952 ( .B1(n14609), .B2(n16062), .A(n14608), .ZN(P2_U3240) );
  XOR2_X1 U15953 ( .A(n14610), .B(n14613), .Z(n14828) );
  AOI21_X1 U15954 ( .B1(n14613), .B2(n14612), .A(n14611), .ZN(n14616) );
  AOI22_X1 U15955 ( .A1(n14614), .A2(n14791), .B1(n14647), .B2(n14646), .ZN(
        n14615) );
  OAI21_X1 U15956 ( .B1(n14616), .B2(n14719), .A(n14615), .ZN(n14617) );
  AOI21_X1 U15957 ( .B1(n14884), .B2(n14828), .A(n14617), .ZN(n14832) );
  INV_X1 U15958 ( .A(n14618), .ZN(n14619) );
  AOI211_X1 U15959 ( .C1(n14830), .C2(n14637), .A(n14300), .B(n14619), .ZN(
        n14829) );
  NOR2_X1 U15960 ( .A1(n14620), .A2(n16085), .ZN(n14625) );
  OAI22_X1 U15961 ( .A1(n14623), .A2(n14622), .B1(n14621), .B2(n14697), .ZN(
        n14624) );
  AOI211_X1 U15962 ( .C1(n14829), .C2(n16088), .A(n14625), .B(n14624), .ZN(
        n14627) );
  NAND2_X1 U15963 ( .A1(n14828), .A2(n16089), .ZN(n14626) );
  OAI211_X1 U15964 ( .C1(n14832), .C2(n16082), .A(n14627), .B(n14626), .ZN(
        P2_U3241) );
  XNOR2_X1 U15965 ( .A(n14628), .B(n14629), .ZN(n14918) );
  XNOR2_X1 U15966 ( .A(n14631), .B(n14630), .ZN(n14635) );
  AOI22_X1 U15967 ( .A1(n14633), .A2(n14791), .B1(n14647), .B2(n14632), .ZN(
        n14634) );
  OAI21_X1 U15968 ( .B1(n14635), .B2(n14719), .A(n14634), .ZN(n14636) );
  AOI21_X1 U15969 ( .B1(n14884), .B2(n14918), .A(n14636), .ZN(n14835) );
  OAI211_X1 U15970 ( .C1(n14914), .C2(n14651), .A(n14267), .B(n14637), .ZN(
        n14834) );
  OAI22_X1 U15971 ( .A1(n14805), .A2(n14639), .B1(n14638), .B2(n14697), .ZN(
        n14640) );
  AOI21_X1 U15972 ( .B1(n14641), .B2(n14747), .A(n14640), .ZN(n14642) );
  OAI21_X1 U15973 ( .B1(n14834), .B2(n14751), .A(n14642), .ZN(n14643) );
  AOI21_X1 U15974 ( .B1(n14918), .B2(n16089), .A(n14643), .ZN(n14644) );
  OAI21_X1 U15975 ( .B1(n14835), .B2(n16082), .A(n14644), .ZN(P2_U3242) );
  XOR2_X1 U15976 ( .A(n14645), .B(n14655), .Z(n14649) );
  AOI222_X1 U15977 ( .A1(n9112), .A2(n14649), .B1(n14648), .B2(n14647), .C1(
        n14646), .C2(n14791), .ZN(n14842) );
  OAI21_X1 U15978 ( .B1(n14654), .B2(n14662), .A(n14267), .ZN(n14650) );
  NOR2_X1 U15979 ( .A1(n14651), .A2(n14650), .ZN(n14839) );
  AOI22_X1 U15980 ( .A1(n16082), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14652), 
        .B2(n16080), .ZN(n14653) );
  OAI21_X1 U15981 ( .B1(n14654), .B2(n16085), .A(n14653), .ZN(n14658) );
  XNOR2_X1 U15982 ( .A(n14656), .B(n14655), .ZN(n14843) );
  NOR2_X1 U15983 ( .A1(n14843), .A2(n16062), .ZN(n14657) );
  AOI211_X1 U15984 ( .C1(n14839), .C2(n16088), .A(n14658), .B(n14657), .ZN(
        n14659) );
  OAI21_X1 U15985 ( .B1(n14842), .B2(n16082), .A(n14659), .ZN(P2_U3243) );
  XOR2_X1 U15986 ( .A(n14660), .B(n14667), .Z(n14845) );
  INV_X1 U15987 ( .A(n14845), .ZN(n14674) );
  OAI21_X1 U15988 ( .B1(n14925), .B2(n14676), .A(n14267), .ZN(n14661) );
  NOR2_X1 U15989 ( .A1(n14663), .A2(n14697), .ZN(n14664) );
  AOI21_X1 U15990 ( .B1(n16094), .B2(P2_REG2_REG_21__SCAN_IN), .A(n14664), 
        .ZN(n14665) );
  OAI21_X1 U15991 ( .B1(n14925), .B2(n16085), .A(n14665), .ZN(n14666) );
  AOI21_X1 U15992 ( .B1(n7239), .B2(n16088), .A(n14666), .ZN(n14673) );
  XOR2_X1 U15993 ( .A(n14668), .B(n14667), .Z(n14671) );
  INV_X1 U15994 ( .A(n14669), .ZN(n14670) );
  OAI21_X1 U15995 ( .B1(n14671), .B2(n14719), .A(n14670), .ZN(n14844) );
  NAND2_X1 U15996 ( .A1(n14844), .A2(n14805), .ZN(n14672) );
  OAI211_X1 U15997 ( .C1(n14674), .C2(n16062), .A(n14673), .B(n14672), .ZN(
        P2_U3244) );
  XOR2_X1 U15998 ( .A(n14675), .B(n14681), .Z(n14850) );
  INV_X1 U15999 ( .A(n14850), .ZN(n14687) );
  OAI21_X1 U16000 ( .B1(n14929), .B2(n14696), .A(n14267), .ZN(n14677) );
  NOR2_X1 U16001 ( .A1(n14677), .A2(n14676), .ZN(n14849) );
  AOI22_X1 U16002 ( .A1(n16082), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14678), 
        .B2(n16080), .ZN(n14679) );
  OAI21_X1 U16003 ( .B1(n14929), .B2(n16085), .A(n14679), .ZN(n14680) );
  AOI21_X1 U16004 ( .B1(n14849), .B2(n16088), .A(n14680), .ZN(n14686) );
  XOR2_X1 U16005 ( .A(n14682), .B(n14681), .Z(n14684) );
  OAI21_X1 U16006 ( .B1(n14684), .B2(n14719), .A(n14683), .ZN(n14848) );
  NAND2_X1 U16007 ( .A1(n14848), .A2(n14805), .ZN(n14685) );
  OAI211_X1 U16008 ( .C1(n14687), .C2(n16062), .A(n14686), .B(n14685), .ZN(
        P2_U3245) );
  XNOR2_X1 U16009 ( .A(n14689), .B(n14688), .ZN(n14691) );
  AOI21_X1 U16010 ( .B1(n14691), .B2(n9112), .A(n14690), .ZN(n14854) );
  XNOR2_X1 U16011 ( .A(n14692), .B(n14693), .ZN(n14856) );
  NAND2_X1 U16012 ( .A1(n14700), .A2(n14711), .ZN(n14694) );
  NAND2_X1 U16013 ( .A1(n14694), .A2(n14267), .ZN(n14695) );
  OR2_X1 U16014 ( .A1(n14696), .A2(n14695), .ZN(n14853) );
  OAI22_X1 U16015 ( .A1(n14805), .A2(n12052), .B1(n14698), .B2(n14697), .ZN(
        n14699) );
  AOI21_X1 U16016 ( .B1(n14700), .B2(n14747), .A(n14699), .ZN(n14701) );
  OAI21_X1 U16017 ( .B1(n14853), .B2(n14751), .A(n14701), .ZN(n14702) );
  AOI21_X1 U16018 ( .B1(n14856), .B2(n14753), .A(n14702), .ZN(n14703) );
  OAI21_X1 U16019 ( .B1(n16094), .B2(n14854), .A(n14703), .ZN(P2_U3246) );
  XNOR2_X1 U16020 ( .A(n14704), .B(n14707), .ZN(n14706) );
  AOI21_X1 U16021 ( .B1(n14706), .B2(n9112), .A(n14705), .ZN(n14860) );
  XNOR2_X1 U16022 ( .A(n14708), .B(n14707), .ZN(n14863) );
  INV_X1 U16023 ( .A(n14724), .ZN(n14709) );
  AOI21_X1 U16024 ( .B1(n14713), .B2(n14709), .A(n14300), .ZN(n14710) );
  NAND2_X1 U16025 ( .A1(n14711), .A2(n14710), .ZN(n14859) );
  AOI22_X1 U16026 ( .A1(n16094), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14712), 
        .B2(n16080), .ZN(n14715) );
  NAND2_X1 U16027 ( .A1(n14713), .A2(n14747), .ZN(n14714) );
  OAI211_X1 U16028 ( .C1(n14859), .C2(n14751), .A(n14715), .B(n14714), .ZN(
        n14716) );
  AOI21_X1 U16029 ( .B1(n14863), .B2(n14753), .A(n14716), .ZN(n14717) );
  OAI21_X1 U16030 ( .B1(n16094), .B2(n14860), .A(n14717), .ZN(P2_U3247) );
  INV_X1 U16031 ( .A(n14718), .ZN(n14720) );
  AOI21_X1 U16032 ( .B1(n14720), .B2(n14731), .A(n14719), .ZN(n14723) );
  AOI21_X1 U16033 ( .B1(n14723), .B2(n14722), .A(n14721), .ZN(n14869) );
  OAI21_X1 U16034 ( .B1(n14728), .B2(n14745), .A(n14267), .ZN(n14725) );
  NOR2_X1 U16035 ( .A1(n14725), .A2(n14724), .ZN(n14866) );
  AOI22_X1 U16036 ( .A1(n16094), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14726), 
        .B2(n16080), .ZN(n14727) );
  OAI21_X1 U16037 ( .B1(n14728), .B2(n16085), .A(n14727), .ZN(n14734) );
  OAI21_X1 U16038 ( .B1(n14731), .B2(n14730), .A(n14729), .ZN(n14732) );
  INV_X1 U16039 ( .A(n14732), .ZN(n14870) );
  NOR2_X1 U16040 ( .A1(n14870), .A2(n16062), .ZN(n14733) );
  AOI211_X1 U16041 ( .C1(n14866), .C2(n16088), .A(n14734), .B(n14733), .ZN(
        n14735) );
  OAI21_X1 U16042 ( .B1(n16094), .B2(n14869), .A(n14735), .ZN(P2_U3248) );
  OAI211_X1 U16043 ( .C1(n14737), .C2(n14740), .A(n14736), .B(n9112), .ZN(
        n14739) );
  AND2_X1 U16044 ( .A1(n14739), .A2(n14738), .ZN(n14875) );
  NAND2_X1 U16045 ( .A1(n14741), .A2(n14740), .ZN(n14742) );
  NAND2_X1 U16046 ( .A1(n14743), .A2(n14742), .ZN(n14942) );
  INV_X1 U16047 ( .A(n14942), .ZN(n14754) );
  OAI21_X1 U16048 ( .B1(n14872), .B2(n14763), .A(n14267), .ZN(n14744) );
  OR2_X1 U16049 ( .A1(n14745), .A2(n14744), .ZN(n14871) );
  AOI22_X1 U16050 ( .A1(n16094), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n14746), 
        .B2(n16080), .ZN(n14750) );
  NAND2_X1 U16051 ( .A1(n14748), .A2(n14747), .ZN(n14749) );
  OAI211_X1 U16052 ( .C1(n14871), .C2(n14751), .A(n14750), .B(n14749), .ZN(
        n14752) );
  AOI21_X1 U16053 ( .B1(n14754), .B2(n14753), .A(n14752), .ZN(n14755) );
  OAI21_X1 U16054 ( .B1(n16094), .B2(n14875), .A(n14755), .ZN(P2_U3249) );
  XNOR2_X1 U16055 ( .A(n14756), .B(n14757), .ZN(n14885) );
  INV_X1 U16056 ( .A(n14885), .ZN(n14946) );
  NAND2_X1 U16057 ( .A1(n14758), .A2(n14757), .ZN(n14759) );
  NAND3_X1 U16058 ( .A1(n14760), .A2(n9112), .A3(n14759), .ZN(n14762) );
  NAND2_X1 U16059 ( .A1(n14762), .A2(n14761), .ZN(n14882) );
  OAI21_X1 U16060 ( .B1(n14879), .B2(n14774), .A(n14267), .ZN(n14764) );
  NOR2_X1 U16061 ( .A1(n14764), .A2(n14763), .ZN(n14880) );
  NAND2_X1 U16062 ( .A1(n14880), .A2(n16088), .ZN(n14767) );
  AOI22_X1 U16063 ( .A1(n16094), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14765), 
        .B2(n16080), .ZN(n14766) );
  OAI211_X1 U16064 ( .C1(n14879), .C2(n16085), .A(n14767), .B(n14766), .ZN(
        n14768) );
  AOI21_X1 U16065 ( .B1(n14882), .B2(n14805), .A(n14768), .ZN(n14769) );
  OAI21_X1 U16066 ( .B1(n14946), .B2(n16062), .A(n14769), .ZN(P2_U3250) );
  XNOR2_X1 U16067 ( .A(n14771), .B(n14770), .ZN(n14773) );
  AOI21_X1 U16068 ( .B1(n14773), .B2(n9112), .A(n14772), .ZN(n14891) );
  AOI211_X1 U16069 ( .C1(n14889), .C2(n14802), .A(n14300), .B(n14774), .ZN(
        n14888) );
  AOI22_X1 U16070 ( .A1(n16082), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14775), 
        .B2(n16080), .ZN(n14776) );
  OAI21_X1 U16071 ( .B1(n14777), .B2(n16085), .A(n14776), .ZN(n14783) );
  OAI21_X1 U16072 ( .B1(n14780), .B2(n14779), .A(n14778), .ZN(n14781) );
  INV_X1 U16073 ( .A(n14781), .ZN(n14892) );
  NOR2_X1 U16074 ( .A1(n14892), .A2(n16062), .ZN(n14782) );
  AOI211_X1 U16075 ( .C1(n14888), .C2(n16088), .A(n14783), .B(n14782), .ZN(
        n14784) );
  OAI21_X1 U16076 ( .B1(n16094), .B2(n14891), .A(n14784), .ZN(P2_U3251) );
  OAI21_X1 U16077 ( .B1(n14787), .B2(n14786), .A(n14785), .ZN(n14954) );
  OAI21_X1 U16078 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n14797) );
  NAND2_X1 U16079 ( .A1(n14792), .A2(n14791), .ZN(n14793) );
  OAI21_X1 U16080 ( .B1(n14795), .B2(n14794), .A(n14793), .ZN(n14796) );
  AOI21_X1 U16081 ( .B1(n14797), .B2(n9112), .A(n14796), .ZN(n14798) );
  OAI21_X1 U16082 ( .B1(n14954), .B2(n14876), .A(n14798), .ZN(n14894) );
  AOI21_X1 U16083 ( .B1(n14799), .B2(n16080), .A(n14894), .ZN(n14810) );
  AOI21_X1 U16084 ( .B1(n14801), .B2(n14800), .A(n14300), .ZN(n14803) );
  AND2_X1 U16085 ( .A1(n14803), .A2(n14802), .ZN(n14893) );
  OAI22_X1 U16086 ( .A1(n14952), .A2(n16085), .B1(n14805), .B2(n14804), .ZN(
        n14808) );
  NOR2_X1 U16087 ( .A1(n14954), .A2(n14806), .ZN(n14807) );
  AOI211_X1 U16088 ( .C1(n14893), .C2(n16088), .A(n14808), .B(n14807), .ZN(
        n14809) );
  OAI21_X1 U16089 ( .B1(n16094), .B2(n14810), .A(n14809), .ZN(P2_U3252) );
  NAND2_X1 U16090 ( .A1(n14814), .A2(n14813), .ZN(n14903) );
  MUX2_X1 U16091 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14903), .S(n16208), .Z(
        n14815) );
  AOI21_X1 U16092 ( .B1(n14816), .B2(n14905), .A(n14815), .ZN(n14817) );
  INV_X1 U16093 ( .A(n14817), .ZN(P2_U3529) );
  AOI21_X1 U16094 ( .B1(n16134), .B2(n14819), .A(n14818), .ZN(n14820) );
  OAI211_X1 U16095 ( .C1(n16138), .C2(n14822), .A(n14821), .B(n14820), .ZN(
        n14908) );
  MUX2_X1 U16096 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14908), .S(n16208), .Z(
        P2_U3525) );
  INV_X1 U16097 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14826) );
  AOI211_X1 U16098 ( .C1(n16204), .C2(n14825), .A(n14824), .B(n14823), .ZN(
        n14909) );
  MUX2_X1 U16099 ( .A(n14826), .B(n14909), .S(n16208), .Z(n14827) );
  OAI21_X1 U16100 ( .B1(n14912), .B2(n14896), .A(n14827), .ZN(P2_U3524) );
  INV_X1 U16101 ( .A(n14828), .ZN(n14833) );
  AOI21_X1 U16102 ( .B1(n16134), .B2(n14830), .A(n14829), .ZN(n14831) );
  OAI211_X1 U16103 ( .C1(n9243), .C2(n14833), .A(n14832), .B(n14831), .ZN(
        n14913) );
  MUX2_X1 U16104 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14913), .S(n16208), .Z(
        P2_U3523) );
  NAND2_X1 U16105 ( .A1(n14835), .A2(n14834), .ZN(n14915) );
  MUX2_X1 U16106 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14915), .S(n16208), .Z(
        n14838) );
  INV_X1 U16107 ( .A(n14918), .ZN(n14836) );
  OAI22_X1 U16108 ( .A1(n14836), .A2(n14897), .B1(n14914), .B2(n14896), .ZN(
        n14837) );
  OR2_X1 U16109 ( .A1(n14838), .A2(n14837), .ZN(P2_U3522) );
  AOI21_X1 U16110 ( .B1(n16134), .B2(n14840), .A(n14839), .ZN(n14841) );
  OAI211_X1 U16111 ( .C1(n16138), .C2(n14843), .A(n14842), .B(n14841), .ZN(
        n14921) );
  MUX2_X1 U16112 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14921), .S(n16208), .Z(
        P2_U3521) );
  INV_X1 U16113 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14846) );
  AOI211_X1 U16114 ( .C1(n16204), .C2(n14845), .A(n7239), .B(n14844), .ZN(
        n14922) );
  MUX2_X1 U16115 ( .A(n14846), .B(n14922), .S(n16208), .Z(n14847) );
  OAI21_X1 U16116 ( .B1(n14925), .B2(n14896), .A(n14847), .ZN(P2_U3520) );
  INV_X1 U16117 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n14851) );
  AOI211_X1 U16118 ( .C1(n14850), .C2(n16204), .A(n14849), .B(n14848), .ZN(
        n14926) );
  MUX2_X1 U16119 ( .A(n14851), .B(n14926), .S(n16208), .Z(n14852) );
  OAI21_X1 U16120 ( .B1(n14929), .B2(n14896), .A(n14852), .ZN(P2_U3519) );
  INV_X1 U16121 ( .A(n14856), .ZN(n14933) );
  OAI211_X1 U16122 ( .C1(n8126), .C2(n16201), .A(n14854), .B(n14853), .ZN(
        n14855) );
  AOI21_X1 U16123 ( .B1(n14884), .B2(n14856), .A(n14855), .ZN(n14930) );
  MUX2_X1 U16124 ( .A(n14857), .B(n14930), .S(n16208), .Z(n14858) );
  OAI21_X1 U16125 ( .B1(n14933), .B2(n14897), .A(n14858), .ZN(P2_U3518) );
  INV_X1 U16126 ( .A(n14863), .ZN(n14937) );
  OAI211_X1 U16127 ( .C1(n14861), .C2(n16201), .A(n14860), .B(n14859), .ZN(
        n14862) );
  AOI21_X1 U16128 ( .B1(n14884), .B2(n14863), .A(n14862), .ZN(n14935) );
  INV_X1 U16129 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14864) );
  MUX2_X1 U16130 ( .A(n14935), .B(n14864), .S(n16206), .Z(n14865) );
  OAI21_X1 U16131 ( .B1(n14937), .B2(n14897), .A(n14865), .ZN(P2_U3517) );
  AOI21_X1 U16132 ( .B1(n16134), .B2(n14867), .A(n14866), .ZN(n14868) );
  OAI211_X1 U16133 ( .C1(n14870), .C2(n16138), .A(n14869), .B(n14868), .ZN(
        n14938) );
  MUX2_X1 U16134 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14938), .S(n16208), .Z(
        P2_U3516) );
  OAI21_X1 U16135 ( .B1(n14872), .B2(n16201), .A(n14871), .ZN(n14873) );
  INV_X1 U16136 ( .A(n14873), .ZN(n14874) );
  OAI211_X1 U16137 ( .C1(n14942), .C2(n14876), .A(n14875), .B(n14874), .ZN(
        n14939) );
  MUX2_X1 U16138 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14939), .S(n16208), .Z(
        n14877) );
  INV_X1 U16139 ( .A(n14877), .ZN(n14878) );
  OAI21_X1 U16140 ( .B1(n14942), .B2(n14897), .A(n14878), .ZN(P2_U3515) );
  INV_X1 U16141 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14886) );
  NOR2_X1 U16142 ( .A1(n14879), .A2(n16201), .ZN(n14881) );
  AOI21_X1 U16143 ( .B1(n14885), .B2(n14884), .A(n14883), .ZN(n14943) );
  MUX2_X1 U16144 ( .A(n14886), .B(n14943), .S(n16208), .Z(n14887) );
  OAI21_X1 U16145 ( .B1(n14946), .B2(n14897), .A(n14887), .ZN(P2_U3514) );
  AOI21_X1 U16146 ( .B1(n16134), .B2(n14889), .A(n14888), .ZN(n14890) );
  OAI211_X1 U16147 ( .C1(n14892), .C2(n16138), .A(n14891), .B(n14890), .ZN(
        n14947) );
  MUX2_X1 U16148 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14947), .S(n16208), .Z(
        P2_U3513) );
  INV_X1 U16149 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14895) );
  NOR2_X1 U16150 ( .A1(n14894), .A2(n14893), .ZN(n14949) );
  MUX2_X1 U16151 ( .A(n14895), .B(n14949), .S(n16208), .Z(n14900) );
  OAI22_X1 U16152 ( .A1(n14954), .A2(n14897), .B1(n14952), .B2(n14896), .ZN(
        n14898) );
  INV_X1 U16153 ( .A(n14898), .ZN(n14899) );
  NAND2_X1 U16154 ( .A1(n14900), .A2(n14899), .ZN(P2_U3512) );
  INV_X1 U16155 ( .A(n14951), .ZN(n14906) );
  MUX2_X1 U16156 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14903), .S(n14948), .Z(
        n14904) );
  AOI21_X1 U16157 ( .B1(n14906), .B2(n14905), .A(n14904), .ZN(n14907) );
  INV_X1 U16158 ( .A(n14907), .ZN(P2_U3497) );
  MUX2_X1 U16159 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14908), .S(n14948), .Z(
        P2_U3493) );
  INV_X1 U16160 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14910) );
  MUX2_X1 U16161 ( .A(n14910), .B(n14909), .S(n14948), .Z(n14911) );
  OAI21_X1 U16162 ( .B1(n14912), .B2(n14951), .A(n14911), .ZN(P2_U3492) );
  MUX2_X1 U16163 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14913), .S(n14948), .Z(
        P2_U3491) );
  NOR2_X1 U16164 ( .A1(n14914), .A2(n14951), .ZN(n14917) );
  MUX2_X1 U16165 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14915), .S(n14948), .Z(
        n14916) );
  AOI211_X1 U16166 ( .C1(n14919), .C2(n14918), .A(n14917), .B(n14916), .ZN(
        n14920) );
  INV_X1 U16167 ( .A(n14920), .ZN(P2_U3490) );
  MUX2_X1 U16168 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14921), .S(n14948), .Z(
        P2_U3489) );
  INV_X1 U16169 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14923) );
  MUX2_X1 U16170 ( .A(n14923), .B(n14922), .S(n14948), .Z(n14924) );
  OAI21_X1 U16171 ( .B1(n14925), .B2(n14951), .A(n14924), .ZN(P2_U3488) );
  INV_X1 U16172 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14927) );
  MUX2_X1 U16173 ( .A(n14927), .B(n14926), .S(n14948), .Z(n14928) );
  OAI21_X1 U16174 ( .B1(n14929), .B2(n14951), .A(n14928), .ZN(P2_U3487) );
  INV_X1 U16175 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14931) );
  MUX2_X1 U16176 ( .A(n14931), .B(n14930), .S(n14948), .Z(n14932) );
  OAI21_X1 U16177 ( .B1(n14933), .B2(n14953), .A(n14932), .ZN(P2_U3486) );
  INV_X1 U16178 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14934) );
  MUX2_X1 U16179 ( .A(n14935), .B(n14934), .S(n16209), .Z(n14936) );
  OAI21_X1 U16180 ( .B1(n14937), .B2(n14953), .A(n14936), .ZN(P2_U3484) );
  MUX2_X1 U16181 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14938), .S(n14948), .Z(
        P2_U3481) );
  MUX2_X1 U16182 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14939), .S(n14948), .Z(
        n14940) );
  INV_X1 U16183 ( .A(n14940), .ZN(n14941) );
  OAI21_X1 U16184 ( .B1(n14942), .B2(n14953), .A(n14941), .ZN(P2_U3478) );
  INV_X1 U16185 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14944) );
  MUX2_X1 U16186 ( .A(n14944), .B(n14943), .S(n14948), .Z(n14945) );
  OAI21_X1 U16187 ( .B1(n14946), .B2(n14953), .A(n14945), .ZN(P2_U3475) );
  MUX2_X1 U16188 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14947), .S(n14948), .Z(
        P2_U3472) );
  INV_X1 U16189 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14950) );
  MUX2_X1 U16190 ( .A(n14950), .B(n14949), .S(n14948), .Z(n14957) );
  OAI22_X1 U16191 ( .A1(n14954), .A2(n14953), .B1(n14952), .B2(n14951), .ZN(
        n14955) );
  INV_X1 U16192 ( .A(n14955), .ZN(n14956) );
  NAND2_X1 U16193 ( .A1(n14957), .A2(n14956), .ZN(P2_U3469) );
  INV_X1 U16194 ( .A(n14958), .ZN(n15763) );
  OAI222_X1 U16195 ( .A1(n14975), .A2(n15763), .B1(P2_U3088), .B2(n8609), .C1(
        n14959), .C2(n14970), .ZN(P2_U3298) );
  AOI21_X1 U16196 ( .B1(n14973), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14960), 
        .ZN(n14961) );
  OAI21_X1 U16197 ( .B1(n14962), .B2(n14975), .A(n14961), .ZN(P2_U3299) );
  INV_X1 U16198 ( .A(n14963), .ZN(n15767) );
  OAI222_X1 U16199 ( .A1(P2_U3088), .A2(n14965), .B1(n14968), .B2(n15767), 
        .C1(n14964), .C2(n14970), .ZN(P2_U3301) );
  INV_X1 U16200 ( .A(n14966), .ZN(n15770) );
  OAI222_X1 U16201 ( .A1(n14970), .A2(n14969), .B1(n14968), .B2(n15770), .C1(
        P2_U3088), .C2(n14967), .ZN(P2_U3302) );
  INV_X1 U16202 ( .A(n14971), .ZN(n15777) );
  AOI21_X1 U16203 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14973), .A(n14972), 
        .ZN(n14974) );
  OAI21_X1 U16204 ( .B1(n15777), .B2(n14975), .A(n14974), .ZN(P2_U3304) );
  MUX2_X1 U16205 ( .A(n14976), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U16206 ( .A1(n15705), .A2(n15062), .ZN(n14978) );
  NAND2_X1 U16207 ( .A1(n15369), .A2(n11123), .ZN(n14977) );
  NAND2_X1 U16208 ( .A1(n14978), .A2(n14977), .ZN(n14979) );
  XNOR2_X1 U16209 ( .A(n14979), .B(n15065), .ZN(n15002) );
  INV_X1 U16210 ( .A(n15369), .ZN(n15397) );
  OAI22_X1 U16211 ( .A1(n15597), .A2(n15095), .B1(n15397), .B2(n15094), .ZN(
        n15001) );
  NAND2_X1 U16212 ( .A1(n15729), .A2(n15062), .ZN(n14984) );
  NAND2_X1 U16213 ( .A1(n15223), .A2(n11123), .ZN(n14983) );
  NAND2_X1 U16214 ( .A1(n14984), .A2(n14983), .ZN(n14985) );
  XNOR2_X1 U16215 ( .A(n14985), .B(n7251), .ZN(n14986) );
  INV_X1 U16216 ( .A(n14986), .ZN(n14987) );
  XNOR2_X1 U16217 ( .A(n14988), .B(n14986), .ZN(n15208) );
  AOI22_X1 U16218 ( .A1(n15729), .A2(n11123), .B1(n15050), .B2(n15223), .ZN(
        n15209) );
  NAND2_X1 U16219 ( .A1(n15719), .A2(n15062), .ZN(n14990) );
  NAND2_X1 U16220 ( .A1(n15393), .A2(n11123), .ZN(n14989) );
  NAND2_X1 U16221 ( .A1(n14990), .A2(n14989), .ZN(n14991) );
  XNOR2_X1 U16222 ( .A(n14991), .B(n15065), .ZN(n14992) );
  AOI22_X1 U16223 ( .A1(n15719), .A2(n11123), .B1(n15050), .B2(n15393), .ZN(
        n14993) );
  XNOR2_X1 U16224 ( .A(n14992), .B(n14993), .ZN(n15133) );
  INV_X1 U16225 ( .A(n14992), .ZN(n14994) );
  AOI22_X1 U16226 ( .A1(n15711), .A2(n11123), .B1(n15050), .B2(n15581), .ZN(
        n14998) );
  NAND2_X1 U16227 ( .A1(n15711), .A2(n15062), .ZN(n14996) );
  NAND2_X1 U16228 ( .A1(n15581), .A2(n11123), .ZN(n14995) );
  NAND2_X1 U16229 ( .A1(n14996), .A2(n14995), .ZN(n14997) );
  XNOR2_X1 U16230 ( .A(n14997), .B(n15065), .ZN(n15000) );
  XOR2_X1 U16231 ( .A(n14998), .B(n15000), .Z(n15142) );
  INV_X1 U16232 ( .A(n14998), .ZN(n14999) );
  XOR2_X1 U16233 ( .A(n15001), .B(n15002), .Z(n15189) );
  NAND2_X1 U16234 ( .A1(n15698), .A2(n15062), .ZN(n15004) );
  NAND2_X1 U16235 ( .A1(n15584), .A2(n11123), .ZN(n15003) );
  NAND2_X1 U16236 ( .A1(n15004), .A2(n15003), .ZN(n15005) );
  XNOR2_X1 U16237 ( .A(n15005), .B(n15065), .ZN(n15006) );
  AOI22_X1 U16238 ( .A1(n15698), .A2(n11123), .B1(n15050), .B2(n15584), .ZN(
        n15007) );
  XNOR2_X1 U16239 ( .A(n15006), .B(n15007), .ZN(n15081) );
  INV_X1 U16240 ( .A(n15006), .ZN(n15008) );
  NAND2_X1 U16241 ( .A1(n15008), .A2(n15007), .ZN(n15009) );
  AND2_X1 U16242 ( .A1(n15400), .A2(n15050), .ZN(n15011) );
  AOI21_X1 U16243 ( .B1(n15688), .B2(n11123), .A(n15011), .ZN(n15017) );
  NAND2_X1 U16244 ( .A1(n15688), .A2(n15062), .ZN(n15013) );
  NAND2_X1 U16245 ( .A1(n15400), .A2(n11123), .ZN(n15012) );
  NAND2_X1 U16246 ( .A1(n15013), .A2(n15012), .ZN(n15014) );
  XNOR2_X1 U16247 ( .A(n15014), .B(n15065), .ZN(n15019) );
  XOR2_X1 U16248 ( .A(n15017), .B(n15019), .Z(n15164) );
  INV_X1 U16249 ( .A(n15017), .ZN(n15018) );
  NAND2_X1 U16250 ( .A1(n15019), .A2(n15018), .ZN(n15020) );
  AOI22_X1 U16251 ( .A1(n15679), .A2(n15062), .B1(n11123), .B2(n15402), .ZN(
        n15021) );
  XNOR2_X1 U16252 ( .A(n15021), .B(n15065), .ZN(n15024) );
  AOI22_X1 U16253 ( .A1(n15679), .A2(n11123), .B1(n15050), .B2(n15402), .ZN(
        n15023) );
  XNOR2_X1 U16254 ( .A(n15024), .B(n15023), .ZN(n15116) );
  INV_X1 U16255 ( .A(n15116), .ZN(n15022) );
  NAND2_X1 U16256 ( .A1(n15024), .A2(n15023), .ZN(n15025) );
  OAI22_X1 U16257 ( .A1(n15529), .A2(n15096), .B1(n15376), .B2(n15095), .ZN(
        n15026) );
  XNOR2_X1 U16258 ( .A(n15026), .B(n15065), .ZN(n15028) );
  AND2_X1 U16259 ( .A1(n15501), .A2(n15050), .ZN(n15027) );
  AOI21_X1 U16260 ( .B1(n15672), .B2(n11123), .A(n15027), .ZN(n15029) );
  XNOR2_X1 U16261 ( .A(n15028), .B(n15029), .ZN(n15170) );
  INV_X1 U16262 ( .A(n15028), .ZN(n15030) );
  NAND2_X1 U16263 ( .A1(n15030), .A2(n15029), .ZN(n15031) );
  NAND2_X1 U16264 ( .A1(n15667), .A2(n15062), .ZN(n15033) );
  NAND2_X1 U16265 ( .A1(n15406), .A2(n11123), .ZN(n15032) );
  NAND2_X1 U16266 ( .A1(n15033), .A2(n15032), .ZN(n15034) );
  XNOR2_X1 U16267 ( .A(n15034), .B(n15065), .ZN(n15035) );
  AOI22_X1 U16268 ( .A1(n15667), .A2(n11123), .B1(n15050), .B2(n15406), .ZN(
        n15036) );
  XNOR2_X1 U16269 ( .A(n15035), .B(n15036), .ZN(n15074) );
  INV_X1 U16270 ( .A(n15035), .ZN(n15037) );
  NAND2_X1 U16271 ( .A1(n15037), .A2(n15036), .ZN(n15038) );
  NAND2_X1 U16272 ( .A1(n15662), .A2(n15062), .ZN(n15040) );
  NAND2_X1 U16273 ( .A1(n15502), .A2(n11123), .ZN(n15039) );
  NAND2_X1 U16274 ( .A1(n15040), .A2(n15039), .ZN(n15041) );
  XNOR2_X1 U16275 ( .A(n15041), .B(n15065), .ZN(n15042) );
  AOI22_X1 U16276 ( .A1(n15662), .A2(n11123), .B1(n15050), .B2(n15502), .ZN(
        n15043) );
  XNOR2_X1 U16277 ( .A(n15042), .B(n15043), .ZN(n15150) );
  INV_X1 U16278 ( .A(n15042), .ZN(n15044) );
  NAND2_X1 U16279 ( .A1(n15044), .A2(n15043), .ZN(n15045) );
  NAND2_X1 U16280 ( .A1(n15654), .A2(n15062), .ZN(n15048) );
  NAND2_X1 U16281 ( .A1(n15378), .A2(n11123), .ZN(n15047) );
  NAND2_X1 U16282 ( .A1(n15048), .A2(n15047), .ZN(n15049) );
  XNOR2_X1 U16283 ( .A(n15049), .B(n15065), .ZN(n15051) );
  AOI22_X1 U16284 ( .A1(n15654), .A2(n11123), .B1(n15050), .B2(n15378), .ZN(
        n15052) );
  XNOR2_X1 U16285 ( .A(n15051), .B(n15052), .ZN(n15124) );
  INV_X1 U16286 ( .A(n15051), .ZN(n15053) );
  NAND2_X1 U16287 ( .A1(n15053), .A2(n15052), .ZN(n15054) );
  INV_X1 U16288 ( .A(n15439), .ZN(n15409) );
  OAI22_X1 U16289 ( .A1(n15648), .A2(n15095), .B1(n15409), .B2(n15094), .ZN(
        n15059) );
  NAND2_X1 U16290 ( .A1(n15459), .A2(n15062), .ZN(n15056) );
  NAND2_X1 U16291 ( .A1(n15439), .A2(n11123), .ZN(n15055) );
  NAND2_X1 U16292 ( .A1(n15056), .A2(n15055), .ZN(n15057) );
  XNOR2_X1 U16293 ( .A(n15057), .B(n15065), .ZN(n15058) );
  XOR2_X1 U16294 ( .A(n15059), .B(n15058), .Z(n15200) );
  INV_X1 U16295 ( .A(n15058), .ZN(n15061) );
  INV_X1 U16296 ( .A(n15059), .ZN(n15060) );
  OAI22_X1 U16297 ( .A1(n15447), .A2(n15095), .B1(n15410), .B2(n15094), .ZN(
        n15089) );
  NAND2_X1 U16298 ( .A1(n15643), .A2(n15062), .ZN(n15064) );
  NAND2_X1 U16299 ( .A1(n15222), .A2(n11123), .ZN(n15063) );
  NAND2_X1 U16300 ( .A1(n15064), .A2(n15063), .ZN(n15066) );
  XNOR2_X1 U16301 ( .A(n15066), .B(n15065), .ZN(n15088) );
  XOR2_X1 U16302 ( .A(n15089), .B(n15088), .Z(n15092) );
  XNOR2_X1 U16303 ( .A(n15093), .B(n15092), .ZN(n15067) );
  NAND2_X1 U16304 ( .A1(n15067), .A2(n15210), .ZN(n15072) );
  NOR2_X1 U16305 ( .A1(n15193), .A2(n15381), .ZN(n15070) );
  OAI22_X1 U16306 ( .A1(n15191), .A2(n15409), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15068), .ZN(n15069) );
  AOI211_X1 U16307 ( .C1(n15216), .C2(n15445), .A(n15070), .B(n15069), .ZN(
        n15071) );
  OAI211_X1 U16308 ( .C1(n15447), .C2(n15220), .A(n15072), .B(n15071), .ZN(
        P1_U3214) );
  XOR2_X1 U16309 ( .A(n15074), .B(n15073), .Z(n15080) );
  OAI22_X1 U16310 ( .A1(n15191), .A2(n15376), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15075), .ZN(n15078) );
  INV_X1 U16311 ( .A(n15506), .ZN(n15076) );
  OAI22_X1 U16312 ( .A1(n15192), .A2(n15076), .B1(n8118), .B2(n15193), .ZN(
        n15077) );
  AOI211_X1 U16313 ( .C1(n15667), .C2(n15196), .A(n15078), .B(n15077), .ZN(
        n15079) );
  OAI21_X1 U16314 ( .B1(n15080), .B2(n15205), .A(n15079), .ZN(P1_U3216) );
  XOR2_X1 U16315 ( .A(n15082), .B(n15081), .Z(n15087) );
  NOR2_X1 U16316 ( .A1(n15192), .A2(n15569), .ZN(n15085) );
  AND2_X1 U16317 ( .A1(n15369), .A2(n15582), .ZN(n15083) );
  AOI21_X1 U16318 ( .B1(n15400), .B2(n15583), .A(n15083), .ZN(n15696) );
  NAND2_X1 U16319 ( .A1(n7190), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15346) );
  OAI21_X1 U16320 ( .B1(n15696), .B2(n15213), .A(n15346), .ZN(n15084) );
  AOI211_X1 U16321 ( .C1(n15698), .C2(n15196), .A(n15085), .B(n15084), .ZN(
        n15086) );
  OAI21_X1 U16322 ( .B1(n15087), .B2(n15205), .A(n15086), .ZN(P1_U3219) );
  INV_X1 U16323 ( .A(n15088), .ZN(n15091) );
  INV_X1 U16324 ( .A(n15089), .ZN(n15090) );
  OAI22_X1 U16325 ( .A1(n15427), .A2(n15095), .B1(n15381), .B2(n15094), .ZN(
        n15099) );
  OAI22_X1 U16326 ( .A1(n15427), .A2(n15096), .B1(n15381), .B2(n15095), .ZN(
        n15097) );
  XNOR2_X1 U16327 ( .A(n15097), .B(n15065), .ZN(n15098) );
  XOR2_X1 U16328 ( .A(n15099), .B(n15098), .Z(n15100) );
  AOI22_X1 U16329 ( .A1(n15500), .A2(n15222), .B1(n15221), .B2(n15583), .ZN(
        n15421) );
  OAI22_X1 U16330 ( .A1(n15421), .A2(n15213), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15101), .ZN(n15103) );
  NOR2_X1 U16331 ( .A1(n15427), .A2(n15220), .ZN(n15102) );
  AOI211_X1 U16332 ( .C1(n15425), .C2(n15216), .A(n15103), .B(n15102), .ZN(
        n15104) );
  OAI21_X1 U16333 ( .B1(n15107), .B2(n15106), .A(n15105), .ZN(n15108) );
  NAND2_X1 U16334 ( .A1(n15108), .A2(n15210), .ZN(n15112) );
  AOI22_X1 U16335 ( .A1(n15182), .A2(n15236), .B1(n15196), .B2(n15109), .ZN(
        n15111) );
  AOI22_X1 U16336 ( .A1(n15184), .A2(n15238), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n15183), .ZN(n15110) );
  NAND3_X1 U16337 ( .A1(n15112), .A2(n15111), .A3(n15110), .ZN(P1_U3222) );
  INV_X1 U16338 ( .A(n15113), .ZN(n15114) );
  AOI21_X1 U16339 ( .B1(n15116), .B2(n15115), .A(n15114), .ZN(n15122) );
  AND2_X1 U16340 ( .A1(n15501), .A2(n15583), .ZN(n15117) );
  AOI21_X1 U16341 ( .B1(n15400), .B2(n15582), .A(n15117), .ZN(n15677) );
  INV_X1 U16342 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n15118) );
  OAI22_X1 U16343 ( .A1(n15677), .A2(n15213), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15118), .ZN(n15119) );
  AOI21_X1 U16344 ( .B1(n15540), .B2(n15216), .A(n15119), .ZN(n15121) );
  NAND2_X1 U16345 ( .A1(n15679), .A2(n15196), .ZN(n15120) );
  OAI211_X1 U16346 ( .C1(n15122), .C2(n15205), .A(n15121), .B(n15120), .ZN(
        P1_U3223) );
  XOR2_X1 U16347 ( .A(n15124), .B(n15123), .Z(n15131) );
  NAND2_X1 U16348 ( .A1(n15502), .A2(n15500), .ZN(n15126) );
  NAND2_X1 U16349 ( .A1(n15439), .A2(n15583), .ZN(n15125) );
  AND2_X1 U16350 ( .A1(n15126), .A2(n15125), .ZN(n15656) );
  OAI22_X1 U16351 ( .A1(n15656), .A2(n15213), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15127), .ZN(n15129) );
  NOR2_X1 U16352 ( .A1(n15470), .A2(n15220), .ZN(n15128) );
  AOI211_X1 U16353 ( .C1(n15216), .C2(n15473), .A(n15129), .B(n15128), .ZN(
        n15130) );
  OAI21_X1 U16354 ( .B1(n15131), .B2(n15205), .A(n15130), .ZN(P1_U3225) );
  XOR2_X1 U16355 ( .A(n15133), .B(n15132), .Z(n15140) );
  OAI22_X1 U16356 ( .A1(n15135), .A2(n15213), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15134), .ZN(n15136) );
  AOI21_X1 U16357 ( .B1(n15137), .B2(n15216), .A(n15136), .ZN(n15139) );
  NAND2_X1 U16358 ( .A1(n15719), .A2(n15196), .ZN(n15138) );
  OAI211_X1 U16359 ( .C1(n15140), .C2(n15205), .A(n15139), .B(n15138), .ZN(
        P1_U3226) );
  XOR2_X1 U16360 ( .A(n15142), .B(n15141), .Z(n15148) );
  NAND2_X1 U16361 ( .A1(n15369), .A2(n15437), .ZN(n15144) );
  NAND2_X1 U16362 ( .A1(n15393), .A2(n15500), .ZN(n15143) );
  NAND2_X1 U16363 ( .A1(n15144), .A2(n15143), .ZN(n15710) );
  AOI22_X1 U16364 ( .A1(n15710), .A2(n15159), .B1(P1_REG3_REG_17__SCAN_IN), 
        .B2(P1_U3086), .ZN(n15145) );
  OAI21_X1 U16365 ( .B1(n15614), .B2(n15192), .A(n15145), .ZN(n15146) );
  AOI21_X1 U16366 ( .B1(n15711), .B2(n15196), .A(n15146), .ZN(n15147) );
  OAI21_X1 U16367 ( .B1(n15148), .B2(n15205), .A(n15147), .ZN(P1_U3228) );
  XOR2_X1 U16368 ( .A(n15150), .B(n15149), .Z(n15156) );
  OAI22_X1 U16369 ( .A1(n15191), .A2(n7468), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15151), .ZN(n15154) );
  INV_X1 U16370 ( .A(n15492), .ZN(n15152) );
  INV_X1 U16371 ( .A(n15378), .ZN(n15483) );
  OAI22_X1 U16372 ( .A1(n15192), .A2(n15152), .B1(n15483), .B2(n15193), .ZN(
        n15153) );
  AOI211_X1 U16373 ( .C1(n15662), .C2(n15196), .A(n15154), .B(n15153), .ZN(
        n15155) );
  OAI21_X1 U16374 ( .B1(n15156), .B2(n15205), .A(n15155), .ZN(P1_U3229) );
  NAND2_X1 U16375 ( .A1(n15402), .A2(n15437), .ZN(n15158) );
  NAND2_X1 U16376 ( .A1(n15584), .A2(n15500), .ZN(n15157) );
  NAND2_X1 U16377 ( .A1(n15158), .A2(n15157), .ZN(n15687) );
  AOI22_X1 U16378 ( .A1(n15687), .A2(n15159), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(n7190), .ZN(n15160) );
  OAI21_X1 U16379 ( .B1(n15555), .B2(n15192), .A(n15160), .ZN(n15166) );
  INV_X1 U16380 ( .A(n15161), .ZN(n15162) );
  AOI211_X1 U16381 ( .C1(n15164), .C2(n15163), .A(n15205), .B(n15162), .ZN(
        n15165) );
  AOI211_X1 U16382 ( .C1(n15688), .C2(n15196), .A(n15166), .B(n15165), .ZN(
        n15167) );
  INV_X1 U16383 ( .A(n15167), .ZN(P1_U3233) );
  OAI21_X1 U16384 ( .B1(n15170), .B2(n15168), .A(n15169), .ZN(n15171) );
  NAND2_X1 U16385 ( .A1(n15171), .A2(n15210), .ZN(n15176) );
  AND2_X1 U16386 ( .A1(n15406), .A2(n15583), .ZN(n15172) );
  AOI21_X1 U16387 ( .B1(n15402), .B2(n15500), .A(n15172), .ZN(n15517) );
  OAI22_X1 U16388 ( .A1(n15517), .A2(n15213), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15173), .ZN(n15174) );
  AOI21_X1 U16389 ( .B1(n15526), .B2(n15216), .A(n15174), .ZN(n15175) );
  OAI211_X1 U16390 ( .C1(n15220), .C2(n15529), .A(n15176), .B(n15175), .ZN(
        P1_U3235) );
  OAI21_X1 U16391 ( .B1(n15179), .B2(n15178), .A(n15177), .ZN(n15180) );
  NAND2_X1 U16392 ( .A1(n15180), .A2(n15210), .ZN(n15187) );
  AOI22_X1 U16393 ( .A1(n15182), .A2(n15235), .B1(n15196), .B2(n15181), .ZN(
        n15186) );
  AOI22_X1 U16394 ( .A1(n15184), .A2(n12736), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n15183), .ZN(n15185) );
  NAND3_X1 U16395 ( .A1(n15187), .A2(n15186), .A3(n15185), .ZN(P1_U3237) );
  XOR2_X1 U16396 ( .A(n15189), .B(n15188), .Z(n15198) );
  OAI22_X1 U16397 ( .A1(n15191), .A2(n15367), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15190), .ZN(n15195) );
  INV_X1 U16398 ( .A(n15584), .ZN(n15371) );
  OAI22_X1 U16399 ( .A1(n15371), .A2(n15193), .B1(n15192), .B2(n15594), .ZN(
        n15194) );
  AOI211_X1 U16400 ( .C1(n15705), .C2(n15196), .A(n15195), .B(n15194), .ZN(
        n15197) );
  OAI21_X1 U16401 ( .B1(n15198), .B2(n15205), .A(n15197), .ZN(P1_U3238) );
  XOR2_X1 U16402 ( .A(n15200), .B(n15199), .Z(n15206) );
  AOI22_X1 U16403 ( .A1(n15500), .A2(n15378), .B1(n15222), .B2(n15437), .ZN(
        n15452) );
  OAI22_X1 U16404 ( .A1(n15452), .A2(n15213), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15201), .ZN(n15203) );
  NOR2_X1 U16405 ( .A1(n15648), .A2(n15220), .ZN(n15202) );
  AOI211_X1 U16406 ( .C1(n15216), .C2(n15458), .A(n15203), .B(n15202), .ZN(
        n15204) );
  OAI21_X1 U16407 ( .B1(n15206), .B2(n15205), .A(n15204), .ZN(P1_U3240) );
  OAI21_X1 U16408 ( .B1(n15209), .B2(n15208), .A(n15207), .ZN(n15211) );
  NAND2_X1 U16409 ( .A1(n15211), .A2(n15210), .ZN(n15219) );
  OAI21_X1 U16410 ( .B1(n15214), .B2(n15213), .A(n15212), .ZN(n15215) );
  AOI21_X1 U16411 ( .B1(n15217), .B2(n15216), .A(n15215), .ZN(n15218) );
  OAI211_X1 U16412 ( .C1(n8025), .C2(n15220), .A(n15219), .B(n15218), .ZN(
        P1_U3241) );
  MUX2_X1 U16413 ( .A(n15353), .B(P1_DATAO_REG_31__SCAN_IN), .S(n15237), .Z(
        P1_U3591) );
  MUX2_X1 U16414 ( .A(n15385), .B(P1_DATAO_REG_30__SCAN_IN), .S(n15237), .Z(
        P1_U3590) );
  MUX2_X1 U16415 ( .A(n15221), .B(P1_DATAO_REG_29__SCAN_IN), .S(n15237), .Z(
        P1_U3589) );
  MUX2_X1 U16416 ( .A(n15438), .B(P1_DATAO_REG_28__SCAN_IN), .S(n15237), .Z(
        P1_U3588) );
  MUX2_X1 U16417 ( .A(n15222), .B(P1_DATAO_REG_27__SCAN_IN), .S(n15237), .Z(
        P1_U3587) );
  MUX2_X1 U16418 ( .A(n15439), .B(P1_DATAO_REG_26__SCAN_IN), .S(n15237), .Z(
        P1_U3586) );
  MUX2_X1 U16419 ( .A(n15378), .B(P1_DATAO_REG_25__SCAN_IN), .S(n15237), .Z(
        P1_U3585) );
  MUX2_X1 U16420 ( .A(n15502), .B(P1_DATAO_REG_24__SCAN_IN), .S(n15237), .Z(
        P1_U3584) );
  MUX2_X1 U16421 ( .A(n15406), .B(P1_DATAO_REG_23__SCAN_IN), .S(n15237), .Z(
        P1_U3583) );
  MUX2_X1 U16422 ( .A(n15501), .B(P1_DATAO_REG_22__SCAN_IN), .S(n15237), .Z(
        P1_U3582) );
  MUX2_X1 U16423 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15402), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16424 ( .A(n15400), .B(P1_DATAO_REG_20__SCAN_IN), .S(n15237), .Z(
        P1_U3580) );
  MUX2_X1 U16425 ( .A(n15584), .B(P1_DATAO_REG_19__SCAN_IN), .S(n15237), .Z(
        P1_U3579) );
  MUX2_X1 U16426 ( .A(n15369), .B(P1_DATAO_REG_18__SCAN_IN), .S(n15237), .Z(
        P1_U3578) );
  MUX2_X1 U16427 ( .A(n15581), .B(P1_DATAO_REG_17__SCAN_IN), .S(n15237), .Z(
        P1_U3577) );
  MUX2_X1 U16428 ( .A(n15393), .B(P1_DATAO_REG_16__SCAN_IN), .S(n15237), .Z(
        P1_U3576) );
  MUX2_X1 U16429 ( .A(n15223), .B(P1_DATAO_REG_15__SCAN_IN), .S(n15237), .Z(
        P1_U3575) );
  MUX2_X1 U16430 ( .A(n15224), .B(P1_DATAO_REG_14__SCAN_IN), .S(n15237), .Z(
        P1_U3574) );
  MUX2_X1 U16431 ( .A(n15225), .B(P1_DATAO_REG_13__SCAN_IN), .S(n15237), .Z(
        P1_U3573) );
  MUX2_X1 U16432 ( .A(n15226), .B(P1_DATAO_REG_12__SCAN_IN), .S(n15237), .Z(
        P1_U3572) );
  MUX2_X1 U16433 ( .A(n15227), .B(P1_DATAO_REG_11__SCAN_IN), .S(n15237), .Z(
        P1_U3571) );
  MUX2_X1 U16434 ( .A(n15228), .B(P1_DATAO_REG_10__SCAN_IN), .S(n15237), .Z(
        P1_U3570) );
  MUX2_X1 U16435 ( .A(n15229), .B(P1_DATAO_REG_9__SCAN_IN), .S(n15237), .Z(
        P1_U3569) );
  MUX2_X1 U16436 ( .A(n15230), .B(P1_DATAO_REG_8__SCAN_IN), .S(n15237), .Z(
        P1_U3568) );
  MUX2_X1 U16437 ( .A(n15231), .B(P1_DATAO_REG_7__SCAN_IN), .S(n15237), .Z(
        P1_U3567) );
  MUX2_X1 U16438 ( .A(n15232), .B(P1_DATAO_REG_6__SCAN_IN), .S(n15237), .Z(
        P1_U3566) );
  MUX2_X1 U16439 ( .A(n15233), .B(P1_DATAO_REG_5__SCAN_IN), .S(n15237), .Z(
        P1_U3565) );
  MUX2_X1 U16440 ( .A(n15234), .B(P1_DATAO_REG_4__SCAN_IN), .S(n15237), .Z(
        P1_U3564) );
  MUX2_X1 U16441 ( .A(n15235), .B(P1_DATAO_REG_3__SCAN_IN), .S(n15237), .Z(
        P1_U3563) );
  MUX2_X1 U16442 ( .A(n15236), .B(P1_DATAO_REG_2__SCAN_IN), .S(n15237), .Z(
        P1_U3562) );
  MUX2_X1 U16443 ( .A(n12736), .B(P1_DATAO_REG_1__SCAN_IN), .S(n15237), .Z(
        P1_U3561) );
  MUX2_X1 U16444 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15238), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16445 ( .C1(n15241), .C2(n15240), .A(n15927), .B(n15239), .ZN(
        n15248) );
  NAND2_X1 U16446 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n15249) );
  OAI211_X1 U16447 ( .C1(n15243), .C2(n10278), .A(n15931), .B(n15242), .ZN(
        n15247) );
  AOI22_X1 U16448 ( .A1(n15914), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n7190), .ZN(n15246) );
  NAND2_X1 U16449 ( .A1(n15929), .A2(n15244), .ZN(n15245) );
  NAND4_X1 U16450 ( .A1(n15248), .A2(n15247), .A3(n15246), .A4(n15245), .ZN(
        P1_U3244) );
  MUX2_X1 U16451 ( .A(n15250), .B(n15249), .S(n15905), .Z(n15252) );
  NOR2_X1 U16452 ( .A1(n15351), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n15251) );
  OR2_X1 U16453 ( .A1(n10290), .A2(n15251), .ZN(n15906) );
  INV_X1 U16454 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15908) );
  NAND2_X1 U16455 ( .A1(n15906), .A2(n15908), .ZN(n15911) );
  OAI211_X1 U16456 ( .C1(n15252), .C2(n10290), .A(P1_U4016), .B(n15911), .ZN(
        n15294) );
  NOR2_X1 U16457 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11047), .ZN(n15253) );
  AOI21_X1 U16458 ( .B1(n15914), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n15253), .ZN(
        n15254) );
  OAI21_X1 U16459 ( .B1(n15337), .B2(n15255), .A(n15254), .ZN(n15256) );
  INV_X1 U16460 ( .A(n15256), .ZN(n15264) );
  OAI211_X1 U16461 ( .C1(n15258), .C2(n15257), .A(n15931), .B(n15272), .ZN(
        n15263) );
  OAI211_X1 U16462 ( .C1(n15261), .C2(n15260), .A(n15927), .B(n15259), .ZN(
        n15262) );
  NAND4_X1 U16463 ( .A1(n15294), .A2(n15264), .A3(n15263), .A4(n15262), .ZN(
        P1_U3245) );
  AND2_X1 U16464 ( .A1(n7190), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n15266) );
  NOR2_X1 U16465 ( .A1(n15337), .A2(n15270), .ZN(n15265) );
  AOI211_X1 U16466 ( .C1(n15914), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n15266), .B(
        n15265), .ZN(n15277) );
  OAI211_X1 U16467 ( .C1(n15269), .C2(n15268), .A(n15927), .B(n15267), .ZN(
        n15276) );
  MUX2_X1 U16468 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11068), .S(n15270), .Z(
        n15273) );
  NAND3_X1 U16469 ( .A1(n15273), .A2(n15272), .A3(n15271), .ZN(n15274) );
  NAND3_X1 U16470 ( .A1(n15931), .A2(n15281), .A3(n15274), .ZN(n15275) );
  NAND3_X1 U16471 ( .A1(n15277), .A2(n15276), .A3(n15275), .ZN(P1_U3246) );
  INV_X1 U16472 ( .A(n15278), .ZN(n15279) );
  AOI21_X1 U16473 ( .B1(n15914), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n15279), .ZN(
        n15293) );
  MUX2_X1 U16474 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10277), .S(n15286), .Z(
        n15282) );
  NAND3_X1 U16475 ( .A1(n15282), .A2(n15281), .A3(n15280), .ZN(n15283) );
  NAND2_X1 U16476 ( .A1(n15284), .A2(n15283), .ZN(n15285) );
  OAI22_X1 U16477 ( .A1(n15286), .A2(n15337), .B1(n15338), .B2(n15285), .ZN(
        n15287) );
  INV_X1 U16478 ( .A(n15287), .ZN(n15292) );
  OAI211_X1 U16479 ( .C1(n15290), .C2(n15289), .A(n15927), .B(n15288), .ZN(
        n15291) );
  NAND4_X1 U16480 ( .A1(n15294), .A2(n15293), .A3(n15292), .A4(n15291), .ZN(
        P1_U3247) );
  INV_X1 U16481 ( .A(n15295), .ZN(n15298) );
  NOR2_X1 U16482 ( .A1(n15337), .A2(n15296), .ZN(n15297) );
  AOI211_X1 U16483 ( .C1(n15914), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n15298), .B(
        n15297), .ZN(n15311) );
  OAI211_X1 U16484 ( .C1(n15301), .C2(n15300), .A(n15927), .B(n15299), .ZN(
        n15310) );
  INV_X1 U16485 ( .A(n15302), .ZN(n15305) );
  MUX2_X1 U16486 ( .A(n11381), .B(P1_REG2_REG_6__SCAN_IN), .S(n15303), .Z(
        n15304) );
  NAND2_X1 U16487 ( .A1(n15305), .A2(n15304), .ZN(n15307) );
  OAI211_X1 U16488 ( .C1(n15308), .C2(n15307), .A(n15931), .B(n15306), .ZN(
        n15309) );
  NAND3_X1 U16489 ( .A1(n15311), .A2(n15310), .A3(n15309), .ZN(P1_U3249) );
  OAI211_X1 U16490 ( .C1(n15314), .C2(n15313), .A(n15312), .B(n15927), .ZN(
        n15328) );
  INV_X1 U16491 ( .A(n15315), .ZN(n15318) );
  NOR2_X1 U16492 ( .A1(n15337), .A2(n15316), .ZN(n15317) );
  AOI211_X1 U16493 ( .C1(n15914), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n15318), 
        .B(n15317), .ZN(n15327) );
  INV_X1 U16494 ( .A(n15319), .ZN(n15322) );
  MUX2_X1 U16495 ( .A(n10586), .B(P1_REG2_REG_10__SCAN_IN), .S(n15320), .Z(
        n15321) );
  NAND2_X1 U16496 ( .A1(n15322), .A2(n15321), .ZN(n15324) );
  OAI211_X1 U16497 ( .C1(n15325), .C2(n15324), .A(n15323), .B(n15931), .ZN(
        n15326) );
  NAND3_X1 U16498 ( .A1(n15328), .A2(n15327), .A3(n15326), .ZN(P1_U3253) );
  INV_X1 U16499 ( .A(n15342), .ZN(n15340) );
  NAND2_X1 U16500 ( .A1(n15332), .A2(n15331), .ZN(n15335) );
  NAND2_X1 U16501 ( .A1(n15333), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n15334) );
  NAND2_X1 U16502 ( .A1(n15335), .A2(n15334), .ZN(n15336) );
  XOR2_X1 U16503 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n15336), .Z(n15341) );
  OAI21_X1 U16504 ( .B1(n15341), .B2(n15338), .A(n15337), .ZN(n15339) );
  AOI21_X1 U16505 ( .B1(n15340), .B2(n15927), .A(n15339), .ZN(n15345) );
  AOI22_X1 U16506 ( .A1(n15342), .A2(n15927), .B1(n15931), .B2(n15341), .ZN(
        n15344) );
  MUX2_X1 U16507 ( .A(n15345), .B(n15344), .S(n15343), .Z(n15347) );
  OAI211_X1 U16508 ( .C1(n15348), .C2(n15935), .A(n15347), .B(n15346), .ZN(
        P1_U3262) );
  INV_X1 U16509 ( .A(n15688), .ZN(n15550) );
  OR2_X2 U16510 ( .A1(n15667), .A2(n15524), .ZN(n15504) );
  NAND2_X1 U16511 ( .A1(n15383), .A2(n15627), .ZN(n15357) );
  XOR2_X1 U16512 ( .A(n15354), .B(n15357), .Z(n15349) );
  NAND2_X1 U16513 ( .A1(n15349), .A2(n16153), .ZN(n15623) );
  OR2_X1 U16514 ( .A1(n15351), .A2(n15350), .ZN(n15352) );
  AND2_X1 U16515 ( .A1(n15583), .A2(n15352), .ZN(n15384) );
  NAND2_X1 U16516 ( .A1(n15353), .A2(n15384), .ZN(n15625) );
  NOR2_X1 U16517 ( .A1(n16022), .A2(n15625), .ZN(n15359) );
  INV_X1 U16518 ( .A(n15354), .ZN(n15624) );
  NOR2_X1 U16519 ( .A1(n15624), .A2(n16014), .ZN(n15355) );
  AOI211_X1 U16520 ( .C1(n16022), .C2(P1_REG2_REG_31__SCAN_IN), .A(n15359), 
        .B(n15355), .ZN(n15356) );
  OAI21_X1 U16521 ( .B1(n15363), .B2(n15623), .A(n15356), .ZN(P1_U3263) );
  OAI211_X1 U16522 ( .C1(n15383), .C2(n15627), .A(n16153), .B(n15357), .ZN(
        n15626) );
  NOR2_X1 U16523 ( .A1(n15611), .A2(n15358), .ZN(n15360) );
  AOI211_X1 U16524 ( .C1(n15361), .C2(n15617), .A(n15360), .B(n15359), .ZN(
        n15362) );
  OAI21_X1 U16525 ( .B1(n15626), .B2(n15363), .A(n15362), .ZN(P1_U3264) );
  INV_X1 U16526 ( .A(n15393), .ZN(n15364) );
  NAND2_X1 U16527 ( .A1(n15719), .A2(n15364), .ZN(n15365) );
  INV_X1 U16528 ( .A(n15603), .ZN(n15608) );
  AND2_X1 U16529 ( .A1(n15711), .A2(n15367), .ZN(n15368) );
  NAND2_X1 U16530 ( .A1(n15597), .A2(n15369), .ZN(n15370) );
  NAND2_X1 U16531 ( .A1(n15698), .A2(n15371), .ZN(n15372) );
  INV_X1 U16532 ( .A(n15400), .ZN(n15373) );
  INV_X1 U16533 ( .A(n15667), .ZN(n15508) );
  NAND2_X1 U16534 ( .A1(n15385), .A2(n15384), .ZN(n15630) );
  OAI22_X1 U16535 ( .A1(n15387), .A2(n15630), .B1(n15386), .B2(n15615), .ZN(
        n15389) );
  NAND2_X1 U16536 ( .A1(n15438), .A2(n15500), .ZN(n15631) );
  NOR2_X1 U16537 ( .A1(n16022), .A2(n15631), .ZN(n15388) );
  AOI211_X1 U16538 ( .C1(n16022), .C2(P1_REG2_REG_29__SCAN_IN), .A(n15389), 
        .B(n15388), .ZN(n15390) );
  OAI21_X1 U16539 ( .B1(n15391), .B2(n16014), .A(n15390), .ZN(n15392) );
  AOI21_X1 U16540 ( .B1(n15632), .B2(n15429), .A(n15392), .ZN(n15414) );
  OR2_X1 U16541 ( .A1(n15719), .A2(n15393), .ZN(n15394) );
  NAND2_X1 U16542 ( .A1(n15711), .A2(n15581), .ZN(n15396) );
  NAND2_X1 U16543 ( .A1(n15597), .A2(n15397), .ZN(n15398) );
  OR2_X1 U16544 ( .A1(n15698), .A2(n15584), .ZN(n15399) );
  NAND2_X1 U16545 ( .A1(n15688), .A2(n15400), .ZN(n15401) );
  NOR2_X1 U16546 ( .A1(n15679), .A2(n15402), .ZN(n15403) );
  OR2_X1 U16547 ( .A1(n15672), .A2(n15501), .ZN(n15405) );
  INV_X1 U16548 ( .A(n15407), .ZN(n15408) );
  INV_X1 U16549 ( .A(n15420), .ZN(n15415) );
  NAND2_X1 U16550 ( .A1(n15416), .A2(n15415), .ZN(n15418) );
  NAND2_X1 U16551 ( .A1(n15629), .A2(n15620), .ZN(n15413) );
  OAI211_X1 U16552 ( .C1(n15628), .C2(n15622), .A(n15414), .B(n15413), .ZN(
        P1_U3356) );
  OAI211_X1 U16553 ( .C1(n7328), .C2(n15420), .A(n15419), .B(n15723), .ZN(
        n15422) );
  NAND2_X1 U16554 ( .A1(n15635), .A2(n15611), .ZN(n15432) );
  AOI21_X1 U16555 ( .B1(n15443), .B2(n15636), .A(n16096), .ZN(n15424) );
  NAND2_X1 U16556 ( .A1(n15424), .A2(n15423), .ZN(n15638) );
  INV_X1 U16557 ( .A(n15638), .ZN(n15430) );
  AOI22_X1 U16558 ( .A1(n16022), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n15425), 
        .B2(n16011), .ZN(n15426) );
  OAI21_X1 U16559 ( .B1(n15427), .B2(n16014), .A(n15426), .ZN(n15428) );
  AOI21_X1 U16560 ( .B1(n15430), .B2(n15429), .A(n15428), .ZN(n15431) );
  OAI211_X1 U16561 ( .C1(n15577), .C2(n15640), .A(n15432), .B(n15431), .ZN(
        P1_U3265) );
  XNOR2_X1 U16562 ( .A(n15433), .B(n15434), .ZN(n15442) );
  AOI22_X1 U16563 ( .A1(n15582), .A2(n15439), .B1(n15438), .B2(n15437), .ZN(
        n15440) );
  INV_X1 U16564 ( .A(n15457), .ZN(n15444) );
  AOI21_X1 U16565 ( .B1(n15643), .B2(n15444), .A(n7487), .ZN(n15644) );
  AOI22_X1 U16566 ( .A1(n16022), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n15445), 
        .B2(n16011), .ZN(n15446) );
  OAI21_X1 U16567 ( .B1(n15447), .B2(n16014), .A(n15446), .ZN(n15449) );
  NOR2_X1 U16568 ( .A1(n15647), .A2(n15598), .ZN(n15448) );
  AOI211_X1 U16569 ( .C1(n15644), .C2(n15601), .A(n15449), .B(n15448), .ZN(
        n15450) );
  OAI21_X1 U16570 ( .B1(n16022), .B2(n15646), .A(n15450), .ZN(P1_U3266) );
  XOR2_X1 U16571 ( .A(n15455), .B(n15451), .Z(n15453) );
  OAI21_X1 U16572 ( .B1(n15453), .B2(n16074), .A(n15452), .ZN(n15650) );
  INV_X1 U16573 ( .A(n15650), .ZN(n15464) );
  XOR2_X1 U16574 ( .A(n15455), .B(n15454), .Z(n15652) );
  NOR2_X1 U16575 ( .A1(n15472), .A2(n15648), .ZN(n15456) );
  OR2_X1 U16576 ( .A1(n15457), .A2(n15456), .ZN(n15649) );
  AOI22_X1 U16577 ( .A1(n16022), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n15458), 
        .B2(n16011), .ZN(n15461) );
  NAND2_X1 U16578 ( .A1(n15459), .A2(n15617), .ZN(n15460) );
  OAI211_X1 U16579 ( .C1(n15649), .C2(n16015), .A(n15461), .B(n15460), .ZN(
        n15462) );
  AOI21_X1 U16580 ( .B1(n15652), .B2(n15620), .A(n15462), .ZN(n15463) );
  OAI21_X1 U16581 ( .B1(n15464), .B2(n16022), .A(n15463), .ZN(P1_U3267) );
  AOI21_X1 U16582 ( .B1(n15469), .B2(n15466), .A(n15465), .ZN(n15467) );
  INV_X1 U16583 ( .A(n15467), .ZN(n15661) );
  OAI21_X1 U16584 ( .B1(n7322), .B2(n15469), .A(n15468), .ZN(n15659) );
  NOR2_X1 U16585 ( .A1(n15491), .A2(n15470), .ZN(n15471) );
  OR2_X1 U16586 ( .A1(n15472), .A2(n15471), .ZN(n15657) );
  NAND2_X1 U16587 ( .A1(n16011), .A2(n15473), .ZN(n15475) );
  NAND2_X1 U16588 ( .A1(n16022), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n15474) );
  OAI211_X1 U16589 ( .C1(n15656), .C2(n16022), .A(n15475), .B(n15474), .ZN(
        n15476) );
  AOI21_X1 U16590 ( .B1(n15654), .B2(n15617), .A(n15476), .ZN(n15477) );
  OAI21_X1 U16591 ( .B1(n15657), .B2(n16015), .A(n15477), .ZN(n15478) );
  AOI21_X1 U16592 ( .B1(n15659), .B2(n15575), .A(n15478), .ZN(n15479) );
  OAI21_X1 U16593 ( .B1(n15577), .B2(n15661), .A(n15479), .ZN(P1_U3268) );
  OAI21_X1 U16594 ( .B1(n15481), .B2(n15487), .A(n15480), .ZN(n15494) );
  OAI22_X1 U16595 ( .A1(n7468), .A2(n15484), .B1(n15483), .B2(n15482), .ZN(
        n15489) );
  AOI211_X1 U16596 ( .C1(n15487), .C2(n15486), .A(n16074), .B(n15485), .ZN(
        n15488) );
  AOI211_X1 U16597 ( .C1(n15490), .C2(n15494), .A(n15489), .B(n15488), .ZN(
        n15665) );
  AOI21_X1 U16598 ( .B1(n15662), .B2(n15504), .A(n15491), .ZN(n15663) );
  AOI22_X1 U16599 ( .A1(n16022), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n15492), 
        .B2(n16011), .ZN(n15493) );
  OAI21_X1 U16600 ( .B1(n7546), .B2(n16014), .A(n15493), .ZN(n15496) );
  INV_X1 U16601 ( .A(n15494), .ZN(n15666) );
  NOR2_X1 U16602 ( .A1(n15666), .A2(n15598), .ZN(n15495) );
  AOI211_X1 U16603 ( .C1(n15663), .C2(n15601), .A(n15496), .B(n15495), .ZN(
        n15497) );
  OAI21_X1 U16604 ( .B1(n15665), .B2(n16022), .A(n15497), .ZN(P1_U3269) );
  XNOR2_X1 U16605 ( .A(n15499), .B(n15498), .ZN(n15503) );
  AOI222_X1 U16606 ( .A1(n15723), .A2(n15503), .B1(n15502), .B2(n15583), .C1(
        n15501), .C2(n15500), .ZN(n15670) );
  INV_X1 U16607 ( .A(n15504), .ZN(n15505) );
  AOI21_X1 U16608 ( .B1(n15667), .B2(n15524), .A(n15505), .ZN(n15668) );
  AOI22_X1 U16609 ( .A1(n16022), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n15506), 
        .B2(n16011), .ZN(n15507) );
  OAI21_X1 U16610 ( .B1(n15508), .B2(n16014), .A(n15507), .ZN(n15513) );
  AND2_X1 U16611 ( .A1(n15510), .A2(n15509), .ZN(n15511) );
  OR2_X1 U16612 ( .A1(n15511), .A2(n7315), .ZN(n15671) );
  NOR2_X1 U16613 ( .A1(n15671), .A2(n15577), .ZN(n15512) );
  AOI211_X1 U16614 ( .C1(n15668), .C2(n15601), .A(n15513), .B(n15512), .ZN(
        n15514) );
  OAI21_X1 U16615 ( .B1(n15670), .B2(n16022), .A(n15514), .ZN(P1_U3270) );
  AOI21_X1 U16616 ( .B1(n8205), .B2(n15516), .A(n15515), .ZN(n15518) );
  OAI21_X1 U16617 ( .B1(n15518), .B2(n16074), .A(n15517), .ZN(n15519) );
  INV_X1 U16618 ( .A(n15519), .ZN(n15675) );
  INV_X1 U16619 ( .A(n15520), .ZN(n15521) );
  AOI21_X1 U16620 ( .B1(n15523), .B2(n15522), .A(n15521), .ZN(n15676) );
  INV_X1 U16621 ( .A(n15676), .ZN(n15531) );
  INV_X1 U16622 ( .A(n15524), .ZN(n15525) );
  AOI21_X1 U16623 ( .B1(n15672), .B2(n15539), .A(n15525), .ZN(n15673) );
  NAND2_X1 U16624 ( .A1(n15673), .A2(n15601), .ZN(n15528) );
  AOI22_X1 U16625 ( .A1(n16022), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n15526), 
        .B2(n16011), .ZN(n15527) );
  OAI211_X1 U16626 ( .C1(n16014), .C2(n15529), .A(n15528), .B(n15527), .ZN(
        n15530) );
  AOI21_X1 U16627 ( .B1(n15531), .B2(n15620), .A(n15530), .ZN(n15532) );
  OAI21_X1 U16628 ( .B1(n15675), .B2(n16022), .A(n15532), .ZN(P1_U3271) );
  XNOR2_X1 U16629 ( .A(n15533), .B(n15535), .ZN(n15685) );
  OAI21_X1 U16630 ( .B1(n15536), .B2(n15535), .A(n15534), .ZN(n15537) );
  INV_X1 U16631 ( .A(n15537), .ZN(n15683) );
  NAND2_X1 U16632 ( .A1(n15679), .A2(n15552), .ZN(n15538) );
  NAND2_X1 U16633 ( .A1(n15539), .A2(n15538), .ZN(n15681) );
  AOI22_X1 U16634 ( .A1(n15540), .A2(n16011), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n16022), .ZN(n15541) );
  OAI21_X1 U16635 ( .B1(n15677), .B2(n16022), .A(n15541), .ZN(n15542) );
  AOI21_X1 U16636 ( .B1(n15679), .B2(n15617), .A(n15542), .ZN(n15543) );
  OAI21_X1 U16637 ( .B1(n15681), .B2(n16015), .A(n15543), .ZN(n15544) );
  AOI21_X1 U16638 ( .B1(n15683), .B2(n15575), .A(n15544), .ZN(n15545) );
  OAI21_X1 U16639 ( .B1(n15685), .B2(n15577), .A(n15545), .ZN(P1_U3272) );
  INV_X1 U16640 ( .A(n15549), .ZN(n15547) );
  OAI21_X1 U16641 ( .B1(n15548), .B2(n15547), .A(n15546), .ZN(n15695) );
  NOR2_X1 U16642 ( .A1(n7343), .A2(n15549), .ZN(n15686) );
  NOR2_X1 U16643 ( .A1(n15686), .A2(n15622), .ZN(n15559) );
  OR2_X1 U16644 ( .A1(n15550), .A2(n15568), .ZN(n15551) );
  NAND2_X1 U16645 ( .A1(n15552), .A2(n15551), .ZN(n15690) );
  NAND2_X1 U16646 ( .A1(n15687), .A2(n15611), .ZN(n15554) );
  NAND2_X1 U16647 ( .A1(n16022), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n15553) );
  OAI211_X1 U16648 ( .C1(n15615), .C2(n15555), .A(n15554), .B(n15553), .ZN(
        n15556) );
  AOI21_X1 U16649 ( .B1(n15688), .B2(n15617), .A(n15556), .ZN(n15557) );
  OAI21_X1 U16650 ( .B1(n15690), .B2(n16015), .A(n15557), .ZN(n15558) );
  AOI21_X1 U16651 ( .B1(n15559), .B2(n15692), .A(n15558), .ZN(n15560) );
  OAI21_X1 U16652 ( .B1(n15577), .B2(n15695), .A(n15560), .ZN(P1_U3273) );
  OAI21_X1 U16653 ( .B1(n15562), .B2(n8094), .A(n15561), .ZN(n15563) );
  INV_X1 U16654 ( .A(n15563), .ZN(n15704) );
  OAI21_X1 U16655 ( .B1(n15566), .B2(n15565), .A(n15564), .ZN(n15702) );
  AND2_X1 U16656 ( .A1(n15698), .A2(n15592), .ZN(n15567) );
  OR2_X1 U16657 ( .A1(n15568), .A2(n15567), .ZN(n15700) );
  INV_X1 U16658 ( .A(n15569), .ZN(n15570) );
  AOI22_X1 U16659 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(n16022), .B1(n15570), 
        .B2(n16011), .ZN(n15571) );
  OAI21_X1 U16660 ( .B1(n15696), .B2(n16022), .A(n15571), .ZN(n15572) );
  AOI21_X1 U16661 ( .B1(n15698), .B2(n15617), .A(n15572), .ZN(n15573) );
  OAI21_X1 U16662 ( .B1(n15700), .B2(n16015), .A(n15573), .ZN(n15574) );
  AOI21_X1 U16663 ( .B1(n15702), .B2(n15575), .A(n15574), .ZN(n15576) );
  OAI21_X1 U16664 ( .B1(n15704), .B2(n15577), .A(n15576), .ZN(P1_U3274) );
  INV_X1 U16665 ( .A(n15578), .ZN(n15579) );
  AOI21_X1 U16666 ( .B1(n15586), .B2(n15580), .A(n15579), .ZN(n15709) );
  AOI22_X1 U16667 ( .A1(n15584), .A2(n15583), .B1(n15582), .B2(n15581), .ZN(
        n15589) );
  OAI211_X1 U16668 ( .C1(n15587), .C2(n15586), .A(n15585), .B(n15723), .ZN(
        n15588) );
  OAI211_X1 U16669 ( .C1(n15709), .C2(n16002), .A(n15589), .B(n15588), .ZN(
        n15590) );
  INV_X1 U16670 ( .A(n15590), .ZN(n15708) );
  INV_X1 U16671 ( .A(n15591), .ZN(n15610) );
  INV_X1 U16672 ( .A(n15592), .ZN(n15593) );
  AOI21_X1 U16673 ( .B1(n15705), .B2(n15610), .A(n15593), .ZN(n15706) );
  INV_X1 U16674 ( .A(n15594), .ZN(n15595) );
  AOI22_X1 U16675 ( .A1(n16022), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15595), 
        .B2(n16011), .ZN(n15596) );
  OAI21_X1 U16676 ( .B1(n15597), .B2(n16014), .A(n15596), .ZN(n15600) );
  NOR2_X1 U16677 ( .A1(n15709), .A2(n15598), .ZN(n15599) );
  AOI211_X1 U16678 ( .C1(n15706), .C2(n15601), .A(n15600), .B(n15599), .ZN(
        n15602) );
  OAI21_X1 U16679 ( .B1(n16022), .B2(n15708), .A(n15602), .ZN(P1_U3275) );
  XNOR2_X1 U16680 ( .A(n15604), .B(n15603), .ZN(n15717) );
  INV_X1 U16681 ( .A(n15605), .ZN(n15606) );
  AOI21_X1 U16682 ( .B1(n15608), .B2(n15607), .A(n15606), .ZN(n15715) );
  NAND2_X1 U16683 ( .A1(n15711), .A2(n7335), .ZN(n15609) );
  NAND2_X1 U16684 ( .A1(n15610), .A2(n15609), .ZN(n15713) );
  NAND2_X1 U16685 ( .A1(n15710), .A2(n15611), .ZN(n15613) );
  NAND2_X1 U16686 ( .A1(n16022), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n15612) );
  OAI211_X1 U16687 ( .C1(n15615), .C2(n15614), .A(n15613), .B(n15612), .ZN(
        n15616) );
  AOI21_X1 U16688 ( .B1(n15711), .B2(n15617), .A(n15616), .ZN(n15618) );
  OAI21_X1 U16689 ( .B1(n15713), .B2(n16015), .A(n15618), .ZN(n15619) );
  AOI21_X1 U16690 ( .B1(n15715), .B2(n15620), .A(n15619), .ZN(n15621) );
  OAI21_X1 U16691 ( .B1(n15717), .B2(n15622), .A(n15621), .ZN(P1_U3276) );
  OAI211_X1 U16692 ( .C1(n16171), .C2(n15624), .A(n15623), .B(n15625), .ZN(
        n15741) );
  MUX2_X1 U16693 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15741), .S(n16179), .Z(
        P1_U3559) );
  OAI211_X1 U16694 ( .C1(n16171), .C2(n15627), .A(n15626), .B(n15625), .ZN(
        n15742) );
  MUX2_X1 U16695 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15742), .S(n16179), .Z(
        P1_U3558) );
  NAND2_X1 U16696 ( .A1(n15631), .A2(n15630), .ZN(n15633) );
  NAND2_X1 U16697 ( .A1(n15636), .A2(n16151), .ZN(n15637) );
  INV_X1 U16698 ( .A(n15641), .ZN(n15642) );
  MUX2_X1 U16699 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15743), .S(n16179), .Z(
        P1_U3556) );
  AOI22_X1 U16700 ( .A1(n15644), .A2(n16153), .B1(n15643), .B2(n16151), .ZN(
        n15645) );
  MUX2_X1 U16701 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15744), .S(n16179), .Z(
        P1_U3555) );
  OAI22_X1 U16702 ( .A1(n15649), .A2(n16096), .B1(n15648), .B2(n16171), .ZN(
        n15651) );
  AOI211_X1 U16703 ( .C1(n16176), .C2(n15652), .A(n15651), .B(n15650), .ZN(
        n15653) );
  INV_X1 U16704 ( .A(n15653), .ZN(n15745) );
  MUX2_X1 U16705 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15745), .S(n16179), .Z(
        P1_U3554) );
  NAND2_X1 U16706 ( .A1(n15654), .A2(n16151), .ZN(n15655) );
  OAI211_X1 U16707 ( .C1(n15657), .C2(n16096), .A(n15656), .B(n15655), .ZN(
        n15658) );
  AOI21_X1 U16708 ( .B1(n15659), .B2(n15723), .A(n15658), .ZN(n15660) );
  OAI21_X1 U16709 ( .B1(n15732), .B2(n15661), .A(n15660), .ZN(n15746) );
  MUX2_X1 U16710 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15746), .S(n16179), .Z(
        P1_U3553) );
  AOI22_X1 U16711 ( .A1(n15663), .A2(n16153), .B1(n15662), .B2(n16151), .ZN(
        n15664) );
  OAI211_X1 U16712 ( .C1(n15666), .C2(n16116), .A(n15665), .B(n15664), .ZN(
        n15747) );
  MUX2_X1 U16713 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15747), .S(n16179), .Z(
        P1_U3552) );
  AOI22_X1 U16714 ( .A1(n15668), .A2(n16153), .B1(n15667), .B2(n16151), .ZN(
        n15669) );
  OAI211_X1 U16715 ( .C1(n15732), .C2(n15671), .A(n15670), .B(n15669), .ZN(
        n15748) );
  MUX2_X1 U16716 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15748), .S(n16179), .Z(
        P1_U3551) );
  AOI22_X1 U16717 ( .A1(n15673), .A2(n16153), .B1(n15672), .B2(n16151), .ZN(
        n15674) );
  OAI211_X1 U16718 ( .C1(n15732), .C2(n15676), .A(n15675), .B(n15674), .ZN(
        n15749) );
  MUX2_X1 U16719 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15749), .S(n16179), .Z(
        P1_U3550) );
  INV_X1 U16720 ( .A(n15677), .ZN(n15678) );
  AOI21_X1 U16721 ( .B1(n15679), .B2(n16151), .A(n15678), .ZN(n15680) );
  OAI21_X1 U16722 ( .B1(n15681), .B2(n16096), .A(n15680), .ZN(n15682) );
  AOI21_X1 U16723 ( .B1(n15683), .B2(n15723), .A(n15682), .ZN(n15684) );
  OAI21_X1 U16724 ( .B1(n15732), .B2(n15685), .A(n15684), .ZN(n15750) );
  MUX2_X1 U16725 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15750), .S(n16179), .Z(
        P1_U3549) );
  NOR2_X1 U16726 ( .A1(n15686), .A2(n16074), .ZN(n15693) );
  AOI21_X1 U16727 ( .B1(n15688), .B2(n16151), .A(n15687), .ZN(n15689) );
  OAI21_X1 U16728 ( .B1(n15690), .B2(n16096), .A(n15689), .ZN(n15691) );
  AOI21_X1 U16729 ( .B1(n15693), .B2(n15692), .A(n15691), .ZN(n15694) );
  OAI21_X1 U16730 ( .B1(n15732), .B2(n15695), .A(n15694), .ZN(n15751) );
  MUX2_X1 U16731 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15751), .S(n16179), .Z(
        P1_U3548) );
  INV_X1 U16732 ( .A(n15696), .ZN(n15697) );
  AOI21_X1 U16733 ( .B1(n15698), .B2(n16151), .A(n15697), .ZN(n15699) );
  OAI21_X1 U16734 ( .B1(n15700), .B2(n16096), .A(n15699), .ZN(n15701) );
  AOI21_X1 U16735 ( .B1(n15702), .B2(n15723), .A(n15701), .ZN(n15703) );
  OAI21_X1 U16736 ( .B1(n15704), .B2(n15732), .A(n15703), .ZN(n15752) );
  MUX2_X1 U16737 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15752), .S(n16179), .Z(
        P1_U3547) );
  AOI22_X1 U16738 ( .A1(n15706), .A2(n16153), .B1(n15705), .B2(n16151), .ZN(
        n15707) );
  OAI211_X1 U16739 ( .C1(n15709), .C2(n16116), .A(n15708), .B(n15707), .ZN(
        n15753) );
  MUX2_X1 U16740 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15753), .S(n16179), .Z(
        P1_U3546) );
  AOI21_X1 U16741 ( .B1(n15711), .B2(n16151), .A(n15710), .ZN(n15712) );
  OAI21_X1 U16742 ( .B1(n15713), .B2(n16096), .A(n15712), .ZN(n15714) );
  AOI21_X1 U16743 ( .B1(n15715), .B2(n16176), .A(n15714), .ZN(n15716) );
  OAI21_X1 U16744 ( .B1(n16074), .B2(n15717), .A(n15716), .ZN(n15754) );
  MUX2_X1 U16745 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15754), .S(n16179), .Z(
        P1_U3545) );
  AOI21_X1 U16746 ( .B1(n15719), .B2(n16151), .A(n15718), .ZN(n15720) );
  OAI21_X1 U16747 ( .B1(n15721), .B2(n16096), .A(n15720), .ZN(n15722) );
  AOI21_X1 U16748 ( .B1(n15724), .B2(n15723), .A(n15722), .ZN(n15725) );
  OAI21_X1 U16749 ( .B1(n15726), .B2(n15732), .A(n15725), .ZN(n15755) );
  MUX2_X1 U16750 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15755), .S(n16179), .Z(
        P1_U3544) );
  AOI211_X1 U16751 ( .C1(n15729), .C2(n16151), .A(n15728), .B(n15727), .ZN(
        n15730) );
  OAI21_X1 U16752 ( .B1(n15732), .B2(n15731), .A(n15730), .ZN(n15756) );
  MUX2_X1 U16753 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15756), .S(n16179), .Z(
        P1_U3543) );
  NAND2_X1 U16754 ( .A1(n15733), .A2(n16151), .ZN(n15734) );
  OAI211_X1 U16755 ( .C1(n15736), .C2(n16096), .A(n15735), .B(n15734), .ZN(
        n15737) );
  AOI21_X1 U16756 ( .B1(n15738), .B2(n16176), .A(n15737), .ZN(n15739) );
  OAI21_X1 U16757 ( .B1(n16074), .B2(n15740), .A(n15739), .ZN(n15757) );
  MUX2_X1 U16758 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15757), .S(n16179), .Z(
        P1_U3542) );
  MUX2_X1 U16759 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15741), .S(n16183), .Z(
        P1_U3527) );
  MUX2_X1 U16760 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15742), .S(n16183), .Z(
        P1_U3526) );
  MUX2_X1 U16761 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15744), .S(n16183), .Z(
        P1_U3523) );
  MUX2_X1 U16762 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15745), .S(n16183), .Z(
        P1_U3522) );
  MUX2_X1 U16763 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15746), .S(n16183), .Z(
        P1_U3521) );
  MUX2_X1 U16764 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15747), .S(n16183), .Z(
        P1_U3520) );
  MUX2_X1 U16765 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15748), .S(n16183), .Z(
        P1_U3519) );
  MUX2_X1 U16766 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15749), .S(n16183), .Z(
        P1_U3518) );
  MUX2_X1 U16767 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15750), .S(n16183), .Z(
        P1_U3517) );
  MUX2_X1 U16768 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15751), .S(n16183), .Z(
        P1_U3516) );
  MUX2_X1 U16769 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15752), .S(n16183), .Z(
        P1_U3515) );
  MUX2_X1 U16770 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15753), .S(n16183), .Z(
        P1_U3513) );
  MUX2_X1 U16771 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15754), .S(n16183), .Z(
        P1_U3510) );
  MUX2_X1 U16772 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15755), .S(n16183), .Z(
        P1_U3507) );
  MUX2_X1 U16773 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15756), .S(n16183), .Z(
        P1_U3504) );
  MUX2_X1 U16774 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15757), .S(n16183), .Z(
        P1_U3501) );
  INV_X1 U16775 ( .A(n15758), .ZN(n15762) );
  NOR4_X1 U16776 ( .A1(n15759), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8078), .A4(
        P1_U3086), .ZN(n15760) );
  AOI21_X1 U16777 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n15774), .A(n15760), 
        .ZN(n15761) );
  OAI21_X1 U16778 ( .B1(n15762), .B2(n15771), .A(n15761), .ZN(P1_U3324) );
  OAI222_X1 U16779 ( .A1(n15773), .A2(n15765), .B1(n7190), .B2(n15764), .C1(
        n15771), .C2(n15763), .ZN(P1_U3326) );
  OAI222_X1 U16780 ( .A1(n7190), .A2(n15768), .B1(n15771), .B2(n15767), .C1(
        n15766), .C2(n15773), .ZN(P1_U3329) );
  OAI222_X1 U16781 ( .A1(n15773), .A2(n15772), .B1(n15771), .B2(n15770), .C1(
        n7190), .C2(n15769), .ZN(P1_U3330) );
  NAND2_X1 U16782 ( .A1(n15774), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n15776) );
  OAI211_X1 U16783 ( .C1(n15777), .C2(n15771), .A(n15776), .B(n15775), .ZN(
        P1_U3332) );
  MUX2_X1 U16784 ( .A(n15779), .B(n15778), .S(n7190), .Z(P1_U3333) );
  MUX2_X1 U16785 ( .A(n15780), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16786 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15781) );
  NOR2_X1 U16787 ( .A1(n15811), .A2(n15781), .ZN(P1_U3323) );
  INV_X1 U16788 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15782) );
  NOR2_X1 U16789 ( .A1(n15811), .A2(n15782), .ZN(P1_U3322) );
  INV_X1 U16790 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15783) );
  NOR2_X1 U16791 ( .A1(n15811), .A2(n15783), .ZN(P1_U3321) );
  INV_X1 U16792 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15784) );
  NOR2_X1 U16793 ( .A1(n15811), .A2(n15784), .ZN(P1_U3320) );
  INV_X1 U16794 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15785) );
  NOR2_X1 U16795 ( .A1(n15811), .A2(n15785), .ZN(P1_U3319) );
  INV_X1 U16796 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15786) );
  NOR2_X1 U16797 ( .A1(n15811), .A2(n15786), .ZN(P1_U3318) );
  INV_X1 U16798 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15787) );
  NOR2_X1 U16799 ( .A1(n15811), .A2(n15787), .ZN(P1_U3317) );
  INV_X1 U16800 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15788) );
  NOR2_X1 U16801 ( .A1(n15811), .A2(n15788), .ZN(P1_U3316) );
  INV_X1 U16802 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15789) );
  NOR2_X1 U16803 ( .A1(n15811), .A2(n15789), .ZN(P1_U3315) );
  INV_X1 U16804 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15790) );
  NOR2_X1 U16805 ( .A1(n15811), .A2(n15790), .ZN(P1_U3314) );
  INV_X1 U16806 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15791) );
  NOR2_X1 U16807 ( .A1(n15811), .A2(n15791), .ZN(P1_U3313) );
  INV_X1 U16808 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15792) );
  NOR2_X1 U16809 ( .A1(n15811), .A2(n15792), .ZN(P1_U3312) );
  INV_X1 U16810 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15793) );
  NOR2_X1 U16811 ( .A1(n15811), .A2(n15793), .ZN(P1_U3311) );
  INV_X1 U16812 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15794) );
  NOR2_X1 U16813 ( .A1(n15811), .A2(n15794), .ZN(P1_U3310) );
  INV_X1 U16814 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15795) );
  NOR2_X1 U16815 ( .A1(n15811), .A2(n15795), .ZN(P1_U3309) );
  INV_X1 U16816 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15796) );
  NOR2_X1 U16817 ( .A1(n15811), .A2(n15796), .ZN(P1_U3308) );
  INV_X1 U16818 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15797) );
  NOR2_X1 U16819 ( .A1(n15811), .A2(n15797), .ZN(P1_U3307) );
  INV_X1 U16820 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15798) );
  NOR2_X1 U16821 ( .A1(n15811), .A2(n15798), .ZN(P1_U3306) );
  INV_X1 U16822 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15799) );
  NOR2_X1 U16823 ( .A1(n15811), .A2(n15799), .ZN(P1_U3305) );
  INV_X1 U16824 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15800) );
  NOR2_X1 U16825 ( .A1(n15811), .A2(n15800), .ZN(P1_U3304) );
  INV_X1 U16826 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15801) );
  NOR2_X1 U16827 ( .A1(n15811), .A2(n15801), .ZN(P1_U3303) );
  INV_X1 U16828 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15802) );
  NOR2_X1 U16829 ( .A1(n15811), .A2(n15802), .ZN(P1_U3302) );
  INV_X1 U16830 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15803) );
  NOR2_X1 U16831 ( .A1(n15811), .A2(n15803), .ZN(P1_U3301) );
  INV_X1 U16832 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15804) );
  NOR2_X1 U16833 ( .A1(n15811), .A2(n15804), .ZN(P1_U3300) );
  INV_X1 U16834 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15805) );
  NOR2_X1 U16835 ( .A1(n15811), .A2(n15805), .ZN(P1_U3299) );
  INV_X1 U16836 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15806) );
  NOR2_X1 U16837 ( .A1(n15811), .A2(n15806), .ZN(P1_U3298) );
  NOR2_X1 U16838 ( .A1(n15811), .A2(n15807), .ZN(P1_U3297) );
  NOR2_X1 U16839 ( .A1(n15811), .A2(n15808), .ZN(P1_U3296) );
  NOR2_X1 U16840 ( .A1(n15811), .A2(n15809), .ZN(P1_U3295) );
  NOR2_X1 U16841 ( .A1(n15811), .A2(n15810), .ZN(P1_U3294) );
  INV_X1 U16842 ( .A(n15812), .ZN(n15813) );
  AOI21_X1 U16843 ( .B1(n15814), .B2(n15818), .A(n15813), .ZN(P2_U3417) );
  AND2_X1 U16844 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15816), .ZN(P2_U3295) );
  AND2_X1 U16845 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15816), .ZN(P2_U3294) );
  AND2_X1 U16846 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15816), .ZN(P2_U3293) );
  AND2_X1 U16847 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15816), .ZN(P2_U3292) );
  AND2_X1 U16848 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15816), .ZN(P2_U3291) );
  AND2_X1 U16849 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15816), .ZN(P2_U3290) );
  AND2_X1 U16850 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15816), .ZN(P2_U3289) );
  AND2_X1 U16851 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15816), .ZN(P2_U3288) );
  AND2_X1 U16852 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15816), .ZN(P2_U3287) );
  AND2_X1 U16853 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15816), .ZN(P2_U3286) );
  AND2_X1 U16854 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15816), .ZN(P2_U3285) );
  AND2_X1 U16855 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15816), .ZN(P2_U3284) );
  AND2_X1 U16856 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15816), .ZN(P2_U3283) );
  AND2_X1 U16857 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15816), .ZN(P2_U3282) );
  AND2_X1 U16858 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15816), .ZN(P2_U3281) );
  AND2_X1 U16859 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15816), .ZN(P2_U3280) );
  AND2_X1 U16860 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15816), .ZN(P2_U3279) );
  AND2_X1 U16861 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15816), .ZN(P2_U3278) );
  AND2_X1 U16862 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15816), .ZN(P2_U3277) );
  AND2_X1 U16863 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15816), .ZN(P2_U3276) );
  AND2_X1 U16864 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15816), .ZN(P2_U3275) );
  AND2_X1 U16865 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15816), .ZN(P2_U3274) );
  AND2_X1 U16866 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15816), .ZN(P2_U3273) );
  AND2_X1 U16867 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15816), .ZN(P2_U3272) );
  AND2_X1 U16868 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15816), .ZN(P2_U3271) );
  AND2_X1 U16869 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15816), .ZN(P2_U3270) );
  AND2_X1 U16870 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15816), .ZN(P2_U3269) );
  AND2_X1 U16871 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15816), .ZN(P2_U3268) );
  AND2_X1 U16872 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15816), .ZN(P2_U3267) );
  AND2_X1 U16873 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15816), .ZN(P2_U3266) );
  NOR2_X1 U16874 ( .A1(n15858), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16875 ( .A1(P3_U3897), .A2(n15817), .ZN(P3_U3150) );
  INV_X1 U16876 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15819) );
  AOI22_X1 U16877 ( .A1(n15821), .A2(n15820), .B1(n15819), .B2(n15818), .ZN(
        P2_U3416) );
  NAND2_X1 U16878 ( .A1(n15892), .A2(n15822), .ZN(n15825) );
  INV_X1 U16879 ( .A(n15823), .ZN(n15824) );
  OAI211_X1 U16880 ( .C1(n15904), .C2(n15947), .A(n15825), .B(n15824), .ZN(
        n15826) );
  INV_X1 U16881 ( .A(n15826), .ZN(n15835) );
  OAI211_X1 U16882 ( .C1(n15829), .C2(n15828), .A(n15888), .B(n15827), .ZN(
        n15834) );
  OAI211_X1 U16883 ( .C1(n15832), .C2(n15831), .A(n15898), .B(n15830), .ZN(
        n15833) );
  NAND3_X1 U16884 ( .A1(n15835), .A2(n15834), .A3(n15833), .ZN(P2_U3219) );
  OAI22_X1 U16885 ( .A1(n15837), .A2(n15836), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14456), .ZN(n15838) );
  AOI21_X1 U16886 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n15858), .A(n15838), 
        .ZN(n15845) );
  OAI211_X1 U16887 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15840), .A(n15898), 
        .B(n15839), .ZN(n15844) );
  OAI211_X1 U16888 ( .C1(n15842), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15841), 
        .B(n15888), .ZN(n15843) );
  NAND3_X1 U16889 ( .A1(n15845), .A2(n15844), .A3(n15843), .ZN(P2_U3229) );
  AOI22_X1 U16890 ( .A1(n15858), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n15856) );
  OAI211_X1 U16891 ( .C1(n15848), .C2(n15847), .A(n15898), .B(n15846), .ZN(
        n15855) );
  NAND2_X1 U16892 ( .A1(n15849), .A2(n15892), .ZN(n15854) );
  OAI211_X1 U16893 ( .C1(n15852), .C2(n15851), .A(n15888), .B(n15850), .ZN(
        n15853) );
  NAND4_X1 U16894 ( .A1(n15856), .A2(n15855), .A3(n15854), .A4(n15853), .ZN(
        P2_U3230) );
  AOI22_X1 U16895 ( .A1(n15858), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n15871) );
  AOI211_X1 U16896 ( .C1(n15862), .C2(n15861), .A(n15860), .B(n15859), .ZN(
        n15863) );
  INV_X1 U16897 ( .A(n15863), .ZN(n15870) );
  NAND2_X1 U16898 ( .A1(n15892), .A2(n15864), .ZN(n15869) );
  XOR2_X1 U16899 ( .A(n15866), .B(n15865), .Z(n15867) );
  NAND2_X1 U16900 ( .A1(n15888), .A2(n15867), .ZN(n15868) );
  NAND4_X1 U16901 ( .A1(n15871), .A2(n15870), .A3(n15869), .A4(n15868), .ZN(
        P2_U3231) );
  OAI21_X1 U16902 ( .B1(n15874), .B2(n15873), .A(n15872), .ZN(n15883) );
  INV_X1 U16903 ( .A(n15875), .ZN(n15880) );
  NAND3_X1 U16904 ( .A1(n15878), .A2(n15877), .A3(n15876), .ZN(n15879) );
  NAND2_X1 U16905 ( .A1(n15880), .A2(n15879), .ZN(n15881) );
  AOI222_X1 U16906 ( .A1(n15883), .A2(n15888), .B1(n15882), .B2(n15892), .C1(
        n15881), .C2(n15898), .ZN(n15885) );
  OAI211_X1 U16907 ( .C1(n15968), .C2(n15904), .A(n15885), .B(n15884), .ZN(
        P2_U3226) );
  AND2_X1 U16908 ( .A1(n15887), .A2(n15886), .ZN(n15889) );
  OAI21_X1 U16909 ( .B1(n15890), .B2(n15889), .A(n15888), .ZN(n15901) );
  NAND2_X1 U16910 ( .A1(n15892), .A2(n15891), .ZN(n15900) );
  NAND2_X1 U16911 ( .A1(n15894), .A2(n15893), .ZN(n15895) );
  NAND2_X1 U16912 ( .A1(n15896), .A2(n15895), .ZN(n15897) );
  NAND2_X1 U16913 ( .A1(n15898), .A2(n15897), .ZN(n15899) );
  AND3_X1 U16914 ( .A1(n15901), .A2(n15900), .A3(n15899), .ZN(n15903) );
  OAI211_X1 U16915 ( .C1(n7441), .C2(n15904), .A(n15903), .B(n15902), .ZN(
        P2_U3223) );
  NOR2_X1 U16916 ( .A1(n15905), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15907) );
  OR2_X1 U16917 ( .A1(n15906), .A2(n15907), .ZN(n15910) );
  INV_X1 U16918 ( .A(n15907), .ZN(n15909) );
  MUX2_X1 U16919 ( .A(n15910), .B(n15909), .S(n15908), .Z(n15912) );
  NAND2_X1 U16920 ( .A1(n15912), .A2(n15911), .ZN(n15916) );
  AOI22_X1 U16921 ( .A1(n15914), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15915) );
  OAI21_X1 U16922 ( .B1(n15917), .B2(n15916), .A(n15915), .ZN(P1_U3243) );
  OAI21_X1 U16923 ( .B1(n15920), .B2(n15919), .A(n15918), .ZN(n15932) );
  MUX2_X1 U16924 ( .A(n10940), .B(P1_REG1_REG_12__SCAN_IN), .S(n15930), .Z(
        n15923) );
  INV_X1 U16925 ( .A(n15921), .ZN(n15922) );
  NAND2_X1 U16926 ( .A1(n15923), .A2(n15922), .ZN(n15925) );
  OAI21_X1 U16927 ( .B1(n15926), .B2(n15925), .A(n15924), .ZN(n15928) );
  AOI222_X1 U16928 ( .A1(n15932), .A2(n15931), .B1(n15930), .B2(n15929), .C1(
        n15928), .C2(n15927), .ZN(n15934) );
  OAI211_X1 U16929 ( .C1(n15936), .C2(n15935), .A(n15934), .B(n15933), .ZN(
        P1_U3255) );
  XOR2_X1 U16930 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15937), .Z(SUB_1596_U53) );
  AOI21_X1 U16931 ( .B1(n15940), .B2(n15939), .A(n15938), .ZN(SUB_1596_U61) );
  OAI21_X1 U16932 ( .B1(n15943), .B2(n15942), .A(n15941), .ZN(SUB_1596_U60) );
  AOI21_X1 U16933 ( .B1(n15945), .B2(n15944), .A(n7359), .ZN(SUB_1596_U59) );
  AOI21_X1 U16934 ( .B1(n15948), .B2(n15947), .A(n15946), .ZN(SUB_1596_U58) );
  AOI21_X1 U16935 ( .B1(n15951), .B2(n15950), .A(n15949), .ZN(SUB_1596_U56) );
  OAI21_X1 U16936 ( .B1(n15954), .B2(n15953), .A(n15952), .ZN(SUB_1596_U55) );
  AOI21_X1 U16937 ( .B1(n15957), .B2(n15956), .A(n15955), .ZN(n15958) );
  XOR2_X1 U16938 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n15958), .Z(SUB_1596_U54) );
  AOI21_X1 U16939 ( .B1(n15961), .B2(n15960), .A(n15959), .ZN(n15962) );
  XOR2_X1 U16940 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n15962), .Z(SUB_1596_U70)
         );
  AOI21_X1 U16941 ( .B1(n15965), .B2(n15964), .A(n15963), .ZN(n15966) );
  XOR2_X1 U16942 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15966), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16943 ( .B1(n15969), .B2(n15968), .A(n15967), .ZN(SUB_1596_U68) );
  OAI21_X1 U16944 ( .B1(n15972), .B2(n15971), .A(n15970), .ZN(n15973) );
  XNOR2_X1 U16945 ( .A(n15973), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16946 ( .B1(n15976), .B2(n15975), .A(n15974), .ZN(n15977) );
  XNOR2_X1 U16947 ( .A(n15977), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16948 ( .A1(n15982), .A2(n15981), .B1(n15982), .B2(n15980), .C1(
        n15979), .C2(n15978), .ZN(SUB_1596_U65) );
  OAI21_X1 U16949 ( .B1(n15985), .B2(n15984), .A(n15983), .ZN(n15986) );
  XNOR2_X1 U16950 ( .A(n15986), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  AOI21_X1 U16951 ( .B1(n15989), .B2(n15988), .A(n15987), .ZN(SUB_1596_U63) );
  AOI21_X1 U16952 ( .B1(n15994), .B2(n15993), .A(n15992), .ZN(n15995) );
  XOR2_X1 U16953 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n15995), .Z(SUB_1596_U57) );
  AOI21_X1 U16954 ( .B1(n15998), .B2(n15997), .A(n15996), .ZN(SUB_1596_U5) );
  INV_X1 U16955 ( .A(P2_RD_REG_SCAN_IN), .ZN(n16001) );
  OAI221_X1 U16956 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n16001), .C2(n16000), .A(n15999), .ZN(U29) );
  AOI21_X1 U16957 ( .B1(n16074), .B2(n16002), .A(n16012), .ZN(n16004) );
  NOR2_X1 U16958 ( .A1(n16004), .A2(n16003), .ZN(n16021) );
  INV_X1 U16959 ( .A(n16021), .ZN(n16007) );
  OAI22_X1 U16960 ( .A1(n16012), .A2(n16116), .B1(n16013), .B2(n16005), .ZN(
        n16006) );
  NOR2_X1 U16961 ( .A1(n16007), .A2(n16006), .ZN(n16010) );
  INV_X1 U16962 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n16008) );
  AOI22_X1 U16963 ( .A1(n16179), .A2(n16010), .B1(n16008), .B2(n16178), .ZN(
        P1_U3528) );
  INV_X1 U16964 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n16009) );
  AOI22_X1 U16965 ( .A1(n16183), .A2(n16010), .B1(n16009), .B2(n16180), .ZN(
        P1_U3459) );
  AOI22_X1 U16966 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n16011), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(n16022), .ZN(n16020) );
  INV_X1 U16967 ( .A(n16012), .ZN(n16017) );
  AOI21_X1 U16968 ( .B1(n16015), .B2(n16014), .A(n16013), .ZN(n16016) );
  AOI21_X1 U16969 ( .B1(n16018), .B2(n16017), .A(n16016), .ZN(n16019) );
  OAI211_X1 U16970 ( .C1(n16022), .C2(n16021), .A(n16020), .B(n16019), .ZN(
        P1_U3293) );
  AOI211_X1 U16971 ( .C1(n16226), .C2(n16025), .A(n16024), .B(n16023), .ZN(
        n16026) );
  AOI22_X1 U16972 ( .A1(n16228), .A2(n16026), .B1(n10484), .B2(n7687), .ZN(
        P3_U3460) );
  AOI22_X1 U16973 ( .A1(n16232), .A2(n16026), .B1(n8419), .B2(n16229), .ZN(
        P3_U3393) );
  OAI21_X1 U16974 ( .B1(n7707), .B2(n16028), .A(n16027), .ZN(n16049) );
  NOR2_X1 U16975 ( .A1(n16029), .A2(n16222), .ZN(n16043) );
  XNOR2_X1 U16976 ( .A(n16030), .B(n7707), .ZN(n16038) );
  OAI22_X1 U16977 ( .A1(n16035), .A2(n16034), .B1(n16033), .B2(n16032), .ZN(
        n16036) );
  AOI21_X1 U16978 ( .B1(n16049), .B2(n16212), .A(n16036), .ZN(n16037) );
  OAI21_X1 U16979 ( .B1(n16039), .B2(n16038), .A(n16037), .ZN(n16047) );
  AOI211_X1 U16980 ( .C1(n16213), .C2(n16049), .A(n16043), .B(n16047), .ZN(
        n16042) );
  OR2_X1 U16981 ( .A1(n16042), .A2(n7687), .ZN(n16040) );
  OAI21_X1 U16982 ( .B1(n16228), .B2(n10487), .A(n16040), .ZN(P3_U3461) );
  INV_X1 U16983 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n16041) );
  AOI22_X1 U16984 ( .A1(n16232), .A2(n16042), .B1(n16041), .B2(n16229), .ZN(
        P3_U3396) );
  INV_X1 U16985 ( .A(n16043), .ZN(n16046) );
  OAI22_X1 U16986 ( .A1(n16046), .A2(n16045), .B1(n16128), .B2(n16044), .ZN(
        n16048) );
  AOI211_X1 U16987 ( .C1(n16050), .C2(n16049), .A(n16048), .B(n16047), .ZN(
        n16051) );
  AOI22_X1 U16988 ( .A1(n16052), .A2(n10488), .B1(n16051), .B2(n16131), .ZN(
        P3_U3231) );
  AOI22_X1 U16989 ( .A1(n16055), .A2(n16226), .B1(n16054), .B2(n16053), .ZN(
        n16057) );
  AND2_X1 U16990 ( .A1(n16057), .A2(n16056), .ZN(n16059) );
  AOI22_X1 U16991 ( .A1(n16228), .A2(n16059), .B1(n10493), .B2(n7687), .ZN(
        P3_U3462) );
  INV_X1 U16992 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n16058) );
  AOI22_X1 U16993 ( .A1(n16232), .A2(n16059), .B1(n16058), .B2(n16229), .ZN(
        P3_U3399) );
  AOI22_X1 U16994 ( .A1(n16082), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n16080), 
        .B2(n16060), .ZN(n16061) );
  OAI21_X1 U16995 ( .B1(n16085), .B2(n7910), .A(n16061), .ZN(n16065) );
  NOR2_X1 U16996 ( .A1(n16063), .A2(n16062), .ZN(n16064) );
  AOI211_X1 U16997 ( .C1(n16066), .C2(n16088), .A(n16065), .B(n16064), .ZN(
        n16067) );
  OAI21_X1 U16998 ( .B1(n16094), .B2(n16068), .A(n16067), .ZN(P2_U3262) );
  OAI21_X1 U16999 ( .B1(n16070), .B2(n16171), .A(n16069), .ZN(n16071) );
  AOI21_X1 U17000 ( .B1(n16072), .B2(n16153), .A(n16071), .ZN(n16073) );
  OAI21_X1 U17001 ( .B1(n16075), .B2(n16074), .A(n16073), .ZN(n16076) );
  AOI21_X1 U17002 ( .B1(n16077), .B2(n16176), .A(n16076), .ZN(n16079) );
  AOI22_X1 U17003 ( .A1(n16179), .A2(n16079), .B1(n10302), .B2(n16178), .ZN(
        P1_U3532) );
  INV_X1 U17004 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n16078) );
  AOI22_X1 U17005 ( .A1(n16183), .A2(n16079), .B1(n16078), .B2(n16180), .ZN(
        P1_U3471) );
  AOI22_X1 U17006 ( .A1(n16082), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n16081), 
        .B2(n16080), .ZN(n16083) );
  OAI21_X1 U17007 ( .B1(n16085), .B2(n16084), .A(n16083), .ZN(n16086) );
  INV_X1 U17008 ( .A(n16086), .ZN(n16092) );
  AOI22_X1 U17009 ( .A1(n16090), .A2(n16089), .B1(n16088), .B2(n16087), .ZN(
        n16091) );
  OAI211_X1 U17010 ( .C1(n16094), .C2(n16093), .A(n16092), .B(n16091), .ZN(
        P2_U3261) );
  INV_X1 U17011 ( .A(n16116), .ZN(n16149) );
  OAI22_X1 U17012 ( .A1(n16097), .A2(n16096), .B1(n16095), .B2(n16171), .ZN(
        n16100) );
  INV_X1 U17013 ( .A(n16098), .ZN(n16099) );
  AOI211_X1 U17014 ( .C1(n16149), .C2(n16101), .A(n16100), .B(n16099), .ZN(
        n16103) );
  AOI22_X1 U17015 ( .A1(n16179), .A2(n16103), .B1(n10305), .B2(n16178), .ZN(
        P1_U3533) );
  INV_X1 U17016 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n16102) );
  AOI22_X1 U17017 ( .A1(n16183), .A2(n16103), .B1(n16102), .B2(n16180), .ZN(
        P1_U3474) );
  AOI21_X1 U17018 ( .B1(n16123), .B2(n16105), .A(n16104), .ZN(n16107) );
  OAI222_X1 U17019 ( .A1(n16108), .A2(n16126), .B1(n16052), .B2(n16107), .C1(
        n16128), .C2(n16106), .ZN(n16109) );
  INV_X1 U17020 ( .A(n16109), .ZN(n16110) );
  OAI21_X1 U17021 ( .B1(n16131), .B2(n10659), .A(n16110), .ZN(P3_U3226) );
  AOI22_X1 U17022 ( .A1(n16112), .A2(n16153), .B1(n16111), .B2(n16151), .ZN(
        n16113) );
  OAI211_X1 U17023 ( .C1(n16116), .C2(n16115), .A(n16114), .B(n16113), .ZN(
        n16117) );
  INV_X1 U17024 ( .A(n16117), .ZN(n16120) );
  AOI22_X1 U17025 ( .A1(n16179), .A2(n16120), .B1(n16118), .B2(n16178), .ZN(
        P1_U3535) );
  INV_X1 U17026 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n16119) );
  AOI22_X1 U17027 ( .A1(n16183), .A2(n16120), .B1(n16119), .B2(n16180), .ZN(
        P1_U3480) );
  AOI21_X1 U17028 ( .B1(n16123), .B2(n16122), .A(n16121), .ZN(n16124) );
  OAI222_X1 U17029 ( .A1(n16128), .A2(n16127), .B1(n16126), .B2(n16125), .C1(
        n16052), .C2(n16124), .ZN(n16129) );
  INV_X1 U17030 ( .A(n16129), .ZN(n16130) );
  OAI21_X1 U17031 ( .B1(n16131), .B2(n10806), .A(n16130), .ZN(P3_U3225) );
  AOI21_X1 U17032 ( .B1(n16134), .B2(n16133), .A(n16132), .ZN(n16135) );
  OAI211_X1 U17033 ( .C1(n16138), .C2(n16137), .A(n16136), .B(n16135), .ZN(
        n16139) );
  INV_X1 U17034 ( .A(n16139), .ZN(n16141) );
  AOI22_X1 U17035 ( .A1(n16208), .A2(n16141), .B1(n10919), .B2(n16206), .ZN(
        P2_U3507) );
  INV_X1 U17036 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n16140) );
  AOI22_X1 U17037 ( .A1(n14948), .A2(n16141), .B1(n16140), .B2(n16209), .ZN(
        P2_U3454) );
  OAI22_X1 U17038 ( .A1(n16143), .A2(n16163), .B1(n16222), .B2(n16142), .ZN(
        n16144) );
  NOR2_X1 U17039 ( .A1(n16145), .A2(n16144), .ZN(n16148) );
  AOI22_X1 U17040 ( .A1(n16228), .A2(n16148), .B1(n16146), .B2(n7687), .ZN(
        P3_U3468) );
  INV_X1 U17041 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16147) );
  AOI22_X1 U17042 ( .A1(n16232), .A2(n16148), .B1(n16147), .B2(n16229), .ZN(
        P3_U3417) );
  NAND2_X1 U17043 ( .A1(n16150), .A2(n16149), .ZN(n16156) );
  AOI22_X1 U17044 ( .A1(n16154), .A2(n16153), .B1(n16152), .B2(n16151), .ZN(
        n16155) );
  NAND2_X1 U17045 ( .A1(n16156), .A2(n16155), .ZN(n16157) );
  NOR2_X1 U17046 ( .A1(n16158), .A2(n16157), .ZN(n16161) );
  AOI22_X1 U17047 ( .A1(n16179), .A2(n16161), .B1(n16159), .B2(n16178), .ZN(
        P1_U3537) );
  INV_X1 U17048 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n16160) );
  AOI22_X1 U17049 ( .A1(n16183), .A2(n16161), .B1(n16160), .B2(n16180), .ZN(
        P1_U3486) );
  OAI22_X1 U17050 ( .A1(n16164), .A2(n16163), .B1(n16222), .B2(n16162), .ZN(
        n16165) );
  NOR2_X1 U17051 ( .A1(n16166), .A2(n16165), .ZN(n16167) );
  AOI22_X1 U17052 ( .A1(n16228), .A2(n16167), .B1(n11561), .B2(n7687), .ZN(
        P3_U3469) );
  AOI22_X1 U17053 ( .A1(n16232), .A2(n16167), .B1(n9511), .B2(n16229), .ZN(
        P3_U3420) );
  INV_X1 U17054 ( .A(n16168), .ZN(n16177) );
  OAI211_X1 U17055 ( .C1(n16172), .C2(n16171), .A(n16170), .B(n16169), .ZN(
        n16175) );
  INV_X1 U17056 ( .A(n16173), .ZN(n16174) );
  AOI211_X1 U17057 ( .C1(n16177), .C2(n16176), .A(n16175), .B(n16174), .ZN(
        n16182) );
  AOI22_X1 U17058 ( .A1(n16179), .A2(n16182), .B1(n10578), .B2(n16178), .ZN(
        P1_U3538) );
  INV_X1 U17059 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n16181) );
  AOI22_X1 U17060 ( .A1(n16183), .A2(n16182), .B1(n16181), .B2(n16180), .ZN(
        P1_U3489) );
  INV_X1 U17061 ( .A(n16184), .ZN(n16189) );
  OAI21_X1 U17062 ( .B1(n16186), .B2(n16201), .A(n16185), .ZN(n16188) );
  AOI22_X1 U17063 ( .A1(n16208), .A2(n16192), .B1(n10923), .B2(n16206), .ZN(
        P2_U3509) );
  INV_X1 U17064 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n16191) );
  AOI22_X1 U17065 ( .A1(n14948), .A2(n16192), .B1(n16191), .B2(n16209), .ZN(
        P2_U3460) );
  NOR2_X1 U17066 ( .A1(n16193), .A2(n16222), .ZN(n16195) );
  AOI211_X1 U17067 ( .C1(n16226), .C2(n16196), .A(n16195), .B(n16194), .ZN(
        n16198) );
  AOI22_X1 U17068 ( .A1(n16228), .A2(n16198), .B1(n9533), .B2(n7687), .ZN(
        P3_U3470) );
  INV_X1 U17069 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16197) );
  AOI22_X1 U17070 ( .A1(n16232), .A2(n16198), .B1(n16197), .B2(n16229), .ZN(
        P3_U3423) );
  OAI211_X1 U17071 ( .C1(n16202), .C2(n16201), .A(n16200), .B(n16199), .ZN(
        n16203) );
  AOI21_X1 U17072 ( .B1(n16205), .B2(n16204), .A(n16203), .ZN(n16211) );
  AOI22_X1 U17073 ( .A1(n16208), .A2(n16211), .B1(n16207), .B2(n16206), .ZN(
        P2_U3511) );
  INV_X1 U17074 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n16210) );
  AOI22_X1 U17075 ( .A1(n14948), .A2(n16211), .B1(n16210), .B2(n16209), .ZN(
        P2_U3466) );
  NAND2_X1 U17076 ( .A1(n16214), .A2(n16212), .ZN(n16216) );
  NAND2_X1 U17077 ( .A1(n16214), .A2(n16213), .ZN(n16215) );
  OAI211_X1 U17078 ( .C1(n16217), .C2(n16222), .A(n16216), .B(n16215), .ZN(
        n16218) );
  NOR2_X1 U17079 ( .A1(n16219), .A2(n16218), .ZN(n16221) );
  AOI22_X1 U17080 ( .A1(n16228), .A2(n16221), .B1(n9571), .B2(n7687), .ZN(
        P3_U3472) );
  INV_X1 U17081 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n16220) );
  AOI22_X1 U17082 ( .A1(n16232), .A2(n16221), .B1(n16220), .B2(n16229), .ZN(
        P3_U3429) );
  NOR2_X1 U17083 ( .A1(n16223), .A2(n16222), .ZN(n16225) );
  AOI211_X1 U17084 ( .C1(n16227), .C2(n16226), .A(n16225), .B(n16224), .ZN(
        n16231) );
  AOI22_X1 U17085 ( .A1(n16228), .A2(n16231), .B1(n9587), .B2(n7687), .ZN(
        P3_U3473) );
  INV_X1 U17086 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n16230) );
  AOI22_X1 U17087 ( .A1(n16232), .A2(n16231), .B1(n16230), .B2(n16229), .ZN(
        P3_U3432) );
  AOI21_X1 U17088 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16233) );
  OAI21_X1 U17089 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16233), 
        .ZN(U28) );
  AND2_X1 U7342 ( .A1(n15585), .A2(n15370), .ZN(n15566) );
  CLKBUF_X1 U8727 ( .A(n10410), .Z(n16153) );
endmodule

