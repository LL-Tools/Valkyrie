

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601;

  NAND2_X1 U4916 ( .A1(n6840), .A2(n6692), .ZN(n8633) );
  AND2_X1 U4917 ( .A1(n8295), .A2(n5043), .ZN(n8593) );
  AND2_X1 U4918 ( .A1(n10173), .A2(n8225), .ZN(n8213) );
  NAND2_X1 U4919 ( .A1(n6212), .A2(n6211), .ZN(n10028) );
  CLKBUF_X2 U4920 ( .A(n5848), .Z(n7033) );
  NAND2_X1 U4921 ( .A1(n4553), .A2(n6798), .ZN(n10170) );
  AND2_X1 U4922 ( .A1(n6718), .A2(n6719), .ZN(n8002) );
  AND2_X2 U4923 ( .A1(n6251), .A2(n6250), .ZN(n6260) );
  CLKBUF_X2 U4924 ( .A(n6606), .Z(n4414) );
  INV_X1 U4925 ( .A(n6284), .ZN(n6586) );
  CLKBUF_X2 U4926 ( .A(n6606), .Z(n4415) );
  NAND4_X1 U4927 ( .A1(n6255), .A2(n6254), .A3(n6253), .A4(n6252), .ZN(n9624)
         );
  BUF_X1 U4928 ( .A(n5733), .Z(n4726) );
  INV_X2 U4929 ( .A(n6913), .ZN(n5653) );
  NAND2_X1 U4930 ( .A1(n4997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6653) );
  NAND4_X1 U4931 ( .A1(n4958), .A2(n4960), .A3(n4957), .A4(n4956), .ZN(n5270)
         );
  INV_X1 U4932 ( .A(n10438), .ZN(n4409) );
  INV_X2 U4933 ( .A(n4409), .ZN(n4410) );
  INV_X1 U4934 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n10438) );
  MUX2_X1 U4935 ( .A(n6349), .B(n6348), .S(n10210), .Z(n6350) );
  OAI21_X1 U4936 ( .B1(n6542), .B2(n6541), .A(n6540), .ZN(n6552) );
  OAI21_X1 U4937 ( .B1(n6656), .B2(n6655), .A(n6806), .ZN(n6767) );
  INV_X1 U4938 ( .A(n7058), .ZN(n7304) );
  INV_X1 U4939 ( .A(n7058), .ZN(n7274) );
  NAND2_X1 U4940 ( .A1(n8341), .A2(n4490), .ZN(n8585) );
  OAI21_X1 U4941 ( .B1(n7378), .B2(n5324), .A(n5048), .ZN(n5326) );
  OR2_X1 U4942 ( .A1(n5733), .A2(n4666), .ZN(n5300) );
  NAND2_X1 U4943 ( .A1(n7899), .A2(n9248), .ZN(n7819) );
  BUF_X1 U4944 ( .A(n7286), .Z(n4420) );
  AND2_X1 U4945 ( .A1(n6755), .A2(n6844), .ZN(n7346) );
  NAND2_X1 U4946 ( .A1(n9842), .A2(n9843), .ZN(n9841) );
  INV_X1 U4947 ( .A(n6791), .ZN(n8140) );
  AND2_X1 U4949 ( .A1(n7762), .A2(n6100), .ZN(n9203) );
  INV_X1 U4950 ( .A(n8911), .ZN(n8118) );
  NAND2_X1 U4951 ( .A1(n4812), .A2(n5298), .ZN(n9248) );
  INV_X1 U4953 ( .A(n9844), .ZN(n9827) );
  INV_X1 U4954 ( .A(n9621), .ZN(n8005) );
  XNOR2_X1 U4955 ( .A(n6061), .B(n6060), .ZN(n6063) );
  NAND2_X1 U4956 ( .A1(n6136), .A2(n6135), .ZN(n6893) );
  NAND2_X2 U4957 ( .A1(n5401), .A2(n5400), .ZN(n8121) );
  NAND2_X1 U4958 ( .A1(n5373), .A2(n5372), .ZN(n10238) );
  INV_X1 U4959 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5331) );
  OAI21_X1 U4960 ( .B1(n7067), .B2(n7068), .A(n7684), .ZN(n7652) );
  AND2_X1 U4961 ( .A1(n6197), .A2(n6196), .ZN(n9587) );
  NAND2_X1 U4962 ( .A1(n6775), .A2(n6842), .ZN(n9826) );
  MUX2_X1 U4963 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10071), .S(n10225), .Z(
        n9991) );
  MUX2_X1 U4964 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10071), .S(n10218), .Z(
        n10072) );
  NAND2_X1 U4965 ( .A1(n6641), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6642) );
  OR3_X1 U4966 ( .A1(n9796), .A2(n9795), .A3(n9971), .ZN(n9990) );
  OAI21_X1 U4967 ( .B1(n10267), .B2(n10271), .A(n10269), .ZN(n10596) );
  OAI21_X2 U4970 ( .B1(n8585), .B2(n4838), .A(n4678), .ZN(n9950) );
  NAND2_X2 U4971 ( .A1(n7153), .A2(n7154), .ZN(n5011) );
  NAND2_X2 U4972 ( .A1(n7152), .A2(n7151), .ZN(n7155) );
  XNOR2_X2 U4973 ( .A(n10144), .B(n10499), .ZN(n10593) );
  INV_X1 U4974 ( .A(n9240), .ZN(n7913) );
  NAND4_X2 U4975 ( .A1(n5315), .A2(n5314), .A3(n5313), .A4(n5312), .ZN(n9240)
         );
  NAND2_X1 U4976 ( .A1(n6938), .A2(n5848), .ZN(n4412) );
  NAND2_X2 U4977 ( .A1(n10142), .A2(n10143), .ZN(n10144) );
  NAND2_X2 U4978 ( .A1(n6445), .A2(n6444), .ZN(n10058) );
  OAI21_X4 U4979 ( .B1(n5723), .B2(n5722), .A(n5721), .ZN(n5741) );
  OAI21_X2 U4980 ( .B1(n5640), .B2(n5077), .A(n5073), .ZN(n5723) );
  NAND2_X1 U4981 ( .A1(n6009), .A2(n9179), .ZN(n6018) );
  OR2_X2 U4982 ( .A1(n6298), .A2(n5357), .ZN(n5401) );
  NAND3_X2 U4983 ( .A1(n5139), .A2(n6825), .A3(n5138), .ZN(n8625) );
  OAI222_X1 U4984 ( .A1(n10118), .A2(n8662), .B1(n4410), .B2(n8661), .C1(n9417), .C2(n10121), .ZN(P1_U3326) );
  NAND2_X2 U4985 ( .A1(n6309), .A2(n6308), .ZN(n7105) );
  AOI21_X2 U4986 ( .B1(n7351), .B2(n10163), .A(n7350), .ZN(n8637) );
  OAI21_X2 U4987 ( .B1(n6555), .B2(n4440), .A(n4883), .ZN(n6595) );
  INV_X2 U4988 ( .A(n5185), .ZN(n7756) );
  XNOR2_X2 U4989 ( .A(n5399), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6992) );
  AOI21_X2 U4990 ( .B1(n8847), .B2(n8848), .A(n4441), .ZN(n8821) );
  NAND2_X2 U4991 ( .A1(n8708), .A2(n8707), .ZN(n8847) );
  XNOR2_X2 U4992 ( .A(n5680), .B(n5679), .ZN(n8285) );
  NAND2_X2 U4993 ( .A1(n4782), .A2(n5079), .ZN(n5680) );
  XNOR2_X2 U4995 ( .A(n6276), .B(P1_IR_REG_2__SCAN_IN), .ZN(n7582) );
  NAND2_X2 U4996 ( .A1(n5730), .A2(n5729), .ZN(n9344) );
  NOR2_X2 U4997 ( .A1(n8118), .A2(n10238), .ZN(n8054) );
  XOR2_X2 U4998 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10147), .Z(n10594) );
  NAND2_X2 U4999 ( .A1(n10146), .A2(n10145), .ZN(n10147) );
  XNOR2_X2 U5000 ( .A(n5279), .B(n5278), .ZN(n6938) );
  NOR2_X2 U5001 ( .A1(n8633), .A2(n6838), .ZN(n6839) );
  XNOR2_X2 U5002 ( .A(n6642), .B(n6643), .ZN(n6856) );
  NAND2_X2 U5003 ( .A1(n6301), .A2(n6300), .ZN(n10210) );
  INV_X1 U5004 ( .A(n6884), .ZN(n6894) );
  NAND2_X1 U5005 ( .A1(n4667), .A2(n6016), .ZN(n9123) );
  NAND2_X1 U5006 ( .A1(n8668), .A2(n8667), .ZN(n8739) );
  NAND2_X1 U5007 ( .A1(n6581), .A2(n6580), .ZN(n9998) );
  NAND2_X1 U5008 ( .A1(n6570), .A2(n6569), .ZN(n10004) );
  NAND2_X1 U5009 ( .A1(n8115), .A2(n5128), .ZN(n8252) );
  OR2_X1 U5010 ( .A1(n6928), .A2(n8271), .ZN(n4980) );
  NAND2_X1 U5011 ( .A1(n8342), .A2(n4787), .ZN(n8341) );
  INV_X2 U5012 ( .A(n7919), .ZN(n7911) );
  NAND2_X1 U5013 ( .A1(n5556), .A2(n5555), .ZN(n5575) );
  NAND2_X1 U5014 ( .A1(n8020), .A2(n7960), .ZN(n5972) );
  INV_X1 U5015 ( .A(n7847), .ZN(n7850) );
  NAND2_X1 U5016 ( .A1(n7976), .A2(n7913), .ZN(n7904) );
  INV_X2 U5017 ( .A(n7170), .ZN(n7230) );
  INV_X1 U5018 ( .A(n8742), .ZN(n8397) );
  BUF_X1 U5019 ( .A(n7286), .Z(n4421) );
  INV_X1 U5020 ( .A(n9224), .ZN(n8789) );
  INV_X4 U5021 ( .A(n7277), .ZN(n7301) );
  INV_X2 U5022 ( .A(n8020), .ZN(n5157) );
  INV_X1 U5023 ( .A(n9622), .ZN(n8006) );
  INV_X1 U5024 ( .A(n6792), .ZN(n6793) );
  CLKBUF_X3 U5025 ( .A(n7049), .Z(n7369) );
  INV_X8 U5026 ( .A(n6910), .ZN(n6100) );
  NOR2_X1 U5027 ( .A1(n9624), .A2(n6853), .ZN(n8139) );
  CLKBUF_X2 U5028 ( .A(n6259), .Z(n6792) );
  NAND2_X2 U5029 ( .A1(n9781), .A2(n8505), .ZN(n6834) );
  CLKBUF_X1 U5030 ( .A(n7046), .Z(n4422) );
  CLKBUF_X1 U5031 ( .A(n6284), .Z(n6619) );
  INV_X1 U5032 ( .A(n6263), .ZN(n4417) );
  INV_X1 U5033 ( .A(n5544), .ZN(n5842) );
  NAND2_X1 U5034 ( .A1(n6174), .A2(n6175), .ZN(n6282) );
  NAND2_X1 U5035 ( .A1(n6645), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6649) );
  AND2_X2 U5036 ( .A1(n4565), .A2(n4564), .ZN(n5347) );
  INV_X2 U5037 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5267) );
  INV_X1 U5038 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4551) );
  NOR2_X1 U5039 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6367) );
  NAND2_X1 U5040 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6311) );
  INV_X1 U5041 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6648) );
  AOI21_X1 U5042 ( .B1(n8794), .B2(n8795), .A(n5108), .ZN(n8879) );
  NAND2_X1 U5043 ( .A1(n5112), .A2(n8714), .ZN(n8794) );
  NAND2_X1 U5044 ( .A1(n5099), .A2(n5096), .ZN(n8761) );
  NOR2_X1 U5045 ( .A1(n4805), .A2(n4616), .ZN(n10076) );
  NAND2_X1 U5046 ( .A1(n4480), .A2(n4854), .ZN(n4805) );
  XNOR2_X1 U5047 ( .A(n6893), .B(n6894), .ZN(n9035) );
  OAI21_X1 U5048 ( .B1(n9530), .B2(n4560), .A(n4477), .ZN(n4559) );
  AOI21_X1 U5049 ( .B1(n9434), .B2(n4695), .A(n4479), .ZN(n4694) );
  AND2_X1 U5050 ( .A1(n9580), .A2(n5026), .ZN(n9434) );
  AND2_X1 U5051 ( .A1(n4563), .A2(n4562), .ZN(n9530) );
  NAND2_X1 U5052 ( .A1(n9803), .A2(n9804), .ZN(n9802) );
  AND2_X1 U5053 ( .A1(n9995), .A2(n10206), .ZN(n4616) );
  AOI21_X1 U5054 ( .B1(n8621), .B2(n10163), .A(n4713), .ZN(n10000) );
  NAND2_X1 U5055 ( .A1(n4657), .A2(n4655), .ZN(n10006) );
  NAND2_X1 U5056 ( .A1(n9562), .A2(n9560), .ZN(n9559) );
  AOI21_X1 U5057 ( .B1(n5228), .B2(n5230), .A(n5227), .ZN(n5226) );
  AND2_X1 U5058 ( .A1(n8615), .A2(n6829), .ZN(n9812) );
  CLKBUF_X1 U5059 ( .A(n8813), .Z(n4596) );
  MUX2_X1 U5060 ( .A(n9783), .B(n9782), .S(n9781), .Z(n9785) );
  NAND2_X1 U5061 ( .A1(n7239), .A2(n7238), .ZN(n9478) );
  INV_X1 U5062 ( .A(n9994), .ZN(n4854) );
  AOI21_X1 U5063 ( .B1(n4848), .B2(n4851), .A(n4846), .ZN(n4845) );
  NAND2_X1 U5064 ( .A1(n4595), .A2(n4523), .ZN(n10070) );
  NAND2_X1 U5065 ( .A1(n9096), .A2(n9097), .ZN(n5181) );
  OR2_X1 U5066 ( .A1(n9412), .A2(n7378), .ZN(n4595) );
  NAND2_X1 U5067 ( .A1(n6161), .A2(n6160), .ZN(n7352) );
  INV_X1 U5068 ( .A(n8616), .ZN(n4416) );
  XNOR2_X1 U5069 ( .A(n6081), .B(n6080), .ZN(n8610) );
  OAI21_X1 U5070 ( .B1(n8739), .B2(n5121), .A(n5118), .ZN(n8685) );
  OAI21_X1 U5071 ( .B1(n6063), .B2(n10526), .A(n6062), .ZN(n6081) );
  NAND2_X1 U5072 ( .A1(n5819), .A2(n5818), .ZN(n9261) );
  XNOR2_X1 U5073 ( .A(n6063), .B(SI_29_), .ZN(n8660) );
  NAND2_X1 U5074 ( .A1(n5802), .A2(n5801), .ZN(n9327) );
  NAND2_X1 U5075 ( .A1(n6190), .A2(n6189), .ZN(n9816) );
  NAND2_X1 U5076 ( .A1(n9958), .A2(n4548), .ZN(n4799) );
  XNOR2_X1 U5077 ( .A(n5817), .B(n5934), .ZN(n9419) );
  AND2_X1 U5078 ( .A1(n5937), .A2(n5935), .ZN(n5817) );
  NAND2_X1 U5079 ( .A1(n4554), .A2(n6812), .ZN(n9969) );
  AOI21_X1 U5080 ( .B1(n9884), .B2(n4842), .A(n4841), .ZN(n4840) );
  NAND2_X1 U5081 ( .A1(n8252), .A2(n5127), .ZN(n8393) );
  NAND2_X1 U5082 ( .A1(n6558), .A2(n6557), .ZN(n10008) );
  NAND2_X1 U5083 ( .A1(n5672), .A2(n5671), .ZN(n9356) );
  NAND2_X1 U5084 ( .A1(n6235), .A2(n6234), .ZN(n9876) );
  CLKBUF_X1 U5085 ( .A(n9193), .Z(n4625) );
  XNOR2_X1 U5086 ( .A(n10028), .B(n9615), .ZN(n9884) );
  OAI21_X1 U5087 ( .B1(n5492), .B2(n5168), .A(n5164), .ZN(n9187) );
  NAND2_X1 U5088 ( .A1(n6530), .A2(n6529), .ZN(n10011) );
  NAND2_X1 U5089 ( .A1(n5682), .A2(n5681), .ZN(n9124) );
  AND2_X1 U5090 ( .A1(n9475), .A2(n9616), .ZN(n4426) );
  XNOR2_X1 U5091 ( .A(n5758), .B(n5757), .ZN(n8600) );
  NAND2_X1 U5092 ( .A1(n5655), .A2(n5654), .ZN(n9365) );
  NOR2_X1 U5093 ( .A1(n5123), .A2(n8840), .ZN(n5122) );
  AOI21_X1 U5094 ( .B1(n7948), .B2(n8096), .A(n8097), .ZN(n8095) );
  NAND2_X1 U5095 ( .A1(n6221), .A2(n6220), .ZN(n9475) );
  AND4_X1 U5096 ( .A1(n5998), .A2(n6100), .A3(n5997), .A4(n6111), .ZN(n4913)
         );
  NAND2_X1 U5097 ( .A1(n6504), .A2(n6503), .ZN(n10038) );
  AOI21_X1 U5098 ( .B1(n8676), .B2(n8677), .A(n4456), .ZN(n5125) );
  AND2_X1 U5099 ( .A1(n6005), .A2(n6006), .ZN(n9194) );
  NAND2_X1 U5100 ( .A1(n5617), .A2(n5616), .ZN(n9376) );
  NAND2_X1 U5101 ( .A1(n6492), .A2(n6491), .ZN(n10043) );
  NAND2_X1 U5102 ( .A1(n6169), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U5103 ( .A1(n8516), .A2(n9979), .ZN(n6735) );
  AND2_X1 U5104 ( .A1(n6736), .A2(n9947), .ZN(n9977) );
  NAND2_X1 U5105 ( .A1(n8082), .A2(n5983), .ZN(n8048) );
  OAI21_X1 U5106 ( .B1(n5640), .B2(n5083), .A(n5643), .ZN(n5666) );
  NAND2_X1 U5107 ( .A1(n7812), .A2(n7813), .ZN(n7890) );
  NAND2_X2 U5108 ( .A1(n6467), .A2(n6466), .ZN(n10052) );
  NOR2_X1 U5109 ( .A1(n4754), .A2(n4753), .ZN(n4898) );
  NAND2_X1 U5110 ( .A1(n5580), .A2(n5579), .ZN(n9388) );
  NAND2_X1 U5111 ( .A1(n5564), .A2(n5563), .ZN(n9394) );
  NAND2_X1 U5112 ( .A1(n6458), .A2(n6457), .ZN(n9961) );
  NAND2_X1 U5113 ( .A1(n5600), .A2(n5599), .ZN(n9382) );
  NAND2_X1 U5114 ( .A1(n4446), .A2(n5607), .ZN(n5057) );
  NAND2_X1 U5115 ( .A1(n5538), .A2(n5537), .ZN(n9400) );
  NAND2_X1 U5116 ( .A1(n5962), .A2(n8053), .ZN(n5973) );
  OAI21_X1 U5117 ( .B1(n10170), .B2(n6800), .A(n6799), .ZN(n8000) );
  NAND2_X1 U5118 ( .A1(n6398), .A2(n6397), .ZN(n8490) );
  OR2_X1 U5119 ( .A1(n10210), .A2(n8005), .ZN(n6763) );
  NOR2_X1 U5120 ( .A1(n7636), .A2(n6923), .ZN(n6924) );
  NAND2_X1 U5121 ( .A1(n8121), .A2(n8256), .ZN(n5962) );
  NAND2_X1 U5122 ( .A1(n5550), .A2(n5549), .ZN(n5556) );
  AOI21_X1 U5123 ( .B1(n7634), .B2(n7632), .A(n7633), .ZN(n7636) );
  AND2_X2 U5124 ( .A1(n8134), .A2(n9962), .ZN(n10167) );
  NAND3_X1 U5125 ( .A1(n4983), .A2(P2_REG1_REG_5__SCAN_IN), .A3(n7632), .ZN(
        n7634) );
  NAND2_X1 U5126 ( .A1(n5438), .A2(n5437), .ZN(n10248) );
  NAND2_X2 U5127 ( .A1(n6333), .A2(n6332), .ZN(n8246) );
  OR2_X1 U5128 ( .A1(n6298), .A2(n6433), .ZN(n6301) );
  NAND2_X1 U5129 ( .A1(n5360), .A2(n5156), .ZN(n7960) );
  NAND2_X1 U5130 ( .A1(n4544), .A2(n7535), .ZN(n7632) );
  INV_X4 U5131 ( .A(n7170), .ZN(n7240) );
  CLKBUF_X1 U5132 ( .A(n7286), .Z(n4419) );
  XNOR2_X1 U5133 ( .A(n5377), .B(n5376), .ZN(n7387) );
  NAND2_X1 U5134 ( .A1(n5470), .A2(n5466), .ZN(n5450) );
  INV_X1 U5135 ( .A(n8912), .ZN(n7899) );
  INV_X1 U5136 ( .A(n7887), .ZN(n7976) );
  NAND4_X1 U5137 ( .A1(n5463), .A2(n5462), .A3(n5461), .A4(n5460), .ZN(n8742)
         );
  AND4_X2 U5138 ( .A1(n5409), .A2(n5408), .A3(n5407), .A4(n5406), .ZN(n8256)
         );
  AND3_X2 U5139 ( .A1(n5158), .A2(n5344), .A3(n4432), .ZN(n8020) );
  NAND4_X1 U5140 ( .A1(n5366), .A2(n5367), .A3(n5365), .A4(n5364), .ZN(n8911)
         );
  AND2_X1 U5141 ( .A1(n6272), .A2(n6271), .ZN(n7842) );
  INV_X1 U5142 ( .A(n7052), .ZN(n7044) );
  INV_X1 U5143 ( .A(n8333), .ZN(n6377) );
  NAND4_X1 U5144 ( .A1(n6297), .A2(n6296), .A3(n6295), .A4(n6294), .ZN(n9622)
         );
  AND4_X1 U5145 ( .A1(n4675), .A2(n5308), .A3(n5307), .A4(n5309), .ZN(n7766)
         );
  AND2_X1 U5146 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  NAND2_X1 U5147 ( .A1(n7046), .A2(n8445), .ZN(n7052) );
  NAND4_X1 U5148 ( .A1(n5188), .A2(n5187), .A3(n5300), .A4(n5186), .ZN(n5185)
         );
  AND4_X1 U5149 ( .A1(n6363), .A2(n6362), .A3(n6361), .A4(n6360), .ZN(n8438)
         );
  OR2_X1 U5150 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  NAND4_X2 U5151 ( .A1(n6343), .A2(n6342), .A3(n6341), .A4(n6340), .ZN(n8210)
         );
  AND4_X1 U5152 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n6320)
         );
  CLKBUF_X3 U5153 ( .A(n5404), .Z(n6092) );
  NAND2_X1 U5154 ( .A1(n5395), .A2(n5396), .ZN(n4556) );
  NAND3_X1 U5155 ( .A1(n6651), .A2(n6869), .A3(n6650), .ZN(n7049) );
  NAND4_X2 U5156 ( .A1(n6288), .A2(n6287), .A3(n6286), .A4(n6285), .ZN(n10161)
         );
  CLKBUF_X1 U5157 ( .A(n4711), .Z(n4624) );
  OR2_X1 U5158 ( .A1(n4711), .A2(n10256), .ZN(n5188) );
  NAND2_X2 U5159 ( .A1(n6148), .A2(n6144), .ZN(n6910) );
  NAND2_X1 U5160 ( .A1(n4621), .A2(n4620), .ZN(n7631) );
  NAND2_X2 U5161 ( .A1(n8611), .A2(n5270), .ZN(n5404) );
  CLKBUF_X3 U5162 ( .A(n6282), .Z(n6573) );
  AOI21_X1 U5163 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(n9671) );
  NAND2_X1 U5164 ( .A1(n5650), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5652) );
  NOR2_X1 U5165 ( .A1(n10585), .A2(n10140), .ZN(n10141) );
  XNOR2_X1 U5166 ( .A(n6204), .B(n4551), .ZN(n8127) );
  NOR2_X1 U5167 ( .A1(n5665), .A2(n5082), .ZN(n5081) );
  AND2_X1 U5168 ( .A1(n7393), .A2(n7370), .ZN(n6289) );
  NAND2_X1 U5169 ( .A1(n5269), .A2(n5270), .ZN(n5733) );
  CLKBUF_X2 U5170 ( .A(n6258), .Z(n7393) );
  NAND2_X1 U5171 ( .A1(n6501), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6204) );
  INV_X1 U5172 ( .A(n6848), .ZN(n8505) );
  NAND3_X1 U5173 ( .A1(n5323), .A2(n5322), .A3(n5321), .ZN(n5383) );
  XNOR2_X1 U5175 ( .A(n6209), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U5176 ( .A1(n5375), .A2(n10330), .ZN(n5392) );
  XNOR2_X1 U5177 ( .A(n6649), .B(n6648), .ZN(n8601) );
  OR2_X1 U5178 ( .A1(n6653), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U5179 ( .A1(n6653), .A2(n4597), .ZN(n6158) );
  OAI21_X1 U5180 ( .B1(n6208), .B2(n6207), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6209) );
  NAND2_X1 U5181 ( .A1(n5351), .A2(SI_4_), .ZN(n5387) );
  XNOR2_X1 U5182 ( .A(n5472), .B(SI_9_), .ZN(n5469) );
  NAND2_X1 U5183 ( .A1(n5281), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5279) );
  INV_X1 U5184 ( .A(n7382), .ZN(n7524) );
  XNOR2_X1 U5185 ( .A(n5359), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6983) );
  XNOR2_X1 U5186 ( .A(n5003), .B(n4906), .ZN(n8613) );
  NAND2_X2 U5187 ( .A1(n4696), .A2(n4410), .ZN(n10121) );
  AND2_X1 U5188 ( .A1(n5829), .A2(n5828), .ZN(n5837) );
  OR2_X1 U5189 ( .A1(n4427), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5398) );
  OAI211_X1 U5190 ( .C1(n5332), .C2(n5331), .A(n4427), .B(n4745), .ZN(n7382)
         );
  OR2_X1 U5191 ( .A1(n6454), .A2(n4900), .ZN(n4590) );
  NAND2_X1 U5192 ( .A1(n10108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5003) );
  OAI21_X1 U5193 ( .B1(n7378), .B2(P2_DATAO_REG_9__SCAN_IN), .A(n4772), .ZN(
        n5472) );
  NAND2_X1 U5194 ( .A1(n4965), .A2(n4966), .ZN(n5280) );
  OR2_X1 U5195 ( .A1(n5512), .A2(n5266), .ZN(n5860) );
  OAI22_X1 U5196 ( .A1(n6256), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n5347), .ZN(n5293) );
  AND2_X1 U5197 ( .A1(n6634), .A2(n6633), .ZN(n6640) );
  NAND2_X1 U5198 ( .A1(n5348), .A2(n4642), .ZN(n5350) );
  INV_X2 U5199 ( .A(n5347), .ZN(n7370) );
  AND2_X1 U5200 ( .A1(n6200), .A2(n6199), .ZN(n6633) );
  INV_X1 U5201 ( .A(n5347), .ZN(n6256) );
  NAND2_X1 U5202 ( .A1(n4876), .A2(n4875), .ZN(n5333) );
  NAND4_X1 U5203 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6367), .ZN(n6201)
         );
  AND3_X1 U5204 ( .A1(n6437), .A2(n6394), .A3(n6383), .ZN(n6153) );
  AND2_X1 U5205 ( .A1(n4573), .A2(n4572), .ZN(n6154) );
  NAND2_X1 U5206 ( .A1(n6269), .A2(n5025), .ZN(n6290) );
  AND3_X1 U5207 ( .A1(n5265), .A2(n5264), .A3(n5263), .ZN(n5479) );
  INV_X1 U5208 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4906) );
  INV_X2 U5209 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4546) );
  INV_X4 U5210 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5211 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5025) );
  INV_X1 U5212 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5595) );
  INV_X1 U5213 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5613) );
  INV_X1 U5214 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6639) );
  INV_X1 U5215 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5594) );
  NOR2_X1 U5216 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4549) );
  NOR2_X1 U5217 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4550) );
  NOR2_X1 U5218 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5255) );
  NOR2_X1 U5219 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5265) );
  NOR2_X1 U5220 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5264) );
  NOR2_X1 U5221 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5263) );
  INV_X1 U5222 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6199) );
  INV_X1 U5223 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6915) );
  NOR2_X1 U5224 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6152) );
  NOR2_X1 U5225 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4572) );
  NOR2_X1 U5226 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4573) );
  INV_X1 U5227 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6394) );
  INV_X1 U5228 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6437) );
  NOR2_X2 U5229 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6269) );
  INV_X1 U5230 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6202) );
  INV_X2 U5231 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5560) );
  INV_X1 U5232 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6383) );
  XNOR2_X1 U5233 ( .A(n5741), .B(n5740), .ZN(n8509) );
  NAND2_X1 U5234 ( .A1(n7755), .A2(n9242), .ZN(n5094) );
  NAND2_X2 U5235 ( .A1(n8393), .A2(n8392), .ZN(n8549) );
  NAND2_X2 U5236 ( .A1(n5884), .A2(n8287), .ZN(n7751) );
  OAI21_X2 U5237 ( .B1(n9123), .B2(n5903), .A(n6027), .ZN(n9105) );
  NAND3_X1 U5238 ( .A1(n7048), .A2(n7369), .A3(n8136), .ZN(n7286) );
  OAI21_X2 U5239 ( .B1(n8003), .B2(n6720), .A(n6719), .ZN(n8174) );
  XNOR2_X1 U5240 ( .A(n6630), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7046) );
  AND2_X1 U5241 ( .A1(n8661), .A2(n6175), .ZN(n6281) );
  NOR2_X2 U5242 ( .A1(n9443), .A2(n9442), .ZN(n9505) );
  XNOR2_X2 U5243 ( .A(n9440), .B(n9506), .ZN(n9443) );
  OAI22_X2 U5244 ( .A1(n8625), .A2(n6826), .B1(n9827), .B2(n9538), .ZN(n9823)
         );
  OAI21_X2 U5245 ( .B1(n5851), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5881) );
  OAI21_X2 U5246 ( .B1(n9105), .B2(n6036), .A(n6032), .ZN(n9095) );
  OAI21_X2 U5247 ( .B1(n10157), .B2(n6659), .A(n6663), .ZN(n8003) );
  NAND2_X2 U5248 ( .A1(n4654), .A2(n6356), .ZN(n8324) );
  OAI22_X2 U5249 ( .A1(n7930), .A2(n5024), .B1(n5023), .B2(n7931), .ZN(n8152)
         );
  INV_X1 U5250 ( .A(n4413), .ZN(n9781) );
  NOR2_X1 U5251 ( .A1(n7045), .A2(n4413), .ZN(n4592) );
  XNOR2_X2 U5252 ( .A(n5450), .B(n5449), .ZN(n7406) );
  OAI21_X1 U5253 ( .B1(n5959), .B2(n5955), .A(n5958), .ZN(n5979) );
  AOI21_X1 U5254 ( .B1(n5950), .B2(n5951), .A(n4674), .ZN(n5953) );
  INV_X1 U5255 ( .A(n5066), .ZN(n5065) );
  OAI21_X1 U5256 ( .B1(n5740), .B2(n5067), .A(n5757), .ZN(n5066) );
  NAND2_X1 U5257 ( .A1(n5866), .A2(n5865), .ZN(n5921) );
  OR2_X1 U5258 ( .A1(n7400), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U5259 ( .A1(n5868), .A2(n5867), .ZN(n7749) );
  NOR2_X1 U5260 ( .A1(n5812), .A2(n4829), .ZN(n4828) );
  INV_X1 U5261 ( .A(n5790), .ZN(n4829) );
  NOR2_X1 U5262 ( .A1(n5756), .A2(n4822), .ZN(n4821) );
  INV_X1 U5263 ( .A(n5739), .ZN(n4822) );
  INV_X1 U5264 ( .A(n9133), .ZN(n5663) );
  OR2_X1 U5265 ( .A1(n9388), .A2(n8807), .ZN(n6010) );
  AND2_X1 U5266 ( .A1(n5145), .A2(n4485), .ZN(n5143) );
  NAND2_X1 U5267 ( .A1(n6815), .A2(n6816), .ZN(n5136) );
  NAND2_X1 U5268 ( .A1(n5777), .A2(n5776), .ZN(n5793) );
  INV_X1 U5269 ( .A(n5493), .ZN(n5072) );
  OAI21_X1 U5270 ( .B1(n7370), .B2(n4738), .A(n4737), .ZN(n5474) );
  NAND2_X1 U5271 ( .A1(n7370), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U5272 ( .A1(n9160), .A2(n6127), .ZN(n4826) );
  INV_X1 U5273 ( .A(n5214), .ZN(n5213) );
  NAND2_X1 U5275 ( .A1(n5902), .A2(n5208), .ZN(n5210) );
  NOR2_X1 U5276 ( .A1(n6110), .A2(n5209), .ZN(n5208) );
  INV_X1 U5277 ( .A(n6024), .ZN(n5209) );
  NAND2_X1 U5278 ( .A1(n4412), .A2(n7370), .ZN(n5358) );
  NAND2_X1 U5279 ( .A1(n4585), .A2(n7269), .ZN(n4582) );
  NAND2_X1 U5280 ( .A1(n7047), .A2(n8505), .ZN(n7048) );
  INV_X1 U5281 ( .A(n6751), .ZN(n6779) );
  OR2_X1 U5282 ( .A1(n10070), .A2(n9789), .ZN(n6753) );
  AND2_X1 U5283 ( .A1(n10070), .A2(n9789), .ZN(n6751) );
  AND2_X1 U5284 ( .A1(n5134), .A2(n4801), .ZN(n4548) );
  INV_X1 U5285 ( .A(n9074), .ZN(n8829) );
  AND2_X1 U5286 ( .A1(n5963), .A2(n4671), .ZN(n4955) );
  OR2_X1 U5287 ( .A1(n4887), .A2(n6485), .ZN(n4436) );
  AOI21_X1 U5288 ( .B1(n6483), .B2(n6669), .A(n4888), .ZN(n4887) );
  NAND2_X1 U5289 ( .A1(n4893), .A2(n6731), .ZN(n4892) );
  AOI21_X1 U5290 ( .B1(n5083), .B2(n5081), .A(n5080), .ZN(n5079) );
  INV_X1 U5291 ( .A(n5664), .ZN(n5080) );
  INV_X1 U5292 ( .A(n8877), .ZN(n5107) );
  NOR2_X1 U5293 ( .A1(n4441), .A2(n8848), .ZN(n5103) );
  INV_X1 U5294 ( .A(n9111), .ZN(n8709) );
  NAND2_X1 U5295 ( .A1(n6075), .A2(n6099), .ZN(n6141) );
  INV_X1 U5296 ( .A(n5270), .ZN(n5272) );
  NAND2_X1 U5297 ( .A1(n4534), .A2(n6918), .ZN(n6919) );
  NAND2_X1 U5298 ( .A1(n4697), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4533) );
  NOR2_X1 U5299 ( .A1(n6998), .A2(n10264), .ZN(n6925) );
  NOR2_X1 U5300 ( .A1(n8961), .A2(n4521), .ZN(n6975) );
  INV_X1 U5301 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n4764) );
  NOR2_X1 U5302 ( .A1(n10248), .A2(n8556), .ZN(n6121) );
  OAI21_X1 U5303 ( .B1(n7819), .B2(n4725), .A(n7904), .ZN(n4724) );
  INV_X1 U5304 ( .A(n5965), .ZN(n4725) );
  NAND2_X1 U5305 ( .A1(n7807), .A2(n7899), .ZN(n7825) );
  NAND2_X1 U5306 ( .A1(n9050), .A2(n9241), .ZN(n5849) );
  AND2_X1 U5307 ( .A1(n5250), .A2(n5773), .ZN(n5182) );
  OR2_X1 U5308 ( .A1(n5943), .A2(n9079), .ZN(n5906) );
  INV_X1 U5309 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5262) );
  INV_X1 U5310 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5254) );
  AOI22_X1 U5311 ( .A1(n9511), .A2(n9510), .B1(n9507), .B2(n9597), .ZN(n7194)
         );
  INV_X1 U5312 ( .A(n9510), .ZN(n4557) );
  INV_X1 U5313 ( .A(n8661), .ZN(n6174) );
  OR2_X2 U5314 ( .A1(n8652), .A2(n9806), .ZN(n7347) );
  NAND2_X1 U5315 ( .A1(n8652), .A2(n9806), .ZN(n6755) );
  OR2_X1 U5316 ( .A1(n9816), .A2(n9587), .ZN(n6776) );
  AND2_X1 U5317 ( .A1(n4849), .A2(n5237), .ZN(n4848) );
  AND2_X1 U5318 ( .A1(n6841), .A2(n6840), .ZN(n5237) );
  OR2_X1 U5319 ( .A1(n10195), .A2(n10161), .ZN(n6761) );
  AND2_X1 U5320 ( .A1(n5814), .A2(n5781), .ZN(n5792) );
  AOI21_X1 U5321 ( .B1(n5065), .B2(n5067), .A(n5063), .ZN(n5062) );
  INV_X1 U5322 ( .A(n5759), .ZN(n5063) );
  OAI21_X1 U5323 ( .B1(n7370), .B2(n4627), .A(n4626), .ZN(n5505) );
  NAND2_X1 U5324 ( .A1(n7370), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n4626) );
  AND2_X1 U5325 ( .A1(n8253), .A2(n8251), .ZN(n5127) );
  NAND2_X1 U5326 ( .A1(n8868), .A2(n5093), .ZN(n5092) );
  NOR2_X1 U5327 ( .A1(n7893), .A2(n4619), .ZN(n5126) );
  INV_X1 U5328 ( .A(n7889), .ZN(n4619) );
  XNOR2_X1 U5329 ( .A(n7035), .B(n6980), .ZN(n7762) );
  AND3_X1 U5330 ( .A1(n5585), .A2(n5584), .A3(n5583), .ZN(n8807) );
  NAND2_X2 U5331 ( .A1(n8611), .A2(n5272), .ZN(n4711) );
  OR2_X1 U5332 ( .A1(n5404), .A2(n5271), .ZN(n5274) );
  NAND2_X1 U5333 ( .A1(n4698), .A2(n7524), .ZN(n4697) );
  INV_X1 U5334 ( .A(n6919), .ZN(n4698) );
  INV_X1 U5335 ( .A(n7631), .ZN(n4869) );
  OR2_X1 U5336 ( .A1(n4945), .A2(n4943), .ZN(n4942) );
  INV_X1 U5337 ( .A(n4948), .ZN(n4943) );
  INV_X1 U5338 ( .A(n4946), .ZN(n4945) );
  OAI21_X1 U5339 ( .B1(n8936), .B2(n4950), .A(n8950), .ZN(n4946) );
  XNOR2_X1 U5340 ( .A(n8991), .B(n6975), .ZN(n8987) );
  NAND2_X1 U5341 ( .A1(n4949), .A2(n4948), .ZN(n4944) );
  OR2_X1 U5342 ( .A1(n8987), .A2(n10425), .ZN(n4882) );
  OR2_X1 U5343 ( .A1(n9334), .A2(n8829), .ZN(n6048) );
  OR2_X1 U5344 ( .A1(n6052), .A2(n6053), .ZN(n9052) );
  NAND2_X1 U5345 ( .A1(n9050), .A2(n9203), .ZN(n4705) );
  OR2_X1 U5346 ( .A1(n5683), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U5347 ( .A1(n6906), .A2(n5924), .ZN(n5927) );
  AND2_X1 U5348 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  NAND2_X1 U5349 ( .A1(n9039), .A2(n9203), .ZN(n9041) );
  AOI21_X1 U5350 ( .B1(n4819), .B2(n4821), .A(n4469), .ZN(n4818) );
  INV_X1 U5351 ( .A(n5180), .ZN(n4819) );
  NOR2_X1 U5352 ( .A1(n4457), .A2(n4825), .ZN(n4824) );
  INV_X1 U5353 ( .A(n5623), .ZN(n4825) );
  AND2_X1 U5354 ( .A1(n6017), .A2(n5191), .ZN(n5190) );
  INV_X1 U5355 ( .A(n6006), .ZN(n5195) );
  NAND2_X1 U5356 ( .A1(n9394), .A2(n8897), .ZN(n6006) );
  NOR2_X1 U5357 ( .A1(n5527), .A2(n5171), .ZN(n5170) );
  INV_X1 U5358 ( .A(n9145), .ZN(n9241) );
  INV_X2 U5359 ( .A(n5358), .ZN(n6086) );
  BUF_X1 U5360 ( .A(n5827), .Z(n5512) );
  OAI21_X1 U5361 ( .B1(n5628), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U5362 ( .A1(n4586), .A2(n4482), .ZN(n4585) );
  AOI21_X1 U5363 ( .B1(n5008), .B2(n5007), .A(n5006), .ZN(n5005) );
  INV_X1 U5364 ( .A(n7247), .ZN(n5007) );
  NAND2_X1 U5365 ( .A1(n4449), .A2(n7239), .ZN(n4584) );
  INV_X1 U5366 ( .A(n7392), .ZN(n7296) );
  INV_X1 U5367 ( .A(n6281), .ZN(n6310) );
  BUF_X1 U5368 ( .A(n6263), .Z(n6611) );
  NAND2_X1 U5369 ( .A1(n5154), .A2(n6830), .ZN(n5152) );
  AOI21_X1 U5370 ( .B1(n5141), .B2(n5143), .A(n4467), .ZN(n5140) );
  INV_X1 U5371 ( .A(n5146), .ZN(n5141) );
  NAND2_X1 U5372 ( .A1(n4706), .A2(n9904), .ZN(n4843) );
  AOI21_X1 U5373 ( .B1(n4795), .B2(n5134), .A(n4794), .ZN(n4797) );
  OAI21_X1 U5374 ( .B1(n6818), .B2(n4426), .A(n6820), .ZN(n4794) );
  AND2_X1 U5375 ( .A1(n4442), .A2(n4796), .ZN(n4795) );
  AOI21_X1 U5376 ( .B1(n4785), .B2(n4788), .A(n4484), .ZN(n4784) );
  NAND2_X1 U5377 ( .A1(n8324), .A2(n8438), .ZN(n8432) );
  AND2_X1 U5378 ( .A1(n6870), .A2(n10106), .ZN(n8132) );
  OR2_X1 U5379 ( .A1(n10105), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6870) );
  AND2_X1 U5380 ( .A1(n7296), .A2(n7564), .ZN(n10160) );
  INV_X1 U5381 ( .A(n10002), .ZN(n4605) );
  OR2_X1 U5382 ( .A1(n6834), .A2(n7045), .ZN(n10190) );
  AND2_X1 U5383 ( .A1(n7650), .A2(n6874), .ZN(n10211) );
  NAND2_X1 U5384 ( .A1(n6871), .A2(n10107), .ZN(n8131) );
  OR2_X1 U5385 ( .A1(n10105), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6871) );
  NAND2_X1 U5386 ( .A1(n4578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U5387 ( .A1(n5069), .A2(n4454), .ZN(n5529) );
  INV_X1 U5388 ( .A(n5509), .ZN(n5068) );
  NAND2_X1 U5389 ( .A1(n5475), .A2(n5476), .ZN(n5494) );
  XNOR2_X1 U5390 ( .A(n7957), .B(n9240), .ZN(n7893) );
  AND2_X1 U5391 ( .A1(n5789), .A2(n5788), .ZN(n8798) );
  INV_X1 U5392 ( .A(n9050), .ZN(n8884) );
  INV_X1 U5393 ( .A(n8798), .ZN(n9062) );
  NAND2_X1 U5394 ( .A1(n5772), .A2(n5771), .ZN(n9074) );
  OR2_X1 U5395 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  INV_X1 U5396 ( .A(n9458), .ZN(n4562) );
  NAND2_X1 U5397 ( .A1(n9559), .A2(n9561), .ZN(n4563) );
  INV_X1 U5398 ( .A(n9434), .ZN(n4574) );
  NOR2_X1 U5399 ( .A1(n6778), .A2(n4773), .ZN(n6780) );
  NAND2_X1 U5400 ( .A1(n6754), .A2(n4774), .ZN(n4773) );
  OR2_X1 U5401 ( .A1(n9831), .A2(n6573), .ZN(n6579) );
  OR2_X1 U5402 ( .A1(n6320), .A2(n6614), .ZN(n6345) );
  INV_X1 U5403 ( .A(n6365), .ZN(n4899) );
  NAND2_X1 U5404 ( .A1(n6022), .A2(n4969), .ZN(n4968) );
  AND2_X1 U5405 ( .A1(n6016), .A2(n6023), .ZN(n4969) );
  NAND2_X1 U5406 ( .A1(n5206), .A2(n6910), .ZN(n4967) );
  OR3_X1 U5407 ( .A1(n7346), .A2(n6597), .A3(n6834), .ZN(n6598) );
  NAND2_X1 U5408 ( .A1(n4734), .A2(n4733), .ZN(n4732) );
  INV_X1 U5409 ( .A(n8057), .ZN(n4733) );
  INV_X1 U5410 ( .A(n8905), .ZN(n4722) );
  AND2_X1 U5411 ( .A1(n5891), .A2(n5965), .ZN(n5956) );
  AND2_X1 U5412 ( .A1(n6108), .A2(n9080), .ZN(n5905) );
  NOR2_X1 U5413 ( .A1(n4571), .A2(n9520), .ZN(n5019) );
  OR2_X1 U5414 ( .A1(n7352), .A2(n8112), .ZN(n6682) );
  NAND2_X1 U5415 ( .A1(n5941), .A2(n5940), .ZN(n6061) );
  NAND2_X1 U5416 ( .A1(n4631), .A2(n4630), .ZN(n5382) );
  INV_X1 U5417 ( .A(SI_3_), .ZN(n4630) );
  NAND2_X1 U5418 ( .A1(n5107), .A2(n8795), .ZN(n5106) );
  INV_X1 U5419 ( .A(n8676), .ZN(n5120) );
  NAND2_X1 U5420 ( .A1(n4755), .A2(n8905), .ZN(n6142) );
  NAND2_X1 U5421 ( .A1(n6137), .A2(n6076), .ZN(n6099) );
  NAND2_X1 U5422 ( .A1(n5050), .A2(n5049), .ZN(n6097) );
  AND2_X1 U5423 ( .A1(n8904), .A2(n6068), .ZN(n5049) );
  OR2_X1 U5424 ( .A1(n6941), .A2(n6984), .ZN(n6917) );
  NAND2_X1 U5425 ( .A1(n4543), .A2(n6991), .ZN(n4983) );
  INV_X1 U5426 ( .A(n7869), .ZN(n4977) );
  OR2_X1 U5427 ( .A1(n4931), .A2(n7876), .ZN(n4927) );
  INV_X1 U5428 ( .A(n8997), .ZN(n4988) );
  AND2_X1 U5429 ( .A1(n10582), .A2(n4770), .ZN(n4769) );
  INV_X1 U5430 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4770) );
  INV_X1 U5431 ( .A(n5619), .ZN(n5618) );
  INV_X1 U5432 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4760) );
  NOR2_X1 U5433 ( .A1(n5498), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5517) );
  INV_X1 U5434 ( .A(n7960), .ZN(n5155) );
  AND2_X1 U5435 ( .A1(n6904), .A2(n5870), .ZN(n5918) );
  NAND2_X1 U5436 ( .A1(n8610), .A2(n6087), .ZN(n5050) );
  NAND2_X1 U5437 ( .A1(n5217), .A2(n6048), .ZN(n5216) );
  NAND2_X1 U5438 ( .A1(n9339), .A2(n8823), .ZN(n6108) );
  OR2_X1 U5439 ( .A1(n9339), .A2(n8823), .ZN(n6109) );
  OR2_X1 U5440 ( .A1(n9350), .A2(n8709), .ZN(n6037) );
  OR2_X1 U5441 ( .A1(n9365), .A2(n9146), .ZN(n6016) );
  OR2_X1 U5442 ( .A1(n9382), .A2(n8815), .ZN(n6019) );
  INV_X1 U5443 ( .A(n5526), .ZN(n5169) );
  NAND2_X1 U5444 ( .A1(n7038), .A2(n8606), .ZN(n6146) );
  INV_X1 U5445 ( .A(SI_17_), .ZN(n10497) );
  INV_X1 U5446 ( .A(n7268), .ZN(n5006) );
  AOI21_X1 U5447 ( .B1(n9479), .B2(n7247), .A(n4481), .ZN(n5008) );
  NOR2_X1 U5448 ( .A1(n9454), .A2(n9560), .ZN(n5009) );
  INV_X1 U5449 ( .A(n7229), .ZN(n5015) );
  OAI21_X1 U5450 ( .B1(n9478), .B2(n9479), .A(n7247), .ZN(n9455) );
  AOI21_X1 U5451 ( .B1(n5019), .B2(n5017), .A(n4513), .ZN(n5016) );
  INV_X1 U5452 ( .A(n5021), .ZN(n5017) );
  INV_X1 U5453 ( .A(n5019), .ZN(n5018) );
  NOR2_X1 U5454 ( .A1(n4779), .A2(n6773), .ZN(n4778) );
  NAND2_X1 U5455 ( .A1(n4780), .A2(n4416), .ZN(n4779) );
  OR2_X1 U5456 ( .A1(n4417), .A2(n6313), .ZN(n6314) );
  INV_X1 U5457 ( .A(n5231), .ZN(n5230) );
  OAI21_X1 U5458 ( .B1(n9804), .B2(n5232), .A(n7347), .ZN(n5231) );
  AND2_X1 U5459 ( .A1(n5140), .A2(n4448), .ZN(n4547) );
  NOR2_X1 U5460 ( .A1(n6522), .A2(n6521), .ZN(n4720) );
  NOR2_X1 U5461 ( .A1(n6505), .A2(n9572), .ZN(n4721) );
  NOR2_X1 U5462 ( .A1(n5033), .A2(n10043), .ZN(n5031) );
  OR2_X1 U5463 ( .A1(n9961), .A2(n9524), .ZN(n6740) );
  NAND2_X1 U5464 ( .A1(n6854), .A2(n5034), .ZN(n5033) );
  NAND2_X1 U5465 ( .A1(n4718), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6470) );
  INV_X1 U5466 ( .A(n6468), .ZN(n4718) );
  AND2_X1 U5467 ( .A1(n4786), .A2(n8588), .ZN(n4785) );
  NAND2_X1 U5468 ( .A1(n4787), .A2(n6810), .ZN(n4786) );
  INV_X1 U5469 ( .A(n6810), .ZN(n4788) );
  AND2_X1 U5470 ( .A1(n8348), .A2(n5046), .ZN(n5045) );
  NOR2_X1 U5471 ( .A1(n8490), .A2(n8317), .ZN(n5046) );
  NAND2_X1 U5472 ( .A1(n10210), .A2(n8005), .ZN(n8175) );
  AND2_X1 U5473 ( .A1(n8429), .A2(n8431), .ZN(n8295) );
  NAND2_X1 U5474 ( .A1(n6640), .A2(n6639), .ZN(n6645) );
  AND2_X1 U5475 ( .A1(n5759), .A2(n5746), .ZN(n5757) );
  AOI21_X1 U5476 ( .B1(n5076), .B2(n5075), .A(n5074), .ZN(n5073) );
  INV_X1 U5477 ( .A(n5704), .ZN(n5074) );
  INV_X1 U5478 ( .A(n5081), .ZN(n5075) );
  OAI21_X1 U5479 ( .B1(n5680), .B2(n5698), .A(n5699), .ZN(n5668) );
  AND2_X1 U5480 ( .A1(n6202), .A2(n6203), .ZN(n4591) );
  INV_X1 U5481 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6203) );
  OAI21_X1 U5482 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U5483 ( .A1(n5640), .A2(n5081), .ZN(n4782) );
  AOI21_X1 U5484 ( .B1(n5607), .B2(n5059), .A(n4476), .ZN(n5058) );
  INV_X1 U5485 ( .A(n5592), .ZN(n5059) );
  INV_X1 U5486 ( .A(n5589), .ZN(n4568) );
  NAND2_X1 U5487 ( .A1(n5535), .A2(n5534), .ZN(n5550) );
  AND2_X1 U5488 ( .A1(n4488), .A2(n5415), .ZN(n4686) );
  OAI21_X1 U5489 ( .B1(n5053), .B2(n5052), .A(n5473), .ZN(n5051) );
  NOR2_X1 U5490 ( .A1(n5466), .A2(n5054), .ZN(n5053) );
  NAND2_X1 U5491 ( .A1(n5281), .A2(n4951), .ZN(n5848) );
  AOI21_X1 U5492 ( .B1(n5280), .B2(n4461), .A(n4952), .ZN(n4951) );
  NOR2_X1 U5493 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4952) );
  INV_X1 U5494 ( .A(n8714), .ZN(n5105) );
  INV_X1 U5495 ( .A(n5110), .ZN(n5109) );
  OAI21_X1 U5496 ( .B1(n8877), .B2(n5111), .A(n8875), .ZN(n5110) );
  NOR2_X1 U5497 ( .A1(n5106), .A2(n5102), .ZN(n5100) );
  NOR2_X1 U5498 ( .A1(n5106), .A2(n5098), .ZN(n5097) );
  NAND2_X1 U5499 ( .A1(n5101), .A2(n4441), .ZN(n5098) );
  XNOR2_X1 U5500 ( .A(n7809), .B(n9248), .ZN(n7888) );
  INV_X1 U5501 ( .A(n5091), .ZN(n5090) );
  OAI21_X1 U5502 ( .B1(n5092), .B2(n8696), .A(n8698), .ZN(n5091) );
  INV_X1 U5503 ( .A(n8684), .ZN(n8762) );
  NAND2_X1 U5504 ( .A1(n8694), .A2(n8803), .ZN(n8813) );
  NAND2_X1 U5505 ( .A1(n5090), .A2(n5092), .ZN(n5089) );
  NAND2_X1 U5506 ( .A1(n8813), .A2(n5090), .ZN(n4613) );
  INV_X1 U5507 ( .A(n9248), .ZN(n7807) );
  NAND2_X1 U5508 ( .A1(n8716), .A2(n8829), .ZN(n5111) );
  OR3_X1 U5509 ( .A1(n5864), .A2(n5869), .A3(n9430), .ZN(n7038) );
  AND4_X1 U5510 ( .A1(n5489), .A2(n5488), .A3(n5487), .A4(n5486), .ZN(n8781)
         );
  OR2_X1 U5511 ( .A1(n5404), .A2(n5306), .ZN(n5309) );
  OAI21_X1 U5512 ( .B1(n7379), .B2(n6940), .A(n4874), .ZN(n7589) );
  NAND2_X1 U5513 ( .A1(n7379), .A2(n6940), .ZN(n4874) );
  XNOR2_X1 U5514 ( .A(n7379), .B(n10258), .ZN(n7592) );
  INV_X1 U5515 ( .A(n4533), .ZN(n4532) );
  NAND2_X1 U5516 ( .A1(n4932), .A2(n7724), .ZN(n4931) );
  NAND2_X1 U5517 ( .A1(n7627), .A2(n6994), .ZN(n4932) );
  AND2_X1 U5518 ( .A1(n7868), .A2(n4539), .ZN(n7728) );
  NAND2_X1 U5519 ( .A1(n4540), .A2(n7730), .ZN(n7868) );
  INV_X1 U5520 ( .A(n6924), .ZN(n4540) );
  OR2_X1 U5521 ( .A1(n4929), .A2(n7876), .ZN(n4926) );
  INV_X1 U5522 ( .A(n4930), .ZN(n4929) );
  OAI21_X1 U5523 ( .B1(n4931), .B2(n6994), .A(n7877), .ZN(n4930) );
  INV_X1 U5524 ( .A(n4927), .ZN(n4923) );
  AND2_X1 U5525 ( .A1(n6928), .A2(n8271), .ZN(n4982) );
  NAND2_X1 U5526 ( .A1(n8937), .A2(n8936), .ZN(n8935) );
  AND2_X1 U5527 ( .A1(n4989), .A2(n8998), .ZN(n8985) );
  NAND2_X1 U5528 ( .A1(n6933), .A2(n7940), .ZN(n8998) );
  OR2_X1 U5529 ( .A1(n8987), .A2(n4525), .ZN(n4880) );
  NAND2_X1 U5530 ( .A1(n6976), .A2(n4879), .ZN(n4878) );
  INV_X1 U5531 ( .A(n8996), .ZN(n4879) );
  NAND2_X1 U5532 ( .A1(n5804), .A2(n4762), .ZN(n9024) );
  OR2_X1 U5533 ( .A1(n5712), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5731) );
  OR2_X1 U5534 ( .A1(n9376), .A2(n9144), .ZN(n6024) );
  OR2_X1 U5535 ( .A1(n6110), .A2(n5206), .ZN(n9148) );
  OR2_X1 U5536 ( .A1(n5601), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U5537 ( .A1(n5541), .A2(n5540), .ZN(n5565) );
  OR2_X1 U5538 ( .A1(n8554), .A2(n8397), .ZN(n5985) );
  AND2_X1 U5539 ( .A1(n4766), .A2(n5457), .ZN(n4765) );
  NOR2_X1 U5540 ( .A1(n5410), .A2(n4810), .ZN(n4807) );
  INV_X1 U5541 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4771) );
  NAND2_X1 U5542 ( .A1(n4811), .A2(n7910), .ZN(n4809) );
  NAND2_X1 U5543 ( .A1(n7766), .A2(n7753), .ZN(n7848) );
  INV_X1 U5544 ( .A(n5921), .ZN(n6904) );
  AOI21_X1 U5545 ( .B1(n4730), .B2(n5175), .A(n4518), .ZN(n5174) );
  NOR2_X1 U5546 ( .A1(n6885), .A2(n9142), .ZN(n5175) );
  NAND2_X1 U5547 ( .A1(n8905), .A2(n9203), .ZN(n5850) );
  NAND2_X1 U5548 ( .A1(n4831), .A2(n5177), .ZN(n5176) );
  NOR2_X1 U5549 ( .A1(n4730), .A2(n5178), .ZN(n5177) );
  NAND2_X1 U5550 ( .A1(n6885), .A2(n9247), .ZN(n5178) );
  INV_X1 U5551 ( .A(n4821), .ZN(n4820) );
  NAND2_X1 U5552 ( .A1(n6037), .A2(n6038), .ZN(n9097) );
  INV_X1 U5553 ( .A(n5884), .ZN(n6936) );
  AND2_X1 U5554 ( .A1(n6016), .A2(n6026), .ZN(n9133) );
  AOI21_X1 U5555 ( .B1(n4429), .B2(n5163), .A(n4466), .ZN(n5160) );
  OAI21_X1 U5556 ( .B1(n5195), .B2(n6005), .A(n6010), .ZN(n5194) );
  AND2_X1 U5557 ( .A1(n5985), .A2(n6118), .ZN(n5223) );
  OR2_X1 U5558 ( .A1(n8163), .A2(n8164), .ZN(n5224) );
  OR2_X1 U5559 ( .A1(n7751), .A2(n6910), .ZN(n7737) );
  NAND2_X1 U5560 ( .A1(n5868), .A2(n5863), .ZN(n7400) );
  NAND2_X1 U5561 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n4964) );
  INV_X1 U5562 ( .A(n4964), .ZN(n4959) );
  INV_X1 U5563 ( .A(n4966), .ZN(n5266) );
  INV_X1 U5564 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5853) );
  INV_X1 U5565 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5830) );
  INV_X1 U5566 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5648) );
  XNOR2_X1 U5567 ( .A(n5436), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6998) );
  INV_X1 U5568 ( .A(n6941), .ZN(n4876) );
  AND2_X1 U5569 ( .A1(n4558), .A2(n4452), .ZN(n9510) );
  NAND2_X1 U5570 ( .A1(n9961), .A2(n7230), .ZN(n4558) );
  AND2_X1 U5571 ( .A1(n7187), .A2(n7186), .ZN(n9597) );
  AND3_X1 U5572 ( .A1(n7295), .A2(n8132), .A3(n7294), .ZN(n7318) );
  AND2_X1 U5573 ( .A1(n6748), .A2(n6834), .ZN(n4901) );
  AND4_X1 U5574 ( .A1(n6431), .A2(n6430), .A3(n6429), .A4(n6428), .ZN(n9444)
         );
  AND4_X1 U5575 ( .A1(n6376), .A2(n6375), .A3(n6374), .A4(n6373), .ZN(n8333)
         );
  NAND4_X1 U5576 ( .A1(n6246), .A2(n6244), .A3(n6245), .A4(n6247), .ZN(n6259)
         );
  OR2_X1 U5577 ( .A1(n6282), .A2(n9625), .ZN(n6246) );
  OR2_X1 U5578 ( .A1(n6284), .A2(n9629), .ZN(n6244) );
  AND2_X1 U5579 ( .A1(n7390), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7367) );
  AOI21_X1 U5580 ( .B1(n9643), .B2(n7555), .A(n7554), .ZN(n7553) );
  CLKBUF_X1 U5581 ( .A(n6394), .Z(n6436) );
  NOR2_X1 U5582 ( .A1(n9742), .A2(n9741), .ZN(n9752) );
  NOR2_X1 U5583 ( .A1(n9752), .A2(n4676), .ZN(n9767) );
  OR2_X1 U5584 ( .A1(n9750), .A2(n9751), .ZN(n4676) );
  AND2_X1 U5585 ( .A1(n6188), .A2(n6187), .ZN(n9806) );
  OR2_X1 U5586 ( .A1(n8650), .A2(n6573), .ZN(n6188) );
  NOR2_X1 U5587 ( .A1(n9829), .A2(n9998), .ZN(n9813) );
  INV_X1 U5588 ( .A(n4552), .ZN(n8617) );
  NAND2_X1 U5589 ( .A1(n8617), .A2(n8616), .ZN(n8615) );
  NAND2_X1 U5590 ( .A1(n4844), .A2(n4848), .ZN(n9824) );
  NAND2_X1 U5591 ( .A1(n4679), .A2(n6839), .ZN(n4844) );
  INV_X1 U5592 ( .A(n8633), .ZN(n4659) );
  INV_X1 U5593 ( .A(n5143), .ZN(n5142) );
  AND2_X1 U5594 ( .A1(n6756), .A2(n8632), .ZN(n9843) );
  OR2_X1 U5595 ( .A1(n9876), .A2(n9862), .ZN(n5145) );
  NOR2_X1 U5596 ( .A1(n6824), .A2(n5147), .ZN(n5146) );
  INV_X1 U5597 ( .A(n6822), .ZN(n5147) );
  AND2_X1 U5598 ( .A1(n6539), .A2(n6837), .ZN(n9860) );
  AND2_X1 U5599 ( .A1(n4442), .A2(n4801), .ZN(n4793) );
  NAND2_X1 U5600 ( .A1(n9937), .A2(n5236), .ZN(n9912) );
  AND2_X1 U5601 ( .A1(n6743), .A2(n6741), .ZN(n5236) );
  INV_X1 U5602 ( .A(n9915), .ZN(n6743) );
  NAND2_X1 U5603 ( .A1(n5135), .A2(n4471), .ZN(n5134) );
  OR2_X1 U5604 ( .A1(n4492), .A2(n4430), .ZN(n5135) );
  NAND2_X1 U5605 ( .A1(n4717), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6493) );
  INV_X1 U5606 ( .A(n6470), .ZN(n4717) );
  AND2_X1 U5607 ( .A1(n6741), .A2(n6544), .ZN(n9938) );
  NAND2_X1 U5608 ( .A1(n9939), .A2(n9938), .ZN(n9937) );
  OR2_X1 U5609 ( .A1(n9958), .A2(n6815), .ZN(n9956) );
  NAND2_X1 U5610 ( .A1(n6740), .A2(n6737), .ZN(n9948) );
  OAI21_X1 U5611 ( .B1(n4609), .B2(n4788), .A(n4785), .ZN(n8583) );
  BUF_X1 U5612 ( .A(n8585), .Z(n4739) );
  NAND2_X1 U5614 ( .A1(n4609), .A2(n8346), .ZN(n8345) );
  AND2_X1 U5615 ( .A1(n8358), .A2(n6726), .ZN(n5235) );
  NAND2_X1 U5616 ( .A1(n6165), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6387) );
  OAI21_X1 U5617 ( .B1(n5132), .B2(n5131), .A(n5130), .ZN(n8428) );
  AOI21_X1 U5618 ( .B1(n5129), .B2(n8330), .A(n4470), .ZN(n5130) );
  INV_X1 U5619 ( .A(n8330), .ZN(n5131) );
  INV_X1 U5620 ( .A(n10160), .ZN(n9921) );
  AND2_X1 U5621 ( .A1(n6280), .A2(n6279), .ZN(n10195) );
  NOR2_X1 U5622 ( .A1(n8130), .A2(n8132), .ZN(n7338) );
  NAND2_X1 U5623 ( .A1(n6869), .A2(n6858), .ZN(n10105) );
  INV_X1 U5624 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5002) );
  AND2_X1 U5625 ( .A1(n6172), .A2(n5002), .ZN(n5001) );
  NAND2_X1 U5626 ( .A1(n5027), .A2(n4741), .ZN(n4740) );
  INV_X1 U5627 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6643) );
  OR2_X1 U5628 ( .A1(n6409), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6422) );
  AOI21_X1 U5629 ( .B1(n5477), .B2(n5071), .A(n4483), .ZN(n5070) );
  NAND2_X1 U5630 ( .A1(n4685), .A2(n5051), .ZN(n5476) );
  NAND2_X1 U5631 ( .A1(n5095), .A2(n5101), .ZN(n5112) );
  AND4_X1 U5632 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n8556)
         );
  OR2_X1 U5633 ( .A1(n5544), .A2(n8402), .ZN(n5443) );
  NAND2_X1 U5634 ( .A1(n5630), .A2(n5629), .ZN(n9150) );
  AND2_X1 U5635 ( .A1(n8116), .A2(n8114), .ZN(n5128) );
  INV_X1 U5636 ( .A(n8889), .ZN(n8855) );
  NAND2_X1 U5637 ( .A1(n5783), .A2(n5782), .ZN(n9268) );
  NAND2_X1 U5638 ( .A1(n7700), .A2(n9207), .ZN(n8886) );
  OR2_X1 U5639 ( .A1(n7895), .A2(n7894), .ZN(n8899) );
  NAND2_X1 U5640 ( .A1(n5755), .A2(n5754), .ZN(n9089) );
  NAND2_X1 U5641 ( .A1(n5738), .A2(n5737), .ZN(n9099) );
  NAND2_X1 U5642 ( .A1(n5690), .A2(n5689), .ZN(n9136) );
  NAND2_X1 U5643 ( .A1(n5637), .A2(n5636), .ZN(n9161) );
  INV_X1 U5644 ( .A(n8807), .ZN(n9188) );
  INV_X1 U5645 ( .A(n8556), .ZN(n8908) );
  INV_X1 U5646 ( .A(n8256), .ZN(n8910) );
  NAND2_X1 U5647 ( .A1(n6088), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5315) );
  OR2_X1 U5648 ( .A1(n5404), .A2(n5311), .ZN(n5314) );
  NAND3_X2 U5649 ( .A1(n5275), .A2(n5276), .A3(n5277), .ZN(n8912) );
  AND2_X1 U5650 ( .A1(n5274), .A2(n5273), .ZN(n5275) );
  OAI21_X1 U5651 ( .B1(n7529), .B2(n4870), .A(n4868), .ZN(n7629) );
  AOI21_X1 U5652 ( .B1(n6953), .B2(n4872), .A(n4869), .ZN(n4868) );
  INV_X1 U5653 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4872) );
  NOR2_X1 U5654 ( .A1(n9003), .A2(n7035), .ZN(n8980) );
  NAND2_X1 U5655 ( .A1(n8987), .A2(n10425), .ZN(n4744) );
  NAND2_X1 U5656 ( .A1(n8990), .A2(n4689), .ZN(n4688) );
  AOI21_X1 U5657 ( .B1(n9011), .B2(n8991), .A(n4690), .ZN(n4689) );
  INV_X1 U5658 ( .A(n8989), .ZN(n4690) );
  NAND2_X1 U5659 ( .A1(n4939), .A2(n4938), .ZN(n8983) );
  AOI21_X1 U5660 ( .B1(n4439), .B2(n4944), .A(n4947), .ZN(n4938) );
  XNOR2_X1 U5661 ( .A(n6978), .B(n6981), .ZN(n4920) );
  AND3_X1 U5662 ( .A1(n4880), .A2(n4878), .A3(n6977), .ZN(n6978) );
  AND2_X1 U5663 ( .A1(n7414), .A2(n7033), .ZN(n9000) );
  INV_X1 U5664 ( .A(n7041), .ZN(n4919) );
  AND2_X1 U5665 ( .A1(n6899), .A2(n6898), .ZN(n4712) );
  NAND2_X1 U5666 ( .A1(n5218), .A2(n6048), .ZN(n9053) );
  NAND2_X1 U5667 ( .A1(n9067), .A2(n6049), .ZN(n5218) );
  AOI21_X1 U5668 ( .B1(n9051), .B2(n9247), .A(n4703), .ZN(n9271) );
  NAND2_X1 U5669 ( .A1(n4705), .A2(n4704), .ZN(n4703) );
  NAND2_X1 U5670 ( .A1(n9074), .A2(n9241), .ZN(n4704) );
  NOR2_X1 U5671 ( .A1(n9207), .A2(n4653), .ZN(n4652) );
  INV_X1 U5672 ( .A(n9077), .ZN(n4653) );
  NAND2_X1 U5673 ( .A1(n5483), .A2(n5482), .ZN(n8669) );
  INV_X1 U5674 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7896) );
  AND2_X1 U5675 ( .A1(n5928), .A2(n9191), .ZN(n9230) );
  AND2_X1 U5676 ( .A1(n8503), .A2(n8465), .ZN(n10249) );
  NAND2_X2 U5677 ( .A1(n5927), .A2(n9207), .ZN(n9253) );
  OR2_X1 U5678 ( .A1(n5800), .A2(n10410), .ZN(n5818) );
  AND3_X1 U5679 ( .A1(n5176), .A2(n5174), .A3(n5172), .ZN(n9258) );
  AOI21_X1 U5680 ( .B1(n9043), .B2(n9247), .A(n9042), .ZN(n9325) );
  NAND2_X1 U5681 ( .A1(n9062), .A2(n9241), .ZN(n9040) );
  OR2_X1 U5682 ( .A1(n7665), .A2(n5357), .ZN(n5564) );
  NAND2_X1 U5683 ( .A1(n5515), .A2(n5514), .ZN(n9406) );
  INV_X1 U5684 ( .A(n9372), .ZN(n9407) );
  OR2_X1 U5685 ( .A1(n10255), .A2(n10241), .ZN(n9372) );
  OR2_X1 U5686 ( .A1(n6556), .A2(n10429), .ZN(n6189) );
  OR2_X1 U5687 ( .A1(n7665), .A2(n6433), .ZN(n6445) );
  NOR2_X1 U5688 ( .A1(n7292), .A2(n7293), .ZN(n5026) );
  NAND2_X1 U5689 ( .A1(n4581), .A2(n4580), .ZN(n9497) );
  NAND2_X1 U5690 ( .A1(n4582), .A2(n4583), .ZN(n4581) );
  INV_X1 U5691 ( .A(n9498), .ZN(n4583) );
  NAND2_X1 U5692 ( .A1(n5004), .A2(n4561), .ZN(n4560) );
  INV_X1 U5693 ( .A(n9529), .ZN(n4561) );
  AND2_X1 U5694 ( .A1(n7327), .A2(n7326), .ZN(n9603) );
  OR2_X1 U5695 ( .A1(n7316), .A2(n10115), .ZN(n9584) );
  AND2_X1 U5696 ( .A1(n6584), .A2(n6583), .ZN(n9591) );
  INV_X1 U5697 ( .A(n9603), .ZN(n9590) );
  AOI211_X1 U5698 ( .C1(n6781), .C2(n6786), .A(n9781), .B(n6784), .ZN(n6782)
         );
  INV_X1 U5699 ( .A(n9806), .ZN(n9611) );
  INV_X1 U5700 ( .A(n9828), .ZN(n9613) );
  NAND2_X1 U5701 ( .A1(n6566), .A2(n6565), .ZN(n9844) );
  OR2_X1 U5702 ( .A1(n9531), .A2(n6573), .ZN(n6566) );
  NAND2_X1 U5703 ( .A1(n6538), .A2(n6537), .ZN(n9861) );
  NAND2_X1 U5704 ( .A1(n6528), .A2(n6527), .ZN(n9845) );
  INV_X1 U5705 ( .A(n9524), .ZN(n9978) );
  OR2_X1 U5706 ( .A1(n6282), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6287) );
  OR2_X1 U5707 ( .A1(n6282), .A2(n6262), .ZN(n6268) );
  OR2_X1 U5708 ( .A1(n6449), .A2(n6264), .ZN(n6266) );
  NAND2_X1 U5709 ( .A1(n6281), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6254) );
  OR2_X1 U5710 ( .A1(n6282), .A2(n7542), .ZN(n6253) );
  NAND2_X1 U5711 ( .A1(n9644), .A2(n9645), .ZN(n9643) );
  NOR2_X1 U5712 ( .A1(n9787), .A2(n9971), .ZN(n9986) );
  NAND2_X1 U5713 ( .A1(n4715), .A2(n4714), .ZN(n4713) );
  NAND2_X1 U5714 ( .A1(n9614), .A2(n10160), .ZN(n4714) );
  OR2_X1 U5715 ( .A1(n10167), .A2(n8207), .ZN(n9984) );
  OR2_X1 U5716 ( .A1(n10167), .A2(n8135), .ZN(n9976) );
  INV_X1 U5717 ( .A(n9801), .ZN(n10178) );
  NAND2_X1 U5718 ( .A1(n5150), .A2(n5149), .ZN(n5148) );
  NAND2_X1 U5719 ( .A1(n10004), .A2(n10211), .ZN(n4603) );
  INV_X1 U5720 ( .A(n10003), .ZN(n4604) );
  NAND2_X1 U5721 ( .A1(n4710), .A2(n10206), .ZN(n4709) );
  OR2_X1 U5722 ( .A1(n10010), .A2(n10215), .ZN(n4662) );
  NOR2_X1 U5723 ( .A1(n10006), .A2(n4600), .ZN(n10009) );
  OR2_X1 U5724 ( .A1(n10007), .A2(n4601), .ZN(n4600) );
  INV_X1 U5725 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5282) );
  INV_X1 U5726 ( .A(n5952), .ZN(n4674) );
  OAI211_X1 U5727 ( .C1(n6834), .C2(n6658), .A(n4904), .B(n4903), .ZN(n6323)
         );
  NAND2_X1 U5728 ( .A1(n4905), .A2(n6834), .ZN(n4904) );
  INV_X1 U5729 ( .A(n6350), .ZN(n4753) );
  NOR2_X1 U5730 ( .A1(n4673), .A2(n4672), .ZN(n4671) );
  NAND2_X1 U5731 ( .A1(n8053), .A2(n6100), .ZN(n4672) );
  INV_X1 U5732 ( .A(n5962), .ZN(n4673) );
  NAND2_X1 U5733 ( .A1(n5979), .A2(n5978), .ZN(n4954) );
  NAND2_X1 U5734 ( .A1(n5993), .A2(n6910), .ZN(n4636) );
  NOR2_X1 U5735 ( .A1(n4458), .A2(n4752), .ZN(n4751) );
  INV_X1 U5736 ( .A(n4833), .ZN(n4752) );
  NOR2_X1 U5737 ( .A1(n4458), .A2(n4896), .ZN(n4895) );
  INV_X1 U5738 ( .A(n6806), .ZN(n4896) );
  NAND2_X1 U5739 ( .A1(n6003), .A2(n6123), .ZN(n4915) );
  NAND2_X1 U5740 ( .A1(n6011), .A2(n6100), .ZN(n4910) );
  NAND2_X1 U5741 ( .A1(n4886), .A2(n6834), .ZN(n4885) );
  NOR2_X1 U5742 ( .A1(n6475), .A2(n6834), .ZN(n4890) );
  AOI21_X1 U5743 ( .B1(n4617), .B2(n6030), .A(n4474), .ZN(n6035) );
  INV_X1 U5744 ( .A(n4884), .ZN(n4883) );
  AND2_X1 U5745 ( .A1(n8328), .A2(n8432), .ZN(n6655) );
  AND2_X1 U5746 ( .A1(n4973), .A2(n6055), .ZN(n4972) );
  NAND2_X1 U5747 ( .A1(n7807), .A2(n8912), .ZN(n5891) );
  NOR2_X1 U5748 ( .A1(n9826), .A2(n8633), .ZN(n4780) );
  INV_X1 U5749 ( .A(n9843), .ZN(n4850) );
  NAND2_X1 U5750 ( .A1(n4995), .A2(n4598), .ZN(n4597) );
  AND2_X1 U5751 ( .A1(n4598), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4996) );
  INV_X1 U5752 ( .A(n5742), .ZN(n5067) );
  INV_X1 U5753 ( .A(n5705), .ZN(n5078) );
  INV_X1 U5754 ( .A(n5643), .ZN(n5082) );
  INV_X1 U5755 ( .A(n5468), .ZN(n5054) );
  OAI21_X1 U5756 ( .B1(n7370), .B2(n4743), .A(n4742), .ZN(n5467) );
  NAND2_X1 U5757 ( .A1(n7370), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5758 ( .A1(n5283), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5759 ( .A1(n4857), .A2(n5282), .ZN(n4862) );
  NAND2_X1 U5760 ( .A1(n10523), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U5761 ( .A1(n4859), .A2(n4858), .ZN(n4857) );
  NAND2_X1 U5762 ( .A1(n5287), .A2(n5286), .ZN(n5317) );
  NOR2_X1 U5763 ( .A1(n8688), .A2(n5115), .ZN(n5114) );
  INV_X1 U5764 ( .A(n8691), .ZN(n5115) );
  INV_X1 U5765 ( .A(n8802), .ZN(n5117) );
  INV_X1 U5766 ( .A(n8663), .ZN(n5086) );
  NAND2_X1 U5767 ( .A1(n4731), .A2(n4450), .ZN(n6122) );
  NOR2_X1 U5768 ( .A1(n4732), .A2(n8446), .ZN(n4731) );
  INV_X1 U5769 ( .A(n9082), .ZN(n4735) );
  NOR2_X1 U5770 ( .A1(n9088), .A2(n9110), .ZN(n4736) );
  INV_X1 U5771 ( .A(n6077), .ZN(n4970) );
  NAND2_X1 U5772 ( .A1(n6132), .A2(n6100), .ZN(n4701) );
  NAND2_X1 U5773 ( .A1(n6141), .A2(n6910), .ZN(n4702) );
  AND2_X1 U5774 ( .A1(n7868), .A2(n4975), .ZN(n4974) );
  INV_X1 U5775 ( .A(n6925), .ZN(n4975) );
  INV_X1 U5776 ( .A(n8093), .ZN(n4866) );
  NAND2_X1 U5777 ( .A1(n8571), .A2(n5247), .ZN(n4541) );
  NAND2_X1 U5778 ( .A1(n4542), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U5779 ( .A1(n4817), .A2(n4815), .ZN(n5183) );
  AND2_X1 U5780 ( .A1(n9060), .A2(n4816), .ZN(n4815) );
  NAND2_X1 U5781 ( .A1(n4818), .A2(n4820), .ZN(n4816) );
  NAND2_X1 U5782 ( .A1(n5749), .A2(n4757), .ZN(n4756) );
  INV_X1 U5783 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5749) );
  INV_X1 U5784 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n4757) );
  OAI22_X1 U5785 ( .A1(n8043), .A2(n5446), .B1(n10248), .B2(n8908), .ZN(n8165)
         );
  AND2_X1 U5786 ( .A1(n5423), .A2(n4767), .ZN(n4766) );
  INV_X1 U5787 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4767) );
  NOR2_X1 U5788 ( .A1(n5973), .A2(n7915), .ZN(n5893) );
  NAND2_X1 U5789 ( .A1(n7847), .A2(n7849), .ZN(n7824) );
  AND2_X1 U5790 ( .A1(n5215), .A2(n6044), .ZN(n5211) );
  AND2_X1 U5791 ( .A1(n9110), .A2(n5691), .ZN(n5692) );
  OR2_X1 U5792 ( .A1(n9124), .A2(n8776), .ZN(n6031) );
  OR2_X1 U5793 ( .A1(n9356), .A2(n9121), .ZN(n6032) );
  NAND2_X1 U5794 ( .A1(n9179), .A2(n5586), .ZN(n5162) );
  INV_X1 U5795 ( .A(n5586), .ZN(n5163) );
  NAND2_X1 U5796 ( .A1(n5193), .A2(n5195), .ZN(n5191) );
  OR2_X1 U5797 ( .A1(n9406), .A2(n8860), .ZN(n6112) );
  OR2_X1 U5798 ( .A1(n8670), .A2(n8789), .ZN(n9198) );
  OR2_X1 U5799 ( .A1(n7717), .A2(n6146), .ZN(n7708) );
  INV_X1 U5800 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U5801 ( .A1(n4668), .A2(n5419), .ZN(n5433) );
  INV_X1 U5802 ( .A(n5418), .ZN(n4668) );
  NAND2_X1 U5803 ( .A1(n4670), .A2(n4669), .ZN(n5418) );
  INV_X1 U5804 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4669) );
  INV_X1 U5805 ( .A(n5398), .ZN(n4670) );
  INV_X1 U5806 ( .A(SI_29_), .ZN(n10526) );
  AND2_X1 U5807 ( .A1(n4413), .A2(n8445), .ZN(n7047) );
  NOR2_X1 U5808 ( .A1(n7932), .A2(n7130), .ZN(n5024) );
  INV_X1 U5809 ( .A(n7932), .ZN(n5023) );
  OAI21_X1 U5810 ( .B1(n6602), .B2(n6603), .A(n4781), .ZN(n6605) );
  INV_X1 U5811 ( .A(n8613), .ZN(n6175) );
  NAND2_X1 U5812 ( .A1(n5038), .A2(n7303), .ZN(n5037) );
  NOR2_X1 U5813 ( .A1(n6582), .A2(n9583), .ZN(n4719) );
  NOR2_X1 U5814 ( .A1(n9816), .A2(n9998), .ZN(n5038) );
  OR2_X1 U5815 ( .A1(n10004), .A2(n9585), .ZN(n6775) );
  INV_X1 U5816 ( .A(n9842), .ZN(n4679) );
  NOR2_X1 U5817 ( .A1(n10028), .A2(n9876), .ZN(n5041) );
  INV_X1 U5818 ( .A(n6816), .ZN(n5137) );
  INV_X1 U5819 ( .A(n6811), .ZN(n5133) );
  OAI21_X1 U5820 ( .B1(n6758), .B2(n6657), .A(n6721), .ZN(n6722) );
  NAND2_X1 U5821 ( .A1(n8404), .A2(n6760), .ZN(n6658) );
  OR2_X1 U5822 ( .A1(n10105), .A2(n6868), .ZN(n7294) );
  XNOR2_X1 U5823 ( .A(n6260), .B(n6259), .ZN(n6791) );
  INV_X1 U5824 ( .A(n8231), .ZN(n6853) );
  NAND2_X1 U5825 ( .A1(n9887), .A2(n9894), .ZN(n9888) );
  INV_X1 U5826 ( .A(n7047), .ZN(n6874) );
  NAND2_X1 U5827 ( .A1(n5816), .A2(n5815), .ZN(n5937) );
  INV_X1 U5828 ( .A(n5639), .ZN(n5083) );
  AND2_X1 U5829 ( .A1(n5058), .A2(n5060), .ZN(n5056) );
  INV_X1 U5830 ( .A(n5624), .ZN(n5060) );
  NAND2_X1 U5831 ( .A1(n6208), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6627) );
  INV_X1 U5832 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U5833 ( .A1(n5575), .A2(n5574), .ZN(n5590) );
  NAND2_X1 U5834 ( .A1(n5529), .A2(n5528), .ZN(n5535) );
  OR2_X1 U5835 ( .A1(n6369), .A2(n6368), .ZN(n6382) );
  INV_X1 U5836 ( .A(n5414), .ZN(n5415) );
  NAND2_X1 U5837 ( .A1(n6256), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5369) );
  INV_X1 U5838 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4858) );
  AOI21_X1 U5839 ( .B1(n5122), .B2(n5120), .A(n5119), .ZN(n5118) );
  XNOR2_X1 U5840 ( .A(n9344), .B(n8684), .ZN(n8820) );
  NAND2_X1 U5841 ( .A1(n8739), .A2(n8676), .ZN(n5124) );
  OR2_X1 U5842 ( .A1(n8695), .A2(n9171), .ZN(n8696) );
  INV_X1 U5843 ( .A(n7966), .ZN(n7964) );
  INV_X1 U5844 ( .A(n6142), .ZN(n5202) );
  OR2_X1 U5845 ( .A1(n6140), .A2(n6141), .ZN(n5203) );
  NOR2_X1 U5846 ( .A1(n6143), .A2(n8465), .ZN(n5200) );
  NAND2_X1 U5847 ( .A1(n6131), .A2(n4729), .ZN(n4728) );
  NOR2_X1 U5848 ( .A1(n6132), .A2(n4730), .ZN(n4729) );
  INV_X1 U5849 ( .A(n6101), .ZN(n4611) );
  NOR2_X1 U5850 ( .A1(n5544), .A2(n4763), .ZN(n4761) );
  AND3_X1 U5851 ( .A1(n5605), .A2(n5604), .A3(n5603), .ZN(n8815) );
  OR2_X1 U5852 ( .A1(n4711), .A2(n10258), .ZN(n5273) );
  OAI21_X1 U5853 ( .B1(n7512), .B2(n6916), .A(n6917), .ZN(n7506) );
  NAND2_X1 U5854 ( .A1(n4937), .A2(n4936), .ZN(n4935) );
  NAND2_X1 U5855 ( .A1(n7033), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4936) );
  OR2_X1 U5856 ( .A1(n7033), .A2(n4666), .ZN(n4937) );
  NAND2_X1 U5857 ( .A1(n7592), .A2(n7591), .ZN(n4534) );
  NAND2_X1 U5858 ( .A1(n4533), .A2(n7469), .ZN(n6920) );
  NAND2_X1 U5859 ( .A1(n4983), .A2(n7632), .ZN(n7530) );
  NAND2_X1 U5860 ( .A1(n4538), .A2(n4536), .ZN(n7872) );
  NAND2_X1 U5861 ( .A1(n4537), .A2(n4977), .ZN(n4536) );
  NAND2_X1 U5862 ( .A1(n4512), .A2(n4926), .ZN(n7946) );
  OAI21_X1 U5863 ( .B1(n8919), .B2(n4541), .A(n8930), .ZN(n8920) );
  NAND2_X1 U5864 ( .A1(n4541), .A2(n8919), .ZN(n8930) );
  NAND2_X1 U5865 ( .A1(n6929), .A2(n4877), .ZN(n8971) );
  NAND2_X1 U5866 ( .A1(n4990), .A2(n8971), .ZN(n8973) );
  INV_X1 U5867 ( .A(n4991), .ZN(n4990) );
  INV_X1 U5868 ( .A(n8964), .ZN(n4940) );
  AND2_X1 U5869 ( .A1(n4988), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4987) );
  INV_X1 U5870 ( .A(n7033), .ZN(n6980) );
  OR2_X1 U5871 ( .A1(n4425), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5805) );
  OR2_X1 U5872 ( .A1(n5731), .A2(n4756), .ZN(n5766) );
  NAND2_X1 U5873 ( .A1(n5674), .A2(n5673), .ZN(n5712) );
  INV_X1 U5874 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5673) );
  INV_X1 U5875 ( .A(n5685), .ZN(n5674) );
  NOR2_X1 U5876 ( .A1(n5207), .A2(n5206), .ZN(n5205) );
  INV_X1 U5877 ( .A(n6026), .ZN(n5207) );
  INV_X1 U5878 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4768) );
  NAND2_X1 U5879 ( .A1(n5618), .A2(n4769), .ZN(n5656) );
  NAND2_X1 U5880 ( .A1(n5618), .A2(n10582), .ZN(n5631) );
  AND2_X1 U5881 ( .A1(n4438), .A2(n4759), .ZN(n4758) );
  INV_X1 U5882 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U5883 ( .A1(n5541), .A2(n4438), .ZN(n5581) );
  INV_X1 U5884 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5516) );
  OR2_X1 U5885 ( .A1(n5484), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U5886 ( .A1(n6118), .A2(n8531), .ZN(n8446) );
  NAND2_X1 U5887 ( .A1(n5424), .A2(n4766), .ZN(n5458) );
  NAND2_X1 U5888 ( .A1(n5424), .A2(n5423), .ZN(n5439) );
  NAND2_X1 U5889 ( .A1(n7896), .A2(n5340), .ZN(n5362) );
  INV_X1 U5890 ( .A(n4724), .ZN(n5892) );
  NAND2_X1 U5891 ( .A1(n5965), .A2(n7904), .ZN(n7827) );
  INV_X1 U5892 ( .A(n4813), .ZN(n4812) );
  OAI22_X1 U5893 ( .A1(n5800), .A2(n7380), .B1(n5357), .B2(n4814), .ZN(n4813)
         );
  NAND2_X1 U5894 ( .A1(n7749), .A2(n7748), .ZN(n6901) );
  NOR2_X1 U5895 ( .A1(n5918), .A2(n5917), .ZN(n6906) );
  NOR2_X1 U5896 ( .A1(n10243), .A2(n6144), .ZN(n6900) );
  NAND2_X1 U5897 ( .A1(n4629), .A2(n4628), .ZN(n6139) );
  NAND2_X1 U5898 ( .A1(n6086), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U5899 ( .A1(n9412), .A2(n6087), .ZN(n4629) );
  NAND2_X1 U5900 ( .A1(n5050), .A2(n6068), .ZN(n6137) );
  OR2_X1 U5901 ( .A1(n9344), .A2(n8851), .ZN(n9079) );
  AND2_X1 U5902 ( .A1(n5239), .A2(n5720), .ZN(n5180) );
  AOI21_X1 U5903 ( .B1(n5167), .B2(n5169), .A(n5165), .ZN(n5164) );
  INV_X1 U5904 ( .A(n6123), .ZN(n5165) );
  NAND2_X1 U5905 ( .A1(n8527), .A2(n8533), .ZN(n9221) );
  AOI21_X1 U5906 ( .B1(n5223), .B2(n8164), .A(n5221), .ZN(n5220) );
  INV_X1 U5907 ( .A(n5994), .ZN(n5221) );
  INV_X1 U5908 ( .A(n7708), .ZN(n7705) );
  AND2_X1 U5909 ( .A1(n5883), .A2(n7401), .ZN(n7703) );
  INV_X1 U5910 ( .A(n6146), .ZN(n7401) );
  AND2_X1 U5911 ( .A1(n7037), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7894) );
  NAND2_X1 U5912 ( .A1(n5832), .A2(n5831), .ZN(n5851) );
  INV_X1 U5913 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5831) );
  XNOR2_X1 U5914 ( .A(n5839), .B(P2_IR_REG_20__SCAN_IN), .ZN(n7746) );
  AND2_X1 U5915 ( .A1(n5577), .A2(n5562), .ZN(n8927) );
  NAND2_X1 U5916 ( .A1(n4873), .A2(n5333), .ZN(n7379) );
  NAND2_X1 U5917 ( .A1(n4875), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4992) );
  INV_X1 U5918 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5423) );
  INV_X1 U5919 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U5920 ( .A1(n7179), .A2(n7178), .ZN(n9440) );
  AND2_X1 U5921 ( .A1(n7289), .A2(n7288), .ZN(n7310) );
  AND2_X1 U5922 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n6163) );
  NOR2_X1 U5923 ( .A1(n7203), .A2(n5022), .ZN(n5021) );
  INV_X1 U5924 ( .A(n7178), .ZN(n5022) );
  NAND2_X1 U5925 ( .A1(n7201), .A2(n7200), .ZN(n4571) );
  AND2_X1 U5926 ( .A1(n7196), .A2(n4557), .ZN(n7197) );
  INV_X1 U5927 ( .A(n9486), .ZN(n4576) );
  AND2_X1 U5928 ( .A1(n7057), .A2(n7056), .ZN(n9560) );
  INV_X1 U5929 ( .A(n9455), .ZN(n9453) );
  INV_X1 U5930 ( .A(n6237), .ZN(n6169) );
  INV_X1 U5931 ( .A(n4720), .ZN(n6531) );
  NAND2_X1 U5932 ( .A1(n8479), .A2(n8480), .ZN(n8478) );
  OAI21_X1 U5933 ( .B1(n7179), .B2(n5018), .A(n5016), .ZN(n9466) );
  INV_X1 U5934 ( .A(n10104), .ZN(n7656) );
  NAND2_X1 U5935 ( .A1(n4781), .A2(n4776), .ZN(n4775) );
  NOR2_X1 U5936 ( .A1(n6845), .A2(n4777), .ZN(n4776) );
  NAND2_X1 U5937 ( .A1(n9804), .A2(n4778), .ZN(n4777) );
  AND4_X1 U5938 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(n7159)
         );
  NOR3_X1 U5939 ( .A1(n9683), .A2(n9682), .A3(n9681), .ZN(n9680) );
  AOI21_X1 U5940 ( .B1(n9713), .B2(P1_REG1_REG_15__SCAN_IN), .A(n4677), .ZN(
        n9715) );
  NOR2_X1 U5941 ( .A1(n7354), .A2(n7346), .ZN(n5228) );
  NOR2_X1 U5942 ( .A1(n5230), .A2(n4781), .ZN(n5227) );
  NAND2_X1 U5943 ( .A1(n7354), .A2(n7346), .ZN(n5229) );
  OR2_X1 U5944 ( .A1(n9818), .A2(n6573), .ZN(n6197) );
  NAND2_X1 U5945 ( .A1(n7347), .A2(n6755), .ZN(n6845) );
  NAND2_X1 U5946 ( .A1(n4719), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6192) );
  INV_X1 U5947 ( .A(n4719), .ZN(n6584) );
  NOR2_X1 U5948 ( .A1(n9829), .A2(n5036), .ZN(n9814) );
  INV_X1 U5949 ( .A(n5038), .ZN(n5036) );
  INV_X1 U5950 ( .A(n6842), .ZN(n4846) );
  NAND2_X1 U5951 ( .A1(n9612), .A2(n10158), .ZN(n4715) );
  NAND2_X1 U5952 ( .A1(n5140), .A2(n4465), .ZN(n5138) );
  NAND2_X1 U5953 ( .A1(n6823), .A2(n4547), .ZN(n5139) );
  NAND2_X1 U5954 ( .A1(n4720), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6560) );
  AND2_X1 U5955 ( .A1(n4428), .A2(n4606), .ZN(n8626) );
  AND2_X1 U5956 ( .A1(n9887), .A2(n5040), .ZN(n4606) );
  NAND2_X1 U5957 ( .A1(n9887), .A2(n4428), .ZN(n9853) );
  NAND2_X1 U5958 ( .A1(n4721), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6225) );
  INV_X1 U5959 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U5961 ( .A1(n9926), .A2(n5031), .ZN(n5030) );
  INV_X1 U5962 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9572) );
  INV_X1 U5963 ( .A(n4721), .ZN(n6507) );
  NAND2_X1 U5964 ( .A1(n6168), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6505) );
  NOR2_X1 U5965 ( .A1(n9972), .A2(n5029), .ZN(n9931) );
  INV_X1 U5966 ( .A(n5031), .ZN(n5029) );
  AND2_X1 U5967 ( .A1(n4835), .A2(n6739), .ZN(n4678) );
  NOR2_X1 U5968 ( .A1(n5044), .A2(n9555), .ZN(n5043) );
  INV_X1 U5969 ( .A(n5045), .ZN(n5044) );
  NAND2_X1 U5970 ( .A1(n6734), .A2(n4739), .ZN(n8520) );
  NAND2_X1 U5971 ( .A1(n8295), .A2(n8308), .ZN(n8364) );
  NAND2_X1 U5972 ( .A1(n8295), .A2(n5046), .ZN(n8362) );
  NAND2_X1 U5973 ( .A1(n8427), .A2(n6807), .ZN(n8290) );
  NAND2_X1 U5974 ( .A1(n4716), .A2(n4462), .ZN(n6400) );
  INV_X1 U5975 ( .A(n6387), .ZN(n4716) );
  NAND2_X1 U5976 ( .A1(n8428), .A2(n8437), .ZN(n8427) );
  AND2_X1 U5977 ( .A1(n8213), .A2(n4431), .ZN(n8429) );
  NAND2_X1 U5978 ( .A1(n8213), .A2(n4423), .ZN(n8325) );
  NAND2_X1 U5979 ( .A1(n6658), .A2(n6761), .ZN(n10157) );
  NAND2_X1 U5980 ( .A1(n8408), .A2(n8409), .ZN(n4553) );
  INV_X1 U5981 ( .A(n10195), .ZN(n8412) );
  OR2_X1 U5982 ( .A1(n8410), .A2(n8412), .ZN(n10172) );
  INV_X1 U5983 ( .A(n8445), .ZN(n7045) );
  AND2_X1 U5984 ( .A1(n6260), .A2(n6853), .ZN(n8147) );
  AND2_X1 U5985 ( .A1(n10158), .A2(n9790), .ZN(n9985) );
  AND2_X1 U5986 ( .A1(n8644), .A2(n7355), .ZN(n7356) );
  INV_X1 U5987 ( .A(n8639), .ZN(n5150) );
  NOR2_X1 U5988 ( .A1(n7354), .A2(n10215), .ZN(n5149) );
  INV_X1 U5989 ( .A(n10005), .ZN(n4710) );
  AND2_X1 U5990 ( .A1(n10008), .A2(n10211), .ZN(n4601) );
  AND2_X1 U5991 ( .A1(n7650), .A2(n8445), .ZN(n10174) );
  INV_X1 U5992 ( .A(n7311), .ZN(n7650) );
  AND2_X1 U5993 ( .A1(n7369), .A2(n7367), .ZN(n10104) );
  XNOR2_X1 U5994 ( .A(n6652), .B(P1_IR_REG_28__SCAN_IN), .ZN(n7564) );
  XNOR2_X1 U5995 ( .A(n5798), .B(n5797), .ZN(n9422) );
  XNOR2_X1 U5996 ( .A(n5793), .B(n5792), .ZN(n9426) );
  AND2_X1 U5997 ( .A1(n5742), .A2(n5728), .ZN(n5740) );
  XNOR2_X1 U5998 ( .A(n5670), .B(n5669), .ZN(n8424) );
  NAND2_X1 U5999 ( .A1(n4590), .A2(n4588), .ZN(n6631) );
  INV_X1 U6000 ( .A(n4589), .ZN(n4588) );
  OAI21_X1 U6001 ( .B1(n4591), .B2(n4900), .A(n6626), .ZN(n4589) );
  NAND2_X1 U6002 ( .A1(n6629), .A2(n6628), .ZN(n4578) );
  INV_X1 U6003 ( .A(n6631), .ZN(n6629) );
  NAND2_X1 U6004 ( .A1(n5057), .A2(n5058), .ZN(n5625) );
  XNOR2_X1 U6005 ( .A(n4569), .B(n5606), .ZN(n7804) );
  INV_X1 U6006 ( .A(n4567), .ZN(n4566) );
  OR2_X1 U6007 ( .A1(n6439), .A2(n6438), .ZN(n6441) );
  AND2_X1 U6008 ( .A1(n6422), .A2(n6410), .ZN(n7784) );
  NAND2_X1 U6009 ( .A1(n5494), .A2(n5493), .ZN(n5507) );
  NAND2_X1 U6010 ( .A1(n5416), .A2(n5415), .ZN(n5470) );
  AND2_X1 U6011 ( .A1(n6354), .A2(n6331), .ZN(n7613) );
  INV_X1 U6012 ( .A(n5383), .ZN(n5327) );
  NOR2_X1 U6013 ( .A1(n10138), .A2(n10137), .ZN(n10139) );
  AND2_X1 U6014 ( .A1(n8252), .A2(n8251), .ZN(n8254) );
  NOR2_X1 U6015 ( .A1(n4468), .A2(n5097), .ZN(n5096) );
  AND4_X1 U6016 ( .A1(n5548), .A2(n5547), .A3(n5546), .A4(n5545), .ZN(n8729)
         );
  NAND2_X1 U6017 ( .A1(n8892), .A2(n8691), .ZN(n8804) );
  OAI21_X1 U6018 ( .B1(n8549), .B2(n8550), .A(n8553), .ZN(n8664) );
  NAND2_X1 U6019 ( .A1(n4613), .A2(n4455), .ZN(n8701) );
  NAND2_X1 U6020 ( .A1(n5124), .A2(n5125), .ZN(n8841) );
  INV_X1 U6021 ( .A(n9099), .ZN(n8851) );
  INV_X1 U6022 ( .A(n5111), .ZN(n5108) );
  OR2_X1 U6023 ( .A1(n8891), .A2(n8890), .ZN(n8892) );
  XNOR2_X1 U6024 ( .A(n5833), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U6025 ( .A1(n5851), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6026 ( .A1(n5826), .A2(n5825), .ZN(n9039) );
  NAND2_X1 U6027 ( .A1(n5811), .A2(n5810), .ZN(n9050) );
  NAND2_X1 U6028 ( .A1(n5719), .A2(n5718), .ZN(n9111) );
  INV_X1 U6029 ( .A(n8815), .ZN(n9181) );
  OR2_X1 U6030 ( .A1(n7038), .A2(n7720), .ZN(n9003) );
  INV_X1 U6031 ( .A(n8781), .ZN(n8907) );
  CLKBUF_X1 U6032 ( .A(n6915), .Z(n7419) );
  INV_X1 U6033 ( .A(n9014), .ZN(n8988) );
  XNOR2_X1 U6034 ( .A(n4935), .B(n4934), .ZN(n7500) );
  INV_X1 U6035 ( .A(n4639), .ZN(n4934) );
  AOI21_X1 U6036 ( .B1(n7501), .B2(n7500), .A(n4933), .ZN(n7586) );
  AND2_X1 U6037 ( .A1(n4935), .A2(n4639), .ZN(n4933) );
  NAND2_X1 U6038 ( .A1(n4697), .A2(n7469), .ZN(n7518) );
  OR2_X1 U6039 ( .A1(n6992), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U6040 ( .A1(n6992), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U6041 ( .A1(n4871), .A2(n6953), .ZN(n7630) );
  NAND2_X1 U6042 ( .A1(n7529), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4871) );
  OAI21_X1 U6043 ( .B1(n4925), .B2(n4923), .A(n7944), .ZN(n4922) );
  NAND2_X1 U6044 ( .A1(n4864), .A2(n6961), .ZN(n8092) );
  NAND2_X1 U6045 ( .A1(n7943), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4864) );
  NAND2_X1 U6046 ( .A1(n4980), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U6047 ( .A1(n8935), .A2(n4949), .ZN(n8949) );
  NAND2_X1 U6048 ( .A1(n4941), .A2(n4942), .ZN(n8965) );
  OR2_X1 U6049 ( .A1(n8937), .A2(n4944), .ZN(n4941) );
  NAND2_X1 U6050 ( .A1(n4880), .A2(n4878), .ZN(n8995) );
  NAND2_X1 U6051 ( .A1(n4984), .A2(n4985), .ZN(n9002) );
  NAND2_X1 U6052 ( .A1(n4826), .A2(n5623), .ZN(n9141) );
  NAND2_X1 U6053 ( .A1(n5902), .A2(n6024), .ZN(n9149) );
  NAND2_X1 U6054 ( .A1(n4806), .A2(n4445), .ZN(n8084) );
  OR2_X1 U6055 ( .A1(n6913), .A2(n4639), .ZN(n5087) );
  AND2_X1 U6056 ( .A1(n5174), .A2(n10266), .ZN(n5173) );
  INV_X1 U6057 ( .A(n6139), .ZN(n9321) );
  NAND2_X1 U6058 ( .A1(n9271), .A2(n9270), .ZN(n9331) );
  NAND2_X1 U6059 ( .A1(n5765), .A2(n5764), .ZN(n9334) );
  OAI21_X1 U6060 ( .B1(n5181), .B2(n4820), .A(n4818), .ZN(n9061) );
  NAND2_X1 U6061 ( .A1(n8600), .A2(n6087), .ZN(n5748) );
  NAND2_X1 U6062 ( .A1(n5711), .A2(n5710), .ZN(n9350) );
  NAND2_X1 U6063 ( .A1(n5179), .A2(n5638), .ZN(n9132) );
  NAND2_X1 U6064 ( .A1(n5210), .A2(n6013), .ZN(n9130) );
  NAND2_X1 U6065 ( .A1(n5161), .A2(n5586), .ZN(n9169) );
  NAND2_X1 U6066 ( .A1(n9180), .A2(n9178), .ZN(n5161) );
  OAI21_X1 U6067 ( .B1(n4625), .B2(n5195), .A(n5193), .ZN(n9167) );
  NAND2_X1 U6068 ( .A1(n6006), .A2(n5192), .ZN(n9177) );
  NAND2_X1 U6069 ( .A1(n4625), .A2(n6005), .ZN(n5192) );
  NAND2_X1 U6070 ( .A1(n5166), .A2(n5526), .ZN(n9202) );
  NAND2_X1 U6071 ( .A1(n8527), .A2(n5170), .ZN(n5166) );
  NAND2_X1 U6072 ( .A1(n5224), .A2(n5223), .ZN(n8532) );
  INV_X1 U6073 ( .A(n8669), .ZN(n8745) );
  AOI22_X1 U6074 ( .A1(n6086), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6983), .B2(
        n5653), .ZN(n5156) );
  AND2_X1 U6075 ( .A1(n6911), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8606) );
  NAND2_X1 U6076 ( .A1(n7401), .A2(n7400), .ZN(n8609) );
  OR2_X1 U6077 ( .A1(n4966), .A2(n4964), .ZN(n4957) );
  NAND2_X1 U6078 ( .A1(n5280), .A2(n5862), .ZN(n9430) );
  INV_X1 U6079 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10543) );
  INV_X1 U6080 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U6081 ( .A1(n5856), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5858) );
  INV_X1 U6082 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8602) );
  INV_X1 U6083 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8512) );
  INV_X1 U6084 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8504) );
  INV_X1 U6085 ( .A(n6148), .ZN(n8503) );
  INV_X1 U6086 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8466) );
  INV_X1 U6087 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8286) );
  INV_X1 U6088 ( .A(n7746), .ZN(n8287) );
  INV_X1 U6089 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8126) );
  INV_X1 U6090 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5651) );
  INV_X1 U6091 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10441) );
  INV_X1 U6092 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7942) );
  INV_X1 U6093 ( .A(n7017), .ZN(n8919) );
  INV_X1 U6094 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7409) );
  INV_X1 U6095 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6096 ( .A1(n5331), .A2(n5267), .ZN(n4745) );
  CLKBUF_X1 U6097 ( .A(n7379), .Z(n4699) );
  CLKBUF_X1 U6098 ( .A(n7512), .Z(n4639) );
  INV_X1 U6099 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10582) );
  INV_X1 U6100 ( .A(n5011), .ZN(n5010) );
  NAND2_X1 U6101 ( .A1(n7153), .A2(n7155), .ZN(n8304) );
  NAND2_X1 U6102 ( .A1(n7687), .A2(n7086), .ZN(n7771) );
  NAND2_X1 U6103 ( .A1(n8478), .A2(n8482), .ZN(n9487) );
  INV_X1 U6104 ( .A(n4582), .ZN(n4579) );
  AND2_X1 U6105 ( .A1(n7107), .A2(n7106), .ZN(n8029) );
  NAND2_X1 U6106 ( .A1(n5020), .A2(n7202), .ZN(n9522) );
  INV_X1 U6107 ( .A(n4571), .ZN(n7202) );
  NAND2_X1 U6108 ( .A1(n7179), .A2(n5021), .ZN(n5020) );
  AND2_X1 U6109 ( .A1(n5013), .A2(n7228), .ZN(n5012) );
  INV_X1 U6110 ( .A(n9587), .ZN(n9612) );
  OR2_X1 U6111 ( .A1(n6474), .A2(n6473), .ZN(n9952) );
  INV_X1 U6112 ( .A(n8438), .ZN(n9620) );
  NAND2_X1 U6113 ( .A1(n6263), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n4783) );
  INV_X1 U6114 ( .A(n6320), .ZN(n10159) );
  OR2_X2 U6115 ( .A1(n7369), .A2(n7368), .ZN(n9623) );
  AND2_X1 U6116 ( .A1(n7432), .A2(n7431), .ZN(n7547) );
  INV_X1 U6117 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10132) );
  OAI21_X1 U6118 ( .B1(n7553), .B2(n9656), .A(n7428), .ZN(n9674) );
  NOR2_X1 U6119 ( .A1(n7600), .A2(n7601), .ZN(n9683) );
  AOI21_X1 U6120 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9690), .A(n9680), .ZN(
        n7669) );
  OR2_X1 U6121 ( .A1(n9704), .A2(n9703), .ZN(n9705) );
  AND2_X1 U6122 ( .A1(n9715), .A2(n9714), .ZN(n9740) );
  OR2_X1 U6123 ( .A1(n9735), .A2(n9736), .ZN(n9756) );
  NAND2_X1 U6124 ( .A1(n7547), .A2(n7567), .ZN(n9775) );
  NOR2_X1 U6125 ( .A1(n9767), .A2(n4530), .ZN(n9768) );
  AND2_X1 U6126 ( .A1(n7547), .A2(n10117), .ZN(n9779) );
  NAND2_X1 U6127 ( .A1(n8615), .A2(n5153), .ZN(n9810) );
  INV_X1 U6128 ( .A(n4681), .ZN(n4680) );
  OAI22_X1 U6129 ( .A1(n9828), .A2(n9919), .B1(n9921), .B2(n9827), .ZN(n4681)
         );
  AOI21_X1 U6130 ( .B1(n9614), .B2(n10158), .A(n4656), .ZN(n4655) );
  NAND2_X1 U6131 ( .A1(n4658), .A2(n10163), .ZN(n4657) );
  NOR2_X1 U6132 ( .A1(n9533), .A2(n9921), .ZN(n4656) );
  OAI21_X1 U6133 ( .B1(n6823), .B2(n5142), .A(n5140), .ZN(n9838) );
  NAND2_X1 U6134 ( .A1(n5144), .A2(n5145), .ZN(n9851) );
  NAND2_X1 U6135 ( .A1(n6823), .A2(n5146), .ZN(n5144) );
  NAND2_X1 U6136 ( .A1(n6823), .A2(n6822), .ZN(n9867) );
  NAND2_X1 U6137 ( .A1(n6835), .A2(n9884), .ZN(n9872) );
  AOI21_X1 U6138 ( .B1(n4793), .B2(n5134), .A(n4800), .ZN(n4798) );
  NAND2_X1 U6139 ( .A1(n9937), .A2(n6741), .ZN(n9914) );
  OR2_X1 U6140 ( .A1(n9958), .A2(n4442), .ZN(n4802) );
  NAND2_X1 U6141 ( .A1(n9956), .A2(n6816), .ZN(n9930) );
  NAND2_X1 U6142 ( .A1(n8583), .A2(n6811), .ZN(n8513) );
  NAND2_X1 U6143 ( .A1(n8345), .A2(n6810), .ZN(n8584) );
  NAND2_X1 U6144 ( .A1(n8341), .A2(n6730), .ZN(n8587) );
  AND2_X1 U6145 ( .A1(n8291), .A2(n6726), .ZN(n8359) );
  NAND2_X1 U6146 ( .A1(n8322), .A2(n8330), .ZN(n8323) );
  INV_X1 U6147 ( .A(n9984), .ZN(n10179) );
  MUX2_X1 U6148 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10125), .S(n7393), .Z(n8231)
         );
  INV_X1 U6149 ( .A(n9976), .ZN(n10168) );
  NAND2_X1 U6150 ( .A1(n7378), .A2(n4594), .ZN(n4593) );
  INV_X1 U6151 ( .A(n9961), .ZN(n6854) );
  AND2_X1 U6152 ( .A1(n6872), .A2(n8131), .ZN(n6873) );
  NOR2_X1 U6153 ( .A1(n4792), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U6154 ( .A1(n6173), .A2(n4995), .ZN(n4791) );
  NAND2_X1 U6155 ( .A1(n4999), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U6156 ( .A1(n6652), .A2(n5001), .ZN(n5000) );
  INV_X1 U6157 ( .A(n6172), .ZN(n4999) );
  INV_X1 U6158 ( .A(n7564), .ZN(n10115) );
  INV_X1 U6159 ( .A(n6869), .ZN(n10122) );
  INV_X1 U6160 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10359) );
  INV_X1 U6161 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8426) );
  INV_X1 U6162 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10396) );
  INV_X1 U6163 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8129) );
  INV_X1 U6164 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8041) );
  NAND2_X1 U6165 ( .A1(n4608), .A2(n4607), .ZN(n5557) );
  INV_X1 U6166 ( .A(n5555), .ZN(n4607) );
  INV_X1 U6167 ( .A(n5556), .ZN(n4608) );
  NAND2_X1 U6168 ( .A1(n5069), .A2(n5070), .ZN(n5510) );
  INV_X1 U6169 ( .A(n5476), .ZN(n4570) );
  AND2_X1 U6171 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10139), .ZN(n10586) );
  NOR2_X1 U6172 ( .A1(n10151), .A2(n10589), .ZN(n10299) );
  AOI21_X1 U6173 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10294), .ZN(n10292) );
  OAI21_X1 U6174 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10291), .ZN(n10289) );
  NAND2_X1 U6175 ( .A1(n10289), .A2(n10290), .ZN(n10288) );
  NAND2_X1 U6176 ( .A1(n10288), .A2(n4649), .ZN(n10286) );
  NAND2_X1 U6177 ( .A1(n10384), .A2(n4650), .ZN(n4649) );
  INV_X1 U6178 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n4650) );
  OAI21_X1 U6179 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10285), .ZN(n10283) );
  NAND2_X1 U6180 ( .A1(n10283), .A2(n10284), .ZN(n10282) );
  NAND2_X1 U6181 ( .A1(n10282), .A2(n4646), .ZN(n10280) );
  NAND2_X1 U6182 ( .A1(n4648), .A2(n4647), .ZN(n4646) );
  INV_X1 U6183 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n4648) );
  INV_X1 U6184 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n4647) );
  NAND2_X1 U6185 ( .A1(n7890), .A2(n7889), .ZN(n7892) );
  NAND2_X1 U6186 ( .A1(n5094), .A2(n7810), .ZN(n7760) );
  AND2_X1 U6187 ( .A1(n8115), .A2(n8114), .ZN(n8117) );
  AOI21_X1 U6188 ( .B1(n4434), .B2(n8578), .A(n4688), .ZN(n8992) );
  AND2_X1 U6189 ( .A1(n4507), .A2(n4919), .ZN(n4665) );
  INV_X1 U6190 ( .A(n5930), .ZN(n5931) );
  MUX2_X1 U6191 ( .A(n5925), .B(n9258), .S(n9253), .Z(n5932) );
  NAND2_X1 U6192 ( .A1(n9045), .A2(n9044), .ZN(n9048) );
  AND2_X1 U6193 ( .A1(n9338), .A2(n4519), .ZN(n9086) );
  OAI22_X1 U6194 ( .A1(n4755), .A2(n9298), .B1(n10266), .B2(n10483), .ZN(n6907) );
  OAI22_X1 U6195 ( .A1(n4755), .A2(n9372), .B1(n10254), .B2(n7332), .ZN(n7333)
         );
  INV_X1 U6196 ( .A(n5912), .ZN(n5913) );
  NAND2_X1 U6197 ( .A1(n9816), .A2(n9576), .ZN(n4691) );
  NAND2_X1 U6198 ( .A1(n4694), .A2(n4575), .ZN(P1_U3220) );
  NAND2_X1 U6199 ( .A1(n4574), .A2(n4451), .ZN(n4575) );
  NOR2_X1 U6200 ( .A1(n7309), .A2(n9578), .ZN(n4695) );
  NAND2_X1 U6201 ( .A1(n4559), .A2(n9598), .ZN(n9537) );
  NOR2_X1 U6202 ( .A1(n10000), .A2(n10167), .ZN(n8622) );
  AOI21_X1 U6203 ( .B1(n8652), .B2(n9992), .A(n7341), .ZN(n7342) );
  INV_X1 U6204 ( .A(n4853), .ZN(n4852) );
  OAI22_X1 U6205 ( .A1(n10078), .A2(n10066), .B1(n10225), .B2(n9996), .ZN(
        n4853) );
  NAND2_X1 U6206 ( .A1(n4661), .A2(n4660), .ZN(P1_U3546) );
  NAND2_X1 U6207 ( .A1(n10222), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n4660) );
  AOI21_X1 U6208 ( .B1(n7359), .B2(n10074), .A(n7364), .ZN(n7365) );
  INV_X1 U6209 ( .A(n6876), .ZN(n6877) );
  OAI22_X1 U6210 ( .A1(n7303), .A2(n10102), .B1(n10218), .B2(n6875), .ZN(n6876) );
  INV_X1 U6211 ( .A(n4804), .ZN(n4803) );
  OAI22_X1 U6212 ( .A1(n10078), .A2(n10102), .B1(n10218), .B2(n10077), .ZN(
        n4804) );
  NAND2_X1 U6213 ( .A1(n4708), .A2(n4522), .ZN(P1_U3515) );
  INV_X1 U6214 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n4707) );
  INV_X1 U6215 ( .A(n10156), .ZN(n4651) );
  AND2_X1 U6216 ( .A1(n8216), .A2(n8186), .ZN(n4423) );
  AND2_X1 U6217 ( .A1(n9486), .A2(n8480), .ZN(n4424) );
  INV_X1 U6218 ( .A(n8763), .ZN(n4730) );
  OR3_X1 U6219 ( .A1(n5731), .A2(n4756), .A3(P2_REG3_REG_25__SCAN_IN), .ZN(
        n4425) );
  NAND2_X1 U6220 ( .A1(n4837), .A2(n8520), .ZN(n9946) );
  OR2_X1 U6221 ( .A1(n5333), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n4427) );
  NAND2_X2 U6222 ( .A1(n6913), .A2(n7378), .ZN(n5357) );
  NAND2_X1 U6223 ( .A1(n4926), .A2(n7002), .ZN(n4925) );
  AND2_X1 U6224 ( .A1(n5041), .A2(n9857), .ZN(n4428) );
  AND2_X1 U6225 ( .A1(n9170), .A2(n5162), .ZN(n4429) );
  INV_X1 U6226 ( .A(n7352), .ZN(n7362) );
  INV_X1 U6227 ( .A(n7362), .ZN(n7359) );
  AND2_X1 U6228 ( .A1(n10043), .A2(n9953), .ZN(n4430) );
  NAND2_X1 U6229 ( .A1(n10028), .A2(n9907), .ZN(n9868) );
  INV_X1 U6230 ( .A(n9868), .ZN(n4841) );
  AND2_X1 U6231 ( .A1(n4423), .A2(n5028), .ZN(n4431) );
  OR2_X1 U6232 ( .A1(n4726), .A2(n6950), .ZN(n4432) );
  INV_X1 U6233 ( .A(n6757), .ZN(n4893) );
  NOR2_X1 U6234 ( .A1(n8482), .A2(n4576), .ZN(n4433) );
  NAND2_X1 U6235 ( .A1(n4882), .A2(n4744), .ZN(n4434) );
  OR2_X1 U6236 ( .A1(n8259), .A2(n8909), .ZN(n4435) );
  INV_X1 U6237 ( .A(n6659), .ZN(n4903) );
  AND2_X1 U6238 ( .A1(n5008), .A2(n4482), .ZN(n4437) );
  AND2_X1 U6239 ( .A1(n5540), .A2(n4760), .ZN(n4438) );
  AND2_X1 U6240 ( .A1(n4942), .A2(n4940), .ZN(n4439) );
  INV_X1 U6241 ( .A(n9614), .ZN(n9585) );
  OR2_X1 U6242 ( .A1(n8633), .A2(n6567), .ZN(n4440) );
  AND2_X1 U6243 ( .A1(n8710), .A2(n8709), .ZN(n4441) );
  NAND2_X1 U6244 ( .A1(n5136), .A2(n6817), .ZN(n4442) );
  INV_X1 U6245 ( .A(n5404), .ZN(n5714) );
  NAND2_X1 U6246 ( .A1(n4843), .A2(n6746), .ZN(n6835) );
  AND2_X1 U6247 ( .A1(n9898), .A2(n10092), .ZN(n9887) );
  INV_X1 U6248 ( .A(n7077), .ZN(n7058) );
  XNOR2_X1 U6249 ( .A(n5454), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7005) );
  OR2_X1 U6250 ( .A1(n5731), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4443) );
  NOR2_X1 U6251 ( .A1(n10058), .A2(n9979), .ZN(n4444) );
  OR2_X1 U6252 ( .A1(n8910), .A2(n8121), .ZN(n4445) );
  INV_X1 U6253 ( .A(n5168), .ZN(n5167) );
  OAI21_X1 U6254 ( .B1(n5170), .B2(n5169), .A(n6124), .ZN(n5168) );
  AND2_X1 U6255 ( .A1(n5590), .A2(n5589), .ZN(n4446) );
  INV_X1 U6256 ( .A(n4831), .ZN(n6882) );
  NAND2_X1 U6257 ( .A1(n5791), .A2(n4828), .ZN(n4831) );
  AND2_X1 U6258 ( .A1(n6000), .A2(n6001), .ZN(n4447) );
  XNOR2_X1 U6259 ( .A(n9327), .B(n8884), .ZN(n9037) );
  INV_X1 U6260 ( .A(n9037), .ZN(n4973) );
  NAND2_X1 U6261 ( .A1(n10011), .A2(n9861), .ZN(n4448) );
  INV_X1 U6262 ( .A(n8346), .ZN(n4787) );
  INV_X1 U6263 ( .A(n8652), .ZN(n7303) );
  INV_X1 U6264 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U6265 ( .A1(n5181), .A2(n5720), .ZN(n9087) );
  NAND2_X1 U6266 ( .A1(n4802), .A2(n5134), .ZN(n9911) );
  NAND2_X1 U6267 ( .A1(n6700), .A2(n6682), .ZN(n7354) );
  AND2_X1 U6268 ( .A1(n4437), .A2(n7238), .ZN(n4449) );
  AND4_X1 U6269 ( .A1(n6117), .A2(n8083), .A3(n6116), .A4(n7921), .ZN(n4450)
         );
  AND2_X1 U6270 ( .A1(n7309), .A2(n7308), .ZN(n4451) );
  INV_X1 U6271 ( .A(n6013), .ZN(n5206) );
  INV_X1 U6272 ( .A(n6201), .ZN(n4741) );
  AND2_X1 U6273 ( .A1(n6386), .A2(n6385), .ZN(n8308) );
  INV_X2 U6274 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5593) );
  OR2_X1 U6275 ( .A1(n9524), .A2(n4421), .ZN(n4452) );
  INV_X1 U6276 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6299) );
  AND2_X1 U6277 ( .A1(n5387), .A2(n5386), .ZN(n4453) );
  AND2_X1 U6278 ( .A1(n5070), .A2(n5068), .ZN(n4454) );
  NAND2_X1 U6279 ( .A1(n6425), .A2(n6424), .ZN(n9555) );
  AND2_X1 U6280 ( .A1(n5089), .A2(n8751), .ZN(n4455) );
  INV_X1 U6281 ( .A(n6107), .ZN(n6138) );
  AND2_X1 U6282 ( .A1(n8679), .A2(n9205), .ZN(n4456) );
  AND2_X1 U6283 ( .A1(n9150), .A2(n9161), .ZN(n4457) );
  INV_X1 U6284 ( .A(n6839), .ZN(n4851) );
  INV_X1 U6285 ( .A(n6731), .ZN(n4888) );
  NAND2_X1 U6286 ( .A1(n9887), .A2(n5041), .ZN(n5042) );
  AND2_X1 U6287 ( .A1(n6381), .A2(n4899), .ZN(n4458) );
  INV_X1 U6288 ( .A(n7346), .ZN(n5232) );
  AND2_X1 U6289 ( .A1(n5230), .A2(n4781), .ZN(n4459) );
  AND2_X1 U6290 ( .A1(n6023), .A2(n6024), .ZN(n4460) );
  AND2_X1 U6291 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4461) );
  AND2_X1 U6292 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_REG3_REG_9__SCAN_IN), 
        .ZN(n4462) );
  OR2_X1 U6293 ( .A1(n6004), .A2(n6003), .ZN(n4463) );
  AND2_X1 U6294 ( .A1(n6051), .A2(n6050), .ZN(n4464) );
  AND2_X1 U6295 ( .A1(n5142), .A2(n4448), .ZN(n4465) );
  INV_X1 U6296 ( .A(n6127), .ZN(n9159) );
  AND2_X1 U6297 ( .A1(n9382), .A2(n9181), .ZN(n4466) );
  AND2_X1 U6298 ( .A1(n10017), .A2(n9845), .ZN(n4467) );
  NAND2_X1 U6299 ( .A1(n5109), .A2(n5104), .ZN(n4468) );
  NOR2_X1 U6300 ( .A1(n9339), .A2(n9089), .ZN(n4469) );
  NOR2_X1 U6301 ( .A1(n8324), .A2(n9620), .ZN(n4470) );
  OR2_X1 U6302 ( .A1(n5136), .A2(n4430), .ZN(n4471) );
  AND2_X1 U6303 ( .A1(n4834), .A2(n5468), .ZN(n4472) );
  OR2_X1 U6304 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4473) );
  AND2_X1 U6305 ( .A1(n6029), .A2(n6910), .ZN(n4474) );
  AND2_X1 U6306 ( .A1(n9194), .A2(n4463), .ZN(n4475) );
  NAND2_X1 U6307 ( .A1(n5856), .A2(n5855), .ZN(n5869) );
  INV_X1 U6308 ( .A(n5102), .ZN(n5101) );
  OR2_X1 U6309 ( .A1(n8715), .A2(n5103), .ZN(n5102) );
  AND2_X1 U6310 ( .A1(n5608), .A2(SI_16_), .ZN(n4476) );
  AND2_X1 U6311 ( .A1(n4584), .A2(n4585), .ZN(n4477) );
  NAND2_X1 U6312 ( .A1(n6830), .A2(n8616), .ZN(n4478) );
  INV_X1 U6313 ( .A(n4838), .ZN(n4837) );
  NAND2_X1 U6314 ( .A1(n9977), .A2(n6735), .ZN(n4838) );
  NAND2_X1 U6315 ( .A1(n7331), .A2(n7330), .ZN(n4479) );
  INV_X1 U6316 ( .A(n5077), .ZN(n5076) );
  NAND2_X1 U6317 ( .A1(n5079), .A2(n5078), .ZN(n5077) );
  AND2_X1 U6318 ( .A1(n9809), .A2(n9808), .ZN(n4480) );
  INV_X1 U6319 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5451) );
  OR2_X1 U6320 ( .A1(n9457), .A2(n5009), .ZN(n4481) );
  INV_X1 U6321 ( .A(n6818), .ZN(n4800) );
  INV_X1 U6322 ( .A(n5035), .ZN(n7353) );
  NOR2_X1 U6323 ( .A1(n9829), .A2(n5037), .ZN(n5035) );
  AND2_X1 U6324 ( .A1(n7269), .A2(n7267), .ZN(n4482) );
  INV_X1 U6325 ( .A(n4482), .ZN(n5004) );
  NOR2_X1 U6326 ( .A1(n5505), .A2(SI_11_), .ZN(n4483) );
  OR2_X1 U6327 ( .A1(n4444), .A2(n5133), .ZN(n4484) );
  INV_X1 U6328 ( .A(n5154), .ZN(n5153) );
  NAND2_X1 U6329 ( .A1(n9811), .A2(n6829), .ZN(n5154) );
  OAI21_X1 U6330 ( .B1(n7370), .B2(n5370), .A(n5369), .ZN(n5385) );
  OR2_X1 U6331 ( .A1(n10017), .A2(n9845), .ZN(n4485) );
  AND2_X1 U6332 ( .A1(n5016), .A2(n5015), .ZN(n4486) );
  AND3_X1 U6333 ( .A1(n9119), .A2(n9133), .A3(n9094), .ZN(n4487) );
  AND2_X1 U6334 ( .A1(n5468), .A2(n5473), .ZN(n4488) );
  AND2_X1 U6335 ( .A1(n4730), .A2(n9247), .ZN(n4489) );
  AND2_X1 U6336 ( .A1(n6732), .A2(n6730), .ZN(n4490) );
  INV_X1 U6337 ( .A(n8348), .ZN(n9494) );
  AND2_X1 U6338 ( .A1(n6412), .A2(n6411), .ZN(n8348) );
  AND2_X1 U6339 ( .A1(n6727), .A2(n6729), .ZN(n4491) );
  AND2_X1 U6340 ( .A1(n6817), .A2(n5137), .ZN(n4492) );
  AND2_X1 U6341 ( .A1(n4967), .A2(n6026), .ZN(n4493) );
  AND2_X1 U6342 ( .A1(n7148), .A2(n7150), .ZN(n4494) );
  NAND2_X1 U6343 ( .A1(n6520), .A2(n6519), .ZN(n10017) );
  AND2_X1 U6344 ( .A1(n4977), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4495) );
  AND2_X1 U6345 ( .A1(n6019), .A2(n6010), .ZN(n4496) );
  AND2_X1 U6346 ( .A1(n4702), .A2(n4701), .ZN(n4497) );
  AND2_X1 U6347 ( .A1(n5268), .A2(n5267), .ZN(n4498) );
  AND2_X1 U6348 ( .A1(n5663), .A2(n5638), .ZN(n4499) );
  AND2_X1 U6349 ( .A1(n8520), .A2(n6735), .ZN(n4500) );
  AND2_X1 U6350 ( .A1(n4636), .A2(n4635), .ZN(n4501) );
  AND2_X1 U6351 ( .A1(n4445), .A2(n4435), .ZN(n4502) );
  OAI21_X1 U6352 ( .B1(n4977), .B2(n6925), .A(n7951), .ZN(n4976) );
  AND2_X1 U6353 ( .A1(n7272), .A2(n7273), .ZN(n4503) );
  AND2_X1 U6354 ( .A1(n4882), .A2(n4881), .ZN(n4504) );
  AND2_X1 U6355 ( .A1(n4579), .A2(n4584), .ZN(n4505) );
  NOR2_X1 U6356 ( .A1(n4473), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4963) );
  AND2_X1 U6357 ( .A1(n4447), .A2(n4915), .ZN(n4506) );
  INV_X1 U6358 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4598) );
  INV_X1 U6359 ( .A(n4925), .ZN(n4924) );
  NAND2_X1 U6360 ( .A1(n7042), .A2(n8980), .ZN(n4507) );
  INV_X1 U6361 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4995) );
  INV_X1 U6363 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5268) );
  INV_X1 U6364 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5325) );
  INV_X1 U6365 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5285) );
  INV_X1 U6366 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4832) );
  INV_X1 U6367 ( .A(n9207), .ZN(n9250) );
  AND2_X1 U6368 ( .A1(n5124), .A2(n5122), .ZN(n4508) );
  AND2_X1 U6369 ( .A1(n8213), .A2(n8216), .ZN(n4509) );
  AND2_X1 U6370 ( .A1(n7169), .A2(n7168), .ZN(n4510) );
  NOR2_X1 U6371 ( .A1(n7019), .A2(n8940), .ZN(n4950) );
  AND2_X1 U6372 ( .A1(n5224), .A2(n5985), .ZN(n4511) );
  INV_X1 U6373 ( .A(n6746), .ZN(n4842) );
  OR2_X1 U6374 ( .A1(n7628), .A2(n4927), .ZN(n4512) );
  INV_X1 U6375 ( .A(n10011), .ZN(n5040) );
  NOR2_X1 U6376 ( .A1(n9972), .A2(n5030), .ZN(n9898) );
  AND2_X1 U6377 ( .A1(n7212), .A2(n7211), .ZN(n4513) );
  INV_X1 U6378 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6434) );
  AND2_X1 U6379 ( .A1(n4979), .A2(n4980), .ZN(n4514) );
  INV_X1 U6380 ( .A(n4921), .ZN(n8105) );
  INV_X1 U6381 ( .A(n4928), .ZN(n7878) );
  AOI21_X1 U6382 ( .B1(n7628), .B2(n6994), .A(n4931), .ZN(n4928) );
  NAND2_X1 U6383 ( .A1(n8295), .A2(n5045), .ZN(n5047) );
  NOR2_X1 U6384 ( .A1(n9972), .A2(n10052), .ZN(n9959) );
  INV_X1 U6385 ( .A(n5032), .ZN(n9960) );
  NOR2_X1 U6386 ( .A1(n9972), .A2(n5033), .ZN(n5032) );
  AND2_X1 U6387 ( .A1(n5010), .A2(n7155), .ZN(n4515) );
  INV_X1 U6388 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U6389 ( .A1(n7144), .A2(n7143), .ZN(n8194) );
  NAND2_X1 U6390 ( .A1(n6454), .A2(n6202), .ZN(n4516) );
  NOR2_X1 U6391 ( .A1(n4978), .A2(n4982), .ZN(n4517) );
  NAND2_X1 U6392 ( .A1(n5850), .A2(n5849), .ZN(n4518) );
  INV_X1 U6393 ( .A(n4950), .ZN(n4949) );
  NOR2_X1 U6394 ( .A1(n9076), .A2(n4652), .ZN(n4519) );
  AND2_X1 U6395 ( .A1(n4769), .A2(n4768), .ZN(n4520) );
  INV_X1 U6396 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n4666) );
  INV_X1 U6397 ( .A(n8324), .ZN(n5028) );
  INV_X1 U6398 ( .A(n10225), .ZN(n10222) );
  INV_X1 U6399 ( .A(n7022), .ZN(n4877) );
  NAND2_X1 U6400 ( .A1(n7046), .A2(n4592), .ZN(n8136) );
  NAND2_X1 U6401 ( .A1(n10218), .A2(n10211), .ZN(n10102) );
  INV_X1 U6402 ( .A(n10052), .ZN(n5034) );
  NAND2_X1 U6403 ( .A1(n4578), .A2(n6632), .ZN(n8445) );
  AND2_X2 U6404 ( .A1(n7338), .A2(n6873), .ZN(n10218) );
  NAND2_X2 U6405 ( .A1(n5841), .A2(n5840), .ZN(n9247) );
  INV_X1 U6406 ( .A(n9247), .ZN(n9142) );
  AND2_X1 U6407 ( .A1(n8968), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4521) );
  INV_X1 U6408 ( .A(n8533), .ZN(n5171) );
  AND2_X1 U6409 ( .A1(n7318), .A2(n7297), .ZN(n9598) );
  INV_X1 U6410 ( .A(n10158), .ZN(n9919) );
  AND2_X1 U6411 ( .A1(n7296), .A2(n10115), .ZN(n10158) );
  INV_X1 U6412 ( .A(n8047), .ZN(n4734) );
  NAND2_X1 U6413 ( .A1(n6797), .A2(n6796), .ZN(n8408) );
  NAND2_X1 U6414 ( .A1(n7414), .A2(n6980), .ZN(n9020) );
  INV_X1 U6415 ( .A(n8723), .ZN(n5119) );
  INV_X1 U6416 ( .A(n10163), .ZN(n9917) );
  NAND2_X1 U6417 ( .A1(n6850), .A2(n6849), .ZN(n10163) );
  OR2_X1 U6418 ( .A1(n10218), .A2(n4707), .ZN(n4522) );
  NAND2_X1 U6419 ( .A1(n5132), .A2(n6805), .ZN(n8322) );
  AND2_X1 U6420 ( .A1(n7393), .A2(n4593), .ZN(n4523) );
  NAND2_X1 U6421 ( .A1(n4587), .A2(n7686), .ZN(n7687) );
  NOR2_X1 U6422 ( .A1(n5800), .A2(n9418), .ZN(n4524) );
  OR2_X1 U6423 ( .A1(n8996), .A2(n10425), .ZN(n4525) );
  OR2_X1 U6424 ( .A1(n8927), .A2(n10566), .ZN(n4526) );
  AND2_X1 U6425 ( .A1(n8940), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4527) );
  INV_X1 U6426 ( .A(n6114), .ZN(n4810) );
  AND2_X1 U6427 ( .A1(n4877), .A2(n6971), .ZN(n4528) );
  INV_X1 U6428 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n4743) );
  AND2_X1 U6429 ( .A1(n4532), .A2(n7469), .ZN(n4529) );
  XNOR2_X1 U6430 ( .A(n5296), .B(n5295), .ZN(n7374) );
  INV_X1 U6431 ( .A(n7374), .ZN(n4814) );
  INV_X1 U6432 ( .A(n8465), .ZN(n6144) );
  NAND2_X1 U6433 ( .A1(n5851), .A2(n5836), .ZN(n8465) );
  AND2_X1 U6434 ( .A1(n9769), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4530) );
  INV_X1 U6435 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n4981) );
  INV_X1 U6436 ( .A(n4763), .ZN(n4762) );
  NAND2_X1 U6437 ( .A1(n5803), .A2(n4764), .ZN(n4763) );
  AND2_X1 U6438 ( .A1(n7894), .A2(n7746), .ZN(n4531) );
  INV_X1 U6439 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n4594) );
  INV_X1 U6440 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4861) );
  INV_X1 U6441 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n4627) );
  INV_X1 U6442 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4643) );
  INV_X1 U6443 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n4738) );
  INV_X1 U6444 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4859) );
  OAI21_X1 U6445 ( .B1(n7592), .B2(n7591), .A(n4534), .ZN(n7593) );
  NAND3_X1 U6446 ( .A1(n9019), .A2(n4535), .A3(n9018), .ZN(P2_U3200) );
  OR2_X1 U6447 ( .A1(n9021), .A2(n9020), .ZN(n4535) );
  INV_X1 U6448 ( .A(n7868), .ZN(n4537) );
  NAND2_X1 U6449 ( .A1(n7728), .A2(n4495), .ZN(n4538) );
  NAND2_X1 U6450 ( .A1(n6924), .A2(n6955), .ZN(n4539) );
  NAND3_X1 U6451 ( .A1(n4748), .A2(n8568), .A3(n4747), .ZN(n8571) );
  AND2_X1 U6452 ( .A1(n8971), .A2(n4542), .ZN(n8948) );
  NAND2_X1 U6453 ( .A1(n6930), .A2(n7022), .ZN(n4542) );
  INV_X1 U6454 ( .A(n4544), .ZN(n4543) );
  NAND2_X1 U6455 ( .A1(n7468), .A2(n6921), .ZN(n4544) );
  OAI211_X1 U6456 ( .C1(n5301), .C2(n4546), .A(n6941), .B(n4545), .ZN(n7512)
         );
  NAND2_X1 U6457 ( .A1(n5267), .A2(n4546), .ZN(n4545) );
  NAND2_X2 U6458 ( .A1(n6915), .A2(n4546), .ZN(n6941) );
  OR2_X2 U6459 ( .A1(n9883), .A2(n6821), .ZN(n6823) );
  OAI21_X2 U6460 ( .B1(n4799), .B2(n4426), .A(n4797), .ZN(n9883) );
  NAND4_X2 U6461 ( .A1(n6206), .A2(n4550), .A3(n4549), .A4(n6202), .ZN(n4792)
         );
  AND2_X2 U6462 ( .A1(n6628), .A2(n4551), .ZN(n6206) );
  NAND2_X1 U6463 ( .A1(n6802), .A2(n8202), .ZN(n5132) );
  NAND2_X2 U6464 ( .A1(n6831), .A2(n6845), .ZN(n8639) );
  OAI21_X2 U6465 ( .B1(n4552), .B2(n4478), .A(n5152), .ZN(n6831) );
  OR2_X2 U6466 ( .A1(n6828), .A2(n5249), .ZN(n4552) );
  NAND2_X1 U6467 ( .A1(n4555), .A2(n4784), .ZN(n4554) );
  NAND2_X1 U6468 ( .A1(n8347), .A2(n4785), .ZN(n4555) );
  NAND2_X1 U6469 ( .A1(n8369), .A2(n6809), .ZN(n8347) );
  OAI211_X2 U6470 ( .C1(n5002), .C2(n6652), .A(n5000), .B(n4998), .ZN(n8661)
         );
  NAND2_X2 U6471 ( .A1(n6174), .A2(n8613), .ZN(n6284) );
  NAND2_X2 U6472 ( .A1(n4556), .A2(n5411), .ZN(n5416) );
  NAND2_X1 U6473 ( .A1(n5397), .A2(n4556), .ZN(n6298) );
  NAND3_X1 U6474 ( .A1(n4859), .A2(n5282), .A3(n4858), .ZN(n4565) );
  NAND3_X1 U6475 ( .A1(n10523), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4564) );
  OAI21_X1 U6476 ( .B1(n5575), .B2(n4568), .A(n4566), .ZN(n4569) );
  OAI21_X1 U6477 ( .B1(n4568), .B2(n5574), .A(n5592), .ZN(n4567) );
  NAND3_X1 U6478 ( .A1(n4685), .A2(n5051), .A3(n5071), .ZN(n5069) );
  NAND2_X1 U6479 ( .A1(n4570), .A2(n5477), .ZN(n5478) );
  AOI211_X2 U6480 ( .C1(n8479), .C2(n4424), .A(n4433), .B(n4510), .ZN(n4577)
         );
  INV_X1 U6481 ( .A(n4577), .ZN(n9549) );
  NAND3_X1 U6482 ( .A1(n7239), .A2(n4449), .A3(n4583), .ZN(n4580) );
  INV_X1 U6483 ( .A(n5005), .ZN(n4586) );
  NAND2_X1 U6484 ( .A1(n7653), .A2(n7684), .ZN(n4587) );
  OR2_X2 U6485 ( .A1(n7652), .A2(n7655), .ZN(n7653) );
  NAND2_X1 U6486 ( .A1(n6454), .A2(n4591), .ZN(n6208) );
  NAND2_X1 U6487 ( .A1(n8194), .A2(n7148), .ZN(n7152) );
  NAND2_X1 U6488 ( .A1(n8194), .A2(n4494), .ZN(n7153) );
  NAND2_X1 U6489 ( .A1(n5014), .A2(n5012), .ZN(n9542) );
  NOR2_X1 U6490 ( .A1(n9497), .A2(n4503), .ZN(n9582) );
  NAND2_X1 U6491 ( .A1(n9582), .A2(n9581), .ZN(n9580) );
  OR2_X1 U6492 ( .A1(n7083), .A2(n7084), .ZN(n7085) );
  NAND2_X1 U6493 ( .A1(n7771), .A2(n7772), .ZN(n7770) );
  NAND2_X2 U6494 ( .A1(n7044), .A2(n7369), .ZN(n7170) );
  NAND2_X1 U6495 ( .A1(n8292), .A2(n8293), .ZN(n8291) );
  NAND2_X1 U6496 ( .A1(n9859), .A2(n9860), .ZN(n9858) );
  NAND2_X1 U6497 ( .A1(n7839), .A2(n7840), .ZN(n7838) );
  NAND2_X1 U6498 ( .A1(n8620), .A2(n4416), .ZN(n8619) );
  INV_X1 U6499 ( .A(n4632), .ZN(n7361) );
  AND2_X1 U6500 ( .A1(n6779), .A2(n6621), .ZN(n5240) );
  NAND2_X1 U6501 ( .A1(n7063), .A2(n7064), .ZN(n4615) );
  NAND2_X2 U6502 ( .A1(n7068), .A2(n7067), .ZN(n7684) );
  NAND3_X1 U6503 ( .A1(n4727), .A2(n8465), .A3(n6130), .ZN(n5204) );
  NAND2_X1 U6504 ( .A1(n5126), .A2(n7890), .ZN(n7959) );
  NAND2_X1 U6505 ( .A1(n8725), .A2(n8687), .ZN(n8891) );
  NAND2_X1 U6506 ( .A1(n8704), .A2(n8703), .ZN(n8773) );
  NAND2_X1 U6507 ( .A1(n8290), .A2(n8289), .ZN(n8288) );
  OAI21_X2 U6508 ( .B1(n9969), .B2(n6814), .A(n6813), .ZN(n9958) );
  NAND3_X1 U6509 ( .A1(n8649), .A2(n4599), .A3(n8655), .ZN(n7339) );
  XNOR2_X1 U6511 ( .A(n8634), .B(n4659), .ZN(n4658) );
  NAND2_X1 U6512 ( .A1(n9912), .A2(n6744), .ZN(n9903) );
  AOI21_X2 U6513 ( .B1(n6852), .B2(n10163), .A(n6851), .ZN(n8649) );
  NAND2_X1 U6514 ( .A1(n9950), .A2(n6740), .ZN(n9939) );
  XNOR2_X1 U6515 ( .A(n6273), .B(n7842), .ZN(n7837) );
  NAND2_X1 U6516 ( .A1(n4602), .A2(n9869), .ZN(n9870) );
  NAND2_X1 U6517 ( .A1(n8140), .A2(n8139), .ZN(n8138) );
  OAI21_X1 U6518 ( .B1(n8174), .B2(n6723), .A(n6722), .ZN(n6724) );
  NAND2_X1 U6519 ( .A1(n4633), .A2(n4840), .ZN(n4602) );
  OAI21_X4 U6520 ( .B1(n4740), .B2(n4789), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6652) );
  NAND4_X1 U6521 ( .A1(n4709), .A2(n4605), .A3(n4604), .A4(n4603), .ZN(n10080)
         );
  AOI21_X2 U6522 ( .B1(n10074), .B2(n10073), .A(n10072), .ZN(n10075) );
  NOR2_X2 U6523 ( .A1(n9830), .A2(n10004), .ZN(n6855) );
  NAND2_X1 U6524 ( .A1(n4723), .A2(n4722), .ZN(n6075) );
  AOI21_X2 U6525 ( .B1(n4916), .B2(n6078), .A(n4640), .ZN(n6102) );
  NAND2_X2 U6526 ( .A1(n5904), .A2(n6037), .ZN(n9078) );
  NAND2_X1 U6527 ( .A1(n5842), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5186) );
  OAI21_X2 U6528 ( .B1(n8048), .B2(n6121), .A(n6119), .ZN(n8163) );
  NAND2_X1 U6529 ( .A1(n4623), .A2(n6019), .ZN(n9158) );
  OAI21_X1 U6530 ( .B1(n10076), .B2(n10217), .A(n4803), .ZN(P1_U3517) );
  OAI21_X1 U6531 ( .B1(n10076), .B2(n10222), .A(n4852), .ZN(P1_U3549) );
  OAI21_X1 U6532 ( .B1(n7361), .B2(n10222), .A(n7360), .ZN(P1_U3551) );
  AOI21_X2 U6533 ( .B1(n6104), .B2(n4610), .A(n6107), .ZN(n6105) );
  NAND2_X1 U6534 ( .A1(n4612), .A2(n4611), .ZN(n4610) );
  INV_X1 U6535 ( .A(n6102), .ZN(n4612) );
  NOR2_X1 U6536 ( .A1(n5114), .A2(n5117), .ZN(n5113) );
  AOI21_X1 U6537 ( .B1(n8550), .B2(n8553), .A(n5086), .ZN(n5085) );
  AOI21_X2 U6538 ( .B1(n4614), .B2(n6753), .A(n4901), .ZN(n6783) );
  NAND2_X1 U6539 ( .A1(n4902), .A2(n6624), .ZN(n4614) );
  XNOR2_X2 U6540 ( .A(n4615), .B(n7301), .ZN(n7068) );
  NOR2_X1 U6541 ( .A1(n4426), .A2(n6819), .ZN(n4796) );
  NAND2_X1 U6542 ( .A1(n4683), .A2(n10163), .ZN(n4682) );
  NAND2_X1 U6543 ( .A1(n9825), .A2(n9826), .ZN(n4684) );
  OAI21_X1 U6544 ( .B1(n4914), .B2(n4913), .A(n4475), .ZN(n6008) );
  NAND2_X1 U6545 ( .A1(n6792), .A2(n7230), .ZN(n7063) );
  NAND2_X1 U6546 ( .A1(n6056), .A2(n4972), .ZN(n4622) );
  NAND2_X1 U6547 ( .A1(n5992), .A2(n6100), .ZN(n4635) );
  NAND3_X1 U6548 ( .A1(n4912), .A2(n4911), .A3(n4493), .ZN(n4617) );
  AOI21_X1 U6549 ( .B1(n7870), .B2(n4974), .A(n4976), .ZN(n6927) );
  NOR2_X1 U6550 ( .A1(n8934), .A2(n4527), .ZN(n6930) );
  OR2_X1 U6551 ( .A1(n6699), .A2(n6698), .ZN(n6701) );
  NAND2_X1 U6552 ( .A1(n4993), .A2(n4992), .ZN(n4873) );
  INV_X1 U6553 ( .A(n4618), .ZN(n6711) );
  NOR3_X2 U6554 ( .A1(n6710), .A2(n7326), .A3(n6874), .ZN(n4618) );
  NAND2_X1 U6555 ( .A1(n7629), .A2(n6954), .ZN(n6956) );
  NAND2_X1 U6556 ( .A1(n4634), .A2(n4526), .ZN(n6972) );
  NAND2_X1 U6557 ( .A1(n6970), .A2(n6969), .ZN(n8929) );
  NAND2_X2 U6558 ( .A1(n6960), .A2(n7951), .ZN(n6961) );
  AOI21_X2 U6559 ( .B1(n8962), .B2(n8960), .A(n8959), .ZN(n8961) );
  NAND2_X1 U6560 ( .A1(n9903), .A2(n4839), .ZN(n4633) );
  NAND2_X1 U6561 ( .A1(n7838), .A2(n6274), .ZN(n8404) );
  NOR3_X1 U6562 ( .A1(n9698), .A2(n9697), .A3(n9696), .ZN(n9695) );
  XNOR2_X2 U6563 ( .A(n6248), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9628) );
  AOI211_X1 U6564 ( .C1(n6334), .C2(n7618), .A(n7430), .B(n7429), .ZN(n7626)
         );
  AND3_X2 U6565 ( .A1(n6894), .A2(n4622), .A3(n6059), .ZN(n4971) );
  NAND2_X1 U6566 ( .A1(n5189), .A2(n5190), .ZN(n4623) );
  NAND2_X1 U6567 ( .A1(n7845), .A2(n5950), .ZN(n9235) );
  NAND2_X1 U6568 ( .A1(n5901), .A2(n5900), .ZN(n9193) );
  OAI21_X2 U6569 ( .B1(n4909), .B2(n6127), .A(n6015), .ZN(n6022) );
  INV_X2 U6570 ( .A(n4711), .ZN(n5843) );
  OAI21_X1 U6571 ( .B1(n4955), .B2(n4953), .A(n4501), .ZN(n5996) );
  INV_X4 U6572 ( .A(n5733), .ZN(n6088) );
  NAND2_X1 U6573 ( .A1(n6088), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4675) );
  NAND2_X1 U6574 ( .A1(n4644), .A2(n4497), .ZN(n4640) );
  AOI21_X2 U6575 ( .B1(n9506), .B2(n9440), .A(n9505), .ZN(n9509) );
  AOI21_X1 U6576 ( .B1(n6018), .B2(n4496), .A(n4910), .ZN(n4909) );
  NOR2_X1 U6577 ( .A1(n7766), .A2(n7753), .ZN(n5951) );
  OAI21_X1 U6578 ( .B1(n6081), .B2(n6080), .A(n6079), .ZN(n6085) );
  NOR2_X1 U6579 ( .A1(n5506), .A2(n5072), .ZN(n5071) );
  OAI21_X1 U6580 ( .B1(n6622), .B2(n10073), .A(n5240), .ZN(n4902) );
  AOI21_X2 U6581 ( .B1(n8660), .B2(n6087), .A(n4524), .ZN(n4755) );
  NOR2_X1 U6582 ( .A1(n6077), .A2(n6884), .ZN(n4917) );
  NAND2_X1 U6583 ( .A1(n5837), .A2(n5830), .ZN(n5834) );
  NAND2_X1 U6584 ( .A1(n5854), .A2(n5853), .ZN(n5856) );
  NAND2_X1 U6585 ( .A1(n8371), .A2(n8370), .ZN(n8369) );
  INV_X1 U6586 ( .A(n5326), .ZN(n4631) );
  NAND2_X1 U6587 ( .A1(n4632), .A2(n10218), .ZN(n7366) );
  NAND3_X1 U6588 ( .A1(n5148), .A2(n7357), .A3(n5151), .ZN(n4632) );
  NAND2_X1 U6589 ( .A1(n8357), .A2(n6728), .ZN(n8342) );
  NAND2_X2 U6590 ( .A1(n8619), .A2(n6843), .ZN(n9803) );
  NAND2_X1 U6591 ( .A1(n8291), .A2(n5235), .ZN(n8357) );
  INV_X1 U6592 ( .A(n5194), .ZN(n5193) );
  NOR2_X1 U6593 ( .A1(n6941), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U6594 ( .A1(n4682), .A2(n4680), .ZN(n10002) );
  NAND2_X1 U6595 ( .A1(n9824), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U6596 ( .A1(n5908), .A2(n6058), .ZN(n6134) );
  XNOR2_X1 U6597 ( .A(n6952), .B(n6991), .ZN(n7529) );
  NAND2_X1 U6598 ( .A1(n7464), .A2(n6951), .ZN(n6952) );
  INV_X1 U6599 ( .A(n8929), .ZN(n4634) );
  NAND2_X1 U6600 ( .A1(n7587), .A2(n6946), .ZN(n6947) );
  NAND2_X1 U6601 ( .A1(n8576), .A2(n8577), .ZN(n8575) );
  NAND2_X2 U6602 ( .A1(n7865), .A2(n6959), .ZN(n6960) );
  OAI21_X1 U6603 ( .B1(n7943), .B2(n4867), .A(n4865), .ZN(n6963) );
  NAND2_X1 U6604 ( .A1(n6941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4994) );
  NAND2_X2 U6605 ( .A1(n5960), .A2(n5972), .ZN(n7919) );
  NAND2_X1 U6606 ( .A1(n4920), .A2(n8578), .ZN(n4687) );
  NAND2_X1 U6607 ( .A1(n4663), .A2(n4973), .ZN(n5908) );
  NAND2_X1 U6608 ( .A1(n4637), .A2(n4464), .ZN(n6056) );
  OAI211_X1 U6609 ( .C1(n6046), .C2(n6047), .A(n6045), .B(n9068), .ZN(n4637)
         );
  NAND2_X1 U6610 ( .A1(n4980), .A2(n4981), .ZN(n4747) );
  INV_X1 U6611 ( .A(n6933), .ZN(n4749) );
  NOR2_X1 U6612 ( .A1(n7872), .A2(n6925), .ZN(n6926) );
  AND2_X1 U6613 ( .A1(n7356), .A2(n8637), .ZN(n5151) );
  NAND2_X1 U6614 ( .A1(n5389), .A2(n5388), .ZN(n4641) );
  AND2_X1 U6615 ( .A1(n4641), .A2(n4453), .ZN(n5390) );
  NAND2_X1 U6616 ( .A1(n5347), .A2(n4643), .ZN(n4642) );
  NAND2_X2 U6617 ( .A1(n6075), .A2(n6142), .ZN(n6884) );
  NAND2_X1 U6618 ( .A1(n4971), .A2(n4970), .ZN(n4644) );
  NAND2_X1 U6619 ( .A1(n4645), .A2(n5383), .ZN(n5391) );
  AND2_X1 U6620 ( .A1(n5382), .A2(n5388), .ZN(n4645) );
  XNOR2_X1 U6621 ( .A(n10155), .B(n4651), .ZN(ADD_1068_U4) );
  XNOR2_X1 U6622 ( .A(n10275), .B(n9013), .ZN(ADD_1068_U55) );
  NAND2_X1 U6623 ( .A1(n8985), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8999) );
  AOI21_X1 U6624 ( .B1(n8932), .B2(n8930), .A(n8931), .ZN(n8934) );
  OR2_X1 U6625 ( .A1(n7074), .A2(n7071), .ZN(n7563) );
  NAND2_X1 U6626 ( .A1(n9542), .A2(n7235), .ZN(n7239) );
  NAND2_X1 U6627 ( .A1(n5573), .A2(n5572), .ZN(n9180) );
  NAND2_X1 U6628 ( .A1(n4823), .A2(n5739), .ZN(n9073) );
  NAND3_X1 U6629 ( .A1(n4809), .A2(n4808), .A3(n4807), .ZN(n4806) );
  NAND2_X1 U6630 ( .A1(n7124), .A2(n7123), .ZN(n7930) );
  NAND2_X1 U6631 ( .A1(n6421), .A2(n4491), .ZN(n6432) );
  NAND3_X1 U6632 ( .A1(n6596), .A2(n7346), .A3(n6834), .ZN(n6599) );
  NAND2_X1 U6633 ( .A1(n7406), .A2(n4414), .ZN(n4654) );
  NAND2_X1 U6634 ( .A1(n4833), .A2(n8433), .ZN(n6656) );
  NAND2_X1 U6635 ( .A1(n4897), .A2(n4751), .ZN(n6393) );
  NAND2_X1 U6636 ( .A1(n6381), .A2(n6351), .ZN(n4754) );
  NOR2_X1 U6637 ( .A1(n5248), .A2(n6715), .ZN(n6790) );
  OAI21_X1 U6638 ( .B1(n4894), .B2(n4892), .A(n6476), .ZN(n4891) );
  NAND2_X1 U6639 ( .A1(n10081), .A2(n10225), .ZN(n4661) );
  NAND2_X1 U6640 ( .A1(n10009), .A2(n4662), .ZN(n10081) );
  NAND2_X1 U6641 ( .A1(n6634), .A2(n5027), .ZN(n4997) );
  INV_X1 U6642 ( .A(n9036), .ZN(n4663) );
  NAND2_X1 U6643 ( .A1(n5212), .A2(n5213), .ZN(n9036) );
  NAND2_X1 U6644 ( .A1(n9078), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U6645 ( .A1(n4664), .A2(n4531), .ZN(n6150) );
  XNOR2_X1 U6646 ( .A(n6145), .B(n5884), .ZN(n4664) );
  NAND2_X1 U6647 ( .A1(n9158), .A2(n6012), .ZN(n5902) );
  NAND2_X1 U6648 ( .A1(n4986), .A2(n4988), .ZN(n4985) );
  NAND2_X1 U6649 ( .A1(n6920), .A2(n7470), .ZN(n7468) );
  NAND2_X1 U6650 ( .A1(n4700), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8932) );
  OAI21_X1 U6651 ( .B1(n9434), .B2(n9435), .A(n9598), .ZN(n4692) );
  NAND2_X1 U6652 ( .A1(n5387), .A2(n5368), .ZN(n5377) );
  NAND3_X1 U6653 ( .A1(n4687), .A2(n7043), .A3(n4665), .ZN(P2_U3201) );
  NAND2_X1 U6654 ( .A1(n7179), .A2(n4486), .ZN(n5014) );
  NAND3_X1 U6655 ( .A1(n4965), .A2(n4966), .A3(n4832), .ZN(n5281) );
  NAND2_X1 U6656 ( .A1(n5329), .A2(n5383), .ZN(n5346) );
  NAND2_X1 U6657 ( .A1(n7850), .A2(n5890), .ZN(n7845) );
  NAND2_X1 U6658 ( .A1(n5210), .A2(n5205), .ZN(n4667) );
  INV_X1 U6659 ( .A(n5834), .ZN(n5832) );
  INV_X1 U6660 ( .A(n5125), .ZN(n5123) );
  NAND2_X1 U6661 ( .A1(n5852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5854) );
  INV_X1 U6662 ( .A(n5122), .ZN(n5121) );
  NAND2_X1 U6663 ( .A1(n5346), .A2(n5384), .ZN(n5355) );
  NAND2_X1 U6664 ( .A1(n6025), .A2(n4460), .ZN(n4912) );
  NAND2_X1 U6665 ( .A1(n4968), .A2(n6100), .ZN(n4911) );
  AND2_X1 U6666 ( .A1(n9712), .A2(n9720), .ZN(n4677) );
  XNOR2_X1 U6667 ( .A(n9712), .B(n7995), .ZN(n9713) );
  NAND2_X2 U6668 ( .A1(n9858), .A2(n6837), .ZN(n9842) );
  NAND2_X1 U6669 ( .A1(n5416), .A2(n4686), .ZN(n4685) );
  OAI21_X1 U6670 ( .B1(n5284), .B2(n5347), .A(n4750), .ZN(n5288) );
  NAND3_X1 U6671 ( .A1(n4985), .A2(n6935), .A3(n4984), .ZN(n6937) );
  NAND3_X1 U6672 ( .A1(n4989), .A2(n8998), .A3(n4987), .ZN(n4984) );
  INV_X1 U6673 ( .A(n8920), .ZN(n4700) );
  AND2_X2 U6674 ( .A1(n4741), .A2(n6633), .ZN(n6454) );
  NAND3_X1 U6675 ( .A1(n4692), .A2(n9439), .A3(n4691), .ZN(P1_U3214) );
  NAND2_X1 U6676 ( .A1(n5185), .A2(n5184), .ZN(n5952) );
  AND2_X2 U6677 ( .A1(n5828), .A2(n5244), .ZN(n4966) );
  NOR2_X1 U6678 ( .A1(n6893), .A2(n5202), .ZN(n5201) );
  NAND3_X1 U6679 ( .A1(n5316), .A2(n5317), .A3(n5319), .ZN(n5323) );
  BUF_X1 U6680 ( .A(n7370), .Z(n4696) );
  NAND2_X1 U6681 ( .A1(n4907), .A2(n5479), .ZN(n5827) );
  NAND2_X1 U6682 ( .A1(n5881), .A2(n5882), .ZN(n5852) );
  NOR3_X1 U6683 ( .A1(n6133), .A2(n4728), .A3(n6107), .ZN(n4727) );
  NAND2_X1 U6684 ( .A1(n4749), .A2(n8991), .ZN(n4989) );
  OAI21_X1 U6685 ( .B1(n6932), .B2(n9302), .A(n8976), .ZN(n6933) );
  NAND2_X1 U6686 ( .A1(n7949), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7948) );
  AOI21_X1 U6687 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7404), .A(n8095), .ZN(
        n6928) );
  OR2_X1 U6688 ( .A1(n7506), .A2(n10256), .ZN(n7504) );
  NAND2_X1 U6689 ( .A1(n7504), .A2(n6917), .ZN(n7591) );
  NAND2_X1 U6690 ( .A1(n4994), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4993) );
  AOI21_X1 U6691 ( .B1(n6926), .B2(n7005), .A(n6927), .ZN(n7949) );
  INV_X1 U6692 ( .A(n4755), .ZN(n4723) );
  NAND2_X1 U6693 ( .A1(n6761), .A2(n6760), .ZN(n8409) );
  NAND2_X1 U6694 ( .A1(n5183), .A2(n5773), .ZN(n9049) );
  NAND2_X1 U6695 ( .A1(n4806), .A2(n4502), .ZN(n5432) );
  NAND2_X1 U6696 ( .A1(n6972), .A2(n6971), .ZN(n6973) );
  NAND2_X1 U6697 ( .A1(n6952), .A2(n7535), .ZN(n6953) );
  INV_X1 U6698 ( .A(n6961), .ZN(n4867) );
  NAND2_X1 U6699 ( .A1(n9841), .A2(n6839), .ZN(n5238) );
  NAND2_X1 U6700 ( .A1(n10080), .A2(n10218), .ZN(n4708) );
  NAND2_X1 U6701 ( .A1(n5222), .A2(n5220), .ZN(n9197) );
  NAND2_X1 U6702 ( .A1(n6897), .A2(n4712), .ZN(n9029) );
  NOR2_X2 U6703 ( .A1(n9029), .A2(n5242), .ZN(n7335) );
  INV_X1 U6704 ( .A(n8998), .ZN(n4986) );
  OR2_X2 U6705 ( .A1(n10008), .A2(n9827), .ZN(n6840) );
  OAI21_X1 U6706 ( .B1(n9197), .B2(n5899), .A(n5898), .ZN(n5901) );
  NAND2_X1 U6707 ( .A1(n5064), .A2(n5742), .ZN(n5758) );
  NAND2_X1 U6708 ( .A1(n4847), .A2(n4845), .ZN(n8620) );
  INV_X4 U6709 ( .A(n5357), .ZN(n6087) );
  NAND2_X1 U6710 ( .A1(n6839), .A2(n4850), .ZN(n4849) );
  NAND2_X1 U6711 ( .A1(n6170), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6571) );
  BUF_X4 U6712 ( .A(n5347), .Z(n7378) );
  OAI21_X1 U6713 ( .B1(n5203), .B2(n5201), .A(n5200), .ZN(n5199) );
  NOR2_X2 U6714 ( .A1(n6201), .A2(n4792), .ZN(n6634) );
  NAND4_X1 U6715 ( .A1(n6128), .A2(n4487), .A3(n4736), .A4(n4735), .ZN(n6129)
         );
  NAND2_X1 U6716 ( .A1(n4837), .A2(n4836), .ZN(n4835) );
  NAND2_X2 U6717 ( .A1(n9549), .A2(n9548), .ZN(n7179) );
  INV_X1 U6718 ( .A(n6290), .ZN(n6200) );
  NAND2_X1 U6719 ( .A1(n5011), .A2(n7155), .ZN(n8479) );
  NAND2_X1 U6720 ( .A1(n5238), .A2(n6840), .ZN(n9825) );
  NAND3_X1 U6721 ( .A1(n6974), .A2(P2_REG2_REG_15__SCAN_IN), .A3(n8960), .ZN(
        n8962) );
  NAND2_X1 U6722 ( .A1(n4746), .A2(n5895), .ZN(n8080) );
  OAI211_X1 U6723 ( .C1(n5198), .C2(n7919), .A(n5197), .B(n5893), .ZN(n4746)
         );
  INV_X1 U6724 ( .A(n9035), .ZN(n6896) );
  NAND2_X1 U6725 ( .A1(n4982), .A2(n4980), .ZN(n4748) );
  NAND2_X1 U6726 ( .A1(n4991), .A2(n8971), .ZN(n6931) );
  NAND2_X1 U6727 ( .A1(n7728), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7870) );
  NAND2_X1 U6728 ( .A1(n5355), .A2(n5354), .ZN(n5368) );
  NAND2_X1 U6729 ( .A1(n5347), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4750) );
  AOI21_X1 U6730 ( .B1(n6432), .B2(n6730), .A(n6733), .ZN(n4894) );
  NAND2_X1 U6731 ( .A1(n4891), .A2(n4890), .ZN(n4889) );
  NAND2_X1 U6732 ( .A1(n4889), .A2(n4885), .ZN(n6489) );
  NAND2_X1 U6733 ( .A1(n5204), .A2(n5199), .ZN(n6145) );
  NAND2_X1 U6734 ( .A1(n5541), .A2(n4758), .ZN(n5601) );
  NAND2_X1 U6735 ( .A1(n5804), .A2(n4761), .ZN(n6096) );
  NAND2_X1 U6736 ( .A1(n5804), .A2(n5803), .ZN(n5820) );
  NAND2_X1 U6737 ( .A1(n5424), .A2(n4765), .ZN(n5484) );
  NAND2_X1 U6738 ( .A1(n5618), .A2(n4520), .ZN(n5683) );
  NAND3_X1 U6739 ( .A1(n7896), .A2(n5361), .A3(n5340), .ZN(n5402) );
  NAND4_X1 U6740 ( .A1(n7896), .A2(n5340), .A3(n5361), .A4(n4771), .ZN(n5425)
         );
  NAND2_X1 U6741 ( .A1(n7378), .A2(n7409), .ZN(n4772) );
  NOR2_X1 U6742 ( .A1(n6777), .A2(n4775), .ZN(n4774) );
  INV_X2 U6743 ( .A(n7354), .ZN(n4781) );
  NAND2_X2 U6744 ( .A1(n5627), .A2(n5626), .ZN(n5640) );
  NAND4_X2 U6745 ( .A1(n6305), .A2(n6303), .A3(n6304), .A4(n4783), .ZN(n9621)
         );
  OR2_X2 U6746 ( .A1(n4792), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4789) );
  NAND3_X1 U6747 ( .A1(n5027), .A2(n4790), .A3(n4741), .ZN(n10108) );
  INV_X1 U6748 ( .A(n6819), .ZN(n4801) );
  NAND2_X1 U6749 ( .A1(n4799), .A2(n4798), .ZN(n9897) );
  NAND2_X1 U6750 ( .A1(n4811), .A2(n7911), .ZN(n4808) );
  AND2_X1 U6751 ( .A1(n5374), .A2(n6115), .ZN(n4811) );
  NAND3_X1 U6752 ( .A1(n4809), .A2(n4808), .A3(n6114), .ZN(n8058) );
  NAND2_X1 U6753 ( .A1(n5181), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U6754 ( .A1(n5181), .A2(n5180), .ZN(n4823) );
  NAND2_X1 U6755 ( .A1(n4826), .A2(n4824), .ZN(n5179) );
  INV_X1 U6756 ( .A(n5492), .ZN(n8527) );
  NAND2_X1 U6757 ( .A1(n9187), .A2(n5571), .ZN(n5573) );
  NAND2_X1 U6758 ( .A1(n6883), .A2(n4827), .ZN(n6891) );
  NAND2_X1 U6759 ( .A1(n4831), .A2(n4830), .ZN(n4827) );
  NAND2_X1 U6760 ( .A1(n5791), .A2(n5790), .ZN(n9038) );
  NOR2_X1 U6761 ( .A1(n6884), .A2(n6881), .ZN(n4830) );
  NAND2_X1 U6762 ( .A1(n4833), .A2(n6806), .ZN(n8437) );
  NAND2_X1 U6763 ( .A1(n6654), .A2(n4833), .ZN(n6758) );
  NAND2_X2 U6764 ( .A1(n6378), .A2(n6377), .ZN(n4833) );
  NAND3_X1 U6765 ( .A1(n5414), .A2(n5234), .A3(n5466), .ZN(n4834) );
  INV_X1 U6766 ( .A(n6734), .ZN(n4836) );
  AND2_X1 U6767 ( .A1(n9884), .A2(n9904), .ZN(n4839) );
  NAND2_X1 U6768 ( .A1(n9842), .A2(n4848), .ZN(n4847) );
  NAND3_X1 U6769 ( .A1(n4856), .A2(n4860), .A3(n4855), .ZN(n5412) );
  NAND3_X1 U6770 ( .A1(n5283), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_DATAO_REG_7__SCAN_IN), .ZN(n4855) );
  NAND3_X1 U6771 ( .A1(n4862), .A2(n4863), .A3(P2_DATAO_REG_7__SCAN_IN), .ZN(
        n4856) );
  NAND3_X1 U6772 ( .A1(n4857), .A2(n5282), .A3(P1_DATAO_REG_7__SCAN_IN), .ZN(
        n4860) );
  AOI21_X2 U6773 ( .B1(n6961), .B2(n10315), .A(n4866), .ZN(n4865) );
  XNOR2_X2 U6774 ( .A(n6960), .B(n7005), .ZN(n7943) );
  INV_X1 U6775 ( .A(n6953), .ZN(n4870) );
  NAND2_X1 U6776 ( .A1(n7588), .A2(n7589), .ZN(n7587) );
  INV_X1 U6777 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U6778 ( .A1(n6974), .A2(n8960), .ZN(n8947) );
  NAND2_X1 U6779 ( .A1(n6972), .A2(n4528), .ZN(n8960) );
  INV_X1 U6780 ( .A(n6976), .ZN(n4881) );
  INV_X1 U6781 ( .A(n6595), .ZN(n6592) );
  OAI21_X1 U6782 ( .B1(n4440), .B2(n6554), .A(n6568), .ZN(n4884) );
  NAND3_X1 U6783 ( .A1(n6676), .A2(n4436), .A3(n6735), .ZN(n4886) );
  NAND2_X1 U6784 ( .A1(n4897), .A2(n4895), .ZN(n6478) );
  NAND3_X1 U6785 ( .A1(n6352), .A2(n6353), .A3(n4898), .ZN(n4897) );
  OAI21_X1 U6786 ( .B1(n8404), .B2(n6319), .A(n6663), .ZN(n4905) );
  INV_X2 U6787 ( .A(n6449), .ZN(n6263) );
  NAND2_X1 U6788 ( .A1(n8613), .A2(n8661), .ZN(n6449) );
  NOR2_X2 U6789 ( .A1(n5827), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4965) );
  NAND3_X1 U6790 ( .A1(n5262), .A2(n5331), .A3(n4875), .ZN(n4908) );
  NAND2_X1 U6791 ( .A1(n6002), .A2(n4506), .ZN(n4914) );
  OR2_X1 U6792 ( .A1(n4971), .A2(n4917), .ZN(n4916) );
  XNOR2_X2 U6793 ( .A(n4918), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5269) );
  OR2_X2 U6794 ( .A1(n9413), .A2(n5267), .ZN(n4918) );
  AOI21_X1 U6795 ( .B1(n7628), .B2(n4924), .A(n4922), .ZN(n4921) );
  NOR2_X1 U6796 ( .A1(n7628), .A2(n7627), .ZN(n7726) );
  NAND2_X1 U6797 ( .A1(n8937), .A2(n4439), .ZN(n4939) );
  NOR2_X1 U6798 ( .A1(n7023), .A2(n8968), .ZN(n4947) );
  NAND2_X1 U6799 ( .A1(n7021), .A2(n7022), .ZN(n4948) );
  NAND4_X1 U6800 ( .A1(n5977), .A2(n4954), .A3(n8083), .A4(n5982), .ZN(n4953)
         );
  NAND2_X1 U6801 ( .A1(n4962), .A2(n4959), .ZN(n4956) );
  AOI21_X1 U6802 ( .B1(n5512), .B2(n4959), .A(n4498), .ZN(n4958) );
  NAND3_X1 U6803 ( .A1(n4963), .A2(n4966), .A3(n4961), .ZN(n4960) );
  NOR2_X1 U6804 ( .A1(n5512), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4961) );
  INV_X1 U6805 ( .A(n4963), .ZN(n4962) );
  INV_X1 U6806 ( .A(n4980), .ZN(n8569) );
  INV_X1 U6807 ( .A(n4982), .ZN(n4979) );
  NAND2_X1 U6808 ( .A1(n4997), .A2(n4996), .ZN(n6157) );
  AND2_X1 U6809 ( .A1(n4997), .A2(n6647), .ZN(n6869) );
  NAND3_X1 U6810 ( .A1(n5016), .A2(n5018), .A3(n5015), .ZN(n5013) );
  NAND2_X1 U6811 ( .A1(n8152), .A2(n7135), .ZN(n7144) );
  NOR2_X2 U6812 ( .A1(n6290), .A2(n6156), .ZN(n5027) );
  NOR3_X2 U6813 ( .A1(n9829), .A2(n5037), .A3(n7359), .ZN(n5039) );
  INV_X1 U6814 ( .A(n5039), .ZN(n9794) );
  INV_X1 U6815 ( .A(n5042), .ZN(n9852) );
  INV_X1 U6816 ( .A(n5047), .ZN(n8592) );
  NAND2_X1 U6817 ( .A1(n7378), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6818 ( .A1(n5469), .A2(n5055), .ZN(n5052) );
  NAND2_X1 U6819 ( .A1(n5467), .A2(SI_8_), .ZN(n5055) );
  NAND2_X1 U6820 ( .A1(n5057), .A2(n5056), .ZN(n5627) );
  NAND2_X1 U6821 ( .A1(n5741), .A2(n5065), .ZN(n5061) );
  NAND2_X1 U6822 ( .A1(n5061), .A2(n5062), .ZN(n5775) );
  NAND2_X1 U6823 ( .A1(n5741), .A2(n5740), .ZN(n5064) );
  NAND2_X1 U6824 ( .A1(n5084), .A2(n5085), .ZN(n8668) );
  NAND2_X1 U6825 ( .A1(n8549), .A2(n8553), .ZN(n5084) );
  OAI211_X2 U6826 ( .C1(n5357), .C2(n7381), .A(n5088), .B(n5087), .ZN(n7857)
         );
  OR2_X1 U6827 ( .A1(n5358), .A2(n5285), .ZN(n5088) );
  NAND2_X2 U6828 ( .A1(n6938), .A2(n5848), .ZN(n6913) );
  OAI21_X1 U6829 ( .B1(n4596), .B2(n5092), .A(n5090), .ZN(n8750) );
  OAI21_X1 U6830 ( .B1(n4596), .B2(n8812), .A(n8696), .ZN(n8869) );
  NAND2_X1 U6831 ( .A1(n8812), .A2(n8696), .ZN(n5093) );
  NAND3_X1 U6832 ( .A1(n5094), .A2(n7758), .A3(n7810), .ZN(n7811) );
  NAND2_X1 U6833 ( .A1(n7757), .A2(n7756), .ZN(n7810) );
  OR2_X1 U6834 ( .A1(n8847), .A2(n4441), .ZN(n5095) );
  NAND2_X1 U6835 ( .A1(n8847), .A2(n5100), .ZN(n5099) );
  NAND3_X1 U6836 ( .A1(n5107), .A2(n8795), .A3(n5105), .ZN(n5104) );
  NAND2_X1 U6837 ( .A1(n8891), .A2(n8691), .ZN(n5116) );
  NAND2_X1 U6838 ( .A1(n5116), .A2(n5113), .ZN(n8694) );
  NAND2_X1 U6839 ( .A1(n6281), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6267) );
  INV_X1 U6840 ( .A(n6805), .ZN(n5129) );
  NAND2_X1 U6841 ( .A1(n5157), .A2(n5155), .ZN(n5960) );
  AND2_X1 U6842 ( .A1(n5345), .A2(n5343), .ZN(n5158) );
  NAND2_X1 U6843 ( .A1(n9180), .A2(n4429), .ZN(n5159) );
  NAND2_X1 U6844 ( .A1(n5159), .A2(n5160), .ZN(n9160) );
  NAND2_X1 U6845 ( .A1(n6882), .A2(n4489), .ZN(n5172) );
  NAND3_X1 U6846 ( .A1(n5176), .A2(n5173), .A3(n5172), .ZN(n9260) );
  NAND2_X1 U6847 ( .A1(n5179), .A2(n4499), .ZN(n9106) );
  NAND2_X1 U6848 ( .A1(n5183), .A2(n5182), .ZN(n5791) );
  NAND2_X2 U6849 ( .A1(n5952), .A2(n5950), .ZN(n7847) );
  NAND2_X2 U6850 ( .A1(n7756), .A2(n7857), .ZN(n5950) );
  INV_X1 U6851 ( .A(n7857), .ZN(n5184) );
  OR2_X1 U6852 ( .A1(n5404), .A2(n5299), .ZN(n5187) );
  NAND2_X1 U6853 ( .A1(n9193), .A2(n5193), .ZN(n5189) );
  NAND2_X1 U6854 ( .A1(n5196), .A2(n7911), .ZN(n7906) );
  NAND2_X1 U6855 ( .A1(n5198), .A2(n5892), .ZN(n5196) );
  NAND2_X1 U6856 ( .A1(n4724), .A2(n7911), .ZN(n5197) );
  NAND2_X1 U6857 ( .A1(n9235), .A2(n5956), .ZN(n5198) );
  NAND2_X1 U6858 ( .A1(n5907), .A2(n5211), .ZN(n5212) );
  INV_X1 U6859 ( .A(n6052), .ZN(n5217) );
  INV_X1 U6860 ( .A(n5216), .ZN(n5215) );
  NAND2_X1 U6861 ( .A1(n5907), .A2(n6044), .ZN(n9067) );
  OAI21_X1 U6862 ( .B1(n5216), .B2(n6049), .A(n5942), .ZN(n5214) );
  NOR2_X2 U6863 ( .A1(n5280), .A2(n5219), .ZN(n9413) );
  NAND3_X1 U6864 ( .A1(n5278), .A2(n4832), .A3(n5268), .ZN(n5219) );
  NAND2_X1 U6865 ( .A1(n8163), .A2(n5223), .ZN(n5222) );
  NAND2_X1 U6866 ( .A1(n9803), .A2(n4459), .ZN(n5225) );
  OAI211_X1 U6867 ( .C1(n9803), .C2(n5229), .A(n5226), .B(n5225), .ZN(n7351)
         );
  INV_X1 U6868 ( .A(n5449), .ZN(n5234) );
  NAND2_X1 U6869 ( .A1(n5234), .A2(n5466), .ZN(n5233) );
  OAI21_X2 U6870 ( .B1(n5416), .B2(n5233), .A(n4472), .ZN(n5452) );
  INV_X1 U6871 ( .A(n6724), .ZN(n8292) );
  INV_X1 U6872 ( .A(n9826), .ZN(n6841) );
  NAND2_X1 U6873 ( .A1(n9325), .A2(n9253), .ZN(n9045) );
  AND2_X1 U6874 ( .A1(n5550), .A2(n5536), .ZN(n7644) );
  CLKBUF_X1 U6875 ( .A(n7653), .Z(n7689) );
  NAND2_X1 U6876 ( .A1(n6793), .A2(n6260), .ZN(n6794) );
  OR2_X1 U6877 ( .A1(n7105), .A2(n6320), .ZN(n6718) );
  INV_X1 U6878 ( .A(n9959), .ZN(n9970) );
  INV_X1 U6879 ( .A(n6607), .ZN(n6556) );
  NAND2_X1 U6880 ( .A1(n7339), .A2(n10225), .ZN(n7343) );
  NAND2_X1 U6881 ( .A1(n9260), .A2(n9259), .ZN(n9263) );
  INV_X1 U6882 ( .A(n7756), .ZN(n9242) );
  INV_X1 U6883 ( .A(n5416), .ZN(n5413) );
  NAND2_X1 U6884 ( .A1(n5380), .A2(SI_6_), .ZN(n5411) );
  OAI21_X1 U6885 ( .B1(n7370), .B2(n5379), .A(n5378), .ZN(n5380) );
  NAND2_X1 U6886 ( .A1(n7370), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5378) );
  INV_X1 U6887 ( .A(n8471), .ZN(n6378) );
  NOR2_X1 U6888 ( .A1(n10190), .A2(n4422), .ZN(n7336) );
  INV_X1 U6889 ( .A(n4422), .ZN(n8425) );
  OR2_X1 U6890 ( .A1(n9344), .A2(n9099), .ZN(n5239) );
  AND2_X1 U6891 ( .A1(n8206), .A2(n10190), .ZN(n10215) );
  OR2_X1 U6892 ( .A1(n10254), .A2(n10337), .ZN(n5241) );
  AND2_X1 U6893 ( .A1(n6896), .A2(n10234), .ZN(n5242) );
  AND2_X1 U6894 ( .A1(n6785), .A2(n9781), .ZN(n5243) );
  AND3_X1 U6895 ( .A1(n5261), .A2(n5260), .A3(n5259), .ZN(n5244) );
  AND2_X1 U6896 ( .A1(n7825), .A2(n7823), .ZN(n5245) );
  INV_X1 U6897 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5379) );
  AND2_X1 U6898 ( .A1(n7354), .A2(n7345), .ZN(n5246) );
  OR2_X1 U6899 ( .A1(n8574), .A2(n9314), .ZN(n5247) );
  AND2_X1 U6900 ( .A1(n6783), .A2(n6638), .ZN(n5248) );
  INV_X1 U6901 ( .A(n9948), .ZN(n6815) );
  INV_X1 U6902 ( .A(SI_19_), .ZN(n5644) );
  NOR2_X1 U6903 ( .A1(n10004), .A2(n9614), .ZN(n5249) );
  INV_X1 U6904 ( .A(n6855), .ZN(n9829) );
  OR2_X1 U6905 ( .A1(n9268), .A2(n9062), .ZN(n5250) );
  NOR4_X1 U6906 ( .A1(n9915), .A2(n9929), .A3(n9948), .A4(n6770), .ZN(n5251)
         );
  INV_X1 U6907 ( .A(n8588), .ZN(n6732) );
  AND2_X1 U6908 ( .A1(n7894), .A2(n8287), .ZN(n5252) );
  AND2_X2 U6909 ( .A1(n6906), .A2(n6905), .ZN(n10266) );
  INV_X1 U6910 ( .A(n10266), .ZN(n6909) );
  NAND2_X1 U6911 ( .A1(n7737), .A2(n5910), .ZN(n9244) );
  INV_X2 U6912 ( .A(n10255), .ZN(n10254) );
  INV_X1 U6913 ( .A(n8638), .ZN(n7344) );
  AND2_X1 U6914 ( .A1(n5911), .A2(n5241), .ZN(n5253) );
  AND2_X1 U6915 ( .A1(n9122), .A2(n9107), .ZN(n5691) );
  INV_X1 U6916 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5256) );
  INV_X1 U6917 ( .A(n9039), .ZN(n6879) );
  NAND4_X1 U6918 ( .A1(n5560), .A2(n5593), .A3(n5595), .A4(n5256), .ZN(n5257)
         );
  INV_X1 U6919 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6922) );
  AND2_X1 U6920 ( .A1(n7748), .A2(n7747), .ZN(n7750) );
  NOR2_X1 U6921 ( .A1(n6992), .A2(n6922), .ZN(n6923) );
  NAND2_X1 U6922 ( .A1(n6885), .A2(n6880), .ZN(n6881) );
  AND2_X1 U6923 ( .A1(n8208), .A2(n6804), .ZN(n6802) );
  INV_X1 U6924 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5609) );
  INV_X1 U6925 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5540) );
  INV_X1 U6926 ( .A(n7309), .ZN(n7307) );
  INV_X1 U6927 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6413) );
  INV_X1 U6928 ( .A(SI_26_), .ZN(n5778) );
  INV_X1 U6929 ( .A(SI_20_), .ZN(n5698) );
  INV_X1 U6930 ( .A(n7809), .ZN(n8684) );
  AND2_X1 U6931 ( .A1(n8785), .A2(n8675), .ZN(n8676) );
  INV_X1 U6932 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10410) );
  OR2_X1 U6933 ( .A1(n7400), .A2(n5880), .ZN(n5916) );
  INV_X1 U6934 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5799) );
  OR2_X1 U6935 ( .A1(n7766), .A2(n7745), .ZN(n7849) );
  INV_X1 U6936 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5278) );
  INV_X1 U6937 ( .A(n8305), .ZN(n7154) );
  NOR2_X1 U6938 ( .A1(n7310), .A2(n9578), .ZN(n7308) );
  INV_X1 U6939 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6521) );
  INV_X1 U6940 ( .A(n4421), .ZN(n7298) );
  OR2_X1 U6941 ( .A1(n10211), .A2(n7296), .ZN(n7320) );
  NOR2_X1 U6942 ( .A1(n10172), .A2(n10169), .ZN(n10173) );
  AND2_X1 U6943 ( .A1(n5549), .A2(n5533), .ZN(n5534) );
  INV_X1 U6944 ( .A(n5477), .ZN(n5475) );
  INV_X1 U6945 ( .A(n6633), .ZN(n6306) );
  INV_X1 U6946 ( .A(n9161), .ZN(n8754) );
  INV_X1 U6947 ( .A(n9136), .ZN(n8776) );
  INV_X1 U6948 ( .A(n9089), .ZN(n8823) );
  NAND2_X1 U6949 ( .A1(n8681), .A2(n8729), .ZN(n8723) );
  INV_X1 U6950 ( .A(n8894), .ZN(n8883) );
  OR2_X1 U6951 ( .A1(n4711), .A2(n5339), .ZN(n5345) );
  OR2_X1 U6952 ( .A1(P2_U3150), .A2(n7039), .ZN(n9014) );
  INV_X1 U6953 ( .A(n8906), .ZN(n9146) );
  AND2_X1 U6954 ( .A1(n5983), .A2(n5988), .ZN(n8083) );
  NAND2_X1 U6955 ( .A1(n6936), .A2(n8287), .ZN(n9249) );
  AND2_X1 U6956 ( .A1(n5919), .A2(n6910), .ZN(n6902) );
  NAND2_X1 U6957 ( .A1(n9041), .A2(n9040), .ZN(n9042) );
  OR2_X1 U6958 ( .A1(n7762), .A2(n6910), .ZN(n9145) );
  OR2_X1 U6959 ( .A1(n9249), .A2(n6148), .ZN(n10243) );
  XNOR2_X1 U6960 ( .A(n6636), .B(n6639), .ZN(n7390) );
  INV_X1 U6961 ( .A(n9619), .ZN(n8486) );
  INV_X1 U6962 ( .A(n6573), .ZN(n6585) );
  INV_X1 U6963 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7782) );
  AND2_X1 U6964 ( .A1(n7394), .A2(n7393), .ZN(n7432) );
  AND2_X1 U6965 ( .A1(n6771), .A2(n6836), .ZN(n9869) );
  AND2_X1 U6966 ( .A1(n6745), .A2(n6746), .ZN(n9904) );
  INV_X1 U6967 ( .A(n9618), .ZN(n8591) );
  NAND2_X1 U6968 ( .A1(n8138), .A2(n6261), .ZN(n7839) );
  OR2_X1 U6969 ( .A1(n8234), .A2(n6833), .ZN(n8206) );
  INV_X1 U6970 ( .A(n8210), .ZN(n8332) );
  INV_X1 U6971 ( .A(n7105), .ZN(n8225) );
  NAND2_X1 U6972 ( .A1(n8425), .A2(n8505), .ZN(n7311) );
  AND2_X1 U6973 ( .A1(n5776), .A2(n5763), .ZN(n5774) );
  AND2_X1 U6974 ( .A1(n5574), .A2(n5554), .ZN(n5555) );
  INV_X1 U6975 ( .A(n5355), .ZN(n5352) );
  NAND2_X1 U6976 ( .A1(n7764), .A2(n7763), .ZN(n8896) );
  AND2_X1 U6977 ( .A1(n7764), .A2(n7762), .ZN(n8894) );
  INV_X1 U6978 ( .A(n8896), .ZN(n8880) );
  AOI21_X1 U6979 ( .B1(n9114), .B2(n4411), .A(n5678), .ZN(n9121) );
  INV_X1 U6980 ( .A(n6938), .ZN(n7035) );
  AND2_X1 U6981 ( .A1(n7034), .A2(n9420), .ZN(n7414) );
  OAI21_X1 U6982 ( .B1(n9264), .B2(n9233), .A(n5929), .ZN(n5930) );
  INV_X1 U6983 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10566) );
  INV_X1 U6984 ( .A(n9233), .ZN(n9155) );
  NAND2_X1 U6985 ( .A1(n7401), .A2(n6900), .ZN(n9207) );
  XNOR2_X1 U6986 ( .A(n9261), .B(n9039), .ZN(n8763) );
  INV_X1 U6987 ( .A(n9298), .ZN(n9315) );
  OAI21_X1 U6988 ( .B1(n9264), .B2(n9403), .A(n5253), .ZN(n5912) );
  INV_X1 U6989 ( .A(n10249), .ZN(n10241) );
  NAND2_X1 U6990 ( .A1(n9244), .A2(n10243), .ZN(n10250) );
  XNOR2_X1 U6991 ( .A(n5881), .B(n5882), .ZN(n6911) );
  OR2_X1 U6992 ( .A1(n7390), .A2(n4410), .ZN(n7326) );
  INV_X1 U6993 ( .A(n9609), .ZN(n9576) );
  INV_X1 U6994 ( .A(n9584), .ZN(n9606) );
  OR2_X1 U6995 ( .A1(n9460), .A2(n6573), .ZN(n6538) );
  AND3_X1 U6996 ( .A1(n6463), .A2(n6462), .A3(n6461), .ZN(n9524) );
  INV_X1 U6997 ( .A(n9775), .ZN(n9773) );
  INV_X1 U6998 ( .A(n9786), .ZN(n9762) );
  INV_X1 U6999 ( .A(n10174), .ZN(n9971) );
  INV_X1 U7000 ( .A(n9938), .ZN(n9929) );
  INV_X1 U7001 ( .A(n7159), .ZN(n9489) );
  AND2_X1 U7002 ( .A1(n8206), .A2(n8136), .ZN(n8207) );
  NAND2_X1 U7003 ( .A1(n7336), .A2(n10104), .ZN(n9962) );
  INV_X1 U7004 ( .A(n7842), .ZN(n8280) );
  NOR2_X1 U7005 ( .A1(n10225), .A2(n10381), .ZN(n7358) );
  NOR2_X1 U7006 ( .A1(n8131), .A2(n7336), .ZN(n7337) );
  INV_X1 U7007 ( .A(n10215), .ZN(n10206) );
  OR2_X1 U7008 ( .A1(n6441), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6464) );
  AND2_X1 U7009 ( .A1(n5346), .A2(n5330), .ZN(n7372) );
  INV_X1 U7010 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10397) );
  INV_X1 U7011 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10439) );
  INV_X1 U7012 ( .A(n8899), .ZN(n8862) );
  AND2_X1 U7013 ( .A1(n7707), .A2(n7706), .ZN(n8889) );
  INV_X1 U7014 ( .A(n8729), .ZN(n9225) );
  MUX2_X1 U7015 ( .A(n7036), .B(n9003), .S(n7035), .Z(n8969) );
  INV_X1 U7016 ( .A(n8980), .ZN(n9006) );
  INV_X1 U7017 ( .A(n9253), .ZN(n9213) );
  NAND2_X1 U7018 ( .A1(n9253), .A2(n5926), .ZN(n9233) );
  INV_X1 U7019 ( .A(n9230), .ZN(n9153) );
  NAND2_X1 U7020 ( .A1(n10266), .A2(n10250), .ZN(n9313) );
  NAND2_X1 U7021 ( .A1(n10266), .A2(n10249), .ZN(n9298) );
  INV_X1 U7022 ( .A(n6137), .ZN(n9324) );
  OR2_X1 U7023 ( .A1(n10255), .A2(n8060), .ZN(n9403) );
  AND2_X1 U7024 ( .A1(n10253), .A2(n10252), .ZN(n10265) );
  AND2_X1 U7025 ( .A1(n5889), .A2(n5888), .ZN(n10255) );
  INV_X1 U7026 ( .A(n8609), .ZN(n7411) );
  INV_X1 U7027 ( .A(n6991), .ZN(n7535) );
  INV_X1 U7028 ( .A(n10008), .ZN(n9538) );
  INV_X1 U7029 ( .A(n9598), .ZN(n9578) );
  AND2_X1 U7030 ( .A1(n7313), .A2(n9962), .ZN(n9609) );
  AND2_X1 U7031 ( .A1(n6180), .A2(n6179), .ZN(n8112) );
  INV_X1 U7032 ( .A(n9779), .ZN(n9743) );
  NAND2_X1 U7033 ( .A1(n7395), .A2(n7431), .ZN(n9786) );
  OR2_X1 U7034 ( .A1(n10167), .A2(n9781), .ZN(n9801) );
  AOI21_X1 U7035 ( .B1(n7359), .B2(n9992), .A(n7358), .ZN(n7360) );
  NAND2_X1 U7036 ( .A1(n10225), .A2(n10211), .ZN(n10066) );
  AND2_X2 U7037 ( .A1(n7338), .A2(n7337), .ZN(n10225) );
  INV_X1 U7038 ( .A(n9816), .ZN(n10078) );
  INV_X1 U7039 ( .A(n9475), .ZN(n10092) );
  INV_X1 U7040 ( .A(n9555), .ZN(n10103) );
  INV_X1 U7041 ( .A(n10218), .ZN(n10217) );
  INV_X1 U7042 ( .A(n10182), .ZN(n10183) );
  AND2_X1 U7043 ( .A1(n10105), .A2(n10104), .ZN(n10182) );
  INV_X1 U7044 ( .A(n7433), .ZN(n10117) );
  INV_X1 U7045 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8507) );
  INV_X1 U7046 ( .A(n9720), .ZN(n7995) );
  INV_X1 U7047 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10591) );
  INV_X2 U7048 ( .A(n9003), .ZN(P2_U3893) );
  OAI21_X1 U7049 ( .B1(n7335), .B2(n6909), .A(n6908), .ZN(P2_U3488) );
  OAI21_X1 U7050 ( .B1(n7335), .B2(n10255), .A(n7334), .ZN(P2_U3456) );
  OAI21_X1 U7051 ( .B1(n9258), .B2(n10255), .A(n5913), .ZN(P2_U3455) );
  INV_X1 U7052 ( .A(n9623), .ZN(P1_U3973) );
  NAND4_X1 U7053 ( .A1(n5255), .A2(n5613), .A3(n5254), .A4(n5594), .ZN(n5258)
         );
  NOR2_X2 U7054 ( .A1(n5258), .A2(n5257), .ZN(n5828) );
  NOR2_X1 U7055 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5261) );
  NOR2_X1 U7056 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5260) );
  NOR2_X1 U7057 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5259) );
  INV_X1 U7058 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6940) );
  OR2_X1 U7059 ( .A1(n4726), .A2(n6940), .ZN(n5277) );
  NAND2_X2 U7060 ( .A1(n5269), .A2(n5272), .ZN(n5544) );
  NAND2_X1 U7061 ( .A1(n5842), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5276) );
  INV_X1 U7063 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5271) );
  INV_X1 U7064 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10258) );
  INV_X1 U7065 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7380) );
  INV_X1 U7066 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5284) );
  INV_X1 U7067 ( .A(n5288), .ZN(n5287) );
  INV_X1 U7068 ( .A(SI_1_), .ZN(n5286) );
  NAND2_X1 U7069 ( .A1(n5288), .A2(SI_1_), .ZN(n5318) );
  NAND2_X1 U7070 ( .A1(n5317), .A2(n5318), .ZN(n5303) );
  INV_X1 U7071 ( .A(n5303), .ZN(n5291) );
  OR2_X1 U7072 ( .A1(n5347), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5289) );
  OAI21_X1 U7073 ( .B1(n6256), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n5289), .ZN(
        n5290) );
  NOR2_X2 U7074 ( .A1(n5290), .A2(n10413), .ZN(n5316) );
  NAND2_X1 U7075 ( .A1(n5291), .A2(n5316), .ZN(n5305) );
  NAND2_X1 U7076 ( .A1(n5305), .A2(n5318), .ZN(n5296) );
  INV_X1 U7077 ( .A(SI_2_), .ZN(n5292) );
  NAND2_X1 U7078 ( .A1(n5293), .A2(n5292), .ZN(n5319) );
  INV_X1 U7079 ( .A(n5293), .ZN(n5294) );
  NAND2_X1 U7080 ( .A1(n5294), .A2(SI_2_), .ZN(n5321) );
  NAND2_X1 U7081 ( .A1(n5319), .A2(n5321), .ZN(n5295) );
  INV_X1 U7082 ( .A(n4699), .ZN(n7597) );
  NAND2_X1 U7083 ( .A1(n5653), .A2(n7597), .ZN(n5298) );
  NAND2_X1 U7084 ( .A1(n7819), .A2(n5891), .ZN(n5955) );
  INV_X1 U7085 ( .A(n7825), .ZN(n5338) );
  INV_X1 U7086 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5299) );
  INV_X1 U7087 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10331) );
  INV_X1 U7088 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U7089 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5301) );
  INV_X1 U7090 ( .A(n5316), .ZN(n5302) );
  NAND2_X1 U7091 ( .A1(n5303), .A2(n5302), .ZN(n5304) );
  AND2_X1 U7092 ( .A1(n5305), .A2(n5304), .ZN(n6249) );
  INV_X1 U7093 ( .A(n6249), .ZN(n7381) );
  INV_X1 U7094 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5306) );
  INV_X1 U7095 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7416) );
  OR2_X1 U7096 ( .A1(n5544), .A2(n7416), .ZN(n5308) );
  INV_X1 U7097 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6984) );
  OR2_X1 U7098 ( .A1(n4711), .A2(n6984), .ZN(n5307) );
  NAND2_X1 U7099 ( .A1(n7378), .A2(SI_0_), .ZN(n5310) );
  XNOR2_X1 U7100 ( .A(n5310), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9431) );
  MUX2_X1 U7101 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9431), .S(n6913), .Z(n7753) );
  INV_X1 U7102 ( .A(n7753), .ZN(n7745) );
  NAND2_X1 U7103 ( .A1(n7756), .A2(n5184), .ZN(n7823) );
  NAND2_X1 U7104 ( .A1(n7824), .A2(n5245), .ZN(n5337) );
  INV_X1 U7105 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5311) );
  OR2_X1 U7106 ( .A1(n5544), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5313) );
  INV_X1 U7107 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7519) );
  OR2_X1 U7108 ( .A1(n4711), .A2(n7519), .ZN(n5312) );
  INV_X1 U7109 ( .A(n5318), .ZN(n5320) );
  NAND2_X1 U7110 ( .A1(n5320), .A2(n5319), .ZN(n5322) );
  INV_X1 U7111 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U7112 ( .A1(n5326), .A2(SI_3_), .ZN(n5384) );
  NAND2_X1 U7113 ( .A1(n5384), .A2(n5382), .ZN(n5328) );
  NAND2_X1 U7114 ( .A1(n5327), .A2(n5328), .ZN(n5330) );
  INV_X1 U7115 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U7116 ( .A1(n6087), .A2(n7372), .ZN(n5336) );
  NAND2_X1 U7117 ( .A1(n5333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U7118 ( .A1(n5653), .A2(n7524), .ZN(n5335) );
  OR2_X1 U7119 ( .A1(n5358), .A2(n5325), .ZN(n5334) );
  AND3_X2 U7120 ( .A1(n5336), .A2(n5335), .A3(n5334), .ZN(n7887) );
  NAND2_X1 U7121 ( .A1(n9240), .A2(n7887), .ZN(n5965) );
  OAI211_X1 U7122 ( .C1(n5955), .C2(n5338), .A(n5337), .B(n7827), .ZN(n7910)
         );
  INV_X1 U7123 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5339) );
  INV_X1 U7124 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6950) );
  INV_X1 U7125 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U7126 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5341) );
  AND2_X1 U7127 ( .A1(n5362), .A2(n5341), .ZN(n8074) );
  OR2_X1 U7128 ( .A1(n5544), .A2(n8074), .ZN(n5344) );
  INV_X1 U7129 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5342) );
  OR2_X1 U7130 ( .A1(n5404), .A2(n5342), .ZN(n5343) );
  OR2_X1 U7131 ( .A1(n5347), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5348) );
  INV_X1 U7132 ( .A(SI_4_), .ZN(n5349) );
  NAND2_X1 U7133 ( .A1(n5350), .A2(n5349), .ZN(n5388) );
  INV_X1 U7134 ( .A(n5350), .ZN(n5351) );
  NAND2_X1 U7135 ( .A1(n5388), .A2(n5387), .ZN(n5353) );
  NAND2_X1 U7136 ( .A1(n5352), .A2(n5353), .ZN(n5356) );
  INV_X1 U7137 ( .A(n5353), .ZN(n5354) );
  NAND2_X1 U7138 ( .A1(n5356), .A2(n5368), .ZN(n7398) );
  OR2_X1 U7139 ( .A1(n7398), .A2(n5357), .ZN(n5360) );
  NAND2_X1 U7140 ( .A1(n4427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5359) );
  NOR2_X1 U7141 ( .A1(n9240), .A2(n7976), .ZN(n7908) );
  AND2_X1 U7142 ( .A1(n8020), .A2(n5155), .ZN(n7918) );
  AOI21_X1 U7143 ( .B1(n7919), .B2(n7908), .A(n7918), .ZN(n5374) );
  NAND2_X1 U7144 ( .A1(n6088), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U7145 ( .A1(n5714), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5366) );
  INV_X1 U7146 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10260) );
  OR2_X1 U7147 ( .A1(n4711), .A2(n10260), .ZN(n5365) );
  INV_X1 U7148 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U7149 ( .A1(n5362), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5363) );
  AND2_X1 U7150 ( .A1(n5402), .A2(n5363), .ZN(n8025) );
  OR2_X1 U7151 ( .A1(n5544), .A2(n8025), .ZN(n5364) );
  XNOR2_X1 U7152 ( .A(n5385), .B(SI_5_), .ZN(n5376) );
  NAND2_X1 U7153 ( .A1(n7387), .A2(n6087), .ZN(n5373) );
  NAND2_X1 U7154 ( .A1(n5398), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5371) );
  XNOR2_X1 U7155 ( .A(n5371), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6991) );
  AOI22_X1 U7156 ( .A1(n6086), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5653), .B2(
        n6991), .ZN(n5372) );
  OR2_X1 U7157 ( .A1(n8911), .A2(n10238), .ZN(n6115) );
  NAND2_X1 U7158 ( .A1(n10238), .A2(n8911), .ZN(n6114) );
  INV_X1 U7159 ( .A(n5385), .ZN(n5375) );
  INV_X1 U7160 ( .A(SI_5_), .ZN(n10330) );
  OAI21_X1 U7161 ( .B1(n5377), .B2(n5376), .A(n5392), .ZN(n5381) );
  OAI21_X1 U7162 ( .B1(n5380), .B2(SI_6_), .A(n5411), .ZN(n5394) );
  NAND2_X1 U7163 ( .A1(n5381), .A2(n5394), .ZN(n5397) );
  INV_X1 U7164 ( .A(n5384), .ZN(n5389) );
  NAND2_X1 U7165 ( .A1(n5385), .A2(SI_5_), .ZN(n5386) );
  NAND2_X1 U7166 ( .A1(n5391), .A2(n5390), .ZN(n5396) );
  INV_X1 U7167 ( .A(n5392), .ZN(n5393) );
  NOR2_X1 U7168 ( .A1(n5394), .A2(n5393), .ZN(n5395) );
  NAND2_X1 U7169 ( .A1(n5418), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5399) );
  AOI22_X1 U7170 ( .A1(n6086), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5653), .B2(
        n6992), .ZN(n5400) );
  NAND2_X1 U7171 ( .A1(n6088), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U7172 ( .A1(n5843), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U7173 ( .A1(n5402), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5403) );
  AND2_X1 U7174 ( .A1(n5425), .A2(n5403), .ZN(n8124) );
  OR2_X1 U7175 ( .A1(n5544), .A2(n8124), .ZN(n5407) );
  INV_X1 U7176 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5405) );
  OR2_X1 U7177 ( .A1(n6092), .A2(n5405), .ZN(n5406) );
  AND2_X1 U7178 ( .A1(n8121), .A2(n8910), .ZN(n5410) );
  NAND2_X1 U7179 ( .A1(n5412), .A2(SI_7_), .ZN(n5466) );
  OAI21_X1 U7180 ( .B1(n5412), .B2(SI_7_), .A(n5466), .ZN(n5414) );
  NAND2_X1 U7181 ( .A1(n5413), .A2(n5414), .ZN(n5417) );
  NAND2_X1 U7182 ( .A1(n5417), .A2(n5470), .ZN(n7385) );
  OR2_X1 U7183 ( .A1(n7385), .A2(n5357), .ZN(n5422) );
  INV_X1 U7184 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U7185 ( .A1(n5433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5420) );
  XNOR2_X1 U7186 ( .A(n5420), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6955) );
  AOI22_X1 U7187 ( .A1(n6086), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5653), .B2(
        n6955), .ZN(n5421) );
  NAND2_X1 U7188 ( .A1(n5422), .A2(n5421), .ZN(n8259) );
  NAND2_X1 U7189 ( .A1(n6088), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7190 ( .A1(n5714), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5429) );
  INV_X1 U7191 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10262) );
  OR2_X1 U7192 ( .A1(n4711), .A2(n10262), .ZN(n5428) );
  INV_X1 U7193 ( .A(n5425), .ZN(n5424) );
  NAND2_X1 U7194 ( .A1(n5425), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5426) );
  AND2_X1 U7195 ( .A1(n5439), .A2(n5426), .ZN(n8262) );
  OR2_X1 U7196 ( .A1(n5544), .A2(n8262), .ZN(n5427) );
  NAND4_X1 U7197 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n8909)
         );
  NAND2_X1 U7198 ( .A1(n8259), .A2(n8909), .ZN(n5431) );
  NAND2_X1 U7199 ( .A1(n5432), .A2(n5431), .ZN(n8043) );
  XNOR2_X1 U7200 ( .A(n5467), .B(SI_8_), .ZN(n5449) );
  NAND2_X1 U7201 ( .A1(n7406), .A2(n6087), .ZN(n5438) );
  INV_X1 U7202 ( .A(n5433), .ZN(n5435) );
  INV_X1 U7203 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U7204 ( .A1(n5435), .A2(n5434), .ZN(n5453) );
  NAND2_X1 U7205 ( .A1(n5453), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5436) );
  AOI22_X1 U7206 ( .A1(n6086), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5653), .B2(
        n6998), .ZN(n5437) );
  NAND2_X1 U7207 ( .A1(n5843), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5445) );
  INV_X1 U7208 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6997) );
  OR2_X1 U7209 ( .A1(n4726), .A2(n6997), .ZN(n5444) );
  NAND2_X1 U7210 ( .A1(n5439), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5440) );
  AND2_X1 U7211 ( .A1(n5458), .A2(n5440), .ZN(n8402) );
  INV_X1 U7212 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5441) );
  OR2_X1 U7213 ( .A1(n6092), .A2(n5441), .ZN(n5442) );
  AND2_X1 U7214 ( .A1(n10248), .A2(n8908), .ZN(n5446) );
  INV_X1 U7215 ( .A(n5467), .ZN(n5448) );
  INV_X1 U7216 ( .A(SI_8_), .ZN(n5447) );
  NAND2_X1 U7217 ( .A1(n5448), .A2(n5447), .ZN(n5468) );
  XNOR2_X2 U7218 ( .A(n5452), .B(n5469), .ZN(n6366) );
  NAND2_X1 U7219 ( .A1(n6366), .A2(n6087), .ZN(n5456) );
  OAI21_X1 U7220 ( .B1(n5453), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5454) );
  AOI22_X1 U7221 ( .A1(n6086), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7005), .B2(
        n5653), .ZN(n5455) );
  NAND2_X1 U7222 ( .A1(n5456), .A2(n5455), .ZN(n8554) );
  INV_X1 U7223 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10495) );
  OR2_X1 U7224 ( .A1(n4711), .A2(n10495), .ZN(n5463) );
  NAND2_X1 U7225 ( .A1(n5714), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5462) );
  INV_X1 U7226 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10315) );
  OR2_X1 U7227 ( .A1(n4726), .A2(n10315), .ZN(n5461) );
  NAND2_X1 U7228 ( .A1(n5458), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5459) );
  AND2_X1 U7229 ( .A1(n5484), .A2(n5459), .ZN(n8562) );
  OR2_X1 U7230 ( .A1(n5544), .A2(n8562), .ZN(n5460) );
  NOR2_X1 U7231 ( .A1(n8554), .A2(n8742), .ZN(n5465) );
  NAND2_X1 U7232 ( .A1(n8554), .A2(n8742), .ZN(n5464) );
  OAI21_X1 U7233 ( .B1(n8165), .B2(n5465), .A(n5464), .ZN(n8448) );
  INV_X1 U7234 ( .A(SI_9_), .ZN(n5471) );
  NAND2_X1 U7235 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  NAND2_X1 U7236 ( .A1(n5474), .A2(SI_10_), .ZN(n5493) );
  OAI21_X1 U7237 ( .B1(n5474), .B2(SI_10_), .A(n5493), .ZN(n5477) );
  NAND2_X1 U7238 ( .A1(n5494), .A2(n5478), .ZN(n7405) );
  OR2_X1 U7239 ( .A1(n7405), .A2(n5357), .ZN(n5483) );
  INV_X1 U7240 ( .A(n5479), .ZN(n5480) );
  OAI21_X1 U7241 ( .B1(n4427), .B2(n5480), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5481) );
  XNOR2_X1 U7242 ( .A(n5481), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8102) );
  AOI22_X1 U7243 ( .A1(n6086), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5653), .B2(
        n8102), .ZN(n5482) );
  NAND2_X1 U7244 ( .A1(n5843), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5489) );
  INV_X1 U7245 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7007) );
  OR2_X1 U7246 ( .A1(n4726), .A2(n7007), .ZN(n5488) );
  NAND2_X1 U7247 ( .A1(n5484), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5485) );
  AND2_X1 U7248 ( .A1(n5498), .A2(n5485), .ZN(n8453) );
  OR2_X1 U7249 ( .A1(n5544), .A2(n8453), .ZN(n5487) );
  INV_X1 U7250 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8459) );
  OR2_X1 U7251 ( .A1(n6092), .A2(n8459), .ZN(n5486) );
  AND2_X1 U7252 ( .A1(n8669), .A2(n8907), .ZN(n5491) );
  NAND2_X1 U7253 ( .A1(n8745), .A2(n8781), .ZN(n5490) );
  OAI21_X1 U7254 ( .B1(n8448), .B2(n5491), .A(n5490), .ZN(n5492) );
  XNOR2_X1 U7255 ( .A(n5505), .B(SI_11_), .ZN(n5506) );
  XNOR2_X1 U7256 ( .A(n5507), .B(n5506), .ZN(n7454) );
  NAND2_X1 U7257 ( .A1(n7454), .A2(n6087), .ZN(n5497) );
  NAND2_X1 U7258 ( .A1(n5512), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5495) );
  XNOR2_X1 U7259 ( .A(n5495), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8271) );
  AOI22_X1 U7260 ( .A1(n6086), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5653), .B2(
        n8271), .ZN(n5496) );
  NAND2_X1 U7261 ( .A1(n5497), .A2(n5496), .ZN(n8670) );
  NAND2_X1 U7262 ( .A1(n6088), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7263 ( .A1(n5843), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5503) );
  INV_X1 U7264 ( .A(n5517), .ZN(n5518) );
  NAND2_X1 U7265 ( .A1(n5498), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5499) );
  AND2_X1 U7266 ( .A1(n5518), .A2(n5499), .ZN(n8861) );
  OR2_X1 U7267 ( .A1(n5544), .A2(n8861), .ZN(n5502) );
  INV_X1 U7268 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5500) );
  OR2_X1 U7269 ( .A1(n6092), .A2(n5500), .ZN(n5501) );
  NAND4_X1 U7270 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n9224)
         );
  NAND2_X1 U7271 ( .A1(n8670), .A2(n8789), .ZN(n5997) );
  NAND2_X1 U7272 ( .A1(n9198), .A2(n5997), .ZN(n8533) );
  MUX2_X1 U7273 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7370), .Z(n5508) );
  NAND2_X1 U7274 ( .A1(n5508), .A2(SI_12_), .ZN(n5528) );
  OAI21_X1 U7275 ( .B1(n5508), .B2(SI_12_), .A(n5528), .ZN(n5509) );
  NAND2_X1 U7276 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  NAND2_X1 U7277 ( .A1(n5529), .A2(n5511), .ZN(n7481) );
  OR2_X1 U7278 ( .A1(n7481), .A2(n5357), .ZN(n5515) );
  OR2_X2 U7279 ( .A1(n5512), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7280 ( .A1(n5597), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5513) );
  XNOR2_X1 U7281 ( .A(n5513), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8574) );
  AOI22_X1 U7282 ( .A1(n6086), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5653), .B2(
        n8574), .ZN(n5514) );
  NAND2_X1 U7283 ( .A1(n5843), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5523) );
  INV_X1 U7284 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9227) );
  OR2_X1 U7285 ( .A1(n4726), .A2(n9227), .ZN(n5522) );
  NAND2_X1 U7286 ( .A1(n5517), .A2(n5516), .ZN(n5542) );
  NAND2_X1 U7287 ( .A1(n5518), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5519) );
  AND2_X1 U7288 ( .A1(n5542), .A2(n5519), .ZN(n9228) );
  OR2_X1 U7289 ( .A1(n5544), .A2(n9228), .ZN(n5521) );
  INV_X1 U7290 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10386) );
  OR2_X1 U7291 ( .A1(n6092), .A2(n10386), .ZN(n5520) );
  NAND4_X1 U7292 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n9205)
         );
  NOR2_X1 U7293 ( .A1(n9406), .A2(n9205), .ZN(n5527) );
  NAND2_X1 U7294 ( .A1(n8670), .A2(n9224), .ZN(n9220) );
  INV_X1 U7295 ( .A(n9205), .ZN(n8860) );
  NAND2_X1 U7296 ( .A1(n9220), .A2(n8860), .ZN(n5525) );
  INV_X1 U7297 ( .A(n9220), .ZN(n5524) );
  AOI22_X1 U7298 ( .A1(n9406), .A2(n5525), .B1(n5524), .B2(n9205), .ZN(n5526)
         );
  MUX2_X1 U7299 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7370), .Z(n5530) );
  NAND2_X1 U7300 ( .A1(n5530), .A2(SI_13_), .ZN(n5549) );
  INV_X1 U7301 ( .A(n5530), .ZN(n5532) );
  INV_X1 U7302 ( .A(SI_13_), .ZN(n5531) );
  NAND2_X1 U7303 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  OR2_X1 U7304 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  NAND2_X1 U7305 ( .A1(n7644), .A2(n6087), .ZN(n5538) );
  OAI21_X1 U7306 ( .B1(n5597), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5558) );
  XNOR2_X1 U7307 ( .A(n5558), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7017) );
  AOI22_X1 U7308 ( .A1(n6086), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5653), .B2(
        n7017), .ZN(n5537) );
  NAND2_X1 U7309 ( .A1(n5843), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5548) );
  INV_X1 U7310 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5539) );
  OR2_X1 U7311 ( .A1(n4726), .A2(n5539), .ZN(n5547) );
  INV_X1 U7312 ( .A(n5542), .ZN(n5541) );
  NAND2_X1 U7313 ( .A1(n5542), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5543) );
  AND2_X1 U7314 ( .A1(n5565), .A2(n5543), .ZN(n9208) );
  OR2_X1 U7315 ( .A1(n5544), .A2(n9208), .ZN(n5546) );
  INV_X1 U7316 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9399) );
  OR2_X1 U7317 ( .A1(n6092), .A2(n9399), .ZN(n5545) );
  OR2_X1 U7318 ( .A1(n9400), .A2(n9225), .ZN(n6124) );
  NAND2_X1 U7319 ( .A1(n9400), .A2(n9225), .ZN(n6123) );
  MUX2_X1 U7320 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4696), .Z(n5551) );
  NAND2_X1 U7321 ( .A1(n5551), .A2(SI_14_), .ZN(n5574) );
  INV_X1 U7322 ( .A(n5551), .ZN(n5553) );
  INV_X1 U7323 ( .A(SI_14_), .ZN(n5552) );
  NAND2_X1 U7324 ( .A1(n5553), .A2(n5552), .ZN(n5554) );
  NAND2_X1 U7325 ( .A1(n5575), .A2(n5557), .ZN(n7665) );
  NAND2_X1 U7326 ( .A1(n5558), .A2(n5594), .ZN(n5559) );
  NAND2_X1 U7327 ( .A1(n5559), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7328 ( .A1(n5561), .A2(n5560), .ZN(n5577) );
  OR2_X1 U7329 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  AOI22_X1 U7330 ( .A1(n6086), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5653), .B2(
        n8927), .ZN(n5563) );
  INV_X1 U7331 ( .A(n9394), .ZN(n8733) );
  NAND2_X1 U7332 ( .A1(n5565), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7333 ( .A1(n5581), .A2(n5566), .ZN(n9190) );
  NAND2_X1 U7334 ( .A1(n4411), .A2(n9190), .ZN(n5570) );
  NAND2_X1 U7335 ( .A1(n5714), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5569) );
  INV_X1 U7336 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10533) );
  OR2_X1 U7337 ( .A1(n4624), .A2(n10533), .ZN(n5568) );
  OR2_X1 U7338 ( .A1(n4726), .A2(n10566), .ZN(n5567) );
  NAND4_X1 U7339 ( .A1(n5570), .A2(n5569), .A3(n5568), .A4(n5567), .ZN(n9204)
         );
  INV_X1 U7340 ( .A(n9204), .ZN(n8897) );
  NAND2_X1 U7341 ( .A1(n8733), .A2(n8897), .ZN(n5571) );
  NAND2_X1 U7342 ( .A1(n9394), .A2(n9204), .ZN(n5572) );
  MUX2_X1 U7343 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4696), .Z(n5591) );
  XNOR2_X1 U7344 ( .A(n5591), .B(SI_15_), .ZN(n5576) );
  XNOR2_X1 U7345 ( .A(n5590), .B(n5576), .ZN(n7778) );
  NAND2_X1 U7346 ( .A1(n7778), .A2(n6087), .ZN(n5580) );
  NAND2_X1 U7347 ( .A1(n5577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5578) );
  XNOR2_X1 U7348 ( .A(n5578), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7022) );
  AOI22_X1 U7349 ( .A1(n6086), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7022), .B2(
        n5653), .ZN(n5579) );
  NAND2_X1 U7350 ( .A1(n5581), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7351 ( .A1(n5601), .A2(n5582), .ZN(n9184) );
  NAND2_X1 U7352 ( .A1(n9184), .A2(n4411), .ZN(n5585) );
  AOI22_X1 U7353 ( .A1(n5843), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n6088), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7354 ( .A1(n5714), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U7355 ( .A1(n9388), .A2(n8807), .ZN(n9166) );
  NAND2_X1 U7356 ( .A1(n6010), .A2(n9166), .ZN(n9178) );
  NAND2_X1 U7357 ( .A1(n9388), .A2(n9188), .ZN(n5586) );
  INV_X1 U7358 ( .A(n5591), .ZN(n5588) );
  INV_X1 U7359 ( .A(SI_15_), .ZN(n5587) );
  NAND2_X1 U7360 ( .A1(n5588), .A2(n5587), .ZN(n5589) );
  NAND2_X1 U7361 ( .A1(n5591), .A2(SI_15_), .ZN(n5592) );
  MUX2_X1 U7362 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4696), .Z(n5608) );
  XNOR2_X1 U7363 ( .A(n5608), .B(SI_16_), .ZN(n5606) );
  NAND2_X1 U7364 ( .A1(n7804), .A2(n6087), .ZN(n5600) );
  NAND4_X1 U7365 ( .A1(n5593), .A2(n5560), .A3(n5595), .A4(n5594), .ZN(n5596)
         );
  NOR2_X2 U7366 ( .A1(n5597), .A2(n5596), .ZN(n5614) );
  OR2_X1 U7367 ( .A1(n5614), .A2(n5267), .ZN(n5598) );
  XNOR2_X1 U7368 ( .A(n5598), .B(n5613), .ZN(n8968) );
  INV_X1 U7369 ( .A(n8968), .ZN(n6932) );
  AOI22_X1 U7370 ( .A1(n6086), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5653), .B2(
        n6932), .ZN(n5599) );
  NAND2_X1 U7371 ( .A1(n5601), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7372 ( .A1(n5619), .A2(n5602), .ZN(n9174) );
  NAND2_X1 U7373 ( .A1(n9174), .A2(n4411), .ZN(n5605) );
  AOI22_X1 U7374 ( .A1(n5843), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n6088), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7375 ( .A1(n5714), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7376 ( .A1(n9382), .A2(n8815), .ZN(n6011) );
  NAND2_X1 U7377 ( .A1(n6019), .A2(n6011), .ZN(n9170) );
  INV_X1 U7378 ( .A(n5606), .ZN(n5607) );
  MUX2_X1 U7379 ( .A(n7942), .B(n5609), .S(n4696), .Z(n5610) );
  NAND2_X1 U7380 ( .A1(n5610), .A2(n10497), .ZN(n5626) );
  INV_X1 U7381 ( .A(n5610), .ZN(n5611) );
  NAND2_X1 U7382 ( .A1(n5611), .A2(SI_17_), .ZN(n5612) );
  NAND2_X1 U7383 ( .A1(n5626), .A2(n5612), .ZN(n5624) );
  XNOR2_X1 U7384 ( .A(n5625), .B(n5624), .ZN(n7902) );
  NAND2_X1 U7385 ( .A1(n7902), .A2(n6087), .ZN(n5617) );
  NAND2_X1 U7386 ( .A1(n5614), .A2(n5613), .ZN(n5628) );
  NAND2_X1 U7387 ( .A1(n5628), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5615) );
  XNOR2_X1 U7388 ( .A(n5615), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8991) );
  AOI22_X1 U7389 ( .A1(n6086), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5653), .B2(
        n8991), .ZN(n5616) );
  INV_X1 U7390 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U7391 ( .A1(n5619), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U7392 ( .A1(n5631), .A2(n5620), .ZN(n9163) );
  NAND2_X1 U7393 ( .A1(n9163), .A2(n4411), .ZN(n5622) );
  AOI22_X1 U7394 ( .A1(n5714), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n6088), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n5621) );
  OAI211_X1 U7395 ( .C1(n4624), .C2(n9299), .A(n5622), .B(n5621), .ZN(n9171)
         );
  INV_X1 U7396 ( .A(n9171), .ZN(n9144) );
  NAND2_X1 U7397 ( .A1(n9376), .A2(n9144), .ZN(n6012) );
  NAND2_X1 U7398 ( .A1(n6024), .A2(n6012), .ZN(n6127) );
  NAND2_X1 U7399 ( .A1(n9376), .A2(n9171), .ZN(n5623) );
  MUX2_X1 U7400 ( .A(n10441), .B(n8041), .S(n4696), .Z(n5641) );
  XNOR2_X1 U7401 ( .A(n5641), .B(SI_18_), .ZN(n5639) );
  XNOR2_X1 U7402 ( .A(n5640), .B(n5639), .ZN(n8040) );
  NAND2_X1 U7403 ( .A1(n8040), .A2(n6087), .ZN(n5630) );
  XNOR2_X1 U7404 ( .A(n5649), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7026) );
  AOI22_X1 U7405 ( .A1(n6086), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5653), .B2(
        n7026), .ZN(n5629) );
  NAND2_X1 U7406 ( .A1(n5631), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7407 ( .A1(n5656), .A2(n5632), .ZN(n9151) );
  NAND2_X1 U7408 ( .A1(n9151), .A2(n4411), .ZN(n5637) );
  INV_X1 U7409 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U7410 ( .A1(n6088), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7411 ( .A1(n5843), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5633) );
  OAI211_X1 U7412 ( .C1(n9370), .C2(n6092), .A(n5634), .B(n5633), .ZN(n5635)
         );
  INV_X1 U7413 ( .A(n5635), .ZN(n5636) );
  OR2_X1 U7414 ( .A1(n9150), .A2(n9161), .ZN(n5638) );
  INV_X1 U7415 ( .A(n5641), .ZN(n5642) );
  NAND2_X1 U7416 ( .A1(n5642), .A2(SI_18_), .ZN(n5643) );
  MUX2_X1 U7417 ( .A(n8126), .B(n8129), .S(n4696), .Z(n5645) );
  NAND2_X1 U7418 ( .A1(n5645), .A2(n5644), .ZN(n5664) );
  INV_X1 U7419 ( .A(n5645), .ZN(n5646) );
  NAND2_X1 U7420 ( .A1(n5646), .A2(SI_19_), .ZN(n5647) );
  NAND2_X1 U7421 ( .A1(n5664), .A2(n5647), .ZN(n5665) );
  XNOR2_X1 U7422 ( .A(n5666), .B(n5665), .ZN(n8125) );
  NAND2_X1 U7423 ( .A1(n8125), .A2(n6087), .ZN(n5655) );
  NAND2_X1 U7424 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  XNOR2_X2 U7425 ( .A(n5652), .B(n5651), .ZN(n5884) );
  AOI22_X1 U7426 ( .A1(n6086), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6936), .B2(
        n5653), .ZN(n5654) );
  NAND2_X1 U7427 ( .A1(n5656), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7428 ( .A1(n5683), .A2(n5657), .ZN(n9138) );
  NAND2_X1 U7429 ( .A1(n9138), .A2(n4411), .ZN(n5662) );
  INV_X1 U7430 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n10510) );
  NAND2_X1 U7431 ( .A1(n6088), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7432 ( .A1(n5843), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5658) );
  OAI211_X1 U7433 ( .C1(n6092), .C2(n10510), .A(n5659), .B(n5658), .ZN(n5660)
         );
  INV_X1 U7434 ( .A(n5660), .ZN(n5661) );
  NAND2_X1 U7435 ( .A1(n5662), .A2(n5661), .ZN(n8906) );
  NAND2_X1 U7436 ( .A1(n9365), .A2(n9146), .ZN(n6026) );
  MUX2_X1 U7437 ( .A(n8286), .B(n10396), .S(n4696), .Z(n5699) );
  NAND2_X1 U7438 ( .A1(n5680), .A2(n5698), .ZN(n5667) );
  NAND2_X1 U7439 ( .A1(n5668), .A2(n5667), .ZN(n5670) );
  MUX2_X1 U7440 ( .A(n8466), .B(n8426), .S(n4696), .Z(n5696) );
  XNOR2_X1 U7441 ( .A(n5696), .B(SI_21_), .ZN(n5669) );
  NAND2_X1 U7442 ( .A1(n8424), .A2(n6087), .ZN(n5672) );
  OR2_X1 U7443 ( .A1(n5800), .A2(n8466), .ZN(n5671) );
  NAND2_X1 U7444 ( .A1(n5685), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7445 ( .A1(n5712), .A2(n5675), .ZN(n9114) );
  INV_X1 U7446 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9355) );
  NAND2_X1 U7447 ( .A1(n5843), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7448 ( .A1(n6088), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5676) );
  OAI211_X1 U7449 ( .C1(n9355), .C2(n6092), .A(n5677), .B(n5676), .ZN(n5678)
         );
  NAND2_X1 U7450 ( .A1(n9356), .A2(n9121), .ZN(n6028) );
  NAND2_X1 U7451 ( .A1(n6032), .A2(n6028), .ZN(n9110) );
  XNOR2_X1 U7452 ( .A(n5699), .B(SI_20_), .ZN(n5679) );
  NAND2_X1 U7453 ( .A1(n8285), .A2(n6087), .ZN(n5682) );
  OR2_X1 U7454 ( .A1(n5800), .A2(n8286), .ZN(n5681) );
  NAND2_X1 U7455 ( .A1(n5683), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7456 ( .A1(n5685), .A2(n5684), .ZN(n9125) );
  NAND2_X1 U7457 ( .A1(n9125), .A2(n4411), .ZN(n5690) );
  INV_X1 U7458 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U7459 ( .A1(n5843), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7460 ( .A1(n6088), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5686) );
  OAI211_X1 U7461 ( .C1(n9361), .C2(n6092), .A(n5687), .B(n5686), .ZN(n5688)
         );
  INV_X1 U7462 ( .A(n5688), .ZN(n5689) );
  NAND2_X1 U7463 ( .A1(n9124), .A2(n8776), .ZN(n6027) );
  NAND2_X1 U7464 ( .A1(n6031), .A2(n6027), .ZN(n9122) );
  NAND2_X1 U7465 ( .A1(n9365), .A2(n8906), .ZN(n9107) );
  NAND2_X1 U7466 ( .A1(n9106), .A2(n5692), .ZN(n5695) );
  NOR2_X1 U7467 ( .A1(n9124), .A2(n9136), .ZN(n9108) );
  INV_X1 U7468 ( .A(n9356), .ZN(n5693) );
  AOI22_X1 U7469 ( .A1(n9110), .A2(n9108), .B1(n9121), .B2(n5693), .ZN(n5694)
         );
  NAND2_X1 U7470 ( .A1(n5695), .A2(n5694), .ZN(n9096) );
  INV_X1 U7471 ( .A(n5699), .ZN(n5701) );
  INV_X1 U7472 ( .A(n5696), .ZN(n5702) );
  OAI22_X1 U7473 ( .A1(SI_20_), .A2(n5701), .B1(n5702), .B2(SI_21_), .ZN(n5705) );
  INV_X1 U7474 ( .A(SI_21_), .ZN(n5697) );
  OAI21_X1 U7475 ( .B1(n5699), .B2(n5698), .A(n5697), .ZN(n5703) );
  AND2_X1 U7476 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5700) );
  AOI22_X1 U7477 ( .A1(n5703), .A2(n5702), .B1(n5701), .B2(n5700), .ZN(n5704)
         );
  MUX2_X1 U7478 ( .A(n8504), .B(n8507), .S(n4696), .Z(n5707) );
  INV_X1 U7479 ( .A(SI_22_), .ZN(n5706) );
  NAND2_X1 U7480 ( .A1(n5707), .A2(n5706), .ZN(n5721) );
  INV_X1 U7481 ( .A(n5707), .ZN(n5708) );
  NAND2_X1 U7482 ( .A1(n5708), .A2(SI_22_), .ZN(n5709) );
  NAND2_X1 U7483 ( .A1(n5721), .A2(n5709), .ZN(n5722) );
  XNOR2_X1 U7484 ( .A(n5723), .B(n5722), .ZN(n8502) );
  NAND2_X1 U7485 ( .A1(n8502), .A2(n6087), .ZN(n5711) );
  OR2_X1 U7486 ( .A1(n5800), .A2(n8504), .ZN(n5710) );
  NAND2_X1 U7487 ( .A1(n5712), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7488 ( .A1(n5731), .A2(n5713), .ZN(n9102) );
  NAND2_X1 U7489 ( .A1(n9102), .A2(n4411), .ZN(n5719) );
  INV_X1 U7490 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U7491 ( .A1(n5714), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5716) );
  INV_X1 U7492 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9101) );
  OR2_X1 U7493 ( .A1(n4726), .A2(n9101), .ZN(n5715) );
  OAI211_X1 U7494 ( .C1(n4624), .C2(n9281), .A(n5716), .B(n5715), .ZN(n5717)
         );
  INV_X1 U7495 ( .A(n5717), .ZN(n5718) );
  NAND2_X1 U7496 ( .A1(n9350), .A2(n8709), .ZN(n6038) );
  OR2_X1 U7497 ( .A1(n9350), .A2(n9111), .ZN(n5720) );
  INV_X1 U7498 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5724) );
  MUX2_X1 U7499 ( .A(n8512), .B(n5724), .S(n4696), .Z(n5726) );
  INV_X1 U7500 ( .A(SI_23_), .ZN(n5725) );
  NAND2_X1 U7501 ( .A1(n5726), .A2(n5725), .ZN(n5742) );
  INV_X1 U7502 ( .A(n5726), .ZN(n5727) );
  NAND2_X1 U7503 ( .A1(n5727), .A2(SI_23_), .ZN(n5728) );
  NAND2_X1 U7504 ( .A1(n8509), .A2(n6087), .ZN(n5730) );
  OR2_X1 U7505 ( .A1(n5800), .A2(n8512), .ZN(n5729) );
  NAND2_X1 U7506 ( .A1(n5731), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U7507 ( .A1(n4443), .A2(n5732), .ZN(n9091) );
  NAND2_X1 U7508 ( .A1(n9091), .A2(n4411), .ZN(n5738) );
  INV_X1 U7509 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10336) );
  NAND2_X1 U7510 ( .A1(n5843), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5735) );
  INV_X1 U7511 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n10442) );
  OR2_X1 U7512 ( .A1(n4726), .A2(n10442), .ZN(n5734) );
  OAI211_X1 U7513 ( .C1(n10336), .C2(n6092), .A(n5735), .B(n5734), .ZN(n5736)
         );
  INV_X1 U7514 ( .A(n5736), .ZN(n5737) );
  NAND2_X1 U7515 ( .A1(n9344), .A2(n9099), .ZN(n5739) );
  MUX2_X1 U7516 ( .A(n8602), .B(n10359), .S(n4696), .Z(n5744) );
  INV_X1 U7517 ( .A(SI_24_), .ZN(n5743) );
  NAND2_X1 U7518 ( .A1(n5744), .A2(n5743), .ZN(n5759) );
  INV_X1 U7519 ( .A(n5744), .ZN(n5745) );
  NAND2_X1 U7520 ( .A1(n5745), .A2(SI_24_), .ZN(n5746) );
  OR2_X1 U7521 ( .A1(n5800), .A2(n8602), .ZN(n5747) );
  NAND2_X2 U7522 ( .A1(n5748), .A2(n5747), .ZN(n9339) );
  NAND2_X1 U7523 ( .A1(n4443), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7524 ( .A1(n5766), .A2(n5750), .ZN(n9077) );
  NAND2_X1 U7525 ( .A1(n9077), .A2(n4411), .ZN(n5755) );
  INV_X1 U7526 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U7527 ( .A1(n5843), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7528 ( .A1(n6088), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5751) );
  OAI211_X1 U7529 ( .C1(n10511), .C2(n6092), .A(n5752), .B(n5751), .ZN(n5753)
         );
  INV_X1 U7530 ( .A(n5753), .ZN(n5754) );
  AND2_X1 U7531 ( .A1(n9339), .A2(n9089), .ZN(n5756) );
  INV_X1 U7532 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10123) );
  MUX2_X1 U7533 ( .A(n10543), .B(n10123), .S(n4696), .Z(n5761) );
  INV_X1 U7534 ( .A(SI_25_), .ZN(n5760) );
  NAND2_X1 U7535 ( .A1(n5761), .A2(n5760), .ZN(n5776) );
  INV_X1 U7536 ( .A(n5761), .ZN(n5762) );
  NAND2_X1 U7537 ( .A1(n5762), .A2(SI_25_), .ZN(n5763) );
  XNOR2_X1 U7538 ( .A(n5775), .B(n5774), .ZN(n8604) );
  NAND2_X1 U7539 ( .A1(n8604), .A2(n6087), .ZN(n5765) );
  OR2_X1 U7540 ( .A1(n5800), .A2(n10543), .ZN(n5764) );
  NAND2_X1 U7541 ( .A1(n5766), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7542 ( .A1(n4425), .A2(n5767), .ZN(n9066) );
  NAND2_X1 U7543 ( .A1(n9066), .A2(n4411), .ZN(n5772) );
  INV_X1 U7544 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U7545 ( .A1(n6088), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7546 ( .A1(n5843), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5768) );
  OAI211_X1 U7547 ( .C1(n9333), .C2(n6092), .A(n5769), .B(n5768), .ZN(n5770)
         );
  INV_X1 U7548 ( .A(n5770), .ZN(n5771) );
  NAND2_X1 U7549 ( .A1(n9334), .A2(n8829), .ZN(n6049) );
  NAND2_X1 U7550 ( .A1(n6048), .A2(n6049), .ZN(n9060) );
  OR2_X1 U7551 ( .A1(n9334), .A2(n9074), .ZN(n5773) );
  NAND2_X1 U7552 ( .A1(n5775), .A2(n5774), .ZN(n5777) );
  INV_X1 U7553 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9428) );
  INV_X1 U7554 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10119) );
  MUX2_X1 U7555 ( .A(n9428), .B(n10119), .S(n4696), .Z(n5779) );
  NAND2_X1 U7556 ( .A1(n5779), .A2(n5778), .ZN(n5814) );
  INV_X1 U7557 ( .A(n5779), .ZN(n5780) );
  NAND2_X1 U7558 ( .A1(n5780), .A2(SI_26_), .ZN(n5781) );
  NAND2_X1 U7559 ( .A1(n9426), .A2(n6087), .ZN(n5783) );
  OR2_X1 U7560 ( .A1(n5800), .A2(n9428), .ZN(n5782) );
  NAND2_X1 U7561 ( .A1(n4425), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7562 ( .A1(n5805), .A2(n5784), .ZN(n9054) );
  NAND2_X1 U7563 ( .A1(n9054), .A2(n4411), .ZN(n5789) );
  INV_X1 U7564 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10554) );
  NAND2_X1 U7565 ( .A1(n5843), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U7566 ( .A1(n6088), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5785) );
  OAI211_X1 U7567 ( .C1(n10554), .C2(n6092), .A(n5786), .B(n5785), .ZN(n5787)
         );
  INV_X1 U7568 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U7569 ( .A1(n9268), .A2(n9062), .ZN(n5790) );
  NAND2_X1 U7570 ( .A1(n5793), .A2(n5792), .ZN(n5816) );
  NAND2_X1 U7571 ( .A1(n5816), .A2(n5814), .ZN(n5798) );
  INV_X1 U7572 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10429) );
  MUX2_X1 U7573 ( .A(n5799), .B(n10429), .S(n4696), .Z(n5795) );
  INV_X1 U7574 ( .A(SI_27_), .ZN(n5794) );
  NAND2_X1 U7575 ( .A1(n5795), .A2(n5794), .ZN(n5813) );
  INV_X1 U7576 ( .A(n5795), .ZN(n5796) );
  NAND2_X1 U7577 ( .A1(n5796), .A2(SI_27_), .ZN(n5935) );
  AND2_X1 U7578 ( .A1(n5813), .A2(n5935), .ZN(n5797) );
  NAND2_X1 U7579 ( .A1(n9422), .A2(n6087), .ZN(n5802) );
  INV_X1 U7580 ( .A(n5805), .ZN(n5804) );
  INV_X1 U7581 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U7582 ( .A1(n5805), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U7583 ( .A1(n5820), .A2(n5806), .ZN(n9046) );
  NAND2_X1 U7584 ( .A1(n9046), .A2(n4411), .ZN(n5811) );
  INV_X1 U7585 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U7586 ( .A1(n6088), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7587 ( .A1(n5843), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5807) );
  OAI211_X1 U7588 ( .C1(n6092), .C2(n9326), .A(n5808), .B(n5807), .ZN(n5809)
         );
  INV_X1 U7589 ( .A(n5809), .ZN(n5810) );
  AND2_X1 U7590 ( .A1(n9327), .A2(n9050), .ZN(n5812) );
  OR2_X1 U7591 ( .A1(n9327), .A2(n9050), .ZN(n6885) );
  INV_X1 U7592 ( .A(n6885), .ZN(n6887) );
  AND2_X1 U7593 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  INV_X1 U7594 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10113) );
  MUX2_X1 U7595 ( .A(n10410), .B(n10113), .S(n4696), .Z(n5939) );
  XNOR2_X1 U7596 ( .A(n5939), .B(SI_28_), .ZN(n5934) );
  NAND2_X1 U7597 ( .A1(n9419), .A2(n6087), .ZN(n5819) );
  NAND2_X1 U7598 ( .A1(n5820), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7599 ( .A1(n9024), .A2(n5821), .ZN(n8766) );
  NAND2_X1 U7600 ( .A1(n8766), .A2(n4411), .ZN(n5826) );
  INV_X1 U7601 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U7602 ( .A1(n6088), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5823) );
  INV_X1 U7603 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10525) );
  OR2_X1 U7604 ( .A1(n4624), .A2(n10525), .ZN(n5822) );
  OAI211_X1 U7605 ( .C1(n6092), .C2(n10337), .A(n5823), .B(n5822), .ZN(n5824)
         );
  INV_X1 U7606 ( .A(n5824), .ZN(n5825) );
  INV_X1 U7607 ( .A(n5827), .ZN(n5829) );
  OR2_X1 U7608 ( .A1(n5884), .A2(n8503), .ZN(n5841) );
  NAND2_X1 U7609 ( .A1(n5834), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5835) );
  MUX2_X1 U7610 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5835), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5836) );
  INV_X1 U7611 ( .A(n5837), .ZN(n5838) );
  NAND2_X1 U7612 ( .A1(n5838), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7613 ( .A1(n6144), .A2(n7746), .ZN(n5840) );
  INV_X1 U7614 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7332) );
  NAND2_X1 U7615 ( .A1(n6088), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7616 ( .A1(n5843), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5844) );
  OAI211_X1 U7617 ( .C1(n6092), .C2(n7332), .A(n5845), .B(n5844), .ZN(n5846)
         );
  INV_X1 U7618 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U7619 ( .A1(n6096), .A2(n5847), .ZN(n8905) );
  XNOR2_X1 U7620 ( .A(n5869), .B(P2_B_REG_SCAN_IN), .ZN(n5859) );
  XNOR2_X2 U7621 ( .A(n5858), .B(n5857), .ZN(n5864) );
  NAND2_X1 U7622 ( .A1(n5859), .A2(n5864), .ZN(n5868) );
  NAND2_X1 U7623 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  MUX2_X1 U7624 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5861), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5862) );
  INV_X1 U7625 ( .A(n9430), .ZN(n5863) );
  NAND2_X1 U7626 ( .A1(n5864), .A2(n9430), .ZN(n5865) );
  NOR2_X1 U7627 ( .A1(n9430), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7628 ( .A1(n5869), .A2(n9430), .ZN(n7748) );
  INV_X1 U7629 ( .A(n6901), .ZN(n5870) );
  NOR4_X1 U7630 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n10304) );
  NOR2_X1 U7631 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n5873) );
  NOR4_X1 U7632 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n5872) );
  NOR4_X1 U7633 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n5871) );
  NAND4_X1 U7634 ( .A1(n10304), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n5879)
         );
  NOR4_X1 U7635 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5877) );
  NOR4_X1 U7636 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5876) );
  NOR4_X1 U7637 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5875) );
  NOR4_X1 U7638 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5874) );
  NAND4_X1 U7639 ( .A1(n5877), .A2(n5876), .A3(n5875), .A4(n5874), .ZN(n5878)
         );
  NOR2_X1 U7640 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  NAND2_X1 U7641 ( .A1(n5918), .A2(n5916), .ZN(n7710) );
  INV_X1 U7642 ( .A(n7710), .ZN(n5883) );
  AND3_X1 U7643 ( .A1(n6148), .A2(n7746), .A3(n8465), .ZN(n5885) );
  NAND2_X1 U7644 ( .A1(n6936), .A2(n5885), .ZN(n7704) );
  NAND2_X1 U7645 ( .A1(n7737), .A2(n7704), .ZN(n5886) );
  NAND2_X1 U7646 ( .A1(n7703), .A2(n5886), .ZN(n5889) );
  NAND3_X1 U7647 ( .A1(n5921), .A2(n6901), .A3(n5916), .ZN(n7717) );
  NAND2_X1 U7648 ( .A1(n9249), .A2(n10249), .ZN(n9209) );
  AND2_X1 U7649 ( .A1(n6910), .A2(n10241), .ZN(n5887) );
  NAND2_X1 U7650 ( .A1(n7704), .A2(n5887), .ZN(n7701) );
  NAND2_X1 U7651 ( .A1(n9209), .A2(n7701), .ZN(n7709) );
  NAND2_X1 U7652 ( .A1(n7705), .A2(n7709), .ZN(n5888) );
  INV_X1 U7653 ( .A(n7848), .ZN(n5890) );
  NAND2_X1 U7654 ( .A1(n8118), .A2(n10238), .ZN(n8053) );
  INV_X1 U7655 ( .A(n5972), .ZN(n7915) );
  INV_X1 U7656 ( .A(n5973), .ZN(n5894) );
  NOR2_X1 U7657 ( .A1(n8121), .A2(n8256), .ZN(n5964) );
  AOI21_X1 U7658 ( .B1(n5894), .B2(n8054), .A(n5964), .ZN(n5895) );
  INV_X1 U7659 ( .A(n8259), .ZN(n10242) );
  NAND2_X1 U7660 ( .A1(n10242), .A2(n8909), .ZN(n5983) );
  INV_X1 U7661 ( .A(n8909), .ZN(n8396) );
  NAND2_X1 U7662 ( .A1(n8396), .A2(n8259), .ZN(n5988) );
  NAND2_X1 U7663 ( .A1(n8080), .A2(n8083), .ZN(n8082) );
  NAND2_X1 U7664 ( .A1(n10248), .A2(n8556), .ZN(n6119) );
  NAND2_X1 U7665 ( .A1(n8554), .A2(n8397), .ZN(n5989) );
  NAND2_X1 U7666 ( .A1(n5985), .A2(n5989), .ZN(n8164) );
  NAND2_X1 U7667 ( .A1(n8745), .A2(n8907), .ZN(n6118) );
  NAND2_X1 U7668 ( .A1(n8669), .A2(n8781), .ZN(n8531) );
  AND2_X1 U7669 ( .A1(n5997), .A2(n8531), .ZN(n5994) );
  NAND2_X1 U7670 ( .A1(n9406), .A2(n8860), .ZN(n6111) );
  INV_X1 U7671 ( .A(n6111), .ZN(n5899) );
  INV_X1 U7672 ( .A(n9198), .ZN(n9216) );
  NAND2_X1 U7673 ( .A1(n6111), .A2(n9216), .ZN(n5896) );
  OAI211_X1 U7674 ( .C1(n9400), .C2(n8729), .A(n5896), .B(n6112), .ZN(n5897)
         );
  INV_X1 U7675 ( .A(n5897), .ZN(n5898) );
  NAND2_X1 U7676 ( .A1(n9400), .A2(n8729), .ZN(n5900) );
  NAND2_X1 U7677 ( .A1(n8733), .A2(n9204), .ZN(n6005) );
  AND2_X1 U7678 ( .A1(n6011), .A2(n9166), .ZN(n6017) );
  NOR2_X1 U7679 ( .A1(n9150), .A2(n8754), .ZN(n6110) );
  NAND2_X1 U7680 ( .A1(n9150), .A2(n8754), .ZN(n6013) );
  INV_X1 U7681 ( .A(n6031), .ZN(n5903) );
  INV_X1 U7682 ( .A(n6028), .ZN(n6036) );
  NAND2_X1 U7683 ( .A1(n9095), .A2(n6038), .ZN(n5904) );
  NAND2_X1 U7684 ( .A1(n9344), .A2(n8851), .ZN(n9080) );
  INV_X1 U7685 ( .A(n5905), .ZN(n5943) );
  AND2_X1 U7686 ( .A1(n5906), .A2(n6109), .ZN(n6044) );
  NOR2_X1 U7687 ( .A1(n9268), .A2(n8798), .ZN(n6052) );
  NAND2_X1 U7688 ( .A1(n9268), .A2(n8798), .ZN(n5942) );
  OR2_X1 U7689 ( .A1(n9327), .A2(n8884), .ZN(n6058) );
  XNOR2_X1 U7690 ( .A(n6134), .B(n8763), .ZN(n9264) );
  OAI211_X1 U7691 ( .C1(n6148), .C2(n8287), .A(n5884), .B(n10241), .ZN(n5909)
         );
  INV_X1 U7692 ( .A(n5909), .ZN(n5910) );
  INV_X1 U7693 ( .A(n10250), .ZN(n8060) );
  NAND2_X1 U7694 ( .A1(n9261), .A2(n9407), .ZN(n5911) );
  INV_X1 U7695 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7696 ( .A1(n7751), .A2(n6100), .ZN(n5914) );
  NAND2_X1 U7697 ( .A1(n7038), .A2(n5914), .ZN(n7711) );
  INV_X1 U7698 ( .A(n7711), .ZN(n5915) );
  NAND3_X1 U7699 ( .A1(n5916), .A2(n8606), .A3(n5915), .ZN(n5917) );
  NAND3_X1 U7700 ( .A1(n5884), .A2(n6148), .A3(n7746), .ZN(n5919) );
  INV_X1 U7701 ( .A(n6902), .ZN(n5920) );
  NAND2_X1 U7702 ( .A1(n6901), .A2(n5920), .ZN(n5923) );
  NAND2_X1 U7703 ( .A1(n5921), .A2(n6902), .ZN(n5922) );
  OR2_X1 U7704 ( .A1(n9249), .A2(n8465), .ZN(n9252) );
  NAND2_X1 U7705 ( .A1(n9244), .A2(n9252), .ZN(n5926) );
  INV_X1 U7706 ( .A(n5927), .ZN(n5928) );
  INV_X1 U7707 ( .A(n9209), .ZN(n9191) );
  AOI22_X1 U7708 ( .A1(n9261), .A2(n9230), .B1(n9250), .B2(n8766), .ZN(n5929)
         );
  NAND2_X1 U7709 ( .A1(n5932), .A2(n5931), .ZN(P2_U3205) );
  INV_X1 U7710 ( .A(n9261), .ZN(n5933) );
  MUX2_X1 U7711 ( .A(n6879), .B(n5933), .S(n6100), .Z(n6078) );
  MUX2_X1 U7712 ( .A(n6879), .B(n5933), .S(n6910), .Z(n6077) );
  AND2_X1 U7713 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  NAND2_X1 U7714 ( .A1(n5937), .A2(n5936), .ZN(n5941) );
  INV_X1 U7715 ( .A(SI_28_), .ZN(n5938) );
  NAND2_X1 U7716 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  INV_X1 U7717 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9418) );
  INV_X1 U7718 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8662) );
  MUX2_X1 U7719 ( .A(n9418), .B(n8662), .S(n4696), .Z(n6060) );
  INV_X1 U7720 ( .A(n5942), .ZN(n6053) );
  INV_X1 U7721 ( .A(n9052), .ZN(n6051) );
  NAND2_X1 U7722 ( .A1(n6109), .A2(n9079), .ZN(n5944) );
  MUX2_X1 U7723 ( .A(n5944), .B(n5943), .S(n6100), .Z(n6047) );
  AND2_X1 U7724 ( .A1(n6027), .A2(n6026), .ZN(n5947) );
  INV_X1 U7725 ( .A(n6016), .ZN(n5945) );
  NOR2_X1 U7726 ( .A1(n9122), .A2(n5945), .ZN(n5946) );
  MUX2_X1 U7727 ( .A(n5947), .B(n5946), .S(n6910), .Z(n6030) );
  INV_X1 U7728 ( .A(n5951), .ZN(n6113) );
  NAND2_X1 U7729 ( .A1(n6113), .A2(n6144), .ZN(n5948) );
  NAND3_X1 U7730 ( .A1(n5948), .A2(n5950), .A3(n7848), .ZN(n5949) );
  NAND2_X1 U7731 ( .A1(n5949), .A2(n5952), .ZN(n5954) );
  MUX2_X1 U7732 ( .A(n5954), .B(n5953), .S(n6100), .Z(n5959) );
  AND2_X1 U7733 ( .A1(n7819), .A2(n7904), .ZN(n5957) );
  MUX2_X1 U7734 ( .A(n5957), .B(n5956), .S(n6100), .Z(n5958) );
  NAND3_X1 U7735 ( .A1(n5979), .A2(n7911), .A3(n7904), .ZN(n5961) );
  INV_X1 U7736 ( .A(n8054), .ZN(n5966) );
  NAND3_X1 U7737 ( .A1(n5961), .A2(n5960), .A3(n5966), .ZN(n5963) );
  INV_X1 U7738 ( .A(n5964), .ZN(n5968) );
  AND2_X1 U7739 ( .A1(n5965), .A2(n6910), .ZN(n5967) );
  AND4_X1 U7740 ( .A1(n5968), .A2(n7911), .A3(n5967), .A4(n5966), .ZN(n5978)
         );
  NAND2_X1 U7741 ( .A1(n8256), .A2(n6910), .ZN(n5970) );
  NAND2_X1 U7742 ( .A1(n8910), .A2(n6100), .ZN(n5969) );
  OAI22_X1 U7743 ( .A1(n8054), .A2(n5970), .B1(n5969), .B2(n8121), .ZN(n5976)
         );
  NAND2_X1 U7744 ( .A1(n8121), .A2(n6910), .ZN(n5971) );
  AOI21_X1 U7745 ( .B1(n8054), .B2(n8910), .A(n5971), .ZN(n5975) );
  NAND2_X1 U7746 ( .A1(n5972), .A2(n6910), .ZN(n5974) );
  OAI22_X1 U7747 ( .A1(n5976), .A2(n5975), .B1(n5974), .B2(n5973), .ZN(n5977)
         );
  INV_X1 U7748 ( .A(n6121), .ZN(n5980) );
  NAND2_X1 U7749 ( .A1(n5980), .A2(n5985), .ZN(n5991) );
  AND2_X1 U7750 ( .A1(n6119), .A2(n6910), .ZN(n5981) );
  NAND2_X1 U7751 ( .A1(n5989), .A2(n5981), .ZN(n5987) );
  OAI21_X1 U7752 ( .B1(n5991), .B2(n6910), .A(n5987), .ZN(n5982) );
  INV_X1 U7753 ( .A(n5983), .ZN(n5984) );
  NOR2_X1 U7754 ( .A1(n6121), .A2(n5984), .ZN(n5986) );
  OAI211_X1 U7755 ( .C1(n5987), .C2(n5986), .A(n5985), .B(n6118), .ZN(n5993)
         );
  AND2_X1 U7756 ( .A1(n6119), .A2(n5988), .ZN(n5990) );
  OAI211_X1 U7757 ( .C1(n5991), .C2(n5990), .A(n8531), .B(n5989), .ZN(n5992)
         );
  NAND2_X1 U7758 ( .A1(n5996), .A2(n5994), .ZN(n5995) );
  NAND4_X1 U7759 ( .A1(n5995), .A2(n6910), .A3(n9198), .A4(n6112), .ZN(n6002)
         );
  NAND2_X1 U7760 ( .A1(n5996), .A2(n6118), .ZN(n5998) );
  INV_X1 U7761 ( .A(n6112), .ZN(n9199) );
  NAND2_X1 U7762 ( .A1(n9199), .A2(n6100), .ZN(n6001) );
  OAI21_X1 U7763 ( .B1(n9198), .B2(n6910), .A(n6111), .ZN(n5999) );
  OAI21_X1 U7764 ( .B1(n6111), .B2(n6910), .A(n5999), .ZN(n6000) );
  MUX2_X1 U7765 ( .A(n9400), .B(n9225), .S(n6100), .Z(n6003) );
  INV_X1 U7766 ( .A(n6124), .ZN(n6004) );
  MUX2_X1 U7767 ( .A(n6006), .B(n6005), .S(n6100), .Z(n6007) );
  NAND2_X1 U7768 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  INV_X1 U7769 ( .A(n9178), .ZN(n9179) );
  NAND2_X1 U7770 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  NAND2_X1 U7771 ( .A1(n6014), .A2(n6100), .ZN(n6015) );
  INV_X1 U7772 ( .A(n6110), .ZN(n6023) );
  NAND2_X1 U7773 ( .A1(n6018), .A2(n6017), .ZN(n6020) );
  NAND3_X1 U7774 ( .A1(n6020), .A2(n6910), .A3(n6019), .ZN(n6021) );
  NAND2_X1 U7775 ( .A1(n6022), .A2(n6021), .ZN(n6025) );
  NAND2_X1 U7776 ( .A1(n6028), .A2(n6027), .ZN(n6029) );
  INV_X1 U7777 ( .A(n6032), .ZN(n6034) );
  AND2_X1 U7778 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  OAI22_X1 U7779 ( .A1(n6035), .A2(n6034), .B1(n6033), .B2(n6910), .ZN(n6043)
         );
  AOI21_X1 U7780 ( .B1(n6100), .B2(n6036), .A(n9097), .ZN(n6042) );
  INV_X1 U7781 ( .A(n6037), .ZN(n6040) );
  NAND2_X1 U7782 ( .A1(n9080), .A2(n6038), .ZN(n6039) );
  MUX2_X1 U7783 ( .A(n6040), .B(n6039), .S(n6910), .Z(n6041) );
  AOI21_X1 U7784 ( .B1(n6043), .B2(n6042), .A(n6041), .ZN(n6046) );
  MUX2_X1 U7785 ( .A(n6044), .B(n6108), .S(n6910), .Z(n6045) );
  INV_X1 U7786 ( .A(n9060), .ZN(n9068) );
  MUX2_X1 U7787 ( .A(n6049), .B(n6048), .S(n6910), .Z(n6050) );
  MUX2_X1 U7788 ( .A(n6053), .B(n6052), .S(n6100), .Z(n6054) );
  INV_X1 U7789 ( .A(n6054), .ZN(n6055) );
  NAND2_X1 U7790 ( .A1(n9327), .A2(n8884), .ZN(n6057) );
  MUX2_X1 U7791 ( .A(n6058), .B(n6057), .S(n6100), .Z(n6059) );
  OR2_X1 U7792 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  INV_X1 U7793 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10362) );
  INV_X1 U7794 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8612) );
  MUX2_X1 U7795 ( .A(n10362), .B(n8612), .S(n7378), .Z(n6065) );
  INV_X1 U7796 ( .A(SI_30_), .ZN(n6064) );
  NAND2_X1 U7797 ( .A1(n6065), .A2(n6064), .ZN(n6079) );
  INV_X1 U7798 ( .A(n6065), .ZN(n6066) );
  NAND2_X1 U7799 ( .A1(n6066), .A2(SI_30_), .ZN(n6067) );
  NAND2_X1 U7800 ( .A1(n6079), .A2(n6067), .ZN(n6080) );
  OR2_X1 U7801 ( .A1(n5800), .A2(n8612), .ZN(n6068) );
  INV_X1 U7802 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7803 ( .A1(n6088), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6071) );
  INV_X1 U7804 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6069) );
  OR2_X1 U7805 ( .A1(n4624), .A2(n6069), .ZN(n6070) );
  OAI211_X1 U7806 ( .C1(n6072), .C2(n6092), .A(n6071), .B(n6070), .ZN(n6073)
         );
  INV_X1 U7807 ( .A(n6073), .ZN(n6074) );
  NAND2_X1 U7808 ( .A1(n6096), .A2(n6074), .ZN(n8904) );
  INV_X1 U7809 ( .A(n8904), .ZN(n6076) );
  NAND2_X1 U7810 ( .A1(n6097), .A2(n6142), .ZN(n6132) );
  INV_X1 U7811 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6082) );
  MUX2_X1 U7812 ( .A(n4594), .B(n6082), .S(n5347), .Z(n6083) );
  XNOR2_X1 U7813 ( .A(n6083), .B(SI_31_), .ZN(n6084) );
  XNOR2_X1 U7814 ( .A(n6085), .B(n6084), .ZN(n9412) );
  INV_X1 U7815 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7816 ( .A1(n6088), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6091) );
  INV_X1 U7817 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6089) );
  OR2_X1 U7818 ( .A1(n4624), .A2(n6089), .ZN(n6090) );
  OAI211_X1 U7819 ( .C1(n6093), .C2(n6092), .A(n6091), .B(n6090), .ZN(n6094)
         );
  INV_X1 U7820 ( .A(n6094), .ZN(n6095) );
  NAND2_X1 U7821 ( .A1(n6096), .A2(n6095), .ZN(n9023) );
  NOR2_X1 U7822 ( .A1(n9321), .A2(n9023), .ZN(n6133) );
  AOI21_X1 U7823 ( .B1(n6102), .B2(n6910), .A(n6133), .ZN(n6104) );
  INV_X1 U7824 ( .A(n6097), .ZN(n6098) );
  AOI21_X1 U7825 ( .B1(n6100), .B2(n6099), .A(n6098), .ZN(n6101) );
  INV_X1 U7826 ( .A(n9023), .ZN(n6103) );
  NOR2_X1 U7827 ( .A1(n6139), .A2(n6103), .ZN(n6107) );
  XNOR2_X1 U7828 ( .A(n6105), .B(n6936), .ZN(n6106) );
  INV_X1 U7829 ( .A(n6911), .ZN(n7037) );
  NAND2_X1 U7830 ( .A1(n6106), .A2(n5252), .ZN(n6151) );
  INV_X1 U7831 ( .A(n6141), .ZN(n6131) );
  NAND2_X1 U7832 ( .A1(n6109), .A2(n6108), .ZN(n9082) );
  INV_X1 U7833 ( .A(n9097), .ZN(n9094) );
  INV_X1 U7834 ( .A(n9122), .ZN(n9119) );
  NAND2_X1 U7835 ( .A1(n6112), .A2(n6111), .ZN(n9223) );
  NOR3_X1 U7836 ( .A1(n5955), .A2(n7847), .A3(n7827), .ZN(n6117) );
  NAND2_X1 U7837 ( .A1(n6113), .A2(n7848), .ZN(n7736) );
  NOR2_X1 U7838 ( .A1(n7919), .A2(n7736), .ZN(n6116) );
  NAND2_X1 U7839 ( .A1(n6115), .A2(n6114), .ZN(n7921) );
  INV_X1 U7840 ( .A(n6119), .ZN(n6120) );
  OR2_X1 U7841 ( .A1(n6121), .A2(n6120), .ZN(n8047) );
  XNOR2_X1 U7842 ( .A(n8121), .B(n8256), .ZN(n8057) );
  NOR4_X1 U7843 ( .A1(n9223), .A2(n8533), .A3(n8164), .A4(n6122), .ZN(n6125)
         );
  NAND2_X1 U7844 ( .A1(n6124), .A2(n6123), .ZN(n9201) );
  NAND4_X1 U7845 ( .A1(n9179), .A2(n9194), .A3(n6125), .A4(n9201), .ZN(n6126)
         );
  NOR4_X1 U7846 ( .A1(n9148), .A2(n6127), .A3(n9170), .A4(n6126), .ZN(n6128)
         );
  NAND2_X1 U7847 ( .A1(n9079), .A2(n9080), .ZN(n9088) );
  NOR4_X1 U7848 ( .A1(n9037), .A2(n9052), .A3(n9060), .A4(n6129), .ZN(n6130)
         );
  NAND2_X1 U7849 ( .A1(n6134), .A2(n8763), .ZN(n6136) );
  OR2_X1 U7850 ( .A1(n9261), .A2(n6879), .ZN(n6135) );
  OAI21_X1 U7851 ( .B1(n9324), .B2(n6139), .A(n6138), .ZN(n6140) );
  AOI21_X1 U7852 ( .B1(n9023), .B2(n6097), .A(n9321), .ZN(n6143) );
  INV_X1 U7853 ( .A(n7894), .ZN(n8510) );
  NOR2_X1 U7854 ( .A1(n6146), .A2(n7737), .ZN(n7716) );
  NAND3_X1 U7855 ( .A1(n7716), .A2(n7035), .A3(n7033), .ZN(n6147) );
  OAI211_X1 U7856 ( .C1(n6148), .C2(n8510), .A(n6147), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6149) );
  NAND3_X1 U7857 ( .A1(n6151), .A2(n6150), .A3(n6149), .ZN(P2_U3296) );
  NOR2_X1 U7858 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n6155) );
  NAND4_X1 U7859 ( .A1(n6155), .A2(n6199), .A3(n6648), .A4(n6639), .ZN(n6156)
         );
  NAND3_X2 U7860 ( .A1(n6159), .A2(n6158), .A3(n6157), .ZN(n6258) );
  NAND2_X1 U7861 ( .A1(n8660), .A2(n4415), .ZN(n6161) );
  AND2_X4 U7862 ( .A1(n6258), .A2(n7378), .ZN(n6607) );
  NAND2_X1 U7863 ( .A1(n6607), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6160) );
  INV_X1 U7864 ( .A(n6311), .ZN(n6162) );
  NAND2_X1 U7865 ( .A1(n6162), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6337) );
  INV_X1 U7866 ( .A(n6337), .ZN(n6164) );
  NAND2_X1 U7867 ( .A1(n6164), .A2(n6163), .ZN(n6358) );
  INV_X1 U7868 ( .A(n6358), .ZN(n6165) );
  INV_X1 U7869 ( .A(n6400), .ZN(n6166) );
  NAND2_X1 U7870 ( .A1(n6166), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6414) );
  OR2_X2 U7871 ( .A1(n6414), .A2(n6413), .ZN(n6426) );
  INV_X1 U7872 ( .A(n6426), .ZN(n6167) );
  NAND2_X1 U7873 ( .A1(n6167), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6446) );
  OR2_X2 U7874 ( .A1(n6446), .A2(n7782), .ZN(n6468) );
  INV_X1 U7875 ( .A(n6493), .ZN(n6168) );
  OR2_X2 U7876 ( .A1(n6225), .A2(n6213), .ZN(n6237) );
  INV_X1 U7877 ( .A(n6560), .ZN(n6170) );
  INV_X1 U7878 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9499) );
  OR2_X2 U7879 ( .A1(n6571), .A2(n9499), .ZN(n6582) );
  INV_X1 U7880 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9583) );
  INV_X1 U7881 ( .A(n6192), .ZN(n6171) );
  NAND2_X1 U7882 ( .A1(n6171), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U7883 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n6172) );
  NOR2_X1 U7884 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6173) );
  OR2_X1 U7885 ( .A1(n8643), .A2(n6573), .ZN(n6180) );
  INV_X1 U7886 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10381) );
  NAND2_X1 U7887 ( .A1(n6263), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6177) );
  INV_X1 U7888 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8642) );
  OR2_X1 U7889 ( .A1(n6310), .A2(n8642), .ZN(n6176) );
  OAI211_X1 U7890 ( .C1(n6619), .C2(n10381), .A(n6177), .B(n6176), .ZN(n6178)
         );
  INV_X1 U7891 ( .A(n6178), .ZN(n6179) );
  NAND2_X1 U7892 ( .A1(n7352), .A2(n8112), .ZN(n6700) );
  NAND2_X1 U7893 ( .A1(n9419), .A2(n4414), .ZN(n6182) );
  NAND2_X1 U7894 ( .A1(n6607), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6181) );
  NAND2_X2 U7895 ( .A1(n6182), .A2(n6181), .ZN(n8652) );
  INV_X1 U7896 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7315) );
  NAND2_X1 U7897 ( .A1(n6192), .A2(n7315), .ZN(n6183) );
  NAND2_X1 U7898 ( .A1(n8643), .A2(n6183), .ZN(n8650) );
  INV_X1 U7899 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U7900 ( .A1(n6615), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7901 ( .A1(n6263), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6184) );
  OAI211_X1 U7902 ( .C1(n6619), .C2(n7340), .A(n6185), .B(n6184), .ZN(n6186)
         );
  INV_X1 U7903 ( .A(n6186), .ZN(n6187) );
  NAND2_X1 U7904 ( .A1(n9422), .A2(n4415), .ZN(n6190) );
  INV_X1 U7905 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U7906 ( .A1(n6584), .A2(n9436), .ZN(n6191) );
  NAND2_X1 U7907 ( .A1(n6192), .A2(n6191), .ZN(n9818) );
  INV_X1 U7908 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U7909 ( .A1(n6586), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7910 ( .A1(n6263), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6193) );
  OAI211_X1 U7911 ( .C1(n6310), .C2(n9817), .A(n6194), .B(n6193), .ZN(n6195)
         );
  INV_X1 U7912 ( .A(n6195), .ZN(n6196) );
  NAND2_X1 U7913 ( .A1(n9816), .A2(n9587), .ZN(n6844) );
  INV_X1 U7914 ( .A(n6776), .ZN(n6198) );
  NAND2_X1 U7915 ( .A1(n7346), .A2(n6198), .ZN(n6210) );
  NAND2_X1 U7916 ( .A1(n6627), .A2(n6499), .ZN(n6501) );
  INV_X1 U7917 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6205) );
  NAND3_X1 U7918 ( .A1(n6206), .A2(n6205), .A3(n6499), .ZN(n6207) );
  INV_X1 U7919 ( .A(n6834), .ZN(n6614) );
  AOI21_X1 U7920 ( .B1(n6210), .B2(n7347), .A(n6614), .ZN(n6603) );
  NAND2_X1 U7921 ( .A1(n8285), .A2(n4414), .ZN(n6212) );
  OR2_X1 U7922 ( .A1(n6556), .A2(n10396), .ZN(n6211) );
  NAND2_X1 U7923 ( .A1(n6225), .A2(n6213), .ZN(n6214) );
  AND2_X1 U7924 ( .A1(n6237), .A2(n6214), .ZN(n9891) );
  NAND2_X1 U7925 ( .A1(n9891), .A2(n6585), .ZN(n6219) );
  INV_X1 U7926 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10471) );
  NAND2_X1 U7927 ( .A1(n6611), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7928 ( .A1(n6615), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6215) );
  OAI211_X1 U7929 ( .C1(n6619), .C2(n10471), .A(n6216), .B(n6215), .ZN(n6217)
         );
  INV_X1 U7930 ( .A(n6217), .ZN(n6218) );
  NAND2_X1 U7931 ( .A1(n6219), .A2(n6218), .ZN(n9615) );
  INV_X1 U7932 ( .A(n9615), .ZN(n9907) );
  NAND2_X1 U7933 ( .A1(n8125), .A2(n4415), .ZN(n6221) );
  INV_X2 U7934 ( .A(n6258), .ZN(n6502) );
  AOI22_X1 U7935 ( .A1(n9781), .A2(n6502), .B1(n6607), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7936 ( .A1(n9868), .A2(n10092), .ZN(n6222) );
  NAND2_X1 U7937 ( .A1(n6222), .A2(n6834), .ZN(n6231) );
  INV_X1 U7938 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7939 ( .A1(n6507), .A2(n6223), .ZN(n6224) );
  NAND2_X1 U7940 ( .A1(n6225), .A2(n6224), .ZN(n9900) );
  OR2_X1 U7941 ( .A1(n9900), .A2(n6573), .ZN(n6230) );
  INV_X1 U7942 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10341) );
  NAND2_X1 U7943 ( .A1(n6586), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7944 ( .A1(n6611), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6226) );
  OAI211_X1 U7945 ( .C1(n6310), .C2(n10341), .A(n6227), .B(n6226), .ZN(n6228)
         );
  INV_X1 U7946 ( .A(n6228), .ZN(n6229) );
  NAND2_X1 U7947 ( .A1(n6230), .A2(n6229), .ZN(n9616) );
  INV_X1 U7948 ( .A(n9616), .ZN(n9918) );
  OR2_X1 U7949 ( .A1(n9475), .A2(n9918), .ZN(n6745) );
  OR2_X1 U7950 ( .A1(n10028), .A2(n9907), .ZN(n6547) );
  NAND3_X1 U7951 ( .A1(n6231), .A2(n6745), .A3(n6547), .ZN(n6233) );
  NAND3_X1 U7952 ( .A1(n9868), .A2(n6834), .A3(n9616), .ZN(n6232) );
  NAND2_X1 U7953 ( .A1(n6233), .A2(n6232), .ZN(n6543) );
  NAND2_X1 U7954 ( .A1(n8424), .A2(n4415), .ZN(n6235) );
  NAND2_X1 U7955 ( .A1(n6607), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6234) );
  INV_X1 U7956 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7957 ( .A1(n6237), .A2(n6236), .ZN(n6238) );
  NAND2_X1 U7958 ( .A1(n6522), .A2(n6238), .ZN(n9480) );
  OR2_X1 U7959 ( .A1(n9480), .A2(n6573), .ZN(n6243) );
  INV_X1 U7960 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10024) );
  NAND2_X1 U7961 ( .A1(n6615), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7962 ( .A1(n6611), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6239) );
  OAI211_X1 U7963 ( .C1(n10024), .C2(n6619), .A(n6240), .B(n6239), .ZN(n6241)
         );
  INV_X1 U7964 ( .A(n6241), .ZN(n6242) );
  NAND2_X1 U7965 ( .A1(n6243), .A2(n6242), .ZN(n9862) );
  INV_X1 U7966 ( .A(n9862), .ZN(n9886) );
  OR2_X1 U7967 ( .A1(n9876), .A2(n9886), .ZN(n6771) );
  NAND2_X1 U7968 ( .A1(n6263), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6247) );
  INV_X1 U7969 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9625) );
  NAND2_X1 U7970 ( .A1(n6281), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6245) );
  INV_X1 U7971 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U7972 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6248) );
  AOI22_X1 U7973 ( .A1(n6607), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n6502), .B2(
        n9628), .ZN(n6251) );
  NAND2_X1 U7974 ( .A1(n6249), .A2(n6289), .ZN(n6250) );
  NAND2_X1 U7975 ( .A1(n6263), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6255) );
  INV_X1 U7976 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7542) );
  INV_X1 U7977 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7540) );
  OR2_X1 U7978 ( .A1(n6284), .A2(n7540), .ZN(n6252) );
  NAND2_X1 U7979 ( .A1(n7370), .A2(SI_0_), .ZN(n6257) );
  XNOR2_X1 U7980 ( .A(n6257), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10125) );
  OR2_X1 U7981 ( .A1(n6792), .A2(n6260), .ZN(n6261) );
  INV_X1 U7982 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6262) );
  INV_X1 U7983 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8277) );
  INV_X1 U7984 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6264) );
  INV_X1 U7985 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n7420) );
  OR2_X1 U7986 ( .A1(n6284), .A2(n7420), .ZN(n6265) );
  NAND4_X2 U7987 ( .A1(n6268), .A2(n6267), .A3(n6266), .A4(n6265), .ZN(n6273)
         );
  NAND2_X1 U7988 ( .A1(n7374), .A2(n6289), .ZN(n6272) );
  INV_X1 U7989 ( .A(n6269), .ZN(n6270) );
  NAND2_X1 U7990 ( .A1(n6270), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6276) );
  AOI22_X1 U7991 ( .A1(n6607), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n6502), .B2(
        n7582), .ZN(n6271) );
  INV_X1 U7992 ( .A(n7837), .ZN(n7840) );
  OR2_X1 U7993 ( .A1(n6273), .A2(n7842), .ZN(n6274) );
  NAND2_X1 U7994 ( .A1(n7372), .A2(n6289), .ZN(n6280) );
  INV_X1 U7995 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7996 ( .A1(n6276), .A2(n6275), .ZN(n6277) );
  NAND2_X1 U7997 ( .A1(n6277), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6278) );
  XNOR2_X1 U7998 ( .A(n6278), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9639) );
  AOI22_X1 U7999 ( .A1(n6607), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n6502), .B2(
        n9639), .ZN(n6279) );
  NAND2_X1 U8000 ( .A1(n6281), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6288) );
  INV_X1 U8001 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6283) );
  OR2_X1 U8002 ( .A1(n6449), .A2(n6283), .ZN(n6286) );
  INV_X1 U8003 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7424) );
  OR2_X1 U8004 ( .A1(n6284), .A2(n7424), .ZN(n6285) );
  INV_X1 U8005 ( .A(n6761), .ZN(n6319) );
  INV_X1 U8006 ( .A(n6289), .ZN(n6433) );
  OR2_X1 U8007 ( .A1(n7398), .A2(n6433), .ZN(n6293) );
  NAND2_X1 U8008 ( .A1(n6290), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6291) );
  XNOR2_X1 U8009 ( .A(n6291), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7561) );
  AOI22_X1 U8010 ( .A1(n6607), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6502), .B2(
        n7561), .ZN(n6292) );
  NAND2_X1 U8011 ( .A1(n6293), .A2(n6292), .ZN(n10169) );
  INV_X1 U8012 ( .A(n10169), .ZN(n10202) );
  NAND2_X1 U8013 ( .A1(n6611), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6297) );
  INV_X1 U8014 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7441) );
  OR2_X1 U8015 ( .A1(n6310), .A2(n7441), .ZN(n6296) );
  OAI21_X1 U8016 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n6311), .ZN(n10164) );
  OR2_X1 U8017 ( .A1(n6573), .A2(n10164), .ZN(n6295) );
  INV_X1 U8018 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7425) );
  OR2_X1 U8019 ( .A1(n6284), .A2(n7425), .ZN(n6294) );
  NAND2_X1 U8020 ( .A1(n10202), .A2(n9622), .ZN(n6663) );
  NAND2_X1 U8021 ( .A1(n10161), .A2(n10195), .ZN(n6760) );
  AND2_X1 U8022 ( .A1(n8006), .A2(n10169), .ZN(n6659) );
  NAND2_X1 U8023 ( .A1(n6633), .A2(n6299), .ZN(n6369) );
  NAND2_X1 U8024 ( .A1(n6369), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6328) );
  XNOR2_X1 U8025 ( .A(n6328), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7444) );
  AOI22_X1 U8026 ( .A1(n6607), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6502), .B2(
        n7444), .ZN(n6300) );
  NAND2_X1 U8027 ( .A1(n6586), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6305) );
  INV_X1 U8028 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8212) );
  OR2_X1 U8029 ( .A1(n6310), .A2(n8212), .ZN(n6304) );
  INV_X1 U8030 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6336) );
  XNOR2_X1 U8031 ( .A(n6337), .B(n6336), .ZN(n8215) );
  OR2_X1 U8032 ( .A1(n6573), .A2(n8215), .ZN(n6303) );
  INV_X1 U8033 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U8034 ( .A1(n7387), .A2(n4415), .ZN(n6309) );
  NAND2_X1 U8035 ( .A1(n6306), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6307) );
  XNOR2_X1 U8036 ( .A(n6307), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9657) );
  AOI22_X1 U8037 ( .A1(n6607), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6502), .B2(
        n9657), .ZN(n6308) );
  NAND2_X1 U8038 ( .A1(n6586), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6317) );
  INV_X1 U8039 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n8223) );
  OR2_X1 U8040 ( .A1(n6310), .A2(n8223), .ZN(n6316) );
  INV_X1 U8041 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10527) );
  NAND2_X1 U8042 ( .A1(n6311), .A2(n10527), .ZN(n6312) );
  NAND2_X1 U8043 ( .A1(n6337), .A2(n6312), .ZN(n8224) );
  OR2_X1 U8044 ( .A1(n6573), .A2(n8224), .ZN(n6315) );
  INV_X1 U8045 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6313) );
  AND4_X1 U8046 ( .A1(n6763), .A2(n6614), .A3(n6718), .A4(n6663), .ZN(n6318)
         );
  OAI21_X1 U8047 ( .B1(n6323), .B2(n6319), .A(n6318), .ZN(n6353) );
  INV_X1 U8048 ( .A(n6760), .ZN(n6322) );
  NAND2_X1 U8049 ( .A1(n7105), .A2(n6320), .ZN(n6719) );
  AND4_X1 U8050 ( .A1(n8175), .A2(n6834), .A3(n4903), .A4(n6719), .ZN(n6321)
         );
  OAI21_X1 U8051 ( .B1(n6323), .B2(n6322), .A(n6321), .ZN(n6352) );
  NOR2_X1 U8052 ( .A1(n6345), .A2(n8005), .ZN(n6326) );
  AND2_X1 U8053 ( .A1(n6320), .A2(n6614), .ZN(n6347) );
  INV_X1 U8054 ( .A(n6347), .ZN(n6324) );
  OAI21_X1 U8055 ( .B1(n6324), .B2(n9621), .A(n7105), .ZN(n6325) );
  OAI21_X1 U8056 ( .B1(n6326), .B2(n7105), .A(n6325), .ZN(n6344) );
  OR2_X1 U8057 ( .A1(n7385), .A2(n6433), .ZN(n6333) );
  INV_X1 U8058 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U8059 ( .A1(n6328), .A2(n6327), .ZN(n6329) );
  NAND2_X1 U8060 ( .A1(n6329), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6330) );
  INV_X1 U8061 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U8062 ( .A1(n6330), .A2(n10310), .ZN(n6354) );
  OR2_X1 U8063 ( .A1(n6330), .A2(n10310), .ZN(n6331) );
  AOI22_X1 U8064 ( .A1(n6607), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6502), .B2(
        n7613), .ZN(n6332) );
  NAND2_X1 U8065 ( .A1(n6615), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6343) );
  INV_X1 U8066 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6334) );
  OR2_X1 U8067 ( .A1(n6284), .A2(n6334), .ZN(n6342) );
  INV_X1 U8068 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6335) );
  OAI21_X1 U8069 ( .B1(n6337), .B2(n6336), .A(n6335), .ZN(n6338) );
  NAND2_X1 U8070 ( .A1(n6338), .A2(n6358), .ZN(n8243) );
  OR2_X1 U8071 ( .A1(n6573), .A2(n8243), .ZN(n6341) );
  INV_X1 U8072 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6339) );
  OR2_X1 U8073 ( .A1(n4417), .A2(n6339), .ZN(n6340) );
  XNOR2_X1 U8074 ( .A(n8246), .B(n8210), .ZN(n8176) );
  AND2_X1 U8075 ( .A1(n6344), .A2(n8176), .ZN(n6351) );
  OAI22_X1 U8076 ( .A1(n7105), .A2(n6345), .B1(n6614), .B2(n8005), .ZN(n6346)
         );
  INV_X1 U8077 ( .A(n6346), .ZN(n6349) );
  AOI22_X1 U8078 ( .A1(n7105), .A2(n6347), .B1(n6614), .B2(n8005), .ZN(n6348)
         );
  NAND2_X1 U8079 ( .A1(n6354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6355) );
  INV_X1 U8080 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10335) );
  XNOR2_X1 U8081 ( .A(n6355), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7488) );
  AOI22_X1 U8082 ( .A1(n7488), .A2(n6502), .B1(n6607), .B2(
        P2_DATAO_REG_8__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8083 ( .A1(n6586), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6363) );
  INV_X1 U8084 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8378) );
  OR2_X1 U8085 ( .A1(n6310), .A2(n8378), .ZN(n6362) );
  INV_X1 U8086 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U8087 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  NAND2_X1 U8088 ( .A1(n6387), .A2(n6359), .ZN(n8379) );
  OR2_X1 U8089 ( .A1(n6573), .A2(n8379), .ZN(n6361) );
  INV_X1 U8090 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n8337) );
  OR2_X1 U8091 ( .A1(n4417), .A2(n8337), .ZN(n6360) );
  OR2_X1 U8092 ( .A1(n8324), .A2(n8438), .ZN(n8433) );
  INV_X1 U8093 ( .A(n8246), .ZN(n8186) );
  NAND2_X1 U8094 ( .A1(n8186), .A2(n8210), .ZN(n6364) );
  AND2_X1 U8095 ( .A1(n8433), .A2(n6364), .ZN(n6654) );
  NAND2_X1 U8096 ( .A1(n8246), .A2(n8332), .ZN(n8328) );
  MUX2_X1 U8097 ( .A(n6654), .B(n6655), .S(n6834), .Z(n6365) );
  NAND2_X1 U8098 ( .A1(n6366), .A2(n4415), .ZN(n6372) );
  NAND2_X1 U8099 ( .A1(n6367), .A2(n10335), .ZN(n6368) );
  NAND2_X1 U8100 ( .A1(n6382), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6370) );
  XNOR2_X1 U8101 ( .A(n6370), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7491) );
  AOI22_X1 U8102 ( .A1(n6607), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6502), .B2(
        n7491), .ZN(n6371) );
  NAND2_X2 U8103 ( .A1(n6372), .A2(n6371), .ZN(n8471) );
  NAND2_X1 U8104 ( .A1(n6586), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6376) );
  INV_X1 U8105 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8469) );
  OR2_X1 U8106 ( .A1(n6310), .A2(n8469), .ZN(n6375) );
  INV_X1 U8107 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7602) );
  XNOR2_X1 U8108 ( .A(n6387), .B(n7602), .ZN(n8468) );
  OR2_X1 U8109 ( .A1(n6573), .A2(n8468), .ZN(n6374) );
  INV_X1 U8110 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10551) );
  OR2_X1 U8111 ( .A1(n4417), .A2(n10551), .ZN(n6373) );
  NAND2_X1 U8112 ( .A1(n8471), .A2(n8333), .ZN(n6806) );
  NAND2_X1 U8113 ( .A1(n6806), .A2(n8432), .ZN(n6379) );
  MUX2_X1 U8114 ( .A(n6379), .B(n6656), .S(n6834), .Z(n6380) );
  INV_X1 U8115 ( .A(n6380), .ZN(n6381) );
  OR2_X1 U8116 ( .A1(n7405), .A2(n6433), .ZN(n6386) );
  INV_X1 U8117 ( .A(n6382), .ZN(n6384) );
  NAND2_X1 U8118 ( .A1(n6384), .A2(n6383), .ZN(n6439) );
  NAND2_X1 U8119 ( .A1(n6439), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6408) );
  XNOR2_X1 U8120 ( .A(n6408), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9690) );
  AOI22_X1 U8121 ( .A1(n6502), .A2(n9690), .B1(n6607), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n6385) );
  INV_X1 U8122 ( .A(n8308), .ZN(n8317) );
  NAND2_X1 U8123 ( .A1(n6586), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6392) );
  INV_X1 U8124 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7493) );
  OR2_X1 U8125 ( .A1(n6310), .A2(n7493), .ZN(n6391) );
  INV_X1 U8126 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10430) );
  OAI21_X1 U8127 ( .B1(n6387), .B2(n7602), .A(n10430), .ZN(n6388) );
  NAND2_X1 U8128 ( .A1(n6388), .A2(n6400), .ZN(n8313) );
  OR2_X1 U8129 ( .A1(n6573), .A2(n8313), .ZN(n6390) );
  INV_X1 U8130 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8300) );
  OR2_X1 U8131 ( .A1(n4417), .A2(n8300), .ZN(n6389) );
  NAND4_X1 U8132 ( .A1(n6392), .A2(n6391), .A3(n6390), .A4(n6389), .ZN(n9619)
         );
  NAND2_X1 U8133 ( .A1(n8317), .A2(n8486), .ZN(n6726) );
  NAND2_X1 U8134 ( .A1(n6393), .A2(n6726), .ZN(n6406) );
  NAND2_X1 U8135 ( .A1(n7454), .A2(n4414), .ZN(n6398) );
  NAND2_X1 U8136 ( .A1(n6408), .A2(n6436), .ZN(n6395) );
  NAND2_X1 U8137 ( .A1(n6395), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6396) );
  XNOR2_X1 U8138 ( .A(n6396), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7674) );
  AOI22_X1 U8139 ( .A1(n7674), .A2(n6502), .B1(n6607), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U8140 ( .A1(n6615), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6405) );
  INV_X1 U8141 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10468) );
  OR2_X1 U8142 ( .A1(n6619), .A2(n10468), .ZN(n6404) );
  INV_X1 U8143 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8144 ( .A1(n6400), .A2(n6399), .ZN(n6401) );
  NAND2_X1 U8145 ( .A1(n6414), .A2(n6401), .ZN(n8487) );
  OR2_X1 U8146 ( .A1(n6573), .A2(n8487), .ZN(n6403) );
  INV_X1 U8147 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10469) );
  OR2_X1 U8148 ( .A1(n4417), .A2(n10469), .ZN(n6402) );
  OR2_X1 U8149 ( .A1(n8490), .A2(n7159), .ZN(n6728) );
  NAND2_X1 U8150 ( .A1(n8308), .A2(n9619), .ZN(n6725) );
  NAND3_X1 U8151 ( .A1(n6406), .A2(n6728), .A3(n6725), .ZN(n6421) );
  OR2_X1 U8152 ( .A1(n7481), .A2(n6433), .ZN(n6412) );
  OAI21_X1 U8153 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8154 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  NAND2_X1 U8155 ( .A1(n6409), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6410) );
  AOI22_X1 U8156 ( .A1(n7784), .A2(n6502), .B1(n6607), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U8157 ( .A1(n6611), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6420) );
  INV_X1 U8158 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8349) );
  OR2_X1 U8159 ( .A1(n6310), .A2(n8349), .ZN(n6419) );
  NAND2_X1 U8160 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  NAND2_X1 U8161 ( .A1(n6426), .A2(n6415), .ZN(n9492) );
  OR2_X1 U8162 ( .A1(n6573), .A2(n9492), .ZN(n6418) );
  INV_X1 U8163 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6416) );
  OR2_X1 U8164 ( .A1(n6619), .A2(n6416), .ZN(n6417) );
  NAND4_X1 U8165 ( .A1(n6420), .A2(n6419), .A3(n6418), .A4(n6417), .ZN(n9618)
         );
  NAND2_X1 U8166 ( .A1(n9494), .A2(n8591), .ZN(n6729) );
  NAND2_X1 U8167 ( .A1(n8490), .A2(n7159), .ZN(n6727) );
  NAND2_X1 U8168 ( .A1(n8348), .A2(n9618), .ZN(n6730) );
  NAND2_X1 U8169 ( .A1(n7644), .A2(n4414), .ZN(n6425) );
  NAND2_X1 U8170 ( .A1(n6422), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6423) );
  XNOR2_X1 U8171 ( .A(n6423), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9707) );
  AOI22_X1 U8172 ( .A1(n9707), .A2(n6502), .B1(n6607), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8173 ( .A1(n6615), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6431) );
  INV_X1 U8174 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10340) );
  OR2_X1 U8175 ( .A1(n4417), .A2(n10340), .ZN(n6430) );
  INV_X1 U8176 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9701) );
  NAND2_X1 U8177 ( .A1(n6426), .A2(n9701), .ZN(n6427) );
  NAND2_X1 U8178 ( .A1(n6446), .A2(n6427), .ZN(n9553) );
  OR2_X1 U8179 ( .A1(n6573), .A2(n9553), .ZN(n6429) );
  INV_X1 U8180 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10064) );
  OR2_X1 U8181 ( .A1(n6619), .A2(n10064), .ZN(n6428) );
  NAND2_X1 U8182 ( .A1(n9555), .A2(n9444), .ZN(n8521) );
  INV_X1 U8183 ( .A(n8521), .ZN(n6733) );
  OR2_X1 U8184 ( .A1(n9555), .A2(n9444), .ZN(n6731) );
  INV_X1 U8185 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6435) );
  NAND4_X1 U8186 ( .A1(n6437), .A2(n6436), .A3(n6435), .A4(n6434), .ZN(n6438)
         );
  NAND2_X1 U8187 ( .A1(n6441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6440) );
  MUX2_X1 U8188 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6440), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6442) );
  NAND2_X1 U8189 ( .A1(n6442), .A2(n6464), .ZN(n7991) );
  INV_X1 U8190 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7664) );
  OAI22_X1 U8191 ( .A1(n7991), .A2(n7393), .B1(n6556), .B2(n7664), .ZN(n6443)
         );
  INV_X1 U8192 ( .A(n6443), .ZN(n6444) );
  INV_X1 U8193 ( .A(n10058), .ZN(n8516) );
  NAND2_X1 U8194 ( .A1(n6615), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6453) );
  INV_X1 U8195 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10361) );
  OR2_X1 U8196 ( .A1(n6619), .A2(n10361), .ZN(n6452) );
  NAND2_X1 U8197 ( .A1(n6446), .A2(n7782), .ZN(n6447) );
  NAND2_X1 U8198 ( .A1(n6468), .A2(n6447), .ZN(n9448) );
  OR2_X1 U8199 ( .A1(n6573), .A2(n9448), .ZN(n6451) );
  INV_X1 U8200 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n6448) );
  OR2_X1 U8201 ( .A1(n4417), .A2(n6448), .ZN(n6450) );
  NAND4_X1 U8202 ( .A1(n6453), .A2(n6452), .A3(n6451), .A4(n6450), .ZN(n9979)
         );
  INV_X1 U8203 ( .A(n9979), .ZN(n8590) );
  NAND2_X1 U8204 ( .A1(n10058), .A2(n8590), .ZN(n6484) );
  NAND2_X1 U8205 ( .A1(n6735), .A2(n6484), .ZN(n6757) );
  NAND2_X1 U8206 ( .A1(n7804), .A2(n4414), .ZN(n6458) );
  INV_X1 U8207 ( .A(n6454), .ZN(n6455) );
  NAND2_X1 U8208 ( .A1(n6455), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6456) );
  XNOR2_X1 U8209 ( .A(n6456), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9731) );
  AOI22_X1 U8210 ( .A1(n6607), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6502), .B2(
        n9731), .ZN(n6457) );
  INV_X1 U8211 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U8212 ( .A1(n6470), .A2(n6459), .ZN(n6460) );
  NAND2_X1 U8213 ( .A1(n6493), .A2(n6460), .ZN(n9963) );
  OR2_X1 U8214 ( .A1(n9963), .A2(n6573), .ZN(n6463) );
  AOI22_X1 U8215 ( .A1(n6586), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6615), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8216 ( .A1(n6611), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U8217 ( .A1(n9961), .A2(n9524), .ZN(n6737) );
  NAND2_X1 U8218 ( .A1(n7778), .A2(n4415), .ZN(n6467) );
  NAND2_X1 U8219 ( .A1(n6464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6465) );
  XNOR2_X1 U8220 ( .A(n6465), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9720) );
  AOI22_X1 U8221 ( .A1(n9720), .A2(n6502), .B1(n6607), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8222 ( .A1(n6468), .A2(n9602), .ZN(n6469) );
  NAND2_X1 U8223 ( .A1(n6470), .A2(n6469), .ZN(n9973) );
  INV_X1 U8224 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10411) );
  OAI22_X1 U8225 ( .A1(n9973), .A2(n6573), .B1(n4417), .B2(n10411), .ZN(n6474)
         );
  INV_X1 U8226 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U8227 ( .A1(n6586), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6471) );
  OAI21_X1 U8228 ( .B1(n6310), .B2(n6472), .A(n6471), .ZN(n6473) );
  INV_X1 U8229 ( .A(n9952), .ZN(n9515) );
  NAND2_X1 U8230 ( .A1(n10052), .A2(n9515), .ZN(n9947) );
  AND2_X1 U8231 ( .A1(n9947), .A2(n6484), .ZN(n6673) );
  AND2_X1 U8232 ( .A1(n6737), .A2(n6673), .ZN(n6476) );
  INV_X1 U8233 ( .A(n6740), .ZN(n6475) );
  OR2_X1 U8234 ( .A1(n10052), .A2(n9515), .ZN(n6736) );
  AND2_X1 U8235 ( .A1(n6740), .A2(n6736), .ZN(n6676) );
  NAND2_X1 U8236 ( .A1(n6730), .A2(n6728), .ZN(n6479) );
  INV_X1 U8237 ( .A(n6725), .ZN(n6477) );
  NOR2_X1 U8238 ( .A1(n6479), .A2(n6477), .ZN(n6668) );
  NAND2_X1 U8239 ( .A1(n6478), .A2(n6668), .ZN(n6483) );
  INV_X1 U8240 ( .A(n6479), .ZN(n6482) );
  NAND2_X1 U8241 ( .A1(n6727), .A2(n6726), .ZN(n6481) );
  INV_X1 U8242 ( .A(n6729), .ZN(n6480) );
  AOI21_X1 U8243 ( .B1(n6482), .B2(n6481), .A(n6480), .ZN(n6669) );
  NAND2_X1 U8244 ( .A1(n6484), .A2(n8521), .ZN(n6485) );
  INV_X1 U8245 ( .A(n9947), .ZN(n6738) );
  NAND3_X1 U8246 ( .A1(n6740), .A2(n6738), .A3(n6834), .ZN(n6488) );
  OR3_X1 U8247 ( .A1(n10052), .A2(n9515), .A3(n6834), .ZN(n6486) );
  MUX2_X1 U8248 ( .A(n6614), .B(n6486), .S(n6737), .Z(n6487) );
  NAND3_X1 U8249 ( .A1(n6489), .A2(n6488), .A3(n6487), .ZN(n6498) );
  NAND2_X1 U8250 ( .A1(n7902), .A2(n4415), .ZN(n6492) );
  NAND2_X1 U8251 ( .A1(n4516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6490) );
  XNOR2_X1 U8252 ( .A(n6490), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9749) );
  AOI22_X1 U8253 ( .A1(n6607), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6502), .B2(
        n9749), .ZN(n6491) );
  INV_X1 U8254 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n6497) );
  INV_X1 U8255 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10498) );
  NAND2_X1 U8256 ( .A1(n6493), .A2(n10498), .ZN(n6494) );
  NAND2_X1 U8257 ( .A1(n6505), .A2(n6494), .ZN(n9933) );
  OR2_X1 U8258 ( .A1(n9933), .A2(n6573), .ZN(n6496) );
  AOI22_X1 U8259 ( .A1(n6586), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n6615), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n6495) );
  OAI211_X1 U8260 ( .C1(n4417), .C2(n6497), .A(n6496), .B(n6495), .ZN(n9953)
         );
  INV_X1 U8261 ( .A(n9953), .ZN(n9920) );
  OR2_X1 U8262 ( .A1(n10043), .A2(n9920), .ZN(n6741) );
  NAND2_X1 U8263 ( .A1(n10043), .A2(n9920), .ZN(n6544) );
  NAND2_X1 U8264 ( .A1(n6498), .A2(n9938), .ZN(n6546) );
  NAND2_X1 U8265 ( .A1(n8040), .A2(n4414), .ZN(n6504) );
  OR2_X1 U8266 ( .A1(n6627), .A2(n6499), .ZN(n6500) );
  AND2_X1 U8267 ( .A1(n6501), .A2(n6500), .ZN(n9769) );
  AOI22_X1 U8268 ( .A1(n6502), .A2(n9769), .B1(n6607), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U8269 ( .A1(n6505), .A2(n9572), .ZN(n6506) );
  AND2_X1 U8270 ( .A1(n6507), .A2(n6506), .ZN(n9923) );
  NAND2_X1 U8271 ( .A1(n9923), .A2(n6585), .ZN(n6513) );
  INV_X1 U8272 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U8273 ( .A1(n6611), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8274 ( .A1(n6615), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6508) );
  OAI211_X1 U8275 ( .C1(n6619), .C2(n6510), .A(n6509), .B(n6508), .ZN(n6511)
         );
  INV_X1 U8276 ( .A(n6511), .ZN(n6512) );
  NAND2_X1 U8277 ( .A1(n6513), .A2(n6512), .ZN(n9940) );
  INV_X1 U8278 ( .A(n9940), .ZN(n9906) );
  OR2_X1 U8279 ( .A1(n10038), .A2(n9906), .ZN(n6742) );
  NAND2_X1 U8280 ( .A1(n6742), .A2(n6741), .ZN(n6679) );
  INV_X1 U8281 ( .A(n6679), .ZN(n6514) );
  NAND2_X1 U8282 ( .A1(n6546), .A2(n6514), .ZN(n6515) );
  NAND2_X1 U8283 ( .A1(n9475), .A2(n9918), .ZN(n6746) );
  NAND2_X1 U8284 ( .A1(n10038), .A2(n9906), .ZN(n6744) );
  NAND3_X1 U8285 ( .A1(n6515), .A2(n6746), .A3(n6744), .ZN(n6516) );
  NAND3_X1 U8286 ( .A1(n6543), .A2(n6771), .A3(n6516), .ZN(n6518) );
  NAND2_X1 U8287 ( .A1(n9876), .A2(n9886), .ZN(n6836) );
  NAND2_X1 U8288 ( .A1(n6836), .A2(n9868), .ZN(n6517) );
  NAND2_X1 U8289 ( .A1(n6517), .A2(n6771), .ZN(n6690) );
  AOI21_X1 U8290 ( .B1(n6518), .B2(n6690), .A(n6834), .ZN(n6542) );
  NAND2_X1 U8291 ( .A1(n8502), .A2(n4414), .ZN(n6520) );
  NAND2_X1 U8292 ( .A1(n6607), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6519) );
  INV_X1 U8293 ( .A(n10017), .ZN(n9857) );
  NAND2_X1 U8294 ( .A1(n6522), .A2(n6521), .ZN(n6523) );
  AND2_X1 U8295 ( .A1(n6531), .A2(n6523), .ZN(n9855) );
  NAND2_X1 U8296 ( .A1(n9855), .A2(n6585), .ZN(n6528) );
  INV_X1 U8297 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10544) );
  NAND2_X1 U8298 ( .A1(n6586), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U8299 ( .A1(n6615), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6524) );
  OAI211_X1 U8300 ( .C1(n10544), .C2(n4417), .A(n6525), .B(n6524), .ZN(n6526)
         );
  INV_X1 U8301 ( .A(n6526), .ZN(n6527) );
  NAND2_X1 U8302 ( .A1(n9857), .A2(n9845), .ZN(n6539) );
  INV_X1 U8303 ( .A(n9845), .ZN(n9875) );
  NAND2_X1 U8304 ( .A1(n10017), .A2(n9875), .ZN(n6837) );
  INV_X1 U8305 ( .A(n9860), .ZN(n6541) );
  NAND2_X1 U8306 ( .A1(n8509), .A2(n4415), .ZN(n6530) );
  NAND2_X1 U8307 ( .A1(n6607), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6529) );
  INV_X1 U8308 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U8309 ( .A1(n6531), .A2(n10565), .ZN(n6532) );
  NAND2_X1 U8310 ( .A1(n6560), .A2(n6532), .ZN(n9460) );
  INV_X1 U8311 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U8312 ( .A1(n6611), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U8313 ( .A1(n6615), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6533) );
  OAI211_X1 U8314 ( .C1(n6619), .C2(n6535), .A(n6534), .B(n6533), .ZN(n6536)
         );
  INV_X1 U8315 ( .A(n6536), .ZN(n6537) );
  INV_X1 U8316 ( .A(n9861), .ZN(n9533) );
  OR2_X1 U8317 ( .A1(n10011), .A2(n9533), .ZN(n6756) );
  NAND2_X1 U8318 ( .A1(n6756), .A2(n6539), .ZN(n6683) );
  NAND2_X1 U8319 ( .A1(n6683), .A2(n6614), .ZN(n6540) );
  NAND2_X1 U8320 ( .A1(n10011), .A2(n9533), .ZN(n8632) );
  INV_X1 U8321 ( .A(n6543), .ZN(n6549) );
  AND2_X1 U8322 ( .A1(n6744), .A2(n6544), .ZN(n6677) );
  AND2_X1 U8323 ( .A1(n6745), .A2(n6742), .ZN(n6681) );
  INV_X1 U8324 ( .A(n6681), .ZN(n6545) );
  AOI21_X1 U8325 ( .B1(n6677), .B2(n6546), .A(n6545), .ZN(n6548) );
  AND2_X1 U8326 ( .A1(n6771), .A2(n6547), .ZN(n6688) );
  OAI21_X1 U8327 ( .B1(n6549), .B2(n6548), .A(n6688), .ZN(n6550) );
  NAND3_X1 U8328 ( .A1(n6550), .A2(n6834), .A3(n6836), .ZN(n6551) );
  NAND3_X1 U8329 ( .A1(n6552), .A2(n8632), .A3(n6551), .ZN(n6555) );
  AND2_X1 U8330 ( .A1(n8632), .A2(n6837), .ZN(n6691) );
  INV_X1 U8331 ( .A(n6691), .ZN(n6553) );
  NAND2_X1 U8332 ( .A1(n6553), .A2(n6834), .ZN(n6554) );
  NAND2_X1 U8333 ( .A1(n8600), .A2(n4414), .ZN(n6558) );
  OR2_X1 U8334 ( .A1(n6556), .A2(n10359), .ZN(n6557) );
  INV_X1 U8335 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U8336 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  NAND2_X1 U8337 ( .A1(n6571), .A2(n6561), .ZN(n9531) );
  INV_X1 U8338 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U8339 ( .A1(n6586), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U8340 ( .A1(n6611), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6562) );
  OAI211_X1 U8341 ( .C1(n6310), .C2(n8629), .A(n6563), .B(n6562), .ZN(n6564)
         );
  INV_X1 U8342 ( .A(n6564), .ZN(n6565) );
  NAND2_X1 U8343 ( .A1(n10008), .A2(n9827), .ZN(n6692) );
  NOR2_X1 U8344 ( .A1(n6756), .A2(n6614), .ZN(n6567) );
  MUX2_X1 U8345 ( .A(n6840), .B(n6692), .S(n6834), .Z(n6568) );
  NAND2_X1 U8346 ( .A1(n8604), .A2(n4415), .ZN(n6570) );
  NAND2_X1 U8347 ( .A1(n6607), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6569) );
  NAND2_X1 U8348 ( .A1(n6571), .A2(n9499), .ZN(n6572) );
  NAND2_X1 U8349 ( .A1(n6582), .A2(n6572), .ZN(n9831) );
  INV_X1 U8350 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U8351 ( .A1(n6611), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6575) );
  NAND2_X1 U8352 ( .A1(n6615), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6574) );
  OAI211_X1 U8353 ( .C1(n6619), .C2(n6576), .A(n6575), .B(n6574), .ZN(n6577)
         );
  INV_X1 U8354 ( .A(n6577), .ZN(n6578) );
  NAND2_X2 U8355 ( .A1(n6579), .A2(n6578), .ZN(n9614) );
  NAND2_X1 U8356 ( .A1(n9426), .A2(n4414), .ZN(n6581) );
  NAND2_X1 U8357 ( .A1(n6607), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U8358 ( .A1(n6582), .A2(n9583), .ZN(n6583) );
  NAND2_X1 U8359 ( .A1(n9591), .A2(n6585), .ZN(n6591) );
  INV_X1 U8360 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10451) );
  NAND2_X1 U8361 ( .A1(n6615), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U8362 ( .A1(n6586), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6587) );
  OAI211_X1 U8363 ( .C1(n4417), .C2(n10451), .A(n6588), .B(n6587), .ZN(n6589)
         );
  INV_X1 U8364 ( .A(n6589), .ZN(n6590) );
  AND2_X2 U8365 ( .A1(n6591), .A2(n6590), .ZN(n9828) );
  NAND2_X1 U8366 ( .A1(n9998), .A2(n9828), .ZN(n6843) );
  NAND2_X1 U8367 ( .A1(n10004), .A2(n9585), .ZN(n6842) );
  NAND2_X1 U8368 ( .A1(n6843), .A2(n6842), .ZN(n6696) );
  AOI21_X1 U8369 ( .B1(n6592), .B2(n6775), .A(n6696), .ZN(n6601) );
  OR2_X2 U8370 ( .A1(n9998), .A2(n9828), .ZN(n6774) );
  NAND4_X1 U8371 ( .A1(n7347), .A2(n6614), .A3(n6776), .A4(n6774), .ZN(n6600)
         );
  NAND2_X1 U8372 ( .A1(n6774), .A2(n6775), .ZN(n6593) );
  NAND2_X1 U8373 ( .A1(n6593), .A2(n6843), .ZN(n6594) );
  OAI21_X1 U8374 ( .B1(n6595), .B2(n6696), .A(n6594), .ZN(n6596) );
  INV_X1 U8375 ( .A(n7347), .ZN(n6597) );
  OAI211_X1 U8376 ( .C1(n6601), .C2(n6600), .A(n6599), .B(n6598), .ZN(n6602)
         );
  MUX2_X1 U8377 ( .A(n6700), .B(n6682), .S(n6834), .Z(n6604) );
  NAND2_X1 U8378 ( .A1(n6605), .A2(n6604), .ZN(n6622) );
  NAND2_X1 U8379 ( .A1(n8610), .A2(n4414), .ZN(n6609) );
  NAND2_X1 U8380 ( .A1(n6607), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6608) );
  NAND2_X2 U8381 ( .A1(n6609), .A2(n6608), .ZN(n10073) );
  INV_X1 U8382 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9987) );
  INV_X1 U8383 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6610) );
  OR2_X1 U8384 ( .A1(n6310), .A2(n6610), .ZN(n6613) );
  NAND2_X1 U8385 ( .A1(n6263), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6612) );
  OAI211_X1 U8386 ( .C1(n6619), .C2(n9987), .A(n6613), .B(n6612), .ZN(n9789)
         );
  INV_X1 U8387 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U8388 ( .A1(n6615), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U8389 ( .A1(n6263), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6616) );
  OAI211_X1 U8390 ( .C1(n6619), .C2(n6618), .A(n6617), .B(n6616), .ZN(n9610)
         );
  NAND2_X1 U8391 ( .A1(n9789), .A2(n9610), .ZN(n6717) );
  INV_X1 U8392 ( .A(n6717), .ZN(n6620) );
  AOI21_X1 U8393 ( .B1(n10073), .B2(n6834), .A(n6620), .ZN(n6621) );
  INV_X1 U8394 ( .A(n10070), .ZN(n6623) );
  NAND4_X1 U8395 ( .A1(n6623), .A2(n9610), .A3(n6622), .A4(n10073), .ZN(n6624)
         );
  INV_X1 U8396 ( .A(n9610), .ZN(n6702) );
  OR2_X1 U8397 ( .A1(n10073), .A2(n6702), .ZN(n6754) );
  OR2_X1 U8398 ( .A1(n10070), .A2(n6754), .ZN(n6625) );
  NAND2_X1 U8399 ( .A1(n6753), .A2(n6625), .ZN(n6748) );
  NOR2_X1 U8400 ( .A1(n6779), .A2(n4413), .ZN(n6637) );
  INV_X1 U8401 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U8402 ( .A1(n6631), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6632) );
  INV_X1 U8403 ( .A(n6640), .ZN(n6635) );
  NAND2_X1 U8404 ( .A1(n6635), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6636) );
  INV_X1 U8405 ( .A(n7326), .ZN(n8493) );
  NAND2_X1 U8406 ( .A1(n7045), .A2(n8493), .ZN(n6784) );
  NOR4_X1 U8407 ( .A1(n6637), .A2(n6848), .A3(n8425), .A4(n6784), .ZN(n6638)
         );
  NAND2_X1 U8408 ( .A1(n4422), .A2(n6848), .ZN(n7392) );
  OR2_X1 U8409 ( .A1(n7392), .A2(n6874), .ZN(n6832) );
  NAND2_X1 U8410 ( .A1(n6649), .A2(n6648), .ZN(n6641) );
  INV_X1 U8411 ( .A(n6856), .ZN(n6651) );
  NAND2_X1 U8412 ( .A1(n6648), .A2(n6643), .ZN(n6644) );
  OAI21_X1 U8413 ( .B1(n6645), .B2(n6644), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6646) );
  MUX2_X1 U8414 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6646), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6647) );
  INV_X1 U8415 ( .A(n8601), .ZN(n6650) );
  OR2_X1 U8416 ( .A1(n6832), .A2(n7656), .ZN(n7319) );
  XNOR2_X1 U8417 ( .A(n6653), .B(P1_IR_REG_27__SCAN_IN), .ZN(n7433) );
  NAND2_X1 U8418 ( .A1(n7564), .A2(n7433), .ZN(n7447) );
  NOR2_X1 U8419 ( .A1(n7319), .A2(n7447), .ZN(n6714) );
  OAI21_X1 U8420 ( .B1(n6848), .B2(n7326), .A(P1_B_REG_SCAN_IN), .ZN(n6713) );
  INV_X1 U8421 ( .A(n6763), .ZN(n6657) );
  NAND2_X1 U8422 ( .A1(n8003), .A2(n6719), .ZN(n6660) );
  NAND2_X1 U8423 ( .A1(n6660), .A2(n6718), .ZN(n6666) );
  INV_X1 U8424 ( .A(n6767), .ZN(n6721) );
  INV_X1 U8425 ( .A(n6273), .ZN(n8142) );
  AOI21_X1 U8426 ( .B1(n6792), .B2(n6260), .A(n8425), .ZN(n6662) );
  AND2_X1 U8427 ( .A1(n9624), .A2(n6853), .ZN(n6759) );
  INV_X1 U8428 ( .A(n6759), .ZN(n6661) );
  AND4_X1 U8429 ( .A1(n6663), .A2(n6662), .A3(n6760), .A4(n6661), .ZN(n6664)
         );
  OAI211_X1 U8430 ( .C1(n8142), .C2(n8280), .A(n6718), .B(n6664), .ZN(n6665)
         );
  NAND4_X1 U8431 ( .A1(n6666), .A2(n6721), .A3(n8175), .A4(n6665), .ZN(n6667)
         );
  NAND3_X1 U8432 ( .A1(n6668), .A2(n6722), .A3(n6667), .ZN(n6670) );
  NAND3_X1 U8433 ( .A1(n6670), .A2(n6669), .A3(n8521), .ZN(n6671) );
  NAND3_X1 U8434 ( .A1(n6671), .A2(n6731), .A3(n6735), .ZN(n6672) );
  NAND2_X1 U8435 ( .A1(n6673), .A2(n6672), .ZN(n6675) );
  INV_X1 U8436 ( .A(n6737), .ZN(n6674) );
  AOI21_X1 U8437 ( .B1(n6676), .B2(n6675), .A(n6674), .ZN(n6678) );
  OAI21_X1 U8438 ( .B1(n6679), .B2(n6678), .A(n6677), .ZN(n6680) );
  AOI21_X1 U8439 ( .B1(n6681), .B2(n6680), .A(n4842), .ZN(n6706) );
  NAND2_X1 U8440 ( .A1(n6682), .A2(n7347), .ZN(n6699) );
  NAND2_X1 U8441 ( .A1(n6683), .A2(n8632), .ZN(n6684) );
  NAND2_X1 U8442 ( .A1(n6684), .A2(n6840), .ZN(n6685) );
  NAND2_X1 U8443 ( .A1(n6685), .A2(n6692), .ZN(n6686) );
  NAND2_X1 U8444 ( .A1(n6775), .A2(n6686), .ZN(n6694) );
  INV_X1 U8445 ( .A(n6694), .ZN(n6687) );
  NAND4_X1 U8446 ( .A1(n6776), .A2(n6688), .A3(n6687), .A4(n6774), .ZN(n6689)
         );
  NOR2_X1 U8447 ( .A1(n6699), .A2(n6689), .ZN(n6747) );
  INV_X1 U8448 ( .A(n6747), .ZN(n6705) );
  AND3_X1 U8449 ( .A1(n6692), .A2(n6691), .A3(n6690), .ZN(n6693) );
  NOR2_X1 U8450 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  OAI211_X1 U8451 ( .C1(n6696), .C2(n6695), .A(n6776), .B(n6774), .ZN(n6697)
         );
  AND2_X1 U8452 ( .A1(n7346), .A2(n6697), .ZN(n6698) );
  NAND2_X1 U8453 ( .A1(n6701), .A2(n6700), .ZN(n6716) );
  INV_X1 U8454 ( .A(n6716), .ZN(n6704) );
  AND2_X1 U8455 ( .A1(n10073), .A2(n6702), .ZN(n6777) );
  INV_X1 U8456 ( .A(n6777), .ZN(n6703) );
  OAI211_X1 U8457 ( .C1(n6706), .C2(n6705), .A(n6704), .B(n6703), .ZN(n6707)
         );
  NAND2_X1 U8458 ( .A1(n6707), .A2(n6754), .ZN(n6708) );
  NAND2_X1 U8459 ( .A1(n6708), .A2(n6779), .ZN(n6709) );
  NAND2_X1 U8460 ( .A1(n6709), .A2(n6753), .ZN(n6710) );
  NAND4_X1 U8461 ( .A1(n6710), .A2(n9781), .A3(n8493), .A4(n8445), .ZN(n6712)
         );
  OAI211_X1 U8462 ( .C1(n6714), .C2(n6713), .A(n6712), .B(n6711), .ZN(n6715)
         );
  AOI21_X1 U8463 ( .B1(n10073), .B2(n6717), .A(n6716), .ZN(n6750) );
  INV_X1 U8464 ( .A(n8002), .ZN(n6720) );
  NAND2_X1 U8465 ( .A1(n6721), .A2(n8175), .ZN(n6723) );
  NAND2_X1 U8466 ( .A1(n6725), .A2(n6726), .ZN(n8289) );
  INV_X1 U8467 ( .A(n8289), .ZN(n8293) );
  NAND2_X1 U8468 ( .A1(n6728), .A2(n6727), .ZN(n8370) );
  INV_X1 U8469 ( .A(n8370), .ZN(n8358) );
  NAND2_X1 U8470 ( .A1(n6730), .A2(n6729), .ZN(n8346) );
  NAND2_X1 U8471 ( .A1(n6731), .A2(n8521), .ZN(n8588) );
  NOR2_X1 U8472 ( .A1(n6757), .A2(n6733), .ZN(n6734) );
  NOR2_X1 U8473 ( .A1(n9948), .A2(n6738), .ZN(n6739) );
  NAND2_X1 U8474 ( .A1(n6742), .A2(n6744), .ZN(n9915) );
  NAND2_X1 U8475 ( .A1(n6747), .A2(n6835), .ZN(n6749) );
  AOI21_X1 U8476 ( .B1(n6750), .B2(n6749), .A(n6748), .ZN(n6752) );
  OAI21_X1 U8477 ( .B1(n6752), .B2(n6751), .A(n7296), .ZN(n6781) );
  INV_X1 U8478 ( .A(n6753), .ZN(n6778) );
  INV_X1 U8479 ( .A(n6758), .ZN(n6766) );
  OR2_X1 U8480 ( .A1(n8139), .A2(n6759), .ZN(n7648) );
  NOR3_X1 U8481 ( .A1(n7648), .A2(n8409), .A3(n4422), .ZN(n6762) );
  XNOR2_X1 U8482 ( .A(n10169), .B(n9622), .ZN(n10171) );
  NAND4_X1 U8483 ( .A1(n6762), .A2(n8140), .A3(n7840), .A4(n10171), .ZN(n6764)
         );
  NAND2_X2 U8484 ( .A1(n8175), .A2(n6763), .ZN(n8208) );
  NOR2_X1 U8485 ( .A1(n6764), .A2(n8208), .ZN(n6765) );
  NAND4_X1 U8486 ( .A1(n8293), .A2(n6766), .A3(n8002), .A4(n6765), .ZN(n6768)
         );
  NOR4_X1 U8487 ( .A1(n8346), .A2(n6768), .A3(n8370), .A4(n6767), .ZN(n6769)
         );
  NAND4_X1 U8488 ( .A1(n9977), .A2(n4893), .A3(n6732), .A4(n6769), .ZN(n6770)
         );
  AND3_X1 U8489 ( .A1(n9860), .A2(n9904), .A3(n5251), .ZN(n6772) );
  NAND4_X1 U8490 ( .A1(n9843), .A2(n6772), .A3(n9869), .A4(n9884), .ZN(n6773)
         );
  NAND2_X1 U8491 ( .A1(n6774), .A2(n6843), .ZN(n8616) );
  NAND2_X1 U8492 ( .A1(n6776), .A2(n6844), .ZN(n9811) );
  NAND2_X1 U8493 ( .A1(n6780), .A2(n6779), .ZN(n6786) );
  INV_X1 U8494 ( .A(n6782), .ZN(n6789) );
  OAI21_X1 U8495 ( .B1(n6783), .B2(n8505), .A(n4422), .ZN(n6787) );
  INV_X1 U8496 ( .A(n6784), .ZN(n6785) );
  NAND3_X1 U8497 ( .A1(n6787), .A2(n6786), .A3(n5243), .ZN(n6788) );
  NAND3_X1 U8498 ( .A1(n6790), .A2(n6789), .A3(n6788), .ZN(P1_U3242) );
  AND2_X1 U8499 ( .A1(n10004), .A2(n9614), .ZN(n6827) );
  NAND2_X1 U8500 ( .A1(n9624), .A2(n8231), .ZN(n8137) );
  NAND2_X1 U8501 ( .A1(n6791), .A2(n8137), .ZN(n6795) );
  NAND2_X1 U8502 ( .A1(n6795), .A2(n6794), .ZN(n7836) );
  NAND2_X1 U8503 ( .A1(n7836), .A2(n7837), .ZN(n6797) );
  OR2_X1 U8504 ( .A1(n6273), .A2(n8280), .ZN(n6796) );
  OR2_X1 U8505 ( .A1(n10161), .A2(n8412), .ZN(n6798) );
  NOR2_X1 U8506 ( .A1(n10169), .A2(n9622), .ZN(n6800) );
  NAND2_X1 U8507 ( .A1(n10169), .A2(n9622), .ZN(n6799) );
  OR2_X1 U8508 ( .A1(n7105), .A2(n10159), .ZN(n6801) );
  OAI21_X2 U8509 ( .B1(n8000), .B2(n8002), .A(n6801), .ZN(n8202) );
  NAND2_X1 U8510 ( .A1(n8246), .A2(n8210), .ZN(n6804) );
  NOR2_X1 U8511 ( .A1(n10210), .A2(n9621), .ZN(n8172) );
  NOR2_X1 U8512 ( .A1(n8246), .A2(n8210), .ZN(n6803) );
  AOI21_X1 U8513 ( .B1(n8172), .B2(n6804), .A(n6803), .ZN(n6805) );
  NAND2_X1 U8514 ( .A1(n8433), .A2(n8432), .ZN(n8330) );
  OR2_X1 U8515 ( .A1(n8471), .A2(n6377), .ZN(n6807) );
  NAND2_X1 U8516 ( .A1(n8308), .A2(n8486), .ZN(n6808) );
  NAND2_X1 U8517 ( .A1(n8288), .A2(n6808), .ZN(n8371) );
  OR2_X1 U8518 ( .A1(n8490), .A2(n9489), .ZN(n6809) );
  NAND2_X1 U8519 ( .A1(n8348), .A2(n8591), .ZN(n6810) );
  NAND2_X1 U8520 ( .A1(n10103), .A2(n9444), .ZN(n6811) );
  NAND2_X1 U8521 ( .A1(n10058), .A2(n9979), .ZN(n6812) );
  AND2_X1 U8522 ( .A1(n10052), .A2(n9952), .ZN(n6814) );
  OR2_X1 U8523 ( .A1(n10052), .A2(n9952), .ZN(n6813) );
  NAND2_X1 U8524 ( .A1(n9961), .A2(n9978), .ZN(n6816) );
  OR2_X1 U8525 ( .A1(n10043), .A2(n9953), .ZN(n6817) );
  AND2_X1 U8526 ( .A1(n10038), .A2(n9940), .ZN(n6819) );
  OR2_X1 U8527 ( .A1(n10038), .A2(n9940), .ZN(n6818) );
  OR2_X1 U8528 ( .A1(n9475), .A2(n9616), .ZN(n6820) );
  NOR2_X1 U8529 ( .A1(n10028), .A2(n9615), .ZN(n6821) );
  NAND2_X1 U8530 ( .A1(n10028), .A2(n9615), .ZN(n6822) );
  AND2_X1 U8531 ( .A1(n9876), .A2(n9862), .ZN(n6824) );
  OR2_X1 U8532 ( .A1(n10011), .A2(n9861), .ZN(n6825) );
  NOR2_X1 U8533 ( .A1(n10008), .A2(n9844), .ZN(n6826) );
  NOR2_X1 U8534 ( .A1(n6827), .A2(n9823), .ZN(n6828) );
  NAND2_X1 U8535 ( .A1(n9998), .A2(n9613), .ZN(n6829) );
  OR2_X1 U8536 ( .A1(n9816), .A2(n9612), .ZN(n6830) );
  OAI21_X1 U8537 ( .B1(n6831), .B2(n6845), .A(n8639), .ZN(n8659) );
  NAND2_X1 U8538 ( .A1(n6832), .A2(n7311), .ZN(n8234) );
  NAND2_X1 U8539 ( .A1(n4413), .A2(n6848), .ZN(n7050) );
  AND2_X1 U8540 ( .A1(n6874), .A2(n7050), .ZN(n6833) );
  NAND2_X1 U8541 ( .A1(n9870), .A2(n6836), .ZN(n9859) );
  INV_X1 U8542 ( .A(n8632), .ZN(n6838) );
  INV_X1 U8543 ( .A(n9811), .ZN(n9804) );
  NAND2_X1 U8544 ( .A1(n9802), .A2(n6844), .ZN(n6847) );
  INV_X1 U8545 ( .A(n6845), .ZN(n6846) );
  XNOR2_X1 U8546 ( .A(n6847), .B(n6846), .ZN(n6852) );
  NAND2_X1 U8547 ( .A1(n4422), .A2(n7045), .ZN(n6850) );
  NAND2_X1 U8548 ( .A1(n9781), .A2(n6848), .ZN(n6849) );
  OAI22_X1 U8549 ( .A1(n8112), .A2(n9919), .B1(n9587), .B2(n9921), .ZN(n6851)
         );
  INV_X1 U8550 ( .A(n10028), .ZN(n9894) );
  NAND2_X1 U8551 ( .A1(n7842), .A2(n8147), .ZN(n8410) );
  INV_X1 U8552 ( .A(n10210), .ZN(n8216) );
  INV_X1 U8553 ( .A(n8471), .ZN(n8431) );
  NAND2_X1 U8554 ( .A1(n8593), .A2(n8516), .ZN(n9972) );
  INV_X1 U8555 ( .A(n10038), .ZN(n9926) );
  NAND2_X1 U8556 ( .A1(n8626), .A2(n9538), .ZN(n9830) );
  OAI211_X1 U8557 ( .C1(n7303), .C2(n9814), .A(n10174), .B(n7353), .ZN(n8655)
         );
  INV_X1 U8558 ( .A(n7339), .ZN(n6878) );
  NAND2_X1 U8559 ( .A1(n6856), .A2(P1_B_REG_SCAN_IN), .ZN(n6857) );
  MUX2_X1 U8560 ( .A(P1_B_REG_SCAN_IN), .B(n6857), .S(n8601), .Z(n6858) );
  NOR4_X1 U8561 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10303) );
  NOR2_X1 U8562 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n6861) );
  NOR4_X1 U8563 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6860) );
  NOR4_X1 U8564 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6859) );
  NAND4_X1 U8565 ( .A1(n10303), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6867)
         );
  NOR4_X1 U8566 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6865) );
  NOR4_X1 U8567 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6864) );
  NOR4_X1 U8568 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6863) );
  NOR4_X1 U8569 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6862) );
  NAND4_X1 U8570 ( .A1(n6865), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(n6866)
         );
  NOR2_X1 U8571 ( .A1(n6867), .A2(n6866), .ZN(n6868) );
  OR2_X1 U8572 ( .A1(n7392), .A2(n7047), .ZN(n7323) );
  NAND3_X1 U8573 ( .A1(n7294), .A2(n10104), .A3(n7323), .ZN(n8130) );
  NAND2_X1 U8574 ( .A1(n6856), .A2(n10122), .ZN(n10106) );
  INV_X1 U8575 ( .A(n7336), .ZN(n6872) );
  NAND2_X1 U8576 ( .A1(n10122), .A2(n8601), .ZN(n10107) );
  INV_X1 U8577 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6875) );
  OAI21_X1 U8578 ( .B1(n6878), .B2(n10217), .A(n6877), .ZN(P1_U3518) );
  NAND2_X1 U8579 ( .A1(n5933), .A2(n6879), .ZN(n6880) );
  NAND2_X1 U8580 ( .A1(n9261), .A2(n9039), .ZN(n6889) );
  NAND3_X1 U8581 ( .A1(n6882), .A2(n6884), .A3(n6889), .ZN(n6883) );
  AOI21_X1 U8582 ( .B1(n9039), .B2(n6885), .A(n9261), .ZN(n6886) );
  AOI211_X1 U8583 ( .C1(n6879), .C2(n6887), .A(n6886), .B(n6894), .ZN(n6888)
         );
  AOI21_X1 U8584 ( .B1(n6894), .B2(n6889), .A(n6888), .ZN(n6890) );
  OAI21_X1 U8585 ( .B1(n6891), .B2(n6890), .A(n9247), .ZN(n6899) );
  NAND2_X1 U8586 ( .A1(n6913), .A2(P2_B_REG_SCAN_IN), .ZN(n6892) );
  AND2_X1 U8587 ( .A1(n9203), .A2(n6892), .ZN(n9022) );
  AOI22_X1 U8588 ( .A1(n9241), .A2(n9039), .B1(n8904), .B2(n9022), .ZN(n6898)
         );
  INV_X1 U8589 ( .A(n9244), .ZN(n6895) );
  NAND2_X1 U8590 ( .A1(n6896), .A2(n6895), .ZN(n6897) );
  INV_X1 U8591 ( .A(n10243), .ZN(n10234) );
  NOR2_X1 U8592 ( .A1(n6901), .A2(n6900), .ZN(n6903) );
  MUX2_X1 U8593 ( .A(n6904), .B(n6903), .S(n6902), .Z(n6905) );
  INV_X1 U8594 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n10483) );
  INV_X1 U8595 ( .A(n6907), .ZN(n6908) );
  NAND2_X1 U8596 ( .A1(n7038), .A2(n6910), .ZN(n6912) );
  NAND2_X1 U8597 ( .A1(n6912), .A2(n6911), .ZN(n7034) );
  NAND2_X1 U8598 ( .A1(n7034), .A2(n4412), .ZN(n6914) );
  NAND2_X1 U8599 ( .A1(n6914), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8600 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9302) );
  INV_X1 U8601 ( .A(n8927), .ZN(n8940) );
  INV_X1 U8602 ( .A(n8102), .ZN(n7404) );
  AND2_X1 U8603 ( .A1(n7419), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U8604 ( .A1(n4699), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U8605 ( .A1(n6919), .A2(n7382), .ZN(n7469) );
  XNOR2_X1 U8606 ( .A(n6983), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n7470) );
  OR2_X1 U8607 ( .A1(n6983), .A2(n5339), .ZN(n6921) );
  XNOR2_X1 U8608 ( .A(n6992), .B(n6922), .ZN(n7633) );
  INV_X1 U8609 ( .A(n6992), .ZN(n7639) );
  XNOR2_X1 U8610 ( .A(n6998), .B(n10264), .ZN(n7869) );
  INV_X1 U8611 ( .A(n6998), .ZN(n7875) );
  INV_X1 U8612 ( .A(n6927), .ZN(n8096) );
  INV_X1 U8613 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U8614 ( .A(n8102), .B(n8462), .ZN(n8097) );
  XNOR2_X1 U8615 ( .A(n8574), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n8568) );
  INV_X1 U8616 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9314) );
  INV_X1 U8617 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9310) );
  XNOR2_X1 U8618 ( .A(n8927), .B(n10533), .ZN(n8931) );
  INV_X1 U8619 ( .A(n6930), .ZN(n6929) );
  XNOR2_X1 U8620 ( .A(n8968), .B(n9302), .ZN(n8970) );
  NAND2_X1 U8621 ( .A1(n6931), .A2(n8970), .ZN(n8976) );
  INV_X1 U8622 ( .A(n8991), .ZN(n7940) );
  INV_X1 U8623 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9296) );
  OR2_X1 U8624 ( .A1(n7026), .A2(n9296), .ZN(n6935) );
  NAND2_X1 U8625 ( .A1(n7026), .A2(n9296), .ZN(n6934) );
  NAND2_X1 U8626 ( .A1(n6935), .A2(n6934), .ZN(n8997) );
  XNOR2_X1 U8627 ( .A(n6936), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6979) );
  XNOR2_X1 U8628 ( .A(n6937), .B(n6979), .ZN(n6939) );
  NOR2_X1 U8629 ( .A1(n6938), .A2(P2_U3151), .ZN(n9420) );
  NAND2_X1 U8630 ( .A1(n6939), .A2(n9000), .ZN(n7043) );
  XNOR2_X1 U8631 ( .A(n5884), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6981) );
  INV_X1 U8632 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7743) );
  OR2_X1 U8633 ( .A1(n6941), .A2(n7743), .ZN(n6944) );
  NAND2_X1 U8634 ( .A1(n7512), .A2(n6944), .ZN(n6943) );
  NAND3_X1 U8635 ( .A1(n6941), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n7419), .ZN(
        n6942) );
  NAND2_X1 U8636 ( .A1(n6943), .A2(n6942), .ZN(n7502) );
  NAND2_X1 U8637 ( .A1(n7502), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6945) );
  NAND2_X1 U8638 ( .A1(n6945), .A2(n6944), .ZN(n7588) );
  NAND2_X1 U8639 ( .A1(n7379), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6946) );
  XNOR2_X1 U8640 ( .A(n6947), .B(n7524), .ZN(n7516) );
  NAND2_X1 U8641 ( .A1(n7516), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8642 ( .A1(n6947), .A2(n7382), .ZN(n6948) );
  NAND2_X1 U8643 ( .A1(n6949), .A2(n6948), .ZN(n7465) );
  MUX2_X1 U8644 ( .A(n6950), .B(P2_REG2_REG_4__SCAN_IN), .S(n6983), .Z(n7466)
         );
  NAND2_X1 U8645 ( .A1(n7465), .A2(n7466), .ZN(n7464) );
  OR2_X1 U8646 ( .A1(n6983), .A2(n6950), .ZN(n6951) );
  INV_X1 U8647 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8066) );
  NAND2_X1 U8648 ( .A1(n7639), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6954) );
  XNOR2_X1 U8649 ( .A(n6956), .B(n6955), .ZN(n7723) );
  NAND2_X1 U8650 ( .A1(n7723), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6958) );
  INV_X1 U8651 ( .A(n6955), .ZN(n7730) );
  NAND2_X1 U8652 ( .A1(n6956), .A2(n7730), .ZN(n6957) );
  NAND2_X1 U8653 ( .A1(n6958), .A2(n6957), .ZN(n7866) );
  MUX2_X1 U8654 ( .A(n6997), .B(P2_REG2_REG_8__SCAN_IN), .S(n6998), .Z(n7867)
         );
  NAND2_X1 U8655 ( .A1(n7866), .A2(n7867), .ZN(n7865) );
  OR2_X1 U8656 ( .A1(n6998), .A2(n6997), .ZN(n6959) );
  INV_X1 U8657 ( .A(n7005), .ZN(n7951) );
  XNOR2_X1 U8658 ( .A(n8102), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n8093) );
  OR2_X1 U8659 ( .A1(n8102), .A2(n7007), .ZN(n6962) );
  NAND2_X1 U8660 ( .A1(n6963), .A2(n6962), .ZN(n6964) );
  XNOR2_X1 U8661 ( .A(n6964), .B(n8271), .ZN(n8263) );
  NAND2_X1 U8662 ( .A1(n8263), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6966) );
  INV_X1 U8663 ( .A(n8271), .ZN(n7455) );
  NAND2_X1 U8664 ( .A1(n6964), .A2(n7455), .ZN(n6965) );
  NAND2_X1 U8665 ( .A1(n6966), .A2(n6965), .ZN(n8576) );
  MUX2_X1 U8666 ( .A(n9227), .B(P2_REG2_REG_12__SCAN_IN), .S(n8574), .Z(n8577)
         );
  OR2_X1 U8667 ( .A1(n8574), .A2(n9227), .ZN(n6967) );
  NAND2_X1 U8668 ( .A1(n8575), .A2(n6967), .ZN(n6968) );
  XNOR2_X1 U8669 ( .A(n6968), .B(n7017), .ZN(n8913) );
  NAND2_X1 U8670 ( .A1(n8913), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6970) );
  NAND2_X1 U8671 ( .A1(n6968), .A2(n8919), .ZN(n6969) );
  NAND2_X1 U8672 ( .A1(n8927), .A2(n10566), .ZN(n6971) );
  NAND2_X1 U8673 ( .A1(n6973), .A2(n7022), .ZN(n6974) );
  INV_X1 U8674 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9183) );
  XNOR2_X1 U8675 ( .A(n8968), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8959) );
  NOR2_X1 U8676 ( .A1(n8991), .A2(n6975), .ZN(n6976) );
  INV_X1 U8677 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10425) );
  INV_X1 U8678 ( .A(n7026), .ZN(n9009) );
  NAND2_X1 U8679 ( .A1(n9009), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6977) );
  OAI21_X1 U8680 ( .B1(n9009), .B2(P2_REG2_REG_18__SCAN_IN), .A(n6977), .ZN(
        n8996) );
  INV_X1 U8681 ( .A(n6979), .ZN(n6982) );
  MUX2_X1 U8682 ( .A(n6982), .B(n6981), .S(n6980), .Z(n7032) );
  MUX2_X1 U8683 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n7033), .Z(n7019) );
  MUX2_X1 U8684 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n7033), .Z(n7018) );
  MUX2_X1 U8685 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n7033), .Z(n7013) );
  INV_X1 U8686 ( .A(n7013), .ZN(n7014) );
  MUX2_X1 U8687 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n7033), .Z(n6988) );
  INV_X1 U8688 ( .A(n6983), .ZN(n7478) );
  MUX2_X1 U8689 ( .A(n7743), .B(n6984), .S(n7033), .Z(n7412) );
  NAND2_X1 U8690 ( .A1(n7412), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7501) );
  MUX2_X1 U8691 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n7033), .Z(n6985) );
  XNOR2_X1 U8692 ( .A(n6985), .B(n4699), .ZN(n7585) );
  INV_X1 U8693 ( .A(n6985), .ZN(n6986) );
  OAI22_X1 U8694 ( .A1(n7586), .A2(n7585), .B1(n7597), .B2(n6986), .ZN(n7514)
         );
  MUX2_X1 U8695 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n7033), .Z(n6987) );
  XOR2_X1 U8696 ( .A(n7524), .B(n6987), .Z(n7515) );
  NOR2_X1 U8697 ( .A1(n7514), .A2(n7515), .ZN(n7513) );
  NOR2_X1 U8698 ( .A1(n6987), .A2(n7382), .ZN(n7461) );
  XNOR2_X1 U8699 ( .A(n6988), .B(n7478), .ZN(n7460) );
  NOR3_X1 U8700 ( .A1(n7513), .A2(n7461), .A3(n7460), .ZN(n7459) );
  AOI21_X1 U8701 ( .B1(n6988), .B2(n7478), .A(n7459), .ZN(n7528) );
  MUX2_X1 U8702 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n7033), .Z(n6989) );
  XNOR2_X1 U8703 ( .A(n6989), .B(n7535), .ZN(n7527) );
  INV_X1 U8704 ( .A(n6989), .ZN(n6990) );
  OAI22_X1 U8705 ( .A1(n7528), .A2(n7527), .B1(n6991), .B2(n6990), .ZN(n7628)
         );
  MUX2_X1 U8706 ( .A(n8066), .B(n6922), .S(n7033), .Z(n6993) );
  NAND2_X1 U8707 ( .A1(n6993), .A2(n6992), .ZN(n6994) );
  OAI21_X1 U8708 ( .B1(n6993), .B2(n6992), .A(n6994), .ZN(n7627) );
  INV_X1 U8709 ( .A(n6994), .ZN(n7725) );
  MUX2_X1 U8710 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n7033), .Z(n6995) );
  NOR2_X1 U8711 ( .A1(n6995), .A2(n7730), .ZN(n6996) );
  AOI21_X1 U8712 ( .B1(n6995), .B2(n7730), .A(n6996), .ZN(n7724) );
  INV_X1 U8713 ( .A(n6996), .ZN(n7877) );
  MUX2_X1 U8714 ( .A(n6997), .B(n10264), .S(n7033), .Z(n6999) );
  NAND2_X1 U8715 ( .A1(n6999), .A2(n6998), .ZN(n7002) );
  INV_X1 U8716 ( .A(n6999), .ZN(n7000) );
  NAND2_X1 U8717 ( .A1(n7000), .A2(n7875), .ZN(n7001) );
  NAND2_X1 U8718 ( .A1(n7002), .A2(n7001), .ZN(n7876) );
  INV_X1 U8719 ( .A(n7002), .ZN(n7945) );
  MUX2_X1 U8720 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n7033), .Z(n7003) );
  NAND2_X1 U8721 ( .A1(n7951), .A2(n7003), .ZN(n7006) );
  INV_X1 U8722 ( .A(n7003), .ZN(n7004) );
  NAND2_X1 U8723 ( .A1(n7005), .A2(n7004), .ZN(n8104) );
  AND2_X1 U8724 ( .A1(n7006), .A2(n8104), .ZN(n7944) );
  MUX2_X1 U8725 ( .A(n7007), .B(n8462), .S(n7033), .Z(n7008) );
  NAND2_X1 U8726 ( .A1(n7008), .A2(n8102), .ZN(n7011) );
  INV_X1 U8727 ( .A(n7008), .ZN(n7009) );
  NAND2_X1 U8728 ( .A1(n7009), .A2(n7404), .ZN(n7010) );
  NAND2_X1 U8729 ( .A1(n7011), .A2(n7010), .ZN(n8103) );
  AOI21_X1 U8730 ( .B1(n8105), .B2(n8104), .A(n8103), .ZN(n8107) );
  INV_X1 U8731 ( .A(n7011), .ZN(n7012) );
  NOR2_X1 U8732 ( .A1(n8107), .A2(n7012), .ZN(n8267) );
  XOR2_X1 U8733 ( .A(n8271), .B(n7013), .Z(n8266) );
  NOR2_X1 U8734 ( .A1(n8267), .A2(n8266), .ZN(n8265) );
  AOI21_X1 U8735 ( .B1(n8271), .B2(n7014), .A(n8265), .ZN(n8567) );
  MUX2_X1 U8736 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n7033), .Z(n7016) );
  INV_X1 U8737 ( .A(n7016), .ZN(n7015) );
  NAND2_X1 U8738 ( .A1(n7015), .A2(n8574), .ZN(n8563) );
  INV_X1 U8739 ( .A(n8574), .ZN(n7479) );
  AND2_X1 U8740 ( .A1(n7016), .A2(n7479), .ZN(n8564) );
  AOI21_X1 U8741 ( .B1(n8567), .B2(n8563), .A(n8564), .ZN(n8916) );
  XNOR2_X1 U8742 ( .A(n7018), .B(n7017), .ZN(n8915) );
  NAND2_X1 U8743 ( .A1(n8916), .A2(n8915), .ZN(n8914) );
  OAI21_X1 U8744 ( .B1(n7018), .B2(n8919), .A(n8914), .ZN(n8937) );
  XNOR2_X1 U8745 ( .A(n7019), .B(n8927), .ZN(n8936) );
  MUX2_X1 U8746 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n7033), .Z(n7020) );
  XNOR2_X1 U8747 ( .A(n7020), .B(n7022), .ZN(n8950) );
  INV_X1 U8748 ( .A(n7020), .ZN(n7021) );
  MUX2_X1 U8749 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n7033), .Z(n7023) );
  XNOR2_X1 U8750 ( .A(n7023), .B(n8968), .ZN(n8964) );
  MUX2_X1 U8751 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n7033), .Z(n7024) );
  XNOR2_X1 U8752 ( .A(n7024), .B(n8991), .ZN(n8984) );
  INV_X1 U8753 ( .A(n7024), .ZN(n7025) );
  AOI22_X1 U8754 ( .A1(n8983), .A2(n8984), .B1(n8991), .B2(n7025), .ZN(n7027)
         );
  MUX2_X1 U8755 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n7033), .Z(n7028) );
  NAND2_X1 U8756 ( .A1(n7027), .A2(n7028), .ZN(n9008) );
  NAND2_X1 U8757 ( .A1(n9008), .A2(n7026), .ZN(n9005) );
  INV_X1 U8758 ( .A(n7027), .ZN(n7030) );
  INV_X1 U8759 ( .A(n7028), .ZN(n7029) );
  NAND2_X1 U8760 ( .A1(n7030), .A2(n7029), .ZN(n9007) );
  NAND2_X1 U8761 ( .A1(n9005), .A2(n9007), .ZN(n7031) );
  XOR2_X1 U8762 ( .A(n7032), .B(n7031), .Z(n7042) );
  INV_X1 U8763 ( .A(n8606), .ZN(n7720) );
  NOR2_X1 U8764 ( .A1(n7033), .A2(P2_U3151), .ZN(n9423) );
  NAND2_X1 U8765 ( .A1(n7034), .A2(n9423), .ZN(n7036) );
  NOR2_X1 U8766 ( .A1(n7038), .A2(n7037), .ZN(n7039) );
  NAND2_X1 U8767 ( .A1(n8988), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U8768 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8752) );
  OAI211_X1 U8769 ( .C1(n8969), .C2(n5884), .A(n7040), .B(n8752), .ZN(n7041)
         );
  INV_X1 U8770 ( .A(n10004), .ZN(n9835) );
  OAI22_X1 U8771 ( .A1(n9835), .A2(n7170), .B1(n9585), .B2(n4420), .ZN(n7270)
         );
  INV_X1 U8772 ( .A(n7270), .ZN(n7273) );
  NAND2_X4 U8773 ( .A1(n7052), .A2(n7051), .ZN(n7277) );
  NAND2_X2 U8774 ( .A1(n4419), .A2(n7277), .ZN(n7077) );
  NAND2_X1 U8775 ( .A1(n10004), .A2(n7274), .ZN(n7054) );
  NAND2_X1 U8776 ( .A1(n9614), .A2(n7240), .ZN(n7053) );
  NAND2_X1 U8777 ( .A1(n7054), .A2(n7053), .ZN(n7055) );
  XNOR2_X1 U8778 ( .A(n7055), .B(n7277), .ZN(n7271) );
  INV_X1 U8779 ( .A(n7271), .ZN(n7272) );
  NAND2_X1 U8780 ( .A1(n10017), .A2(n7240), .ZN(n7057) );
  NAND2_X1 U8781 ( .A1(n9845), .A2(n7298), .ZN(n7056) );
  NAND2_X1 U8782 ( .A1(n10017), .A2(n7304), .ZN(n7060) );
  NAND2_X1 U8783 ( .A1(n9845), .A2(n7188), .ZN(n7059) );
  NAND2_X1 U8784 ( .A1(n7060), .A2(n7059), .ZN(n7061) );
  XNOR2_X1 U8785 ( .A(n7061), .B(n7301), .ZN(n9454) );
  INV_X1 U8786 ( .A(n6260), .ZN(n7062) );
  NAND2_X1 U8787 ( .A1(n7077), .A2(n7062), .ZN(n7064) );
  OR2_X1 U8788 ( .A1(n6793), .A2(n4420), .ZN(n7066) );
  NAND2_X1 U8789 ( .A1(n7240), .A2(n7062), .ZN(n7065) );
  AND2_X1 U8790 ( .A1(n7066), .A2(n7065), .ZN(n7067) );
  NAND2_X1 U8791 ( .A1(n7077), .A2(n8231), .ZN(n7070) );
  NAND2_X1 U8792 ( .A1(n7188), .A2(n9624), .ZN(n7069) );
  NAND2_X1 U8793 ( .A1(n7070), .A2(n7069), .ZN(n7074) );
  NOR2_X1 U8794 ( .A1(n7369), .A2(n7540), .ZN(n7071) );
  INV_X1 U8795 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7565) );
  INV_X1 U8796 ( .A(n9624), .ZN(n8141) );
  OR2_X1 U8797 ( .A1(n8141), .A2(n4420), .ZN(n7073) );
  NAND2_X1 U8798 ( .A1(n7240), .A2(n8231), .ZN(n7072) );
  OAI211_X1 U8799 ( .C1(n7369), .C2(n7565), .A(n7073), .B(n7072), .ZN(n7562)
         );
  NAND2_X1 U8800 ( .A1(n7563), .A2(n7562), .ZN(n7076) );
  OR2_X1 U8801 ( .A1(n7074), .A2(n7277), .ZN(n7075) );
  NAND2_X1 U8802 ( .A1(n7076), .A2(n7075), .ZN(n7655) );
  NAND2_X1 U8803 ( .A1(n7077), .A2(n8280), .ZN(n7079) );
  NAND2_X1 U8804 ( .A1(n7240), .A2(n6273), .ZN(n7078) );
  NAND2_X1 U8805 ( .A1(n7079), .A2(n7078), .ZN(n7080) );
  XNOR2_X1 U8806 ( .A(n7080), .B(n7301), .ZN(n7083) );
  OR2_X1 U8807 ( .A1(n8142), .A2(n4420), .ZN(n7082) );
  INV_X2 U8808 ( .A(n7170), .ZN(n7188) );
  NAND2_X1 U8809 ( .A1(n7240), .A2(n8280), .ZN(n7081) );
  AND2_X1 U8810 ( .A1(n7082), .A2(n7081), .ZN(n7084) );
  NAND2_X1 U8811 ( .A1(n7083), .A2(n7084), .ZN(n7086) );
  AND2_X1 U8812 ( .A1(n7086), .A2(n7085), .ZN(n7686) );
  NAND2_X1 U8813 ( .A1(n7304), .A2(n8412), .ZN(n7088) );
  NAND2_X1 U8814 ( .A1(n7188), .A2(n10161), .ZN(n7087) );
  NAND2_X1 U8815 ( .A1(n7088), .A2(n7087), .ZN(n7089) );
  XNOR2_X1 U8816 ( .A(n7089), .B(n7301), .ZN(n7100) );
  INV_X1 U8817 ( .A(n10161), .ZN(n7090) );
  OR2_X1 U8818 ( .A1(n7090), .A2(n4421), .ZN(n7092) );
  NAND2_X1 U8819 ( .A1(n7188), .A2(n8412), .ZN(n7091) );
  NAND2_X1 U8820 ( .A1(n7092), .A2(n7091), .ZN(n7098) );
  XNOR2_X1 U8821 ( .A(n7100), .B(n7098), .ZN(n7772) );
  NAND2_X1 U8822 ( .A1(n7304), .A2(n10169), .ZN(n7094) );
  NAND2_X1 U8823 ( .A1(n7240), .A2(n9622), .ZN(n7093) );
  NAND2_X1 U8824 ( .A1(n7094), .A2(n7093), .ZN(n7095) );
  XNOR2_X1 U8825 ( .A(n7095), .B(n7301), .ZN(n7113) );
  OR2_X1 U8826 ( .A1(n8006), .A2(n4420), .ZN(n7097) );
  NAND2_X1 U8827 ( .A1(n7240), .A2(n10169), .ZN(n7096) );
  NAND2_X1 U8828 ( .A1(n7097), .A2(n7096), .ZN(n7114) );
  XNOR2_X1 U8829 ( .A(n7113), .B(n7114), .ZN(n7794) );
  INV_X1 U8830 ( .A(n7098), .ZN(n7099) );
  NAND2_X1 U8831 ( .A1(n7100), .A2(n7099), .ZN(n7795) );
  AND2_X1 U8832 ( .A1(n7794), .A2(n7795), .ZN(n7101) );
  NAND2_X1 U8833 ( .A1(n7770), .A2(n7101), .ZN(n7793) );
  NAND2_X1 U8834 ( .A1(n7105), .A2(n7274), .ZN(n7103) );
  NAND2_X1 U8835 ( .A1(n10159), .A2(n7188), .ZN(n7102) );
  NAND2_X1 U8836 ( .A1(n7103), .A2(n7102), .ZN(n7104) );
  XNOR2_X1 U8837 ( .A(n7104), .B(n7301), .ZN(n7979) );
  NAND2_X1 U8838 ( .A1(n7105), .A2(n7240), .ZN(n7107) );
  OR2_X1 U8839 ( .A1(n6320), .A2(n4420), .ZN(n7106) );
  NAND2_X1 U8840 ( .A1(n10210), .A2(n7274), .ZN(n7109) );
  NAND2_X1 U8841 ( .A1(n9621), .A2(n7240), .ZN(n7108) );
  NAND2_X1 U8842 ( .A1(n7109), .A2(n7108), .ZN(n7110) );
  XNOR2_X1 U8843 ( .A(n7110), .B(n7277), .ZN(n8031) );
  NAND2_X1 U8844 ( .A1(n10210), .A2(n7240), .ZN(n7112) );
  OR2_X1 U8845 ( .A1(n8005), .A2(n4420), .ZN(n7111) );
  NAND2_X1 U8846 ( .A1(n7112), .A2(n7111), .ZN(n8032) );
  NAND2_X1 U8847 ( .A1(n8031), .A2(n8032), .ZN(n8030) );
  INV_X1 U8848 ( .A(n7113), .ZN(n7115) );
  NAND2_X1 U8849 ( .A1(n7115), .A2(n7114), .ZN(n7978) );
  OAI211_X1 U8850 ( .C1(n7979), .C2(n8029), .A(n8030), .B(n7978), .ZN(n7116)
         );
  INV_X1 U8851 ( .A(n7116), .ZN(n7117) );
  NAND2_X1 U8852 ( .A1(n7793), .A2(n7117), .ZN(n7124) );
  INV_X1 U8853 ( .A(n7979), .ZN(n7118) );
  INV_X1 U8854 ( .A(n8029), .ZN(n7119) );
  OAI21_X1 U8855 ( .B1(n7118), .B2(n7119), .A(n8032), .ZN(n7122) );
  INV_X1 U8856 ( .A(n8031), .ZN(n7121) );
  NOR2_X1 U8857 ( .A1(n8032), .A2(n7119), .ZN(n7120) );
  AOI22_X1 U8858 ( .A1(n7122), .A2(n7121), .B1(n7979), .B2(n7120), .ZN(n7123)
         );
  NAND2_X1 U8859 ( .A1(n8246), .A2(n7188), .ZN(n7126) );
  OR2_X1 U8860 ( .A1(n8332), .A2(n4421), .ZN(n7125) );
  AND2_X1 U8861 ( .A1(n7126), .A2(n7125), .ZN(n7931) );
  NAND2_X1 U8862 ( .A1(n8246), .A2(n7274), .ZN(n7128) );
  NAND2_X1 U8863 ( .A1(n7188), .A2(n8210), .ZN(n7127) );
  NAND2_X1 U8864 ( .A1(n7128), .A2(n7127), .ZN(n7129) );
  XNOR2_X1 U8865 ( .A(n7129), .B(n7277), .ZN(n7932) );
  INV_X1 U8866 ( .A(n7931), .ZN(n7130) );
  NAND2_X1 U8867 ( .A1(n8324), .A2(n7274), .ZN(n7132) );
  NAND2_X1 U8868 ( .A1(n9620), .A2(n7230), .ZN(n7131) );
  NAND2_X1 U8869 ( .A1(n7132), .A2(n7131), .ZN(n7133) );
  XNOR2_X1 U8870 ( .A(n7133), .B(n7301), .ZN(n8153) );
  NOR2_X1 U8871 ( .A1(n4420), .A2(n8438), .ZN(n7134) );
  AOI21_X1 U8872 ( .B1(n8324), .B2(n7188), .A(n7134), .ZN(n7140) );
  NAND2_X1 U8873 ( .A1(n8153), .A2(n7140), .ZN(n7135) );
  NAND2_X1 U8874 ( .A1(n8471), .A2(n7274), .ZN(n7137) );
  NAND2_X1 U8875 ( .A1(n6377), .A2(n7240), .ZN(n7136) );
  NAND2_X1 U8876 ( .A1(n7137), .A2(n7136), .ZN(n7138) );
  XNOR2_X1 U8877 ( .A(n7138), .B(n7277), .ZN(n7145) );
  NOR2_X1 U8878 ( .A1(n4420), .A2(n8333), .ZN(n7139) );
  AOI21_X1 U8879 ( .B1(n8471), .B2(n7240), .A(n7139), .ZN(n7146) );
  XNOR2_X1 U8880 ( .A(n7145), .B(n7146), .ZN(n8192) );
  INV_X1 U8881 ( .A(n8153), .ZN(n7141) );
  INV_X1 U8882 ( .A(n7140), .ZN(n8156) );
  NAND2_X1 U8883 ( .A1(n7141), .A2(n8156), .ZN(n7142) );
  AND2_X1 U8884 ( .A1(n8192), .A2(n7142), .ZN(n7143) );
  INV_X1 U8885 ( .A(n7145), .ZN(n7147) );
  NAND2_X1 U8886 ( .A1(n7147), .A2(n7146), .ZN(n7148) );
  OAI22_X1 U8887 ( .A1(n8308), .A2(n7058), .B1(n8486), .B2(n7170), .ZN(n7149)
         );
  XNOR2_X1 U8888 ( .A(n7149), .B(n7301), .ZN(n7151) );
  INV_X1 U8889 ( .A(n7151), .ZN(n7150) );
  OAI22_X1 U8890 ( .A1(n8308), .A2(n7170), .B1(n8486), .B2(n4421), .ZN(n8305)
         );
  NAND2_X1 U8891 ( .A1(n8490), .A2(n7304), .ZN(n7157) );
  NAND2_X1 U8892 ( .A1(n9489), .A2(n7188), .ZN(n7156) );
  NAND2_X1 U8893 ( .A1(n7157), .A2(n7156), .ZN(n7158) );
  XNOR2_X1 U8894 ( .A(n7158), .B(n7277), .ZN(n7162) );
  NAND2_X1 U8895 ( .A1(n8490), .A2(n7188), .ZN(n7161) );
  OR2_X1 U8896 ( .A1(n7159), .A2(n4420), .ZN(n7160) );
  NAND2_X1 U8897 ( .A1(n7161), .A2(n7160), .ZN(n7163) );
  NAND2_X1 U8898 ( .A1(n7162), .A2(n7163), .ZN(n8480) );
  INV_X1 U8899 ( .A(n7162), .ZN(n7165) );
  INV_X1 U8900 ( .A(n7163), .ZN(n7164) );
  NAND2_X1 U8901 ( .A1(n7165), .A2(n7164), .ZN(n8482) );
  OAI22_X1 U8902 ( .A1(n8348), .A2(n7058), .B1(n8591), .B2(n7170), .ZN(n7166)
         );
  XNOR2_X1 U8903 ( .A(n7166), .B(n7301), .ZN(n7169) );
  OAI22_X1 U8904 ( .A1(n8348), .A2(n7170), .B1(n8591), .B2(n4421), .ZN(n7167)
         );
  XNOR2_X1 U8905 ( .A(n7169), .B(n7167), .ZN(n9486) );
  INV_X1 U8906 ( .A(n7167), .ZN(n7168) );
  NAND2_X1 U8907 ( .A1(n9555), .A2(n7274), .ZN(n7172) );
  OR2_X1 U8908 ( .A1(n7170), .A2(n9444), .ZN(n7171) );
  NAND2_X1 U8909 ( .A1(n7172), .A2(n7171), .ZN(n7173) );
  XNOR2_X1 U8910 ( .A(n7173), .B(n7277), .ZN(n7175) );
  NOR2_X1 U8911 ( .A1(n4420), .A2(n9444), .ZN(n7174) );
  AOI21_X1 U8912 ( .B1(n9555), .B2(n7230), .A(n7174), .ZN(n7176) );
  XNOR2_X1 U8913 ( .A(n7175), .B(n7176), .ZN(n9548) );
  INV_X1 U8914 ( .A(n7175), .ZN(n7177) );
  NAND2_X1 U8915 ( .A1(n7177), .A2(n7176), .ZN(n7178) );
  NAND2_X1 U8916 ( .A1(n9961), .A2(n7304), .ZN(n7181) );
  NAND2_X1 U8917 ( .A1(n9978), .A2(n7240), .ZN(n7180) );
  NAND2_X1 U8918 ( .A1(n7181), .A2(n7180), .ZN(n7182) );
  XNOR2_X1 U8919 ( .A(n7182), .B(n7301), .ZN(n9511) );
  NAND2_X1 U8920 ( .A1(n10052), .A2(n7274), .ZN(n7184) );
  NAND2_X1 U8921 ( .A1(n7240), .A2(n9952), .ZN(n7183) );
  NAND2_X1 U8922 ( .A1(n7184), .A2(n7183), .ZN(n7185) );
  XNOR2_X1 U8923 ( .A(n7185), .B(n7301), .ZN(n9507) );
  NAND2_X1 U8924 ( .A1(n10052), .A2(n7188), .ZN(n7187) );
  NAND2_X1 U8925 ( .A1(n7298), .A2(n9952), .ZN(n7186) );
  NAND2_X1 U8926 ( .A1(n10058), .A2(n7274), .ZN(n7190) );
  NAND2_X1 U8927 ( .A1(n7240), .A2(n9979), .ZN(n7189) );
  NAND2_X1 U8928 ( .A1(n7190), .A2(n7189), .ZN(n7191) );
  XNOR2_X1 U8929 ( .A(n7191), .B(n7301), .ZN(n9506) );
  NOR2_X1 U8930 ( .A1(n8590), .A2(n4421), .ZN(n7192) );
  AOI21_X1 U8931 ( .B1(n10058), .B2(n7188), .A(n7192), .ZN(n9441) );
  NAND2_X1 U8932 ( .A1(n9506), .A2(n9441), .ZN(n7193) );
  NAND2_X1 U8933 ( .A1(n7194), .A2(n7193), .ZN(n7203) );
  INV_X1 U8934 ( .A(n7194), .ZN(n7195) );
  OR3_X1 U8935 ( .A1(n7195), .A2(n9506), .A3(n9441), .ZN(n7201) );
  OAI21_X1 U8936 ( .B1(n9507), .B2(n9597), .A(n9510), .ZN(n7199) );
  INV_X1 U8937 ( .A(n9511), .ZN(n7198) );
  INV_X1 U8938 ( .A(n9597), .ZN(n7196) );
  INV_X1 U8939 ( .A(n9507), .ZN(n9508) );
  AOI22_X1 U8940 ( .A1(n7199), .A2(n7198), .B1(n7197), .B2(n9508), .ZN(n7200)
         );
  NAND2_X1 U8941 ( .A1(n10043), .A2(n7304), .ZN(n7205) );
  NAND2_X1 U8942 ( .A1(n9953), .A2(n7240), .ZN(n7204) );
  NAND2_X1 U8943 ( .A1(n7205), .A2(n7204), .ZN(n7206) );
  XNOR2_X1 U8944 ( .A(n7206), .B(n7277), .ZN(n7209) );
  NAND2_X1 U8945 ( .A1(n10043), .A2(n7240), .ZN(n7208) );
  NAND2_X1 U8946 ( .A1(n9953), .A2(n7298), .ZN(n7207) );
  NAND2_X1 U8947 ( .A1(n7208), .A2(n7207), .ZN(n7210) );
  AND2_X1 U8948 ( .A1(n7209), .A2(n7210), .ZN(n9520) );
  INV_X1 U8949 ( .A(n7209), .ZN(n7212) );
  INV_X1 U8950 ( .A(n7210), .ZN(n7211) );
  NAND2_X1 U8951 ( .A1(n9475), .A2(n7274), .ZN(n7214) );
  NAND2_X1 U8952 ( .A1(n9616), .A2(n7230), .ZN(n7213) );
  NAND2_X1 U8953 ( .A1(n7214), .A2(n7213), .ZN(n7215) );
  XNOR2_X1 U8954 ( .A(n7215), .B(n7277), .ZN(n9469) );
  NAND2_X1 U8955 ( .A1(n9475), .A2(n7188), .ZN(n7217) );
  NAND2_X1 U8956 ( .A1(n9616), .A2(n7298), .ZN(n7216) );
  NAND2_X1 U8957 ( .A1(n7217), .A2(n7216), .ZN(n7224) );
  NAND2_X1 U8958 ( .A1(n10038), .A2(n7274), .ZN(n7219) );
  NAND2_X1 U8959 ( .A1(n9940), .A2(n7188), .ZN(n7218) );
  NAND2_X1 U8960 ( .A1(n7219), .A2(n7218), .ZN(n7220) );
  XNOR2_X1 U8961 ( .A(n7220), .B(n7277), .ZN(n7225) );
  NAND2_X1 U8962 ( .A1(n10038), .A2(n7240), .ZN(n7222) );
  NAND2_X1 U8963 ( .A1(n9940), .A2(n7298), .ZN(n7221) );
  NAND2_X1 U8964 ( .A1(n7222), .A2(n7221), .ZN(n9570) );
  OAI22_X1 U8965 ( .A1(n9469), .A2(n7224), .B1(n7225), .B2(n9570), .ZN(n7229)
         );
  INV_X1 U8966 ( .A(n7225), .ZN(n9467) );
  INV_X1 U8967 ( .A(n9570), .ZN(n7223) );
  INV_X1 U8968 ( .A(n7224), .ZN(n9468) );
  OAI21_X1 U8969 ( .B1(n9467), .B2(n7223), .A(n9468), .ZN(n7227) );
  AND2_X1 U8970 ( .A1(n7224), .A2(n9570), .ZN(n7226) );
  AOI22_X1 U8971 ( .A1(n9469), .A2(n7227), .B1(n7226), .B2(n7225), .ZN(n7228)
         );
  NAND2_X1 U8972 ( .A1(n10028), .A2(n7274), .ZN(n7232) );
  NAND2_X1 U8973 ( .A1(n9615), .A2(n7230), .ZN(n7231) );
  NAND2_X1 U8974 ( .A1(n7232), .A2(n7231), .ZN(n7233) );
  XNOR2_X1 U8975 ( .A(n7233), .B(n7301), .ZN(n9540) );
  AND2_X1 U8976 ( .A1(n9615), .A2(n7298), .ZN(n7234) );
  AOI21_X1 U8977 ( .B1(n10028), .B2(n7240), .A(n7234), .ZN(n7236) );
  NAND2_X1 U8978 ( .A1(n9540), .A2(n7236), .ZN(n7235) );
  INV_X1 U8979 ( .A(n9540), .ZN(n7237) );
  INV_X1 U8980 ( .A(n7236), .ZN(n9539) );
  NAND2_X1 U8981 ( .A1(n7237), .A2(n9539), .ZN(n7238) );
  NAND2_X1 U8982 ( .A1(n9876), .A2(n7304), .ZN(n7242) );
  NAND2_X1 U8983 ( .A1(n9862), .A2(n7188), .ZN(n7241) );
  NAND2_X1 U8984 ( .A1(n7242), .A2(n7241), .ZN(n7243) );
  XNOR2_X1 U8985 ( .A(n7243), .B(n7301), .ZN(n7246) );
  AND2_X1 U8986 ( .A1(n9862), .A2(n7298), .ZN(n7244) );
  AOI21_X1 U8987 ( .B1(n9876), .B2(n7188), .A(n7244), .ZN(n7245) );
  XNOR2_X1 U8988 ( .A(n7246), .B(n7245), .ZN(n9479) );
  NAND2_X1 U8989 ( .A1(n7246), .A2(n7245), .ZN(n7247) );
  NAND2_X1 U8990 ( .A1(n10011), .A2(n7304), .ZN(n7249) );
  NAND2_X1 U8991 ( .A1(n9861), .A2(n7240), .ZN(n7248) );
  NAND2_X1 U8992 ( .A1(n7249), .A2(n7248), .ZN(n7250) );
  XNOR2_X1 U8993 ( .A(n7250), .B(n7277), .ZN(n7254) );
  NAND2_X1 U8994 ( .A1(n10011), .A2(n7230), .ZN(n7252) );
  NAND2_X1 U8995 ( .A1(n9861), .A2(n7298), .ZN(n7251) );
  NAND2_X1 U8996 ( .A1(n7252), .A2(n7251), .ZN(n7255) );
  NAND2_X1 U8997 ( .A1(n7254), .A2(n7255), .ZN(n9456) );
  INV_X1 U8998 ( .A(n9454), .ZN(n9452) );
  INV_X1 U8999 ( .A(n9560), .ZN(n7253) );
  NOR2_X1 U9000 ( .A1(n9452), .A2(n7253), .ZN(n7258) );
  INV_X1 U9001 ( .A(n7254), .ZN(n7257) );
  INV_X1 U9002 ( .A(n7255), .ZN(n7256) );
  AND2_X1 U9003 ( .A1(n7257), .A2(n7256), .ZN(n9529) );
  AOI21_X1 U9004 ( .B1(n7258), .B2(n9456), .A(n9529), .ZN(n7268) );
  NAND2_X1 U9005 ( .A1(n10008), .A2(n7304), .ZN(n7260) );
  NAND2_X1 U9006 ( .A1(n9844), .A2(n7240), .ZN(n7259) );
  NAND2_X1 U9007 ( .A1(n7260), .A2(n7259), .ZN(n7261) );
  XNOR2_X1 U9008 ( .A(n7261), .B(n7301), .ZN(n7263) );
  AND2_X1 U9009 ( .A1(n9844), .A2(n7298), .ZN(n7262) );
  AOI21_X1 U9010 ( .B1(n10008), .B2(n7188), .A(n7262), .ZN(n7264) );
  NAND2_X1 U9011 ( .A1(n7263), .A2(n7264), .ZN(n7269) );
  INV_X1 U9012 ( .A(n7263), .ZN(n7266) );
  INV_X1 U9013 ( .A(n7264), .ZN(n7265) );
  NAND2_X1 U9014 ( .A1(n7266), .A2(n7265), .ZN(n7267) );
  XNOR2_X1 U9015 ( .A(n7271), .B(n7270), .ZN(n9498) );
  NAND2_X1 U9016 ( .A1(n9998), .A2(n7274), .ZN(n7276) );
  NAND2_X1 U9017 ( .A1(n9613), .A2(n7188), .ZN(n7275) );
  NAND2_X1 U9018 ( .A1(n7276), .A2(n7275), .ZN(n7278) );
  XNOR2_X1 U9019 ( .A(n7278), .B(n7277), .ZN(n7282) );
  NOR2_X1 U9020 ( .A1(n9828), .A2(n4420), .ZN(n7279) );
  AOI21_X1 U9021 ( .B1(n9998), .B2(n7240), .A(n7279), .ZN(n7280) );
  XNOR2_X1 U9022 ( .A(n7282), .B(n7280), .ZN(n9581) );
  INV_X1 U9023 ( .A(n7280), .ZN(n7281) );
  NAND2_X1 U9024 ( .A1(n7282), .A2(n7281), .ZN(n9433) );
  INV_X1 U9025 ( .A(n9433), .ZN(n7293) );
  NAND2_X1 U9026 ( .A1(n9816), .A2(n7304), .ZN(n7284) );
  NAND2_X1 U9027 ( .A1(n9612), .A2(n7230), .ZN(n7283) );
  NAND2_X1 U9028 ( .A1(n7284), .A2(n7283), .ZN(n7285) );
  XNOR2_X1 U9029 ( .A(n7285), .B(n7301), .ZN(n7289) );
  INV_X1 U9030 ( .A(n7289), .ZN(n7291) );
  NOR2_X1 U9031 ( .A1(n9587), .A2(n4421), .ZN(n7287) );
  AOI21_X1 U9032 ( .B1(n9816), .B2(n7240), .A(n7287), .ZN(n7288) );
  INV_X1 U9033 ( .A(n7288), .ZN(n7290) );
  AOI21_X1 U9034 ( .B1(n7291), .B2(n7290), .A(n7310), .ZN(n9432) );
  INV_X1 U9035 ( .A(n9432), .ZN(n7292) );
  INV_X1 U9036 ( .A(n8131), .ZN(n7295) );
  NOR2_X1 U9037 ( .A1(n7320), .A2(n7656), .ZN(n7297) );
  NAND2_X1 U9038 ( .A1(n8652), .A2(n7230), .ZN(n7300) );
  NAND2_X1 U9039 ( .A1(n9611), .A2(n7298), .ZN(n7299) );
  NAND2_X1 U9040 ( .A1(n7300), .A2(n7299), .ZN(n7302) );
  XNOR2_X1 U9041 ( .A(n7302), .B(n7301), .ZN(n7306) );
  AOI22_X1 U9042 ( .A1(n8652), .A2(n7274), .B1(n7188), .B2(n9611), .ZN(n7305)
         );
  XNOR2_X1 U9043 ( .A(n7306), .B(n7305), .ZN(n7309) );
  NAND3_X1 U9044 ( .A1(n7307), .A2(n9598), .A3(n7310), .ZN(n7331) );
  OR2_X1 U9045 ( .A1(n7311), .A2(n8445), .ZN(n8135) );
  NOR2_X1 U9046 ( .A1(n8135), .A2(n7656), .ZN(n7312) );
  NAND2_X1 U9047 ( .A1(n7318), .A2(n7312), .ZN(n7313) );
  INV_X1 U9048 ( .A(n7319), .ZN(n7314) );
  NAND2_X1 U9049 ( .A1(n7318), .A2(n7314), .ZN(n7316) );
  OAI22_X1 U9050 ( .A1(n9587), .A2(n9584), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7315), .ZN(n7329) );
  INV_X1 U9051 ( .A(n7316), .ZN(n7317) );
  AND2_X2 U9052 ( .A1(n7317), .A2(n10115), .ZN(n9600) );
  INV_X1 U9053 ( .A(n9600), .ZN(n9586) );
  INV_X1 U9054 ( .A(n7318), .ZN(n7322) );
  NAND3_X1 U9055 ( .A1(n7320), .A2(n7319), .A3(n8135), .ZN(n7321) );
  NAND2_X1 U9056 ( .A1(n7322), .A2(n7321), .ZN(n7324) );
  NAND2_X1 U9057 ( .A1(n7324), .A2(n7323), .ZN(n7657) );
  INV_X1 U9058 ( .A(n7369), .ZN(n7325) );
  OAI21_X1 U9059 ( .B1(n7657), .B2(n7325), .A(P1_STATE_REG_SCAN_IN), .ZN(n7327) );
  OAI22_X1 U9060 ( .A1(n8112), .A2(n9586), .B1(n9603), .B2(n8650), .ZN(n7328)
         );
  AOI211_X1 U9061 ( .C1(n8652), .C2(n9576), .A(n7329), .B(n7328), .ZN(n7330)
         );
  INV_X1 U9062 ( .A(n7333), .ZN(n7334) );
  NOR2_X1 U9063 ( .A1(n10225), .A2(n7340), .ZN(n7341) );
  NAND2_X1 U9064 ( .A1(n7343), .A2(n7342), .ZN(P1_U3550) );
  NAND2_X1 U9065 ( .A1(n8652), .A2(n9611), .ZN(n8638) );
  NOR2_X1 U9066 ( .A1(n7344), .A2(n10215), .ZN(n7345) );
  NAND2_X1 U9067 ( .A1(n8639), .A2(n5246), .ZN(n7357) );
  NAND2_X1 U9068 ( .A1(n9611), .A2(n10160), .ZN(n7349) );
  NAND2_X1 U9069 ( .A1(n7433), .A2(P1_B_REG_SCAN_IN), .ZN(n9788) );
  NAND3_X1 U9070 ( .A1(n10158), .A2(n9610), .A3(n9788), .ZN(n7348) );
  NAND2_X1 U9071 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  OAI211_X1 U9072 ( .C1(n7362), .C2(n5035), .A(n10174), .B(n9794), .ZN(n8644)
         );
  NAND3_X1 U9073 ( .A1(n4781), .A2(n7344), .A3(n10206), .ZN(n7355) );
  INV_X1 U9074 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7363) );
  NOR2_X1 U9075 ( .A1(n10218), .A2(n7363), .ZN(n7364) );
  NAND2_X1 U9076 ( .A1(n7366), .A2(n7365), .ZN(P1_U3519) );
  INV_X1 U9077 ( .A(n7367), .ZN(n7368) );
  NAND2_X1 U9078 ( .A1(n5347), .A2(n4410), .ZN(n10118) );
  INV_X1 U9079 ( .A(n10118), .ZN(n10110) );
  AOI22_X1 U9080 ( .A1(n10110), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n9628), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n7371) );
  OAI21_X1 U9081 ( .B1(n7381), .B2(n10121), .A(n7371), .ZN(P1_U3354) );
  INV_X1 U9082 ( .A(n7372), .ZN(n7383) );
  AOI22_X1 U9083 ( .A1(n9639), .A2(P1_STATE_REG_SCAN_IN), .B1(n10110), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n7373) );
  OAI21_X1 U9084 ( .B1(n7383), .B2(n10121), .A(n7373), .ZN(P1_U3352) );
  INV_X1 U9085 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7376) );
  INV_X1 U9086 ( .A(n7582), .ZN(n7375) );
  OAI222_X1 U9087 ( .A1(n10118), .A2(n7376), .B1(n10121), .B2(n4814), .C1(
        n4410), .C2(n7375), .ZN(P1_U3353) );
  INV_X1 U9088 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7377) );
  INV_X1 U9089 ( .A(n7561), .ZN(n7426) );
  OAI222_X1 U9090 ( .A1(n10118), .A2(n7377), .B1(n10121), .B2(n7398), .C1(
        n7426), .C2(n4410), .ZN(P1_U3351) );
  NOR2_X1 U9091 ( .A1(n7378), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9424) );
  INV_X2 U9092 ( .A(n9424), .ZN(n9427) );
  NAND2_X1 U9093 ( .A1(n7378), .A2(P2_U3151), .ZN(n9429) );
  OAI222_X1 U9094 ( .A1(n9427), .A2(n7380), .B1(n9429), .B2(n4814), .C1(
        P2_U3151), .C2(n4699), .ZN(P2_U3293) );
  OAI222_X1 U9095 ( .A1(n9427), .A2(n5285), .B1(n9429), .B2(n7381), .C1(n4639), 
        .C2(P2_U3151), .ZN(P2_U3294) );
  OAI222_X1 U9096 ( .A1(n9427), .A2(n5325), .B1(n9429), .B2(n7383), .C1(n7382), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  INV_X1 U9097 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7384) );
  INV_X1 U9098 ( .A(n7613), .ZN(n7618) );
  OAI222_X1 U9099 ( .A1(n10118), .A2(n7384), .B1(n10121), .B2(n7385), .C1(
        n7618), .C2(n4410), .ZN(P1_U3348) );
  OAI222_X1 U9100 ( .A1(P2_U3151), .A2(n7730), .B1(n9427), .B2(n4861), .C1(
        n7385), .C2(n9429), .ZN(P2_U3288) );
  INV_X1 U9101 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7386) );
  INV_X1 U9102 ( .A(n7444), .ZN(n9665) );
  OAI222_X1 U9103 ( .A1(n10118), .A2(n7386), .B1(n10121), .B2(n6298), .C1(
        n9665), .C2(n4410), .ZN(P1_U3349) );
  INV_X1 U9104 ( .A(n7387), .ZN(n7396) );
  AOI22_X1 U9105 ( .A1(n9657), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10110), .ZN(n7388) );
  OAI21_X1 U9106 ( .B1(n7396), .B2(n10121), .A(n7388), .ZN(P1_U3350) );
  NAND2_X1 U9107 ( .A1(P1_U3973), .A2(n9789), .ZN(n7389) );
  OAI21_X1 U9108 ( .B1(P1_U3973), .B2(n6082), .A(n7389), .ZN(P1_U3585) );
  INV_X1 U9109 ( .A(n7390), .ZN(n7391) );
  OR2_X1 U9110 ( .A1(n7392), .A2(n7391), .ZN(n7394) );
  INV_X1 U9111 ( .A(n7432), .ZN(n7395) );
  OR2_X1 U9112 ( .A1(n10104), .A2(n8493), .ZN(n7431) );
  AND2_X1 U9113 ( .A1(n9786), .A2(n9623), .ZN(P1_U3085) );
  OAI222_X1 U9114 ( .A1(n9427), .A2(n5370), .B1(n9429), .B2(n7396), .C1(
        P2_U3151), .C2(n7535), .ZN(P2_U3290) );
  NAND2_X1 U9115 ( .A1(n8210), .A2(P1_U3973), .ZN(n7397) );
  OAI21_X1 U9116 ( .B1(P1_U3973), .B2(n4861), .A(n7397), .ZN(P1_U3561) );
  INV_X1 U9117 ( .A(n9429), .ZN(n8508) );
  INV_X1 U9118 ( .A(n8508), .ZN(n8605) );
  OAI222_X1 U9119 ( .A1(n9427), .A2(n5379), .B1(n8605), .B2(n6298), .C1(n7639), 
        .C2(P2_U3151), .ZN(P2_U3289) );
  OAI222_X1 U9120 ( .A1(n9427), .A2(n4643), .B1(n8605), .B2(n7398), .C1(n7478), 
        .C2(P2_U3151), .ZN(P2_U3291) );
  AOI22_X1 U9121 ( .A1(n9690), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10110), .ZN(n7399) );
  OAI21_X1 U9122 ( .B1(n7405), .B2(n10121), .A(n7399), .ZN(P1_U3345) );
  INV_X1 U9123 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7403) );
  INV_X1 U9124 ( .A(n7748), .ZN(n7402) );
  AOI22_X1 U9125 ( .A1(n8609), .A2(n7403), .B1(n8606), .B2(n7402), .ZN(
        P2_U3376) );
  OAI222_X1 U9126 ( .A1(n9427), .A2(n4738), .B1(n9429), .B2(n7405), .C1(n7404), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U9127 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10371) );
  INV_X1 U9128 ( .A(n7406), .ZN(n7407) );
  INV_X1 U9129 ( .A(n7488), .ZN(n7483) );
  OAI222_X1 U9130 ( .A1(n10118), .A2(n10371), .B1(n10121), .B2(n7407), .C1(
        n4410), .C2(n7483), .ZN(P1_U3347) );
  OAI222_X1 U9131 ( .A1(n9427), .A2(n4743), .B1(n9429), .B2(n7407), .C1(
        P2_U3151), .C2(n7875), .ZN(P2_U3287) );
  NAND2_X1 U9132 ( .A1(n9489), .A2(P1_U3973), .ZN(n7408) );
  OAI21_X1 U9133 ( .B1(P1_U3973), .B2(n4627), .A(n7408), .ZN(P1_U3565) );
  AND2_X1 U9134 ( .A1(n8609), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U9135 ( .A1(n8609), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U9136 ( .A1(n8609), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U9137 ( .A1(n8609), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U9138 ( .A1(n8609), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U9139 ( .A1(n8609), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U9140 ( .A1(n8609), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U9141 ( .A1(n8609), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U9142 ( .A1(n8609), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U9143 ( .A1(n8609), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U9144 ( .A1(n8609), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U9145 ( .A1(n8609), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U9146 ( .A1(n8609), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U9147 ( .A1(n8609), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U9148 ( .A1(n8609), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U9149 ( .A1(n8609), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U9150 ( .A1(n8609), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U9151 ( .A1(n8609), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U9152 ( .A1(n8609), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U9153 ( .A1(n8609), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U9154 ( .A1(n8609), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U9155 ( .A1(n8609), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U9156 ( .A1(n8609), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U9157 ( .A(n6366), .ZN(n7410) );
  OAI222_X1 U9158 ( .A1(n9427), .A2(n7409), .B1(n9429), .B2(n7410), .C1(n7951), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U9159 ( .A(n7491), .ZN(n7603) );
  OAI222_X1 U9160 ( .A1(n4410), .A2(n7603), .B1(n10118), .B2(n5451), .C1(n7410), .C2(n10121), .ZN(P1_U3346) );
  INV_X1 U9161 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10490) );
  NOR2_X1 U9162 ( .A1(n7411), .A2(n10490), .ZN(P2_U3261) );
  INV_X1 U9163 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10415) );
  NOR2_X1 U9164 ( .A1(n7411), .A2(n10415), .ZN(P2_U3256) );
  INV_X1 U9165 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10418) );
  NOR2_X1 U9166 ( .A1(n7411), .A2(n10418), .ZN(P2_U3255) );
  INV_X1 U9167 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10454) );
  NOR2_X1 U9168 ( .A1(n7411), .A2(n10454), .ZN(P2_U3262) );
  INV_X1 U9169 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10358) );
  NOR2_X1 U9170 ( .A1(n7411), .A2(n10358), .ZN(P2_U3243) );
  INV_X1 U9171 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10453) );
  NOR2_X1 U9172 ( .A1(n7411), .A2(n10453), .ZN(P2_U3249) );
  INV_X1 U9173 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10534) );
  NOR2_X1 U9174 ( .A1(n7411), .A2(n10534), .ZN(P2_U3253) );
  OAI21_X1 U9175 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7412), .A(n7501), .ZN(n7413) );
  OAI21_X1 U9176 ( .B1(n8980), .B2(n7414), .A(n7413), .ZN(n7415) );
  OAI21_X1 U9177 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7416), .A(n7415), .ZN(n7417) );
  AOI21_X1 U9178 ( .B1(n8988), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n7417), .ZN(
        n7418) );
  OAI21_X1 U9179 ( .B1(n7419), .B2(n8969), .A(n7418), .ZN(P2_U3182) );
  AND2_X1 U9180 ( .A1(n7613), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7430) );
  XNOR2_X1 U9181 ( .A(n7582), .B(n7420), .ZN(n7576) );
  AND2_X1 U9182 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9632) );
  NAND2_X1 U9183 ( .A1(n9628), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7421) );
  OAI211_X1 U9184 ( .C1(n9628), .C2(P1_REG1_REG_1__SCAN_IN), .A(n9632), .B(
        n7421), .ZN(n9630) );
  NAND2_X1 U9185 ( .A1(n9630), .A2(n7421), .ZN(n7574) );
  NAND2_X1 U9186 ( .A1(n7576), .A2(n7574), .ZN(n7423) );
  NAND2_X1 U9187 ( .A1(n7582), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7422) );
  NAND2_X1 U9188 ( .A1(n7423), .A2(n7422), .ZN(n9644) );
  MUX2_X1 U9189 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n7424), .S(n9639), .Z(n9645)
         );
  NAND2_X1 U9190 ( .A1(n9639), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7555) );
  MUX2_X1 U9191 ( .A(n7425), .B(P1_REG1_REG_4__SCAN_IN), .S(n7561), .Z(n7554)
         );
  NOR2_X1 U9192 ( .A1(n7426), .A2(n7425), .ZN(n9656) );
  INV_X1 U9193 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7427) );
  MUX2_X1 U9194 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7427), .S(n9657), .Z(n7428)
         );
  NAND2_X1 U9195 ( .A1(n9657), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9673) );
  INV_X1 U9196 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10223) );
  MUX2_X1 U9197 ( .A(n10223), .B(P1_REG1_REG_6__SCAN_IN), .S(n7444), .Z(n9672)
         );
  NOR2_X1 U9198 ( .A1(n9665), .A2(n10223), .ZN(n7614) );
  NOR2_X1 U9199 ( .A1(n9671), .A2(n7614), .ZN(n7429) );
  NOR2_X1 U9200 ( .A1(n7626), .A2(n7430), .ZN(n7485) );
  XNOR2_X1 U9201 ( .A(n7488), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7484) );
  XNOR2_X1 U9202 ( .A(n7485), .B(n7484), .ZN(n7452) );
  INV_X1 U9203 ( .A(n7547), .ZN(n7434) );
  NOR2_X2 U9204 ( .A1(n7434), .A2(n7564), .ZN(n9777) );
  INV_X1 U9205 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U9206 ( .A1(n4410), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8157) );
  OAI21_X1 U9207 ( .B1(n9786), .B2(n7435), .A(n8157), .ZN(n7436) );
  AOI21_X1 U9208 ( .B1(n9777), .B2(n7488), .A(n7436), .ZN(n7451) );
  MUX2_X1 U9209 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n8378), .S(n7488), .Z(n7449)
         );
  XNOR2_X1 U9210 ( .A(n7582), .B(n8277), .ZN(n7573) );
  INV_X1 U9211 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10482) );
  XNOR2_X1 U9212 ( .A(n9628), .B(n10482), .ZN(n9635) );
  AND2_X1 U9213 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9634) );
  NAND2_X1 U9214 ( .A1(n9635), .A2(n9634), .ZN(n9633) );
  NAND2_X1 U9215 ( .A1(n9628), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9216 ( .A1(n9633), .A2(n7437), .ZN(n7572) );
  NAND2_X1 U9217 ( .A1(n7573), .A2(n7572), .ZN(n7571) );
  NAND2_X1 U9218 ( .A1(n7582), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7438) );
  NAND2_X1 U9219 ( .A1(n7571), .A2(n7438), .ZN(n9641) );
  INV_X1 U9220 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7439) );
  XNOR2_X1 U9221 ( .A(n9639), .B(n7439), .ZN(n9642) );
  NAND2_X1 U9222 ( .A1(n9641), .A2(n9642), .ZN(n9640) );
  NAND2_X1 U9223 ( .A1(n9639), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U9224 ( .A1(n9640), .A2(n7440), .ZN(n7551) );
  XNOR2_X1 U9225 ( .A(n7561), .B(n7441), .ZN(n7552) );
  NAND2_X1 U9226 ( .A1(n7551), .A2(n7552), .ZN(n7550) );
  NAND2_X1 U9227 ( .A1(n7561), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U9228 ( .A1(n7550), .A2(n7442), .ZN(n9654) );
  MUX2_X1 U9229 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n8223), .S(n9657), .Z(n9655)
         );
  NAND2_X1 U9230 ( .A1(n9654), .A2(n9655), .ZN(n9653) );
  NAND2_X1 U9231 ( .A1(n9657), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7443) );
  NAND2_X1 U9232 ( .A1(n9653), .A2(n7443), .ZN(n9669) );
  MUX2_X1 U9233 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n8212), .S(n7444), .Z(n9670)
         );
  NAND2_X1 U9234 ( .A1(n9669), .A2(n9670), .ZN(n9668) );
  NAND2_X1 U9235 ( .A1(n7444), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7445) );
  NAND2_X1 U9236 ( .A1(n9668), .A2(n7445), .ZN(n7621) );
  INV_X1 U9237 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8244) );
  XNOR2_X1 U9238 ( .A(n7613), .B(n8244), .ZN(n7622) );
  NAND2_X1 U9239 ( .A1(n7621), .A2(n7622), .ZN(n7620) );
  NAND2_X1 U9240 ( .A1(n7613), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7446) );
  NAND2_X1 U9241 ( .A1(n7620), .A2(n7446), .ZN(n7448) );
  INV_X1 U9242 ( .A(n7447), .ZN(n7567) );
  NAND2_X1 U9243 ( .A1(n7448), .A2(n7449), .ZN(n7490) );
  OAI211_X1 U9244 ( .C1(n7449), .C2(n7448), .A(n9773), .B(n7490), .ZN(n7450)
         );
  OAI211_X1 U9245 ( .C1(n7452), .C2(n9743), .A(n7451), .B(n7450), .ZN(P1_U3251) );
  NAND2_X1 U9246 ( .A1(P2_U3893), .A2(n8742), .ZN(n7453) );
  OAI21_X1 U9247 ( .B1(P2_U3893), .B2(n5451), .A(n7453), .ZN(P2_U3500) );
  INV_X1 U9248 ( .A(n7454), .ZN(n7456) );
  OAI222_X1 U9249 ( .A1(P2_U3151), .A2(n7455), .B1(n8605), .B2(n7456), .C1(
        n9427), .C2(n4627), .ZN(P2_U3284) );
  INV_X1 U9250 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7457) );
  INV_X1 U9251 ( .A(n7674), .ZN(n7667) );
  OAI222_X1 U9252 ( .A1(n10118), .A2(n7457), .B1(n10121), .B2(n7456), .C1(
        n4410), .C2(n7667), .ZN(P1_U3344) );
  INV_X1 U9253 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10541) );
  INV_X1 U9254 ( .A(n7766), .ZN(n7852) );
  NAND2_X1 U9255 ( .A1(n7852), .A2(P2_U3893), .ZN(n7458) );
  OAI21_X1 U9256 ( .B1(P2_U3893), .B2(n10541), .A(n7458), .ZN(P2_U3491) );
  INV_X1 U9257 ( .A(n7459), .ZN(n7463) );
  OAI21_X1 U9258 ( .B1(n7513), .B2(n7461), .A(n7460), .ZN(n7462) );
  NAND3_X1 U9259 ( .A1(n7463), .A2(n8980), .A3(n7462), .ZN(n7477) );
  INV_X1 U9260 ( .A(n9020), .ZN(n8578) );
  OAI21_X1 U9261 ( .B1(n7466), .B2(n7465), .A(n7464), .ZN(n7467) );
  AOI22_X1 U9262 ( .A1(n8988), .A2(P2_ADDR_REG_4__SCAN_IN), .B1(n8578), .B2(
        n7467), .ZN(n7475) );
  NAND2_X1 U9263 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7968) );
  INV_X1 U9264 ( .A(n7468), .ZN(n7473) );
  INV_X1 U9265 ( .A(n7469), .ZN(n7471) );
  NOR3_X1 U9266 ( .A1(n4529), .A2(n7471), .A3(n7470), .ZN(n7472) );
  OAI21_X1 U9267 ( .B1(n7473), .B2(n7472), .A(n9000), .ZN(n7474) );
  AND3_X1 U9268 ( .A1(n7475), .A2(n7968), .A3(n7474), .ZN(n7476) );
  OAI211_X1 U9269 ( .C1(n8969), .C2(n7478), .A(n7477), .B(n7476), .ZN(P2_U3186) );
  INV_X1 U9270 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7480) );
  OAI222_X1 U9271 ( .A1(n9427), .A2(n7480), .B1(n8605), .B2(n7481), .C1(n7479), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U9272 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7482) );
  INV_X1 U9273 ( .A(n7784), .ZN(n7672) );
  OAI222_X1 U9274 ( .A1(n10118), .A2(n7482), .B1(n10121), .B2(n7481), .C1(
        n7672), .C2(n4410), .ZN(P1_U3343) );
  INV_X1 U9275 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n8334) );
  OAI22_X1 U9276 ( .A1(n7485), .A2(n7484), .B1(n7483), .B2(n8334), .ZN(n7600)
         );
  XNOR2_X1 U9277 ( .A(n7491), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7601) );
  NOR2_X1 U9278 ( .A1(n7491), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9682) );
  XNOR2_X1 U9279 ( .A(n9690), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n9681) );
  XNOR2_X1 U9280 ( .A(n7674), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7668) );
  XNOR2_X1 U9281 ( .A(n7669), .B(n7668), .ZN(n7499) );
  INV_X1 U9282 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7486) );
  NAND2_X1 U9283 ( .A1(n4410), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8484) );
  OAI21_X1 U9284 ( .B1(n9786), .B2(n7486), .A(n8484), .ZN(n7487) );
  AOI21_X1 U9285 ( .B1(n9777), .B2(n7674), .A(n7487), .ZN(n7498) );
  NAND2_X1 U9286 ( .A1(n7488), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7489) );
  NAND2_X1 U9287 ( .A1(n7490), .A2(n7489), .ZN(n7607) );
  XNOR2_X1 U9288 ( .A(n7491), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7608) );
  OR2_X1 U9289 ( .A1(n7607), .A2(n7608), .ZN(n7605) );
  OR2_X1 U9290 ( .A1(n7491), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U9291 ( .A1(n7605), .A2(n7492), .ZN(n9687) );
  MUX2_X1 U9292 ( .A(n7493), .B(P1_REG2_REG_10__SCAN_IN), .S(n9690), .Z(n9686)
         );
  OR2_X1 U9293 ( .A1(n9687), .A2(n9686), .ZN(n9688) );
  NAND2_X1 U9294 ( .A1(n9690), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U9295 ( .A1(n9688), .A2(n7494), .ZN(n7496) );
  INV_X1 U9296 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8366) );
  XNOR2_X1 U9297 ( .A(n7674), .B(n8366), .ZN(n7495) );
  NAND2_X1 U9298 ( .A1(n7496), .A2(n7495), .ZN(n7676) );
  OAI211_X1 U9299 ( .C1(n7496), .C2(n7495), .A(n7676), .B(n9773), .ZN(n7497)
         );
  OAI211_X1 U9300 ( .C1(n7499), .C2(n9743), .A(n7498), .B(n7497), .ZN(P1_U3254) );
  XOR2_X1 U9301 ( .A(n7501), .B(n7500), .Z(n7510) );
  XNOR2_X1 U9302 ( .A(n7502), .B(n4666), .ZN(n7503) );
  OAI22_X1 U9303 ( .A1(n9020), .A2(n7503), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10331), .ZN(n7509) );
  INV_X1 U9304 ( .A(n9000), .ZN(n8974) );
  INV_X1 U9305 ( .A(n7504), .ZN(n7505) );
  AOI21_X1 U9306 ( .B1(n10256), .B2(n7506), .A(n7505), .ZN(n7507) );
  INV_X1 U9307 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10271) );
  OAI22_X1 U9308 ( .A1(n8974), .A2(n7507), .B1(n10271), .B2(n9014), .ZN(n7508)
         );
  AOI211_X1 U9309 ( .C1(n8980), .C2(n7510), .A(n7509), .B(n7508), .ZN(n7511)
         );
  OAI21_X1 U9310 ( .B1(n4639), .B2(n8969), .A(n7511), .ZN(P2_U3183) );
  AOI21_X1 U9311 ( .B1(n7515), .B2(n7514), .A(n7513), .ZN(n7526) );
  INV_X1 U9312 ( .A(n8969), .ZN(n9011) );
  INV_X1 U9313 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7832) );
  XNOR2_X1 U9314 ( .A(n7516), .B(n7832), .ZN(n7517) );
  OAI22_X1 U9315 ( .A1(n9020), .A2(n7517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7896), .ZN(n7523) );
  AOI21_X1 U9316 ( .B1(n7519), .B2(n7518), .A(n4529), .ZN(n7521) );
  INV_X1 U9317 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7520) );
  OAI22_X1 U9318 ( .A1(n8974), .A2(n7521), .B1(n9014), .B2(n7520), .ZN(n7522)
         );
  AOI211_X1 U9319 ( .C1(n7524), .C2(n9011), .A(n7523), .B(n7522), .ZN(n7525)
         );
  OAI21_X1 U9320 ( .B1(n7526), .B2(n9006), .A(n7525), .ZN(P2_U3185) );
  XNOR2_X1 U9321 ( .A(n7528), .B(n7527), .ZN(n7539) );
  XNOR2_X1 U9322 ( .A(n7529), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7537) );
  AND2_X1 U9323 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8022) );
  AOI21_X1 U9324 ( .B1(n8988), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8022), .ZN(
        n7534) );
  NAND2_X1 U9325 ( .A1(n7530), .A2(n10260), .ZN(n7531) );
  NAND2_X1 U9326 ( .A1(n7634), .A2(n7531), .ZN(n7532) );
  NAND2_X1 U9327 ( .A1(n9000), .A2(n7532), .ZN(n7533) );
  OAI211_X1 U9328 ( .C1(n8969), .C2(n7535), .A(n7534), .B(n7533), .ZN(n7536)
         );
  AOI21_X1 U9329 ( .B1(n8578), .B2(n7537), .A(n7536), .ZN(n7538) );
  OAI21_X1 U9330 ( .B1(n7539), .B2(n9006), .A(n7538), .ZN(P2_U3187) );
  OAI21_X1 U9331 ( .B1(n10117), .B2(P1_REG2_REG_0__SCAN_IN), .A(n7564), .ZN(
        n7566) );
  AOI21_X1 U9332 ( .B1(n7540), .B2(n10117), .A(n7566), .ZN(n7541) );
  MUX2_X1 U9333 ( .A(n7566), .B(n7541), .S(n7565), .Z(n7546) );
  INV_X1 U9334 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7543) );
  OAI22_X1 U9335 ( .A1(n9786), .A2(n7543), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7542), .ZN(n7545) );
  NOR3_X1 U9336 ( .A1(n9743), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n7565), .ZN(
        n7544) );
  AOI211_X1 U9337 ( .C1(n7547), .C2(n7546), .A(n7545), .B(n7544), .ZN(n7548)
         );
  INV_X1 U9338 ( .A(n7548), .ZN(P1_U3243) );
  INV_X1 U9339 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7549) );
  NAND2_X1 U9340 ( .A1(n4410), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7798) );
  OAI21_X1 U9341 ( .B1(n9786), .B2(n7549), .A(n7798), .ZN(n7560) );
  OAI21_X1 U9342 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(n7558) );
  INV_X1 U9343 ( .A(n7553), .ZN(n9660) );
  NAND3_X1 U9344 ( .A1(n9643), .A2(n7555), .A3(n7554), .ZN(n7556) );
  NAND3_X1 U9345 ( .A1(n9779), .A2(n9660), .A3(n7556), .ZN(n7557) );
  OAI21_X1 U9346 ( .B1(n7558), .B2(n9775), .A(n7557), .ZN(n7559) );
  AOI211_X1 U9347 ( .C1(n7561), .C2(n9777), .A(n7560), .B(n7559), .ZN(n7570)
         );
  XNOR2_X1 U9348 ( .A(n7563), .B(n7562), .ZN(n7663) );
  NAND3_X1 U9349 ( .A1(n7663), .A2(n7564), .A3(n10117), .ZN(n7569) );
  AOI22_X1 U9350 ( .A1(n7567), .A2(n9634), .B1(n7566), .B2(n7565), .ZN(n7568)
         );
  NAND3_X1 U9351 ( .A1(n7569), .A2(P1_U3973), .A3(n7568), .ZN(n7583) );
  NAND2_X1 U9352 ( .A1(n7570), .A2(n7583), .ZN(P1_U3247) );
  OAI22_X1 U9353 ( .A1(n9786), .A2(n10132), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6262), .ZN(n7581) );
  OAI21_X1 U9354 ( .B1(n7573), .B2(n7572), .A(n7571), .ZN(n7579) );
  INV_X1 U9355 ( .A(n7574), .ZN(n7575) );
  XNOR2_X1 U9356 ( .A(n7576), .B(n7575), .ZN(n7577) );
  NAND2_X1 U9357 ( .A1(n9779), .A2(n7577), .ZN(n7578) );
  OAI21_X1 U9358 ( .B1(n9775), .B2(n7579), .A(n7578), .ZN(n7580) );
  AOI211_X1 U9359 ( .C1(n7582), .C2(n9777), .A(n7581), .B(n7580), .ZN(n7584)
         );
  NAND2_X1 U9360 ( .A1(n7584), .A2(n7583), .ZN(P1_U3245) );
  XNOR2_X1 U9361 ( .A(n7586), .B(n7585), .ZN(n7599) );
  INV_X1 U9362 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10563) );
  OAI21_X1 U9363 ( .B1(n7589), .B2(n7588), .A(n7587), .ZN(n7590) );
  AOI22_X1 U9364 ( .A1(n8988), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8578), .B2(
        n7590), .ZN(n7595) );
  NAND2_X1 U9365 ( .A1(n9000), .A2(n7593), .ZN(n7594) );
  OAI211_X1 U9366 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10563), .A(n7595), .B(
        n7594), .ZN(n7596) );
  AOI21_X1 U9367 ( .B1(n7597), .B2(n9011), .A(n7596), .ZN(n7598) );
  OAI21_X1 U9368 ( .B1(n9006), .B2(n7599), .A(n7598), .ZN(P2_U3184) );
  AOI21_X1 U9369 ( .B1(n7601), .B2(n7600), .A(n9683), .ZN(n7612) );
  NOR2_X1 U9370 ( .A1(n7602), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8197) );
  INV_X1 U9371 ( .A(n9777), .ZN(n9766) );
  NOR2_X1 U9372 ( .A1(n9766), .A2(n7603), .ZN(n7604) );
  AOI211_X1 U9373 ( .C1(n9762), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n8197), .B(
        n7604), .ZN(n7611) );
  INV_X1 U9374 ( .A(n7605), .ZN(n7606) );
  AOI21_X1 U9375 ( .B1(n7608), .B2(n7607), .A(n7606), .ZN(n7609) );
  OR2_X1 U9376 ( .A1(n7609), .A2(n9775), .ZN(n7610) );
  OAI211_X1 U9377 ( .C1(n7612), .C2(n9743), .A(n7611), .B(n7610), .ZN(P1_U3252) );
  MUX2_X1 U9378 ( .A(n6334), .B(P1_REG1_REG_7__SCAN_IN), .S(n7613), .Z(n7616)
         );
  INV_X1 U9379 ( .A(n7614), .ZN(n7615) );
  NAND2_X1 U9380 ( .A1(n7616), .A2(n7615), .ZN(n7617) );
  OAI21_X1 U9381 ( .B1(n9671), .B2(n7617), .A(n9779), .ZN(n7625) );
  AND2_X1 U9382 ( .A1(n4410), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7934) );
  NOR2_X1 U9383 ( .A1(n9766), .A2(n7618), .ZN(n7619) );
  AOI211_X1 U9384 ( .C1(n9762), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7934), .B(
        n7619), .ZN(n7624) );
  OAI211_X1 U9385 ( .C1(n7622), .C2(n7621), .A(n9773), .B(n7620), .ZN(n7623)
         );
  OAI211_X1 U9386 ( .C1(n7626), .C2(n7625), .A(n7624), .B(n7623), .ZN(P1_U3250) );
  AOI21_X1 U9387 ( .B1(n7628), .B2(n7627), .A(n7726), .ZN(n7643) );
  OAI21_X1 U9388 ( .B1(n7631), .B2(n7630), .A(n7629), .ZN(n7641) );
  AND2_X1 U9389 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8120) );
  AOI21_X1 U9390 ( .B1(n8988), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8120), .ZN(
        n7638) );
  AND3_X1 U9391 ( .A1(n7634), .A2(n7633), .A3(n7632), .ZN(n7635) );
  OAI21_X1 U9392 ( .B1(n7636), .B2(n7635), .A(n9000), .ZN(n7637) );
  OAI211_X1 U9393 ( .C1(n8969), .C2(n7639), .A(n7638), .B(n7637), .ZN(n7640)
         );
  AOI21_X1 U9394 ( .B1(n8578), .B2(n7641), .A(n7640), .ZN(n7642) );
  OAI21_X1 U9395 ( .B1(n7643), .B2(n9006), .A(n7642), .ZN(P2_U3188) );
  INV_X1 U9396 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10475) );
  INV_X1 U9397 ( .A(n7644), .ZN(n7646) );
  INV_X1 U9398 ( .A(n9707), .ZN(n7645) );
  OAI222_X1 U9399 ( .A1(n10118), .A2(n10475), .B1(n10121), .B2(n7646), .C1(
        n7645), .C2(n4410), .ZN(P1_U3342) );
  INV_X1 U9400 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7647) );
  OAI222_X1 U9401 ( .A1(n9427), .A2(n7647), .B1(n8605), .B2(n7646), .C1(n8919), 
        .C2(P2_U3151), .ZN(P2_U3282) );
  NOR2_X1 U9402 ( .A1(n9919), .A2(n6793), .ZN(n8232) );
  INV_X1 U9403 ( .A(n7648), .ZN(n8235) );
  AOI21_X1 U9404 ( .B1(n10215), .B2(n9917), .A(n8235), .ZN(n7649) );
  AOI211_X1 U9405 ( .C1(n7650), .C2(n8231), .A(n8232), .B(n7649), .ZN(n10185)
         );
  NAND2_X1 U9406 ( .A1(n10222), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7651) );
  OAI21_X1 U9407 ( .B1(n10185), .B2(n10222), .A(n7651), .ZN(P1_U3522) );
  INV_X1 U9408 ( .A(n7689), .ZN(n7654) );
  AOI21_X1 U9409 ( .B1(n7655), .B2(n7652), .A(n7654), .ZN(n7660) );
  AOI22_X1 U9410 ( .A1(n7062), .A2(n9576), .B1(n9606), .B2(n9624), .ZN(n7659)
         );
  OR2_X1 U9411 ( .A1(n7657), .A2(n7656), .ZN(n7691) );
  AOI22_X1 U9412 ( .A1(n9600), .A2(n6273), .B1(n7691), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7658) );
  OAI211_X1 U9413 ( .C1(n7660), .C2(n9578), .A(n7659), .B(n7658), .ZN(P1_U3222) );
  AOI22_X1 U9414 ( .A1(n8231), .A2(n9576), .B1(n9600), .B2(n6792), .ZN(n7662)
         );
  NAND2_X1 U9415 ( .A1(n7691), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7661) );
  OAI211_X1 U9416 ( .C1(n7663), .C2(n9578), .A(n7662), .B(n7661), .ZN(P1_U3232) );
  OAI222_X1 U9417 ( .A1(n10118), .A2(n7664), .B1(n10121), .B2(n7665), .C1(
        n7991), .C2(n4410), .ZN(P1_U3341) );
  INV_X1 U9418 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7666) );
  OAI222_X1 U9419 ( .A1(n9427), .A2(n7666), .B1(n8605), .B2(n7665), .C1(n8940), 
        .C2(P2_U3151), .ZN(P2_U3281) );
  XNOR2_X1 U9420 ( .A(n7784), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7671) );
  OAI22_X1 U9421 ( .A1(n7669), .A2(n7668), .B1(n10468), .B2(n7667), .ZN(n7670)
         );
  NOR2_X1 U9422 ( .A1(n7670), .A2(n7671), .ZN(n9698) );
  AOI21_X1 U9423 ( .B1(n7671), .B2(n7670), .A(n9698), .ZN(n7683) );
  AND2_X1 U9424 ( .A1(n4410), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9488) );
  NOR2_X1 U9425 ( .A1(n9766), .A2(n7672), .ZN(n7673) );
  AOI211_X1 U9426 ( .C1(n9762), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9488), .B(
        n7673), .ZN(n7682) );
  XNOR2_X1 U9427 ( .A(n7784), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U9428 ( .A1(n7674), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9429 ( .A1(n7676), .A2(n7675), .ZN(n7678) );
  OR2_X1 U9430 ( .A1(n7678), .A2(n7679), .ZN(n7786) );
  INV_X1 U9431 ( .A(n7786), .ZN(n7677) );
  AOI21_X1 U9432 ( .B1(n7679), .B2(n7678), .A(n7677), .ZN(n7680) );
  OR2_X1 U9433 ( .A1(n7680), .A2(n9775), .ZN(n7681) );
  OAI211_X1 U9434 ( .C1(n7683), .C2(n9743), .A(n7682), .B(n7681), .ZN(P1_U3255) );
  INV_X1 U9435 ( .A(n7684), .ZN(n7685) );
  NOR2_X1 U9436 ( .A1(n7686), .A2(n7685), .ZN(n7690) );
  INV_X1 U9437 ( .A(n7687), .ZN(n7688) );
  AOI21_X1 U9438 ( .B1(n7690), .B2(n7689), .A(n7688), .ZN(n7694) );
  AOI22_X1 U9439 ( .A1(n8280), .A2(n9576), .B1(n9606), .B2(n6792), .ZN(n7693)
         );
  AOI22_X1 U9440 ( .A1(n9600), .A2(n10161), .B1(n7691), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7692) );
  OAI211_X1 U9441 ( .C1(n7694), .C2(n9578), .A(n7693), .B(n7692), .ZN(P1_U3237) );
  OAI21_X1 U9442 ( .B1(n9247), .B2(n10250), .A(n7736), .ZN(n7696) );
  INV_X1 U9443 ( .A(n9203), .ZN(n9147) );
  NOR2_X1 U9444 ( .A1(n7756), .A2(n9147), .ZN(n7741) );
  INV_X1 U9445 ( .A(n7741), .ZN(n7695) );
  OAI211_X1 U9446 ( .C1(n10241), .C2(n7745), .A(n7696), .B(n7695), .ZN(n7698)
         );
  NAND2_X1 U9447 ( .A1(n10266), .A2(n7698), .ZN(n7697) );
  OAI21_X1 U9448 ( .B1(n10266), .B2(n6984), .A(n7697), .ZN(P2_U3459) );
  NAND2_X1 U9449 ( .A1(n10254), .A2(n7698), .ZN(n7699) );
  OAI21_X1 U9450 ( .B1(n10254), .B2(n5306), .A(n7699), .ZN(P2_U3390) );
  NAND2_X1 U9451 ( .A1(n7703), .A2(n10249), .ZN(n7700) );
  INV_X1 U9452 ( .A(n8886), .ZN(n8902) );
  INV_X1 U9453 ( .A(n7701), .ZN(n7702) );
  NAND2_X1 U9454 ( .A1(n7703), .A2(n7702), .ZN(n7707) );
  INV_X1 U9455 ( .A(n7704), .ZN(n7712) );
  NAND2_X1 U9456 ( .A1(n7705), .A2(n7712), .ZN(n7706) );
  NOR2_X1 U9457 ( .A1(n7708), .A2(n7737), .ZN(n7764) );
  AOI22_X1 U9458 ( .A1(n8855), .A2(n7736), .B1(n8894), .B2(n9242), .ZN(n7722)
         );
  NAND2_X1 U9459 ( .A1(n7710), .A2(n7709), .ZN(n7714) );
  AOI21_X1 U9460 ( .B1(n7717), .B2(n7712), .A(n7711), .ZN(n7713) );
  NAND2_X1 U9461 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  NAND2_X1 U9462 ( .A1(n7715), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7719) );
  NAND2_X1 U9463 ( .A1(n7717), .A2(n7716), .ZN(n7718) );
  NAND2_X1 U9464 ( .A1(n7719), .A2(n7718), .ZN(n7895) );
  OR2_X1 U9465 ( .A1(n7895), .A2(n7720), .ZN(n7806) );
  NAND2_X1 U9466 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n7806), .ZN(n7721) );
  OAI211_X1 U9467 ( .C1(n8902), .C2(n7745), .A(n7722), .B(n7721), .ZN(P2_U3172) );
  INV_X1 U9468 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8088) );
  XNOR2_X1 U9469 ( .A(n7723), .B(n8088), .ZN(n7735) );
  NOR3_X1 U9470 ( .A1(n7726), .A2(n7725), .A3(n7724), .ZN(n7727) );
  OAI21_X1 U9471 ( .B1(n4928), .B2(n7727), .A(n8980), .ZN(n7734) );
  OAI21_X1 U9472 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n7728), .A(n7870), .ZN(
        n7732) );
  NOR2_X1 U9473 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5423), .ZN(n8258) );
  AOI21_X1 U9474 ( .B1(n8988), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8258), .ZN(
        n7729) );
  OAI21_X1 U9475 ( .B1(n7730), .B2(n8969), .A(n7729), .ZN(n7731) );
  AOI21_X1 U9476 ( .B1(n7732), .B2(n9000), .A(n7731), .ZN(n7733) );
  OAI211_X1 U9477 ( .C1(n7735), .C2(n9020), .A(n7734), .B(n7733), .ZN(P2_U3189) );
  INV_X1 U9478 ( .A(n7736), .ZN(n7739) );
  INV_X1 U9479 ( .A(n7737), .ZN(n7738) );
  NOR3_X1 U9480 ( .A1(n7739), .A2(n7738), .A3(n10249), .ZN(n7740) );
  AOI211_X1 U9481 ( .C1(n9250), .C2(P2_REG3_REG_0__SCAN_IN), .A(n7741), .B(
        n7740), .ZN(n7742) );
  MUX2_X1 U9482 ( .A(n7743), .B(n7742), .S(n9253), .Z(n7744) );
  OAI21_X1 U9483 ( .B1(n9153), .B2(n7745), .A(n7744), .ZN(P2_U3233) );
  XNOR2_X1 U9484 ( .A(n8465), .B(n7746), .ZN(n7747) );
  NAND2_X1 U9485 ( .A1(n7750), .A2(n7749), .ZN(n7752) );
  NAND2_X2 U9486 ( .A1(n7752), .A2(n7751), .ZN(n7809) );
  OR2_X1 U9487 ( .A1(n7809), .A2(n7753), .ZN(n7754) );
  AND2_X1 U9488 ( .A1(n7754), .A2(n7848), .ZN(n7761) );
  XNOR2_X1 U9489 ( .A(n7809), .B(n7857), .ZN(n7757) );
  INV_X1 U9490 ( .A(n7757), .ZN(n7755) );
  INV_X1 U9491 ( .A(n7761), .ZN(n7758) );
  INV_X1 U9492 ( .A(n7811), .ZN(n7759) );
  AOI21_X1 U9493 ( .B1(n7761), .B2(n7760), .A(n7759), .ZN(n7769) );
  INV_X1 U9494 ( .A(n7762), .ZN(n7763) );
  AOI22_X1 U9495 ( .A1(n8886), .A2(n7857), .B1(n8894), .B2(n8912), .ZN(n7765)
         );
  OAI21_X1 U9496 ( .B1(n7766), .B2(n8896), .A(n7765), .ZN(n7767) );
  AOI21_X1 U9497 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7806), .A(n7767), .ZN(
        n7768) );
  OAI21_X1 U9498 ( .B1(n8889), .B2(n7769), .A(n7768), .ZN(P2_U3162) );
  OAI21_X1 U9499 ( .B1(n7772), .B2(n7771), .A(n7770), .ZN(n7776) );
  MUX2_X1 U9500 ( .A(n9603), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7774) );
  AOI22_X1 U9501 ( .A1(n8412), .A2(n9576), .B1(n9606), .B2(n6273), .ZN(n7773)
         );
  OAI211_X1 U9502 ( .C1(n8006), .C2(n9586), .A(n7774), .B(n7773), .ZN(n7775)
         );
  AOI21_X1 U9503 ( .B1(n7776), .B2(n9598), .A(n7775), .ZN(n7777) );
  INV_X1 U9504 ( .A(n7777), .ZN(P1_U3218) );
  INV_X1 U9505 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7779) );
  INV_X1 U9506 ( .A(n7778), .ZN(n7780) );
  OAI222_X1 U9507 ( .A1(n10118), .A2(n7779), .B1(n10121), .B2(n7780), .C1(
        n4410), .C2(n7995), .ZN(P1_U3340) );
  INV_X1 U9508 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7781) );
  OAI222_X1 U9509 ( .A1(n9427), .A2(n7781), .B1(n8605), .B2(n7780), .C1(
        P2_U3151), .C2(n4877), .ZN(P2_U3280) );
  NOR2_X1 U9510 ( .A1(n7784), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9697) );
  XNOR2_X1 U9511 ( .A(n9707), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9696) );
  AOI21_X1 U9512 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n9707), .A(n9695), .ZN(
        n7988) );
  XNOR2_X1 U9513 ( .A(n7991), .B(n10361), .ZN(n7987) );
  XNOR2_X1 U9514 ( .A(n7988), .B(n7987), .ZN(n7792) );
  NOR2_X1 U9515 ( .A1(n7782), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9446) );
  NOR2_X1 U9516 ( .A1(n9766), .A2(n7991), .ZN(n7783) );
  AOI211_X1 U9517 ( .C1(n9762), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9446), .B(
        n7783), .ZN(n7791) );
  OR2_X1 U9518 ( .A1(n7784), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7785) );
  NAND2_X1 U9519 ( .A1(n7786), .A2(n7785), .ZN(n9704) );
  XNOR2_X1 U9520 ( .A(n9707), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U9521 ( .A1(n9707), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U9522 ( .A1(n9705), .A2(n7787), .ZN(n7789) );
  XNOR2_X1 U9523 ( .A(n7991), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U9524 ( .A1(n7789), .A2(n7788), .ZN(n7994) );
  OAI211_X1 U9525 ( .C1(n7789), .C2(n7788), .A(n7994), .B(n9773), .ZN(n7790)
         );
  OAI211_X1 U9526 ( .C1(n7792), .C2(n9743), .A(n7791), .B(n7790), .ZN(P1_U3257) );
  INV_X1 U9527 ( .A(n7793), .ZN(n7797) );
  AOI21_X1 U9528 ( .B1(n7770), .B2(n7795), .A(n7794), .ZN(n7796) );
  NOR3_X1 U9529 ( .A1(n7797), .A2(n7796), .A3(n9578), .ZN(n7803) );
  AOI22_X1 U9530 ( .A1(n9606), .A2(n10161), .B1(n9600), .B2(n10159), .ZN(n7801) );
  OAI21_X1 U9531 ( .B1(n9609), .B2(n10202), .A(n7798), .ZN(n7799) );
  INV_X1 U9532 ( .A(n7799), .ZN(n7800) );
  OAI211_X1 U9533 ( .C1(n9603), .C2(n10164), .A(n7801), .B(n7800), .ZN(n7802)
         );
  OR2_X1 U9534 ( .A1(n7803), .A2(n7802), .ZN(P1_U3230) );
  INV_X1 U9535 ( .A(n7804), .ZN(n7885) );
  AOI22_X1 U9536 ( .A1(n9731), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10110), .ZN(n7805) );
  OAI21_X1 U9537 ( .B1(n7885), .B2(n10121), .A(n7805), .ZN(P1_U3339) );
  INV_X1 U9538 ( .A(n7806), .ZN(n7817) );
  OAI22_X1 U9539 ( .A1(n8902), .A2(n7807), .B1(n8883), .B2(n7913), .ZN(n7808)
         );
  AOI21_X1 U9540 ( .B1(n8880), .B2(n9242), .A(n7808), .ZN(n7816) );
  XNOR2_X1 U9541 ( .A(n7888), .B(n8912), .ZN(n7813) );
  NAND2_X1 U9542 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  OAI21_X1 U9543 ( .B1(n7813), .B2(n7812), .A(n7890), .ZN(n7814) );
  NAND2_X1 U9544 ( .A1(n8855), .A2(n7814), .ZN(n7815) );
  OAI211_X1 U9545 ( .C1(n7817), .C2(n10563), .A(n7816), .B(n7815), .ZN(
        P2_U3177) );
  INV_X1 U9546 ( .A(n5955), .ZN(n7818) );
  NAND2_X1 U9547 ( .A1(n9235), .A2(n7818), .ZN(n9236) );
  NAND2_X1 U9548 ( .A1(n9236), .A2(n7819), .ZN(n7821) );
  INV_X1 U9549 ( .A(n7827), .ZN(n7820) );
  NAND2_X1 U9550 ( .A1(n7821), .A2(n7820), .ZN(n7905) );
  OR2_X1 U9551 ( .A1(n7821), .A2(n7820), .ZN(n7822) );
  NAND2_X1 U9552 ( .A1(n7905), .A2(n7822), .ZN(n7860) );
  INV_X1 U9553 ( .A(n7860), .ZN(n7835) );
  NAND2_X1 U9554 ( .A1(n7824), .A2(n7823), .ZN(n9239) );
  NAND2_X1 U9555 ( .A1(n9239), .A2(n5955), .ZN(n7826) );
  NAND2_X1 U9556 ( .A1(n7826), .A2(n7825), .ZN(n7828) );
  XNOR2_X1 U9557 ( .A(n7828), .B(n7827), .ZN(n7831) );
  NAND2_X1 U9558 ( .A1(n8912), .A2(n9241), .ZN(n7829) );
  OAI21_X1 U9559 ( .B1(n8020), .B2(n9147), .A(n7829), .ZN(n7830) );
  AOI21_X1 U9560 ( .B1(n7831), .B2(n9247), .A(n7830), .ZN(n7861) );
  MUX2_X1 U9561 ( .A(n7861), .B(n7832), .S(n9213), .Z(n7834) );
  AOI22_X1 U9562 ( .A1(n9230), .A2(n7976), .B1(n9250), .B2(n7896), .ZN(n7833)
         );
  OAI211_X1 U9563 ( .C1(n7835), .C2(n9233), .A(n7834), .B(n7833), .ZN(P2_U3230) );
  XNOR2_X1 U9564 ( .A(n7837), .B(n7836), .ZN(n8281) );
  INV_X1 U9565 ( .A(n10211), .ZN(n10201) );
  OAI21_X1 U9566 ( .B1(n7840), .B2(n7839), .A(n7838), .ZN(n7841) );
  AOI222_X1 U9567 ( .A1(n10163), .A2(n7841), .B1(n10161), .B2(n10158), .C1(
        n6792), .C2(n10160), .ZN(n8284) );
  OAI211_X1 U9568 ( .C1(n7842), .C2(n8147), .A(n10174), .B(n8410), .ZN(n8276)
         );
  OAI211_X1 U9569 ( .C1(n7842), .C2(n10201), .A(n8284), .B(n8276), .ZN(n7843)
         );
  AOI21_X1 U9570 ( .B1(n8281), .B2(n10206), .A(n7843), .ZN(n10193) );
  NAND2_X1 U9571 ( .A1(n10222), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7844) );
  OAI21_X1 U9572 ( .B1(n10193), .B2(n10222), .A(n7844), .ZN(P1_U3524) );
  INV_X1 U9573 ( .A(n7845), .ZN(n7846) );
  AOI21_X1 U9574 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(n10226) );
  OAI22_X1 U9575 ( .A1(n10226), .A2(n9252), .B1(n10331), .B2(n9207), .ZN(n7856) );
  XNOR2_X1 U9576 ( .A(n7850), .B(n7849), .ZN(n7855) );
  INV_X1 U9577 ( .A(n10226), .ZN(n7851) );
  NAND2_X1 U9578 ( .A1(n7851), .A2(n6895), .ZN(n7854) );
  AOI22_X1 U9579 ( .A1(n7852), .A2(n9241), .B1(n9203), .B2(n8912), .ZN(n7853)
         );
  OAI211_X1 U9580 ( .C1(n7855), .C2(n9142), .A(n7854), .B(n7853), .ZN(n10227)
         );
  OAI21_X1 U9581 ( .B1(n7856), .B2(n10227), .A(n9253), .ZN(n7859) );
  NAND2_X1 U9582 ( .A1(n9230), .A2(n7857), .ZN(n7858) );
  OAI211_X1 U9583 ( .C1(n4666), .C2(n9253), .A(n7859), .B(n7858), .ZN(P2_U3232) );
  NAND2_X1 U9584 ( .A1(n7860), .A2(n10250), .ZN(n7862) );
  NAND2_X1 U9585 ( .A1(n7862), .A2(n7861), .ZN(n7974) );
  OAI22_X1 U9586 ( .A1(n7887), .A2(n9372), .B1(n10254), .B2(n5311), .ZN(n7863)
         );
  AOI21_X1 U9587 ( .B1(n10254), .B2(n7974), .A(n7863), .ZN(n7864) );
  INV_X1 U9588 ( .A(n7864), .ZN(P2_U3399) );
  OAI21_X1 U9589 ( .B1(n7867), .B2(n7866), .A(n7865), .ZN(n7883) );
  AND3_X1 U9590 ( .A1(n7870), .A2(n7869), .A3(n7868), .ZN(n7871) );
  OAI21_X1 U9591 ( .B1(n7872), .B2(n7871), .A(n9000), .ZN(n7874) );
  AND2_X1 U9592 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8399) );
  AOI21_X1 U9593 ( .B1(n8988), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8399), .ZN(
        n7873) );
  OAI211_X1 U9594 ( .C1(n8969), .C2(n7875), .A(n7874), .B(n7873), .ZN(n7882)
         );
  INV_X1 U9595 ( .A(n7946), .ZN(n7880) );
  NAND3_X1 U9596 ( .A1(n7878), .A2(n7877), .A3(n7876), .ZN(n7879) );
  AOI21_X1 U9597 ( .B1(n7880), .B2(n7879), .A(n9006), .ZN(n7881) );
  AOI211_X1 U9598 ( .C1(n8578), .C2(n7883), .A(n7882), .B(n7881), .ZN(n7884)
         );
  INV_X1 U9599 ( .A(n7884), .ZN(P2_U3190) );
  INV_X1 U9600 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7886) );
  OAI222_X1 U9601 ( .A1(n9427), .A2(n7886), .B1(n8605), .B2(n7885), .C1(
        P2_U3151), .C2(n8968), .ZN(P2_U3279) );
  XNOR2_X1 U9602 ( .A(n7809), .B(n7887), .ZN(n7957) );
  NAND2_X1 U9603 ( .A1(n7888), .A2(n7899), .ZN(n7889) );
  INV_X1 U9604 ( .A(n7959), .ZN(n7891) );
  AOI211_X1 U9605 ( .C1(n7893), .C2(n7892), .A(n8889), .B(n7891), .ZN(n7901)
         );
  MUX2_X1 U9606 ( .A(P2_STATE_REG_SCAN_IN), .B(n8862), .S(n7896), .Z(n7898) );
  AOI22_X1 U9607 ( .A1(n8886), .A2(n7976), .B1(n8894), .B2(n5157), .ZN(n7897)
         );
  OAI211_X1 U9608 ( .C1(n7899), .C2(n8896), .A(n7898), .B(n7897), .ZN(n7900)
         );
  OR2_X1 U9609 ( .A1(n7901), .A2(n7900), .ZN(P2_U3158) );
  INV_X1 U9610 ( .A(n7902), .ZN(n7941) );
  AOI22_X1 U9611 ( .A1(n9749), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10110), .ZN(n7903) );
  OAI21_X1 U9612 ( .B1(n7941), .B2(n10121), .A(n7903), .ZN(P1_U3338) );
  NAND3_X1 U9613 ( .A1(n7905), .A2(n7904), .A3(n7919), .ZN(n7907) );
  NAND2_X1 U9614 ( .A1(n7907), .A2(n7906), .ZN(n8078) );
  INV_X1 U9615 ( .A(n7908), .ZN(n7909) );
  NAND2_X1 U9616 ( .A1(n7910), .A2(n7909), .ZN(n7920) );
  XNOR2_X1 U9617 ( .A(n7920), .B(n7911), .ZN(n7912) );
  OAI222_X1 U9618 ( .A1(n9145), .A2(n7913), .B1(n9147), .B2(n8118), .C1(n9142), 
        .C2(n7912), .ZN(n8075) );
  AOI21_X1 U9619 ( .B1(n10250), .B2(n8078), .A(n8075), .ZN(n8063) );
  AOI22_X1 U9620 ( .A1(n9407), .A2(n7960), .B1(n10255), .B2(
        P2_REG0_REG_4__SCAN_IN), .ZN(n7914) );
  OAI21_X1 U9621 ( .B1(n8063), .B2(n10255), .A(n7914), .ZN(P2_U3402) );
  INV_X1 U9622 ( .A(n7906), .ZN(n7916) );
  NOR2_X1 U9623 ( .A1(n7916), .A2(n7915), .ZN(n8055) );
  XNOR2_X1 U9624 ( .A(n8055), .B(n7921), .ZN(n10235) );
  INV_X1 U9625 ( .A(n9252), .ZN(n7917) );
  NAND2_X1 U9626 ( .A1(n9253), .A2(n7917), .ZN(n9034) );
  AOI21_X1 U9627 ( .B1(n7920), .B2(n7919), .A(n7918), .ZN(n7922) );
  XNOR2_X1 U9628 ( .A(n7922), .B(n7921), .ZN(n7924) );
  OAI22_X1 U9629 ( .A1(n8256), .A2(n9147), .B1(n8020), .B2(n9145), .ZN(n7923)
         );
  AOI21_X1 U9630 ( .B1(n7924), .B2(n9247), .A(n7923), .ZN(n7925) );
  OAI21_X1 U9631 ( .B1(n10235), .B2(n9244), .A(n7925), .ZN(n10236) );
  NAND2_X1 U9632 ( .A1(n10236), .A2(n9253), .ZN(n7929) );
  INV_X1 U9633 ( .A(n10238), .ZN(n7926) );
  OAI22_X1 U9634 ( .A1(n9153), .A2(n7926), .B1(n8025), .B2(n9207), .ZN(n7927)
         );
  AOI21_X1 U9635 ( .B1(n9213), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7927), .ZN(
        n7928) );
  OAI211_X1 U9636 ( .C1(n10235), .C2(n9034), .A(n7929), .B(n7928), .ZN(
        P2_U3228) );
  XNOR2_X1 U9637 ( .A(n7932), .B(n7931), .ZN(n7933) );
  XNOR2_X1 U9638 ( .A(n7930), .B(n7933), .ZN(n7938) );
  AOI22_X1 U9639 ( .A1(n9606), .A2(n9621), .B1(n9600), .B2(n9620), .ZN(n7936)
         );
  AOI21_X1 U9640 ( .B1(n9576), .B2(n8246), .A(n7934), .ZN(n7935) );
  OAI211_X1 U9641 ( .C1(n9603), .C2(n8243), .A(n7936), .B(n7935), .ZN(n7937)
         );
  AOI21_X1 U9642 ( .B1(n7938), .B2(n9598), .A(n7937), .ZN(n7939) );
  INV_X1 U9643 ( .A(n7939), .ZN(P1_U3213) );
  OAI222_X1 U9644 ( .A1(n9427), .A2(n7942), .B1(n8605), .B2(n7941), .C1(
        P2_U3151), .C2(n7940), .ZN(P2_U3278) );
  XOR2_X1 U9645 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7943), .Z(n7956) );
  NOR3_X1 U9646 ( .A1(n7946), .A2(n7945), .A3(n7944), .ZN(n7947) );
  OAI21_X1 U9647 ( .B1(n4921), .B2(n7947), .A(n8980), .ZN(n7955) );
  OAI21_X1 U9648 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7949), .A(n7948), .ZN(
        n7953) );
  NOR2_X1 U9649 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5457), .ZN(n8559) );
  AOI21_X1 U9650 ( .B1(n8988), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8559), .ZN(
        n7950) );
  OAI21_X1 U9651 ( .B1(n7951), .B2(n8969), .A(n7950), .ZN(n7952) );
  AOI21_X1 U9652 ( .B1(n7953), .B2(n9000), .A(n7952), .ZN(n7954) );
  OAI211_X1 U9653 ( .C1(n7956), .C2(n9020), .A(n7955), .B(n7954), .ZN(P2_U3191) );
  NAND2_X1 U9654 ( .A1(n7957), .A2(n9240), .ZN(n7958) );
  NAND2_X1 U9655 ( .A1(n7959), .A2(n7958), .ZN(n7967) );
  INV_X2 U9656 ( .A(n8684), .ZN(n8680) );
  XNOR2_X1 U9657 ( .A(n8680), .B(n7960), .ZN(n7961) );
  NAND2_X1 U9658 ( .A1(n7961), .A2(n8020), .ZN(n8014) );
  INV_X1 U9659 ( .A(n7961), .ZN(n7962) );
  NAND2_X1 U9660 ( .A1(n7962), .A2(n5157), .ZN(n7963) );
  NAND2_X1 U9661 ( .A1(n8014), .A2(n7963), .ZN(n7966) );
  INV_X1 U9662 ( .A(n7967), .ZN(n7965) );
  NAND2_X1 U9663 ( .A1(n7965), .A2(n7964), .ZN(n8015) );
  INV_X1 U9664 ( .A(n8015), .ZN(n8013) );
  AOI21_X1 U9665 ( .B1(n7967), .B2(n7966), .A(n8013), .ZN(n7973) );
  INV_X1 U9666 ( .A(n8074), .ZN(n7971) );
  AOI22_X1 U9667 ( .A1(n8880), .A2(n9240), .B1(n8894), .B2(n8911), .ZN(n7969)
         );
  OAI211_X1 U9668 ( .C1(n8902), .C2(n5155), .A(n7969), .B(n7968), .ZN(n7970)
         );
  AOI21_X1 U9669 ( .B1(n7971), .B2(n8899), .A(n7970), .ZN(n7972) );
  OAI21_X1 U9670 ( .B1(n7973), .B2(n8889), .A(n7972), .ZN(P2_U3170) );
  MUX2_X1 U9671 ( .A(n7974), .B(P2_REG1_REG_3__SCAN_IN), .S(n6909), .Z(n7975)
         );
  AOI21_X1 U9672 ( .B1(n9315), .B2(n7976), .A(n7975), .ZN(n7977) );
  INV_X1 U9673 ( .A(n7977), .ZN(P2_U3462) );
  AOI21_X1 U9674 ( .B1(n7793), .B2(n7978), .A(n7979), .ZN(n8026) );
  AND3_X1 U9675 ( .A1(n7793), .A2(n7979), .A3(n7978), .ZN(n8028) );
  NOR2_X1 U9676 ( .A1(n8026), .A2(n8028), .ZN(n7980) );
  XNOR2_X1 U9677 ( .A(n7980), .B(n8029), .ZN(n7985) );
  AOI22_X1 U9678 ( .A1(n9606), .A2(n9622), .B1(n9600), .B2(n9621), .ZN(n7983)
         );
  NAND2_X1 U9679 ( .A1(n4410), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9650) );
  OAI21_X1 U9680 ( .B1(n9609), .B2(n8225), .A(n9650), .ZN(n7981) );
  INV_X1 U9681 ( .A(n7981), .ZN(n7982) );
  OAI211_X1 U9682 ( .C1(n9603), .C2(n8224), .A(n7983), .B(n7982), .ZN(n7984)
         );
  AOI21_X1 U9683 ( .B1(n7985), .B2(n9598), .A(n7984), .ZN(n7986) );
  INV_X1 U9684 ( .A(n7986), .ZN(P1_U3227) );
  OAI22_X1 U9685 ( .A1(n7988), .A2(n7987), .B1(n10361), .B2(n7991), .ZN(n9712)
         );
  XNOR2_X1 U9686 ( .A(n9713), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n7999) );
  NOR2_X1 U9687 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9602), .ZN(n7990) );
  NOR2_X1 U9688 ( .A1(n9766), .A2(n7995), .ZN(n7989) );
  AOI211_X1 U9689 ( .C1(n9762), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7990), .B(
        n7989), .ZN(n7998) );
  INV_X1 U9690 ( .A(n7991), .ZN(n7992) );
  NAND2_X1 U9691 ( .A1(n7992), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U9692 ( .A1(n7994), .A2(n7993), .ZN(n9721) );
  XNOR2_X1 U9693 ( .A(n9721), .B(n7995), .ZN(n7996) );
  NAND2_X1 U9694 ( .A1(n7996), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9723) );
  OAI211_X1 U9695 ( .C1(n7996), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9723), .B(
        n9773), .ZN(n7997) );
  OAI211_X1 U9696 ( .C1(n7999), .C2(n9743), .A(n7998), .B(n7997), .ZN(P1_U3258) );
  XNOR2_X1 U9697 ( .A(n8000), .B(n8002), .ZN(n8220) );
  OAI21_X1 U9698 ( .B1(n10173), .B2(n8225), .A(n10174), .ZN(n8001) );
  NOR2_X1 U9699 ( .A1(n8001), .A2(n8213), .ZN(n8227) );
  XNOR2_X1 U9700 ( .A(n8003), .B(n8002), .ZN(n8004) );
  OAI222_X1 U9701 ( .A1(n9921), .A2(n8006), .B1(n9919), .B2(n8005), .C1(n9917), 
        .C2(n8004), .ZN(n8221) );
  AOI211_X1 U9702 ( .C1(n8220), .C2(n10206), .A(n8227), .B(n8221), .ZN(n8011)
         );
  OAI22_X1 U9703 ( .A1(n10066), .A2(n8225), .B1(n10225), .B2(n7427), .ZN(n8007) );
  INV_X1 U9704 ( .A(n8007), .ZN(n8008) );
  OAI21_X1 U9705 ( .B1(n8011), .B2(n10222), .A(n8008), .ZN(P1_U3527) );
  OAI22_X1 U9706 ( .A1(n10102), .A2(n8225), .B1(n10218), .B2(n6313), .ZN(n8009) );
  INV_X1 U9707 ( .A(n8009), .ZN(n8010) );
  OAI21_X1 U9708 ( .B1(n8011), .B2(n10217), .A(n8010), .ZN(P1_U3468) );
  INV_X1 U9709 ( .A(n8014), .ZN(n8012) );
  XNOR2_X1 U9710 ( .A(n8680), .B(n10238), .ZN(n8113) );
  XNOR2_X1 U9711 ( .A(n8113), .B(n8911), .ZN(n8016) );
  NOR3_X1 U9712 ( .A1(n8013), .A2(n8012), .A3(n8016), .ZN(n8019) );
  NAND2_X1 U9713 ( .A1(n8015), .A2(n8014), .ZN(n8017) );
  NAND2_X1 U9714 ( .A1(n8017), .A2(n8016), .ZN(n8115) );
  INV_X1 U9715 ( .A(n8115), .ZN(n8018) );
  OAI21_X1 U9716 ( .B1(n8019), .B2(n8018), .A(n8855), .ZN(n8024) );
  OAI22_X1 U9717 ( .A1(n8883), .A2(n8256), .B1(n8020), .B2(n8896), .ZN(n8021)
         );
  AOI211_X1 U9718 ( .C1(n10238), .C2(n8886), .A(n8022), .B(n8021), .ZN(n8023)
         );
  OAI211_X1 U9719 ( .C1(n8025), .C2(n8862), .A(n8024), .B(n8023), .ZN(P2_U3167) );
  INV_X1 U9720 ( .A(n8026), .ZN(n8027) );
  OAI21_X1 U9721 ( .B1(n8029), .B2(n8028), .A(n8027), .ZN(n8034) );
  OAI21_X1 U9722 ( .B1(n8032), .B2(n8031), .A(n8030), .ZN(n8033) );
  XNOR2_X1 U9723 ( .A(n8034), .B(n8033), .ZN(n8038) );
  AOI22_X1 U9724 ( .A1(n9606), .A2(n10159), .B1(n9600), .B2(n8210), .ZN(n8036)
         );
  AND2_X1 U9725 ( .A1(n4410), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9667) );
  AOI21_X1 U9726 ( .B1(n9576), .B2(n10210), .A(n9667), .ZN(n8035) );
  OAI211_X1 U9727 ( .C1(n9603), .C2(n8215), .A(n8036), .B(n8035), .ZN(n8037)
         );
  AOI21_X1 U9728 ( .B1(n8038), .B2(n9598), .A(n8037), .ZN(n8039) );
  INV_X1 U9729 ( .A(n8039), .ZN(P1_U3239) );
  INV_X1 U9730 ( .A(n8040), .ZN(n8042) );
  INV_X1 U9731 ( .A(n9769), .ZN(n9765) );
  OAI222_X1 U9732 ( .A1(n10118), .A2(n8041), .B1(n10121), .B2(n8042), .C1(
        n9765), .C2(n4410), .ZN(P1_U3337) );
  OAI222_X1 U9733 ( .A1(P2_U3151), .A2(n9009), .B1(n8605), .B2(n8042), .C1(
        n10441), .C2(n9427), .ZN(P2_U3277) );
  XNOR2_X1 U9734 ( .A(n8043), .B(n4734), .ZN(n8044) );
  NAND2_X1 U9735 ( .A1(n8044), .A2(n9247), .ZN(n8046) );
  AOI22_X1 U9736 ( .A1(n9203), .A2(n8742), .B1(n8909), .B2(n9241), .ZN(n8045)
         );
  AND2_X1 U9737 ( .A1(n8046), .A2(n8045), .ZN(n10253) );
  XNOR2_X1 U9738 ( .A(n8048), .B(n8047), .ZN(n10251) );
  NOR2_X1 U9739 ( .A1(n9253), .A2(n6997), .ZN(n8051) );
  INV_X1 U9740 ( .A(n10248), .ZN(n8049) );
  OAI22_X1 U9741 ( .A1(n9153), .A2(n8049), .B1(n8402), .B2(n9207), .ZN(n8050)
         );
  AOI211_X1 U9742 ( .C1(n10251), .C2(n9155), .A(n8051), .B(n8050), .ZN(n8052)
         );
  OAI21_X1 U9743 ( .B1(n10253), .B2(n9213), .A(n8052), .ZN(P2_U3225) );
  OAI21_X1 U9744 ( .B1(n8055), .B2(n8054), .A(n8053), .ZN(n8056) );
  XNOR2_X1 U9745 ( .A(n8056), .B(n8057), .ZN(n8070) );
  XOR2_X1 U9746 ( .A(n8058), .B(n8057), .Z(n8059) );
  AOI222_X1 U9747 ( .A1(n9247), .A2(n8059), .B1(n8909), .B2(n9203), .C1(n8911), 
        .C2(n9241), .ZN(n8065) );
  OAI21_X1 U9748 ( .B1(n8060), .B2(n8070), .A(n8065), .ZN(n8071) );
  INV_X1 U9749 ( .A(n8071), .ZN(n8062) );
  AOI22_X1 U9750 ( .A1(n9315), .A2(n8121), .B1(n6909), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n8061) );
  OAI21_X1 U9751 ( .B1(n8062), .B2(n6909), .A(n8061), .ZN(P2_U3465) );
  MUX2_X1 U9752 ( .A(n5339), .B(n8063), .S(n10266), .Z(n8064) );
  OAI21_X1 U9753 ( .B1(n5155), .B2(n9298), .A(n8064), .ZN(P2_U3463) );
  MUX2_X1 U9754 ( .A(n8066), .B(n8065), .S(n9253), .Z(n8069) );
  INV_X1 U9755 ( .A(n8124), .ZN(n8067) );
  AOI22_X1 U9756 ( .A1(n9230), .A2(n8121), .B1(n9250), .B2(n8067), .ZN(n8068)
         );
  OAI211_X1 U9757 ( .C1(n8070), .C2(n9233), .A(n8069), .B(n8068), .ZN(P2_U3227) );
  NAND2_X1 U9758 ( .A1(n8071), .A2(n10254), .ZN(n8073) );
  NAND2_X1 U9759 ( .A1(n9407), .A2(n8121), .ZN(n8072) );
  OAI211_X1 U9760 ( .C1(n5405), .C2(n10254), .A(n8073), .B(n8072), .ZN(
        P2_U3408) );
  OAI22_X1 U9761 ( .A1(n9153), .A2(n5155), .B1(n8074), .B2(n9207), .ZN(n8077)
         );
  MUX2_X1 U9762 ( .A(n8075), .B(P2_REG2_REG_4__SCAN_IN), .S(n9213), .Z(n8076)
         );
  AOI211_X1 U9763 ( .C1(n9155), .C2(n8078), .A(n8077), .B(n8076), .ZN(n8079)
         );
  INV_X1 U9764 ( .A(n8079), .ZN(P2_U3229) );
  OR2_X1 U9765 ( .A1(n8080), .A2(n8083), .ZN(n8081) );
  NAND2_X1 U9766 ( .A1(n8082), .A2(n8081), .ZN(n10244) );
  XOR2_X1 U9767 ( .A(n8084), .B(n8083), .Z(n8087) );
  AOI22_X1 U9768 ( .A1(n8908), .A2(n9203), .B1(n9241), .B2(n8910), .ZN(n8085)
         );
  OAI21_X1 U9769 ( .B1(n10244), .B2(n9244), .A(n8085), .ZN(n8086) );
  AOI21_X1 U9770 ( .B1(n8087), .B2(n9247), .A(n8086), .ZN(n10240) );
  MUX2_X1 U9771 ( .A(n8088), .B(n10240), .S(n9253), .Z(n8091) );
  INV_X1 U9772 ( .A(n8262), .ZN(n8089) );
  AOI22_X1 U9773 ( .A1(n9230), .A2(n8259), .B1(n9250), .B2(n8089), .ZN(n8090)
         );
  OAI211_X1 U9774 ( .C1(n10244), .C2(n9034), .A(n8091), .B(n8090), .ZN(
        P2_U3226) );
  XOR2_X1 U9775 ( .A(n8093), .B(n8092), .Z(n8110) );
  INV_X1 U9776 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U9777 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8743) );
  OAI21_X1 U9778 ( .B1(n9014), .B2(n8094), .A(n8743), .ZN(n8101) );
  INV_X1 U9779 ( .A(n8095), .ZN(n8099) );
  NAND3_X1 U9780 ( .A1(n7948), .A2(n8097), .A3(n8096), .ZN(n8098) );
  AOI21_X1 U9781 ( .B1(n8099), .B2(n8098), .A(n8974), .ZN(n8100) );
  AOI211_X1 U9782 ( .C1(n9011), .C2(n8102), .A(n8101), .B(n8100), .ZN(n8109)
         );
  AND3_X1 U9783 ( .A1(n8105), .A2(n8104), .A3(n8103), .ZN(n8106) );
  OAI21_X1 U9784 ( .B1(n8107), .B2(n8106), .A(n8980), .ZN(n8108) );
  OAI211_X1 U9785 ( .C1(n8110), .C2(n9020), .A(n8109), .B(n8108), .ZN(P2_U3192) );
  NAND2_X1 U9786 ( .A1(n9623), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8111) );
  OAI21_X1 U9787 ( .B1(n8112), .B2(n9623), .A(n8111), .ZN(P1_U3583) );
  NAND2_X1 U9788 ( .A1(n8113), .A2(n8118), .ZN(n8114) );
  XNOR2_X1 U9789 ( .A(n8121), .B(n8680), .ZN(n8250) );
  XNOR2_X1 U9790 ( .A(n8250), .B(n8910), .ZN(n8116) );
  OAI211_X1 U9791 ( .C1(n8117), .C2(n8116), .A(n8252), .B(n8855), .ZN(n8123)
         );
  OAI22_X1 U9792 ( .A1(n8883), .A2(n8396), .B1(n8118), .B2(n8896), .ZN(n8119)
         );
  AOI211_X1 U9793 ( .C1(n8121), .C2(n8886), .A(n8120), .B(n8119), .ZN(n8122)
         );
  OAI211_X1 U9794 ( .C1(n8124), .C2(n8862), .A(n8123), .B(n8122), .ZN(P2_U3179) );
  INV_X1 U9795 ( .A(n8125), .ZN(n8128) );
  OAI222_X1 U9796 ( .A1(n9427), .A2(n8126), .B1(n8605), .B2(n8128), .C1(n5884), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U9797 ( .A1(n10118), .A2(n8129), .B1(n10121), .B2(n8128), .C1(
        n4410), .C2(n4413), .ZN(P1_U3336) );
  INV_X1 U9798 ( .A(n8130), .ZN(n8133) );
  NAND3_X1 U9799 ( .A1(n8133), .A2(n8132), .A3(n8131), .ZN(n8134) );
  XNOR2_X1 U9800 ( .A(n8140), .B(n8137), .ZN(n10189) );
  OAI21_X1 U9801 ( .B1(n8140), .B2(n8139), .A(n8138), .ZN(n8145) );
  OAI22_X1 U9802 ( .A1(n8142), .A2(n9919), .B1(n9921), .B2(n8141), .ZN(n8144)
         );
  NOR2_X1 U9803 ( .A1(n10189), .A2(n8206), .ZN(n8143) );
  AOI211_X1 U9804 ( .C1(n10163), .C2(n8145), .A(n8144), .B(n8143), .ZN(n10188)
         );
  OAI21_X1 U9805 ( .B1(n8136), .B2(n10189), .A(n10188), .ZN(n8146) );
  INV_X2 U9806 ( .A(n10167), .ZN(n9943) );
  NAND2_X1 U9807 ( .A1(n8146), .A2(n9943), .ZN(n8150) );
  AOI211_X1 U9808 ( .C1(n8231), .C2(n7062), .A(n8147), .B(n9971), .ZN(n10186)
         );
  OAI22_X1 U9809 ( .A1(n9943), .A2(n10482), .B1(n9625), .B2(n9962), .ZN(n8148)
         );
  AOI21_X1 U9810 ( .B1(n10178), .B2(n10186), .A(n8148), .ZN(n8149) );
  OAI211_X1 U9811 ( .C1(n6260), .C2(n9976), .A(n8150), .B(n8149), .ZN(P1_U3292) );
  INV_X1 U9812 ( .A(n8152), .ZN(n8154) );
  NAND2_X1 U9813 ( .A1(n8154), .A2(n8153), .ZN(n8190) );
  OAI21_X1 U9814 ( .B1(n8154), .B2(n8153), .A(n8190), .ZN(n8155) );
  NOR2_X1 U9815 ( .A1(n8155), .A2(n8156), .ZN(n8193) );
  AOI21_X1 U9816 ( .B1(n8156), .B2(n8155), .A(n8193), .ZN(n8162) );
  INV_X1 U9817 ( .A(n8379), .ZN(n8160) );
  AOI22_X1 U9818 ( .A1(n9606), .A2(n8210), .B1(n9600), .B2(n6377), .ZN(n8158)
         );
  OAI211_X1 U9819 ( .C1(n5028), .C2(n9609), .A(n8158), .B(n8157), .ZN(n8159)
         );
  AOI21_X1 U9820 ( .B1(n8160), .B2(n9590), .A(n8159), .ZN(n8161) );
  OAI21_X1 U9821 ( .B1(n8162), .B2(n9578), .A(n8161), .ZN(P1_U3221) );
  XNOR2_X1 U9822 ( .A(n8163), .B(n8164), .ZN(n8170) );
  INV_X1 U9823 ( .A(n8170), .ZN(n8422) );
  XNOR2_X1 U9824 ( .A(n8165), .B(n8164), .ZN(n8166) );
  NAND2_X1 U9825 ( .A1(n8166), .A2(n9247), .ZN(n8169) );
  OAI22_X1 U9826 ( .A1(n8556), .A2(n9145), .B1(n8781), .B2(n9147), .ZN(n8167)
         );
  INV_X1 U9827 ( .A(n8167), .ZN(n8168) );
  OAI211_X1 U9828 ( .C1(n8170), .C2(n9244), .A(n8169), .B(n8168), .ZN(n8418)
         );
  AOI21_X1 U9829 ( .B1(n10234), .B2(n8422), .A(n8418), .ZN(n8355) );
  AOI22_X1 U9830 ( .A1(n9407), .A2(n8554), .B1(P2_REG0_REG_9__SCAN_IN), .B2(
        n10255), .ZN(n8171) );
  OAI21_X1 U9831 ( .B1(n8355), .B2(n10255), .A(n8171), .ZN(P2_U3417) );
  AND2_X1 U9832 ( .A1(n8202), .A2(n8208), .ZN(n8203) );
  NOR2_X1 U9833 ( .A1(n8203), .A2(n8172), .ZN(n8173) );
  XOR2_X1 U9834 ( .A(n8176), .B(n8173), .Z(n8240) );
  INV_X1 U9835 ( .A(n8174), .ZN(n8209) );
  NOR2_X1 U9836 ( .A1(n8209), .A2(n8208), .ZN(n8178) );
  INV_X1 U9837 ( .A(n8175), .ZN(n8177) );
  OAI21_X1 U9838 ( .B1(n8178), .B2(n8177), .A(n8176), .ZN(n8329) );
  INV_X1 U9839 ( .A(n8329), .ZN(n8180) );
  NOR3_X1 U9840 ( .A1(n8178), .A2(n8177), .A3(n8176), .ZN(n8179) );
  OAI21_X1 U9841 ( .B1(n8180), .B2(n8179), .A(n10163), .ZN(n8182) );
  AOI22_X1 U9842 ( .A1(n10160), .A2(n9621), .B1(n9620), .B2(n10158), .ZN(n8181) );
  OAI211_X1 U9843 ( .C1(n8240), .C2(n8206), .A(n8182), .B(n8181), .ZN(n8242)
         );
  INV_X1 U9844 ( .A(n8242), .ZN(n8183) );
  OAI211_X1 U9845 ( .C1(n8186), .C2(n4509), .A(n8325), .B(n10174), .ZN(n8249)
         );
  OAI211_X1 U9846 ( .C1(n8240), .C2(n10190), .A(n8183), .B(n8249), .ZN(n8188)
         );
  OAI22_X1 U9847 ( .A1(n10066), .A2(n8186), .B1(n10225), .B2(n6334), .ZN(n8184) );
  AOI21_X1 U9848 ( .B1(n8188), .B2(n10225), .A(n8184), .ZN(n8185) );
  INV_X1 U9849 ( .A(n8185), .ZN(P1_U3529) );
  OAI22_X1 U9850 ( .A1(n10102), .A2(n8186), .B1(n10218), .B2(n6339), .ZN(n8187) );
  AOI21_X1 U9851 ( .B1(n8188), .B2(n10218), .A(n8187), .ZN(n8189) );
  INV_X1 U9852 ( .A(n8189), .ZN(P1_U3474) );
  INV_X1 U9853 ( .A(n8190), .ZN(n8191) );
  NOR3_X1 U9854 ( .A1(n8193), .A2(n8192), .A3(n8191), .ZN(n8196) );
  INV_X1 U9855 ( .A(n8194), .ZN(n8195) );
  OAI21_X1 U9856 ( .B1(n8196), .B2(n8195), .A(n9598), .ZN(n8201) );
  AOI21_X1 U9857 ( .B1(n9606), .B2(n9620), .A(n8197), .ZN(n8198) );
  OAI21_X1 U9858 ( .B1(n9586), .B2(n8486), .A(n8198), .ZN(n8199) );
  AOI21_X1 U9859 ( .B1(n8471), .B2(n9576), .A(n8199), .ZN(n8200) );
  OAI211_X1 U9860 ( .C1(n9603), .C2(n8468), .A(n8201), .B(n8200), .ZN(P1_U3231) );
  INV_X1 U9861 ( .A(n8202), .ZN(n8205) );
  INV_X1 U9862 ( .A(n8208), .ZN(n8204) );
  AOI21_X1 U9863 ( .B1(n8205), .B2(n8204), .A(n8203), .ZN(n10214) );
  XNOR2_X1 U9864 ( .A(n8209), .B(n8208), .ZN(n8211) );
  AOI222_X1 U9865 ( .A1(n10163), .A2(n8211), .B1(n8210), .B2(n10158), .C1(
        n10159), .C2(n10160), .ZN(n10213) );
  MUX2_X1 U9866 ( .A(n8212), .B(n10213), .S(n9943), .Z(n8219) );
  INV_X1 U9867 ( .A(n8213), .ZN(n8214) );
  AOI211_X1 U9868 ( .C1(n10210), .C2(n8214), .A(n9971), .B(n4509), .ZN(n10209)
         );
  OAI22_X1 U9869 ( .A1(n9976), .A2(n8216), .B1(n9962), .B2(n8215), .ZN(n8217)
         );
  AOI21_X1 U9870 ( .B1(n10209), .B2(n10178), .A(n8217), .ZN(n8218) );
  OAI211_X1 U9871 ( .C1(n10214), .C2(n9984), .A(n8219), .B(n8218), .ZN(
        P1_U3287) );
  INV_X1 U9872 ( .A(n8220), .ZN(n8230) );
  INV_X1 U9873 ( .A(n8221), .ZN(n8222) );
  MUX2_X1 U9874 ( .A(n8223), .B(n8222), .S(n9943), .Z(n8229) );
  OAI22_X1 U9875 ( .A1(n9976), .A2(n8225), .B1(n9962), .B2(n8224), .ZN(n8226)
         );
  AOI21_X1 U9876 ( .B1(n10178), .B2(n8227), .A(n8226), .ZN(n8228) );
  OAI211_X1 U9877 ( .C1(n9984), .C2(n8230), .A(n8229), .B(n8228), .ZN(P1_U3288) );
  INV_X1 U9878 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8239) );
  NOR2_X1 U9879 ( .A1(n9801), .A2(n9971), .ZN(n9849) );
  OAI21_X1 U9880 ( .B1(n9849), .B2(n10168), .A(n8231), .ZN(n8238) );
  INV_X1 U9881 ( .A(n9962), .ZN(n10166) );
  AOI21_X1 U9882 ( .B1(n10166), .B2(P1_REG3_REG_0__SCAN_IN), .A(n8232), .ZN(
        n8233) );
  OAI21_X1 U9883 ( .B1(n8235), .B2(n8234), .A(n8233), .ZN(n8236) );
  NAND2_X1 U9884 ( .A1(n8236), .A2(n9943), .ZN(n8237) );
  OAI211_X1 U9885 ( .C1(n9943), .C2(n8239), .A(n8238), .B(n8237), .ZN(P1_U3293) );
  NOR2_X1 U9886 ( .A1(n8240), .A2(n8136), .ZN(n8241) );
  OAI21_X1 U9887 ( .B1(n8242), .B2(n8241), .A(n9943), .ZN(n8248) );
  OAI22_X1 U9888 ( .A1(n9943), .A2(n8244), .B1(n8243), .B2(n9962), .ZN(n8245)
         );
  AOI21_X1 U9889 ( .B1(n10168), .B2(n8246), .A(n8245), .ZN(n8247) );
  OAI211_X1 U9890 ( .C1(n8249), .C2(n9801), .A(n8248), .B(n8247), .ZN(P1_U3286) );
  OR2_X1 U9891 ( .A1(n8250), .A2(n8256), .ZN(n8251) );
  XNOR2_X1 U9892 ( .A(n8680), .B(n8259), .ZN(n8391) );
  XNOR2_X1 U9893 ( .A(n8391), .B(n8909), .ZN(n8253) );
  OAI21_X1 U9894 ( .B1(n8254), .B2(n8253), .A(n8393), .ZN(n8255) );
  NAND2_X1 U9895 ( .A1(n8255), .A2(n8855), .ZN(n8261) );
  OAI22_X1 U9896 ( .A1(n8883), .A2(n8556), .B1(n8256), .B2(n8896), .ZN(n8257)
         );
  AOI211_X1 U9897 ( .C1(n8259), .C2(n8886), .A(n8258), .B(n8257), .ZN(n8260)
         );
  OAI211_X1 U9898 ( .C1(n8262), .C2(n8862), .A(n8261), .B(n8260), .ZN(P2_U3153) );
  XOR2_X1 U9899 ( .A(n8263), .B(P2_REG2_REG_11__SCAN_IN), .Z(n8275) );
  INV_X1 U9900 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U9901 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8859) );
  OAI21_X1 U9902 ( .B1(n9014), .B2(n8264), .A(n8859), .ZN(n8270) );
  AOI21_X1 U9903 ( .B1(n8267), .B2(n8266), .A(n8265), .ZN(n8268) );
  NOR2_X1 U9904 ( .A1(n8268), .A2(n9006), .ZN(n8269) );
  AOI211_X1 U9905 ( .C1(n9011), .C2(n8271), .A(n8270), .B(n8269), .ZN(n8274)
         );
  NOR2_X1 U9906 ( .A1(n4514), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8272) );
  OAI21_X1 U9907 ( .B1(n8272), .B2(n4517), .A(n9000), .ZN(n8273) );
  OAI211_X1 U9908 ( .C1(n8275), .C2(n9020), .A(n8274), .B(n8273), .ZN(P2_U3193) );
  NOR2_X1 U9909 ( .A1(n9801), .A2(n8276), .ZN(n8279) );
  OAI22_X1 U9910 ( .A1(n9943), .A2(n8277), .B1(n6262), .B2(n9962), .ZN(n8278)
         );
  AOI211_X1 U9911 ( .C1(n10168), .C2(n8280), .A(n8279), .B(n8278), .ZN(n8283)
         );
  NAND2_X1 U9912 ( .A1(n10179), .A2(n8281), .ZN(n8282) );
  OAI211_X1 U9913 ( .C1(n10167), .C2(n8284), .A(n8283), .B(n8282), .ZN(
        P1_U3291) );
  INV_X1 U9914 ( .A(n8285), .ZN(n8444) );
  OAI222_X1 U9915 ( .A1(P2_U3151), .A2(n8287), .B1(n8605), .B2(n8444), .C1(
        n8286), .C2(n9427), .ZN(P2_U3275) );
  OAI21_X1 U9916 ( .B1(n8290), .B2(n8289), .A(n8288), .ZN(n8318) );
  INV_X1 U9917 ( .A(n8318), .ZN(n8296) );
  OAI21_X1 U9918 ( .B1(n8293), .B2(n8292), .A(n8291), .ZN(n8294) );
  AOI222_X1 U9919 ( .A1(n10163), .A2(n8294), .B1(n9489), .B2(n10158), .C1(
        n6377), .C2(n10160), .ZN(n8321) );
  OAI211_X1 U9920 ( .C1(n8295), .C2(n8308), .A(n10174), .B(n8364), .ZN(n8314)
         );
  OAI211_X1 U9921 ( .C1(n8296), .C2(n10215), .A(n8321), .B(n8314), .ZN(n8302)
         );
  INV_X1 U9922 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8297) );
  OAI22_X1 U9923 ( .A1(n10066), .A2(n8308), .B1(n10225), .B2(n8297), .ZN(n8298) );
  AOI21_X1 U9924 ( .B1(n8302), .B2(n10225), .A(n8298), .ZN(n8299) );
  INV_X1 U9925 ( .A(n8299), .ZN(P1_U3532) );
  OAI22_X1 U9926 ( .A1(n10102), .A2(n8308), .B1(n10218), .B2(n8300), .ZN(n8301) );
  AOI21_X1 U9927 ( .B1(n8302), .B2(n10218), .A(n8301), .ZN(n8303) );
  INV_X1 U9928 ( .A(n8303), .ZN(P1_U3483) );
  AOI21_X1 U9929 ( .B1(n8305), .B2(n8304), .A(n4515), .ZN(n8312) );
  INV_X1 U9930 ( .A(n8313), .ZN(n8310) );
  AOI22_X1 U9931 ( .A1(n9606), .A2(n6377), .B1(n9600), .B2(n9489), .ZN(n8307)
         );
  AND2_X1 U9932 ( .A1(n4410), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10309) );
  INV_X1 U9933 ( .A(n10309), .ZN(n8306) );
  OAI211_X1 U9934 ( .C1(n8308), .C2(n9609), .A(n8307), .B(n8306), .ZN(n8309)
         );
  AOI21_X1 U9935 ( .B1(n8310), .B2(n9590), .A(n8309), .ZN(n8311) );
  OAI21_X1 U9936 ( .B1(n8312), .B2(n9578), .A(n8311), .ZN(P1_U3217) );
  OAI22_X1 U9937 ( .A1(n9943), .A2(n7493), .B1(n8313), .B2(n9962), .ZN(n8316)
         );
  NOR2_X1 U9938 ( .A1(n8314), .A2(n9801), .ZN(n8315) );
  AOI211_X1 U9939 ( .C1(n10168), .C2(n8317), .A(n8316), .B(n8315), .ZN(n8320)
         );
  NAND2_X1 U9940 ( .A1(n8318), .A2(n10179), .ZN(n8319) );
  OAI211_X1 U9941 ( .C1(n8321), .C2(n10167), .A(n8320), .B(n8319), .ZN(
        P1_U3283) );
  OAI21_X1 U9942 ( .B1(n8322), .B2(n8330), .A(n8323), .ZN(n8375) );
  NAND2_X1 U9943 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  NAND2_X1 U9944 ( .A1(n8326), .A2(n10174), .ZN(n8327) );
  NOR2_X1 U9945 ( .A1(n8429), .A2(n8327), .ZN(n8381) );
  NAND2_X1 U9946 ( .A1(n8329), .A2(n8328), .ZN(n8435) );
  XNOR2_X1 U9947 ( .A(n8435), .B(n8330), .ZN(n8331) );
  OAI222_X1 U9948 ( .A1(n9919), .A2(n8333), .B1(n9921), .B2(n8332), .C1(n8331), 
        .C2(n9917), .ZN(n8376) );
  AOI211_X1 U9949 ( .C1(n10206), .C2(n8375), .A(n8381), .B(n8376), .ZN(n8340)
         );
  OAI22_X1 U9950 ( .A1(n10066), .A2(n5028), .B1(n10225), .B2(n8334), .ZN(n8335) );
  INV_X1 U9951 ( .A(n8335), .ZN(n8336) );
  OAI21_X1 U9952 ( .B1(n8340), .B2(n10222), .A(n8336), .ZN(P1_U3530) );
  OAI22_X1 U9953 ( .A1(n10102), .A2(n5028), .B1(n10218), .B2(n8337), .ZN(n8338) );
  INV_X1 U9954 ( .A(n8338), .ZN(n8339) );
  OAI21_X1 U9955 ( .B1(n8340), .B2(n10217), .A(n8339), .ZN(P1_U3477) );
  OAI211_X1 U9956 ( .C1(n8342), .C2(n4787), .A(n8341), .B(n10163), .ZN(n8344)
         );
  INV_X1 U9957 ( .A(n9444), .ZN(n9617) );
  AOI22_X1 U9958 ( .A1(n10160), .A2(n9489), .B1(n9617), .B2(n10158), .ZN(n8343) );
  NAND2_X1 U9959 ( .A1(n8344), .A2(n8343), .ZN(n8496) );
  INV_X1 U9960 ( .A(n8496), .ZN(n8354) );
  OAI21_X1 U9961 ( .B1(n4609), .B2(n8346), .A(n8345), .ZN(n8498) );
  NAND2_X1 U9962 ( .A1(n8498), .A2(n10179), .ZN(n8353) );
  AOI211_X1 U9963 ( .C1(n9494), .C2(n8362), .A(n9971), .B(n8592), .ZN(n8497)
         );
  NOR2_X1 U9964 ( .A1(n8348), .A2(n9976), .ZN(n8351) );
  OAI22_X1 U9965 ( .A1(n9943), .A2(n8349), .B1(n9492), .B2(n9962), .ZN(n8350)
         );
  AOI211_X1 U9966 ( .C1(n8497), .C2(n10178), .A(n8351), .B(n8350), .ZN(n8352)
         );
  OAI211_X1 U9967 ( .C1(n8354), .C2(n10167), .A(n8353), .B(n8352), .ZN(
        P1_U3281) );
  INV_X1 U9968 ( .A(n8554), .ZN(n8557) );
  MUX2_X1 U9969 ( .A(n10495), .B(n8355), .S(n10266), .Z(n8356) );
  OAI21_X1 U9970 ( .B1(n8557), .B2(n9298), .A(n8356), .ZN(P2_U3468) );
  OAI211_X1 U9971 ( .C1(n8359), .C2(n8358), .A(n8357), .B(n10163), .ZN(n8361)
         );
  AOI22_X1 U9972 ( .A1(n10160), .A2(n9619), .B1(n10158), .B2(n9618), .ZN(n8360) );
  NAND2_X1 U9973 ( .A1(n8361), .A2(n8360), .ZN(n8385) );
  INV_X1 U9974 ( .A(n8385), .ZN(n8374) );
  INV_X1 U9975 ( .A(n8362), .ZN(n8363) );
  AOI211_X1 U9976 ( .C1(n8490), .C2(n8364), .A(n9971), .B(n8363), .ZN(n8386)
         );
  INV_X1 U9977 ( .A(n8490), .ZN(n8365) );
  NOR2_X1 U9978 ( .A1(n8365), .A2(n9976), .ZN(n8368) );
  OAI22_X1 U9979 ( .A1(n9943), .A2(n8366), .B1(n8487), .B2(n9962), .ZN(n8367)
         );
  AOI211_X1 U9980 ( .C1(n8386), .C2(n10178), .A(n8368), .B(n8367), .ZN(n8373)
         );
  OAI21_X1 U9981 ( .B1(n8371), .B2(n8370), .A(n8369), .ZN(n8387) );
  NAND2_X1 U9982 ( .A1(n8387), .A2(n10179), .ZN(n8372) );
  OAI211_X1 U9983 ( .C1(n10167), .C2(n8374), .A(n8373), .B(n8372), .ZN(
        P1_U3282) );
  INV_X1 U9984 ( .A(n8375), .ZN(n8384) );
  INV_X1 U9985 ( .A(n8376), .ZN(n8377) );
  MUX2_X1 U9986 ( .A(n8378), .B(n8377), .S(n9943), .Z(n8383) );
  OAI22_X1 U9987 ( .A1(n9976), .A2(n5028), .B1(n9962), .B2(n8379), .ZN(n8380)
         );
  AOI21_X1 U9988 ( .B1(n8381), .B2(n10178), .A(n8380), .ZN(n8382) );
  OAI211_X1 U9989 ( .C1(n8384), .C2(n9984), .A(n8383), .B(n8382), .ZN(P1_U3285) );
  AOI211_X1 U9990 ( .C1(n10206), .C2(n8387), .A(n8386), .B(n8385), .ZN(n8390)
         );
  INV_X1 U9991 ( .A(n10102), .ZN(n10074) );
  AOI22_X1 U9992 ( .A1(n8490), .A2(n10074), .B1(P1_REG0_REG_11__SCAN_IN), .B2(
        n10217), .ZN(n8388) );
  OAI21_X1 U9993 ( .B1(n8390), .B2(n10217), .A(n8388), .ZN(P1_U3486) );
  INV_X1 U9994 ( .A(n10066), .ZN(n9992) );
  AOI22_X1 U9995 ( .A1(n8490), .A2(n9992), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n10222), .ZN(n8389) );
  OAI21_X1 U9996 ( .B1(n8390), .B2(n10222), .A(n8389), .ZN(P1_U3533) );
  NAND2_X1 U9997 ( .A1(n8391), .A2(n8396), .ZN(n8392) );
  XNOR2_X1 U9998 ( .A(n10248), .B(n8680), .ZN(n8551) );
  XNOR2_X1 U9999 ( .A(n8551), .B(n8908), .ZN(n8394) );
  XNOR2_X1 U10000 ( .A(n8549), .B(n8394), .ZN(n8395) );
  NAND2_X1 U10001 ( .A1(n8395), .A2(n8855), .ZN(n8401) );
  OAI22_X1 U10002 ( .A1(n8883), .A2(n8397), .B1(n8396), .B2(n8896), .ZN(n8398)
         );
  AOI211_X1 U10003 ( .C1(n10248), .C2(n8886), .A(n8399), .B(n8398), .ZN(n8400)
         );
  OAI211_X1 U10004 ( .C1(n8402), .C2(n8862), .A(n8401), .B(n8400), .ZN(
        P2_U3161) );
  INV_X1 U10005 ( .A(n8409), .ZN(n8403) );
  XNOR2_X1 U10006 ( .A(n8404), .B(n8403), .ZN(n8405) );
  NAND2_X1 U10007 ( .A1(n8405), .A2(n10163), .ZN(n8407) );
  AOI22_X1 U10008 ( .A1(n10160), .A2(n6273), .B1(n10158), .B2(n9622), .ZN(
        n8406) );
  AND2_X1 U10009 ( .A1(n8407), .A2(n8406), .ZN(n10199) );
  XNOR2_X1 U10010 ( .A(n8408), .B(n8409), .ZN(n10197) );
  NAND2_X1 U10011 ( .A1(n8410), .A2(n8412), .ZN(n8411) );
  NAND3_X1 U10012 ( .A1(n10172), .A2(n10174), .A3(n8411), .ZN(n10194) );
  NAND2_X1 U10013 ( .A1(n10168), .A2(n8412), .ZN(n8415) );
  NOR2_X1 U10014 ( .A1(n9962), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8413) );
  AOI21_X1 U10015 ( .B1(n10167), .B2(P1_REG2_REG_3__SCAN_IN), .A(n8413), .ZN(
        n8414) );
  OAI211_X1 U10016 ( .C1(n10194), .C2(n9801), .A(n8415), .B(n8414), .ZN(n8416)
         );
  AOI21_X1 U10017 ( .B1(n10179), .B2(n10197), .A(n8416), .ZN(n8417) );
  OAI21_X1 U10018 ( .B1(n10167), .B2(n10199), .A(n8417), .ZN(P1_U3290) );
  INV_X1 U10019 ( .A(n9034), .ZN(n8421) );
  OAI22_X1 U10020 ( .A1(n9153), .A2(n8557), .B1(n8562), .B2(n9207), .ZN(n8420)
         );
  MUX2_X1 U10021 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8418), .S(n9253), .Z(n8419)
         );
  AOI211_X1 U10022 ( .C1(n8422), .C2(n8421), .A(n8420), .B(n8419), .ZN(n8423)
         );
  INV_X1 U10023 ( .A(n8423), .ZN(P2_U3224) );
  INV_X1 U10024 ( .A(n8424), .ZN(n8464) );
  OAI222_X1 U10025 ( .A1(n10118), .A2(n8426), .B1(n10121), .B2(n8464), .C1(
        n8425), .C2(n4410), .ZN(P1_U3334) );
  OAI21_X1 U10026 ( .B1(n8428), .B2(n8437), .A(n8427), .ZN(n8475) );
  XNOR2_X1 U10027 ( .A(n8429), .B(n8471), .ZN(n8430) );
  AOI22_X1 U10028 ( .A1(n8430), .A2(n10174), .B1(n10158), .B2(n9619), .ZN(
        n8473) );
  OAI21_X1 U10029 ( .B1(n8431), .B2(n10201), .A(n8473), .ZN(n8440) );
  INV_X1 U10030 ( .A(n8432), .ZN(n8434) );
  OAI21_X1 U10031 ( .B1(n8435), .B2(n8434), .A(n8433), .ZN(n8436) );
  XOR2_X1 U10032 ( .A(n8437), .B(n8436), .Z(n8439) );
  OAI22_X1 U10033 ( .A1(n8439), .A2(n9917), .B1(n8438), .B2(n9921), .ZN(n8467)
         );
  AOI211_X1 U10034 ( .C1(n10206), .C2(n8475), .A(n8440), .B(n8467), .ZN(n8443)
         );
  NAND2_X1 U10035 ( .A1(n10217), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8441) );
  OAI21_X1 U10036 ( .B1(n8443), .B2(n10217), .A(n8441), .ZN(P1_U3480) );
  NAND2_X1 U10037 ( .A1(n10222), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8442) );
  OAI21_X1 U10038 ( .B1(n8443), .B2(n10222), .A(n8442), .ZN(P1_U3531) );
  OAI222_X1 U10039 ( .A1(n4410), .A2(n8445), .B1(n10121), .B2(n8444), .C1(
        n10396), .C2(n10118), .ZN(P1_U3335) );
  XNOR2_X1 U10040 ( .A(n4511), .B(n8446), .ZN(n8456) );
  AOI22_X1 U10041 ( .A1(n9241), .A2(n8742), .B1(n9224), .B2(n9203), .ZN(n8451)
         );
  INV_X1 U10042 ( .A(n8446), .ZN(n8447) );
  XNOR2_X1 U10043 ( .A(n8448), .B(n8447), .ZN(n8449) );
  NAND2_X1 U10044 ( .A1(n8449), .A2(n9247), .ZN(n8450) );
  OAI211_X1 U10045 ( .C1(n8456), .C2(n9244), .A(n8451), .B(n8450), .ZN(n8457)
         );
  MUX2_X1 U10046 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8457), .S(n9253), .Z(n8452) );
  INV_X1 U10047 ( .A(n8452), .ZN(n8455) );
  INV_X1 U10048 ( .A(n8453), .ZN(n8747) );
  AOI22_X1 U10049 ( .A1(n9230), .A2(n8669), .B1(n9250), .B2(n8747), .ZN(n8454)
         );
  OAI211_X1 U10050 ( .C1(n8456), .C2(n9034), .A(n8455), .B(n8454), .ZN(
        P2_U3223) );
  INV_X1 U10051 ( .A(n8456), .ZN(n8458) );
  AOI21_X1 U10052 ( .B1(n10234), .B2(n8458), .A(n8457), .ZN(n8461) );
  MUX2_X1 U10053 ( .A(n8459), .B(n8461), .S(n10254), .Z(n8460) );
  OAI21_X1 U10054 ( .B1(n8745), .B2(n9372), .A(n8460), .ZN(P2_U3420) );
  MUX2_X1 U10055 ( .A(n8462), .B(n8461), .S(n10266), .Z(n8463) );
  OAI21_X1 U10056 ( .B1(n8745), .B2(n9298), .A(n8463), .ZN(P2_U3469) );
  OAI222_X1 U10057 ( .A1(n9427), .A2(n8466), .B1(P2_U3151), .B2(n8465), .C1(
        n9429), .C2(n8464), .ZN(P2_U3274) );
  INV_X1 U10058 ( .A(n8467), .ZN(n8477) );
  OAI22_X1 U10059 ( .A1(n9943), .A2(n8469), .B1(n8468), .B2(n9962), .ZN(n8470)
         );
  AOI21_X1 U10060 ( .B1(n10168), .B2(n8471), .A(n8470), .ZN(n8472) );
  OAI21_X1 U10061 ( .B1(n8473), .B2(n9801), .A(n8472), .ZN(n8474) );
  AOI21_X1 U10062 ( .B1(n8475), .B2(n10179), .A(n8474), .ZN(n8476) );
  OAI21_X1 U10063 ( .B1(n8477), .B2(n10167), .A(n8476), .ZN(P1_U3284) );
  INV_X1 U10064 ( .A(n8478), .ZN(n8483) );
  AOI21_X1 U10065 ( .B1(n8480), .B2(n8482), .A(n8479), .ZN(n8481) );
  AOI21_X1 U10066 ( .B1(n8483), .B2(n8482), .A(n8481), .ZN(n8492) );
  NAND2_X1 U10067 ( .A1(n9600), .A2(n9618), .ZN(n8485) );
  OAI211_X1 U10068 ( .C1(n8486), .C2(n9584), .A(n8485), .B(n8484), .ZN(n8489)
         );
  NOR2_X1 U10069 ( .A1(n9603), .A2(n8487), .ZN(n8488) );
  AOI211_X1 U10070 ( .C1(n8490), .C2(n9576), .A(n8489), .B(n8488), .ZN(n8491)
         );
  OAI21_X1 U10071 ( .B1(n8492), .B2(n9578), .A(n8491), .ZN(P1_U3236) );
  INV_X1 U10072 ( .A(n8509), .ZN(n8495) );
  AOI21_X1 U10073 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10110), .A(n8493), 
        .ZN(n8494) );
  OAI21_X1 U10074 ( .B1(n8495), .B2(n10121), .A(n8494), .ZN(P1_U3332) );
  AOI211_X1 U10075 ( .C1(n10206), .C2(n8498), .A(n8497), .B(n8496), .ZN(n8501)
         );
  AOI22_X1 U10076 ( .A1(n9494), .A2(n9992), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n10222), .ZN(n8499) );
  OAI21_X1 U10077 ( .B1(n8501), .B2(n10222), .A(n8499), .ZN(P1_U3534) );
  AOI22_X1 U10078 ( .A1(n9494), .A2(n10074), .B1(P1_REG0_REG_12__SCAN_IN), 
        .B2(n10217), .ZN(n8500) );
  OAI21_X1 U10079 ( .B1(n8501), .B2(n10217), .A(n8500), .ZN(P1_U3489) );
  INV_X1 U10080 ( .A(n8502), .ZN(n8506) );
  OAI222_X1 U10081 ( .A1(n9427), .A2(n8504), .B1(n8605), .B2(n8506), .C1(n8503), .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U10082 ( .A1(n10118), .A2(n8507), .B1(n10121), .B2(n8506), .C1(
        n4410), .C2(n8505), .ZN(P1_U3333) );
  NAND2_X1 U10083 ( .A1(n8509), .A2(n8508), .ZN(n8511) );
  OAI211_X1 U10084 ( .C1(n8512), .C2(n9427), .A(n8511), .B(n8510), .ZN(
        P2_U3272) );
  XNOR2_X1 U10085 ( .A(n8513), .B(n4893), .ZN(n10060) );
  INV_X1 U10086 ( .A(n8593), .ZN(n8515) );
  INV_X1 U10087 ( .A(n9972), .ZN(n8514) );
  AOI211_X1 U10088 ( .C1(n10058), .C2(n8515), .A(n9971), .B(n8514), .ZN(n10057) );
  NOR2_X1 U10089 ( .A1(n8516), .A2(n9976), .ZN(n8519) );
  INV_X1 U10090 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8517) );
  OAI22_X1 U10091 ( .A1(n9943), .A2(n8517), .B1(n9448), .B2(n9962), .ZN(n8518)
         );
  AOI211_X1 U10092 ( .C1(n10057), .C2(n10178), .A(n8519), .B(n8518), .ZN(n8526) );
  NAND2_X1 U10093 ( .A1(n8520), .A2(n10163), .ZN(n8524) );
  AOI21_X1 U10094 ( .B1(n4739), .B2(n8521), .A(n4893), .ZN(n8523) );
  AOI22_X1 U10095 ( .A1(n9617), .A2(n10160), .B1(n10158), .B2(n9952), .ZN(
        n8522) );
  OAI21_X1 U10096 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n10056) );
  NAND2_X1 U10097 ( .A1(n10056), .A2(n9943), .ZN(n8525) );
  OAI211_X1 U10098 ( .C1(n10060), .C2(n9984), .A(n8526), .B(n8525), .ZN(
        P1_U3279) );
  OAI211_X1 U10099 ( .C1(n8527), .C2(n8533), .A(n9221), .B(n9247), .ZN(n8529)
         );
  AOI22_X1 U10100 ( .A1(n8907), .A2(n9241), .B1(n9203), .B2(n9205), .ZN(n8528)
         );
  NAND2_X1 U10101 ( .A1(n8529), .A2(n8528), .ZN(n8543) );
  MUX2_X1 U10102 ( .A(n8543), .B(P2_REG2_REG_11__SCAN_IN), .S(n9213), .Z(n8530) );
  INV_X1 U10103 ( .A(n8530), .ZN(n8538) );
  NAND2_X1 U10104 ( .A1(n8532), .A2(n8531), .ZN(n8534) );
  XNOR2_X1 U10105 ( .A(n8534), .B(n5171), .ZN(n8546) );
  NAND2_X1 U10106 ( .A1(n9230), .A2(n8670), .ZN(n8535) );
  OAI21_X1 U10107 ( .B1(n8861), .B2(n9207), .A(n8535), .ZN(n8536) );
  AOI21_X1 U10108 ( .B1(n8546), .B2(n9155), .A(n8536), .ZN(n8537) );
  NAND2_X1 U10109 ( .A1(n8538), .A2(n8537), .ZN(P2_U3222) );
  MUX2_X1 U10110 ( .A(n8543), .B(P2_REG0_REG_11__SCAN_IN), .S(n10255), .Z(
        n8539) );
  INV_X1 U10111 ( .A(n8539), .ZN(n8542) );
  INV_X1 U10112 ( .A(n9403), .ZN(n9408) );
  INV_X1 U10113 ( .A(n8670), .ZN(n8867) );
  NOR2_X1 U10114 ( .A1(n9372), .A2(n8867), .ZN(n8540) );
  AOI21_X1 U10115 ( .B1(n8546), .B2(n9408), .A(n8540), .ZN(n8541) );
  NAND2_X1 U10116 ( .A1(n8542), .A2(n8541), .ZN(P2_U3423) );
  MUX2_X1 U10117 ( .A(n8543), .B(P2_REG1_REG_11__SCAN_IN), .S(n6909), .Z(n8544) );
  INV_X1 U10118 ( .A(n8544), .ZN(n8548) );
  INV_X1 U10119 ( .A(n9313), .ZN(n9316) );
  NOR2_X1 U10120 ( .A1(n9298), .A2(n8867), .ZN(n8545) );
  AOI21_X1 U10121 ( .B1(n8546), .B2(n9316), .A(n8545), .ZN(n8547) );
  NAND2_X1 U10122 ( .A1(n8548), .A2(n8547), .ZN(P2_U3470) );
  AND2_X1 U10123 ( .A1(n8551), .A2(n8556), .ZN(n8550) );
  INV_X1 U10124 ( .A(n8551), .ZN(n8552) );
  NAND2_X1 U10125 ( .A1(n8552), .A2(n8908), .ZN(n8553) );
  XNOR2_X1 U10126 ( .A(n8554), .B(n8680), .ZN(n8665) );
  XNOR2_X1 U10127 ( .A(n8665), .B(n8742), .ZN(n8663) );
  XOR2_X1 U10128 ( .A(n8664), .B(n8663), .Z(n8555) );
  NAND2_X1 U10129 ( .A1(n8555), .A2(n8855), .ZN(n8561) );
  OAI22_X1 U10130 ( .A1(n8902), .A2(n8557), .B1(n8556), .B2(n8896), .ZN(n8558)
         );
  AOI211_X1 U10131 ( .C1(n8894), .C2(n8907), .A(n8559), .B(n8558), .ZN(n8560)
         );
  OAI211_X1 U10132 ( .C1(n8562), .C2(n8862), .A(n8561), .B(n8560), .ZN(
        P2_U3171) );
  INV_X1 U10133 ( .A(n8563), .ZN(n8565) );
  NOR2_X1 U10134 ( .A1(n8565), .A2(n8564), .ZN(n8566) );
  XNOR2_X1 U10135 ( .A(n8567), .B(n8566), .ZN(n8582) );
  INV_X1 U10136 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U10137 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8787) );
  OAI21_X1 U10138 ( .B1(n9014), .B2(n10131), .A(n8787), .ZN(n8573) );
  OR3_X1 U10139 ( .A1(n4517), .A2(n8569), .A3(n8568), .ZN(n8570) );
  AOI21_X1 U10140 ( .B1(n8571), .B2(n8570), .A(n8974), .ZN(n8572) );
  AOI211_X1 U10141 ( .C1(n9011), .C2(n8574), .A(n8573), .B(n8572), .ZN(n8581)
         );
  OAI21_X1 U10142 ( .B1(n8577), .B2(n8576), .A(n8575), .ZN(n8579) );
  NAND2_X1 U10143 ( .A1(n8579), .A2(n8578), .ZN(n8580) );
  OAI211_X1 U10144 ( .C1(n9006), .C2(n8582), .A(n8581), .B(n8580), .ZN(
        P2_U3194) );
  OAI21_X1 U10145 ( .B1(n8584), .B2(n8588), .A(n8583), .ZN(n10063) );
  INV_X1 U10146 ( .A(n10063), .ZN(n8599) );
  INV_X1 U10147 ( .A(n4739), .ZN(n8586) );
  AOI21_X1 U10148 ( .B1(n8588), .B2(n8587), .A(n8586), .ZN(n8589) );
  OAI222_X1 U10149 ( .A1(n9921), .A2(n8591), .B1(n9919), .B2(n8590), .C1(n9917), .C2(n8589), .ZN(n10061) );
  AOI211_X1 U10150 ( .C1(n9555), .C2(n5047), .A(n9971), .B(n8593), .ZN(n10062)
         );
  NAND2_X1 U10151 ( .A1(n10062), .A2(n10178), .ZN(n8596) );
  INV_X1 U10152 ( .A(n9553), .ZN(n8594) );
  AOI22_X1 U10153 ( .A1(n10167), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8594), 
        .B2(n10166), .ZN(n8595) );
  OAI211_X1 U10154 ( .C1(n10103), .C2(n9976), .A(n8596), .B(n8595), .ZN(n8597)
         );
  AOI21_X1 U10155 ( .B1(n10061), .B2(n9943), .A(n8597), .ZN(n8598) );
  OAI21_X1 U10156 ( .B1(n8599), .B2(n9984), .A(n8598), .ZN(P1_U3280) );
  INV_X1 U10157 ( .A(n8600), .ZN(n8603) );
  OAI222_X1 U10158 ( .A1(n8601), .A2(n4410), .B1(n10121), .B2(n8603), .C1(
        n10359), .C2(n10118), .ZN(P1_U3331) );
  OAI222_X1 U10159 ( .A1(n5869), .A2(P2_U3151), .B1(n9429), .B2(n8603), .C1(
        n8602), .C2(n9427), .ZN(P2_U3271) );
  INV_X1 U10160 ( .A(n8604), .ZN(n10124) );
  OAI222_X1 U10161 ( .A1(n5864), .A2(P2_U3151), .B1(n8605), .B2(n10124), .C1(
        n10543), .C2(n9427), .ZN(P2_U3270) );
  INV_X1 U10162 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8608) );
  AND2_X1 U10163 ( .A1(n8606), .A2(n9430), .ZN(n8607) );
  AOI22_X1 U10164 ( .A1(n8609), .A2(n8608), .B1(n8607), .B2(n5864), .ZN(
        P2_U3377) );
  INV_X1 U10165 ( .A(n8610), .ZN(n8614) );
  OAI222_X1 U10166 ( .A1(n9427), .A2(n8612), .B1(n9429), .B2(n8614), .C1(n8611), .C2(P2_U3151), .ZN(P2_U3265) );
  OAI222_X1 U10167 ( .A1(n10118), .A2(n10362), .B1(n10121), .B2(n8614), .C1(
        n4410), .C2(n8613), .ZN(P1_U3325) );
  OAI21_X1 U10168 ( .B1(n8617), .B2(n8616), .A(n8615), .ZN(n10001) );
  AOI211_X1 U10169 ( .C1(n9998), .C2(n9829), .A(n9971), .B(n9813), .ZN(n9997)
         );
  INV_X1 U10170 ( .A(n9998), .ZN(n9594) );
  AOI22_X1 U10171 ( .A1(n9591), .A2(n10166), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10167), .ZN(n8618) );
  OAI21_X1 U10172 ( .B1(n9594), .B2(n9976), .A(n8618), .ZN(n8623) );
  OAI21_X1 U10173 ( .B1(n4416), .B2(n8620), .A(n8619), .ZN(n8621) );
  AOI211_X1 U10174 ( .C1(n9997), .C2(n10178), .A(n8623), .B(n8622), .ZN(n8624)
         );
  OAI21_X1 U10175 ( .B1(n9984), .B2(n10001), .A(n8624), .ZN(P1_U3267) );
  XOR2_X1 U10176 ( .A(n8625), .B(n8633), .Z(n10010) );
  INV_X1 U10177 ( .A(n8626), .ZN(n8628) );
  INV_X1 U10178 ( .A(n9830), .ZN(n8627) );
  AOI211_X1 U10179 ( .C1(n10008), .C2(n8628), .A(n9971), .B(n8627), .ZN(n10007) );
  NOR2_X1 U10180 ( .A1(n9538), .A2(n9976), .ZN(n8631) );
  OAI22_X1 U10181 ( .A1(n9531), .A2(n9962), .B1(n8629), .B2(n9943), .ZN(n8630)
         );
  AOI211_X1 U10182 ( .C1(n10007), .C2(n10178), .A(n8631), .B(n8630), .ZN(n8636) );
  NAND2_X1 U10183 ( .A1(n9841), .A2(n8632), .ZN(n8634) );
  NAND2_X1 U10184 ( .A1(n10006), .A2(n9943), .ZN(n8635) );
  OAI211_X1 U10185 ( .C1(n10010), .C2(n9984), .A(n8636), .B(n8635), .ZN(
        P1_U3269) );
  NAND2_X1 U10186 ( .A1(n8639), .A2(n8638), .ZN(n8640) );
  XNOR2_X1 U10187 ( .A(n8640), .B(n4781), .ZN(n8641) );
  NAND2_X1 U10188 ( .A1(n8641), .A2(n10179), .ZN(n8648) );
  OAI22_X1 U10189 ( .A1(n8643), .A2(n9962), .B1(n8642), .B2(n9943), .ZN(n8646)
         );
  NOR2_X1 U10190 ( .A1(n8644), .A2(n9801), .ZN(n8645) );
  AOI211_X1 U10191 ( .C1(n10168), .C2(n7359), .A(n8646), .B(n8645), .ZN(n8647)
         );
  OAI211_X1 U10192 ( .C1(n8637), .C2(n10167), .A(n8648), .B(n8647), .ZN(
        P1_U3356) );
  INV_X1 U10193 ( .A(n8649), .ZN(n8657) );
  INV_X1 U10194 ( .A(n8650), .ZN(n8651) );
  AOI22_X1 U10195 ( .A1(n8651), .A2(n10166), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10167), .ZN(n8654) );
  NAND2_X1 U10196 ( .A1(n8652), .A2(n10168), .ZN(n8653) );
  OAI211_X1 U10197 ( .C1(n8655), .C2(n9801), .A(n8654), .B(n8653), .ZN(n8656)
         );
  AOI21_X1 U10198 ( .B1(n8657), .B2(n9943), .A(n8656), .ZN(n8658) );
  OAI21_X1 U10199 ( .B1(n8659), .B2(n9984), .A(n8658), .ZN(P1_U3265) );
  INV_X1 U10200 ( .A(n8660), .ZN(n9417) );
  INV_X1 U10201 ( .A(n8665), .ZN(n8666) );
  NAND2_X1 U10202 ( .A1(n8666), .A2(n8742), .ZN(n8667) );
  XNOR2_X1 U10203 ( .A(n8669), .B(n8680), .ZN(n8671) );
  XNOR2_X1 U10204 ( .A(n8670), .B(n8684), .ZN(n8783) );
  NAND2_X1 U10205 ( .A1(n8783), .A2(n9224), .ZN(n8784) );
  OAI21_X1 U10206 ( .B1(n8781), .B2(n8671), .A(n8784), .ZN(n8677) );
  XNOR2_X1 U10207 ( .A(n9406), .B(n8680), .ZN(n8678) );
  XNOR2_X1 U10208 ( .A(n8678), .B(n9205), .ZN(n8785) );
  INV_X1 U10209 ( .A(n8783), .ZN(n8674) );
  INV_X1 U10210 ( .A(n8671), .ZN(n8741) );
  OAI21_X1 U10211 ( .B1(n8741), .B2(n8907), .A(n9224), .ZN(n8673) );
  NOR2_X1 U10212 ( .A1(n8907), .A2(n9224), .ZN(n8672) );
  AOI22_X1 U10213 ( .A1(n8674), .A2(n8673), .B1(n8672), .B2(n8671), .ZN(n8675)
         );
  INV_X1 U10214 ( .A(n8678), .ZN(n8679) );
  XNOR2_X1 U10215 ( .A(n9400), .B(n8680), .ZN(n8681) );
  INV_X1 U10216 ( .A(n8681), .ZN(n8682) );
  NAND2_X1 U10217 ( .A1(n8682), .A2(n9225), .ZN(n8683) );
  NAND2_X1 U10218 ( .A1(n8723), .A2(n8683), .ZN(n8840) );
  XNOR2_X1 U10219 ( .A(n9394), .B(n8762), .ZN(n8686) );
  XNOR2_X1 U10220 ( .A(n8686), .B(n9204), .ZN(n8724) );
  NAND2_X1 U10221 ( .A1(n8685), .A2(n8724), .ZN(n8725) );
  NAND2_X1 U10222 ( .A1(n8686), .A2(n8897), .ZN(n8687) );
  XNOR2_X1 U10223 ( .A(n9388), .B(n8762), .ZN(n8689) );
  XNOR2_X1 U10224 ( .A(n8689), .B(n8807), .ZN(n8890) );
  INV_X1 U10225 ( .A(n8890), .ZN(n8688) );
  INV_X1 U10226 ( .A(n8689), .ZN(n8690) );
  NAND2_X1 U10227 ( .A1(n8690), .A2(n9188), .ZN(n8691) );
  XNOR2_X1 U10228 ( .A(n9382), .B(n8762), .ZN(n8692) );
  NAND2_X1 U10229 ( .A1(n8692), .A2(n8815), .ZN(n8802) );
  INV_X1 U10230 ( .A(n8692), .ZN(n8693) );
  NAND2_X1 U10231 ( .A1(n8693), .A2(n9181), .ZN(n8803) );
  XNOR2_X1 U10232 ( .A(n9376), .B(n8684), .ZN(n8695) );
  XNOR2_X1 U10233 ( .A(n8695), .B(n9171), .ZN(n8812) );
  XNOR2_X1 U10234 ( .A(n9150), .B(n8762), .ZN(n8697) );
  XNOR2_X1 U10235 ( .A(n8697), .B(n9161), .ZN(n8868) );
  NAND2_X1 U10236 ( .A1(n8697), .A2(n8754), .ZN(n8698) );
  XNOR2_X1 U10237 ( .A(n9365), .B(n8762), .ZN(n8699) );
  XNOR2_X1 U10238 ( .A(n8699), .B(n8906), .ZN(n8751) );
  NAND2_X1 U10239 ( .A1(n8699), .A2(n9146), .ZN(n8700) );
  NAND2_X1 U10240 ( .A1(n8701), .A2(n8700), .ZN(n8833) );
  XNOR2_X1 U10241 ( .A(n9124), .B(n8762), .ZN(n8702) );
  XNOR2_X1 U10242 ( .A(n8702), .B(n9136), .ZN(n8834) );
  NAND2_X1 U10243 ( .A1(n8833), .A2(n8834), .ZN(n8704) );
  NAND2_X1 U10244 ( .A1(n8702), .A2(n8776), .ZN(n8703) );
  XNOR2_X1 U10245 ( .A(n9356), .B(n8684), .ZN(n8705) );
  XNOR2_X1 U10246 ( .A(n8705), .B(n9121), .ZN(n8772) );
  NAND2_X1 U10247 ( .A1(n8773), .A2(n8772), .ZN(n8708) );
  INV_X1 U10248 ( .A(n8705), .ZN(n8706) );
  NAND2_X1 U10249 ( .A1(n8706), .A2(n9121), .ZN(n8707) );
  XNOR2_X1 U10250 ( .A(n9350), .B(n8762), .ZN(n8710) );
  XNOR2_X1 U10251 ( .A(n8710), .B(n9111), .ZN(n8848) );
  XNOR2_X1 U10252 ( .A(n9339), .B(n8762), .ZN(n8824) );
  INV_X1 U10253 ( .A(n8820), .ZN(n8711) );
  OAI22_X1 U10254 ( .A1(n8824), .A2(n8823), .B1(n8851), .B2(n8711), .ZN(n8715)
         );
  OAI21_X1 U10255 ( .B1(n8820), .B2(n9099), .A(n9089), .ZN(n8713) );
  NOR2_X1 U10256 ( .A1(n9089), .A2(n9099), .ZN(n8712) );
  AOI22_X1 U10257 ( .A1(n8713), .A2(n8824), .B1(n8712), .B2(n8711), .ZN(n8714)
         );
  XNOR2_X1 U10258 ( .A(n9334), .B(n8762), .ZN(n8716) );
  XNOR2_X1 U10259 ( .A(n8716), .B(n9074), .ZN(n8795) );
  XNOR2_X1 U10260 ( .A(n9268), .B(n8762), .ZN(n8717) );
  NOR2_X1 U10261 ( .A1(n8717), .A2(n8798), .ZN(n8877) );
  NAND2_X1 U10262 ( .A1(n8717), .A2(n8798), .ZN(n8875) );
  XNOR2_X1 U10263 ( .A(n9327), .B(n8762), .ZN(n8759) );
  XOR2_X1 U10264 ( .A(n9050), .B(n8759), .Z(n8760) );
  XNOR2_X1 U10265 ( .A(n8761), .B(n8760), .ZN(n8722) );
  AOI22_X1 U10266 ( .A1(n9062), .A2(n8880), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8719) );
  NAND2_X1 U10267 ( .A1(n9046), .A2(n8899), .ZN(n8718) );
  OAI211_X1 U10268 ( .C1(n6879), .C2(n8883), .A(n8719), .B(n8718), .ZN(n8720)
         );
  AOI21_X1 U10269 ( .B1(n9327), .B2(n8886), .A(n8720), .ZN(n8721) );
  OAI21_X1 U10270 ( .B1(n8722), .B2(n8889), .A(n8721), .ZN(P2_U3154) );
  NOR3_X1 U10271 ( .A1(n4508), .A2(n5119), .A3(n8724), .ZN(n8727) );
  INV_X1 U10272 ( .A(n8725), .ZN(n8726) );
  OAI21_X1 U10273 ( .B1(n8727), .B2(n8726), .A(n8855), .ZN(n8732) );
  NAND2_X1 U10274 ( .A1(n8894), .A2(n9188), .ZN(n8728) );
  NAND2_X1 U10275 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8938) );
  OAI211_X1 U10276 ( .C1(n8729), .C2(n8896), .A(n8728), .B(n8938), .ZN(n8730)
         );
  AOI21_X1 U10277 ( .B1(n9190), .B2(n8899), .A(n8730), .ZN(n8731) );
  OAI211_X1 U10278 ( .C1(n8733), .C2(n8902), .A(n8732), .B(n8731), .ZN(
        P2_U3155) );
  XNOR2_X1 U10279 ( .A(n8821), .B(n8820), .ZN(n8822) );
  XNOR2_X1 U10280 ( .A(n8822), .B(n8851), .ZN(n8738) );
  AOI22_X1 U10281 ( .A1(n9111), .A2(n8880), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8735) );
  NAND2_X1 U10282 ( .A1(n9091), .A2(n8899), .ZN(n8734) );
  OAI211_X1 U10283 ( .C1(n8823), .C2(n8883), .A(n8735), .B(n8734), .ZN(n8736)
         );
  AOI21_X1 U10284 ( .B1(n9344), .B2(n8886), .A(n8736), .ZN(n8737) );
  OAI21_X1 U10285 ( .B1(n8738), .B2(n8889), .A(n8737), .ZN(P2_U3156) );
  XNOR2_X1 U10286 ( .A(n8739), .B(n8907), .ZN(n8740) );
  NOR2_X1 U10287 ( .A1(n8740), .A2(n8741), .ZN(n8780) );
  AOI21_X1 U10288 ( .B1(n8741), .B2(n8740), .A(n8780), .ZN(n8749) );
  AOI22_X1 U10289 ( .A1(n8880), .A2(n8742), .B1(n8894), .B2(n9224), .ZN(n8744)
         );
  OAI211_X1 U10290 ( .C1(n8902), .C2(n8745), .A(n8744), .B(n8743), .ZN(n8746)
         );
  AOI21_X1 U10291 ( .B1(n8747), .B2(n8899), .A(n8746), .ZN(n8748) );
  OAI21_X1 U10292 ( .B1(n8749), .B2(n8889), .A(n8748), .ZN(P2_U3157) );
  XOR2_X1 U10293 ( .A(n8750), .B(n8751), .Z(n8758) );
  NAND2_X1 U10294 ( .A1(n8894), .A2(n9136), .ZN(n8753) );
  OAI211_X1 U10295 ( .C1(n8754), .C2(n8896), .A(n8753), .B(n8752), .ZN(n8755)
         );
  AOI21_X1 U10296 ( .B1(n9138), .B2(n8899), .A(n8755), .ZN(n8757) );
  NAND2_X1 U10297 ( .A1(n9365), .A2(n8886), .ZN(n8756) );
  OAI211_X1 U10298 ( .C1(n8758), .C2(n8889), .A(n8757), .B(n8756), .ZN(
        P2_U3159) );
  OAI22_X1 U10299 ( .A1(n8761), .A2(n8760), .B1(n8884), .B2(n8759), .ZN(n8765)
         );
  XNOR2_X1 U10300 ( .A(n8763), .B(n8762), .ZN(n8764) );
  XNOR2_X1 U10301 ( .A(n8765), .B(n8764), .ZN(n8771) );
  NAND2_X1 U10302 ( .A1(n8905), .A2(n8894), .ZN(n8768) );
  AOI22_X1 U10303 ( .A1(n8766), .A2(n8899), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8767) );
  OAI211_X1 U10304 ( .C1(n8884), .C2(n8896), .A(n8768), .B(n8767), .ZN(n8769)
         );
  AOI21_X1 U10305 ( .B1(n9261), .B2(n8886), .A(n8769), .ZN(n8770) );
  OAI21_X1 U10306 ( .B1(n8771), .B2(n8889), .A(n8770), .ZN(P2_U3160) );
  XOR2_X1 U10307 ( .A(n8773), .B(n8772), .Z(n8779) );
  AOI22_X1 U10308 ( .A1(n9111), .A2(n8894), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8775) );
  NAND2_X1 U10309 ( .A1(n8899), .A2(n9114), .ZN(n8774) );
  OAI211_X1 U10310 ( .C1(n8776), .C2(n8896), .A(n8775), .B(n8774), .ZN(n8777)
         );
  AOI21_X1 U10311 ( .B1(n9356), .B2(n8886), .A(n8777), .ZN(n8778) );
  OAI21_X1 U10312 ( .B1(n8779), .B2(n8889), .A(n8778), .ZN(P2_U3163) );
  INV_X1 U10313 ( .A(n8739), .ZN(n8782) );
  AOI21_X1 U10314 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8858) );
  XNOR2_X1 U10315 ( .A(n8783), .B(n8789), .ZN(n8857) );
  NAND2_X1 U10316 ( .A1(n8858), .A2(n8857), .ZN(n8856) );
  NAND2_X1 U10317 ( .A1(n8856), .A2(n8784), .ZN(n8786) );
  XNOR2_X1 U10318 ( .A(n8786), .B(n8785), .ZN(n8793) );
  NAND2_X1 U10319 ( .A1(n8894), .A2(n9225), .ZN(n8788) );
  OAI211_X1 U10320 ( .C1(n8789), .C2(n8896), .A(n8788), .B(n8787), .ZN(n8791)
         );
  NOR2_X1 U10321 ( .A1(n8862), .A2(n9228), .ZN(n8790) );
  AOI211_X1 U10322 ( .C1(n9406), .C2(n8886), .A(n8791), .B(n8790), .ZN(n8792)
         );
  OAI21_X1 U10323 ( .B1(n8793), .B2(n8889), .A(n8792), .ZN(P2_U3164) );
  XOR2_X1 U10324 ( .A(n8795), .B(n8794), .Z(n8801) );
  AOI22_X1 U10325 ( .A1(n9089), .A2(n8880), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8797) );
  NAND2_X1 U10326 ( .A1(n9066), .A2(n8899), .ZN(n8796) );
  OAI211_X1 U10327 ( .C1(n8798), .C2(n8883), .A(n8797), .B(n8796), .ZN(n8799)
         );
  AOI21_X1 U10328 ( .B1(n9334), .B2(n8886), .A(n8799), .ZN(n8800) );
  OAI21_X1 U10329 ( .B1(n8801), .B2(n8889), .A(n8800), .ZN(P2_U3165) );
  NAND2_X1 U10330 ( .A1(n8803), .A2(n8802), .ZN(n8805) );
  XOR2_X1 U10331 ( .A(n8805), .B(n8804), .Z(n8811) );
  NAND2_X1 U10332 ( .A1(n8894), .A2(n9171), .ZN(n8806) );
  NAND2_X1 U10333 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8966) );
  OAI211_X1 U10334 ( .C1(n8807), .C2(n8896), .A(n8806), .B(n8966), .ZN(n8808)
         );
  AOI21_X1 U10335 ( .B1(n9174), .B2(n8899), .A(n8808), .ZN(n8810) );
  NAND2_X1 U10336 ( .A1(n9382), .A2(n8886), .ZN(n8809) );
  OAI211_X1 U10337 ( .C1(n8811), .C2(n8889), .A(n8810), .B(n8809), .ZN(
        P2_U3166) );
  XOR2_X1 U10338 ( .A(n4596), .B(n8812), .Z(n8819) );
  NAND2_X1 U10339 ( .A1(n8894), .A2(n9161), .ZN(n8814) );
  NAND2_X1 U10340 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8989) );
  OAI211_X1 U10341 ( .C1(n8815), .C2(n8896), .A(n8814), .B(n8989), .ZN(n8816)
         );
  AOI21_X1 U10342 ( .B1(n9163), .B2(n8899), .A(n8816), .ZN(n8818) );
  NAND2_X1 U10343 ( .A1(n9376), .A2(n8886), .ZN(n8817) );
  OAI211_X1 U10344 ( .C1(n8819), .C2(n8889), .A(n8818), .B(n8817), .ZN(
        P2_U3168) );
  OAI22_X1 U10345 ( .A1(n8822), .A2(n9099), .B1(n8821), .B2(n8820), .ZN(n8826)
         );
  XNOR2_X1 U10346 ( .A(n8824), .B(n8823), .ZN(n8825) );
  XNOR2_X1 U10347 ( .A(n8826), .B(n8825), .ZN(n8832) );
  AOI22_X1 U10348 ( .A1(n9099), .A2(n8880), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8828) );
  NAND2_X1 U10349 ( .A1(n9077), .A2(n8899), .ZN(n8827) );
  OAI211_X1 U10350 ( .C1(n8829), .C2(n8883), .A(n8828), .B(n8827), .ZN(n8830)
         );
  AOI21_X1 U10351 ( .B1(n9339), .B2(n8886), .A(n8830), .ZN(n8831) );
  OAI21_X1 U10352 ( .B1(n8832), .B2(n8889), .A(n8831), .ZN(P2_U3169) );
  XOR2_X1 U10353 ( .A(n8833), .B(n8834), .Z(n8839) );
  INV_X1 U10354 ( .A(n9121), .ZN(n9098) );
  AOI22_X1 U10355 ( .A1(n9098), .A2(n8894), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8836) );
  NAND2_X1 U10356 ( .A1(n8899), .A2(n9125), .ZN(n8835) );
  OAI211_X1 U10357 ( .C1(n9146), .C2(n8896), .A(n8836), .B(n8835), .ZN(n8837)
         );
  AOI21_X1 U10358 ( .B1(n9124), .B2(n8886), .A(n8837), .ZN(n8838) );
  OAI21_X1 U10359 ( .B1(n8839), .B2(n8889), .A(n8838), .ZN(P2_U3173) );
  AOI21_X1 U10360 ( .B1(n8841), .B2(n8840), .A(n4508), .ZN(n8846) );
  NAND2_X1 U10361 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8917) );
  OAI21_X1 U10362 ( .B1(n8883), .B2(n8897), .A(n8917), .ZN(n8842) );
  AOI21_X1 U10363 ( .B1(n8880), .B2(n9205), .A(n8842), .ZN(n8843) );
  OAI21_X1 U10364 ( .B1(n9208), .B2(n8862), .A(n8843), .ZN(n8844) );
  AOI21_X1 U10365 ( .B1(n9400), .B2(n8886), .A(n8844), .ZN(n8845) );
  OAI21_X1 U10366 ( .B1(n8846), .B2(n8889), .A(n8845), .ZN(P2_U3174) );
  XOR2_X1 U10367 ( .A(n8848), .B(n8847), .Z(n8854) );
  AOI22_X1 U10368 ( .A1(n9098), .A2(n8880), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8850) );
  NAND2_X1 U10369 ( .A1(n8899), .A2(n9102), .ZN(n8849) );
  OAI211_X1 U10370 ( .C1(n8851), .C2(n8883), .A(n8850), .B(n8849), .ZN(n8852)
         );
  AOI21_X1 U10371 ( .B1(n9350), .B2(n8886), .A(n8852), .ZN(n8853) );
  OAI21_X1 U10372 ( .B1(n8854), .B2(n8889), .A(n8853), .ZN(P2_U3175) );
  OAI211_X1 U10373 ( .C1(n8858), .C2(n8857), .A(n8856), .B(n8855), .ZN(n8866)
         );
  OAI21_X1 U10374 ( .B1(n8883), .B2(n8860), .A(n8859), .ZN(n8864) );
  NOR2_X1 U10375 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  AOI211_X1 U10376 ( .C1(n8880), .C2(n8907), .A(n8864), .B(n8863), .ZN(n8865)
         );
  OAI211_X1 U10377 ( .C1(n8867), .C2(n8902), .A(n8866), .B(n8865), .ZN(
        P2_U3176) );
  XOR2_X1 U10378 ( .A(n8869), .B(n8868), .Z(n8874) );
  NAND2_X1 U10379 ( .A1(n8894), .A2(n8906), .ZN(n8870) );
  NAND2_X1 U10380 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9012) );
  OAI211_X1 U10381 ( .C1(n9144), .C2(n8896), .A(n8870), .B(n9012), .ZN(n8871)
         );
  AOI21_X1 U10382 ( .B1(n9151), .B2(n8899), .A(n8871), .ZN(n8873) );
  NAND2_X1 U10383 ( .A1(n9150), .A2(n8886), .ZN(n8872) );
  OAI211_X1 U10384 ( .C1(n8874), .C2(n8889), .A(n8873), .B(n8872), .ZN(
        P2_U3178) );
  INV_X1 U10385 ( .A(n8875), .ZN(n8876) );
  NOR2_X1 U10386 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  XNOR2_X1 U10387 ( .A(n8879), .B(n8878), .ZN(n8888) );
  AOI22_X1 U10388 ( .A1(n9074), .A2(n8880), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8882) );
  NAND2_X1 U10389 ( .A1(n9054), .A2(n8899), .ZN(n8881) );
  OAI211_X1 U10390 ( .C1(n8884), .C2(n8883), .A(n8882), .B(n8881), .ZN(n8885)
         );
  AOI21_X1 U10391 ( .B1(n9268), .B2(n8886), .A(n8885), .ZN(n8887) );
  OAI21_X1 U10392 ( .B1(n8888), .B2(n8889), .A(n8887), .ZN(P2_U3180) );
  INV_X1 U10393 ( .A(n9388), .ZN(n8903) );
  AOI21_X1 U10394 ( .B1(n8891), .B2(n8890), .A(n8889), .ZN(n8893) );
  NAND2_X1 U10395 ( .A1(n8893), .A2(n8892), .ZN(n8901) );
  NAND2_X1 U10396 ( .A1(n8894), .A2(n9181), .ZN(n8895) );
  NAND2_X1 U10397 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8952) );
  OAI211_X1 U10398 ( .C1(n8897), .C2(n8896), .A(n8895), .B(n8952), .ZN(n8898)
         );
  AOI21_X1 U10399 ( .B1(n9184), .B2(n8899), .A(n8898), .ZN(n8900) );
  OAI211_X1 U10400 ( .C1(n8903), .C2(n8902), .A(n8901), .B(n8900), .ZN(
        P2_U3181) );
  MUX2_X1 U10401 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9023), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10402 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8904), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10403 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8905), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10404 ( .A(n9039), .B(P2_DATAO_REG_28__SCAN_IN), .S(n9003), .Z(
        P2_U3519) );
  MUX2_X1 U10405 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9050), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10406 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n9062), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10407 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9074), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10408 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9089), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10409 ( .A(n9099), .B(P2_DATAO_REG_23__SCAN_IN), .S(n9003), .Z(
        P2_U3514) );
  MUX2_X1 U10410 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9111), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10411 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9098), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10412 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9136), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10413 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8906), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10414 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9161), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10415 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9171), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10416 ( .A(n9181), .B(P2_DATAO_REG_16__SCAN_IN), .S(n9003), .Z(
        P2_U3507) );
  MUX2_X1 U10417 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9188), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10418 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n9204), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10419 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9225), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10420 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n9205), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10421 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9224), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10422 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8907), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10423 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8908), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10424 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8909), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10425 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8910), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10426 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8911), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10427 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n5157), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10428 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9240), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10429 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8912), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10430 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9242), .S(P2_U3893), .Z(
        P2_U3492) );
  XOR2_X1 U10431 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n8913), .Z(n8926) );
  OAI21_X1 U10432 ( .B1(n8916), .B2(n8915), .A(n8914), .ZN(n8924) );
  NAND2_X1 U10433 ( .A1(n8988), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8918) );
  OAI211_X1 U10434 ( .C1(n8969), .C2(n8919), .A(n8918), .B(n8917), .ZN(n8923)
         );
  NAND2_X1 U10435 ( .A1(n8920), .A2(n9310), .ZN(n8921) );
  AOI21_X1 U10436 ( .B1(n8932), .B2(n8921), .A(n8974), .ZN(n8922) );
  AOI211_X1 U10437 ( .C1(n8980), .C2(n8924), .A(n8923), .B(n8922), .ZN(n8925)
         );
  OAI21_X1 U10438 ( .B1(n8926), .B2(n9020), .A(n8925), .ZN(P2_U3195) );
  XNOR2_X1 U10439 ( .A(n8927), .B(n10566), .ZN(n8928) );
  XNOR2_X1 U10440 ( .A(n8929), .B(n8928), .ZN(n8945) );
  AND3_X1 U10441 ( .A1(n8932), .A2(n8931), .A3(n8930), .ZN(n8933) );
  OAI21_X1 U10442 ( .B1(n8934), .B2(n8933), .A(n9000), .ZN(n8944) );
  OAI21_X1 U10443 ( .B1(n8937), .B2(n8936), .A(n8935), .ZN(n8942) );
  NAND2_X1 U10444 ( .A1(n8988), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8939) );
  OAI211_X1 U10445 ( .C1(n8969), .C2(n8940), .A(n8939), .B(n8938), .ZN(n8941)
         );
  AOI21_X1 U10446 ( .B1(n8942), .B2(n8980), .A(n8941), .ZN(n8943) );
  OAI211_X1 U10447 ( .C1(n8945), .C2(n9020), .A(n8944), .B(n8943), .ZN(
        P2_U3196) );
  INV_X1 U10448 ( .A(n8962), .ZN(n8946) );
  AOI21_X1 U10449 ( .B1(n9183), .B2(n8947), .A(n8946), .ZN(n8958) );
  OAI21_X1 U10450 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8948), .A(n8973), .ZN(
        n8956) );
  XOR2_X1 U10451 ( .A(n8950), .B(n8949), .Z(n8951) );
  NOR2_X1 U10452 ( .A1(n8951), .A2(n9006), .ZN(n8955) );
  NAND2_X1 U10453 ( .A1(n8988), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8953) );
  OAI211_X1 U10454 ( .C1(n8969), .C2(n4877), .A(n8953), .B(n8952), .ZN(n8954)
         );
  AOI211_X1 U10455 ( .C1(n8956), .C2(n9000), .A(n8955), .B(n8954), .ZN(n8957)
         );
  OAI21_X1 U10456 ( .B1(n8958), .B2(n9020), .A(n8957), .ZN(P2_U3197) );
  AND2_X1 U10457 ( .A1(n8960), .A2(n8959), .ZN(n8963) );
  AOI21_X1 U10458 ( .B1(n8963), .B2(n8962), .A(n8961), .ZN(n8982) );
  XNOR2_X1 U10459 ( .A(n8965), .B(n8964), .ZN(n8979) );
  NAND2_X1 U10460 ( .A1(n8988), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8967) );
  OAI211_X1 U10461 ( .C1(n8969), .C2(n8968), .A(n8967), .B(n8966), .ZN(n8978)
         );
  INV_X1 U10462 ( .A(n8970), .ZN(n8972) );
  NAND3_X1 U10463 ( .A1(n8973), .A2(n8972), .A3(n8971), .ZN(n8975) );
  AOI21_X1 U10464 ( .B1(n8976), .B2(n8975), .A(n8974), .ZN(n8977) );
  AOI211_X1 U10465 ( .C1(n8980), .C2(n8979), .A(n8978), .B(n8977), .ZN(n8981)
         );
  OAI21_X1 U10466 ( .B1(n8982), .B2(n9020), .A(n8981), .ZN(P2_U3198) );
  XOR2_X1 U10467 ( .A(n8984), .B(n8983), .Z(n8994) );
  OAI21_X1 U10468 ( .B1(n8985), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8999), .ZN(
        n8986) );
  NAND2_X1 U10469 ( .A1(n8986), .A2(n9000), .ZN(n8993) );
  NAND2_X1 U10470 ( .A1(n8988), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8990) );
  OAI211_X1 U10471 ( .C1(n8994), .C2(n9006), .A(n8993), .B(n8992), .ZN(
        P2_U3199) );
  AOI21_X1 U10472 ( .B1(n4504), .B2(n8996), .A(n8995), .ZN(n9021) );
  AND3_X1 U10473 ( .A1(n8999), .A2(n8998), .A3(n8997), .ZN(n9001) );
  OAI21_X1 U10474 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9019) );
  INV_X1 U10475 ( .A(n9007), .ZN(n9004) );
  NOR3_X1 U10476 ( .A1(n9005), .A2(n9004), .A3(n9003), .ZN(n9017) );
  AOI21_X1 U10477 ( .B1(n9008), .B2(n9007), .A(n9006), .ZN(n9010) );
  MUX2_X1 U10478 ( .A(n9011), .B(n9010), .S(n9009), .Z(n9016) );
  INV_X1 U10479 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9013) );
  OAI21_X1 U10480 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(n9015) );
  NOR3_X1 U10481 ( .A1(n9017), .A2(n9016), .A3(n9015), .ZN(n9018) );
  NAND2_X1 U10482 ( .A1(n9023), .A2(n9022), .ZN(n9319) );
  INV_X1 U10483 ( .A(n9319), .ZN(n9025) );
  NOR2_X1 U10484 ( .A1(n9024), .A2(n9207), .ZN(n9031) );
  AOI21_X1 U10485 ( .B1(n9025), .B2(n9253), .A(n9031), .ZN(n9028) );
  NAND2_X1 U10486 ( .A1(n9213), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9026) );
  OAI211_X1 U10487 ( .C1(n9321), .C2(n9153), .A(n9028), .B(n9026), .ZN(
        P2_U3202) );
  NAND2_X1 U10488 ( .A1(n9213), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9027) );
  OAI211_X1 U10489 ( .C1(n9324), .C2(n9153), .A(n9028), .B(n9027), .ZN(
        P2_U3203) );
  NAND2_X1 U10490 ( .A1(n9029), .A2(n9253), .ZN(n9033) );
  NOR2_X1 U10491 ( .A1(n4755), .A2(n9153), .ZN(n9030) );
  AOI211_X1 U10492 ( .C1(n9213), .C2(P2_REG2_REG_29__SCAN_IN), .A(n9031), .B(
        n9030), .ZN(n9032) );
  OAI211_X1 U10493 ( .C1(n9035), .C2(n9034), .A(n9033), .B(n9032), .ZN(
        P2_U3204) );
  XNOR2_X1 U10494 ( .A(n9036), .B(n9037), .ZN(n9330) );
  XOR2_X1 U10495 ( .A(n9038), .B(n9037), .Z(n9043) );
  OR2_X1 U10496 ( .A1(n9253), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9044) );
  AOI22_X1 U10497 ( .A1(n9327), .A2(n9230), .B1(n9250), .B2(n9046), .ZN(n9047)
         );
  OAI211_X1 U10498 ( .C1(n9330), .C2(n9233), .A(n9048), .B(n9047), .ZN(
        P2_U3206) );
  XNOR2_X1 U10499 ( .A(n9049), .B(n9052), .ZN(n9051) );
  XNOR2_X1 U10500 ( .A(n9053), .B(n9052), .ZN(n9269) );
  NAND2_X1 U10501 ( .A1(n9268), .A2(n9230), .ZN(n9056) );
  AOI22_X1 U10502 ( .A1(n9054), .A2(n9250), .B1(n9213), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U10503 ( .A1(n9056), .A2(n9055), .ZN(n9057) );
  AOI21_X1 U10504 ( .B1(n9269), .B2(n9155), .A(n9057), .ZN(n9058) );
  OAI21_X1 U10505 ( .B1(n9271), .B2(n9213), .A(n9058), .ZN(P2_U3207) );
  INV_X1 U10506 ( .A(n9334), .ZN(n9059) );
  NOR2_X1 U10507 ( .A1(n9059), .A2(n9209), .ZN(n9065) );
  XNOR2_X1 U10508 ( .A(n9061), .B(n9060), .ZN(n9063) );
  AOI222_X1 U10509 ( .A1(n9247), .A2(n9063), .B1(n9062), .B2(n9203), .C1(n9089), .C2(n9241), .ZN(n9332) );
  INV_X1 U10510 ( .A(n9332), .ZN(n9064) );
  AOI211_X1 U10511 ( .C1(n9250), .C2(n9066), .A(n9065), .B(n9064), .ZN(n9071)
         );
  XNOR2_X1 U10512 ( .A(n9067), .B(n9068), .ZN(n9337) );
  INV_X1 U10513 ( .A(n9337), .ZN(n9069) );
  AOI22_X1 U10514 ( .A1(n9069), .A2(n9155), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9213), .ZN(n9070) );
  OAI21_X1 U10515 ( .B1(n9071), .B2(n9213), .A(n9070), .ZN(P2_U3208) );
  INV_X1 U10516 ( .A(n9339), .ZN(n9072) );
  NOR2_X1 U10517 ( .A1(n9072), .A2(n9209), .ZN(n9076) );
  XOR2_X1 U10518 ( .A(n9082), .B(n9073), .Z(n9075) );
  AOI222_X1 U10519 ( .A1(n9247), .A2(n9075), .B1(n9099), .B2(n9241), .C1(n9074), .C2(n9203), .ZN(n9338) );
  INV_X1 U10520 ( .A(n9079), .ZN(n9081) );
  OAI21_X1 U10521 ( .B1(n9078), .B2(n9081), .A(n9080), .ZN(n9083) );
  XNOR2_X1 U10522 ( .A(n9083), .B(n9082), .ZN(n9342) );
  INV_X1 U10523 ( .A(n9342), .ZN(n9084) );
  AOI22_X1 U10524 ( .A1(n9084), .A2(n9155), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9213), .ZN(n9085) );
  OAI21_X1 U10525 ( .B1(n9086), .B2(n9213), .A(n9085), .ZN(P2_U3209) );
  XOR2_X1 U10526 ( .A(n9078), .B(n9088), .Z(n9347) );
  XNOR2_X1 U10527 ( .A(n9087), .B(n9088), .ZN(n9090) );
  AOI222_X1 U10528 ( .A1(n9247), .A2(n9090), .B1(n9089), .B2(n9203), .C1(n9111), .C2(n9241), .ZN(n9343) );
  MUX2_X1 U10529 ( .A(n10442), .B(n9343), .S(n9253), .Z(n9093) );
  AOI22_X1 U10530 ( .A1(n9344), .A2(n9230), .B1(n9250), .B2(n9091), .ZN(n9092)
         );
  OAI211_X1 U10531 ( .C1(n9347), .C2(n9233), .A(n9093), .B(n9092), .ZN(
        P2_U3210) );
  XNOR2_X1 U10532 ( .A(n9095), .B(n9094), .ZN(n9353) );
  XNOR2_X1 U10533 ( .A(n9096), .B(n9097), .ZN(n9100) );
  AOI222_X1 U10534 ( .A1(n9247), .A2(n9100), .B1(n9099), .B2(n9203), .C1(n9098), .C2(n9241), .ZN(n9348) );
  MUX2_X1 U10535 ( .A(n9101), .B(n9348), .S(n9253), .Z(n9104) );
  AOI22_X1 U10536 ( .A1(n9350), .A2(n9230), .B1(n9250), .B2(n9102), .ZN(n9103)
         );
  OAI211_X1 U10537 ( .C1(n9353), .C2(n9233), .A(n9104), .B(n9103), .ZN(
        P2_U3211) );
  XNOR2_X1 U10538 ( .A(n9105), .B(n9110), .ZN(n9359) );
  INV_X1 U10539 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U10540 ( .A1(n9106), .A2(n9107), .ZN(n9118) );
  NOR2_X1 U10541 ( .A1(n9118), .A2(n9119), .ZN(n9117) );
  NOR2_X1 U10542 ( .A1(n9117), .A2(n9108), .ZN(n9109) );
  XOR2_X1 U10543 ( .A(n9110), .B(n9109), .Z(n9112) );
  AOI222_X1 U10544 ( .A1(n9247), .A2(n9112), .B1(n9136), .B2(n9241), .C1(n9111), .C2(n9203), .ZN(n9354) );
  MUX2_X1 U10545 ( .A(n9113), .B(n9354), .S(n9253), .Z(n9116) );
  AOI22_X1 U10546 ( .A1(n9356), .A2(n9230), .B1(n9250), .B2(n9114), .ZN(n9115)
         );
  OAI211_X1 U10547 ( .C1(n9359), .C2(n9233), .A(n9116), .B(n9115), .ZN(
        P2_U3212) );
  AOI21_X1 U10548 ( .B1(n9119), .B2(n9118), .A(n9117), .ZN(n9120) );
  OAI222_X1 U10549 ( .A1(n9147), .A2(n9121), .B1(n9145), .B2(n9146), .C1(n9142), .C2(n9120), .ZN(n9287) );
  INV_X1 U10550 ( .A(n9287), .ZN(n9129) );
  XNOR2_X1 U10551 ( .A(n9123), .B(n9122), .ZN(n9288) );
  INV_X1 U10552 ( .A(n9124), .ZN(n9363) );
  AOI22_X1 U10553 ( .A1(n9213), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9250), .B2(
        n9125), .ZN(n9126) );
  OAI21_X1 U10554 ( .B1(n9363), .B2(n9153), .A(n9126), .ZN(n9127) );
  AOI21_X1 U10555 ( .B1(n9288), .B2(n9155), .A(n9127), .ZN(n9128) );
  OAI21_X1 U10556 ( .B1(n9129), .B2(n9213), .A(n9128), .ZN(P2_U3213) );
  XOR2_X1 U10557 ( .A(n9130), .B(n9133), .Z(n9368) );
  INV_X1 U10558 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9137) );
  AND2_X1 U10559 ( .A1(n9161), .A2(n9241), .ZN(n9135) );
  INV_X1 U10560 ( .A(n9106), .ZN(n9131) );
  AOI211_X1 U10561 ( .C1(n9133), .C2(n9132), .A(n9142), .B(n9131), .ZN(n9134)
         );
  AOI211_X1 U10562 ( .C1(n9203), .C2(n9136), .A(n9135), .B(n9134), .ZN(n9364)
         );
  MUX2_X1 U10563 ( .A(n9137), .B(n9364), .S(n9253), .Z(n9140) );
  AOI22_X1 U10564 ( .A1(n9365), .A2(n9230), .B1(n9250), .B2(n9138), .ZN(n9139)
         );
  OAI211_X1 U10565 ( .C1(n9368), .C2(n9233), .A(n9140), .B(n9139), .ZN(
        P2_U3214) );
  XNOR2_X1 U10566 ( .A(n9141), .B(n9148), .ZN(n9143) );
  OAI222_X1 U10567 ( .A1(n9147), .A2(n9146), .B1(n9145), .B2(n9144), .C1(n9143), .C2(n9142), .ZN(n9294) );
  INV_X1 U10568 ( .A(n9294), .ZN(n9157) );
  XNOR2_X1 U10569 ( .A(n9149), .B(n9148), .ZN(n9295) );
  INV_X1 U10570 ( .A(n9150), .ZN(n9373) );
  AOI22_X1 U10571 ( .A1(n9213), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9250), .B2(
        n9151), .ZN(n9152) );
  OAI21_X1 U10572 ( .B1(n9373), .B2(n9153), .A(n9152), .ZN(n9154) );
  AOI21_X1 U10573 ( .B1(n9295), .B2(n9155), .A(n9154), .ZN(n9156) );
  OAI21_X1 U10574 ( .B1(n9157), .B2(n9213), .A(n9156), .ZN(P2_U3215) );
  XNOR2_X1 U10575 ( .A(n9158), .B(n9159), .ZN(n9379) );
  XNOR2_X1 U10576 ( .A(n9160), .B(n9159), .ZN(n9162) );
  AOI222_X1 U10577 ( .A1(n9247), .A2(n9162), .B1(n9161), .B2(n9203), .C1(n9181), .C2(n9241), .ZN(n9374) );
  MUX2_X1 U10578 ( .A(n10425), .B(n9374), .S(n9253), .Z(n9165) );
  AOI22_X1 U10579 ( .A1(n9376), .A2(n9230), .B1(n9250), .B2(n9163), .ZN(n9164)
         );
  OAI211_X1 U10580 ( .C1(n9379), .C2(n9233), .A(n9165), .B(n9164), .ZN(
        P2_U3216) );
  NAND2_X1 U10581 ( .A1(n9167), .A2(n9166), .ZN(n9168) );
  XNOR2_X1 U10582 ( .A(n9168), .B(n9170), .ZN(n9385) );
  INV_X1 U10583 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9173) );
  XOR2_X1 U10584 ( .A(n9170), .B(n9169), .Z(n9172) );
  AOI222_X1 U10585 ( .A1(n9247), .A2(n9172), .B1(n9171), .B2(n9203), .C1(n9188), .C2(n9241), .ZN(n9380) );
  MUX2_X1 U10586 ( .A(n9173), .B(n9380), .S(n9253), .Z(n9176) );
  AOI22_X1 U10587 ( .A1(n9382), .A2(n9230), .B1(n9250), .B2(n9174), .ZN(n9175)
         );
  OAI211_X1 U10588 ( .C1(n9385), .C2(n9233), .A(n9176), .B(n9175), .ZN(
        P2_U3217) );
  XNOR2_X1 U10589 ( .A(n9177), .B(n9178), .ZN(n9391) );
  XNOR2_X1 U10590 ( .A(n9180), .B(n9179), .ZN(n9182) );
  AOI222_X1 U10591 ( .A1(n9247), .A2(n9182), .B1(n9204), .B2(n9241), .C1(n9181), .C2(n9203), .ZN(n9386) );
  MUX2_X1 U10592 ( .A(n9183), .B(n9386), .S(n9253), .Z(n9186) );
  AOI22_X1 U10593 ( .A1(n9388), .A2(n9230), .B1(n9250), .B2(n9184), .ZN(n9185)
         );
  OAI211_X1 U10594 ( .C1(n9391), .C2(n9233), .A(n9186), .B(n9185), .ZN(
        P2_U3218) );
  XNOR2_X1 U10595 ( .A(n9187), .B(n9194), .ZN(n9189) );
  AOI222_X1 U10596 ( .A1(n9247), .A2(n9189), .B1(n9188), .B2(n9203), .C1(n9225), .C2(n9241), .ZN(n9392) );
  AOI22_X1 U10597 ( .A1(n9394), .A2(n9191), .B1(n9250), .B2(n9190), .ZN(n9192)
         );
  AOI21_X1 U10598 ( .B1(n9392), .B2(n9192), .A(n9213), .ZN(n9196) );
  XOR2_X1 U10599 ( .A(n4625), .B(n9194), .Z(n9397) );
  OAI22_X1 U10600 ( .A1(n9397), .A2(n9233), .B1(n10566), .B2(n9253), .ZN(n9195) );
  OR2_X1 U10601 ( .A1(n9196), .A2(n9195), .ZN(P2_U3219) );
  AOI21_X1 U10602 ( .B1(n9197), .B2(n9198), .A(n9223), .ZN(n9218) );
  NOR2_X1 U10603 ( .A1(n9218), .A2(n9199), .ZN(n9200) );
  XOR2_X1 U10604 ( .A(n9201), .B(n9200), .Z(n9404) );
  XNOR2_X1 U10605 ( .A(n9202), .B(n9201), .ZN(n9206) );
  AOI222_X1 U10606 ( .A1(n9247), .A2(n9206), .B1(n9205), .B2(n9241), .C1(n9204), .C2(n9203), .ZN(n9398) );
  INV_X1 U10607 ( .A(n9398), .ZN(n9212) );
  INV_X1 U10608 ( .A(n9400), .ZN(n9210) );
  OAI22_X1 U10609 ( .A1(n9210), .A2(n9209), .B1(n9208), .B2(n9207), .ZN(n9211)
         );
  OAI21_X1 U10610 ( .B1(n9212), .B2(n9211), .A(n9253), .ZN(n9215) );
  NAND2_X1 U10611 ( .A1(n9213), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9214) );
  OAI211_X1 U10612 ( .C1(n9404), .C2(n9233), .A(n9215), .B(n9214), .ZN(
        P2_U3220) );
  INV_X1 U10613 ( .A(n9223), .ZN(n9217) );
  NOR2_X1 U10614 ( .A1(n9217), .A2(n9216), .ZN(n9219) );
  AOI21_X1 U10615 ( .B1(n9219), .B2(n9197), .A(n9218), .ZN(n9409) );
  INV_X1 U10616 ( .A(n9409), .ZN(n9234) );
  NAND2_X1 U10617 ( .A1(n9221), .A2(n9220), .ZN(n9222) );
  XOR2_X1 U10618 ( .A(n9223), .B(n9222), .Z(n9226) );
  AOI222_X1 U10619 ( .A1(n9247), .A2(n9226), .B1(n9225), .B2(n9203), .C1(n9224), .C2(n9241), .ZN(n9405) );
  MUX2_X1 U10620 ( .A(n9227), .B(n9405), .S(n9253), .Z(n9232) );
  INV_X1 U10621 ( .A(n9228), .ZN(n9229) );
  AOI22_X1 U10622 ( .A1(n9230), .A2(n9406), .B1(n9250), .B2(n9229), .ZN(n9231)
         );
  OAI211_X1 U10623 ( .C1(n9234), .C2(n9233), .A(n9232), .B(n9231), .ZN(
        P2_U3221) );
  INV_X1 U10624 ( .A(n9235), .ZN(n9238) );
  INV_X1 U10625 ( .A(n9236), .ZN(n9237) );
  AOI21_X1 U10626 ( .B1(n9238), .B2(n5955), .A(n9237), .ZN(n10229) );
  XNOR2_X1 U10627 ( .A(n9239), .B(n5955), .ZN(n9246) );
  AOI22_X1 U10628 ( .A1(n9242), .A2(n9241), .B1(n9203), .B2(n9240), .ZN(n9243)
         );
  OAI21_X1 U10629 ( .B1(n10229), .B2(n9244), .A(n9243), .ZN(n9245) );
  AOI21_X1 U10630 ( .B1(n9247), .B2(n9246), .A(n9245), .ZN(n10230) );
  AND2_X1 U10631 ( .A1(n9248), .A2(n10249), .ZN(n10232) );
  AOI22_X1 U10632 ( .A1(n9250), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n10232), .B2(
        n9249), .ZN(n9251) );
  OAI211_X1 U10633 ( .C1(n10229), .C2(n9252), .A(n10230), .B(n9251), .ZN(n9254) );
  MUX2_X1 U10634 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9254), .S(n9253), .Z(
        P2_U3231) );
  NOR2_X1 U10635 ( .A1(n9319), .A2(n6909), .ZN(n9256) );
  AOI21_X1 U10636 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n6909), .A(n9256), .ZN(
        n9255) );
  OAI21_X1 U10637 ( .B1(n9321), .B2(n9298), .A(n9255), .ZN(P2_U3490) );
  AOI21_X1 U10638 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n6909), .A(n9256), .ZN(
        n9257) );
  OAI21_X1 U10639 ( .B1(n9324), .B2(n9298), .A(n9257), .ZN(P2_U3489) );
  NAND2_X1 U10640 ( .A1(n6909), .A2(n10525), .ZN(n9259) );
  NAND2_X1 U10641 ( .A1(n9261), .A2(n9315), .ZN(n9262) );
  OAI211_X1 U10642 ( .C1(n9264), .C2(n9313), .A(n9263), .B(n9262), .ZN(
        P2_U3487) );
  INV_X1 U10643 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9265) );
  MUX2_X1 U10644 ( .A(n9265), .B(n9325), .S(n10266), .Z(n9267) );
  NAND2_X1 U10645 ( .A1(n9327), .A2(n9315), .ZN(n9266) );
  OAI211_X1 U10646 ( .C1(n9330), .C2(n9313), .A(n9267), .B(n9266), .ZN(
        P2_U3486) );
  AOI22_X1 U10647 ( .A1(n9269), .A2(n10250), .B1(n10249), .B2(n9268), .ZN(
        n9270) );
  MUX2_X1 U10648 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9331), .S(n10266), .Z(
        P2_U3485) );
  INV_X1 U10649 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9272) );
  MUX2_X1 U10650 ( .A(n9272), .B(n9332), .S(n10266), .Z(n9274) );
  NAND2_X1 U10651 ( .A1(n9334), .A2(n9315), .ZN(n9273) );
  OAI211_X1 U10652 ( .C1(n9337), .C2(n9313), .A(n9274), .B(n9273), .ZN(
        P2_U3484) );
  INV_X1 U10653 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9275) );
  MUX2_X1 U10654 ( .A(n9275), .B(n9338), .S(n10266), .Z(n9277) );
  NAND2_X1 U10655 ( .A1(n9339), .A2(n9315), .ZN(n9276) );
  OAI211_X1 U10656 ( .C1(n9313), .C2(n9342), .A(n9277), .B(n9276), .ZN(
        P2_U3483) );
  INV_X1 U10657 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9278) );
  MUX2_X1 U10658 ( .A(n9278), .B(n9343), .S(n10266), .Z(n9280) );
  NAND2_X1 U10659 ( .A1(n9344), .A2(n9315), .ZN(n9279) );
  OAI211_X1 U10660 ( .C1(n9347), .C2(n9313), .A(n9280), .B(n9279), .ZN(
        P2_U3482) );
  MUX2_X1 U10661 ( .A(n9281), .B(n9348), .S(n10266), .Z(n9283) );
  NAND2_X1 U10662 ( .A1(n9350), .A2(n9315), .ZN(n9282) );
  OAI211_X1 U10663 ( .C1(n9353), .C2(n9313), .A(n9283), .B(n9282), .ZN(
        P2_U3481) );
  INV_X1 U10664 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9284) );
  MUX2_X1 U10665 ( .A(n9284), .B(n9354), .S(n10266), .Z(n9286) );
  NAND2_X1 U10666 ( .A1(n9356), .A2(n9315), .ZN(n9285) );
  OAI211_X1 U10667 ( .C1(n9313), .C2(n9359), .A(n9286), .B(n9285), .ZN(
        P2_U3480) );
  INV_X1 U10668 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9289) );
  AOI21_X1 U10669 ( .B1(n10250), .B2(n9288), .A(n9287), .ZN(n9360) );
  MUX2_X1 U10670 ( .A(n9289), .B(n9360), .S(n10266), .Z(n9290) );
  OAI21_X1 U10671 ( .B1(n9363), .B2(n9298), .A(n9290), .ZN(P2_U3479) );
  INV_X1 U10672 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9291) );
  MUX2_X1 U10673 ( .A(n9291), .B(n9364), .S(n10266), .Z(n9293) );
  NAND2_X1 U10674 ( .A1(n9365), .A2(n9315), .ZN(n9292) );
  OAI211_X1 U10675 ( .C1(n9313), .C2(n9368), .A(n9293), .B(n9292), .ZN(
        P2_U3478) );
  AOI21_X1 U10676 ( .B1(n10250), .B2(n9295), .A(n9294), .ZN(n9369) );
  MUX2_X1 U10677 ( .A(n9296), .B(n9369), .S(n10266), .Z(n9297) );
  OAI21_X1 U10678 ( .B1(n9373), .B2(n9298), .A(n9297), .ZN(P2_U3477) );
  MUX2_X1 U10679 ( .A(n9299), .B(n9374), .S(n10266), .Z(n9301) );
  NAND2_X1 U10680 ( .A1(n9376), .A2(n9315), .ZN(n9300) );
  OAI211_X1 U10681 ( .C1(n9379), .C2(n9313), .A(n9301), .B(n9300), .ZN(
        P2_U3476) );
  MUX2_X1 U10682 ( .A(n9302), .B(n9380), .S(n10266), .Z(n9304) );
  NAND2_X1 U10683 ( .A1(n9382), .A2(n9315), .ZN(n9303) );
  OAI211_X1 U10684 ( .C1(n9313), .C2(n9385), .A(n9304), .B(n9303), .ZN(
        P2_U3475) );
  INV_X1 U10685 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9305) );
  MUX2_X1 U10686 ( .A(n9305), .B(n9386), .S(n10266), .Z(n9307) );
  NAND2_X1 U10687 ( .A1(n9388), .A2(n9315), .ZN(n9306) );
  OAI211_X1 U10688 ( .C1(n9313), .C2(n9391), .A(n9307), .B(n9306), .ZN(
        P2_U3474) );
  MUX2_X1 U10689 ( .A(n10533), .B(n9392), .S(n10266), .Z(n9309) );
  NAND2_X1 U10690 ( .A1(n9394), .A2(n9315), .ZN(n9308) );
  OAI211_X1 U10691 ( .C1(n9313), .C2(n9397), .A(n9309), .B(n9308), .ZN(
        P2_U3473) );
  MUX2_X1 U10692 ( .A(n9310), .B(n9398), .S(n10266), .Z(n9312) );
  NAND2_X1 U10693 ( .A1(n9400), .A2(n9315), .ZN(n9311) );
  OAI211_X1 U10694 ( .C1(n9313), .C2(n9404), .A(n9312), .B(n9311), .ZN(
        P2_U3472) );
  MUX2_X1 U10695 ( .A(n9314), .B(n9405), .S(n10266), .Z(n9318) );
  AOI22_X1 U10696 ( .A1(n9409), .A2(n9316), .B1(n9315), .B2(n9406), .ZN(n9317)
         );
  NAND2_X1 U10697 ( .A1(n9318), .A2(n9317), .ZN(P2_U3471) );
  NOR2_X1 U10698 ( .A1(n9319), .A2(n10255), .ZN(n9322) );
  AOI21_X1 U10699 ( .B1(n10255), .B2(P2_REG0_REG_31__SCAN_IN), .A(n9322), .ZN(
        n9320) );
  OAI21_X1 U10700 ( .B1(n9321), .B2(n9372), .A(n9320), .ZN(P2_U3458) );
  AOI21_X1 U10701 ( .B1(n10255), .B2(P2_REG0_REG_30__SCAN_IN), .A(n9322), .ZN(
        n9323) );
  OAI21_X1 U10702 ( .B1(n9324), .B2(n9372), .A(n9323), .ZN(P2_U3457) );
  MUX2_X1 U10703 ( .A(n9326), .B(n9325), .S(n10254), .Z(n9329) );
  NAND2_X1 U10704 ( .A1(n9327), .A2(n9407), .ZN(n9328) );
  OAI211_X1 U10705 ( .C1(n9330), .C2(n9403), .A(n9329), .B(n9328), .ZN(
        P2_U3454) );
  MUX2_X1 U10706 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9331), .S(n10254), .Z(
        P2_U3453) );
  MUX2_X1 U10707 ( .A(n9333), .B(n9332), .S(n10254), .Z(n9336) );
  NAND2_X1 U10708 ( .A1(n9334), .A2(n9407), .ZN(n9335) );
  OAI211_X1 U10709 ( .C1(n9337), .C2(n9403), .A(n9336), .B(n9335), .ZN(
        P2_U3452) );
  MUX2_X1 U10710 ( .A(n10511), .B(n9338), .S(n10254), .Z(n9341) );
  NAND2_X1 U10711 ( .A1(n9339), .A2(n9407), .ZN(n9340) );
  OAI211_X1 U10712 ( .C1(n9342), .C2(n9403), .A(n9341), .B(n9340), .ZN(
        P2_U3451) );
  MUX2_X1 U10713 ( .A(n10336), .B(n9343), .S(n10254), .Z(n9346) );
  NAND2_X1 U10714 ( .A1(n9344), .A2(n9407), .ZN(n9345) );
  OAI211_X1 U10715 ( .C1(n9347), .C2(n9403), .A(n9346), .B(n9345), .ZN(
        P2_U3450) );
  INV_X1 U10716 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9349) );
  MUX2_X1 U10717 ( .A(n9349), .B(n9348), .S(n10254), .Z(n9352) );
  NAND2_X1 U10718 ( .A1(n9350), .A2(n9407), .ZN(n9351) );
  OAI211_X1 U10719 ( .C1(n9353), .C2(n9403), .A(n9352), .B(n9351), .ZN(
        P2_U3449) );
  MUX2_X1 U10720 ( .A(n9355), .B(n9354), .S(n10254), .Z(n9358) );
  NAND2_X1 U10721 ( .A1(n9356), .A2(n9407), .ZN(n9357) );
  OAI211_X1 U10722 ( .C1(n9359), .C2(n9403), .A(n9358), .B(n9357), .ZN(
        P2_U3448) );
  MUX2_X1 U10723 ( .A(n9361), .B(n9360), .S(n10254), .Z(n9362) );
  OAI21_X1 U10724 ( .B1(n9363), .B2(n9372), .A(n9362), .ZN(P2_U3447) );
  MUX2_X1 U10725 ( .A(n10510), .B(n9364), .S(n10254), .Z(n9367) );
  NAND2_X1 U10726 ( .A1(n9365), .A2(n9407), .ZN(n9366) );
  OAI211_X1 U10727 ( .C1(n9368), .C2(n9403), .A(n9367), .B(n9366), .ZN(
        P2_U3446) );
  MUX2_X1 U10728 ( .A(n9370), .B(n9369), .S(n10254), .Z(n9371) );
  OAI21_X1 U10729 ( .B1(n9373), .B2(n9372), .A(n9371), .ZN(P2_U3444) );
  INV_X1 U10730 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9375) );
  MUX2_X1 U10731 ( .A(n9375), .B(n9374), .S(n10254), .Z(n9378) );
  NAND2_X1 U10732 ( .A1(n9376), .A2(n9407), .ZN(n9377) );
  OAI211_X1 U10733 ( .C1(n9379), .C2(n9403), .A(n9378), .B(n9377), .ZN(
        P2_U3441) );
  INV_X1 U10734 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9381) );
  MUX2_X1 U10735 ( .A(n9381), .B(n9380), .S(n10254), .Z(n9384) );
  NAND2_X1 U10736 ( .A1(n9382), .A2(n9407), .ZN(n9383) );
  OAI211_X1 U10737 ( .C1(n9385), .C2(n9403), .A(n9384), .B(n9383), .ZN(
        P2_U3438) );
  INV_X1 U10738 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9387) );
  MUX2_X1 U10739 ( .A(n9387), .B(n9386), .S(n10254), .Z(n9390) );
  NAND2_X1 U10740 ( .A1(n9388), .A2(n9407), .ZN(n9389) );
  OAI211_X1 U10741 ( .C1(n9391), .C2(n9403), .A(n9390), .B(n9389), .ZN(
        P2_U3435) );
  INV_X1 U10742 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9393) );
  MUX2_X1 U10743 ( .A(n9393), .B(n9392), .S(n10254), .Z(n9396) );
  NAND2_X1 U10744 ( .A1(n9394), .A2(n9407), .ZN(n9395) );
  OAI211_X1 U10745 ( .C1(n9397), .C2(n9403), .A(n9396), .B(n9395), .ZN(
        P2_U3432) );
  MUX2_X1 U10746 ( .A(n9399), .B(n9398), .S(n10254), .Z(n9402) );
  NAND2_X1 U10747 ( .A1(n9407), .A2(n9400), .ZN(n9401) );
  OAI211_X1 U10748 ( .C1(n9404), .C2(n9403), .A(n9402), .B(n9401), .ZN(
        P2_U3429) );
  MUX2_X1 U10749 ( .A(n10386), .B(n9405), .S(n10254), .Z(n9411) );
  AOI22_X1 U10750 ( .A1(n9409), .A2(n9408), .B1(n9407), .B2(n9406), .ZN(n9410)
         );
  NAND2_X1 U10751 ( .A1(n9411), .A2(n9410), .ZN(P2_U3426) );
  INV_X1 U10752 ( .A(n9412), .ZN(n10112) );
  INV_X1 U10753 ( .A(n9413), .ZN(n9414) );
  NOR4_X1 U10754 ( .A1(n9414), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5267), .A4(
        P2_U3151), .ZN(n9415) );
  AOI21_X1 U10755 ( .B1(n9424), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9415), .ZN(
        n9416) );
  OAI21_X1 U10756 ( .B1(n10112), .B2(n9429), .A(n9416), .ZN(P2_U3264) );
  OAI222_X1 U10757 ( .A1(n9427), .A2(n9418), .B1(P2_U3151), .B2(n5270), .C1(
        n9429), .C2(n9417), .ZN(P2_U3266) );
  INV_X1 U10758 ( .A(n9419), .ZN(n10114) );
  AOI21_X1 U10759 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9424), .A(n9420), .ZN(
        n9421) );
  OAI21_X1 U10760 ( .B1(n10114), .B2(n9429), .A(n9421), .ZN(P2_U3267) );
  INV_X1 U10761 ( .A(n9422), .ZN(n10116) );
  AOI21_X1 U10762 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9424), .A(n9423), .ZN(
        n9425) );
  OAI21_X1 U10763 ( .B1(n10116), .B2(n9429), .A(n9425), .ZN(P2_U3268) );
  INV_X1 U10764 ( .A(n9426), .ZN(n10120) );
  OAI222_X1 U10765 ( .A1(n9430), .A2(P2_U3151), .B1(n9429), .B2(n10120), .C1(
        n9428), .C2(n9427), .ZN(P2_U3269) );
  MUX2_X1 U10766 ( .A(n9431), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10767 ( .B1(n9580), .B2(n9433), .A(n9432), .ZN(n9435) );
  NOR2_X1 U10768 ( .A1(n9818), .A2(n9603), .ZN(n9438) );
  OAI22_X1 U10769 ( .A1(n9828), .A2(n9584), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9436), .ZN(n9437) );
  AOI211_X1 U10770 ( .C1(n9611), .C2(n9600), .A(n9438), .B(n9437), .ZN(n9439)
         );
  INV_X1 U10771 ( .A(n9441), .ZN(n9442) );
  AOI21_X1 U10772 ( .B1(n9443), .B2(n9442), .A(n9505), .ZN(n9451) );
  NOR2_X1 U10773 ( .A1(n9584), .A2(n9444), .ZN(n9445) );
  AOI211_X1 U10774 ( .C1(n9600), .C2(n9952), .A(n9446), .B(n9445), .ZN(n9447)
         );
  OAI21_X1 U10775 ( .B1(n9603), .B2(n9448), .A(n9447), .ZN(n9449) );
  AOI21_X1 U10776 ( .B1(n10058), .B2(n9576), .A(n9449), .ZN(n9450) );
  OAI21_X1 U10777 ( .B1(n9451), .B2(n9578), .A(n9450), .ZN(P1_U3215) );
  NAND2_X1 U10778 ( .A1(n9453), .A2(n9452), .ZN(n9562) );
  NAND2_X1 U10779 ( .A1(n9455), .A2(n9454), .ZN(n9561) );
  INV_X1 U10780 ( .A(n9456), .ZN(n9457) );
  OR2_X1 U10781 ( .A1(n9457), .A2(n9529), .ZN(n9458) );
  AND3_X1 U10782 ( .A1(n9559), .A2(n9561), .A3(n9458), .ZN(n9459) );
  OAI21_X1 U10783 ( .B1(n9530), .B2(n9459), .A(n9598), .ZN(n9465) );
  AOI22_X1 U10784 ( .A1(n9844), .A2(n9600), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        n4410), .ZN(n9462) );
  INV_X1 U10785 ( .A(n9460), .ZN(n9839) );
  NAND2_X1 U10786 ( .A1(n9839), .A2(n9590), .ZN(n9461) );
  OAI211_X1 U10787 ( .C1(n9875), .C2(n9584), .A(n9462), .B(n9461), .ZN(n9463)
         );
  AOI21_X1 U10788 ( .B1(n10011), .B2(n9576), .A(n9463), .ZN(n9464) );
  NAND2_X1 U10789 ( .A1(n9465), .A2(n9464), .ZN(P1_U3216) );
  XNOR2_X1 U10790 ( .A(n9466), .B(n9467), .ZN(n9571) );
  NOR2_X1 U10791 ( .A1(n9571), .A2(n9570), .ZN(n9569) );
  AOI21_X1 U10792 ( .B1(n9467), .B2(n9466), .A(n9569), .ZN(n9471) );
  XNOR2_X1 U10793 ( .A(n9469), .B(n9468), .ZN(n9470) );
  XNOR2_X1 U10794 ( .A(n9471), .B(n9470), .ZN(n9477) );
  NOR2_X1 U10795 ( .A1(n9603), .A2(n9900), .ZN(n9474) );
  AOI22_X1 U10796 ( .A1(n9600), .A2(n9615), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        n4410), .ZN(n9472) );
  OAI21_X1 U10797 ( .B1(n9906), .B2(n9584), .A(n9472), .ZN(n9473) );
  AOI211_X1 U10798 ( .C1(n9475), .C2(n9576), .A(n9474), .B(n9473), .ZN(n9476)
         );
  OAI21_X1 U10799 ( .B1(n9477), .B2(n9578), .A(n9476), .ZN(P1_U3219) );
  XOR2_X1 U10800 ( .A(n9478), .B(n9479), .Z(n9485) );
  AOI22_X1 U10801 ( .A1(n9845), .A2(n9600), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        n4410), .ZN(n9482) );
  INV_X1 U10802 ( .A(n9480), .ZN(n9877) );
  NAND2_X1 U10803 ( .A1(n9590), .A2(n9877), .ZN(n9481) );
  OAI211_X1 U10804 ( .C1(n9907), .C2(n9584), .A(n9482), .B(n9481), .ZN(n9483)
         );
  AOI21_X1 U10805 ( .B1(n9876), .B2(n9576), .A(n9483), .ZN(n9484) );
  OAI21_X1 U10806 ( .B1(n9485), .B2(n9578), .A(n9484), .ZN(P1_U3223) );
  XOR2_X1 U10807 ( .A(n9487), .B(n9486), .Z(n9496) );
  AOI21_X1 U10808 ( .B1(n9600), .B2(n9617), .A(n9488), .ZN(n9491) );
  NAND2_X1 U10809 ( .A1(n9606), .A2(n9489), .ZN(n9490) );
  OAI211_X1 U10810 ( .C1(n9603), .C2(n9492), .A(n9491), .B(n9490), .ZN(n9493)
         );
  AOI21_X1 U10811 ( .B1(n9494), .B2(n9576), .A(n9493), .ZN(n9495) );
  OAI21_X1 U10812 ( .B1(n9496), .B2(n9578), .A(n9495), .ZN(P1_U3224) );
  AOI21_X1 U10813 ( .B1(n4505), .B2(n9498), .A(n9497), .ZN(n9504) );
  OAI22_X1 U10814 ( .A1(n9827), .A2(n9584), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9499), .ZN(n9500) );
  AOI21_X1 U10815 ( .B1(n9613), .B2(n9600), .A(n9500), .ZN(n9501) );
  OAI21_X1 U10816 ( .B1(n9603), .B2(n9831), .A(n9501), .ZN(n9502) );
  AOI21_X1 U10817 ( .B1(n10004), .B2(n9576), .A(n9502), .ZN(n9503) );
  OAI21_X1 U10818 ( .B1(n9504), .B2(n9578), .A(n9503), .ZN(P1_U3225) );
  XNOR2_X1 U10819 ( .A(n9509), .B(n9507), .ZN(n9596) );
  NAND2_X1 U10820 ( .A1(n9596), .A2(n9597), .ZN(n9595) );
  OAI21_X1 U10821 ( .B1(n9509), .B2(n9508), .A(n9595), .ZN(n9513) );
  XNOR2_X1 U10822 ( .A(n9511), .B(n9510), .ZN(n9512) );
  XNOR2_X1 U10823 ( .A(n9513), .B(n9512), .ZN(n9519) );
  NOR2_X1 U10824 ( .A1(n9603), .A2(n9963), .ZN(n9517) );
  NAND2_X1 U10825 ( .A1(n9600), .A2(n9953), .ZN(n9514) );
  NAND2_X1 U10826 ( .A1(n4410), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9717) );
  OAI211_X1 U10827 ( .C1(n9515), .C2(n9584), .A(n9514), .B(n9717), .ZN(n9516)
         );
  AOI211_X1 U10828 ( .C1(n9961), .C2(n9576), .A(n9517), .B(n9516), .ZN(n9518)
         );
  OAI21_X1 U10829 ( .B1(n9519), .B2(n9578), .A(n9518), .ZN(P1_U3226) );
  NOR2_X1 U10830 ( .A1(n4513), .A2(n9520), .ZN(n9521) );
  XNOR2_X1 U10831 ( .A(n9522), .B(n9521), .ZN(n9528) );
  NOR2_X1 U10832 ( .A1(n9603), .A2(n9933), .ZN(n9526) );
  NAND2_X1 U10833 ( .A1(n9600), .A2(n9940), .ZN(n9523) );
  NAND2_X1 U10834 ( .A1(n4410), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9737) );
  OAI211_X1 U10835 ( .C1(n9524), .C2(n9584), .A(n9523), .B(n9737), .ZN(n9525)
         );
  AOI211_X1 U10836 ( .C1(n10043), .C2(n9576), .A(n9526), .B(n9525), .ZN(n9527)
         );
  OAI21_X1 U10837 ( .B1(n9528), .B2(n9578), .A(n9527), .ZN(P1_U3228) );
  INV_X1 U10838 ( .A(n9531), .ZN(n9535) );
  AOI22_X1 U10839 ( .A1(n9614), .A2(n9600), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        n4410), .ZN(n9532) );
  OAI21_X1 U10840 ( .B1(n9533), .B2(n9584), .A(n9532), .ZN(n9534) );
  AOI21_X1 U10841 ( .B1(n9535), .B2(n9590), .A(n9534), .ZN(n9536) );
  OAI211_X1 U10842 ( .C1(n9538), .C2(n9609), .A(n9537), .B(n9536), .ZN(
        P1_U3229) );
  XNOR2_X1 U10843 ( .A(n9540), .B(n9539), .ZN(n9541) );
  XNOR2_X1 U10844 ( .A(n9542), .B(n9541), .ZN(n9547) );
  NAND2_X1 U10845 ( .A1(n9590), .A2(n9891), .ZN(n9544) );
  AOI22_X1 U10846 ( .A1(n9862), .A2(n9600), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        n4410), .ZN(n9543) );
  OAI211_X1 U10847 ( .C1(n9918), .C2(n9584), .A(n9544), .B(n9543), .ZN(n9545)
         );
  AOI21_X1 U10848 ( .B1(n10028), .B2(n9576), .A(n9545), .ZN(n9546) );
  OAI21_X1 U10849 ( .B1(n9547), .B2(n9578), .A(n9546), .ZN(P1_U3233) );
  XOR2_X1 U10850 ( .A(n9549), .B(n9548), .Z(n9557) );
  NAND2_X1 U10851 ( .A1(n9600), .A2(n9979), .ZN(n9550) );
  OAI21_X1 U10852 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9701), .A(n9550), .ZN(
        n9551) );
  AOI21_X1 U10853 ( .B1(n9606), .B2(n9618), .A(n9551), .ZN(n9552) );
  OAI21_X1 U10854 ( .B1(n9603), .B2(n9553), .A(n9552), .ZN(n9554) );
  AOI21_X1 U10855 ( .B1(n9555), .B2(n9576), .A(n9554), .ZN(n9556) );
  OAI21_X1 U10856 ( .B1(n9557), .B2(n9578), .A(n9556), .ZN(P1_U3234) );
  INV_X1 U10857 ( .A(n9561), .ZN(n9558) );
  NOR2_X1 U10858 ( .A1(n9559), .A2(n9558), .ZN(n9564) );
  AOI21_X1 U10859 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9563) );
  OAI21_X1 U10860 ( .B1(n9564), .B2(n9563), .A(n9598), .ZN(n9568) );
  AOI22_X1 U10861 ( .A1(n9861), .A2(n9600), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        n4410), .ZN(n9565) );
  OAI21_X1 U10862 ( .B1(n9886), .B2(n9584), .A(n9565), .ZN(n9566) );
  AOI21_X1 U10863 ( .B1(n9855), .B2(n9590), .A(n9566), .ZN(n9567) );
  OAI211_X1 U10864 ( .C1(n9857), .C2(n9609), .A(n9568), .B(n9567), .ZN(
        P1_U3235) );
  AOI21_X1 U10865 ( .B1(n9571), .B2(n9570), .A(n9569), .ZN(n9579) );
  NAND2_X1 U10866 ( .A1(n9590), .A2(n9923), .ZN(n9574) );
  NOR2_X1 U10867 ( .A1(n9572), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9761) );
  AOI21_X1 U10868 ( .B1(n9600), .B2(n9616), .A(n9761), .ZN(n9573) );
  OAI211_X1 U10869 ( .C1(n9920), .C2(n9584), .A(n9574), .B(n9573), .ZN(n9575)
         );
  AOI21_X1 U10870 ( .B1(n10038), .B2(n9576), .A(n9575), .ZN(n9577) );
  OAI21_X1 U10871 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(P1_U3238) );
  OAI211_X1 U10872 ( .C1(n9582), .C2(n9581), .A(n9580), .B(n9598), .ZN(n9593)
         );
  OAI22_X1 U10873 ( .A1(n9585), .A2(n9584), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9583), .ZN(n9589) );
  NOR2_X1 U10874 ( .A1(n9587), .A2(n9586), .ZN(n9588) );
  AOI211_X1 U10875 ( .C1(n9591), .C2(n9590), .A(n9589), .B(n9588), .ZN(n9592)
         );
  OAI211_X1 U10876 ( .C1(n9594), .C2(n9609), .A(n9593), .B(n9592), .ZN(
        P1_U3240) );
  OAI21_X1 U10877 ( .B1(n9597), .B2(n9596), .A(n9595), .ZN(n9599) );
  NAND2_X1 U10878 ( .A1(n9599), .A2(n9598), .ZN(n9608) );
  NAND2_X1 U10879 ( .A1(n9600), .A2(n9978), .ZN(n9601) );
  OAI21_X1 U10880 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9602), .A(n9601), .ZN(
        n9605) );
  NOR2_X1 U10881 ( .A1(n9603), .A2(n9973), .ZN(n9604) );
  AOI211_X1 U10882 ( .C1(n9606), .C2(n9979), .A(n9605), .B(n9604), .ZN(n9607)
         );
  OAI211_X1 U10883 ( .C1(n5034), .C2(n9609), .A(n9608), .B(n9607), .ZN(
        P1_U3241) );
  MUX2_X1 U10884 ( .A(n9610), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9623), .Z(
        P1_U3584) );
  MUX2_X1 U10885 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9611), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10886 ( .A(n9612), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9623), .Z(
        P1_U3581) );
  MUX2_X1 U10887 ( .A(n9613), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9623), .Z(
        P1_U3580) );
  MUX2_X1 U10888 ( .A(n9614), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9623), .Z(
        P1_U3579) );
  MUX2_X1 U10889 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9844), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10890 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9861), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10891 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9845), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10892 ( .A(n9862), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9623), .Z(
        P1_U3575) );
  MUX2_X1 U10893 ( .A(n9615), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9623), .Z(
        P1_U3574) );
  MUX2_X1 U10894 ( .A(n9616), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9623), .Z(
        P1_U3573) );
  MUX2_X1 U10895 ( .A(n9940), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9623), .Z(
        P1_U3572) );
  MUX2_X1 U10896 ( .A(n9953), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9623), .Z(
        P1_U3571) );
  MUX2_X1 U10897 ( .A(n9978), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9623), .Z(
        P1_U3570) );
  MUX2_X1 U10898 ( .A(n9952), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9623), .Z(
        P1_U3569) );
  MUX2_X1 U10899 ( .A(n9979), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9623), .Z(
        P1_U3568) );
  MUX2_X1 U10900 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9617), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10901 ( .A(n9618), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9623), .Z(
        P1_U3566) );
  MUX2_X1 U10902 ( .A(n9619), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9623), .Z(
        P1_U3564) );
  MUX2_X1 U10903 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n6377), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10904 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9620), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10905 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9621), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10906 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n10159), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10907 ( .A(n9622), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9623), .Z(
        P1_U3558) );
  MUX2_X1 U10908 ( .A(n10161), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9623), .Z(
        P1_U3557) );
  MUX2_X1 U10909 ( .A(n6273), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9623), .Z(
        P1_U3556) );
  MUX2_X1 U10910 ( .A(n6792), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9623), .Z(
        P1_U3555) );
  MUX2_X1 U10911 ( .A(n9624), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9623), .Z(
        P1_U3554) );
  INV_X1 U10912 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9626) );
  OAI22_X1 U10913 ( .A1(n9786), .A2(n9626), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9625), .ZN(n9627) );
  AOI21_X1 U10914 ( .B1(n9777), .B2(n9628), .A(n9627), .ZN(n9638) );
  MUX2_X1 U10915 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9629), .S(n9628), .Z(n9631)
         );
  OAI211_X1 U10916 ( .C1(n9632), .C2(n9631), .A(n9779), .B(n9630), .ZN(n9637)
         );
  OAI211_X1 U10917 ( .C1(n9635), .C2(n9634), .A(n9773), .B(n9633), .ZN(n9636)
         );
  NAND3_X1 U10918 ( .A1(n9638), .A2(n9637), .A3(n9636), .ZN(P1_U3244) );
  NAND2_X1 U10919 ( .A1(n9777), .A2(n9639), .ZN(n9649) );
  AOI22_X1 U10920 ( .A1(n9762), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(n4410), .ZN(n9648) );
  OAI211_X1 U10921 ( .C1(n9642), .C2(n9641), .A(n9773), .B(n9640), .ZN(n9647)
         );
  OAI211_X1 U10922 ( .C1(n9645), .C2(n9644), .A(n9779), .B(n9643), .ZN(n9646)
         );
  NAND4_X1 U10923 ( .A1(n9649), .A2(n9648), .A3(n9647), .A4(n9646), .ZN(
        P1_U3246) );
  INV_X1 U10924 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9651) );
  OAI21_X1 U10925 ( .B1(n9786), .B2(n9651), .A(n9650), .ZN(n9652) );
  AOI21_X1 U10926 ( .B1(n9777), .B2(n9657), .A(n9652), .ZN(n9664) );
  OAI211_X1 U10927 ( .C1(n9655), .C2(n9654), .A(n9773), .B(n9653), .ZN(n9663)
         );
  INV_X1 U10928 ( .A(n9656), .ZN(n9659) );
  MUX2_X1 U10929 ( .A(n7427), .B(P1_REG1_REG_5__SCAN_IN), .S(n9657), .Z(n9658)
         );
  NAND3_X1 U10930 ( .A1(n9660), .A2(n9659), .A3(n9658), .ZN(n9661) );
  NAND3_X1 U10931 ( .A1(n9779), .A2(n9674), .A3(n9661), .ZN(n9662) );
  NAND3_X1 U10932 ( .A1(n9664), .A2(n9663), .A3(n9662), .ZN(P1_U3248) );
  NOR2_X1 U10933 ( .A1(n9766), .A2(n9665), .ZN(n9666) );
  AOI211_X1 U10934 ( .C1(n9762), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9667), .B(
        n9666), .ZN(n9679) );
  OAI211_X1 U10935 ( .C1(n9670), .C2(n9669), .A(n9773), .B(n9668), .ZN(n9678)
         );
  INV_X1 U10936 ( .A(n9671), .ZN(n9676) );
  NAND3_X1 U10937 ( .A1(n9674), .A2(n9673), .A3(n9672), .ZN(n9675) );
  NAND3_X1 U10938 ( .A1(n9779), .A2(n9676), .A3(n9675), .ZN(n9677) );
  NAND3_X1 U10939 ( .A1(n9679), .A2(n9678), .A3(n9677), .ZN(P1_U3249) );
  INV_X1 U10940 ( .A(n9680), .ZN(n9685) );
  OAI21_X1 U10941 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n9684) );
  NAND3_X1 U10942 ( .A1(n9685), .A2(n9779), .A3(n9684), .ZN(n9694) );
  AOI21_X1 U10943 ( .B1(n9762), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10309), .ZN(
        n9693) );
  AOI21_X1 U10944 ( .B1(n9687), .B2(n9686), .A(n9775), .ZN(n9689) );
  NAND2_X1 U10945 ( .A1(n9689), .A2(n9688), .ZN(n9692) );
  NAND2_X1 U10946 ( .A1(n9777), .A2(n9690), .ZN(n9691) );
  NAND4_X1 U10947 ( .A1(n9694), .A2(n9693), .A3(n9692), .A4(n9691), .ZN(
        P1_U3253) );
  INV_X1 U10948 ( .A(n9695), .ZN(n9700) );
  OAI21_X1 U10949 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9699) );
  NAND3_X1 U10950 ( .A1(n9700), .A2(n9779), .A3(n9699), .ZN(n9711) );
  NOR2_X1 U10951 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9701), .ZN(n9702) );
  AOI21_X1 U10952 ( .B1(n9762), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n9702), .ZN(
        n9710) );
  AOI21_X1 U10953 ( .B1(n9704), .B2(n9703), .A(n9775), .ZN(n9706) );
  NAND2_X1 U10954 ( .A1(n9706), .A2(n9705), .ZN(n9709) );
  NAND2_X1 U10955 ( .A1(n9777), .A2(n9707), .ZN(n9708) );
  NAND4_X1 U10956 ( .A1(n9711), .A2(n9710), .A3(n9709), .A4(n9708), .ZN(
        P1_U3256) );
  NOR2_X1 U10957 ( .A1(n9731), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9739) );
  AOI21_X1 U10958 ( .B1(n9731), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9739), .ZN(
        n9714) );
  NOR2_X1 U10959 ( .A1(n9715), .A2(n9714), .ZN(n9716) );
  OAI21_X1 U10960 ( .B1(n9716), .B2(n9740), .A(n9779), .ZN(n9729) );
  INV_X1 U10961 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9718) );
  OAI21_X1 U10962 ( .B1(n9786), .B2(n9718), .A(n9717), .ZN(n9719) );
  AOI21_X1 U10963 ( .B1(n9777), .B2(n9731), .A(n9719), .ZN(n9728) );
  NAND2_X1 U10964 ( .A1(n9721), .A2(n9720), .ZN(n9722) );
  NAND2_X1 U10965 ( .A1(n9723), .A2(n9722), .ZN(n9726) );
  INV_X1 U10966 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9724) );
  MUX2_X1 U10967 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n9724), .S(n9731), .Z(n9725) );
  NAND2_X1 U10968 ( .A1(n9726), .A2(n9725), .ZN(n9733) );
  OAI211_X1 U10969 ( .C1(n9726), .C2(n9725), .A(n9733), .B(n9773), .ZN(n9727)
         );
  NAND3_X1 U10970 ( .A1(n9729), .A2(n9728), .A3(n9727), .ZN(P1_U3259) );
  OR2_X1 U10971 ( .A1(n9749), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9755) );
  NAND2_X1 U10972 ( .A1(n9749), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U10973 ( .A1(n9755), .A2(n9730), .ZN(n9736) );
  NAND2_X1 U10974 ( .A1(n9731), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U10975 ( .A1(n9733), .A2(n9732), .ZN(n9735) );
  INV_X1 U10976 ( .A(n9756), .ZN(n9734) );
  AOI21_X1 U10977 ( .B1(n9736), .B2(n9735), .A(n9734), .ZN(n9748) );
  INV_X1 U10978 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9738) );
  OAI21_X1 U10979 ( .B1(n9786), .B2(n9738), .A(n9737), .ZN(n9746) );
  NOR2_X1 U10980 ( .A1(n9740), .A2(n9739), .ZN(n9742) );
  XNOR2_X1 U10981 ( .A(n9749), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9741) );
  AOI21_X1 U10982 ( .B1(n9742), .B2(n9741), .A(n9752), .ZN(n9744) );
  NOR2_X1 U10983 ( .A1(n9744), .A2(n9743), .ZN(n9745) );
  AOI211_X1 U10984 ( .C1(n9777), .C2(n9749), .A(n9746), .B(n9745), .ZN(n9747)
         );
  OAI21_X1 U10985 ( .B1(n9748), .B2(n9775), .A(n9747), .ZN(P1_U3260) );
  NOR2_X1 U10986 ( .A1(n9749), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9751) );
  XNOR2_X1 U10987 ( .A(n9769), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9750) );
  INV_X1 U10988 ( .A(n9767), .ZN(n9754) );
  OAI21_X1 U10989 ( .B1(n9752), .B2(n9751), .A(n9750), .ZN(n9753) );
  NAND3_X1 U10990 ( .A1(n9754), .A2(n9779), .A3(n9753), .ZN(n9764) );
  NAND2_X1 U10991 ( .A1(n9756), .A2(n9755), .ZN(n9759) );
  INV_X1 U10992 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9757) );
  MUX2_X1 U10993 ( .A(n9757), .B(P1_REG2_REG_18__SCAN_IN), .S(n9769), .Z(n9758) );
  NOR2_X1 U10994 ( .A1(n9759), .A2(n9758), .ZN(n9771) );
  AOI211_X1 U10995 ( .C1(n9759), .C2(n9758), .A(n9771), .B(n9775), .ZN(n9760)
         );
  AOI211_X1 U10996 ( .C1(n9762), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9761), .B(
        n9760), .ZN(n9763) );
  OAI211_X1 U10997 ( .C1(n9766), .C2(n9765), .A(n9764), .B(n9763), .ZN(
        P1_U3261) );
  INV_X1 U10998 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10034) );
  XNOR2_X1 U10999 ( .A(n9768), .B(n10034), .ZN(n9780) );
  INV_X1 U11000 ( .A(n9780), .ZN(n9774) );
  AND2_X1 U11001 ( .A1(n9769), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9770) );
  OR2_X1 U11002 ( .A1(n9771), .A2(n9770), .ZN(n9772) );
  XNOR2_X1 U11003 ( .A(n9772), .B(n10341), .ZN(n9776) );
  AOI22_X1 U11004 ( .A1(n9774), .A2(n9779), .B1(n9773), .B2(n9776), .ZN(n9783)
         );
  NOR2_X1 U11005 ( .A1(n9776), .A2(n9775), .ZN(n9778) );
  AOI211_X1 U11006 ( .C1(n9780), .C2(n9779), .A(n9778), .B(n9777), .ZN(n9782)
         );
  NAND2_X1 U11007 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(n4410), .ZN(n9784) );
  OAI211_X1 U11008 ( .C1(n4859), .C2(n9786), .A(n9785), .B(n9784), .ZN(
        P1_U3262) );
  NOR2_X2 U11009 ( .A1(n10073), .A2(n9794), .ZN(n9796) );
  XNOR2_X1 U11010 ( .A(n9796), .B(n10070), .ZN(n9787) );
  AND2_X1 U11011 ( .A1(n9789), .A2(n9788), .ZN(n9790) );
  INV_X1 U11012 ( .A(n9985), .ZN(n9989) );
  OR2_X1 U11013 ( .A1(n10167), .A2(n9989), .ZN(n9797) );
  NAND2_X1 U11014 ( .A1(n10167), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9791) );
  OAI211_X1 U11015 ( .C1(n10070), .C2(n9976), .A(n9797), .B(n9791), .ZN(n9792)
         );
  AOI21_X1 U11016 ( .B1(n9986), .B2(n10178), .A(n9792), .ZN(n9793) );
  INV_X1 U11017 ( .A(n9793), .ZN(P1_U3263) );
  AND2_X1 U11018 ( .A1(n10073), .A2(n9794), .ZN(n9795) );
  INV_X1 U11019 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9798) );
  OAI21_X1 U11020 ( .B1(n9943), .B2(n9798), .A(n9797), .ZN(n9799) );
  AOI21_X1 U11021 ( .B1(n10073), .B2(n10168), .A(n9799), .ZN(n9800) );
  OAI21_X1 U11022 ( .B1(n9990), .B2(n9801), .A(n9800), .ZN(P1_U3264) );
  OAI21_X1 U11023 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(n9805) );
  NAND2_X1 U11024 ( .A1(n9805), .A2(n10163), .ZN(n9809) );
  OAI22_X1 U11025 ( .A1(n9806), .A2(n9919), .B1(n9828), .B2(n9921), .ZN(n9807)
         );
  INV_X1 U11026 ( .A(n9807), .ZN(n9808) );
  OAI21_X1 U11027 ( .B1(n9812), .B2(n9811), .A(n9810), .ZN(n9995) );
  NAND2_X1 U11028 ( .A1(n9995), .A2(n10179), .ZN(n9822) );
  INV_X1 U11029 ( .A(n9813), .ZN(n9815) );
  AOI211_X1 U11030 ( .C1(n9816), .C2(n9815), .A(n9971), .B(n9814), .ZN(n9994)
         );
  NOR2_X1 U11031 ( .A1(n10078), .A2(n9976), .ZN(n9820) );
  OAI22_X1 U11032 ( .A1(n9818), .A2(n9962), .B1(n9817), .B2(n9943), .ZN(n9819)
         );
  AOI211_X1 U11033 ( .C1(n9994), .C2(n10178), .A(n9820), .B(n9819), .ZN(n9821)
         );
  OAI211_X1 U11034 ( .C1(n10167), .C2(n4480), .A(n9822), .B(n9821), .ZN(
        P1_U3266) );
  XNOR2_X1 U11035 ( .A(n9823), .B(n9826), .ZN(n10005) );
  AOI211_X1 U11036 ( .C1(n10004), .C2(n9830), .A(n9971), .B(n6855), .ZN(n10003) );
  NAND2_X1 U11037 ( .A1(n10003), .A2(n10178), .ZN(n9834) );
  INV_X1 U11038 ( .A(n9831), .ZN(n9832) );
  AOI22_X1 U11039 ( .A1(n9832), .A2(n10166), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10167), .ZN(n9833) );
  OAI211_X1 U11040 ( .C1(n9835), .C2(n9976), .A(n9834), .B(n9833), .ZN(n9836)
         );
  AOI21_X1 U11041 ( .B1(n10002), .B2(n9943), .A(n9836), .ZN(n9837) );
  OAI21_X1 U11042 ( .B1(n9984), .B2(n10005), .A(n9837), .ZN(P1_U3268) );
  XOR2_X1 U11043 ( .A(n9838), .B(n9843), .Z(n10015) );
  AOI21_X1 U11044 ( .B1(n10011), .B2(n9853), .A(n8626), .ZN(n10012) );
  AOI22_X1 U11045 ( .A1(n9839), .A2(n10166), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10167), .ZN(n9840) );
  OAI21_X1 U11046 ( .B1(n5040), .B2(n9976), .A(n9840), .ZN(n9848) );
  OAI21_X1 U11047 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(n9846) );
  AOI222_X1 U11048 ( .A1(n10163), .A2(n9846), .B1(n9845), .B2(n10160), .C1(
        n9844), .C2(n10158), .ZN(n10014) );
  NOR2_X1 U11049 ( .A1(n10014), .A2(n10167), .ZN(n9847) );
  AOI211_X1 U11050 ( .C1(n10012), .C2(n9849), .A(n9848), .B(n9847), .ZN(n9850)
         );
  OAI21_X1 U11051 ( .B1(n9984), .B2(n10015), .A(n9850), .ZN(P1_U3270) );
  XNOR2_X1 U11052 ( .A(n9851), .B(n9860), .ZN(n10020) );
  INV_X1 U11053 ( .A(n9853), .ZN(n9854) );
  AOI211_X1 U11054 ( .C1(n10017), .C2(n5042), .A(n9971), .B(n9854), .ZN(n10016) );
  AOI22_X1 U11055 ( .A1(n9855), .A2(n10166), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10167), .ZN(n9856) );
  OAI21_X1 U11056 ( .B1(n9857), .B2(n9976), .A(n9856), .ZN(n9865) );
  OAI21_X1 U11057 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(n9863) );
  AOI222_X1 U11058 ( .A1(n10163), .A2(n9863), .B1(n9862), .B2(n10160), .C1(
        n9861), .C2(n10158), .ZN(n10019) );
  NOR2_X1 U11059 ( .A1(n10019), .A2(n10167), .ZN(n9864) );
  AOI211_X1 U11060 ( .C1(n10016), .C2(n10178), .A(n9865), .B(n9864), .ZN(n9866) );
  OAI21_X1 U11061 ( .B1(n10020), .B2(n9984), .A(n9866), .ZN(P1_U3271) );
  XNOR2_X1 U11062 ( .A(n9867), .B(n9869), .ZN(n10023) );
  INV_X1 U11063 ( .A(n10023), .ZN(n9882) );
  NOR2_X1 U11064 ( .A1(n9869), .A2(n4841), .ZN(n9873) );
  INV_X1 U11065 ( .A(n9870), .ZN(n9871) );
  AOI21_X1 U11066 ( .B1(n9873), .B2(n9872), .A(n9871), .ZN(n9874) );
  OAI222_X1 U11067 ( .A1(n9919), .A2(n9875), .B1(n9921), .B2(n9907), .C1(n9917), .C2(n9874), .ZN(n10021) );
  INV_X1 U11068 ( .A(n9876), .ZN(n10087) );
  AOI211_X1 U11069 ( .C1(n9876), .C2(n9888), .A(n9971), .B(n9852), .ZN(n10022)
         );
  NAND2_X1 U11070 ( .A1(n10022), .A2(n10178), .ZN(n9879) );
  AOI22_X1 U11071 ( .A1(n9877), .A2(n10166), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10167), .ZN(n9878) );
  OAI211_X1 U11072 ( .C1(n10087), .C2(n9976), .A(n9879), .B(n9878), .ZN(n9880)
         );
  AOI21_X1 U11073 ( .B1(n10021), .B2(n9943), .A(n9880), .ZN(n9881) );
  OAI21_X1 U11074 ( .B1(n9984), .B2(n9882), .A(n9881), .ZN(P1_U3272) );
  XNOR2_X1 U11075 ( .A(n9883), .B(n9884), .ZN(n10030) );
  XOR2_X1 U11076 ( .A(n6835), .B(n9884), .Z(n9885) );
  OAI222_X1 U11077 ( .A1(n9919), .A2(n9886), .B1(n9921), .B2(n9918), .C1(n9917), .C2(n9885), .ZN(n10026) );
  INV_X1 U11078 ( .A(n9887), .ZN(n9890) );
  INV_X1 U11079 ( .A(n9888), .ZN(n9889) );
  AOI211_X1 U11080 ( .C1(n10028), .C2(n9890), .A(n9971), .B(n9889), .ZN(n10027) );
  NAND2_X1 U11081 ( .A1(n10027), .A2(n10178), .ZN(n9893) );
  AOI22_X1 U11082 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n10167), .B1(n9891), 
        .B2(n10166), .ZN(n9892) );
  OAI211_X1 U11083 ( .C1(n9894), .C2(n9976), .A(n9893), .B(n9892), .ZN(n9895)
         );
  AOI21_X1 U11084 ( .B1(n10026), .B2(n9943), .A(n9895), .ZN(n9896) );
  OAI21_X1 U11085 ( .B1(n9984), .B2(n10030), .A(n9896), .ZN(P1_U3273) );
  XOR2_X1 U11086 ( .A(n9897), .B(n9904), .Z(n10033) );
  INV_X1 U11087 ( .A(n10033), .ZN(n9910) );
  OAI21_X1 U11088 ( .B1(n10092), .B2(n9898), .A(n10174), .ZN(n9899) );
  NOR2_X1 U11089 ( .A1(n9899), .A2(n9887), .ZN(n10032) );
  NOR2_X1 U11090 ( .A1(n10092), .A2(n9976), .ZN(n9902) );
  OAI22_X1 U11091 ( .A1(n9943), .A2(n10341), .B1(n9900), .B2(n9962), .ZN(n9901) );
  AOI211_X1 U11092 ( .C1(n10032), .C2(n10178), .A(n9902), .B(n9901), .ZN(n9909) );
  XOR2_X1 U11093 ( .A(n4706), .B(n9904), .Z(n9905) );
  OAI222_X1 U11094 ( .A1(n9919), .A2(n9907), .B1(n9921), .B2(n9906), .C1(n9905), .C2(n9917), .ZN(n10031) );
  NAND2_X1 U11095 ( .A1(n10031), .A2(n9943), .ZN(n9908) );
  OAI211_X1 U11096 ( .C1(n9910), .C2(n9984), .A(n9909), .B(n9908), .ZN(
        P1_U3274) );
  XNOR2_X1 U11097 ( .A(n9911), .B(n9915), .ZN(n10040) );
  INV_X1 U11098 ( .A(n9912), .ZN(n9913) );
  AOI21_X1 U11099 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9916) );
  OAI222_X1 U11100 ( .A1(n9921), .A2(n9920), .B1(n9919), .B2(n9918), .C1(n9917), .C2(n9916), .ZN(n10036) );
  INV_X1 U11101 ( .A(n9931), .ZN(n9922) );
  AOI211_X1 U11102 ( .C1(n10038), .C2(n9922), .A(n9971), .B(n9898), .ZN(n10037) );
  NAND2_X1 U11103 ( .A1(n10037), .A2(n10178), .ZN(n9925) );
  AOI22_X1 U11104 ( .A1(n10167), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9923), 
        .B2(n10166), .ZN(n9924) );
  OAI211_X1 U11105 ( .C1(n9926), .C2(n9976), .A(n9925), .B(n9924), .ZN(n9927)
         );
  AOI21_X1 U11106 ( .B1(n10036), .B2(n9943), .A(n9927), .ZN(n9928) );
  OAI21_X1 U11107 ( .B1(n9984), .B2(n10040), .A(n9928), .ZN(P1_U3275) );
  XNOR2_X1 U11108 ( .A(n9930), .B(n9929), .ZN(n10045) );
  AOI211_X1 U11109 ( .C1(n10043), .C2(n9960), .A(n9971), .B(n9931), .ZN(n10042) );
  INV_X1 U11110 ( .A(n10043), .ZN(n9932) );
  NOR2_X1 U11111 ( .A1(n9932), .A2(n9976), .ZN(n9936) );
  INV_X1 U11112 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9934) );
  OAI22_X1 U11113 ( .A1(n9943), .A2(n9934), .B1(n9933), .B2(n9962), .ZN(n9935)
         );
  AOI211_X1 U11114 ( .C1(n10042), .C2(n10178), .A(n9936), .B(n9935), .ZN(n9945) );
  OAI211_X1 U11115 ( .C1(n9939), .C2(n9938), .A(n9937), .B(n10163), .ZN(n9942)
         );
  AOI22_X1 U11116 ( .A1(n9940), .A2(n10158), .B1(n9978), .B2(n10160), .ZN(
        n9941) );
  NAND2_X1 U11117 ( .A1(n9942), .A2(n9941), .ZN(n10041) );
  NAND2_X1 U11118 ( .A1(n10041), .A2(n9943), .ZN(n9944) );
  OAI211_X1 U11119 ( .C1(n10045), .C2(n9984), .A(n9945), .B(n9944), .ZN(
        P1_U3276) );
  NAND2_X1 U11120 ( .A1(n9946), .A2(n9947), .ZN(n9949) );
  NAND2_X1 U11121 ( .A1(n9949), .A2(n9948), .ZN(n9951) );
  NAND3_X1 U11122 ( .A1(n9951), .A2(n9950), .A3(n10163), .ZN(n9955) );
  AOI22_X1 U11123 ( .A1(n9953), .A2(n10158), .B1(n10160), .B2(n9952), .ZN(
        n9954) );
  NAND2_X1 U11124 ( .A1(n9955), .A2(n9954), .ZN(n10046) );
  INV_X1 U11125 ( .A(n10046), .ZN(n9968) );
  INV_X1 U11126 ( .A(n9956), .ZN(n9957) );
  AOI21_X1 U11127 ( .B1(n6815), .B2(n9958), .A(n9957), .ZN(n10048) );
  NAND2_X1 U11128 ( .A1(n10048), .A2(n10179), .ZN(n9967) );
  AOI211_X1 U11129 ( .C1(n9961), .C2(n9970), .A(n9971), .B(n5032), .ZN(n10047)
         );
  NOR2_X1 U11130 ( .A1(n6854), .A2(n9976), .ZN(n9965) );
  OAI22_X1 U11131 ( .A1(n9943), .A2(n9724), .B1(n9963), .B2(n9962), .ZN(n9964)
         );
  AOI211_X1 U11132 ( .C1(n10047), .C2(n10178), .A(n9965), .B(n9964), .ZN(n9966) );
  OAI211_X1 U11133 ( .C1(n10167), .C2(n9968), .A(n9967), .B(n9966), .ZN(
        P1_U3277) );
  XOR2_X1 U11134 ( .A(n9977), .B(n9969), .Z(n10055) );
  AOI211_X1 U11135 ( .C1(n10052), .C2(n9972), .A(n9971), .B(n9959), .ZN(n10051) );
  INV_X1 U11136 ( .A(n9973), .ZN(n9974) );
  AOI22_X1 U11137 ( .A1(n10167), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9974), 
        .B2(n10166), .ZN(n9975) );
  OAI21_X1 U11138 ( .B1(n5034), .B2(n9976), .A(n9975), .ZN(n9982) );
  OAI21_X1 U11139 ( .B1(n9977), .B2(n4500), .A(n9946), .ZN(n9980) );
  AOI222_X1 U11140 ( .A1(n10163), .A2(n9980), .B1(n9979), .B2(n10160), .C1(
        n9978), .C2(n10158), .ZN(n10054) );
  NOR2_X1 U11141 ( .A1(n10054), .A2(n10167), .ZN(n9981) );
  AOI211_X1 U11142 ( .C1(n10051), .C2(n10178), .A(n9982), .B(n9981), .ZN(n9983) );
  OAI21_X1 U11143 ( .B1(n9984), .B2(n10055), .A(n9983), .ZN(P1_U3278) );
  NOR2_X1 U11144 ( .A1(n9986), .A2(n9985), .ZN(n10067) );
  MUX2_X1 U11145 ( .A(n9987), .B(n10067), .S(n10225), .Z(n9988) );
  OAI21_X1 U11146 ( .B1(n10070), .B2(n10066), .A(n9988), .ZN(P1_U3553) );
  NAND2_X1 U11147 ( .A1(n9990), .A2(n9989), .ZN(n10071) );
  AOI21_X1 U11148 ( .B1(n9992), .B2(n10073), .A(n9991), .ZN(n9993) );
  INV_X1 U11149 ( .A(n9993), .ZN(P1_U3552) );
  INV_X1 U11150 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9996) );
  AOI21_X1 U11151 ( .B1(n10211), .B2(n9998), .A(n9997), .ZN(n9999) );
  OAI211_X1 U11152 ( .C1(n10001), .C2(n10215), .A(n10000), .B(n9999), .ZN(
        n10079) );
  MUX2_X1 U11153 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10079), .S(n10225), .Z(
        P1_U3548) );
  MUX2_X1 U11154 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10080), .S(n10225), .Z(
        P1_U3547) );
  AOI22_X1 U11155 ( .A1(n10012), .A2(n10174), .B1(n10211), .B2(n10011), .ZN(
        n10013) );
  OAI211_X1 U11156 ( .C1(n10015), .C2(n10215), .A(n10014), .B(n10013), .ZN(
        n10082) );
  MUX2_X1 U11157 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10082), .S(n10225), .Z(
        P1_U3545) );
  AOI21_X1 U11158 ( .B1(n10211), .B2(n10017), .A(n10016), .ZN(n10018) );
  OAI211_X1 U11159 ( .C1(n10215), .C2(n10020), .A(n10019), .B(n10018), .ZN(
        n10083) );
  MUX2_X1 U11160 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10083), .S(n10225), .Z(
        P1_U3544) );
  AOI211_X1 U11161 ( .C1(n10023), .C2(n10206), .A(n10022), .B(n10021), .ZN(
        n10084) );
  MUX2_X1 U11162 ( .A(n10024), .B(n10084), .S(n10225), .Z(n10025) );
  OAI21_X1 U11163 ( .B1(n10087), .B2(n10066), .A(n10025), .ZN(P1_U3543) );
  AOI211_X1 U11164 ( .C1(n10211), .C2(n10028), .A(n10027), .B(n10026), .ZN(
        n10029) );
  OAI21_X1 U11165 ( .B1(n10215), .B2(n10030), .A(n10029), .ZN(n10088) );
  MUX2_X1 U11166 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10088), .S(n10225), .Z(
        P1_U3542) );
  AOI211_X1 U11167 ( .C1(n10206), .C2(n10033), .A(n10032), .B(n10031), .ZN(
        n10089) );
  MUX2_X1 U11168 ( .A(n10034), .B(n10089), .S(n10225), .Z(n10035) );
  OAI21_X1 U11169 ( .B1(n10092), .B2(n10066), .A(n10035), .ZN(P1_U3541) );
  AOI211_X1 U11170 ( .C1(n10211), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10039) );
  OAI21_X1 U11171 ( .B1(n10215), .B2(n10040), .A(n10039), .ZN(n10093) );
  MUX2_X1 U11172 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10093), .S(n10225), .Z(
        P1_U3540) );
  AOI211_X1 U11173 ( .C1(n10211), .C2(n10043), .A(n10042), .B(n10041), .ZN(
        n10044) );
  OAI21_X1 U11174 ( .B1(n10215), .B2(n10045), .A(n10044), .ZN(n10094) );
  MUX2_X1 U11175 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10094), .S(n10225), .Z(
        P1_U3539) );
  INV_X1 U11176 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10049) );
  AOI211_X1 U11177 ( .C1(n10048), .C2(n10206), .A(n10047), .B(n10046), .ZN(
        n10095) );
  MUX2_X1 U11178 ( .A(n10049), .B(n10095), .S(n10225), .Z(n10050) );
  OAI21_X1 U11179 ( .B1(n6854), .B2(n10066), .A(n10050), .ZN(P1_U3538) );
  AOI21_X1 U11180 ( .B1(n10211), .B2(n10052), .A(n10051), .ZN(n10053) );
  OAI211_X1 U11181 ( .C1(n10055), .C2(n10215), .A(n10054), .B(n10053), .ZN(
        n10098) );
  MUX2_X1 U11182 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10098), .S(n10225), .Z(
        P1_U3537) );
  AOI211_X1 U11183 ( .C1(n10211), .C2(n10058), .A(n10057), .B(n10056), .ZN(
        n10059) );
  OAI21_X1 U11184 ( .B1(n10215), .B2(n10060), .A(n10059), .ZN(n10099) );
  MUX2_X1 U11185 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10099), .S(n10225), .Z(
        P1_U3536) );
  AOI211_X1 U11186 ( .C1(n10206), .C2(n10063), .A(n10062), .B(n10061), .ZN(
        n10100) );
  MUX2_X1 U11187 ( .A(n10064), .B(n10100), .S(n10225), .Z(n10065) );
  OAI21_X1 U11188 ( .B1(n10103), .B2(n10066), .A(n10065), .ZN(P1_U3535) );
  INV_X1 U11189 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10068) );
  MUX2_X1 U11190 ( .A(n10068), .B(n10067), .S(n10218), .Z(n10069) );
  OAI21_X1 U11191 ( .B1(n10070), .B2(n10102), .A(n10069), .ZN(P1_U3521) );
  INV_X1 U11192 ( .A(n10075), .ZN(P1_U3520) );
  INV_X1 U11193 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10077) );
  MUX2_X1 U11194 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10079), .S(n10218), .Z(
        P1_U3516) );
  MUX2_X1 U11195 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10081), .S(n10218), .Z(
        P1_U3514) );
  MUX2_X1 U11196 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10082), .S(n10218), .Z(
        P1_U3513) );
  MUX2_X1 U11197 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10083), .S(n10218), .Z(
        P1_U3512) );
  INV_X1 U11198 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10085) );
  MUX2_X1 U11199 ( .A(n10085), .B(n10084), .S(n10218), .Z(n10086) );
  OAI21_X1 U11200 ( .B1(n10087), .B2(n10102), .A(n10086), .ZN(P1_U3511) );
  MUX2_X1 U11201 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10088), .S(n10218), .Z(
        P1_U3510) );
  INV_X1 U11202 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10090) );
  MUX2_X1 U11203 ( .A(n10090), .B(n10089), .S(n10218), .Z(n10091) );
  OAI21_X1 U11204 ( .B1(n10092), .B2(n10102), .A(n10091), .ZN(P1_U3509) );
  MUX2_X1 U11205 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10093), .S(n10218), .Z(
        P1_U3507) );
  MUX2_X1 U11206 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10094), .S(n10218), .Z(
        P1_U3504) );
  INV_X1 U11207 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10096) );
  MUX2_X1 U11208 ( .A(n10096), .B(n10095), .S(n10218), .Z(n10097) );
  OAI21_X1 U11209 ( .B1(n6854), .B2(n10102), .A(n10097), .ZN(P1_U3501) );
  MUX2_X1 U11210 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10098), .S(n10218), .Z(
        P1_U3498) );
  MUX2_X1 U11211 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10099), .S(n10218), .Z(
        P1_U3495) );
  MUX2_X1 U11212 ( .A(n10340), .B(n10100), .S(n10218), .Z(n10101) );
  OAI21_X1 U11213 ( .B1(n10103), .B2(n10102), .A(n10101), .ZN(P1_U3492) );
  MUX2_X1 U11214 ( .A(P1_D_REG_1__SCAN_IN), .B(n10106), .S(n10182), .Z(
        P1_U3440) );
  MUX2_X1 U11215 ( .A(P1_D_REG_0__SCAN_IN), .B(n10107), .S(n10182), .Z(
        P1_U3439) );
  NOR4_X1 U11216 ( .A1(n10108), .A2(P1_IR_REG_30__SCAN_IN), .A3(n4900), .A4(
        n4410), .ZN(n10109) );
  AOI21_X1 U11217 ( .B1(n10110), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10109), 
        .ZN(n10111) );
  OAI21_X1 U11218 ( .B1(n10112), .B2(n10121), .A(n10111), .ZN(P1_U3324) );
  OAI222_X1 U11219 ( .A1(n10115), .A2(n4410), .B1(n10121), .B2(n10114), .C1(
        n10113), .C2(n10118), .ZN(P1_U3327) );
  OAI222_X1 U11220 ( .A1(n10117), .A2(n4410), .B1(n10121), .B2(n10116), .C1(
        n10429), .C2(n10118), .ZN(P1_U3328) );
  OAI222_X1 U11221 ( .A1(n10122), .A2(n4410), .B1(n10121), .B2(n10120), .C1(
        n10119), .C2(n10118), .ZN(P1_U3329) );
  OAI222_X1 U11222 ( .A1(n6856), .A2(n4410), .B1(n10121), .B2(n10124), .C1(
        n10123), .C2(n10118), .ZN(P1_U3330) );
  MUX2_X1 U11223 ( .A(n10125), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  MUX2_X1 U11224 ( .A(n5282), .B(P2_ADDR_REG_19__SCAN_IN), .S(
        P1_ADDR_REG_19__SCAN_IN), .Z(n10156) );
  INV_X1 U11225 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U11226 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10126) );
  AOI21_X1 U11227 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10126), .ZN(n10278) );
  NOR2_X1 U11228 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10127) );
  AOI21_X1 U11229 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10127), .ZN(n10281) );
  NOR2_X1 U11230 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10128) );
  AOI21_X1 U11231 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10128), .ZN(n10284) );
  NOR2_X1 U11232 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10129) );
  AOI21_X1 U11233 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10129), .ZN(n10287) );
  NOR2_X1 U11234 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10130) );
  AOI21_X1 U11235 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10130), .ZN(n10290) );
  INV_X1 U11236 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U11237 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .B1(n10455), .B2(n10131), .ZN(n10293) );
  NOR2_X1 U11238 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10138) );
  XNOR2_X1 U11239 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10601) );
  NAND2_X1 U11240 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10136) );
  XNOR2_X1 U11241 ( .A(n10397), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U11242 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10134) );
  XNOR2_X1 U11243 ( .A(n10132), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(n10597) );
  AOI21_X1 U11244 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10267) );
  NAND3_X1 U11245 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U11246 ( .A1(n10597), .A2(n10596), .ZN(n10133) );
  NAND2_X1 U11247 ( .A1(n10134), .A2(n10133), .ZN(n10598) );
  NAND2_X1 U11248 ( .A1(n10599), .A2(n10598), .ZN(n10135) );
  NAND2_X1 U11249 ( .A1(n10136), .A2(n10135), .ZN(n10600) );
  NOR2_X1 U11250 ( .A1(n10601), .A2(n10600), .ZN(n10137) );
  NOR2_X1 U11251 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10139), .ZN(n10585) );
  NOR2_X1 U11252 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10586), .ZN(n10140) );
  NAND2_X1 U11253 ( .A1(n10141), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10143) );
  XNOR2_X1 U11254 ( .A(n10141), .B(n10439), .ZN(n10588) );
  NAND2_X1 U11255 ( .A1(n10588), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10142) );
  NAND2_X1 U11256 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10144), .ZN(n10146) );
  INV_X1 U11257 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10499) );
  NAND2_X1 U11258 ( .A1(n10593), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U11259 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10147), .ZN(n10149) );
  NAND2_X1 U11260 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10594), .ZN(n10148) );
  NAND2_X1 U11261 ( .A1(n10149), .A2(n10148), .ZN(n10150) );
  AND2_X1 U11262 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n10150), .ZN(n10151) );
  XNOR2_X1 U11263 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n10150), .ZN(n10590) );
  NOR2_X1 U11264 ( .A1(n10591), .A2(n10590), .ZN(n10589) );
  NAND2_X1 U11265 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10152) );
  OAI21_X1 U11266 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10152), .ZN(n10298) );
  NOR2_X1 U11267 ( .A1(n10299), .A2(n10298), .ZN(n10297) );
  AOI21_X1 U11268 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10297), .ZN(n10296) );
  NAND2_X1 U11269 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10153) );
  OAI21_X1 U11270 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10153), .ZN(n10295) );
  NOR2_X1 U11271 ( .A1(n10296), .A2(n10295), .ZN(n10294) );
  NAND2_X1 U11272 ( .A1(n10293), .A2(n10292), .ZN(n10291) );
  NAND2_X1 U11273 ( .A1(n10287), .A2(n10286), .ZN(n10285) );
  NAND2_X1 U11274 ( .A1(n10281), .A2(n10280), .ZN(n10279) );
  OAI21_X1 U11275 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10279), .ZN(n10277) );
  NAND2_X1 U11276 ( .A1(n10278), .A2(n10277), .ZN(n10276) );
  OAI21_X2 U11277 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10276), .ZN(n10273) );
  NAND2_X1 U11278 ( .A1(n10274), .A2(n10273), .ZN(n10154) );
  NOR2_X1 U11279 ( .A1(n10274), .A2(n10273), .ZN(n10272) );
  AOI21_X1 U11280 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10154), .A(n10272), 
        .ZN(n10155) );
  INV_X1 U11281 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10394) );
  XOR2_X1 U11282 ( .A(n10394), .B(P2_WR_REG_SCAN_IN), .Z(U123) );
  INV_X1 U11283 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10523) );
  XOR2_X1 U11284 ( .A(n10523), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  XNOR2_X1 U11285 ( .A(n10157), .B(n10171), .ZN(n10162) );
  AOI222_X1 U11286 ( .A1(n10163), .A2(n10162), .B1(n10161), .B2(n10160), .C1(
        n10159), .C2(n10158), .ZN(n10203) );
  INV_X1 U11287 ( .A(n10164), .ZN(n10165) );
  AOI222_X1 U11288 ( .A1(n10169), .A2(n10168), .B1(P1_REG2_REG_4__SCAN_IN), 
        .B2(n10167), .C1(n10166), .C2(n10165), .ZN(n10181) );
  XOR2_X1 U11289 ( .A(n10170), .B(n10171), .Z(n10207) );
  INV_X1 U11290 ( .A(n10172), .ZN(n10176) );
  INV_X1 U11291 ( .A(n10173), .ZN(n10175) );
  OAI211_X1 U11292 ( .C1(n10202), .C2(n10176), .A(n10175), .B(n10174), .ZN(
        n10200) );
  INV_X1 U11293 ( .A(n10200), .ZN(n10177) );
  AOI22_X1 U11294 ( .A1(n10207), .A2(n10179), .B1(n10178), .B2(n10177), .ZN(
        n10180) );
  OAI211_X1 U11295 ( .C1(n10167), .C2(n10203), .A(n10181), .B(n10180), .ZN(
        P1_U3289) );
  AND2_X1 U11296 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10183), .ZN(P1_U3294) );
  INV_X1 U11297 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10424) );
  NOR2_X1 U11298 ( .A1(n10182), .A2(n10424), .ZN(P1_U3295) );
  AND2_X1 U11299 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10183), .ZN(P1_U3296) );
  AND2_X1 U11300 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10183), .ZN(P1_U3297) );
  AND2_X1 U11301 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10183), .ZN(P1_U3298) );
  AND2_X1 U11302 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10183), .ZN(P1_U3299) );
  AND2_X1 U11303 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10183), .ZN(P1_U3300) );
  AND2_X1 U11304 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10183), .ZN(P1_U3301) );
  AND2_X1 U11305 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10183), .ZN(P1_U3302) );
  AND2_X1 U11306 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10183), .ZN(P1_U3303) );
  AND2_X1 U11307 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10183), .ZN(P1_U3304) );
  AND2_X1 U11308 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10183), .ZN(P1_U3305) );
  AND2_X1 U11309 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10183), .ZN(P1_U3306) );
  INV_X1 U11310 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10481) );
  NOR2_X1 U11311 ( .A1(n10182), .A2(n10481), .ZN(P1_U3307) );
  AND2_X1 U11312 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10183), .ZN(P1_U3308) );
  AND2_X1 U11313 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10183), .ZN(P1_U3309) );
  AND2_X1 U11314 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10183), .ZN(P1_U3310) );
  AND2_X1 U11315 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10183), .ZN(P1_U3311) );
  INV_X1 U11316 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10416) );
  NOR2_X1 U11317 ( .A1(n10182), .A2(n10416), .ZN(P1_U3312) );
  INV_X1 U11318 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10427) );
  NOR2_X1 U11319 ( .A1(n10182), .A2(n10427), .ZN(P1_U3313) );
  INV_X1 U11320 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10540) );
  NOR2_X1 U11321 ( .A1(n10182), .A2(n10540), .ZN(P1_U3314) );
  AND2_X1 U11322 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10183), .ZN(P1_U3315) );
  AND2_X1 U11323 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10183), .ZN(P1_U3316) );
  AND2_X1 U11324 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10183), .ZN(P1_U3317) );
  INV_X1 U11325 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10532) );
  NOR2_X1 U11326 ( .A1(n10182), .A2(n10532), .ZN(P1_U3318) );
  INV_X1 U11327 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10382) );
  NOR2_X1 U11328 ( .A1(n10182), .A2(n10382), .ZN(P1_U3319) );
  AND2_X1 U11329 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10183), .ZN(P1_U3320) );
  AND2_X1 U11330 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10183), .ZN(P1_U3321) );
  AND2_X1 U11331 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10183), .ZN(P1_U3322) );
  AND2_X1 U11332 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10183), .ZN(P1_U3323) );
  INV_X1 U11333 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U11334 ( .A1(n10218), .A2(n10185), .B1(n10184), .B2(n10217), .ZN(
        P1_U3453) );
  AOI21_X1 U11335 ( .B1(n10211), .B2(n7062), .A(n10186), .ZN(n10187) );
  OAI211_X1 U11336 ( .C1(n10190), .C2(n10189), .A(n10188), .B(n10187), .ZN(
        n10191) );
  INV_X1 U11337 ( .A(n10191), .ZN(n10219) );
  INV_X1 U11338 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U11339 ( .A1(n10218), .A2(n10219), .B1(n10192), .B2(n10217), .ZN(
        P1_U3456) );
  AOI22_X1 U11340 ( .A1(n10218), .A2(n10193), .B1(n6264), .B2(n10217), .ZN(
        P1_U3459) );
  OAI21_X1 U11341 ( .B1(n10195), .B2(n10201), .A(n10194), .ZN(n10196) );
  AOI21_X1 U11342 ( .B1(n10197), .B2(n10206), .A(n10196), .ZN(n10198) );
  AND2_X1 U11343 ( .A1(n10199), .A2(n10198), .ZN(n10220) );
  AOI22_X1 U11344 ( .A1(n10218), .A2(n10220), .B1(n6283), .B2(n10217), .ZN(
        P1_U3462) );
  OAI21_X1 U11345 ( .B1(n10202), .B2(n10201), .A(n10200), .ZN(n10205) );
  INV_X1 U11346 ( .A(n10203), .ZN(n10204) );
  AOI211_X1 U11347 ( .C1(n10207), .C2(n10206), .A(n10205), .B(n10204), .ZN(
        n10221) );
  INV_X1 U11348 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U11349 ( .A1(n10218), .A2(n10221), .B1(n10208), .B2(n10217), .ZN(
        P1_U3465) );
  AOI21_X1 U11350 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(n10212) );
  OAI211_X1 U11351 ( .C1(n10215), .C2(n10214), .A(n10213), .B(n10212), .ZN(
        n10216) );
  INV_X1 U11352 ( .A(n10216), .ZN(n10224) );
  AOI22_X1 U11353 ( .A1(n10218), .A2(n10224), .B1(n6302), .B2(n10217), .ZN(
        P1_U3471) );
  AOI22_X1 U11354 ( .A1(n10225), .A2(n10219), .B1(n9629), .B2(n10222), .ZN(
        P1_U3523) );
  AOI22_X1 U11355 ( .A1(n10225), .A2(n10220), .B1(n7424), .B2(n10222), .ZN(
        P1_U3525) );
  AOI22_X1 U11356 ( .A1(n10225), .A2(n10221), .B1(n7425), .B2(n10222), .ZN(
        P1_U3526) );
  AOI22_X1 U11357 ( .A1(n10225), .A2(n10224), .B1(n10223), .B2(n10222), .ZN(
        P1_U3528) );
  OAI22_X1 U11358 ( .A1(n10226), .A2(n10243), .B1(n5184), .B2(n10241), .ZN(
        n10228) );
  NOR2_X1 U11359 ( .A1(n10228), .A2(n10227), .ZN(n10257) );
  AOI22_X1 U11360 ( .A1(n10255), .A2(n5299), .B1(n10257), .B2(n10254), .ZN(
        P2_U3393) );
  INV_X1 U11361 ( .A(n10229), .ZN(n10233) );
  INV_X1 U11362 ( .A(n10230), .ZN(n10231) );
  AOI211_X1 U11363 ( .C1(n10234), .C2(n10233), .A(n10232), .B(n10231), .ZN(
        n10259) );
  AOI22_X1 U11364 ( .A1(n10255), .A2(n5271), .B1(n10259), .B2(n10254), .ZN(
        P2_U3396) );
  INV_X1 U11365 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10239) );
  NOR2_X1 U11366 ( .A1(n10235), .A2(n10243), .ZN(n10237) );
  AOI211_X1 U11367 ( .C1(n10249), .C2(n10238), .A(n10237), .B(n10236), .ZN(
        n10261) );
  AOI22_X1 U11368 ( .A1(n10255), .A2(n10239), .B1(n10261), .B2(n10254), .ZN(
        P2_U3405) );
  INV_X1 U11369 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10247) );
  INV_X1 U11370 ( .A(n10240), .ZN(n10246) );
  OAI22_X1 U11371 ( .A1(n10244), .A2(n10243), .B1(n10242), .B2(n10241), .ZN(
        n10245) );
  NOR2_X1 U11372 ( .A1(n10246), .A2(n10245), .ZN(n10263) );
  AOI22_X1 U11373 ( .A1(n10255), .A2(n10247), .B1(n10263), .B2(n10254), .ZN(
        P2_U3411) );
  AOI22_X1 U11374 ( .A1(n10251), .A2(n10250), .B1(n10249), .B2(n10248), .ZN(
        n10252) );
  AOI22_X1 U11375 ( .A1(n10255), .A2(n5441), .B1(n10265), .B2(n10254), .ZN(
        P2_U3414) );
  AOI22_X1 U11376 ( .A1(n10266), .A2(n10257), .B1(n10256), .B2(n6909), .ZN(
        P2_U3460) );
  AOI22_X1 U11377 ( .A1(n10266), .A2(n10259), .B1(n10258), .B2(n6909), .ZN(
        P2_U3461) );
  AOI22_X1 U11378 ( .A1(n10266), .A2(n10261), .B1(n10260), .B2(n6909), .ZN(
        P2_U3464) );
  AOI22_X1 U11379 ( .A1(n10266), .A2(n10263), .B1(n10262), .B2(n6909), .ZN(
        P2_U3466) );
  INV_X1 U11380 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U11381 ( .A1(n10266), .A2(n10265), .B1(n10264), .B2(n6909), .ZN(
        P2_U3467) );
  INV_X1 U11382 ( .A(n10267), .ZN(n10268) );
  NAND2_X1 U11383 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  XOR2_X1 U11384 ( .A(n10271), .B(n10270), .Z(ADD_1068_U5) );
  XOR2_X1 U11385 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11386 ( .B1(n10274), .B2(n10273), .A(n10272), .ZN(n10275) );
  OAI21_X1 U11387 ( .B1(n10278), .B2(n10277), .A(n10276), .ZN(ADD_1068_U56) );
  OAI21_X1 U11388 ( .B1(n10281), .B2(n10280), .A(n10279), .ZN(ADD_1068_U57) );
  OAI21_X1 U11389 ( .B1(n10284), .B2(n10283), .A(n10282), .ZN(ADD_1068_U58) );
  OAI21_X1 U11390 ( .B1(n10287), .B2(n10286), .A(n10285), .ZN(ADD_1068_U59) );
  OAI21_X1 U11391 ( .B1(n10290), .B2(n10289), .A(n10288), .ZN(ADD_1068_U60) );
  OAI21_X1 U11392 ( .B1(n10293), .B2(n10292), .A(n10291), .ZN(ADD_1068_U61) );
  AOI21_X1 U11393 ( .B1(n10296), .B2(n10295), .A(n10294), .ZN(ADD_1068_U62) );
  AOI21_X1 U11394 ( .B1(n10299), .B2(n10298), .A(n10297), .ZN(ADD_1068_U63) );
  INV_X1 U11395 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10595) );
  NOR4_X1 U11396 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .A3(P1_ADDR_REG_3__SCAN_IN), .A4(n10595), .ZN(n10308) );
  INV_X1 U11397 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10592) );
  NOR4_X1 U11398 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .A3(n9651), .A4(n10592), .ZN(n10300) );
  NAND3_X1 U11399 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), 
        .A3(n10300), .ZN(n10306) );
  NOR4_X1 U11400 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(P1_REG3_REG_5__SCAN_IN), 
        .A3(n10526), .A4(n10525), .ZN(n10302) );
  NOR4_X1 U11401 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n7782), .A3(n10543), .A4(
        n10544), .ZN(n10301) );
  NAND4_X1 U11402 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10305) );
  NOR4_X1 U11403 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10541), .A3(n10306), .A4(
        n10305), .ZN(n10307) );
  NAND4_X1 U11404 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(n10309), .A3(n10308), .A4(
        n10307), .ZN(n10356) );
  NOR4_X1 U11405 ( .A1(n10310), .A2(SI_10_), .A3(P2_REG0_REG_26__SCAN_IN), 
        .A4(P1_REG2_REG_8__SCAN_IN), .ZN(n10314) );
  INV_X1 U11406 ( .A(SI_12_), .ZN(n10473) );
  NOR4_X1 U11407 ( .A1(SI_15_), .A2(P2_DATAO_REG_13__SCAN_IN), .A3(
        P2_REG0_REG_24__SCAN_IN), .A4(n10473), .ZN(n10312) );
  NOR4_X1 U11408 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n10471), .A3(n10469), 
        .A4(n6313), .ZN(n10311) );
  AND4_X1 U11409 ( .A1(n10274), .A2(P2_REG1_REG_29__SCAN_IN), .A3(n10312), 
        .A4(n10311), .ZN(n10313) );
  NAND4_X1 U11410 ( .A1(n10314), .A2(P1_REG2_REG_1__SCAN_IN), .A3(
        P2_DATAO_REG_2__SCAN_IN), .A4(n10313), .ZN(n10355) );
  NOR4_X1 U11411 ( .A1(P2_REG0_REG_1__SCAN_IN), .A2(P1_REG1_REG_18__SCAN_IN), 
        .A3(n6997), .A4(n5423), .ZN(n10320) );
  NOR4_X1 U11412 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(P2_RD_REG_SCAN_IN), .A3(
        n5457), .A4(n10532), .ZN(n10319) );
  NOR4_X1 U11413 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_2__SCAN_IN), 
        .A3(P1_REG2_REG_9__SCAN_IN), .A4(n10315), .ZN(n10316) );
  NAND3_X1 U11414 ( .A1(n10566), .A2(P1_REG1_REG_2__SCAN_IN), .A3(n10316), 
        .ZN(n10317) );
  NOR3_X1 U11415 ( .A1(n10317), .A2(n10565), .A3(P1_REG0_REG_9__SCAN_IN), .ZN(
        n10318) );
  NAND3_X1 U11416 ( .A1(n10320), .A2(n10319), .A3(n10318), .ZN(n10354) );
  NAND4_X1 U11417 ( .A1(P1_REG2_REG_29__SCAN_IN), .A2(n10495), .A3(n4666), 
        .A4(n8517), .ZN(n10329) );
  NOR4_X1 U11418 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_B_REG_SCAN_IN), .A3(
        P1_DATAO_REG_18__SCAN_IN), .A4(n10442), .ZN(n10323) );
  NOR4_X1 U11419 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(P2_REG1_REG_22__SCAN_IN), 
        .A3(n10453), .A4(n10455), .ZN(n10322) );
  AND4_X1 U11420 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(SI_2_), .A3(
        P2_REG0_REG_19__SCAN_IN), .A4(P2_REG2_REG_5__SCAN_IN), .ZN(n10321) );
  AND4_X1 U11421 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(n10323), .A3(n10322), 
        .A4(n10321), .ZN(n10326) );
  NOR2_X1 U11422 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(SI_17_), .ZN(n10325) );
  NOR2_X1 U11423 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(P1_DATAO_REG_8__SCAN_IN), 
        .ZN(n10324) );
  NAND4_X1 U11424 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(
        P2_DATAO_REG_27__SCAN_IN), .ZN(n10328) );
  NAND4_X1 U11425 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), 
        .A3(P1_REG1_REG_14__SCAN_IN), .A4(n10362), .ZN(n10327) );
  NOR3_X1 U11426 ( .A1(n10329), .A2(n10328), .A3(n10327), .ZN(n10348) );
  NAND4_X1 U11427 ( .A1(n10371), .A2(n10330), .A3(n10396), .A4(
        P1_DATAO_REG_0__SCAN_IN), .ZN(n10333) );
  NAND4_X1 U11428 ( .A1(n10331), .A2(n10386), .A3(P2_REG2_REG_17__SCAN_IN), 
        .A4(P2_REG2_REG_0__SCAN_IN), .ZN(n10332) );
  NOR2_X1 U11429 ( .A1(n10333), .A2(n10332), .ZN(n10347) );
  INV_X1 U11430 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10334) );
  NAND4_X1 U11431 ( .A1(n6299), .A2(n10335), .A3(n10334), .A4(n10498), .ZN(
        n10339) );
  NAND4_X1 U11432 ( .A1(n10337), .A2(n10336), .A3(P1_IR_REG_21__SCAN_IN), .A4(
        P1_IR_REG_26__SCAN_IN), .ZN(n10338) );
  NOR2_X1 U11433 ( .A1(n10339), .A2(n10338), .ZN(n10346) );
  NAND4_X1 U11434 ( .A1(SI_0_), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(n6264), .ZN(n10344) );
  NAND4_X1 U11435 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(SI_19_), .A3(
        P1_REG0_REG_15__SCAN_IN), .A4(P1_WR_REG_SCAN_IN), .ZN(n10343) );
  NAND4_X1 U11436 ( .A1(n10341), .A2(n10340), .A3(P1_REG1_REG_26__SCAN_IN), 
        .A4(P1_REG3_REG_28__SCAN_IN), .ZN(n10342) );
  NOR3_X1 U11437 ( .A1(n10344), .A2(n10343), .A3(n10342), .ZN(n10345) );
  AND4_X1 U11438 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10352) );
  INV_X1 U11439 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10388) );
  NOR4_X1 U11440 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(P1_REG2_REG_27__SCAN_IN), 
        .A3(n10388), .A4(n6082), .ZN(n10351) );
  NAND4_X1 U11441 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(P1_REG1_REG_29__SCAN_IN), 
        .A3(P2_ADDR_REG_13__SCAN_IN), .A4(n7424), .ZN(n10349) );
  NOR3_X1 U11442 ( .A1(SI_16_), .A2(n5342), .A3(n10349), .ZN(n10350) );
  NAND3_X1 U11443 ( .A1(n10352), .A2(n10351), .A3(n10350), .ZN(n10353) );
  NOR4_X1 U11444 ( .A1(n10356), .A2(n10355), .A3(n10354), .A4(n10353), .ZN(
        n10583) );
  AOI22_X1 U11445 ( .A1(n10359), .A2(keyinput86), .B1(n10358), .B2(keyinput104), .ZN(n10357) );
  OAI221_X1 U11446 ( .B1(n10359), .B2(keyinput86), .C1(n10358), .C2(
        keyinput104), .A(n10357), .ZN(n10369) );
  AOI22_X1 U11447 ( .A1(n10362), .A2(keyinput64), .B1(n10361), .B2(keyinput66), 
        .ZN(n10360) );
  OAI221_X1 U11448 ( .B1(n10362), .B2(keyinput64), .C1(n10361), .C2(keyinput66), .A(n10360), .ZN(n10368) );
  XOR2_X1 U11449 ( .A(n10331), .B(keyinput120), .Z(n10366) );
  XNOR2_X1 U11450 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput53), .ZN(n10365) );
  XNOR2_X1 U11451 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput6), .ZN(n10364) );
  XNOR2_X1 U11452 ( .A(P1_REG3_REG_28__SCAN_IN), .B(keyinput117), .ZN(n10363)
         );
  NAND4_X1 U11453 ( .A1(n10366), .A2(n10365), .A3(n10364), .A4(n10363), .ZN(
        n10367) );
  NOR3_X1 U11454 ( .A1(n10369), .A2(n10368), .A3(n10367), .ZN(n10408) );
  AOI22_X1 U11455 ( .A1(n5342), .A2(keyinput30), .B1(keyinput38), .B2(n7424), 
        .ZN(n10370) );
  OAI221_X1 U11456 ( .B1(n5342), .B2(keyinput30), .C1(n7424), .C2(keyinput38), 
        .A(n10370), .ZN(n10379) );
  XNOR2_X1 U11457 ( .A(n10371), .B(keyinput63), .ZN(n10378) );
  XOR2_X1 U11458 ( .A(SI_16_), .B(keyinput123), .Z(n10377) );
  XNOR2_X1 U11459 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(keyinput56), .ZN(n10375)
         );
  XNOR2_X1 U11460 ( .A(SI_5_), .B(keyinput96), .ZN(n10374) );
  XNOR2_X1 U11461 ( .A(P2_REG0_REG_23__SCAN_IN), .B(keyinput126), .ZN(n10373)
         );
  XNOR2_X1 U11462 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput82), .ZN(n10372) );
  NAND4_X1 U11463 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        n10376) );
  NOR4_X1 U11464 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10407) );
  AOI22_X1 U11465 ( .A1(n10382), .A2(keyinput21), .B1(keyinput49), .B2(n10381), 
        .ZN(n10380) );
  OAI221_X1 U11466 ( .B1(n10382), .B2(keyinput21), .C1(n10381), .C2(keyinput49), .A(n10380), .ZN(n10392) );
  INV_X1 U11467 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U11468 ( .A1(n8629), .A2(keyinput95), .B1(keyinput72), .B2(n10384), 
        .ZN(n10383) );
  OAI221_X1 U11469 ( .B1(n8629), .B2(keyinput95), .C1(n10384), .C2(keyinput72), 
        .A(n10383), .ZN(n10391) );
  AOI22_X1 U11470 ( .A1(n10386), .A2(keyinput11), .B1(n4743), .B2(keyinput88), 
        .ZN(n10385) );
  OAI221_X1 U11471 ( .B1(n10386), .B2(keyinput11), .C1(n4743), .C2(keyinput88), 
        .A(n10385), .ZN(n10390) );
  AOI22_X1 U11472 ( .A1(n10388), .A2(keyinput103), .B1(keyinput34), .B2(n6082), 
        .ZN(n10387) );
  OAI221_X1 U11473 ( .B1(n10388), .B2(keyinput103), .C1(n6082), .C2(keyinput34), .A(n10387), .ZN(n10389) );
  NOR4_X1 U11474 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10406) );
  AOI22_X1 U11475 ( .A1(n10341), .A2(keyinput94), .B1(keyinput101), .B2(n10394), .ZN(n10393) );
  OAI221_X1 U11476 ( .B1(n10341), .B2(keyinput94), .C1(n10394), .C2(
        keyinput101), .A(n10393), .ZN(n10404) );
  AOI22_X1 U11477 ( .A1(n10397), .A2(keyinput67), .B1(n10396), .B2(keyinput45), 
        .ZN(n10395) );
  OAI221_X1 U11478 ( .B1(n10397), .B2(keyinput67), .C1(n10396), .C2(keyinput45), .A(n10395), .ZN(n10403) );
  XOR2_X1 U11479 ( .A(n9817), .B(keyinput70), .Z(n10401) );
  XNOR2_X1 U11480 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput9), .ZN(n10400) );
  XNOR2_X1 U11481 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput13), .ZN(n10399)
         );
  XNOR2_X1 U11482 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput116), .ZN(n10398)
         );
  NAND4_X1 U11483 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10402) );
  NOR3_X1 U11484 ( .A1(n10404), .A2(n10403), .A3(n10402), .ZN(n10405) );
  NAND4_X1 U11485 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10580) );
  AOI22_X1 U11486 ( .A1(n10411), .A2(keyinput12), .B1(n10410), .B2(keyinput93), 
        .ZN(n10409) );
  OAI221_X1 U11487 ( .B1(n10411), .B2(keyinput12), .C1(n10410), .C2(keyinput93), .A(n10409), .ZN(n10422) );
  INV_X1 U11488 ( .A(SI_0_), .ZN(n10413) );
  AOI22_X1 U11489 ( .A1(n5644), .A2(keyinput62), .B1(keyinput91), .B2(n10413), 
        .ZN(n10412) );
  OAI221_X1 U11490 ( .B1(n5644), .B2(keyinput62), .C1(n10413), .C2(keyinput91), 
        .A(n10412), .ZN(n10421) );
  AOI22_X1 U11491 ( .A1(n10416), .A2(keyinput89), .B1(n10415), .B2(keyinput112), .ZN(n10414) );
  OAI221_X1 U11492 ( .B1(n10416), .B2(keyinput89), .C1(n10415), .C2(
        keyinput112), .A(n10414), .ZN(n10420) );
  AOI22_X1 U11493 ( .A1(n10418), .A2(keyinput27), .B1(keyinput73), .B2(n6264), 
        .ZN(n10417) );
  OAI221_X1 U11494 ( .B1(n10418), .B2(keyinput27), .C1(n6264), .C2(keyinput73), 
        .A(n10417), .ZN(n10419) );
  NOR4_X1 U11495 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n10466) );
  AOI22_X1 U11496 ( .A1(n10425), .A2(keyinput125), .B1(keyinput107), .B2(
        n10424), .ZN(n10423) );
  OAI221_X1 U11497 ( .B1(n10425), .B2(keyinput125), .C1(n10424), .C2(
        keyinput107), .A(n10423), .ZN(n10436) );
  AOI22_X1 U11498 ( .A1(n10427), .A2(keyinput57), .B1(n5593), .B2(keyinput51), 
        .ZN(n10426) );
  OAI221_X1 U11499 ( .B1(n10427), .B2(keyinput57), .C1(n5593), .C2(keyinput51), 
        .A(n10426), .ZN(n10435) );
  AOI22_X1 U11500 ( .A1(n10430), .A2(keyinput97), .B1(n10429), .B2(keyinput25), 
        .ZN(n10428) );
  OAI221_X1 U11501 ( .B1(n10430), .B2(keyinput97), .C1(n10429), .C2(keyinput25), .A(n10428), .ZN(n10434) );
  XNOR2_X1 U11502 ( .A(P1_REG1_REG_26__SCAN_IN), .B(keyinput36), .ZN(n10432)
         );
  XNOR2_X1 U11503 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput19), .ZN(n10431) );
  NAND2_X1 U11504 ( .A1(n10432), .A2(n10431), .ZN(n10433) );
  NOR4_X1 U11505 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n10465) );
  AOI22_X1 U11506 ( .A1(n10439), .A2(keyinput43), .B1(n4410), .B2(keyinput59), 
        .ZN(n10437) );
  OAI221_X1 U11507 ( .B1(n10439), .B2(keyinput43), .C1(n4410), .C2(keyinput59), 
        .A(n10437), .ZN(n10449) );
  AOI22_X1 U11508 ( .A1(n10442), .A2(keyinput106), .B1(n10441), .B2(
        keyinput121), .ZN(n10440) );
  OAI221_X1 U11509 ( .B1(n10442), .B2(keyinput106), .C1(n10441), .C2(
        keyinput121), .A(n10440), .ZN(n10448) );
  XNOR2_X1 U11510 ( .A(P2_B_REG_SCAN_IN), .B(keyinput87), .ZN(n10446) );
  XNOR2_X1 U11511 ( .A(P1_REG0_REG_13__SCAN_IN), .B(keyinput31), .ZN(n10445)
         );
  XNOR2_X1 U11512 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(keyinput110), .ZN(n10444)
         );
  XNOR2_X1 U11513 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput108), .ZN(n10443) );
  NAND4_X1 U11514 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10447) );
  NOR3_X1 U11515 ( .A1(n10449), .A2(n10448), .A3(n10447), .ZN(n10464) );
  AOI22_X1 U11516 ( .A1(n10451), .A2(keyinput14), .B1(keyinput68), .B2(n10595), 
        .ZN(n10450) );
  OAI221_X1 U11517 ( .B1(n10451), .B2(keyinput14), .C1(n10595), .C2(keyinput68), .A(n10450), .ZN(n10462) );
  AOI22_X1 U11518 ( .A1(n10454), .A2(keyinput1), .B1(keyinput114), .B2(n10453), 
        .ZN(n10452) );
  OAI221_X1 U11519 ( .B1(n10454), .B2(keyinput1), .C1(n10453), .C2(keyinput114), .A(n10452), .ZN(n10461) );
  XOR2_X1 U11520 ( .A(n10455), .B(keyinput22), .Z(n10459) );
  XNOR2_X1 U11521 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput98), .ZN(n10458)
         );
  XNOR2_X1 U11522 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput79), .ZN(n10457) );
  XNOR2_X1 U11523 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput8), .ZN(n10456) );
  NAND4_X1 U11524 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        n10460) );
  NOR3_X1 U11525 ( .A1(n10462), .A2(n10461), .A3(n10460), .ZN(n10463) );
  NAND4_X1 U11526 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10579) );
  AOI22_X1 U11527 ( .A1(n10469), .A2(keyinput78), .B1(n10468), .B2(keyinput85), 
        .ZN(n10467) );
  OAI221_X1 U11528 ( .B1(n10469), .B2(keyinput78), .C1(n10468), .C2(keyinput85), .A(n10467), .ZN(n10479) );
  AOI22_X1 U11529 ( .A1(n10471), .A2(keyinput23), .B1(keyinput81), .B2(n6313), 
        .ZN(n10470) );
  OAI221_X1 U11530 ( .B1(n10471), .B2(keyinput23), .C1(n6313), .C2(keyinput81), 
        .A(n10470), .ZN(n10478) );
  AOI22_X1 U11531 ( .A1(n5587), .A2(keyinput26), .B1(keyinput111), .B2(n10473), 
        .ZN(n10472) );
  OAI221_X1 U11532 ( .B1(n5587), .B2(keyinput26), .C1(n10473), .C2(keyinput111), .A(n10472), .ZN(n10477) );
  AOI22_X1 U11533 ( .A1(n9651), .A2(keyinput52), .B1(n10475), .B2(keyinput118), 
        .ZN(n10474) );
  OAI221_X1 U11534 ( .B1(n9651), .B2(keyinput52), .C1(n10475), .C2(keyinput118), .A(n10474), .ZN(n10476) );
  NOR4_X1 U11535 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10521) );
  AOI22_X1 U11536 ( .A1(n10481), .A2(keyinput127), .B1(keyinput99), .B2(n10591), .ZN(n10480) );
  OAI221_X1 U11537 ( .B1(n10481), .B2(keyinput127), .C1(n10591), .C2(
        keyinput99), .A(n10480), .ZN(n10493) );
  XNOR2_X1 U11538 ( .A(n10482), .B(keyinput74), .ZN(n10485) );
  XNOR2_X1 U11539 ( .A(n10483), .B(keyinput84), .ZN(n10484) );
  NOR2_X1 U11540 ( .A1(n10485), .A2(n10484), .ZN(n10489) );
  XNOR2_X1 U11541 ( .A(keyinput75), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(n10488)
         );
  XNOR2_X1 U11542 ( .A(SI_10_), .B(keyinput113), .ZN(n10487) );
  XNOR2_X1 U11543 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput40), .ZN(n10486) );
  NAND4_X1 U11544 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10492) );
  XNOR2_X1 U11545 ( .A(n10490), .B(keyinput124), .ZN(n10491) );
  NOR3_X1 U11546 ( .A1(n10493), .A2(n10492), .A3(n10491), .ZN(n10520) );
  AOI22_X1 U11547 ( .A1(n10495), .A2(keyinput5), .B1(keyinput18), .B2(n4666), 
        .ZN(n10494) );
  OAI221_X1 U11548 ( .B1(n10495), .B2(keyinput5), .C1(n4666), .C2(keyinput18), 
        .A(n10494), .ZN(n10506) );
  AOI22_X1 U11549 ( .A1(n10498), .A2(keyinput83), .B1(n10497), .B2(keyinput92), 
        .ZN(n10496) );
  OAI221_X1 U11550 ( .B1(n10498), .B2(keyinput83), .C1(n10497), .C2(keyinput92), .A(n10496), .ZN(n10505) );
  XOR2_X1 U11551 ( .A(n10499), .B(keyinput102), .Z(n10503) );
  XNOR2_X1 U11552 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput20), .ZN(n10502) );
  XNOR2_X1 U11553 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput65), .ZN(n10501) );
  XNOR2_X1 U11554 ( .A(P2_REG0_REG_28__SCAN_IN), .B(keyinput50), .ZN(n10500)
         );
  NAND4_X1 U11555 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10504) );
  NOR3_X1 U11556 ( .A1(n10506), .A2(n10505), .A3(n10504), .ZN(n10519) );
  AOI22_X1 U11557 ( .A1(n10592), .A2(keyinput15), .B1(n5560), .B2(keyinput122), 
        .ZN(n10507) );
  OAI221_X1 U11558 ( .B1(n10592), .B2(keyinput15), .C1(n5560), .C2(keyinput122), .A(n10507), .ZN(n10517) );
  AOI22_X1 U11559 ( .A1(n8642), .A2(keyinput4), .B1(n8517), .B2(keyinput109), 
        .ZN(n10508) );
  OAI221_X1 U11560 ( .B1(n8642), .B2(keyinput4), .C1(n8517), .C2(keyinput109), 
        .A(n10508), .ZN(n10516) );
  AOI22_X1 U11561 ( .A1(n10511), .A2(keyinput100), .B1(keyinput37), .B2(n10510), .ZN(n10509) );
  OAI221_X1 U11562 ( .B1(n10511), .B2(keyinput100), .C1(n10510), .C2(
        keyinput37), .A(n10509), .ZN(n10515) );
  XNOR2_X1 U11563 ( .A(SI_2_), .B(keyinput39), .ZN(n10513) );
  XNOR2_X1 U11564 ( .A(keyinput105), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n10512)
         );
  NAND2_X1 U11565 ( .A1(n10513), .A2(n10512), .ZN(n10514) );
  NOR4_X1 U11566 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10518) );
  NAND4_X1 U11567 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10578) );
  AOI22_X1 U11568 ( .A1(n6922), .A2(keyinput48), .B1(n10523), .B2(keyinput28), 
        .ZN(n10522) );
  OAI221_X1 U11569 ( .B1(n6922), .B2(keyinput48), .C1(n10523), .C2(keyinput28), 
        .A(n10522), .ZN(n10530) );
  AOI22_X1 U11570 ( .A1(n10526), .A2(keyinput16), .B1(n10525), .B2(keyinput2), 
        .ZN(n10524) );
  OAI221_X1 U11571 ( .B1(n10526), .B2(keyinput16), .C1(n10525), .C2(keyinput2), 
        .A(n10524), .ZN(n10529) );
  XNOR2_X1 U11572 ( .A(n10527), .B(keyinput76), .ZN(n10528) );
  OR3_X1 U11573 ( .A1(n10530), .A2(n10529), .A3(n10528), .ZN(n10537) );
  AOI22_X1 U11574 ( .A1(n10533), .A2(keyinput60), .B1(keyinput10), .B2(n10532), 
        .ZN(n10531) );
  OAI221_X1 U11575 ( .B1(n10533), .B2(keyinput60), .C1(n10532), .C2(keyinput10), .A(n10531), .ZN(n10536) );
  XNOR2_X1 U11576 ( .A(n10534), .B(keyinput90), .ZN(n10535) );
  NOR3_X1 U11577 ( .A1(n10537), .A2(n10536), .A3(n10535), .ZN(n10576) );
  NAND2_X1 U11578 ( .A1(n9101), .A2(keyinput58), .ZN(n10538) );
  OAI221_X1 U11579 ( .B1(n10582), .B2(keyinput69), .C1(n9101), .C2(keyinput58), 
        .A(n10538), .ZN(n10549) );
  AOI22_X1 U11580 ( .A1(n10541), .A2(keyinput33), .B1(keyinput54), .B2(n10540), 
        .ZN(n10539) );
  OAI221_X1 U11581 ( .B1(n10541), .B2(keyinput33), .C1(n10540), .C2(keyinput54), .A(n10539), .ZN(n10548) );
  AOI22_X1 U11582 ( .A1(n10544), .A2(keyinput42), .B1(n10543), .B2(keyinput7), 
        .ZN(n10542) );
  OAI221_X1 U11583 ( .B1(n10544), .B2(keyinput42), .C1(n10543), .C2(keyinput7), 
        .A(n10542), .ZN(n10547) );
  AOI22_X1 U11584 ( .A1(n9625), .A2(keyinput29), .B1(n7782), .B2(keyinput61), 
        .ZN(n10545) );
  OAI221_X1 U11585 ( .B1(n9625), .B2(keyinput29), .C1(n7782), .C2(keyinput61), 
        .A(n10545), .ZN(n10546) );
  NOR4_X1 U11586 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10575) );
  AOI22_X1 U11587 ( .A1(n10551), .A2(keyinput3), .B1(n6997), .B2(keyinput24), 
        .ZN(n10550) );
  OAI221_X1 U11588 ( .B1(n10551), .B2(keyinput3), .C1(n6997), .C2(keyinput24), 
        .A(n10550), .ZN(n10560) );
  AOI22_X1 U11589 ( .A1(n5299), .A2(keyinput77), .B1(n5423), .B2(keyinput44), 
        .ZN(n10552) );
  OAI221_X1 U11590 ( .B1(n5299), .B2(keyinput77), .C1(n5423), .C2(keyinput44), 
        .A(n10552), .ZN(n10559) );
  AOI22_X1 U11591 ( .A1(n8378), .A2(keyinput35), .B1(n10554), .B2(keyinput41), 
        .ZN(n10553) );
  OAI221_X1 U11592 ( .B1(n8378), .B2(keyinput35), .C1(n10554), .C2(keyinput41), 
        .A(n10553), .ZN(n10558) );
  XNOR2_X1 U11593 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput71), .ZN(n10556)
         );
  XNOR2_X1 U11594 ( .A(P1_REG1_REG_18__SCAN_IN), .B(keyinput46), .ZN(n10555)
         );
  NAND2_X1 U11595 ( .A1(n10556), .A2(n10555), .ZN(n10557) );
  NOR4_X1 U11596 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10574) );
  AOI22_X1 U11597 ( .A1(n5457), .A2(keyinput0), .B1(keyinput47), .B2(n8469), 
        .ZN(n10561) );
  OAI221_X1 U11598 ( .B1(n5457), .B2(keyinput0), .C1(n8469), .C2(keyinput47), 
        .A(n10561), .ZN(n10572) );
  AOI22_X1 U11599 ( .A1(n10563), .A2(keyinput32), .B1(keyinput115), .B2(n6521), 
        .ZN(n10562) );
  OAI221_X1 U11600 ( .B1(n10563), .B2(keyinput32), .C1(n6521), .C2(keyinput115), .A(n10562), .ZN(n10571) );
  AOI22_X1 U11601 ( .A1(n10566), .A2(keyinput17), .B1(keyinput119), .B2(n10565), .ZN(n10564) );
  OAI221_X1 U11602 ( .B1(n10566), .B2(keyinput17), .C1(n10565), .C2(
        keyinput119), .A(n10564), .ZN(n10570) );
  XNOR2_X1 U11603 ( .A(P2_REG2_REG_9__SCAN_IN), .B(keyinput55), .ZN(n10568) );
  XNOR2_X1 U11604 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput80), .ZN(n10567) );
  NAND2_X1 U11605 ( .A1(n10568), .A2(n10567), .ZN(n10569) );
  NOR4_X1 U11606 ( .A1(n10572), .A2(n10571), .A3(n10570), .A4(n10569), .ZN(
        n10573) );
  NAND4_X1 U11607 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n10577) );
  OR4_X1 U11608 ( .A1(n10580), .A2(n10579), .A3(n10578), .A4(n10577), .ZN(
        n10581) );
  AOI221_X1 U11609 ( .B1(n10583), .B2(keyinput69), .C1(n10582), .C2(keyinput69), .A(n10581), .ZN(n10584) );
  XOR2_X1 U11610 ( .A(n4410), .B(n10584), .Z(P1_U3086) );
  NOR2_X1 U11611 ( .A1(n10586), .A2(n10585), .ZN(n10587) );
  XOR2_X1 U11612 ( .A(n10587), .B(P2_ADDR_REG_5__SCAN_IN), .Z(ADD_1068_U51) );
  XOR2_X1 U11613 ( .A(n10588), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  AOI21_X1 U11614 ( .B1(n10591), .B2(n10590), .A(n10589), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11615 ( .A(n10593), .B(n10592), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11616 ( .A(n10595), .B(n10594), .ZN(ADD_1068_U48) );
  XOR2_X1 U11617 ( .A(n10597), .B(n10596), .Z(ADD_1068_U54) );
  XOR2_X1 U11618 ( .A(n10599), .B(n10598), .Z(ADD_1068_U53) );
  XNOR2_X1 U11619 ( .A(n10601), .B(n10600), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4948 ( .A(n6289), .Z(n6606) );
  CLKBUF_X1 U4952 ( .A(n5358), .Z(n5800) );
  CLKBUF_X1 U4968 ( .A(n9903), .Z(n4706) );
  CLKBUF_X1 U4969 ( .A(n5842), .Z(n4411) );
  CLKBUF_X1 U4994 ( .A(n6281), .Z(n6615) );
  OR2_X1 U5174 ( .A1(n8659), .A2(n10215), .ZN(n4599) );
  CLKBUF_X1 U5274 ( .A(n8347), .Z(n4609) );
  INV_X1 U5613 ( .A(n5269), .ZN(n8611) );
  CLKBUF_X2 U5960 ( .A(n8127), .Z(n4413) );
endmodule

