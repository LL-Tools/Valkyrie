

module b14_C_SARLock_k_128_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898;

  MUX2_X1 U2399 ( .A(REG1_REG_28__SCAN_IN), .B(n2764), .S(n4898), .Z(n2760) );
  MUX2_X1 U2400 ( .A(REG0_REG_28__SCAN_IN), .B(n2764), .S(n4886), .Z(n2765) );
  INV_X1 U2402 ( .A(n3483), .ZN(n2984) );
  INV_X1 U2403 ( .A(n3835), .ZN(n3358) );
  NAND2_X1 U2405 ( .A1(n3358), .A2(n4801), .ZN(n3753) );
  INV_X1 U2406 ( .A(n3477), .ZN(n3519) );
  INV_X1 U2407 ( .A(n2885), .ZN(n2156) );
  AND4_X2 U2408 ( .A1(n2303), .A2(n2330), .A3(n2229), .A4(n2166), .ZN(n2542)
         );
  OR2_X1 U2409 ( .A1(n2354), .A2(n2686), .ZN(n2372) );
  INV_X1 U2410 ( .A(n3092), .ZN(n3083) );
  INV_X2 U2411 ( .A(n2156), .ZN(n2158) );
  INV_X1 U2412 ( .A(n2156), .ZN(n2159) );
  CLKBUF_X3 U2413 ( .A(n2383), .Z(n3666) );
  INV_X1 U2414 ( .A(n4793), .ZN(n3053) );
  NAND2_X1 U2415 ( .A1(n2542), .A2(n2170), .ZN(n2700) );
  INV_X1 U2416 ( .A(IR_REG_31__SCAN_IN), .ZN(n2686) );
  NAND2_X1 U2417 ( .A1(n2886), .A2(REG2_REG_3__SCAN_IN), .ZN(n2379) );
  OAI21_X1 U2418 ( .B1(n4301), .B2(n3717), .A(n3715), .ZN(n4288) );
  NAND4_X2 U2419 ( .A1(n2382), .A2(n2381), .A3(n2380), .A4(n2379), .ZN(n3835)
         );
  XNOR2_X1 U2420 ( .A(n2755), .B(n3698), .ZN(n3423) );
  XNOR2_X1 U2421 ( .A(n2372), .B(IR_REG_2__SCAN_IN), .ZN(n4647) );
  NAND2_X1 U2422 ( .A1(n2354), .A2(n2328), .ZN(n2384) );
  INV_X1 U2423 ( .A(n2156), .ZN(n2157) );
  NAND2_X1 U2424 ( .A1(n2157), .A2(REG1_REG_3__SCAN_IN), .ZN(n2380) );
  AND2_X2 U2425 ( .A1(n2779), .A2(n2350), .ZN(n2378) );
  INV_X1 U2426 ( .A(n4647), .ZN(n2160) );
  INV_X1 U2427 ( .A(n2160), .ZN(n2161) );
  AOI21_X2 U2428 ( .B1(n4216), .B2(n2609), .A(n2608), .ZN(n4200) );
  AOI21_X2 U2429 ( .B1(n4228), .B2(n2601), .A(n2189), .ZN(n4216) );
  NAND2_X1 U2430 ( .A1(n2212), .A2(n2213), .ZN(n2755) );
  NAND2_X1 U2431 ( .A1(n4273), .A2(n2586), .ZN(n4261) );
  NAND2_X1 U2432 ( .A1(n4275), .A2(n4274), .ZN(n4273) );
  NAND2_X1 U2433 ( .A1(n4352), .A2(n2557), .ZN(n4331) );
  OAI21_X1 U2434 ( .B1(n4422), .B2(n3714), .A(n3712), .ZN(n4406) );
  NAND2_X1 U2435 ( .A1(n2495), .A2(n2494), .ZN(n4422) );
  NAND2_X1 U2436 ( .A1(n2656), .A2(n3771), .ZN(n3123) );
  AND2_X1 U2437 ( .A1(n3753), .A2(n3750), .ZN(n4788) );
  NAND2_X1 U2438 ( .A1(n3748), .A2(n3751), .ZN(n2650) );
  NAND2_X1 U2439 ( .A1(n2431), .A2(n2430), .ZN(n3832) );
  NOR2_X1 U2440 ( .A1(n2811), .A2(n2912), .ZN(n4771) );
  NAND4_X1 U2441 ( .A1(n2371), .A2(n2370), .A3(n2369), .A4(n2368), .ZN(n3537)
         );
  NAND2_X1 U2442 ( .A1(n3817), .A2(n2683), .ZN(n4789) );
  INV_X4 U2443 ( .A(n2176), .ZN(n2162) );
  CLKBUF_X3 U2444 ( .A(n2376), .Z(n2887) );
  AND2_X1 U2445 ( .A1(n2359), .A2(REG1_REG_1__SCAN_IN), .ZN(n2347) );
  XNOR2_X1 U2446 ( .A(n2345), .B(IR_REG_29__SCAN_IN), .ZN(n4638) );
  OR2_X1 U2447 ( .A1(n3424), .A2(n2686), .ZN(n2343) );
  XNOR2_X1 U2448 ( .A(n2642), .B(n2637), .ZN(n3878) );
  OAI211_X1 U2449 ( .C1(n2270), .C2(n2269), .A(n2268), .B(n2168), .ZN(n2836)
         );
  AND2_X1 U2450 ( .A1(n2316), .A2(n2407), .ZN(n2229) );
  AND2_X1 U2451 ( .A1(n2305), .A2(n2304), .ZN(n2303) );
  AND2_X1 U2452 ( .A1(n2332), .A2(n2331), .ZN(n2305) );
  INV_X1 U2453 ( .A(IR_REG_6__SCAN_IN), .ZN(n2331) );
  INV_X1 U2454 ( .A(IR_REG_3__SCAN_IN), .ZN(n2385) );
  INV_X1 U2455 ( .A(IR_REG_15__SCAN_IN), .ZN(n2533) );
  NOR2_X1 U2456 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2332)
         );
  NOR2_X2 U2457 ( .A1(n2700), .A2(n2275), .ZN(n2685) );
  NAND2_X2 U2458 ( .A1(n2649), .A2(n3745), .ZN(n2648) );
  NAND2_X1 U2459 ( .A1(n2349), .A2(n2350), .ZN(n2376) );
  INV_X2 U2460 ( .A(n3537), .ZN(n2374) );
  OAI21_X2 U2461 ( .B1(n3123), .B2(n3766), .A(n3764), .ZN(n3254) );
  NOR2_X1 U2462 ( .A1(n3832), .A2(n2436), .ZN(n2461) );
  NAND2_X1 U2463 ( .A1(n3813), .A2(n3746), .ZN(n2980) );
  INV_X1 U2464 ( .A(IR_REG_23__SCAN_IN), .ZN(n4025) );
  AND2_X1 U2465 ( .A1(n2338), .A2(n2309), .ZN(n2308) );
  INV_X1 U2466 ( .A(IR_REG_17__SCAN_IN), .ZN(n2336) );
  INV_X1 U2467 ( .A(IR_REG_9__SCAN_IN), .ZN(n2304) );
  OAI21_X1 U2468 ( .B1(n3524), .B2(n2284), .A(n2283), .ZN(n2282) );
  AND2_X1 U2469 ( .A1(n3517), .A2(n3516), .ZN(n2284) );
  NAND2_X1 U2470 ( .A1(n3524), .A2(n3516), .ZN(n2283) );
  OR2_X1 U2471 ( .A1(n2610), .A2(n3923), .ZN(n2624) );
  AND2_X1 U2472 ( .A1(n2773), .A2(n4639), .ZN(n2706) );
  AND2_X1 U2473 ( .A1(n3679), .A2(n3682), .ZN(n3698) );
  NOR2_X1 U2474 ( .A1(n4859), .A2(n3746), .ZN(n2736) );
  NAND2_X1 U2475 ( .A1(n2721), .A2(n2720), .ZN(n2861) );
  OAI22_X1 U2476 ( .A1(n3430), .A2(D_REG_0__SCAN_IN), .B1(n2723), .B2(n4639), 
        .ZN(n2735) );
  OR2_X1 U2477 ( .A1(n3896), .A2(n3897), .ZN(n3899) );
  NAND2_X1 U2478 ( .A1(n2853), .A2(n4836), .ZN(n3428) );
  NAND2_X1 U2479 ( .A1(n2341), .A2(n2276), .ZN(n2275) );
  INV_X1 U2480 ( .A(IR_REG_27__SCAN_IN), .ZN(n2341) );
  INV_X1 U2481 ( .A(IR_REG_26__SCAN_IN), .ZN(n2276) );
  NOR2_X2 U2482 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2354)
         );
  OR2_X1 U2483 ( .A1(n2931), .A2(n2324), .ZN(n2797) );
  OR2_X1 U2484 ( .A1(n4699), .A2(n3192), .ZN(n3193) );
  AND2_X1 U2485 ( .A1(n3849), .A2(n2254), .ZN(n2253) );
  AND2_X1 U2486 ( .A1(n2258), .A2(REG2_REG_12__SCAN_IN), .ZN(n2254) );
  INV_X1 U2487 ( .A(n2614), .ZN(n2215) );
  OAI21_X1 U2488 ( .B1(n2219), .B2(n2218), .A(n2167), .ZN(n2495) );
  NAND2_X1 U2489 ( .A1(n3833), .A2(n3150), .ZN(n3758) );
  NAND2_X1 U2490 ( .A1(n3053), .A2(n3017), .ZN(n2652) );
  NAND2_X1 U2491 ( .A1(n4793), .A2(n3069), .ZN(n3756) );
  NOR2_X1 U2492 ( .A1(n3899), .A2(n2724), .ZN(n2725) );
  AND2_X1 U2493 ( .A1(n2870), .A2(n3746), .ZN(n2782) );
  INV_X1 U2494 ( .A(IR_REG_28__SCAN_IN), .ZN(n2355) );
  NAND2_X1 U2495 ( .A1(n2707), .A2(n4025), .ZN(n2709) );
  INV_X1 U2496 ( .A(n4466), .ZN(n3803) );
  OR2_X1 U2497 ( .A1(n3375), .A2(n3374), .ZN(n4658) );
  AND2_X1 U2498 ( .A1(n3477), .A2(n2856), .ZN(n3483) );
  AND2_X1 U2499 ( .A1(n2853), .A2(n2852), .ZN(n2176) );
  XNOR2_X1 U2500 ( .A(n2797), .B(n4646), .ZN(n2843) );
  AND2_X1 U2501 ( .A1(n2799), .A2(n4645), .ZN(n2800) );
  OR2_X1 U2502 ( .A1(n2922), .A2(n4892), .ZN(n2240) );
  NAND2_X1 U2503 ( .A1(n3200), .A2(n3199), .ZN(n3201) );
  NAND2_X1 U2504 ( .A1(n3198), .A2(n4643), .ZN(n3199) );
  INV_X1 U2505 ( .A(n3196), .ZN(n3200) );
  NAND2_X1 U2506 ( .A1(n2266), .A2(n3204), .ZN(n3186) );
  INV_X1 U2507 ( .A(n3184), .ZN(n2266) );
  OR2_X1 U2508 ( .A1(n3193), .A2(n4641), .ZN(n2257) );
  NAND2_X1 U2509 ( .A1(n4703), .A2(n2196), .ZN(n3863) );
  INV_X1 U2510 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4651) );
  OR2_X1 U2511 ( .A1(n4742), .A2(n2247), .ZN(n2244) );
  OR2_X1 U2512 ( .A1(n4751), .A2(REG1_REG_16__SCAN_IN), .ZN(n2247) );
  NAND2_X1 U2513 ( .A1(n3872), .A2(n2246), .ZN(n2245) );
  INV_X1 U2514 ( .A(n4751), .ZN(n2246) );
  OR2_X1 U2515 ( .A1(n2624), .A2(n2623), .ZN(n2740) );
  AOI21_X1 U2516 ( .B1(n4288), .B2(n2577), .A(n2186), .ZN(n4275) );
  NAND2_X1 U2517 ( .A1(n4542), .A2(n4546), .ZN(n2211) );
  AND2_X1 U2518 ( .A1(n3668), .A2(n3669), .ZN(n4405) );
  NOR2_X1 U2519 ( .A1(n3105), .A2(n2458), .ZN(n2465) );
  NAND2_X1 U2520 ( .A1(n2647), .A2(n3878), .ZN(n4435) );
  AND2_X1 U2521 ( .A1(n2725), .A2(n3684), .ZN(n3883) );
  NAND2_X1 U2522 ( .A1(n3899), .A2(n3898), .ZN(n4461) );
  AOI21_X1 U2523 ( .B1(n4200), .B2(n2615), .A(n2614), .ZN(n3891) );
  NAND2_X1 U2524 ( .A1(n2873), .A2(n3813), .ZN(n4878) );
  OR2_X1 U2525 ( .A1(n4808), .A2(n2870), .ZN(n4859) );
  OAI21_X1 U2526 ( .B1(n2645), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2707) );
  NAND2_X1 U2527 ( .A1(n2702), .A2(n4639), .ZN(n3430) );
  INV_X1 U2528 ( .A(IR_REG_22__SCAN_IN), .ZN(n2340) );
  XNOR2_X1 U2529 ( .A(n2696), .B(IR_REG_24__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U2530 ( .A1(n2709), .A2(IR_REG_31__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U2531 ( .A1(n2178), .A2(IR_REG_31__SCAN_IN), .ZN(n2642) );
  INV_X1 U2532 ( .A(n2542), .ZN(n2543) );
  AND2_X1 U2533 ( .A1(n2424), .A2(n2331), .ZN(n2432) );
  NOR2_X1 U2534 ( .A1(n2164), .A2(n3664), .ZN(n2278) );
  INV_X1 U2535 ( .A(n3516), .ZN(n2281) );
  NAND2_X1 U2536 ( .A1(n2282), .A2(n2285), .ZN(n2280) );
  NAND2_X1 U2537 ( .A1(n3524), .A2(n2286), .ZN(n2285) );
  INV_X1 U2538 ( .A(n3517), .ZN(n2286) );
  AND2_X1 U2539 ( .A1(n3473), .A2(n3555), .ZN(n2306) );
  INV_X1 U2540 ( .A(n4668), .ZN(n3661) );
  NAND2_X1 U2541 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2269)
         );
  INV_X1 U2542 ( .A(n2354), .ZN(n2268) );
  OAI21_X1 U2543 ( .B1(n2161), .B2(REG2_REG_2__SCAN_IN), .A(n2803), .ZN(n2929)
         );
  INV_X1 U2544 ( .A(n4646), .ZN(n2389) );
  XNOR2_X1 U2545 ( .A(n2799), .B(n4645), .ZN(n2922) );
  OAI21_X1 U2546 ( .B1(n4744), .B2(n2272), .A(n2271), .ZN(n4752) );
  NAND2_X1 U2547 ( .A1(n2274), .A2(n2273), .ZN(n2272) );
  NAND2_X1 U2548 ( .A1(n3858), .A2(n2274), .ZN(n2271) );
  INV_X1 U2549 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2273) );
  NAND2_X1 U2550 ( .A1(n2812), .A2(n4650), .ZN(n4775) );
  INV_X1 U2551 ( .A(n4762), .ZN(n4754) );
  OR2_X1 U2552 ( .A1(n3428), .A2(n2737), .ZN(n4350) );
  OAI21_X1 U2553 ( .B1(n3423), .B2(n4536), .A(n2216), .ZN(n2764) );
  AND2_X1 U2554 ( .A1(n3418), .A2(n2759), .ZN(n2216) );
  INV_X1 U2555 ( .A(n3369), .ZN(n2295) );
  INV_X1 U2556 ( .A(n2484), .ZN(n2218) );
  OR2_X1 U2557 ( .A1(n3730), .A2(n2218), .ZN(n2217) );
  NOR2_X1 U2558 ( .A1(n2373), .A2(n2200), .ZN(n2204) );
  INV_X1 U2559 ( .A(n2375), .ZN(n2200) );
  AND2_X1 U2560 ( .A1(n2410), .A2(n2962), .ZN(n2205) );
  AND2_X1 U2561 ( .A1(n2300), .A2(n2302), .ZN(n2299) );
  OR2_X1 U2562 ( .A1(n3343), .A2(n2301), .ZN(n2300) );
  AND2_X1 U2563 ( .A1(n2980), .A2(n2979), .ZN(n3480) );
  OAI21_X1 U2564 ( .B1(n3344), .B2(n2294), .A(n2292), .ZN(n3375) );
  INV_X1 U2565 ( .A(n2293), .ZN(n2292) );
  OAI21_X1 U2566 ( .B1(n2297), .B2(n2294), .A(n3368), .ZN(n2293) );
  NAND2_X1 U2567 ( .A1(n2296), .A2(n2295), .ZN(n2294) );
  AND2_X1 U2568 ( .A1(n2853), .A2(n2980), .ZN(n3477) );
  INV_X1 U2569 ( .A(n4638), .ZN(n2350) );
  NAND2_X1 U2570 ( .A1(n4729), .A2(n3870), .ZN(n3871) );
  OR2_X1 U2571 ( .A1(n3798), .A2(n3718), .ZN(n4253) );
  NOR2_X1 U2572 ( .A1(n4345), .A2(n3719), .ZN(n2564) );
  AND2_X1 U2573 ( .A1(n2211), .A2(n2192), .ZN(n2210) );
  OR2_X1 U2574 ( .A1(n3130), .A2(n2463), .ZN(n2458) );
  NAND2_X1 U2575 ( .A1(n2655), .A2(n3758), .ZN(n3106) );
  INV_X1 U2576 ( .A(n4456), .ZN(n3897) );
  NOR2_X1 U2577 ( .A1(n4489), .A2(n2585), .ZN(n2231) );
  AND2_X1 U2578 ( .A1(n2234), .A2(n4333), .ZN(n2233) );
  AND2_X1 U2579 ( .A1(n2556), .A2(n4369), .ZN(n2234) );
  AND2_X1 U2580 ( .A1(n2172), .A2(n4564), .ZN(n2228) );
  NAND2_X1 U2581 ( .A1(n2221), .A2(n2163), .ZN(n3116) );
  INV_X1 U2582 ( .A(n3068), .ZN(n2221) );
  NOR2_X1 U2583 ( .A1(n3031), .A2(n3629), .ZN(n2952) );
  INV_X1 U2584 ( .A(IR_REG_25__SCAN_IN), .ZN(n2339) );
  AND2_X1 U2585 ( .A1(n2336), .A2(n2337), .ZN(n2309) );
  INV_X1 U2586 ( .A(IR_REG_18__SCAN_IN), .ZN(n2337) );
  INV_X1 U2587 ( .A(IR_REG_2__SCAN_IN), .ZN(n2328) );
  NAND2_X1 U2588 ( .A1(n2299), .A2(n2301), .ZN(n2296) );
  OR2_X1 U2589 ( .A1(n2299), .A2(n2298), .ZN(n2297) );
  AND2_X1 U2590 ( .A1(n3343), .A2(n2301), .ZN(n2298) );
  OR2_X1 U2591 ( .A1(n2602), .A2(n3560), .ZN(n2610) );
  AND2_X1 U2592 ( .A1(n2587), .A2(REG3_REG_23__SCAN_IN), .ZN(n2595) );
  AOI21_X1 U2593 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2857), .A(n2978), .ZN(n2860)
         );
  NAND2_X1 U2594 ( .A1(n3557), .A2(n3556), .ZN(n2307) );
  AND2_X1 U2595 ( .A1(n2477), .A2(n2468), .ZN(n3249) );
  NAND2_X1 U2596 ( .A1(n2378), .A2(REG2_REG_0__SCAN_IN), .ZN(n2362) );
  NOR2_X1 U2597 ( .A1(n2830), .A2(n2236), .ZN(n2829) );
  NAND2_X1 U2598 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2236) );
  OR2_X1 U2599 ( .A1(n2930), .A2(n2929), .ZN(n2250) );
  AND2_X1 U2600 ( .A1(n2250), .A2(n2803), .ZN(n2805) );
  OR2_X1 U2601 ( .A1(n2843), .A2(n2844), .ZN(n2841) );
  INV_X1 U2602 ( .A(IR_REG_4__SCAN_IN), .ZN(n2329) );
  OR2_X1 U2603 ( .A1(n2809), .A2(n2810), .ZN(n3182) );
  AND2_X1 U2604 ( .A1(n3841), .A2(n2267), .ZN(n3184) );
  NAND2_X1 U2605 ( .A1(n4642), .A2(REG2_REG_7__SCAN_IN), .ZN(n2267) );
  NAND2_X1 U2606 ( .A1(n2243), .A2(n2242), .ZN(n3203) );
  NAND2_X1 U2607 ( .A1(n3201), .A2(REG1_REG_7__SCAN_IN), .ZN(n2242) );
  OAI21_X1 U2608 ( .B1(n3201), .B2(REG1_REG_7__SCAN_IN), .A(n4642), .ZN(n2243)
         );
  INV_X1 U2609 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4040) );
  NAND2_X1 U2610 ( .A1(n4686), .A2(n3207), .ZN(n3209) );
  INV_X1 U2611 ( .A(IR_REG_12__SCAN_IN), .ZN(n2503) );
  INV_X1 U2612 ( .A(IR_REG_11__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U2613 ( .A1(n2173), .A2(n2257), .ZN(n2256) );
  NAND2_X1 U2614 ( .A1(n4714), .A2(n2195), .ZN(n3866) );
  NAND2_X1 U2615 ( .A1(n3851), .A2(n2258), .ZN(n2255) );
  AOI21_X1 U2616 ( .B1(n2253), .B2(n2257), .A(n2174), .ZN(n2252) );
  INV_X1 U2617 ( .A(n4753), .ZN(n2274) );
  NOR2_X1 U2618 ( .A1(n4752), .A2(n3859), .ZN(n4763) );
  NOR2_X1 U2619 ( .A1(n3873), .A2(REG2_REG_17__SCAN_IN), .ZN(n3859) );
  NAND2_X1 U2620 ( .A1(n2786), .A2(n2785), .ZN(n2811) );
  NAND2_X1 U2621 ( .A1(n4763), .A2(n4764), .ZN(n4761) );
  NAND2_X1 U2622 ( .A1(n2185), .A2(n2214), .ZN(n2213) );
  NAND2_X1 U2623 ( .A1(n4200), .A2(n2191), .ZN(n2212) );
  NAND2_X1 U2624 ( .A1(n2215), .A2(n2622), .ZN(n2214) );
  AND2_X1 U2625 ( .A1(n4483), .A2(n4489), .ZN(n2593) );
  OR2_X1 U2626 ( .A1(n2571), .A2(n2570), .ZN(n2578) );
  AND4_X1 U2627 ( .A1(n2576), .A2(n2575), .A3(n2574), .A4(n2573), .ZN(n4305)
         );
  AND4_X1 U2628 ( .A1(n2569), .A2(n2568), .A3(n2567), .A4(n2566), .ZN(n4326)
         );
  AND2_X1 U2629 ( .A1(n2548), .A2(n2547), .ZN(n2558) );
  NAND2_X1 U2630 ( .A1(n2209), .A2(n2207), .ZN(n4376) );
  AOI21_X1 U2631 ( .B1(n2210), .B2(n4405), .A(n2208), .ZN(n2207) );
  NAND2_X1 U2632 ( .A1(n4406), .A2(n2210), .ZN(n2209) );
  NOR2_X1 U2633 ( .A1(n4652), .A2(n4399), .ZN(n2208) );
  INV_X1 U2634 ( .A(DATAI_12_), .ZN(n4086) );
  AND2_X1 U2635 ( .A1(n3742), .A2(n3779), .ZN(n3221) );
  NAND2_X1 U2636 ( .A1(n2219), .A2(n3730), .ZN(n3223) );
  INV_X1 U2637 ( .A(n3364), .ZN(n4412) );
  NAND2_X1 U2638 ( .A1(n2446), .A2(n3106), .ZN(n3130) );
  INV_X1 U2639 ( .A(n2461), .ZN(n2446) );
  OR2_X1 U2640 ( .A1(n2461), .A2(n2460), .ZN(n3131) );
  AND3_X1 U2641 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2418) );
  INV_X1 U2642 ( .A(n3017), .ZN(n3069) );
  MUX2_X1 U2643 ( .A(n2357), .B(n2356), .S(IR_REG_27__SCAN_IN), .Z(n2383) );
  INV_X1 U2644 ( .A(n3536), .ZN(n3021) );
  INV_X1 U2645 ( .A(n3878), .ZN(n4349) );
  INV_X1 U2646 ( .A(n3029), .ZN(n2854) );
  AND2_X1 U2647 ( .A1(n3820), .A2(n3736), .ZN(n2873) );
  NAND2_X1 U2648 ( .A1(n2757), .A2(n4789), .ZN(n3418) );
  NOR2_X1 U2649 ( .A1(n4462), .A2(n2225), .ZN(n2224) );
  NAND2_X1 U2650 ( .A1(n4460), .A2(n4459), .ZN(n2225) );
  AND2_X1 U2651 ( .A1(n4230), .A2(n4223), .ZN(n4218) );
  AND2_X1 U2652 ( .A1(n4289), .A2(n2230), .ZN(n4230) );
  AND2_X1 U2653 ( .A1(n2231), .A2(n4480), .ZN(n2230) );
  NAND2_X1 U2654 ( .A1(n4289), .A2(n2231), .ZN(n4263) );
  INV_X1 U2655 ( .A(n4268), .ZN(n4489) );
  NAND2_X1 U2656 ( .A1(n4289), .A2(n4283), .ZN(n4496) );
  AND4_X1 U2657 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .ZN(n4502)
         );
  INV_X1 U2658 ( .A(n4501), .ZN(n4290) );
  NOR2_X1 U2659 ( .A1(n4311), .A2(n4290), .ZN(n4289) );
  NAND2_X1 U2660 ( .A1(n4377), .A2(n2232), .ZN(n4311) );
  AND2_X1 U2661 ( .A1(n2233), .A2(n4312), .ZN(n2232) );
  NAND2_X1 U2662 ( .A1(n4377), .A2(n2233), .ZN(n4332) );
  NAND2_X1 U2663 ( .A1(n4377), .A2(n2234), .ZN(n4342) );
  NOR2_X1 U2664 ( .A1(n4394), .A2(n4657), .ZN(n4377) );
  AND4_X1 U2665 ( .A1(n2532), .A2(n2531), .A3(n2530), .A4(n2529), .ZN(n4525)
         );
  INV_X1 U2666 ( .A(n4873), .ZN(n4536) );
  OR2_X1 U2667 ( .A1(n4409), .A2(n4538), .ZN(n4394) );
  AND2_X1 U2668 ( .A1(n3247), .A2(n2227), .ZN(n4408) );
  AND2_X1 U2669 ( .A1(n2228), .A2(n4437), .ZN(n2227) );
  NAND2_X1 U2670 ( .A1(n3247), .A2(n2172), .ZN(n3310) );
  INV_X1 U2671 ( .A(n3302), .ZN(n3291) );
  OR2_X1 U2672 ( .A1(n3116), .A2(n2436), .ZN(n3125) );
  NOR2_X1 U2673 ( .A1(n3125), .A2(n3269), .ZN(n3247) );
  NAND2_X1 U2674 ( .A1(n2221), .A2(n2220), .ZN(n3148) );
  NOR2_X1 U2675 ( .A1(n3091), .A2(n3056), .ZN(n2220) );
  NOR2_X1 U2676 ( .A1(n3068), .A2(n3056), .ZN(n3098) );
  INV_X1 U2677 ( .A(n4563), .ZN(n4791) );
  AND2_X1 U2678 ( .A1(n2952), .A2(n2993), .ZN(n4799) );
  NAND2_X1 U2679 ( .A1(n4435), .A2(n4859), .ZN(n4873) );
  NAND2_X1 U2680 ( .A1(n2873), .A2(n4640), .ZN(n4563) );
  INV_X1 U2681 ( .A(n4836), .ZN(n3431) );
  NAND2_X1 U2682 ( .A1(n2685), .A2(n2355), .ZN(n2344) );
  OAI21_X1 U2683 ( .B1(n2700), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2684) );
  INV_X1 U2684 ( .A(n2707), .ZN(n2708) );
  XNOR2_X1 U2685 ( .A(n2640), .B(n2639), .ZN(n3813) );
  NAND2_X1 U2686 ( .A1(n2638), .A2(IR_REG_31__SCAN_IN), .ZN(n2640) );
  INV_X1 U2687 ( .A(IR_REG_19__SCAN_IN), .ZN(n2637) );
  AND2_X1 U2688 ( .A1(n2542), .A2(n2336), .ZN(n2554) );
  AND2_X1 U2689 ( .A1(n2229), .A2(n2330), .ZN(n2424) );
  AOI22_X1 U2690 ( .A1(n2165), .A2(n3137), .B1(n3138), .B2(n2290), .ZN(n2289)
         );
  NAND2_X1 U2691 ( .A1(n2291), .A2(n2296), .ZN(n3370) );
  NAND2_X1 U2692 ( .A1(n3344), .A2(n2297), .ZN(n2291) );
  AND2_X1 U2693 ( .A1(n3455), .A2(n3454), .ZN(n2319) );
  AND4_X1 U2694 ( .A1(n2483), .A2(n2482), .A3(n2481), .A4(n2480), .ZN(n4568)
         );
  AND2_X1 U2695 ( .A1(n3298), .A2(n3289), .ZN(n2287) );
  NAND2_X1 U2696 ( .A1(n3290), .A2(n3289), .ZN(n3296) );
  OAI21_X1 U2697 ( .B1(n3666), .B2(n2389), .A(n2388), .ZN(n4801) );
  NAND2_X1 U2698 ( .A1(n3666), .A2(DATAI_3_), .ZN(n2388) );
  AND4_X1 U2699 ( .A1(n2541), .A2(n2540), .A3(n2539), .A4(n2538), .ZN(n4654)
         );
  INV_X1 U2700 ( .A(n4410), .ZN(n4652) );
  NAND2_X1 U2701 ( .A1(n3052), .A2(n3051), .ZN(n3079) );
  INV_X1 U2702 ( .A(n3832), .ZN(n3267) );
  AND4_X1 U2703 ( .A1(n2489), .A2(n2488), .A3(n2487), .A4(n2486), .ZN(n4431)
         );
  NAND2_X1 U2704 ( .A1(n3344), .A2(n3343), .ZN(n3599) );
  INV_X1 U2705 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U2706 ( .A1(n3079), .A2(n2313), .ZN(n3139) );
  NAND2_X1 U2707 ( .A1(n2307), .A2(n3555), .ZN(n3646) );
  INV_X1 U2708 ( .A(n3652), .ZN(n4656) );
  NAND2_X1 U2709 ( .A1(n2621), .A2(n2620), .ZN(n4466) );
  INV_X1 U2710 ( .A(n4502), .ZN(n4291) );
  INV_X1 U2711 ( .A(n4326), .ZN(n4504) );
  INV_X1 U2712 ( .A(n4654), .ZN(n4529) );
  INV_X1 U2713 ( .A(n4525), .ZN(n4539) );
  NAND2_X1 U2714 ( .A1(n2455), .A2(n2177), .ZN(n3831) );
  NAND3_X1 U2715 ( .A1(n2181), .A2(n2320), .A3(n2444), .ZN(n3833) );
  NAND4_X1 U2716 ( .A1(n2405), .A2(n2404), .A3(n2403), .A4(n2402), .ZN(n3092)
         );
  NAND3_X1 U2717 ( .A1(n2322), .A2(n2397), .A3(n2396), .ZN(n4793) );
  OR2_X1 U2718 ( .A1(n2887), .A2(n2395), .ZN(n2397) );
  CLKBUF_X1 U2719 ( .A(n2364), .Z(n2872) );
  OR2_X1 U2720 ( .A1(n2853), .A2(n3431), .ZN(n3836) );
  INV_X1 U2721 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2802) );
  NOR2_X1 U2722 ( .A1(n2829), .A2(n2235), .ZN(n2933) );
  NOR2_X1 U2723 ( .A1(n2836), .A2(n2794), .ZN(n2235) );
  NOR2_X1 U2724 ( .A1(n2933), .A2(n2932), .ZN(n2931) );
  XNOR2_X1 U2725 ( .A(n2805), .B(n2389), .ZN(n2839) );
  INV_X1 U2726 ( .A(n2240), .ZN(n2921) );
  XNOR2_X1 U2727 ( .A(n2806), .B(n4645), .ZN(n2919) );
  NOR2_X1 U2728 ( .A1(n2919), .A2(n2920), .ZN(n2918) );
  OAI21_X1 U2729 ( .B1(n2922), .B2(n2238), .A(n2237), .ZN(n2818) );
  NAND2_X1 U2730 ( .A1(n2241), .A2(REG1_REG_4__SCAN_IN), .ZN(n2238) );
  NAND2_X1 U2731 ( .A1(n2800), .A2(n2241), .ZN(n2237) );
  INV_X1 U2732 ( .A(n2819), .ZN(n2241) );
  INV_X1 U2733 ( .A(n2800), .ZN(n2239) );
  OAI21_X1 U2734 ( .B1(n2919), .B2(n2264), .A(n2263), .ZN(n2820) );
  NAND2_X1 U2735 ( .A1(n2265), .A2(REG2_REG_4__SCAN_IN), .ZN(n2264) );
  NAND2_X1 U2736 ( .A1(n2318), .A2(n2265), .ZN(n2263) );
  INV_X1 U2737 ( .A(n2821), .ZN(n2265) );
  INV_X1 U2738 ( .A(n3201), .ZN(n3839) );
  XNOR2_X1 U2739 ( .A(n3203), .B(n4855), .ZN(n4678) );
  NAND2_X1 U2740 ( .A1(n4678), .A2(REG1_REG_8__SCAN_IN), .ZN(n4677) );
  INV_X1 U2741 ( .A(n3186), .ZN(n3187) );
  XNOR2_X1 U2742 ( .A(n3209), .B(n4851), .ZN(n4696) );
  NOR2_X1 U2743 ( .A1(n4692), .A2(n3250), .ZN(n4691) );
  OAI21_X1 U2744 ( .B1(n4692), .B2(n2262), .A(n2260), .ZN(n4699) );
  OR2_X1 U2745 ( .A1(n4700), .A2(n3250), .ZN(n2262) );
  NAND2_X1 U2746 ( .A1(n3191), .A2(n2261), .ZN(n2260) );
  INV_X1 U2747 ( .A(n4700), .ZN(n2261) );
  INV_X1 U2748 ( .A(n2256), .ZN(n3850) );
  NAND2_X1 U2749 ( .A1(n3865), .A2(n3864), .ZN(n4715) );
  NAND2_X1 U2750 ( .A1(n4715), .A2(n4716), .ZN(n4714) );
  XNOR2_X1 U2751 ( .A(n3866), .B(n3852), .ZN(n4726) );
  NOR2_X1 U2752 ( .A1(n3824), .A2(n2811), .ZN(n4762) );
  AND3_X1 U2753 ( .A1(n2245), .A2(n2244), .A3(n2175), .ZN(n4772) );
  AOI211_X1 U2754 ( .C1(n4462), .C2(n4815), .A(n3904), .B(n3903), .ZN(n3905)
         );
  NAND2_X1 U2755 ( .A1(n3666), .A2(DATAI_26_), .ZN(n4464) );
  NAND2_X1 U2756 ( .A1(n3666), .A2(DATAI_25_), .ZN(n4223) );
  NAND2_X1 U2757 ( .A1(n3666), .A2(DATAI_21_), .ZN(n4501) );
  INV_X1 U2758 ( .A(n4538), .ZN(n4399) );
  NAND2_X1 U2759 ( .A1(n2206), .A2(n2211), .ZN(n4393) );
  OR2_X1 U2760 ( .A1(n4406), .A2(n4405), .ZN(n2206) );
  INV_X1 U2761 ( .A(n4802), .ZN(n4441) );
  NAND2_X1 U2762 ( .A1(n2738), .A2(n4350), .ZN(n4815) );
  INV_X1 U2763 ( .A(n4350), .ZN(n4810) );
  INV_X1 U2764 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3998) );
  AOI21_X1 U2765 ( .B1(n4450), .B2(n4449), .A(n4448), .ZN(n4670) );
  AOI21_X1 U2766 ( .B1(n2747), .B2(n2761), .A(n3883), .ZN(n2742) );
  NAND2_X1 U2767 ( .A1(n2226), .A2(n2222), .ZN(n4583) );
  INV_X1 U2768 ( .A(n2223), .ZN(n2222) );
  NAND2_X1 U2769 ( .A1(n4463), .A2(n4873), .ZN(n2226) );
  OAI21_X1 U2770 ( .B1(n4461), .B2(n4878), .A(n2224), .ZN(n2223) );
  INV_X1 U2771 ( .A(n4865), .ZN(n4632) );
  NOR2_X1 U2772 ( .A1(n4885), .A2(n4878), .ZN(n4865) );
  NAND2_X1 U2773 ( .A1(n3430), .A2(n3429), .ZN(n4835) );
  MUX2_X1 U2774 ( .A(n2688), .B(n2687), .S(IR_REG_28__SCAN_IN), .Z(n4650) );
  XNOR2_X1 U2775 ( .A(n2701), .B(IR_REG_26__SCAN_IN), .ZN(n4639) );
  NAND2_X1 U2776 ( .A1(n2700), .A2(IR_REG_31__SCAN_IN), .ZN(n2701) );
  INV_X1 U2777 ( .A(n2705), .ZN(n2773) );
  INV_X1 U2778 ( .A(n2723), .ZN(n3432) );
  AND2_X1 U2779 ( .A1(n2974), .A2(STATE_REG_SCAN_IN), .ZN(n4836) );
  XNOR2_X1 U2780 ( .A(n2646), .B(IR_REG_22__SCAN_IN), .ZN(n2870) );
  XNOR2_X1 U2781 ( .A(n2644), .B(n2643), .ZN(n3746) );
  INV_X1 U2782 ( .A(IR_REG_21__SCAN_IN), .ZN(n2643) );
  INV_X1 U2783 ( .A(n3862), .ZN(n4839) );
  INV_X1 U2784 ( .A(n3211), .ZN(n4849) );
  AND2_X1 U2785 ( .A1(n2398), .A2(n2387), .ZN(n4646) );
  INV_X2 U2786 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U2787 ( .A1(n2280), .A2(n4663), .ZN(n2279) );
  AOI211_X1 U2788 ( .C1(ADDR_REG_17__SCAN_IN), .C2(n4767), .A(n4759), .B(n4758), .ZN(n4760) );
  AND3_X1 U2789 ( .A1(n3049), .A2(n3150), .A3(n3097), .ZN(n2163) );
  AND2_X1 U2790 ( .A1(n2282), .A2(n2187), .ZN(n2164) );
  OR2_X1 U2791 ( .A1(n2290), .A2(n3138), .ZN(n2165) );
  AND4_X1 U2792 ( .A1(n2335), .A2(n2334), .A3(n2333), .A4(n2533), .ZN(n2166)
         );
  AND2_X1 U2793 ( .A1(n2217), .A2(n2493), .ZN(n2167) );
  OR2_X1 U2794 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2168)
         );
  AND2_X1 U2795 ( .A1(n2188), .A2(n3051), .ZN(n2169) );
  AND2_X1 U2796 ( .A1(n2308), .A2(n2180), .ZN(n2170) );
  AND2_X1 U2797 ( .A1(n3849), .A2(n2256), .ZN(n2171) );
  INV_X1 U2798 ( .A(n4542), .ZN(n4429) );
  AND4_X1 U2799 ( .A1(n2513), .A2(n2512), .A3(n2511), .A4(n2510), .ZN(n4542)
         );
  AND2_X1 U2800 ( .A1(n3291), .A2(n3335), .ZN(n2172) );
  NAND2_X1 U2801 ( .A1(n4374), .A2(n2190), .ZN(n4363) );
  AND2_X1 U2802 ( .A1(n3849), .A2(REG2_REG_12__SCAN_IN), .ZN(n2173) );
  AND2_X1 U2803 ( .A1(n2259), .A2(n2258), .ZN(n2174) );
  OR2_X1 U2804 ( .A1(n3873), .A2(REG1_REG_17__SCAN_IN), .ZN(n2175) );
  NAND2_X1 U2805 ( .A1(n2542), .A2(n2308), .ZN(n2645) );
  NAND2_X1 U2806 ( .A1(n2706), .A2(n2723), .ZN(n2853) );
  AND3_X1 U2807 ( .A1(n2454), .A2(n2453), .A3(n2452), .ZN(n2177) );
  NAND2_X1 U2808 ( .A1(n2542), .A2(n2309), .ZN(n2178) );
  OR2_X1 U2809 ( .A1(n3835), .A2(n4801), .ZN(n2179) );
  INV_X1 U2810 ( .A(n2836), .ZN(n4648) );
  NAND2_X1 U2811 ( .A1(n2330), .A2(n2316), .ZN(n2406) );
  INV_X1 U2812 ( .A(n2650), .ZN(n2945) );
  AND4_X1 U2813 ( .A1(n2340), .A2(n2695), .A3(n4025), .A4(n2339), .ZN(n2180)
         );
  INV_X1 U2814 ( .A(IR_REG_0__SCAN_IN), .ZN(n2270) );
  NAND2_X1 U2815 ( .A1(n2159), .A2(REG1_REG_7__SCAN_IN), .ZN(n2181) );
  NOR2_X1 U2816 ( .A1(n4743), .A2(n3858), .ZN(n2182) );
  NAND2_X1 U2817 ( .A1(n3831), .A2(n3269), .ZN(n2183) );
  AND2_X1 U2818 ( .A1(n2249), .A2(n2248), .ZN(n2184) );
  NAND2_X1 U2819 ( .A1(n2161), .A2(REG2_REG_2__SCAN_IN), .ZN(n2803) );
  AND2_X1 U2820 ( .A1(n3334), .A2(n3333), .ZN(n3541) );
  INV_X1 U2821 ( .A(n3596), .ZN(n2301) );
  OR2_X1 U2822 ( .A1(n3803), .A2(n4456), .ZN(n2185) );
  AND2_X1 U2823 ( .A1(n4305), .A2(n4501), .ZN(n2186) );
  OR2_X1 U2824 ( .A1(n3524), .A2(n2281), .ZN(n2187) );
  INV_X1 U2825 ( .A(n3204), .ZN(n4855) );
  INV_X1 U2826 ( .A(n2517), .ZN(n4546) );
  NAND2_X1 U2827 ( .A1(n4376), .A2(n4375), .ZN(n4374) );
  OR2_X1 U2828 ( .A1(n3138), .A2(n3137), .ZN(n2188) );
  AND2_X1 U2829 ( .A1(n4476), .A2(n4480), .ZN(n2189) );
  OR2_X1 U2830 ( .A1(n3078), .A2(n3077), .ZN(n2313) );
  INV_X1 U2831 ( .A(n2313), .ZN(n2290) );
  NAND2_X1 U2832 ( .A1(n2424), .A2(n2305), .ZN(n2456) );
  OR2_X1 U2833 ( .A1(n4525), .A2(n4381), .ZN(n2190) );
  AND2_X1 U2834 ( .A1(n2185), .A2(n2615), .ZN(n2191) );
  INV_X1 U2835 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4892) );
  OR2_X1 U2836 ( .A1(n4410), .A2(n4538), .ZN(n2192) );
  INV_X1 U2837 ( .A(n3049), .ZN(n3056) );
  INV_X1 U2838 ( .A(n4564), .ZN(n3311) );
  NAND2_X1 U2839 ( .A1(n2424), .A2(n2303), .ZN(n2473) );
  NOR2_X1 U2840 ( .A1(n4691), .A2(n3191), .ZN(n2193) );
  INV_X1 U2841 ( .A(n4428), .ZN(n4437) );
  OAI21_X1 U2842 ( .B1(n3089), .B2(n2427), .A(n2426), .ZN(n3105) );
  AND2_X1 U2843 ( .A1(n4377), .A2(n4369), .ZN(n4341) );
  AND2_X1 U2844 ( .A1(n3247), .A2(n2228), .ZN(n2194) );
  NAND2_X1 U2845 ( .A1(n3247), .A2(n3291), .ZN(n3224) );
  NAND2_X1 U2846 ( .A1(n2652), .A2(n3756), .ZN(n2962) );
  NAND2_X1 U2847 ( .A1(n2288), .A2(n2289), .ZN(n3168) );
  NAND2_X1 U2848 ( .A1(n3223), .A2(n2484), .ZN(n3308) );
  NAND2_X1 U2849 ( .A1(n3666), .A2(DATAI_22_), .ZN(n4283) );
  XNOR2_X1 U2850 ( .A(n2698), .B(IR_REG_25__SCAN_IN), .ZN(n2705) );
  INV_X1 U2851 ( .A(n3719), .ZN(n4333) );
  OAI22_X1 U2852 ( .A1(n3246), .A2(n2476), .B1(n3617), .B2(n3291), .ZN(n3220)
         );
  OR2_X1 U2853 ( .A1(n4847), .A2(n4559), .ZN(n2195) );
  OR2_X1 U2854 ( .A1(n4849), .A2(n3951), .ZN(n2196) );
  INV_X1 U2855 ( .A(n4708), .ZN(n2259) );
  NAND2_X1 U2856 ( .A1(n3666), .A2(DATAI_24_), .ZN(n4480) );
  NAND2_X1 U2857 ( .A1(n3666), .A2(DATAI_20_), .ZN(n4312) );
  INV_X1 U2858 ( .A(n4388), .ZN(n4407) );
  INV_X2 U2859 ( .A(n4885), .ZN(n4886) );
  NOR2_X1 U2860 ( .A1(n2918), .A2(n2318), .ZN(n2197) );
  INV_X2 U2861 ( .A(n4895), .ZN(n4898) );
  OR2_X1 U2862 ( .A1(n2729), .A2(n2735), .ZN(n4895) );
  AND2_X1 U2863 ( .A1(n2240), .A2(n2239), .ZN(n2198) );
  INV_X1 U2864 ( .A(IR_REG_20__SCAN_IN), .ZN(n2639) );
  NOR2_X1 U2865 ( .A1(n2344), .A2(IR_REG_29__SCAN_IN), .ZN(n3424) );
  NAND2_X1 U2866 ( .A1(n2199), .A2(n2390), .ZN(n2202) );
  NAND2_X1 U2867 ( .A1(n2945), .A2(n2375), .ZN(n2199) );
  NAND2_X1 U2868 ( .A1(n2203), .A2(n2201), .ZN(n2961) );
  NAND2_X1 U2869 ( .A1(n2179), .A2(n2202), .ZN(n2201) );
  NAND2_X1 U2870 ( .A1(n2179), .A2(n2204), .ZN(n2203) );
  NAND2_X1 U2871 ( .A1(n2940), .A2(n2375), .ZN(n4785) );
  NAND2_X1 U2872 ( .A1(n2373), .A2(n2650), .ZN(n2940) );
  NAND2_X1 U2873 ( .A1(n2961), .A2(n2205), .ZN(n2415) );
  INV_X1 U2874 ( .A(n3220), .ZN(n2219) );
  AOI21_X2 U2875 ( .B1(n4261), .B2(n2594), .A(n2593), .ZN(n4228) );
  NAND2_X1 U2876 ( .A1(n2245), .A2(n2244), .ZN(n4750) );
  OR2_X1 U2877 ( .A1(n4742), .A2(REG1_REG_16__SCAN_IN), .ZN(n2249) );
  INV_X1 U2878 ( .A(n2249), .ZN(n4741) );
  INV_X1 U2879 ( .A(n3872), .ZN(n2248) );
  INV_X1 U2880 ( .A(n2250), .ZN(n2928) );
  NOR2_X1 U2881 ( .A1(n2827), .A2(n2251), .ZN(n2930) );
  AND2_X1 U2882 ( .A1(n4648), .A2(REG2_REG_1__SCAN_IN), .ZN(n2251) );
  NAND2_X1 U2883 ( .A1(n2255), .A2(n2252), .ZN(n3853) );
  NAND2_X1 U2884 ( .A1(n2257), .A2(n3849), .ZN(n3194) );
  NAND2_X1 U2885 ( .A1(n4847), .A2(n4000), .ZN(n2258) );
  XNOR2_X1 U2886 ( .A(n3190), .B(n4851), .ZN(n4692) );
  XNOR2_X1 U2887 ( .A(n2836), .B(n2802), .ZN(n2828) );
  NOR2_X1 U2888 ( .A1(n4744), .A2(REG2_REG_16__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U2889 ( .A1(n3518), .A2(n2278), .ZN(n2277) );
  OAI211_X1 U2890 ( .C1(n3518), .C2(n2279), .A(n2277), .B(n3531), .ZN(U3217)
         );
  NAND2_X2 U2891 ( .A1(n3365), .A2(n3536), .ZN(n2649) );
  INV_X2 U2892 ( .A(n2364), .ZN(n3365) );
  NAND2_X1 U2893 ( .A1(n3290), .A2(n2287), .ZN(n3334) );
  NAND2_X1 U2894 ( .A1(n3052), .A2(n2169), .ZN(n2288) );
  INV_X1 U2895 ( .A(n3597), .ZN(n2302) );
  NAND2_X1 U2896 ( .A1(n2307), .A2(n2306), .ZN(n3476) );
  AOI21_X2 U2897 ( .B1(n2751), .B2(n4873), .A(n2694), .ZN(n2732) );
  OAI21_X2 U2898 ( .B1(n3062), .B2(n2653), .A(n3756), .ZN(n2959) );
  OAI21_X2 U2899 ( .B1(n2959), .B2(n2958), .A(n3768), .ZN(n3090) );
  OR2_X1 U2900 ( .A1(n2684), .A2(n2355), .ZN(n2356) );
  AND2_X2 U2901 ( .A1(n2779), .A2(n4638), .ZN(n2392) );
  NOR2_X2 U2902 ( .A1(n2465), .A2(n2464), .ZN(n3246) );
  OR2_X1 U2903 ( .A1(n2376), .A2(n2358), .ZN(n2361) );
  NOR2_X1 U2904 ( .A1(n2376), .A2(n2346), .ZN(n2348) );
  AND2_X2 U2905 ( .A1(n2349), .A2(n4638), .ZN(n2359) );
  INV_X1 U2906 ( .A(n2745), .ZN(n2754) );
  AOI21_X2 U2907 ( .B1(n4331), .B2(n2565), .A(n2564), .ZN(n4301) );
  AND2_X1 U2908 ( .A1(n2858), .A2(n3029), .ZN(n3020) );
  NAND2_X1 U2909 ( .A1(n2344), .A2(IR_REG_31__SCAN_IN), .ZN(n2345) );
  INV_X1 U2910 ( .A(n2349), .ZN(n2779) );
  AND2_X1 U2911 ( .A1(n4769), .A2(n4768), .ZN(n2310) );
  AND2_X1 U2912 ( .A1(n2731), .A2(n2730), .ZN(n2311) );
  AND2_X1 U2913 ( .A1(n2728), .A2(n2727), .ZN(n2312) );
  AND2_X1 U2914 ( .A1(n2158), .A2(REG1_REG_8__SCAN_IN), .ZN(n2314) );
  INV_X1 U2915 ( .A(n3873), .ZN(n4840) );
  AND2_X1 U2916 ( .A1(n2886), .A2(REG2_REG_8__SCAN_IN), .ZN(n2315) );
  INV_X2 U2917 ( .A(n3836), .ZN(U4043) );
  INV_X1 U2918 ( .A(IR_REG_24__SCAN_IN), .ZN(n2695) );
  AND2_X1 U2919 ( .A1(n2385), .A2(n2329), .ZN(n2316) );
  AND2_X1 U2920 ( .A1(n4529), .A2(n4521), .ZN(n2317) );
  AND2_X1 U2921 ( .A1(n2806), .A2(n4645), .ZN(n2318) );
  INV_X1 U2922 ( .A(n4643), .ZN(n2807) );
  INV_X1 U2923 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2518) );
  INV_X1 U2924 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2448) );
  AND2_X1 U2925 ( .A1(n2439), .A2(n2438), .ZN(n2320) );
  AND2_X1 U2926 ( .A1(n3092), .A2(n3056), .ZN(n2321) );
  AND2_X1 U2927 ( .A1(n2394), .A2(n2393), .ZN(n2322) );
  OR2_X1 U2928 ( .A1(n3181), .A2(n2807), .ZN(n2323) );
  AND2_X1 U2929 ( .A1(n2161), .A2(REG1_REG_2__SCAN_IN), .ZN(n2324) );
  OR2_X1 U2930 ( .A1(n3415), .A2(n4632), .ZN(n2325) );
  OR2_X1 U2931 ( .A1(n3415), .A2(n4561), .ZN(n2326) );
  INV_X1 U2932 ( .A(n4325), .ZN(n4522) );
  AND2_X1 U2933 ( .A1(n2626), .A2(n3177), .ZN(n2327) );
  INV_X1 U2934 ( .A(n4431), .ZN(n3229) );
  INV_X1 U2935 ( .A(n4344), .ZN(n2556) );
  INV_X1 U2936 ( .A(n3106), .ZN(n3107) );
  INV_X1 U2937 ( .A(n4719), .ZN(n3852) );
  INV_X1 U2938 ( .A(n3706), .ZN(n2676) );
  NAND2_X1 U2939 ( .A1(n2677), .A2(n2676), .ZN(n4206) );
  INV_X1 U2940 ( .A(IR_REG_30__SCAN_IN), .ZN(n2342) );
  OAI22_X1 U2941 ( .A1(n3365), .A2(n2162), .B1(n3021), .B2(n3519), .ZN(n2983)
         );
  AND2_X1 U2942 ( .A1(n2986), .A2(n2985), .ZN(n2987) );
  NAND2_X1 U2943 ( .A1(n4732), .A2(n3856), .ZN(n3857) );
  NAND2_X1 U2944 ( .A1(n4431), .A2(n4564), .ZN(n2494) );
  INV_X1 U2945 ( .A(n3297), .ZN(n3298) );
  OR2_X1 U2946 ( .A1(n3515), .A2(n3514), .ZN(n3516) );
  NOR2_X1 U2947 ( .A1(n3460), .A2(n3462), .ZN(n3458) );
  AND2_X1 U2948 ( .A1(n2864), .A2(n2782), .ZN(n2973) );
  NOR2_X1 U2949 ( .A1(n4681), .A2(n3189), .ZN(n3190) );
  NAND2_X1 U2950 ( .A1(n4730), .A2(n4731), .ZN(n4729) );
  NAND2_X1 U2951 ( .A1(n4325), .A2(n2556), .ZN(n2557) );
  INV_X1 U2952 ( .A(n3833), .ZN(n3082) );
  NAND2_X1 U2953 ( .A1(n2679), .A2(n3890), .ZN(n3895) );
  AOI21_X1 U2954 ( .B1(n4363), .B2(n2546), .A(n2317), .ZN(n4354) );
  INV_X1 U2955 ( .A(n3091), .ZN(n3097) );
  INV_X1 U2956 ( .A(n4547), .ZN(n4792) );
  OR2_X1 U2957 ( .A1(n3428), .A2(n2973), .ZN(n2734) );
  OR2_X1 U2958 ( .A1(n2525), .A2(IR_REG_14__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U2959 ( .A1(n3666), .A2(DATAI_27_), .ZN(n4456) );
  OR2_X1 U2960 ( .A1(n2467), .A2(n4040), .ZN(n2477) );
  INV_X1 U2961 ( .A(n3831), .ZN(n3300) );
  INV_X1 U2962 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3560) );
  NAND2_X1 U2963 ( .A1(n3045), .A2(n3046), .ZN(n3047) );
  NOR2_X1 U2964 ( .A1(n2477), .A2(n3616), .ZN(n2497) );
  OR2_X1 U2965 ( .A1(n2519), .A2(n2518), .ZN(n2527) );
  AND3_X1 U2966 ( .A1(n2890), .A2(n2889), .A3(n2888), .ZN(n3692) );
  AND4_X1 U2967 ( .A1(n2607), .A2(n2606), .A3(n2605), .A4(n2604), .ZN(n4481)
         );
  AND4_X1 U2968 ( .A1(n2563), .A2(n2562), .A3(n2561), .A4(n2560), .ZN(n4304)
         );
  INV_X1 U2969 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3616) );
  AOI21_X1 U2970 ( .B1(n4767), .B2(ADDR_REG_18__SCAN_IN), .A(n4766), .ZN(n4768) );
  NAND2_X1 U2971 ( .A1(n3666), .A2(DATAI_28_), .ZN(n3527) );
  AND2_X1 U2972 ( .A1(n3709), .A2(n4319), .ZN(n4364) );
  INV_X1 U2973 ( .A(n4657), .ZN(n4381) );
  INV_X1 U2974 ( .A(n3361), .ZN(n4416) );
  OR2_X1 U2975 ( .A1(n4886), .A2(n2726), .ZN(n2727) );
  INV_X1 U2976 ( .A(n4480), .ZN(n4231) );
  INV_X1 U2977 ( .A(n4789), .ZN(n4551) );
  INV_X1 U2978 ( .A(n4549), .ZN(n4796) );
  AND2_X1 U2979 ( .A1(n3743), .A2(n3744), .ZN(n3701) );
  AND2_X1 U2980 ( .A1(n2740), .A2(n2625), .ZN(n3530) );
  NOR2_X1 U2981 ( .A1(n2527), .A2(n4651), .ZN(n2548) );
  OR2_X1 U2982 ( .A1(n2449), .A2(n2448), .ZN(n2467) );
  AND2_X1 U2983 ( .A1(n2497), .A2(n2496), .ZN(n2508) );
  INV_X1 U2984 ( .A(n3664), .ZN(n4663) );
  INV_X1 U2985 ( .A(n3692), .ZN(n3886) );
  AND4_X1 U2986 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .ZN(n4476)
         );
  AND4_X1 U2987 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n4325)
         );
  INV_X1 U2988 ( .A(n4771), .ZN(n4756) );
  NAND2_X1 U2989 ( .A1(n4704), .A2(n4705), .ZN(n4703) );
  NAND2_X1 U2990 ( .A1(n4726), .A2(REG1_REG_14__SCAN_IN), .ZN(n4725) );
  INV_X1 U2991 ( .A(n4253), .ZN(n4295) );
  OR2_X1 U2992 ( .A1(n3105), .A2(n3107), .ZN(n4874) );
  AND2_X1 U2993 ( .A1(n4815), .A2(n2739), .ZN(n4802) );
  AND2_X1 U2994 ( .A1(n4815), .A2(n3028), .ZN(n4811) );
  NOR2_X1 U2995 ( .A1(n4895), .A2(n4878), .ZN(n4888) );
  NAND2_X1 U2996 ( .A1(n3666), .A2(DATAI_23_), .ZN(n4268) );
  INV_X1 U2997 ( .A(n4859), .ZN(n4883) );
  NAND2_X1 U2998 ( .A1(n2710), .A2(n2709), .ZN(n2974) );
  OR2_X1 U2999 ( .A1(n2473), .A2(IR_REG_10__SCAN_IN), .ZN(n2506) );
  AND2_X1 U3000 ( .A1(n2786), .A2(n2784), .ZN(n4767) );
  NAND2_X1 U3001 ( .A1(n2977), .A2(STATE_REG_SCAN_IN), .ZN(n4668) );
  OR2_X1 U3002 ( .A1(n2875), .A2(n2868), .ZN(n3664) );
  OAI211_X1 U3003 ( .C1(n3651), .C2(n2635), .A(n2613), .B(n2612), .ZN(n4473)
         );
  INV_X1 U3004 ( .A(n4476), .ZN(n4490) );
  INV_X1 U3005 ( .A(n4568), .ZN(n3829) );
  NAND2_X1 U3006 ( .A1(n2751), .A2(n4407), .ZN(n2752) );
  NAND2_X1 U3007 ( .A1(n4815), .A2(n2750), .ZN(n4388) );
  INV_X1 U3009 ( .A(n4888), .ZN(n4561) );
  OR2_X1 U3010 ( .A1(n4408), .A2(n4438), .ZN(n4633) );
  OR2_X1 U3011 ( .A1(n2729), .A2(n2863), .ZN(n4885) );
  INV_X1 U3012 ( .A(D_REG_16__SCAN_IN), .ZN(n4827) );
  INV_X1 U3013 ( .A(n4835), .ZN(n4834) );
  INV_X1 U3014 ( .A(n4709), .ZN(n4847) );
  INV_X1 U3015 ( .A(n2384), .ZN(n2330) );
  NOR2_X1 U3016 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2335)
         );
  NOR2_X1 U3017 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2334)
         );
  NOR2_X1 U3018 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2333)
         );
  NOR3_X1 U3019 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .A3(
        IR_REG_20__SCAN_IN), .ZN(n2338) );
  XNOR2_X2 U3020 ( .A(n2343), .B(n2342), .ZN(n2349) );
  INV_X1 U3021 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2346) );
  NOR2_X1 U3022 ( .A1(n2348), .A2(n2347), .ZN(n2353) );
  NAND2_X1 U3023 ( .A1(n2378), .A2(REG2_REG_1__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U3024 ( .A1(n2392), .A2(REG3_REG_1__SCAN_IN), .ZN(n2351) );
  NAND3_X1 U3025 ( .A1(n2353), .A2(n2352), .A3(n2351), .ZN(n2364) );
  NAND2_X1 U3026 ( .A1(n2684), .A2(n2355), .ZN(n2357) );
  MUX2_X1 U3027 ( .A(n4648), .B(DATAI_1_), .S(n2383), .Z(n3536) );
  NAND2_X1 U3028 ( .A1(n2364), .A2(n3021), .ZN(n3745) );
  NAND2_X1 U3029 ( .A1(n2392), .A2(REG3_REG_0__SCAN_IN), .ZN(n2363) );
  INV_X1 U3030 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2358) );
  NAND2_X1 U3031 ( .A1(n2359), .A2(REG1_REG_0__SCAN_IN), .ZN(n2360) );
  NAND4_X2 U3032 ( .A1(n2363), .A2(n2362), .A3(n2361), .A4(n2360), .ZN(n2858)
         );
  MUX2_X1 U3033 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2383), .Z(n3029) );
  NAND2_X1 U3034 ( .A1(n2648), .A2(n3020), .ZN(n2366) );
  NAND2_X1 U3035 ( .A1(n2872), .A2(n3536), .ZN(n2365) );
  NAND2_X1 U3036 ( .A1(n2366), .A2(n2365), .ZN(n2941) );
  INV_X1 U3037 ( .A(n2941), .ZN(n2373) );
  NAND2_X1 U3038 ( .A1(n2378), .A2(REG2_REG_2__SCAN_IN), .ZN(n2371) );
  INV_X1 U3039 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2367) );
  OR2_X1 U3040 ( .A1(n2376), .A2(n2367), .ZN(n2370) );
  NAND2_X1 U3041 ( .A1(n2359), .A2(REG1_REG_2__SCAN_IN), .ZN(n2369) );
  NAND2_X1 U3042 ( .A1(n2392), .A2(REG3_REG_2__SCAN_IN), .ZN(n2368) );
  MUX2_X1 U3043 ( .A(n2161), .B(DATAI_2_), .S(n2383), .Z(n3629) );
  NAND2_X1 U3044 ( .A1(n2374), .A2(n3629), .ZN(n3748) );
  INV_X1 U3045 ( .A(n3629), .ZN(n2988) );
  NAND2_X1 U3046 ( .A1(n3537), .A2(n2988), .ZN(n3751) );
  NAND2_X1 U3047 ( .A1(n2374), .A2(n2988), .ZN(n2375) );
  INV_X1 U3048 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2377) );
  OR2_X1 U3049 ( .A1(n2887), .A2(n2377), .ZN(n2382) );
  BUF_X4 U3050 ( .A(n2392), .Z(n2626) );
  NAND2_X1 U3051 ( .A1(n2626), .A2(n4798), .ZN(n2381) );
  BUF_X4 U3052 ( .A(n2378), .Z(n2886) );
  NAND2_X1 U3053 ( .A1(n2384), .A2(IR_REG_31__SCAN_IN), .ZN(n2386) );
  NAND2_X1 U3054 ( .A1(n2386), .A2(n2385), .ZN(n2398) );
  OR2_X1 U3055 ( .A1(n2386), .A2(n2385), .ZN(n2387) );
  NAND2_X1 U3056 ( .A1(n3835), .A2(n4801), .ZN(n2390) );
  NAND2_X1 U3057 ( .A1(n2359), .A2(REG1_REG_4__SCAN_IN), .ZN(n2394) );
  INV_X1 U3058 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2391) );
  XNOR2_X1 U3059 ( .A(n2391), .B(REG3_REG_3__SCAN_IN), .ZN(n3004) );
  NAND2_X1 U3060 ( .A1(n2392), .A2(n3004), .ZN(n2393) );
  INV_X1 U3061 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3062 ( .A1(n2886), .A2(REG2_REG_4__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U3063 ( .A1(n2398), .A2(IR_REG_31__SCAN_IN), .ZN(n2399) );
  XNOR2_X1 U3064 ( .A(n2399), .B(IR_REG_4__SCAN_IN), .ZN(n4645) );
  MUX2_X1 U3065 ( .A(n4645), .B(DATAI_4_), .S(n3666), .Z(n3017) );
  NAND2_X1 U3066 ( .A1(n2886), .A2(REG2_REG_5__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3067 ( .A1(n2158), .A2(REG1_REG_5__SCAN_IN), .ZN(n2404) );
  AOI21_X1 U3068 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2400) );
  NOR2_X1 U3069 ( .A1(n2400), .A2(n2418), .ZN(n2966) );
  NAND2_X1 U3070 ( .A1(n2626), .A2(n2966), .ZN(n2403) );
  INV_X1 U3071 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2401) );
  OR2_X1 U3072 ( .A1(n2887), .A2(n2401), .ZN(n2402) );
  NAND2_X1 U3073 ( .A1(n2406), .A2(IR_REG_31__SCAN_IN), .ZN(n2408) );
  INV_X1 U3074 ( .A(IR_REG_5__SCAN_IN), .ZN(n2407) );
  XNOR2_X1 U3075 ( .A(n2408), .B(n2407), .ZN(n2823) );
  INV_X1 U3076 ( .A(DATAI_5_), .ZN(n2409) );
  MUX2_X1 U3077 ( .A(n2823), .B(n2409), .S(n3666), .Z(n3049) );
  NAND2_X1 U3078 ( .A1(n3083), .A2(n3049), .ZN(n2410) );
  INV_X1 U3079 ( .A(n2410), .ZN(n2413) );
  NAND2_X1 U3080 ( .A1(n4793), .A2(n3017), .ZN(n2963) );
  INV_X1 U3081 ( .A(n2963), .ZN(n2411) );
  NOR2_X1 U3082 ( .A1(n2411), .A2(n2321), .ZN(n2412) );
  OR2_X1 U3083 ( .A1(n2413), .A2(n2412), .ZN(n2414) );
  NAND2_X1 U3084 ( .A1(n2415), .A2(n2414), .ZN(n3089) );
  INV_X1 U3085 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2416) );
  OR2_X1 U3086 ( .A1(n2887), .A2(n2416), .ZN(n2423) );
  INV_X1 U3087 ( .A(n2418), .ZN(n2417) );
  INV_X1 U3088 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2813) );
  NAND2_X1 U3089 ( .A1(n2417), .A2(n2813), .ZN(n2419) );
  NAND2_X1 U3090 ( .A1(n2418), .A2(REG3_REG_6__SCAN_IN), .ZN(n2441) );
  AND2_X1 U3091 ( .A1(n2419), .A2(n2441), .ZN(n4776) );
  NAND2_X1 U3092 ( .A1(n2626), .A2(n4776), .ZN(n2422) );
  NAND2_X1 U3093 ( .A1(n2159), .A2(REG1_REG_6__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U3094 ( .A1(n2886), .A2(REG2_REG_6__SCAN_IN), .ZN(n2420) );
  NAND4_X1 U3095 ( .A1(n2423), .A2(n2422), .A3(n2421), .A4(n2420), .ZN(n3834)
         );
  OR2_X1 U3096 ( .A1(n2424), .A2(n2686), .ZN(n2425) );
  XNOR2_X1 U3097 ( .A(n2425), .B(IR_REG_6__SCAN_IN), .ZN(n4643) );
  MUX2_X1 U3098 ( .A(n4643), .B(DATAI_6_), .S(n3666), .Z(n3091) );
  AND2_X1 U3099 ( .A1(n3834), .A2(n3091), .ZN(n2427) );
  INV_X1 U3100 ( .A(n3834), .ZN(n3142) );
  NAND2_X1 U3101 ( .A1(n3142), .A2(n3097), .ZN(n2426) );
  INV_X1 U3102 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2440) );
  NOR2_X1 U3103 ( .A1(n2441), .A2(n2440), .ZN(n2443) );
  NAND2_X1 U3104 ( .A1(n2443), .A2(REG3_REG_8__SCAN_IN), .ZN(n2449) );
  OR2_X1 U3105 ( .A1(n2443), .A2(REG3_REG_8__SCAN_IN), .ZN(n2428) );
  AND2_X1 U3106 ( .A1(n2449), .A2(n2428), .ZN(n3177) );
  NOR3_X1 U3107 ( .A1(n2315), .A2(n2327), .A3(n2314), .ZN(n2431) );
  INV_X1 U3108 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2429) );
  OR2_X1 U3109 ( .A1(n2887), .A2(n2429), .ZN(n2430) );
  OR2_X1 U3110 ( .A1(n2432), .A2(n2686), .ZN(n2445) );
  INV_X1 U3111 ( .A(IR_REG_7__SCAN_IN), .ZN(n2433) );
  NAND2_X1 U3112 ( .A1(n2445), .A2(n2433), .ZN(n2434) );
  NAND2_X1 U3113 ( .A1(n2434), .A2(IR_REG_31__SCAN_IN), .ZN(n2435) );
  XNOR2_X1 U3114 ( .A(n2435), .B(IR_REG_8__SCAN_IN), .ZN(n3204) );
  INV_X1 U3115 ( .A(DATAI_8_), .ZN(n4854) );
  MUX2_X1 U3116 ( .A(n4855), .B(n4854), .S(n3666), .Z(n3170) );
  INV_X1 U3117 ( .A(n3170), .ZN(n2436) );
  INV_X1 U3118 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2437) );
  OR2_X1 U3119 ( .A1(n2887), .A2(n2437), .ZN(n2439) );
  NAND2_X1 U3120 ( .A1(n2886), .A2(REG2_REG_7__SCAN_IN), .ZN(n2438) );
  AND2_X1 U3121 ( .A1(n2441), .A2(n2440), .ZN(n2442) );
  NOR2_X1 U3122 ( .A1(n2443), .A2(n2442), .ZN(n3156) );
  NAND2_X1 U3123 ( .A1(n2626), .A2(n3156), .ZN(n2444) );
  XNOR2_X1 U3124 ( .A(n2445), .B(IR_REG_7__SCAN_IN), .ZN(n4642) );
  MUX2_X1 U3125 ( .A(n4642), .B(DATAI_7_), .S(n3666), .Z(n3149) );
  NAND2_X1 U3126 ( .A1(n3082), .A2(n3149), .ZN(n2655) );
  INV_X1 U3127 ( .A(n3149), .ZN(n3150) );
  NAND2_X1 U3128 ( .A1(n2159), .A2(REG1_REG_9__SCAN_IN), .ZN(n2455) );
  INV_X1 U3129 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2447) );
  OR2_X1 U3130 ( .A1(n2887), .A2(n2447), .ZN(n2454) );
  NAND2_X1 U3131 ( .A1(n2886), .A2(REG2_REG_9__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U3132 ( .A1(n2449), .A2(n2448), .ZN(n2450) );
  NAND2_X1 U3133 ( .A1(n2467), .A2(n2450), .ZN(n3272) );
  INV_X1 U3134 ( .A(n3272), .ZN(n2451) );
  NAND2_X1 U3135 ( .A1(n2626), .A2(n2451), .ZN(n2452) );
  NAND2_X1 U3136 ( .A1(n2456), .A2(IR_REG_31__SCAN_IN), .ZN(n2457) );
  XNOR2_X1 U3137 ( .A(n2457), .B(IR_REG_9__SCAN_IN), .ZN(n3206) );
  MUX2_X1 U3138 ( .A(n3206), .B(DATAI_9_), .S(n3666), .Z(n3269) );
  INV_X1 U3139 ( .A(n3269), .ZN(n3262) );
  AND2_X1 U3140 ( .A1(n3300), .A2(n3262), .ZN(n2463) );
  NAND2_X1 U3141 ( .A1(n3832), .A2(n2436), .ZN(n2459) );
  NAND2_X1 U3142 ( .A1(n3833), .A2(n3149), .ZN(n3108) );
  AND2_X1 U3143 ( .A1(n2459), .A2(n3108), .ZN(n2460) );
  AND2_X1 U3144 ( .A1(n2183), .A2(n3131), .ZN(n2462) );
  NOR2_X1 U3145 ( .A1(n2463), .A2(n2462), .ZN(n2464) );
  INV_X1 U3146 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2466) );
  OR2_X1 U3147 ( .A1(n2887), .A2(n2466), .ZN(n2472) );
  NAND2_X1 U31480 ( .A1(n2159), .A2(REG1_REG_10__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U31490 ( .A1(n2467), .A2(n4040), .ZN(n2468) );
  NAND2_X1 U3150 ( .A1(n2626), .A2(n3249), .ZN(n2470) );
  NAND2_X1 U3151 ( .A1(n2886), .A2(REG2_REG_10__SCAN_IN), .ZN(n2469) );
  NAND4_X1 U3152 ( .A1(n2472), .A2(n2471), .A3(n2470), .A4(n2469), .ZN(n3830)
         );
  NAND2_X1 U3153 ( .A1(n2473), .A2(IR_REG_31__SCAN_IN), .ZN(n2474) );
  MUX2_X1 U3154 ( .A(IR_REG_31__SCAN_IN), .B(n2474), .S(IR_REG_10__SCAN_IN), 
        .Z(n2475) );
  NAND2_X1 U3155 ( .A1(n2475), .A2(n2506), .ZN(n4851) );
  INV_X1 U3156 ( .A(n4851), .ZN(n3208) );
  MUX2_X1 U3157 ( .A(n3208), .B(DATAI_10_), .S(n3666), .Z(n3302) );
  NOR2_X1 U3158 ( .A1(n3830), .A2(n3302), .ZN(n2476) );
  INV_X1 U3159 ( .A(n3830), .ZN(n3617) );
  NAND2_X1 U3160 ( .A1(n2158), .A2(REG1_REG_11__SCAN_IN), .ZN(n2483) );
  AND2_X1 U3161 ( .A1(n2477), .A2(n3616), .ZN(n2478) );
  NOR2_X1 U3162 ( .A1(n2497), .A2(n2478), .ZN(n3620) );
  NAND2_X1 U3163 ( .A1(n2626), .A2(n3620), .ZN(n2482) );
  NAND2_X1 U3164 ( .A1(n2886), .A2(REG2_REG_11__SCAN_IN), .ZN(n2481) );
  INV_X1 U3165 ( .A(REG0_REG_11__SCAN_IN), .ZN(n2479) );
  OR2_X1 U3166 ( .A1(n2887), .A2(n2479), .ZN(n2480) );
  NAND2_X1 U3167 ( .A1(n2506), .A2(IR_REG_31__SCAN_IN), .ZN(n2490) );
  XNOR2_X1 U3168 ( .A(n2490), .B(IR_REG_11__SCAN_IN), .ZN(n3211) );
  MUX2_X1 U3169 ( .A(n3211), .B(DATAI_11_), .S(n3666), .Z(n3619) );
  NAND2_X1 U3170 ( .A1(n4568), .A2(n3619), .ZN(n3742) );
  INV_X1 U3171 ( .A(n3619), .ZN(n3335) );
  NAND2_X1 U3172 ( .A1(n3829), .A2(n3335), .ZN(n3779) );
  NAND2_X1 U3173 ( .A1(n4568), .A2(n3335), .ZN(n2484) );
  NAND2_X1 U3174 ( .A1(n2158), .A2(REG1_REG_12__SCAN_IN), .ZN(n2489) );
  INV_X1 U3175 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2485) );
  XNOR2_X1 U3176 ( .A(n2497), .B(n2485), .ZN(n3552) );
  NAND2_X1 U3177 ( .A1(n2626), .A2(n3552), .ZN(n2488) );
  NAND2_X1 U3178 ( .A1(n2886), .A2(REG2_REG_12__SCAN_IN), .ZN(n2487) );
  INV_X1 U3179 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4074) );
  OR2_X1 U3180 ( .A1(n2887), .A2(n4074), .ZN(n2486) );
  NAND2_X1 U3181 ( .A1(n2490), .A2(n2504), .ZN(n2491) );
  NAND2_X1 U3182 ( .A1(n2491), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  XNOR2_X1 U3183 ( .A(n2492), .B(n2503), .ZN(n3216) );
  MUX2_X1 U3184 ( .A(n3216), .B(n4086), .S(n3666), .Z(n4564) );
  OR2_X1 U3185 ( .A1(n4431), .A2(n4564), .ZN(n2493) );
  INV_X1 U3186 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4630) );
  OR2_X1 U3187 ( .A1(n2887), .A2(n4630), .ZN(n2502) );
  NAND2_X1 U3188 ( .A1(n2158), .A2(REG1_REG_13__SCAN_IN), .ZN(n2501) );
  AND2_X1 U3189 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_13__SCAN_IN), .ZN(
        n2496) );
  AOI21_X1 U3190 ( .B1(n2497), .B2(REG3_REG_12__SCAN_IN), .A(
        REG3_REG_13__SCAN_IN), .ZN(n2498) );
  OR2_X1 U3191 ( .A1(n2508), .A2(n2498), .ZN(n3604) );
  INV_X1 U3192 ( .A(n3604), .ZN(n4439) );
  NAND2_X1 U3193 ( .A1(n2626), .A2(n4439), .ZN(n2500) );
  NAND2_X1 U3194 ( .A1(n2886), .A2(REG2_REG_13__SCAN_IN), .ZN(n2499) );
  NAND4_X1 U3195 ( .A1(n2502), .A2(n2501), .A3(n2500), .A4(n2499), .ZN(n4566)
         );
  NAND2_X1 U3196 ( .A1(n2504), .A2(n2503), .ZN(n2505) );
  NOR2_X1 U3197 ( .A1(n2506), .A2(n2505), .ZN(n2515) );
  OR2_X1 U3198 ( .A1(n2515), .A2(n2686), .ZN(n2507) );
  XNOR2_X1 U3199 ( .A(n2507), .B(IR_REG_13__SCAN_IN), .ZN(n4709) );
  MUX2_X1 U3200 ( .A(n4709), .B(DATAI_13_), .S(n3666), .Z(n4428) );
  NOR2_X1 U3201 ( .A1(n4566), .A2(n4428), .ZN(n3714) );
  NAND2_X1 U3202 ( .A1(n4566), .A2(n4428), .ZN(n3712) );
  NAND2_X1 U3203 ( .A1(n2159), .A2(REG1_REG_14__SCAN_IN), .ZN(n2513) );
  OR2_X1 U3204 ( .A1(n2508), .A2(REG3_REG_14__SCAN_IN), .ZN(n2509) );
  NAND2_X1 U3205 ( .A1(n2508), .A2(REG3_REG_14__SCAN_IN), .ZN(n2519) );
  AND2_X1 U3206 ( .A1(n2509), .A2(n2519), .ZN(n4413) );
  NAND2_X1 U3207 ( .A1(n2626), .A2(n4413), .ZN(n2512) );
  NAND2_X1 U3208 ( .A1(n2886), .A2(REG2_REG_14__SCAN_IN), .ZN(n2511) );
  INV_X1 U3209 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4626) );
  OR2_X1 U32100 ( .A1(n2887), .A2(n4626), .ZN(n2510) );
  INV_X1 U32110 ( .A(IR_REG_13__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U32120 ( .A1(n2515), .A2(n2514), .ZN(n2525) );
  NAND2_X1 U32130 ( .A1(n2525), .A2(IR_REG_31__SCAN_IN), .ZN(n2516) );
  XNOR2_X1 U32140 ( .A(n2516), .B(IR_REG_14__SCAN_IN), .ZN(n4719) );
  MUX2_X1 U32150 ( .A(n4719), .B(DATAI_14_), .S(n3666), .Z(n2517) );
  NAND2_X1 U32160 ( .A1(n4542), .A2(n2517), .ZN(n3668) );
  NAND2_X1 U32170 ( .A1(n4429), .A2(n4546), .ZN(n3669) );
  INV_X1 U32180 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4622) );
  OR2_X1 U32190 ( .A1(n2887), .A2(n4622), .ZN(n2524) );
  NAND2_X1 U32200 ( .A1(n2158), .A2(REG1_REG_15__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32210 ( .A1(n2519), .A2(n2518), .ZN(n2520) );
  AND2_X1 U32220 ( .A1(n2527), .A2(n2520), .ZN(n4396) );
  NAND2_X1 U32230 ( .A1(n2626), .A2(n4396), .ZN(n2522) );
  NAND2_X1 U32240 ( .A1(n2886), .A2(REG2_REG_15__SCAN_IN), .ZN(n2521) );
  NAND4_X1 U32250 ( .A1(n2524), .A2(n2523), .A3(n2522), .A4(n2521), .ZN(n4410)
         );
  NAND2_X1 U32260 ( .A1(n2526), .A2(IR_REG_31__SCAN_IN), .ZN(n2534) );
  XNOR2_X1 U32270 ( .A(n2534), .B(IR_REG_15__SCAN_IN), .ZN(n3869) );
  MUX2_X1 U32280 ( .A(n3869), .B(DATAI_15_), .S(n3666), .Z(n4538) );
  AND2_X1 U32290 ( .A1(n2527), .A2(n4651), .ZN(n2528) );
  OR2_X1 U32300 ( .A1(n2528), .A2(n2548), .ZN(n4667) );
  INV_X1 U32310 ( .A(n4667), .ZN(n4378) );
  NAND2_X1 U32320 ( .A1(n2626), .A2(n4378), .ZN(n2532) );
  NAND2_X1 U32330 ( .A1(n2159), .A2(REG1_REG_16__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32340 ( .A1(n2886), .A2(REG2_REG_16__SCAN_IN), .ZN(n2530) );
  INV_X1 U32350 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4067) );
  OR2_X1 U32360 ( .A1(n2887), .A2(n4067), .ZN(n2529) );
  NAND2_X1 U32370 ( .A1(n2534), .A2(n2533), .ZN(n2535) );
  NAND2_X1 U32380 ( .A1(n2535), .A2(IR_REG_31__SCAN_IN), .ZN(n2536) );
  XNOR2_X1 U32390 ( .A(n2536), .B(IR_REG_16__SCAN_IN), .ZN(n4740) );
  MUX2_X1 U32400 ( .A(n4740), .B(DATAI_16_), .S(n3666), .Z(n4657) );
  NAND2_X1 U32410 ( .A1(n4525), .A2(n4657), .ZN(n3788) );
  NAND2_X1 U32420 ( .A1(n4539), .A2(n4381), .ZN(n3672) );
  NAND2_X1 U32430 ( .A1(n3788), .A2(n3672), .ZN(n4375) );
  INV_X1 U32440 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2537) );
  XNOR2_X1 U32450 ( .A(n2548), .B(n2537), .ZN(n4366) );
  NAND2_X1 U32460 ( .A1(n2626), .A2(n4366), .ZN(n2541) );
  NAND2_X1 U32470 ( .A1(n2158), .A2(REG1_REG_17__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32480 ( .A1(n2886), .A2(REG2_REG_17__SCAN_IN), .ZN(n2539) );
  INV_X1 U32490 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4617) );
  OR2_X1 U32500 ( .A1(n2887), .A2(n4617), .ZN(n2538) );
  NAND2_X1 U32510 ( .A1(n2543), .A2(IR_REG_31__SCAN_IN), .ZN(n2544) );
  XNOR2_X1 U32520 ( .A(n2544), .B(IR_REG_17__SCAN_IN), .ZN(n3873) );
  INV_X1 U32530 ( .A(DATAI_17_), .ZN(n2545) );
  MUX2_X1 U32540 ( .A(n4840), .B(n2545), .S(n3666), .Z(n4369) );
  NAND2_X1 U32550 ( .A1(n4654), .A2(n4369), .ZN(n2546) );
  INV_X1 U32560 ( .A(n4369), .ZN(n4521) );
  NAND2_X1 U32570 ( .A1(n2159), .A2(REG1_REG_18__SCAN_IN), .ZN(n2553) );
  AND2_X1 U32580 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2547) );
  AOI21_X1 U32590 ( .B1(n2548), .B2(REG3_REG_17__SCAN_IN), .A(
        REG3_REG_18__SCAN_IN), .ZN(n2549) );
  OR2_X1 U32600 ( .A1(n2558), .A2(n2549), .ZN(n4351) );
  INV_X1 U32610 ( .A(n4351), .ZN(n3643) );
  NAND2_X1 U32620 ( .A1(n2626), .A2(n3643), .ZN(n2552) );
  NAND2_X1 U32630 ( .A1(n2886), .A2(REG2_REG_18__SCAN_IN), .ZN(n2551) );
  INV_X1 U32640 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4010) );
  OR2_X1 U32650 ( .A1(n2887), .A2(n4010), .ZN(n2550) );
  OR2_X1 U32660 ( .A1(n2554), .A2(n2686), .ZN(n2555) );
  XNOR2_X1 U32670 ( .A(n2555), .B(IR_REG_18__SCAN_IN), .ZN(n3862) );
  MUX2_X1 U32680 ( .A(n3862), .B(DATAI_18_), .S(n3666), .Z(n4344) );
  NAND2_X1 U32690 ( .A1(n4325), .A2(n4344), .ZN(n4321) );
  NAND2_X1 U32700 ( .A1(n4522), .A2(n2556), .ZN(n4322) );
  NAND2_X1 U32710 ( .A1(n4321), .A2(n4322), .ZN(n4353) );
  NAND2_X1 U32720 ( .A1(n4354), .A2(n4353), .ZN(n4352) );
  NAND2_X1 U32730 ( .A1(n2158), .A2(REG1_REG_19__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32740 ( .A1(n2558), .A2(REG3_REG_19__SCAN_IN), .ZN(n2571) );
  OR2_X1 U32750 ( .A1(n2558), .A2(REG3_REG_19__SCAN_IN), .ZN(n2559) );
  AND2_X1 U32760 ( .A1(n2571), .A2(n2559), .ZN(n3500) );
  NAND2_X1 U32770 ( .A1(n2626), .A2(n3500), .ZN(n2562) );
  NAND2_X1 U32780 ( .A1(n2886), .A2(REG2_REG_19__SCAN_IN), .ZN(n2561) );
  INV_X1 U32790 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4612) );
  OR2_X1 U32800 ( .A1(n2887), .A2(n4612), .ZN(n2560) );
  INV_X1 U32810 ( .A(n4304), .ZN(n4345) );
  MUX2_X1 U32820 ( .A(n4349), .B(DATAI_19_), .S(n3666), .Z(n3719) );
  NAND2_X1 U32830 ( .A1(n4345), .A2(n3719), .ZN(n2565) );
  NAND2_X1 U32840 ( .A1(n2159), .A2(REG1_REG_20__SCAN_IN), .ZN(n2569) );
  XNOR2_X1 U32850 ( .A(n2571), .B(REG3_REG_20__SCAN_IN), .ZN(n4314) );
  NAND2_X1 U32860 ( .A1(n2626), .A2(n4314), .ZN(n2568) );
  NAND2_X1 U32870 ( .A1(n2886), .A2(REG2_REG_20__SCAN_IN), .ZN(n2567) );
  INV_X1 U32880 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4608) );
  OR2_X1 U32890 ( .A1(n2887), .A2(n4608), .ZN(n2566) );
  NOR2_X1 U32900 ( .A1(n4326), .A2(n4312), .ZN(n3717) );
  NAND2_X1 U32910 ( .A1(n4326), .A2(n4312), .ZN(n3715) );
  NAND2_X1 U32920 ( .A1(n2158), .A2(REG1_REG_21__SCAN_IN), .ZN(n2576) );
  INV_X1 U32930 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3591) );
  INV_X1 U32940 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3407) );
  OAI21_X1 U32950 ( .B1(n2571), .B2(n3591), .A(n3407), .ZN(n2572) );
  NAND2_X1 U32960 ( .A1(REG3_REG_20__SCAN_IN), .A2(REG3_REG_21__SCAN_IN), .ZN(
        n2570) );
  AND2_X1 U32970 ( .A1(n2572), .A2(n2578), .ZN(n4292) );
  NAND2_X1 U32980 ( .A1(n2626), .A2(n4292), .ZN(n2575) );
  NAND2_X1 U32990 ( .A1(n2886), .A2(REG2_REG_21__SCAN_IN), .ZN(n2574) );
  INV_X1 U33000 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4604) );
  OR2_X1 U33010 ( .A1(n2887), .A2(n4604), .ZN(n2573) );
  INV_X1 U33020 ( .A(n4305), .ZN(n2901) );
  NAND2_X1 U33030 ( .A1(n2901), .A2(n4290), .ZN(n2577) );
  NAND2_X1 U33040 ( .A1(n2159), .A2(REG1_REG_22__SCAN_IN), .ZN(n2584) );
  NOR2_X1 U33050 ( .A1(n2578), .A2(n4035), .ZN(n2587) );
  AND2_X1 U33060 ( .A1(n2578), .A2(n4035), .ZN(n2579) );
  NOR2_X1 U33070 ( .A1(n2587), .A2(n2579), .ZN(n4282) );
  NAND2_X1 U33080 ( .A1(n2626), .A2(n4282), .ZN(n2583) );
  NAND2_X1 U33090 ( .A1(n2886), .A2(REG2_REG_22__SCAN_IN), .ZN(n2582) );
  INV_X1 U33100 ( .A(REG0_REG_22__SCAN_IN), .ZN(n2580) );
  OR2_X1 U33110 ( .A1(n2887), .A2(n2580), .ZN(n2581) );
  INV_X1 U33120 ( .A(n4283), .ZN(n2585) );
  NAND2_X1 U33130 ( .A1(n4502), .A2(n2585), .ZN(n4256) );
  NAND2_X1 U33140 ( .A1(n4291), .A2(n4283), .ZN(n2671) );
  NAND2_X1 U33150 ( .A1(n4256), .A2(n2671), .ZN(n4274) );
  OR2_X1 U33160 ( .A1(n4502), .A2(n4283), .ZN(n2586) );
  INV_X1 U33170 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4597) );
  OR2_X1 U33180 ( .A1(n2887), .A2(n4597), .ZN(n2592) );
  NAND2_X1 U33190 ( .A1(n2158), .A2(REG1_REG_23__SCAN_IN), .ZN(n2591) );
  NOR2_X1 U33200 ( .A1(n2587), .A2(REG3_REG_23__SCAN_IN), .ZN(n2588) );
  NOR2_X1 U33210 ( .A1(n2595), .A2(n2588), .ZN(n4265) );
  NAND2_X1 U33220 ( .A1(n2626), .A2(n4265), .ZN(n2590) );
  NAND2_X1 U33230 ( .A1(n2886), .A2(REG2_REG_23__SCAN_IN), .ZN(n2589) );
  NAND4_X1 U33240 ( .A1(n2592), .A2(n2591), .A3(n2590), .A4(n2589), .ZN(n4483)
         );
  INV_X1 U33250 ( .A(n4483), .ZN(n3608) );
  NAND2_X1 U33260 ( .A1(n3608), .A2(n4268), .ZN(n2594) );
  NAND2_X1 U33270 ( .A1(n2159), .A2(REG1_REG_24__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U33280 ( .A1(n2595), .A2(REG3_REG_24__SCAN_IN), .ZN(n2602) );
  OR2_X1 U33290 ( .A1(n2595), .A2(REG3_REG_24__SCAN_IN), .ZN(n2596) );
  AND2_X1 U33300 ( .A1(n2602), .A2(n2596), .ZN(n4233) );
  NAND2_X1 U33310 ( .A1(n2626), .A2(n4233), .ZN(n2599) );
  NAND2_X1 U33320 ( .A1(n2886), .A2(REG2_REG_24__SCAN_IN), .ZN(n2598) );
  INV_X1 U33330 ( .A(REG0_REG_24__SCAN_IN), .ZN(n3978) );
  OR2_X1 U33340 ( .A1(n2887), .A2(n3978), .ZN(n2597) );
  NAND2_X1 U33350 ( .A1(n4490), .A2(n4231), .ZN(n2601) );
  NAND2_X1 U33360 ( .A1(n2602), .A2(n3560), .ZN(n2603) );
  AND2_X1 U33370 ( .A1(n2610), .A2(n2603), .ZN(n4220) );
  NAND2_X1 U33380 ( .A1(n4220), .A2(n2626), .ZN(n2607) );
  NAND2_X1 U33390 ( .A1(n2159), .A2(REG1_REG_25__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U33400 ( .A1(n2886), .A2(REG2_REG_25__SCAN_IN), .ZN(n2605) );
  INV_X1 U33410 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4589) );
  OR2_X1 U33420 ( .A1(n2887), .A2(n4589), .ZN(n2604) );
  NAND2_X1 U33430 ( .A1(n4481), .A2(n4223), .ZN(n2609) );
  NOR2_X1 U33440 ( .A1(n4481), .A2(n4223), .ZN(n2608) );
  INV_X1 U33450 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3923) );
  NAND2_X1 U33460 ( .A1(n2610), .A2(n3923), .ZN(n2611) );
  NAND2_X1 U33470 ( .A1(n2624), .A2(n2611), .ZN(n3651) );
  INV_X1 U33480 ( .A(n2626), .ZN(n2635) );
  INV_X1 U33490 ( .A(n2887), .ZN(n2632) );
  AOI22_X1 U33500 ( .A1(n2632), .A2(REG0_REG_26__SCAN_IN), .B1(n2158), .B2(
        REG1_REG_26__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U33510 ( .A1(n2886), .A2(REG2_REG_26__SCAN_IN), .ZN(n2612) );
  INV_X1 U33520 ( .A(n4464), .ZN(n3468) );
  NAND2_X1 U3353 ( .A1(n4473), .A2(n3468), .ZN(n2615) );
  NOR2_X1 U33540 ( .A1(n4473), .A2(n3468), .ZN(n2614) );
  XNOR2_X1 U3355 ( .A(n2624), .B(REG3_REG_27__SCAN_IN), .ZN(n3900) );
  NAND2_X1 U3356 ( .A1(n3900), .A2(n2626), .ZN(n2621) );
  INV_X1 U3357 ( .A(REG0_REG_27__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U3358 ( .A1(n2886), .A2(REG2_REG_27__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U3359 ( .A1(n2159), .A2(REG1_REG_27__SCAN_IN), .ZN(n2616) );
  OAI211_X1 U3360 ( .C1(n2887), .C2(n2618), .A(n2617), .B(n2616), .ZN(n2619)
         );
  INV_X1 U3361 ( .A(n2619), .ZN(n2620) );
  NAND2_X1 U3362 ( .A1(n3803), .A2(n4456), .ZN(n2622) );
  NAND2_X1 U3363 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2623) );
  INV_X1 U3364 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4098) );
  INV_X1 U3365 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3526) );
  OAI21_X1 U3366 ( .B1(n2624), .B2(n4098), .A(n3526), .ZN(n2625) );
  NAND2_X1 U3367 ( .A1(n3530), .A2(n2626), .ZN(n2631) );
  INV_X1 U3368 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3962) );
  NAND2_X1 U3369 ( .A1(n2886), .A2(REG2_REG_28__SCAN_IN), .ZN(n2628) );
  NAND2_X1 U3370 ( .A1(n2158), .A2(REG1_REG_28__SCAN_IN), .ZN(n2627) );
  OAI211_X1 U3371 ( .C1(n2887), .C2(n3962), .A(n2628), .B(n2627), .ZN(n2629)
         );
  INV_X1 U3372 ( .A(n2629), .ZN(n2630) );
  NAND2_X1 U3373 ( .A1(n2631), .A2(n2630), .ZN(n4458) );
  OR2_X1 U3374 ( .A1(n4458), .A2(n3527), .ZN(n3679) );
  NAND2_X1 U3375 ( .A1(n4458), .A2(n3527), .ZN(n3682) );
  INV_X1 U3376 ( .A(n4458), .ZN(n3521) );
  OAI22_X1 U3377 ( .A1(n2755), .A2(n3698), .B1(n3521), .B2(n3527), .ZN(n2636)
         );
  AOI22_X1 U3378 ( .A1(REG1_REG_29__SCAN_IN), .A2(n2158), .B1(n2632), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U3379 ( .A1(n2886), .A2(REG2_REG_29__SCAN_IN), .ZN(n2633) );
  OAI211_X1 U3380 ( .C1(n2740), .C2(n2635), .A(n2634), .B(n2633), .ZN(n3828)
         );
  NAND2_X1 U3381 ( .A1(n3666), .A2(DATAI_29_), .ZN(n3684) );
  INV_X1 U3382 ( .A(n3684), .ZN(n2747) );
  XNOR2_X1 U3383 ( .A(n3828), .B(n2747), .ZN(n2681) );
  XNOR2_X1 U3384 ( .A(n2636), .B(n2681), .ZN(n2751) );
  NAND2_X1 U3385 ( .A1(n2642), .A2(n2637), .ZN(n2638) );
  OAI21_X1 U3386 ( .B1(IR_REG_19__SCAN_IN), .B2(IR_REG_20__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U3387 ( .A1(n2642), .A2(n2641), .ZN(n2644) );
  NAND2_X1 U3388 ( .A1(n2645), .A2(IR_REG_31__SCAN_IN), .ZN(n2646) );
  XNOR2_X1 U3389 ( .A(n2980), .B(n2870), .ZN(n2647) );
  NAND2_X1 U3390 ( .A1(n3813), .A2(n4349), .ZN(n4808) );
  INV_X1 U3391 ( .A(n2870), .ZN(n3820) );
  INV_X1 U3392 ( .A(n3746), .ZN(n3736) );
  INV_X1 U3393 ( .A(n3813), .ZN(n4640) );
  INV_X1 U3394 ( .A(n2858), .ZN(n2855) );
  NAND2_X1 U3395 ( .A1(n2855), .A2(n3029), .ZN(n3743) );
  OR2_X1 U3396 ( .A1(n2648), .A2(n3743), .ZN(n3023) );
  NAND2_X1 U3397 ( .A1(n3023), .A2(n2649), .ZN(n2651) );
  NAND2_X1 U3398 ( .A1(n2651), .A2(n2945), .ZN(n2947) );
  NAND2_X1 U3399 ( .A1(n2947), .A2(n3748), .ZN(n4787) );
  INV_X1 U3400 ( .A(n4801), .ZN(n2993) );
  NAND2_X1 U3401 ( .A1(n3835), .A2(n2993), .ZN(n3750) );
  NAND2_X1 U3402 ( .A1(n4787), .A2(n4788), .ZN(n4786) );
  NAND2_X1 U3403 ( .A1(n4786), .A2(n3753), .ZN(n3062) );
  INV_X1 U3404 ( .A(n2652), .ZN(n2653) );
  AND2_X1 U3405 ( .A1(n3092), .A2(n3049), .ZN(n2958) );
  NAND2_X1 U3406 ( .A1(n3083), .A2(n3056), .ZN(n3768) );
  NAND2_X1 U3407 ( .A1(n3834), .A2(n3097), .ZN(n3770) );
  NAND2_X1 U3408 ( .A1(n3090), .A2(n3770), .ZN(n2654) );
  NAND2_X1 U3409 ( .A1(n3142), .A2(n3091), .ZN(n3759) );
  NAND2_X1 U3410 ( .A1(n2654), .A2(n3759), .ZN(n3151) );
  INV_X1 U3411 ( .A(n2655), .ZN(n3761) );
  OAI21_X2 U3412 ( .B1(n3151), .B2(n3761), .A(n3758), .ZN(n3110) );
  NAND2_X1 U3413 ( .A1(n3267), .A2(n2436), .ZN(n3763) );
  NAND2_X1 U3414 ( .A1(n3110), .A2(n3763), .ZN(n2656) );
  NAND2_X1 U3415 ( .A1(n3832), .A2(n3170), .ZN(n3771) );
  AND2_X1 U3416 ( .A1(n3831), .A2(n3262), .ZN(n3766) );
  NAND2_X1 U3417 ( .A1(n3300), .A2(n3269), .ZN(n3764) );
  NAND2_X1 U3418 ( .A1(n3830), .A2(n3291), .ZN(n3780) );
  NAND2_X1 U3419 ( .A1(n3254), .A2(n3780), .ZN(n2657) );
  NAND2_X1 U3420 ( .A1(n3617), .A2(n3302), .ZN(n3774) );
  NAND2_X1 U3421 ( .A1(n2657), .A2(n3774), .ZN(n3219) );
  NAND2_X1 U3422 ( .A1(n3219), .A2(n3779), .ZN(n2658) );
  NAND2_X1 U3423 ( .A1(n2658), .A2(n3742), .ZN(n4425) );
  NAND2_X1 U3424 ( .A1(n3229), .A2(n4564), .ZN(n4423) );
  NAND2_X1 U3425 ( .A1(n4566), .A2(n4437), .ZN(n2659) );
  AND2_X1 U3426 ( .A1(n4423), .A2(n2659), .ZN(n3738) );
  NAND2_X1 U3427 ( .A1(n4425), .A2(n3738), .ZN(n2661) );
  NOR2_X1 U3428 ( .A1(n3229), .A2(n4564), .ZN(n4424) );
  NOR2_X1 U3429 ( .A1(n4566), .A2(n4437), .ZN(n2660) );
  AOI21_X1 U3430 ( .B1(n3738), .B2(n4424), .A(n2660), .ZN(n3741) );
  NAND2_X1 U3431 ( .A1(n2661), .A2(n3741), .ZN(n4404) );
  NAND2_X1 U3432 ( .A1(n4404), .A2(n4405), .ZN(n2662) );
  NAND2_X1 U3433 ( .A1(n2662), .A2(n3668), .ZN(n4389) );
  NAND2_X1 U3434 ( .A1(n4652), .A2(n4538), .ZN(n3671) );
  NAND2_X1 U3435 ( .A1(n4410), .A2(n4399), .ZN(n3670) );
  NAND2_X1 U3436 ( .A1(n3671), .A2(n3670), .ZN(n4392) );
  OR2_X2 U3437 ( .A1(n4389), .A2(n4392), .ZN(n4390) );
  NAND2_X1 U3438 ( .A1(n4390), .A2(n3670), .ZN(n4384) );
  INV_X1 U3439 ( .A(n4375), .ZN(n4383) );
  NAND2_X1 U3440 ( .A1(n4384), .A2(n4383), .ZN(n4382) );
  NAND2_X2 U3441 ( .A1(n4382), .A2(n3672), .ZN(n4361) );
  NAND2_X1 U3442 ( .A1(n4654), .A2(n4521), .ZN(n4319) );
  NAND2_X1 U3443 ( .A1(n4321), .A2(n4319), .ZN(n2664) );
  NAND2_X1 U3444 ( .A1(n4345), .A2(n4333), .ZN(n2663) );
  AND2_X1 U3445 ( .A1(n4322), .A2(n2663), .ZN(n2668) );
  NAND2_X1 U3446 ( .A1(n2664), .A2(n2668), .ZN(n2666) );
  NAND2_X1 U3447 ( .A1(n4304), .A2(n3719), .ZN(n2665) );
  NAND2_X1 U3448 ( .A1(n2666), .A2(n2665), .ZN(n4246) );
  NOR2_X1 U3449 ( .A1(n4504), .A2(n4312), .ZN(n4250) );
  NAND2_X1 U3450 ( .A1(n4504), .A2(n4312), .ZN(n4249) );
  OAI21_X1 U3451 ( .B1(n4246), .B2(n4250), .A(n4249), .ZN(n3791) );
  NAND2_X1 U3452 ( .A1(n4305), .A2(n4290), .ZN(n4254) );
  AND2_X1 U3453 ( .A1(n4256), .A2(n4254), .ZN(n3797) );
  AND2_X1 U3454 ( .A1(n3791), .A2(n3797), .ZN(n2667) );
  NAND2_X1 U3455 ( .A1(n4361), .A2(n2667), .ZN(n2674) );
  INV_X1 U3456 ( .A(n2667), .ZN(n3675) );
  INV_X1 U3457 ( .A(n2668), .ZN(n2669) );
  AND2_X1 U34580 ( .A1(n4529), .A2(n4369), .ZN(n4320) );
  NOR2_X1 U34590 ( .A1(n2669), .A2(n4320), .ZN(n4244) );
  AND2_X1 U3460 ( .A1(n4244), .A2(n4249), .ZN(n3793) );
  OR2_X1 U3461 ( .A1(n3675), .A2(n3793), .ZN(n2673) );
  NOR2_X1 U3462 ( .A1(n4305), .A2(n4290), .ZN(n3798) );
  NAND2_X1 U3463 ( .A1(n4483), .A2(n4268), .ZN(n2670) );
  NAND2_X1 U3464 ( .A1(n2671), .A2(n2670), .ZN(n3795) );
  AOI21_X1 U3465 ( .B1(n3798), .B2(n4256), .A(n3795), .ZN(n2672) );
  AND2_X1 U3466 ( .A1(n2673), .A2(n2672), .ZN(n3674) );
  NAND2_X1 U34670 ( .A1(n2674), .A2(n3674), .ZN(n4237) );
  NAND2_X1 U3468 ( .A1(n3608), .A2(n4489), .ZN(n4236) );
  NAND2_X1 U34690 ( .A1(n4476), .A2(n4231), .ZN(n3708) );
  AND2_X1 U3470 ( .A1(n4236), .A2(n3708), .ZN(n3799) );
  NAND2_X1 U34710 ( .A1(n4237), .A2(n3799), .ZN(n2675) );
  NAND2_X1 U3472 ( .A1(n4490), .A2(n4480), .ZN(n3707) );
  NAND2_X1 U34730 ( .A1(n2675), .A2(n3707), .ZN(n4214) );
  INV_X1 U3474 ( .A(n4214), .ZN(n2677) );
  INV_X1 U34750 ( .A(n4481), .ZN(n4232) );
  AND2_X1 U3476 ( .A1(n4232), .A2(n4223), .ZN(n3706) );
  OR2_X1 U34770 ( .A1(n4473), .A2(n4464), .ZN(n3699) );
  INV_X1 U3478 ( .A(n4223), .ZN(n4472) );
  NAND2_X1 U34790 ( .A1(n4481), .A2(n4472), .ZN(n4205) );
  AND2_X1 U3480 ( .A1(n3699), .A2(n4205), .ZN(n3807) );
  NAND2_X1 U34810 ( .A1(n4206), .A2(n3807), .ZN(n2678) );
  NAND2_X1 U3482 ( .A1(n4473), .A2(n4464), .ZN(n3700) );
  NAND2_X1 U34830 ( .A1(n2678), .A2(n3700), .ZN(n3893) );
  INV_X1 U3484 ( .A(n3893), .ZN(n2679) );
  XNOR2_X1 U34850 ( .A(n4466), .B(n3897), .ZN(n3890) );
  INV_X1 U3486 ( .A(n3890), .ZN(n3892) );
  NAND2_X1 U34870 ( .A1(n3803), .A2(n3897), .ZN(n3678) );
  NAND2_X1 U3488 ( .A1(n3895), .A2(n3678), .ZN(n2756) );
  INV_X1 U34890 ( .A(n3679), .ZN(n2680) );
  AOI21_X1 U3490 ( .B1(n2756), .B2(n3682), .A(n2680), .ZN(n2682) );
  INV_X1 U34910 ( .A(n2681), .ZN(n3704) );
  XNOR2_X1 U3492 ( .A(n2682), .B(n3704), .ZN(n2692) );
  NAND2_X1 U34930 ( .A1(n4640), .A2(n3746), .ZN(n3817) );
  NAND2_X1 U3494 ( .A1(n2870), .A2(n4349), .ZN(n2683) );
  XNOR2_X1 U34950 ( .A(n2684), .B(IR_REG_27__SCAN_IN), .ZN(n2912) );
  NOR2_X1 U3496 ( .A1(n2685), .A2(n2686), .ZN(n2687) );
  INV_X1 U34970 ( .A(n2687), .ZN(n2688) );
  NAND2_X1 U3498 ( .A1(n4650), .A2(n2782), .ZN(n4547) );
  AOI21_X1 U34990 ( .B1(n2912), .B2(B_REG_SCAN_IN), .A(n4547), .ZN(n3885) );
  INV_X1 U3500 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U35010 ( .A1(n2886), .A2(REG2_REG_30__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3502 ( .A1(n2158), .A2(REG1_REG_30__SCAN_IN), .ZN(n2689) );
  OAI211_X1 U35030 ( .C1(n2887), .C2(n2691), .A(n2690), .B(n2689), .ZN(n3680)
         );
  AOI22_X2 U3504 ( .A1(n2692), .A2(n4789), .B1(n3885), .B2(n3680), .ZN(n2744)
         );
  INV_X1 U35050 ( .A(n2782), .ZN(n2866) );
  NOR2_X2 U35060 ( .A1(n4650), .A2(n2866), .ZN(n4549) );
  NAND2_X1 U35070 ( .A1(n4458), .A2(n4549), .ZN(n2693) );
  OAI211_X1 U35080 ( .C1(n3684), .C2(n4563), .A(n2744), .B(n2693), .ZN(n2694)
         );
  OAI21_X1 U35090 ( .B1(IR_REG_24__SCAN_IN), .B2(IR_REG_23__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2697) );
  NAND2_X1 U35100 ( .A1(n2707), .A2(n2697), .ZN(n2698) );
  NAND2_X1 U35110 ( .A1(n3432), .A2(n2705), .ZN(n2699) );
  MUX2_X1 U35120 ( .A(n3432), .B(n2699), .S(B_REG_SCAN_IN), .Z(n2702) );
  INV_X1 U35130 ( .A(n4639), .ZN(n2703) );
  NAND2_X1 U35140 ( .A1(n2705), .A2(n2703), .ZN(n2704) );
  OAI21_X1 U35150 ( .B1(n3430), .B2(D_REG_1__SCAN_IN), .A(n2704), .ZN(n2733)
         );
  NAND2_X1 U35160 ( .A1(n2708), .A2(IR_REG_23__SCAN_IN), .ZN(n2710) );
  NAND2_X1 U35170 ( .A1(n3813), .A2(n3878), .ZN(n2864) );
  NOR2_X1 U35180 ( .A1(n2734), .A2(n2736), .ZN(n2722) );
  INV_X1 U35190 ( .A(n3430), .ZN(n2721) );
  NOR4_X1 U35200 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2719) );
  NOR4_X1 U35210 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2718) );
  INV_X1 U35220 ( .A(D_REG_10__SCAN_IN), .ZN(n4831) );
  INV_X1 U35230 ( .A(D_REG_25__SCAN_IN), .ZN(n4823) );
  INV_X1 U35240 ( .A(D_REG_12__SCAN_IN), .ZN(n4830) );
  NAND4_X1 U35250 ( .A1(n4831), .A2(n4823), .A3(n4827), .A4(n4830), .ZN(n2716)
         );
  NOR4_X1 U35260 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2714) );
  NOR4_X1 U35270 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2713) );
  NOR4_X1 U35280 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2712) );
  NOR4_X1 U35290 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2711) );
  NAND4_X1 U35300 ( .A1(n2714), .A2(n2713), .A3(n2712), .A4(n2711), .ZN(n2715)
         );
  NOR4_X1 U35310 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(n2716), 
        .A4(n2715), .ZN(n2717) );
  NAND3_X1 U35320 ( .A1(n2719), .A2(n2718), .A3(n2717), .ZN(n2720) );
  NAND3_X1 U35330 ( .A1(n2733), .A2(n2722), .A3(n2861), .ZN(n2729) );
  INV_X1 U35340 ( .A(n2735), .ZN(n2863) );
  NAND2_X1 U35350 ( .A1(n3021), .A2(n2854), .ZN(n3031) );
  NAND2_X1 U35360 ( .A1(n4799), .A2(n3069), .ZN(n3068) );
  NAND2_X1 U35370 ( .A1(n4408), .A2(n4546), .ZN(n4409) );
  NAND2_X1 U35380 ( .A1(n4218), .A2(n4464), .ZN(n3896) );
  INV_X1 U35390 ( .A(n3527), .ZN(n2724) );
  INV_X1 U35400 ( .A(n2725), .ZN(n2761) );
  NAND2_X1 U35410 ( .A1(n2742), .A2(n4865), .ZN(n2728) );
  INV_X1 U35420 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2726) );
  OAI21_X1 U35430 ( .B1(n2732), .B2(n4885), .A(n2312), .ZN(U3515) );
  NAND2_X1 U35440 ( .A1(n2742), .A2(n4888), .ZN(n2731) );
  OR2_X1 U35450 ( .A1(n4898), .A2(n3941), .ZN(n2730) );
  OAI21_X1 U35460 ( .B1(n2732), .B2(n4895), .A(n2311), .ZN(U3547) );
  INV_X1 U35470 ( .A(n2733), .ZN(n2862) );
  INV_X1 U35480 ( .A(n2734), .ZN(n2876) );
  NAND4_X1 U35490 ( .A1(n2862), .A2(n2876), .A3(n2735), .A4(n2861), .ZN(n2738)
         );
  INV_X1 U35500 ( .A(n2736), .ZN(n2737) );
  OR2_X1 U35510 ( .A1(n4878), .A2(n4349), .ZN(n2856) );
  INV_X1 U35520 ( .A(n2856), .ZN(n2739) );
  INV_X1 U35530 ( .A(n2740), .ZN(n2741) );
  AOI22_X1 U35540 ( .A1(n2742), .A2(n4802), .B1(n2741), .B2(n4810), .ZN(n2743)
         );
  AOI21_X1 U35550 ( .B1(n2744), .B2(n2743), .A(n4806), .ZN(n2745) );
  NAND2_X1 U35560 ( .A1(n4815), .A2(n4549), .ZN(n3364) );
  INV_X1 U35570 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2746) );
  OAI22_X1 U35580 ( .A1(n3521), .A2(n3364), .B1(n2746), .B2(n4815), .ZN(n2749)
         );
  AND2_X1 U35590 ( .A1(n4815), .A2(n4791), .ZN(n3361) );
  AND2_X1 U35600 ( .A1(n3361), .A2(n2747), .ZN(n2748) );
  NOR2_X1 U35610 ( .A1(n2749), .A2(n2748), .ZN(n2753) );
  OR2_X1 U35620 ( .A1(n2980), .A2(n3878), .ZN(n3027) );
  NAND2_X1 U35630 ( .A1(n4435), .A2(n3027), .ZN(n2750) );
  NAND3_X1 U35640 ( .A1(n2754), .A2(n2753), .A3(n2752), .ZN(U3354) );
  XNOR2_X1 U35650 ( .A(n2756), .B(n3698), .ZN(n2757) );
  INV_X1 U35660 ( .A(n3828), .ZN(n3525) );
  OAI22_X1 U35670 ( .A1(n3525), .A2(n4547), .B1(n4563), .B2(n3527), .ZN(n2758)
         );
  AOI21_X1 U35680 ( .B1(n4549), .B2(n4466), .A(n2758), .ZN(n2759) );
  INV_X1 U35690 ( .A(n2760), .ZN(n2763) );
  INV_X1 U35700 ( .A(n3899), .ZN(n2762) );
  OAI21_X1 U35710 ( .B1(n2762), .B2(n3527), .A(n2761), .ZN(n3415) );
  NAND2_X1 U35720 ( .A1(n2763), .A2(n2326), .ZN(U3546) );
  INV_X1 U35730 ( .A(n2765), .ZN(n2766) );
  NAND2_X1 U35740 ( .A1(n2766), .A2(n2325), .ZN(U3514) );
  INV_X1 U35750 ( .A(DATAI_22_), .ZN(n2768) );
  NAND2_X1 U35760 ( .A1(n2870), .A2(STATE_REG_SCAN_IN), .ZN(n2767) );
  OAI21_X1 U35770 ( .B1(STATE_REG_SCAN_IN), .B2(n2768), .A(n2767), .ZN(U3330)
         );
  INV_X1 U35780 ( .A(DATAI_21_), .ZN(n2770) );
  NAND2_X1 U35790 ( .A1(n3746), .A2(STATE_REG_SCAN_IN), .ZN(n2769) );
  OAI21_X1 U35800 ( .B1(STATE_REG_SCAN_IN), .B2(n2770), .A(n2769), .ZN(U3331)
         );
  INV_X1 U35810 ( .A(DATAI_19_), .ZN(n2771) );
  MUX2_X1 U3582 ( .A(n2771), .B(n3878), .S(STATE_REG_SCAN_IN), .Z(n2772) );
  INV_X1 U3583 ( .A(n2772), .ZN(U3333) );
  INV_X1 U3584 ( .A(DATAI_25_), .ZN(n2775) );
  NAND2_X1 U3585 ( .A1(n2773), .A2(STATE_REG_SCAN_IN), .ZN(n2774) );
  OAI21_X1 U3586 ( .B1(STATE_REG_SCAN_IN), .B2(n2775), .A(n2774), .ZN(U3327)
         );
  INV_X1 U3587 ( .A(DATAI_24_), .ZN(n2776) );
  MUX2_X1 U3588 ( .A(n2776), .B(n3432), .S(STATE_REG_SCAN_IN), .Z(n2777) );
  INV_X1 U3589 ( .A(n2777), .ZN(U3328) );
  INV_X1 U3590 ( .A(DATAI_27_), .ZN(n4054) );
  NAND2_X1 U3591 ( .A1(n2912), .A2(STATE_REG_SCAN_IN), .ZN(n2778) );
  OAI21_X1 U3592 ( .B1(STATE_REG_SCAN_IN), .B2(n4054), .A(n2778), .ZN(U3325)
         );
  INV_X1 U3593 ( .A(DATAI_30_), .ZN(n2781) );
  NAND2_X1 U3594 ( .A1(n2779), .A2(STATE_REG_SCAN_IN), .ZN(n2780) );
  OAI21_X1 U3595 ( .B1(STATE_REG_SCAN_IN), .B2(n2781), .A(n2780), .ZN(U3322)
         );
  NOR2_X1 U3596 ( .A1(n2974), .A2(U3149), .ZN(n3821) );
  INV_X1 U3597 ( .A(n3821), .ZN(n3826) );
  NAND2_X1 U3598 ( .A1(n3428), .A2(n3826), .ZN(n2786) );
  NAND2_X1 U3599 ( .A1(n2782), .A2(n2974), .ZN(n2783) );
  NAND2_X1 U3600 ( .A1(n3666), .A2(n2783), .ZN(n2784) );
  NOR2_X1 U3601 ( .A1(n4767), .A2(U4043), .ZN(U3148) );
  INV_X1 U3602 ( .A(n4767), .ZN(n2793) );
  INV_X1 U3603 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n2792) );
  INV_X1 U3604 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4814) );
  AOI21_X1 U3605 ( .B1(n2912), .B2(n4814), .A(n4650), .ZN(n2915) );
  OAI21_X1 U3606 ( .B1(n2912), .B2(REG1_REG_0__SCAN_IN), .A(n2270), .ZN(n2788)
         );
  INV_X1 U3607 ( .A(n2784), .ZN(n2785) );
  NOR2_X1 U3608 ( .A1(n2915), .A2(IR_REG_0__SCAN_IN), .ZN(n2787) );
  AOI211_X1 U3609 ( .C1(n2915), .C2(n2788), .A(n2811), .B(n2787), .ZN(n2789)
         );
  AOI21_X1 U3610 ( .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .A(n2789), .ZN(n2791)
         );
  INV_X1 U3611 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2795) );
  NAND3_X1 U3612 ( .A1(n4771), .A2(n2795), .A3(IR_REG_0__SCAN_IN), .ZN(n2790)
         );
  OAI211_X1 U3613 ( .C1(n2793), .C2(n2792), .A(n2791), .B(n2790), .ZN(U3240)
         );
  INV_X1 U3614 ( .A(n2823), .ZN(n4644) );
  INV_X1 U3615 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2794) );
  MUX2_X1 U3616 ( .A(REG1_REG_1__SCAN_IN), .B(n2794), .S(n2836), .Z(n2830) );
  INV_X1 U3617 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2796) );
  MUX2_X1 U3618 ( .A(n2796), .B(REG1_REG_2__SCAN_IN), .S(n4647), .Z(n2932) );
  INV_X1 U3619 ( .A(n2797), .ZN(n2798) );
  INV_X1 U3620 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2844) );
  OAI21_X1 U3621 ( .B1(n2798), .B2(n2389), .A(n2841), .ZN(n2799) );
  XOR2_X1 U3622 ( .A(REG1_REG_5__SCAN_IN), .B(n2823), .Z(n2819) );
  AOI21_X1 U3623 ( .B1(REG1_REG_5__SCAN_IN), .B2(n4644), .A(n2818), .ZN(n3197)
         );
  XOR2_X1 U3624 ( .A(n4643), .B(n3197), .Z(n2801) );
  NOR2_X1 U3625 ( .A1(n2801), .A2(n3998), .ZN(n3196) );
  AOI211_X1 U3626 ( .C1(n3998), .C2(n2801), .A(n4756), .B(n3196), .ZN(n2817)
         );
  INV_X1 U3627 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2810) );
  NAND2_X1 U3628 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2914) );
  NOR2_X1 U3629 ( .A1(n2828), .A2(n2914), .ZN(n2827) );
  INV_X1 U3630 ( .A(n2839), .ZN(n2804) );
  INV_X1 U3631 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2840) );
  NAND2_X1 U3632 ( .A1(n2804), .A2(REG2_REG_3__SCAN_IN), .ZN(n2837) );
  OAI21_X1 U3633 ( .B1(n2805), .B2(n2389), .A(n2837), .ZN(n2806) );
  INV_X1 U3634 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2920) );
  INV_X1 U3635 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2967) );
  XNOR2_X1 U3636 ( .A(n2823), .B(n2967), .ZN(n2821) );
  AOI21_X1 U3637 ( .B1(REG2_REG_5__SCAN_IN), .B2(n4644), .A(n2820), .ZN(n3181)
         );
  XNOR2_X1 U3638 ( .A(n3181), .B(n2807), .ZN(n2809) );
  INV_X1 U3639 ( .A(n4650), .ZN(n2998) );
  NAND2_X1 U3640 ( .A1(n2998), .A2(n2912), .ZN(n3824) );
  INV_X1 U3641 ( .A(n3182), .ZN(n2808) );
  AOI211_X1 U3642 ( .C1(n2810), .C2(n2809), .A(n4754), .B(n2808), .ZN(n2816)
         );
  INV_X1 U3643 ( .A(n2811), .ZN(n2812) );
  NOR2_X1 U3644 ( .A1(STATE_REG_SCAN_IN), .A2(n2813), .ZN(n3085) );
  AOI21_X1 U3645 ( .B1(n4767), .B2(ADDR_REG_6__SCAN_IN), .A(n3085), .ZN(n2814)
         );
  OAI21_X1 U3646 ( .B1(n4775), .B2(n2807), .A(n2814), .ZN(n2815) );
  OR3_X1 U3647 ( .A1(n2817), .A2(n2816), .A3(n2815), .ZN(U3246) );
  AOI211_X1 U3648 ( .C1(n2198), .C2(n2819), .A(n4756), .B(n2818), .ZN(n2826)
         );
  AOI211_X1 U3649 ( .C1(n2197), .C2(n2821), .A(n4754), .B(n2820), .ZN(n2825)
         );
  AND2_X1 U3650 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3055) );
  AOI21_X1 U3651 ( .B1(n4767), .B2(ADDR_REG_5__SCAN_IN), .A(n3055), .ZN(n2822)
         );
  OAI21_X1 U3652 ( .B1(n4775), .B2(n2823), .A(n2822), .ZN(n2824) );
  OR3_X1 U3653 ( .A1(n2826), .A2(n2825), .A3(n2824), .ZN(U3245) );
  AOI211_X1 U3654 ( .C1(n2914), .C2(n2828), .A(n2827), .B(n4754), .ZN(n2833)
         );
  NAND2_X1 U3655 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2831) );
  AOI211_X1 U3656 ( .C1(n2831), .C2(n2830), .A(n2829), .B(n4756), .ZN(n2832)
         );
  NOR2_X1 U3657 ( .A1(n2833), .A2(n2832), .ZN(n2835) );
  AOI22_X1 U3658 ( .A1(n4767), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n2834) );
  OAI211_X1 U3659 ( .C1(n2836), .C2(n4775), .A(n2835), .B(n2834), .ZN(U3241)
         );
  INV_X1 U3660 ( .A(n2837), .ZN(n2838) );
  AOI211_X1 U3661 ( .C1(n2840), .C2(n2839), .A(n2838), .B(n4754), .ZN(n2846)
         );
  INV_X1 U3662 ( .A(n2841), .ZN(n2842) );
  AOI211_X1 U3663 ( .C1(n2844), .C2(n2843), .A(n2842), .B(n4756), .ZN(n2845)
         );
  NOR2_X1 U3664 ( .A1(n2846), .A2(n2845), .ZN(n2848) );
  INV_X1 U3665 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4798) );
  NOR2_X1 U3666 ( .A1(STATE_REG_SCAN_IN), .A2(n4798), .ZN(n3001) );
  AOI21_X1 U3667 ( .B1(n4767), .B2(ADDR_REG_3__SCAN_IN), .A(n3001), .ZN(n2847)
         );
  OAI211_X1 U3668 ( .C1(n2389), .C2(n4775), .A(n2848), .B(n2847), .ZN(U3243)
         );
  NAND2_X1 U3669 ( .A1(n2858), .A2(n2854), .ZN(n3744) );
  INV_X1 U3670 ( .A(n3701), .ZN(n4812) );
  INV_X1 U3671 ( .A(n2873), .ZN(n2849) );
  NOR2_X1 U3672 ( .A1(n2854), .A2(n2849), .ZN(n4809) );
  INV_X1 U3673 ( .A(n4435), .ZN(n4797) );
  NOR2_X1 U3674 ( .A1(n4797), .A2(n4789), .ZN(n2850) );
  OAI22_X1 U3675 ( .A1(n3701), .A2(n2850), .B1(n3365), .B2(n4547), .ZN(n4807)
         );
  AOI211_X1 U3676 ( .C1(n4883), .C2(n4812), .A(n4809), .B(n4807), .ZN(n4857)
         );
  NAND2_X1 U3677 ( .A1(n4895), .A2(REG1_REG_0__SCAN_IN), .ZN(n2851) );
  OAI21_X1 U3678 ( .B1(n4857), .B2(n4895), .A(n2851), .ZN(U3518) );
  INV_X1 U3679 ( .A(n2853), .ZN(n2857) );
  INV_X1 U3680 ( .A(n2980), .ZN(n2852) );
  OAI22_X1 U3681 ( .A1(n2855), .A2(n2162), .B1(n3519), .B2(n2854), .ZN(n2978)
         );
  AOI222_X1 U3682 ( .A1(n2858), .A2(n3483), .B1(n3029), .B2(n2176), .C1(
        IR_REG_0__SCAN_IN), .C2(n2857), .ZN(n2859) );
  NOR2_X1 U3683 ( .A1(n2860), .A2(n2859), .ZN(n2981) );
  AOI21_X1 U3684 ( .B1(n2860), .B2(n2859), .A(n2981), .ZN(n2913) );
  NAND3_X1 U3685 ( .A1(n2863), .A2(n2862), .A3(n2861), .ZN(n2875) );
  NAND2_X1 U3686 ( .A1(n2864), .A2(n2873), .ZN(n2865) );
  NAND2_X1 U3687 ( .A1(n2866), .A2(n2865), .ZN(n2867) );
  OR2_X1 U3688 ( .A1(n3428), .A2(n2867), .ZN(n2868) );
  NOR3_X1 U3689 ( .A1(n2875), .A2(n4563), .A3(n3428), .ZN(n2869) );
  NOR2_X2 U3690 ( .A1(n2869), .A2(n4810), .ZN(n3652) );
  AOI22_X1 U3691 ( .A1(n2913), .A2(n4663), .B1(n3029), .B2(n4656), .ZN(n2878)
         );
  NAND2_X1 U3692 ( .A1(n2870), .A2(n3878), .ZN(n2979) );
  INV_X1 U3693 ( .A(n2979), .ZN(n2871) );
  NAND3_X1 U3694 ( .A1(n2176), .A2(n4836), .A3(n2871), .ZN(n3823) );
  NOR2_X1 U3695 ( .A1(n2875), .A2(n3823), .ZN(n2999) );
  NAND2_X2 U3696 ( .A1(n2999), .A2(n4650), .ZN(n3659) );
  INV_X1 U3697 ( .A(n3659), .ZN(n3631) );
  NAND3_X1 U3698 ( .A1(n4563), .A2(n2873), .A3(n4349), .ZN(n2874) );
  NAND2_X1 U3699 ( .A1(n2875), .A2(n2874), .ZN(n2976) );
  NAND2_X1 U3700 ( .A1(n2976), .A2(n2876), .ZN(n3628) );
  AOI22_X1 U3701 ( .A1(n3631), .A2(n2872), .B1(REG3_REG_0__SCAN_IN), .B2(n3628), .ZN(n2877) );
  NAND2_X1 U3702 ( .A1(n2878), .A2(n2877), .ZN(U3229) );
  INV_X1 U3703 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n2880) );
  NAND2_X1 U3704 ( .A1(n4232), .A2(U4043), .ZN(n2879) );
  OAI21_X1 U3705 ( .B1(U4043), .B2(n2880), .A(n2879), .ZN(U3575) );
  INV_X1 U3706 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U3707 ( .A1(n3537), .A2(U4043), .ZN(n2881) );
  OAI21_X1 U3708 ( .B1(U4043), .B2(n2882), .A(n2881), .ZN(U3552) );
  INV_X1 U3709 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n2884) );
  NAND2_X1 U3710 ( .A1(n4429), .A2(U4043), .ZN(n2883) );
  OAI21_X1 U3711 ( .B1(U4043), .B2(n2884), .A(n2883), .ZN(U3564) );
  INV_X1 U3712 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n2892) );
  NAND2_X1 U3713 ( .A1(n2159), .A2(REG1_REG_31__SCAN_IN), .ZN(n2890) );
  NAND2_X1 U3714 ( .A1(n2886), .A2(REG2_REG_31__SCAN_IN), .ZN(n2889) );
  INV_X1 U3715 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4576) );
  OR2_X1 U3716 ( .A1(n2887), .A2(n4576), .ZN(n2888) );
  NAND2_X1 U3717 ( .A1(n3886), .A2(U4043), .ZN(n2891) );
  OAI21_X1 U3718 ( .B1(U4043), .B2(n2892), .A(n2891), .ZN(U3581) );
  INV_X1 U3719 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n2894) );
  NAND2_X1 U3720 ( .A1(n3680), .A2(U4043), .ZN(n2893) );
  OAI21_X1 U3721 ( .B1(U4043), .B2(n2894), .A(n2893), .ZN(U3580) );
  INV_X1 U3722 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n2896) );
  NAND2_X1 U3723 ( .A1(n4466), .A2(U4043), .ZN(n2895) );
  OAI21_X1 U3724 ( .B1(U4043), .B2(n2896), .A(n2895), .ZN(U3577) );
  INV_X1 U3725 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n2898) );
  NAND2_X1 U3726 ( .A1(n4529), .A2(U4043), .ZN(n2897) );
  OAI21_X1 U3727 ( .B1(U4043), .B2(n2898), .A(n2897), .ZN(U3567) );
  INV_X1 U3728 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n2900) );
  NAND2_X1 U3729 ( .A1(n4483), .A2(U4043), .ZN(n2899) );
  OAI21_X1 U3730 ( .B1(U4043), .B2(n2900), .A(n2899), .ZN(U3573) );
  INV_X1 U3731 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U3732 ( .A1(n2901), .A2(U4043), .ZN(n2902) );
  OAI21_X1 U3733 ( .B1(U4043), .B2(n2903), .A(n2902), .ZN(U3571) );
  INV_X1 U3734 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n2905) );
  NAND2_X1 U3735 ( .A1(n3229), .A2(U4043), .ZN(n2904) );
  OAI21_X1 U3736 ( .B1(U4043), .B2(n2905), .A(n2904), .ZN(U3562) );
  INV_X1 U3737 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n2907) );
  NAND2_X1 U3738 ( .A1(n3092), .A2(U4043), .ZN(n2906) );
  OAI21_X1 U3739 ( .B1(U4043), .B2(n2907), .A(n2906), .ZN(U3555) );
  INV_X1 U3740 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n2909) );
  NAND2_X1 U3741 ( .A1(n4539), .A2(U4043), .ZN(n2908) );
  OAI21_X1 U3742 ( .B1(U4043), .B2(n2909), .A(n2908), .ZN(U3566) );
  INV_X1 U3743 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n2911) );
  NAND2_X1 U3744 ( .A1(n4345), .A2(U4043), .ZN(n2910) );
  OAI21_X1 U3745 ( .B1(U4043), .B2(n2911), .A(n2910), .ZN(U3569) );
  NOR3_X1 U3746 ( .A1(n2913), .A2(n2912), .A3(n4650), .ZN(n2917) );
  OAI22_X1 U3747 ( .A1(n2915), .A2(IR_REG_0__SCAN_IN), .B1(n2914), .B2(n3824), 
        .ZN(n2916) );
  NOR3_X1 U3748 ( .A1(n2917), .A2(n3836), .A3(n2916), .ZN(n2939) );
  AOI211_X1 U3749 ( .C1(n2920), .C2(n2919), .A(n2918), .B(n4754), .ZN(n2927)
         );
  AOI211_X1 U3750 ( .C1(n4892), .C2(n2922), .A(n4756), .B(n2921), .ZN(n2926)
         );
  INV_X1 U3751 ( .A(n4645), .ZN(n2924) );
  AND2_X1 U3752 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3016) );
  AOI21_X1 U3753 ( .B1(n4767), .B2(ADDR_REG_4__SCAN_IN), .A(n3016), .ZN(n2923)
         );
  OAI21_X1 U3754 ( .B1(n4775), .B2(n2924), .A(n2923), .ZN(n2925) );
  OR4_X1 U3755 ( .A1(n2939), .A2(n2927), .A3(n2926), .A4(n2925), .ZN(U3244) );
  AOI211_X1 U3756 ( .C1(n2930), .C2(n2929), .A(n2928), .B(n4754), .ZN(n2938)
         );
  AOI211_X1 U3757 ( .C1(n2933), .C2(n2932), .A(n2931), .B(n4756), .ZN(n2937)
         );
  INV_X1 U3758 ( .A(n2161), .ZN(n2935) );
  AOI22_X1 U3759 ( .A1(n4767), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2934) );
  OAI21_X1 U3760 ( .B1(n4775), .B2(n2935), .A(n2934), .ZN(n2936) );
  OR4_X1 U3761 ( .A1(n2939), .A2(n2938), .A3(n2937), .A4(n2936), .ZN(U3242) );
  NAND2_X1 U3762 ( .A1(n2941), .A2(n2945), .ZN(n2942) );
  NAND2_X1 U3763 ( .A1(n2940), .A2(n2942), .ZN(n3360) );
  NOR2_X1 U3764 ( .A1(n2988), .A2(n4563), .ZN(n2943) );
  AOI21_X1 U3765 ( .B1(n3835), .B2(n4792), .A(n2943), .ZN(n2944) );
  OAI21_X1 U3766 ( .B1(n3365), .B2(n4796), .A(n2944), .ZN(n2951) );
  NAND2_X1 U3767 ( .A1(n3360), .A2(n4797), .ZN(n2950) );
  NAND3_X1 U3768 ( .A1(n2650), .A2(n3023), .A3(n2649), .ZN(n2946) );
  NAND2_X1 U3769 ( .A1(n2947), .A2(n2946), .ZN(n2948) );
  NAND2_X1 U3770 ( .A1(n2948), .A2(n4789), .ZN(n2949) );
  NAND2_X1 U3771 ( .A1(n2950), .A2(n2949), .ZN(n3355) );
  AOI211_X1 U3772 ( .C1(n4883), .C2(n3360), .A(n2951), .B(n3355), .ZN(n2957)
         );
  INV_X1 U3773 ( .A(n2952), .ZN(n4800) );
  NAND2_X1 U3774 ( .A1(n3031), .A2(n3629), .ZN(n2953) );
  NAND2_X1 U3775 ( .A1(n4800), .A2(n2953), .ZN(n3356) );
  INV_X1 U3776 ( .A(n3356), .ZN(n2955) );
  AOI22_X1 U3777 ( .A1(n4888), .A2(n2955), .B1(n4895), .B2(REG1_REG_2__SCAN_IN), .ZN(n2954) );
  OAI21_X1 U3778 ( .B1(n2957), .B2(n4895), .A(n2954), .ZN(U3520) );
  AOI22_X1 U3779 ( .A1(n4865), .A2(n2955), .B1(n4885), .B2(REG0_REG_2__SCAN_IN), .ZN(n2956) );
  OAI21_X1 U3780 ( .B1(n2957), .B2(n4885), .A(n2956), .ZN(U3471) );
  INV_X1 U3781 ( .A(n2958), .ZN(n3755) );
  NAND2_X1 U3782 ( .A1(n3755), .A2(n3768), .ZN(n3729) );
  XNOR2_X1 U3783 ( .A(n2959), .B(n3729), .ZN(n2960) );
  NAND2_X1 U3784 ( .A1(n2960), .A2(n4789), .ZN(n3038) );
  NAND2_X1 U3785 ( .A1(n2961), .A2(n2962), .ZN(n3061) );
  NAND2_X1 U3786 ( .A1(n3061), .A2(n2963), .ZN(n2964) );
  XOR2_X1 U3787 ( .A(n3729), .B(n2964), .Z(n3040) );
  AND2_X1 U3788 ( .A1(n3068), .A2(n3056), .ZN(n2965) );
  NOR2_X1 U3789 ( .A1(n3098), .A2(n2965), .ZN(n3042) );
  INV_X1 U3790 ( .A(n2966), .ZN(n3059) );
  OAI22_X1 U3791 ( .A1(n4815), .A2(n2967), .B1(n3059), .B2(n4350), .ZN(n2968)
         );
  AOI21_X1 U3792 ( .B1(n3042), .B2(n4802), .A(n2968), .ZN(n2970) );
  AND2_X1 U3793 ( .A1(n4815), .A2(n4792), .ZN(n4411) );
  AOI22_X1 U3794 ( .A1(n3361), .A2(n3056), .B1(n4411), .B2(n3834), .ZN(n2969)
         );
  OAI211_X1 U3795 ( .C1(n3053), .C2(n3364), .A(n2970), .B(n2969), .ZN(n2971)
         );
  AOI21_X1 U3796 ( .B1(n3040), .B2(n4407), .A(n2971), .ZN(n2972) );
  OAI21_X1 U3797 ( .B1(n4806), .B2(n3038), .A(n2972), .ZN(U3285) );
  INV_X1 U3798 ( .A(n2973), .ZN(n2975) );
  NAND4_X1 U3799 ( .A1(n2976), .A2(n2975), .A3(n2853), .A4(n2974), .ZN(n2977)
         );
  INV_X1 U3800 ( .A(n2978), .ZN(n2982) );
  AOI21_X1 U3801 ( .B1(n2982), .B2(n3480), .A(n2981), .ZN(n3534) );
  INV_X2 U3802 ( .A(n3480), .ZN(n3011) );
  XNOR2_X1 U3803 ( .A(n2983), .B(n3011), .ZN(n2985) );
  OAI22_X1 U3804 ( .A1(n3365), .A2(n2984), .B1(n3021), .B2(n2162), .ZN(n2986)
         );
  XNOR2_X1 U3805 ( .A(n2985), .B(n2986), .ZN(n3533) );
  NOR2_X1 U3806 ( .A1(n3534), .A2(n3533), .ZN(n3532) );
  NOR2_X1 U3807 ( .A1(n3532), .A2(n2987), .ZN(n3624) );
  OAI22_X1 U3808 ( .A1(n2374), .A2(n2984), .B1(n2988), .B2(n2162), .ZN(n2990)
         );
  OAI22_X1 U3809 ( .A1(n2374), .A2(n2162), .B1(n2988), .B2(n3519), .ZN(n2989)
         );
  XNOR2_X1 U3810 ( .A(n2989), .B(n3011), .ZN(n2991) );
  XOR2_X1 U3811 ( .A(n2990), .B(n2991), .Z(n3626) );
  NAND2_X1 U3812 ( .A1(n3624), .A2(n3626), .ZN(n3625) );
  OR2_X1 U3813 ( .A1(n2991), .A2(n2990), .ZN(n2992) );
  NAND2_X1 U3814 ( .A1(n3625), .A2(n2992), .ZN(n3010) );
  OAI22_X1 U3815 ( .A1(n3358), .A2(n2984), .B1(n2162), .B2(n2993), .ZN(n3005)
         );
  NAND2_X1 U3816 ( .A1(n3835), .A2(n2176), .ZN(n2995) );
  NAND2_X1 U3817 ( .A1(n4801), .A2(n3477), .ZN(n2994) );
  NAND2_X1 U3818 ( .A1(n2995), .A2(n2994), .ZN(n2996) );
  XNOR2_X1 U3819 ( .A(n2996), .B(n3011), .ZN(n3006) );
  XOR2_X1 U3820 ( .A(n3005), .B(n3006), .Z(n3009) );
  XNOR2_X1 U3821 ( .A(n3010), .B(n3009), .ZN(n2997) );
  NAND2_X1 U3822 ( .A1(n2997), .A2(n4663), .ZN(n3003) );
  NAND2_X2 U3823 ( .A1(n2999), .A2(n2998), .ZN(n4653) );
  OAI22_X1 U3824 ( .A1(n2374), .A2(n4653), .B1(n3659), .B2(n3053), .ZN(n3000)
         );
  AOI211_X1 U3825 ( .C1(n4801), .C2(n4656), .A(n3001), .B(n3000), .ZN(n3002)
         );
  OAI211_X1 U3826 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4668), .A(n3003), .B(n3002), 
        .ZN(U3215) );
  INV_X1 U3827 ( .A(n3004), .ZN(n3070) );
  INV_X1 U3828 ( .A(n3005), .ZN(n3008) );
  INV_X1 U3829 ( .A(n3006), .ZN(n3007) );
  AOI22_X1 U3830 ( .A1(n3010), .A2(n3009), .B1(n3008), .B2(n3007), .ZN(n3014)
         );
  OAI22_X1 U3831 ( .A1(n3053), .A2(n2984), .B1(n2162), .B2(n3069), .ZN(n3046)
         );
  OAI22_X1 U3832 ( .A1(n3053), .A2(n2162), .B1(n3519), .B2(n3069), .ZN(n3012)
         );
  XNOR2_X1 U3833 ( .A(n3012), .B(n3011), .ZN(n3045) );
  XOR2_X1 U3834 ( .A(n3046), .B(n3045), .Z(n3013) );
  NAND2_X1 U3835 ( .A1(n3014), .A2(n3013), .ZN(n3048) );
  OAI211_X1 U3836 ( .C1(n3014), .C2(n3013), .A(n3048), .B(n4663), .ZN(n3019)
         );
  OAI22_X1 U3837 ( .A1(n3083), .A2(n3659), .B1(n4653), .B2(n3358), .ZN(n3015)
         );
  AOI211_X1 U3838 ( .C1(n3017), .C2(n4656), .A(n3016), .B(n3015), .ZN(n3018)
         );
  OAI211_X1 U3839 ( .C1(n4668), .C2(n3070), .A(n3019), .B(n3018), .ZN(U3227)
         );
  XNOR2_X1 U3840 ( .A(n2648), .B(n3020), .ZN(n4860) );
  OAI22_X1 U3841 ( .A1(n2374), .A2(n4547), .B1(n4563), .B2(n3021), .ZN(n3025)
         );
  NAND2_X1 U3842 ( .A1(n2648), .A2(n3743), .ZN(n3022) );
  AOI21_X1 U3843 ( .B1(n3023), .B2(n3022), .A(n4551), .ZN(n3024) );
  AOI211_X1 U3844 ( .C1(n4549), .C2(n2858), .A(n3025), .B(n3024), .ZN(n3026)
         );
  OAI21_X1 U3845 ( .B1(n4860), .B2(n4435), .A(n3026), .ZN(n4862) );
  INV_X1 U3846 ( .A(n4862), .ZN(n3036) );
  INV_X1 U3847 ( .A(n4860), .ZN(n3034) );
  INV_X1 U3848 ( .A(n3027), .ZN(n3028) );
  NAND2_X1 U3849 ( .A1(n3536), .A2(n3029), .ZN(n3030) );
  NAND2_X1 U3850 ( .A1(n3031), .A2(n3030), .ZN(n4858) );
  AOI22_X1 U3851 ( .A1(n4806), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4810), .ZN(n3032) );
  OAI21_X1 U3852 ( .B1(n4441), .B2(n4858), .A(n3032), .ZN(n3033) );
  AOI21_X1 U3853 ( .B1(n3034), .B2(n4811), .A(n3033), .ZN(n3035) );
  OAI21_X1 U3854 ( .B1(n3036), .B2(n4806), .A(n3035), .ZN(U3289) );
  AOI22_X1 U3855 ( .A1(n3834), .A2(n4792), .B1(n4791), .B2(n3056), .ZN(n3037)
         );
  OAI211_X1 U3856 ( .C1(n3053), .C2(n4796), .A(n3038), .B(n3037), .ZN(n3039)
         );
  AOI21_X1 U3857 ( .B1(n3040), .B2(n4873), .A(n3039), .ZN(n3044) );
  AOI22_X1 U3858 ( .A1(n3042), .A2(n4865), .B1(REG0_REG_5__SCAN_IN), .B2(n4885), .ZN(n3041) );
  OAI21_X1 U3859 ( .B1(n3044), .B2(n4885), .A(n3041), .ZN(U3477) );
  AOI22_X1 U3860 ( .A1(n3042), .A2(n4888), .B1(REG1_REG_5__SCAN_IN), .B2(n4895), .ZN(n3043) );
  OAI21_X1 U3861 ( .B1(n3044), .B2(n4895), .A(n3043), .ZN(U3523) );
  NAND2_X1 U3862 ( .A1(n3048), .A2(n3047), .ZN(n3052) );
  OAI22_X1 U3863 ( .A1(n3083), .A2(n2984), .B1(n3049), .B2(n2162), .ZN(n3076)
         );
  OAI22_X1 U3864 ( .A1(n3083), .A2(n2162), .B1(n3049), .B2(n3519), .ZN(n3050)
         );
  XNOR2_X1 U3865 ( .A(n3050), .B(n3011), .ZN(n3075) );
  XOR2_X1 U3866 ( .A(n3076), .B(n3075), .Z(n3051) );
  OAI211_X1 U3867 ( .C1(n3052), .C2(n3051), .A(n3079), .B(n4663), .ZN(n3058)
         );
  OAI22_X1 U3868 ( .A1(n3053), .A2(n4653), .B1(n3659), .B2(n3142), .ZN(n3054)
         );
  AOI211_X1 U3869 ( .C1(n3056), .C2(n4656), .A(n3055), .B(n3054), .ZN(n3057)
         );
  OAI211_X1 U3870 ( .C1(n4668), .C2(n3059), .A(n3058), .B(n3057), .ZN(U3224)
         );
  OR2_X1 U3871 ( .A1(n2961), .A2(n2962), .ZN(n3060) );
  NAND2_X1 U3872 ( .A1(n3061), .A2(n3060), .ZN(n4867) );
  INV_X1 U3873 ( .A(n4811), .ZN(n3074) );
  XNOR2_X1 U3874 ( .A(n3062), .B(n2962), .ZN(n3067) );
  NAND2_X1 U3875 ( .A1(n3835), .A2(n4549), .ZN(n3063) );
  OAI21_X1 U3876 ( .B1(n4563), .B2(n3069), .A(n3063), .ZN(n3065) );
  NOR2_X1 U3877 ( .A1(n4867), .A2(n4435), .ZN(n3064) );
  AOI211_X1 U3878 ( .C1(n4792), .C2(n3092), .A(n3065), .B(n3064), .ZN(n3066)
         );
  OAI21_X1 U3879 ( .B1(n4551), .B2(n3067), .A(n3066), .ZN(n4869) );
  INV_X1 U3880 ( .A(n4878), .ZN(n4532) );
  OAI211_X1 U3881 ( .C1(n4799), .C2(n3069), .A(n4532), .B(n3068), .ZN(n4868)
         );
  OAI22_X1 U3882 ( .A1(n4868), .A2(n4349), .B1(n4350), .B2(n3070), .ZN(n3071)
         );
  OAI21_X1 U3883 ( .B1(n4869), .B2(n3071), .A(n4815), .ZN(n3073) );
  NAND2_X1 U3884 ( .A1(n4806), .A2(REG2_REG_4__SCAN_IN), .ZN(n3072) );
  OAI211_X1 U3885 ( .C1(n4867), .C2(n3074), .A(n3073), .B(n3072), .ZN(U3286)
         );
  INV_X1 U3886 ( .A(n3075), .ZN(n3078) );
  INV_X1 U3887 ( .A(n3076), .ZN(n3077) );
  OAI22_X1 U3888 ( .A1(n3142), .A2(n2162), .B1(n3519), .B2(n3097), .ZN(n3080)
         );
  XNOR2_X1 U3889 ( .A(n3080), .B(n3011), .ZN(n3137) );
  OAI22_X1 U3890 ( .A1(n3142), .A2(n2984), .B1(n2162), .B2(n3097), .ZN(n3138)
         );
  INV_X1 U3891 ( .A(n3138), .ZN(n3140) );
  XNOR2_X1 U3892 ( .A(n3137), .B(n3140), .ZN(n3081) );
  XNOR2_X1 U3893 ( .A(n3139), .B(n3081), .ZN(n3088) );
  OAI22_X1 U3894 ( .A1(n3083), .A2(n4653), .B1(n3659), .B2(n3082), .ZN(n3084)
         );
  AOI211_X1 U3895 ( .C1(n3091), .C2(n4656), .A(n3085), .B(n3084), .ZN(n3087)
         );
  NAND2_X1 U3896 ( .A1(n3661), .A2(n4776), .ZN(n3086) );
  OAI211_X1 U3897 ( .C1(n3088), .C2(n3664), .A(n3087), .B(n3086), .ZN(U3236)
         );
  NAND2_X1 U3898 ( .A1(n3759), .A2(n3770), .ZN(n3694) );
  XNOR2_X1 U3899 ( .A(n3089), .B(n3694), .ZN(n4777) );
  XOR2_X1 U3900 ( .A(n3694), .B(n3090), .Z(n3096) );
  AOI22_X1 U3901 ( .A1(n3092), .A2(n4549), .B1(n3091), .B2(n4791), .ZN(n3093)
         );
  OAI21_X1 U3902 ( .B1(n3082), .B2(n4547), .A(n3093), .ZN(n3095) );
  NOR2_X1 U3903 ( .A1(n4777), .A2(n4435), .ZN(n3094) );
  AOI211_X1 U3904 ( .C1(n3096), .C2(n4789), .A(n3095), .B(n3094), .ZN(n4783)
         );
  OAI21_X1 U3905 ( .B1(n4859), .B2(n4777), .A(n4783), .ZN(n3103) );
  OR2_X1 U3906 ( .A1(n3098), .A2(n3097), .ZN(n3099) );
  NAND2_X1 U3907 ( .A1(n3148), .A2(n3099), .ZN(n4778) );
  OAI22_X1 U3908 ( .A1(n4778), .A2(n4632), .B1(n4886), .B2(n2416), .ZN(n3100)
         );
  AOI21_X1 U3909 ( .B1(n3103), .B2(n4886), .A(n3100), .ZN(n3101) );
  INV_X1 U3910 ( .A(n3101), .ZN(U3479) );
  OAI22_X1 U3911 ( .A1(n4778), .A2(n4561), .B1(n4898), .B2(n3998), .ZN(n3102)
         );
  AOI21_X1 U3912 ( .B1(n3103), .B2(n4898), .A(n3102), .ZN(n3104) );
  INV_X1 U3913 ( .A(n3104), .ZN(U3524) );
  NAND2_X1 U3914 ( .A1(n4874), .A2(n3108), .ZN(n3109) );
  NAND2_X1 U3915 ( .A1(n3763), .A2(n3771), .ZN(n3695) );
  XNOR2_X1 U3916 ( .A(n3109), .B(n3695), .ZN(n3115) );
  XNOR2_X1 U3917 ( .A(n3110), .B(n3695), .ZN(n3113) );
  AOI22_X1 U3918 ( .A1(n3831), .A2(n4792), .B1(n4791), .B2(n2436), .ZN(n3111)
         );
  OAI21_X1 U3919 ( .B1(n3082), .B2(n4796), .A(n3111), .ZN(n3112) );
  AOI21_X1 U3920 ( .B1(n3113), .B2(n4789), .A(n3112), .ZN(n3114) );
  OAI21_X1 U3921 ( .B1(n3115), .B2(n4435), .A(n3114), .ZN(n4881) );
  INV_X1 U3922 ( .A(n4881), .ZN(n3122) );
  INV_X1 U3923 ( .A(n3115), .ZN(n4884) );
  INV_X1 U3924 ( .A(n3116), .ZN(n3147) );
  NOR2_X1 U3925 ( .A1(n3147), .A2(n3170), .ZN(n4880) );
  INV_X1 U3926 ( .A(n3125), .ZN(n4879) );
  NOR3_X1 U3927 ( .A1(n4880), .A2(n4879), .A3(n4441), .ZN(n3120) );
  INV_X1 U3928 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3118) );
  INV_X1 U3929 ( .A(n3177), .ZN(n3117) );
  OAI22_X1 U3930 ( .A1(n4815), .A2(n3118), .B1(n3117), .B2(n4350), .ZN(n3119)
         );
  AOI211_X1 U3931 ( .C1(n4884), .C2(n4811), .A(n3120), .B(n3119), .ZN(n3121)
         );
  OAI21_X1 U3932 ( .B1(n3122), .B2(n4806), .A(n3121), .ZN(U3282) );
  INV_X1 U3933 ( .A(n3766), .ZN(n3772) );
  NAND2_X1 U3934 ( .A1(n3772), .A2(n3764), .ZN(n3731) );
  XNOR2_X1 U3935 ( .A(n3123), .B(n3731), .ZN(n3124) );
  NAND2_X1 U3936 ( .A1(n3124), .A2(n4789), .ZN(n3237) );
  AOI21_X1 U3937 ( .B1(n3269), .B2(n3125), .A(n3247), .ZN(n3244) );
  AOI22_X1 U3938 ( .A1(n4412), .A2(n3832), .B1(n4411), .B2(n3830), .ZN(n3128)
         );
  NOR2_X1 U3939 ( .A1(n3272), .A2(n4350), .ZN(n3126) );
  AOI21_X1 U3940 ( .B1(n4806), .B2(REG2_REG_9__SCAN_IN), .A(n3126), .ZN(n3127)
         );
  OAI211_X1 U3941 ( .C1(n3262), .C2(n4416), .A(n3128), .B(n3127), .ZN(n3129)
         );
  AOI21_X1 U3942 ( .B1(n3244), .B2(n4802), .A(n3129), .ZN(n3136) );
  OR2_X1 U3943 ( .A1(n3105), .A2(n3130), .ZN(n3132) );
  NAND2_X1 U3944 ( .A1(n3132), .A2(n3131), .ZN(n3134) );
  INV_X1 U3945 ( .A(n3731), .ZN(n3133) );
  XNOR2_X1 U3946 ( .A(n3134), .B(n3133), .ZN(n3234) );
  NAND2_X1 U3947 ( .A1(n3234), .A2(n4407), .ZN(n3135) );
  OAI211_X1 U3948 ( .C1(n3237), .C2(n4806), .A(n3136), .B(n3135), .ZN(U3281)
         );
  OAI22_X1 U3949 ( .A1(n3082), .A2(n2984), .B1(n2162), .B2(n3150), .ZN(n3163)
         );
  OAI22_X1 U3950 ( .A1(n3082), .A2(n2162), .B1(n3519), .B2(n3150), .ZN(n3141)
         );
  XNOR2_X1 U3951 ( .A(n3141), .B(n3011), .ZN(n3162) );
  XOR2_X1 U3952 ( .A(n3163), .B(n3162), .Z(n3167) );
  XNOR2_X1 U3953 ( .A(n3168), .B(n3167), .ZN(n3146) );
  NOR2_X1 U3954 ( .A1(STATE_REG_SCAN_IN), .A2(n2440), .ZN(n3840) );
  OAI22_X1 U3955 ( .A1(n3267), .A2(n3659), .B1(n4653), .B2(n3142), .ZN(n3143)
         );
  AOI211_X1 U3956 ( .C1(n3149), .C2(n4656), .A(n3840), .B(n3143), .ZN(n3145)
         );
  NAND2_X1 U3957 ( .A1(n3661), .A2(n3156), .ZN(n3144) );
  OAI211_X1 U3958 ( .C1(n3146), .C2(n3664), .A(n3145), .B(n3144), .ZN(U3210)
         );
  AOI211_X1 U3959 ( .C1(n3149), .C2(n3148), .A(n4878), .B(n3147), .ZN(n4876)
         );
  OAI22_X1 U3960 ( .A1(n3267), .A2(n4547), .B1(n3150), .B2(n4563), .ZN(n3154)
         );
  XOR2_X1 U3961 ( .A(n3107), .B(n3151), .Z(n3152) );
  NOR2_X1 U3962 ( .A1(n3152), .A2(n4551), .ZN(n3153) );
  AOI211_X1 U3963 ( .C1(n4549), .C2(n3834), .A(n3154), .B(n3153), .ZN(n3155)
         );
  INV_X1 U3964 ( .A(n3155), .ZN(n4877) );
  AOI21_X1 U3965 ( .B1(n4876), .B2(n3878), .A(n4877), .ZN(n3161) );
  INV_X1 U3966 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3183) );
  INV_X1 U3967 ( .A(n3156), .ZN(n3157) );
  OAI22_X1 U3968 ( .A1(n4815), .A2(n3183), .B1(n3157), .B2(n4350), .ZN(n3158)
         );
  INV_X1 U3969 ( .A(n3158), .ZN(n3160) );
  NAND2_X1 U3970 ( .A1(n3105), .A2(n3107), .ZN(n4872) );
  NAND3_X1 U3971 ( .A1(n4874), .A2(n4872), .A3(n4407), .ZN(n3159) );
  OAI211_X1 U3972 ( .C1(n3161), .C2(n4806), .A(n3160), .B(n3159), .ZN(U3283)
         );
  INV_X1 U3973 ( .A(n3162), .ZN(n3165) );
  INV_X1 U3974 ( .A(n3163), .ZN(n3164) );
  NOR2_X1 U3975 ( .A1(n3165), .A2(n3164), .ZN(n3166) );
  AOI21_X1 U3976 ( .B1(n3168), .B2(n3167), .A(n3166), .ZN(n3259) );
  OAI22_X1 U3977 ( .A1(n3267), .A2(n2162), .B1(n3170), .B2(n3519), .ZN(n3169)
         );
  XNOR2_X1 U3978 ( .A(n3169), .B(n3011), .ZN(n3171) );
  OAI22_X1 U3979 ( .A1(n3267), .A2(n2984), .B1(n3170), .B2(n2162), .ZN(n3172)
         );
  NAND2_X1 U3980 ( .A1(n3171), .A2(n3172), .ZN(n3258) );
  INV_X1 U3981 ( .A(n3171), .ZN(n3174) );
  INV_X1 U3982 ( .A(n3172), .ZN(n3173) );
  NAND2_X1 U3983 ( .A1(n3174), .A2(n3173), .ZN(n3260) );
  NAND2_X1 U3984 ( .A1(n3258), .A2(n3260), .ZN(n3175) );
  XNOR2_X1 U3985 ( .A(n3259), .B(n3175), .ZN(n3180) );
  INV_X1 U3986 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4100) );
  NOR2_X1 U3987 ( .A1(STATE_REG_SCAN_IN), .A2(n4100), .ZN(n4675) );
  OAI22_X1 U3988 ( .A1(n3082), .A2(n4653), .B1(n3659), .B2(n3300), .ZN(n3176)
         );
  AOI211_X1 U3989 ( .C1(n2436), .C2(n4656), .A(n4675), .B(n3176), .ZN(n3179)
         );
  NAND2_X1 U3990 ( .A1(n3661), .A2(n3177), .ZN(n3178) );
  OAI211_X1 U3991 ( .C1(n3180), .C2(n3664), .A(n3179), .B(n3178), .ZN(U3218)
         );
  INV_X1 U3992 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3995) );
  NAND2_X1 U3993 ( .A1(n3182), .A2(n2323), .ZN(n3843) );
  XNOR2_X1 U3994 ( .A(n4642), .B(n3183), .ZN(n3842) );
  NAND2_X1 U3995 ( .A1(n3843), .A2(n3842), .ZN(n3841) );
  NAND2_X1 U3996 ( .A1(n3184), .A2(n4855), .ZN(n3185) );
  NAND2_X1 U3997 ( .A1(n3186), .A2(n3185), .ZN(n4674) );
  NOR2_X1 U3998 ( .A1(n3118), .A2(n4674), .ZN(n4673) );
  NOR2_X1 U3999 ( .A1(n3187), .A2(n4673), .ZN(n4683) );
  NAND2_X1 U4000 ( .A1(n3206), .A2(REG2_REG_9__SCAN_IN), .ZN(n3188) );
  OAI21_X1 U4001 ( .B1(n3206), .B2(REG2_REG_9__SCAN_IN), .A(n3188), .ZN(n4682)
         );
  NOR2_X1 U4002 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  INV_X1 U4003 ( .A(n3188), .ZN(n3189) );
  NOR2_X1 U4004 ( .A1(n3190), .A2(n4851), .ZN(n3191) );
  AOI22_X1 U4005 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4849), .B1(n3211), .B2(
        n3227), .ZN(n4700) );
  AND2_X1 U4006 ( .A1(n3211), .A2(REG2_REG_11__SCAN_IN), .ZN(n3192) );
  INV_X1 U4007 ( .A(n3216), .ZN(n4641) );
  NAND2_X1 U4008 ( .A1(n3193), .A2(n4641), .ZN(n3849) );
  AOI211_X1 U4009 ( .C1(n3995), .C2(n3194), .A(n3850), .B(n4754), .ZN(n3218)
         );
  INV_X1 U4010 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3195) );
  INV_X1 U4011 ( .A(n3206), .ZN(n4853) );
  AOI22_X1 U4012 ( .A1(n3206), .A2(REG1_REG_9__SCAN_IN), .B1(n3195), .B2(n4853), .ZN(n4688) );
  INV_X1 U4013 ( .A(n3197), .ZN(n3198) );
  INV_X1 U4014 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4015 ( .A1(n3204), .A2(n3203), .ZN(n3205) );
  NAND2_X1 U4016 ( .A1(n3205), .A2(n4677), .ZN(n4687) );
  NAND2_X1 U4017 ( .A1(n4688), .A2(n4687), .ZN(n4686) );
  NAND2_X1 U4018 ( .A1(n3206), .A2(REG1_REG_9__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U4019 ( .A1(n3208), .A2(n3209), .ZN(n3210) );
  NAND2_X1 U4020 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4696), .ZN(n4695) );
  NAND2_X1 U4021 ( .A1(n3210), .A2(n4695), .ZN(n4704) );
  INV_X1 U4022 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4023 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3211), .B1(n4849), .B2(
        n3951), .ZN(n4705) );
  XNOR2_X1 U4024 ( .A(n3863), .B(n3216), .ZN(n3212) );
  NAND2_X1 U4025 ( .A1(n3212), .A2(REG1_REG_12__SCAN_IN), .ZN(n3865) );
  OAI211_X1 U4026 ( .C1(n3212), .C2(REG1_REG_12__SCAN_IN), .A(n4771), .B(n3865), .ZN(n3215) );
  NAND2_X1 U4027 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n3549) );
  INV_X1 U4028 ( .A(n3549), .ZN(n3213) );
  AOI21_X1 U4029 ( .B1(n4767), .B2(ADDR_REG_12__SCAN_IN), .A(n3213), .ZN(n3214) );
  OAI211_X1 U4030 ( .C1(n4775), .C2(n3216), .A(n3215), .B(n3214), .ZN(n3217)
         );
  OR2_X1 U4031 ( .A1(n3218), .A2(n3217), .ZN(U3252) );
  NAND2_X1 U4032 ( .A1(n4815), .A2(n4789), .ZN(n4421) );
  INV_X1 U4033 ( .A(n3221), .ZN(n3730) );
  XNOR2_X1 U4034 ( .A(n3219), .B(n3730), .ZN(n3323) );
  NAND2_X1 U4035 ( .A1(n3220), .A2(n3221), .ZN(n3222) );
  NAND2_X1 U4036 ( .A1(n3223), .A2(n3222), .ZN(n3317) );
  NAND2_X1 U4037 ( .A1(n3224), .A2(n3619), .ZN(n3225) );
  NAND2_X1 U4038 ( .A1(n3310), .A2(n3225), .ZN(n3329) );
  INV_X1 U4039 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3227) );
  INV_X1 U4040 ( .A(n3620), .ZN(n3226) );
  OAI22_X1 U4041 ( .A1(n4815), .A2(n3227), .B1(n3226), .B2(n4350), .ZN(n3228)
         );
  AOI21_X1 U4042 ( .B1(n3619), .B2(n3361), .A(n3228), .ZN(n3231) );
  AOI22_X1 U40430 ( .A1(n4412), .A2(n3830), .B1(n4411), .B2(n3229), .ZN(n3230)
         );
  OAI211_X1 U4044 ( .C1(n3329), .C2(n4441), .A(n3231), .B(n3230), .ZN(n3232)
         );
  AOI21_X1 U4045 ( .B1(n3317), .B2(n4407), .A(n3232), .ZN(n3233) );
  OAI21_X1 U4046 ( .B1(n4421), .B2(n3323), .A(n3233), .ZN(U3279) );
  NAND2_X1 U4047 ( .A1(n3234), .A2(n4873), .ZN(n3239) );
  NOR2_X1 U4048 ( .A1(n3262), .A2(n4563), .ZN(n3235) );
  AOI21_X1 U4049 ( .B1(n3830), .B2(n4792), .A(n3235), .ZN(n3238) );
  NAND2_X1 U4050 ( .A1(n3832), .A2(n4549), .ZN(n3236) );
  NAND4_X1 U4051 ( .A1(n3239), .A2(n3238), .A3(n3237), .A4(n3236), .ZN(n3242)
         );
  MUX2_X1 U4052 ( .A(REG0_REG_9__SCAN_IN), .B(n3242), .S(n4886), .Z(n3240) );
  AOI21_X1 U4053 ( .B1(n3244), .B2(n4865), .A(n3240), .ZN(n3241) );
  INV_X1 U4054 ( .A(n3241), .ZN(U3485) );
  MUX2_X1 U4055 ( .A(REG1_REG_9__SCAN_IN), .B(n3242), .S(n4898), .Z(n3243) );
  AOI21_X1 U4056 ( .B1(n4888), .B2(n3244), .A(n3243), .ZN(n3245) );
  INV_X1 U4057 ( .A(n3245), .ZN(U3527) );
  NAND2_X1 U4058 ( .A1(n3774), .A2(n3780), .ZN(n3728) );
  XNOR2_X1 U4059 ( .A(n3246), .B(n3728), .ZN(n3277) );
  OR2_X1 U4060 ( .A1(n3247), .A2(n3291), .ZN(n3248) );
  NAND2_X1 U4061 ( .A1(n3224), .A2(n3248), .ZN(n3282) );
  INV_X1 U4062 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3250) );
  INV_X1 U4063 ( .A(n3249), .ZN(n3305) );
  OAI22_X1 U4064 ( .A1(n4815), .A2(n3250), .B1(n3305), .B2(n4350), .ZN(n3251)
         );
  AOI21_X1 U4065 ( .B1(n3302), .B2(n3361), .A(n3251), .ZN(n3253) );
  AOI22_X1 U4066 ( .A1(n4412), .A2(n3831), .B1(n4411), .B2(n3829), .ZN(n3252)
         );
  OAI211_X1 U4067 ( .C1(n3282), .C2(n4441), .A(n3253), .B(n3252), .ZN(n3256)
         );
  XNOR2_X1 U4068 ( .A(n3254), .B(n3728), .ZN(n3275) );
  NOR2_X1 U4069 ( .A1(n3275), .A2(n4421), .ZN(n3255) );
  AOI211_X1 U4070 ( .C1(n4407), .C2(n3277), .A(n3256), .B(n3255), .ZN(n3257)
         );
  INV_X1 U4071 ( .A(n3257), .ZN(U3280) );
  NAND2_X1 U4072 ( .A1(n3259), .A2(n3258), .ZN(n3261) );
  NAND2_X1 U4073 ( .A1(n3261), .A2(n3260), .ZN(n3284) );
  OAI22_X1 U4074 ( .A1(n3300), .A2(n2984), .B1(n3262), .B2(n2162), .ZN(n3286)
         );
  NAND2_X1 U4075 ( .A1(n3831), .A2(n2176), .ZN(n3264) );
  NAND2_X1 U4076 ( .A1(n3269), .A2(n3477), .ZN(n3263) );
  NAND2_X1 U4077 ( .A1(n3264), .A2(n3263), .ZN(n3265) );
  XNOR2_X1 U4078 ( .A(n3265), .B(n3011), .ZN(n3285) );
  XOR2_X1 U4079 ( .A(n3286), .B(n3285), .Z(n3283) );
  XNOR2_X1 U4080 ( .A(n3284), .B(n3283), .ZN(n3266) );
  NAND2_X1 U4081 ( .A1(n3266), .A2(n4663), .ZN(n3271) );
  NOR2_X1 U4082 ( .A1(STATE_REG_SCAN_IN), .A2(n2448), .ZN(n4684) );
  OAI22_X1 U4083 ( .A1(n3267), .A2(n4653), .B1(n3659), .B2(n3617), .ZN(n3268)
         );
  AOI211_X1 U4084 ( .C1(n3269), .C2(n4656), .A(n4684), .B(n3268), .ZN(n3270)
         );
  OAI211_X1 U4085 ( .C1(n4668), .C2(n3272), .A(n3271), .B(n3270), .ZN(U3228)
         );
  OAI22_X1 U4086 ( .A1(n4568), .A2(n4547), .B1(n4563), .B2(n3291), .ZN(n3273)
         );
  AOI21_X1 U4087 ( .B1(n4549), .B2(n3831), .A(n3273), .ZN(n3274) );
  OAI21_X1 U4088 ( .B1(n3275), .B2(n4551), .A(n3274), .ZN(n3276) );
  AOI21_X1 U4089 ( .B1(n4873), .B2(n3277), .A(n3276), .ZN(n3279) );
  MUX2_X1 U4090 ( .A(n2466), .B(n3279), .S(n4886), .Z(n3278) );
  OAI21_X1 U4091 ( .B1(n3282), .B2(n4632), .A(n3278), .ZN(U3487) );
  INV_X1 U4092 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3280) );
  MUX2_X1 U4093 ( .A(n3280), .B(n3279), .S(n4898), .Z(n3281) );
  OAI21_X1 U4094 ( .B1(n3282), .B2(n4561), .A(n3281), .ZN(U3528) );
  NAND2_X1 U4095 ( .A1(n3284), .A2(n3283), .ZN(n3290) );
  INV_X1 U4096 ( .A(n3285), .ZN(n3288) );
  INV_X1 U4097 ( .A(n3286), .ZN(n3287) );
  NAND2_X1 U4098 ( .A1(n3288), .A2(n3287), .ZN(n3289) );
  NOR2_X1 U4099 ( .A1(n3291), .A2(n2162), .ZN(n3292) );
  AOI21_X1 U4100 ( .B1(n3830), .B2(n3483), .A(n3292), .ZN(n3330) );
  NAND2_X1 U4101 ( .A1(n3830), .A2(n2176), .ZN(n3294) );
  NAND2_X1 U4102 ( .A1(n3302), .A2(n3477), .ZN(n3293) );
  NAND2_X1 U4103 ( .A1(n3294), .A2(n3293), .ZN(n3295) );
  XNOR2_X1 U4104 ( .A(n3295), .B(n3011), .ZN(n3332) );
  XOR2_X1 U4105 ( .A(n3330), .B(n3332), .Z(n3297) );
  AOI21_X1 U4106 ( .B1(n3296), .B2(n3297), .A(n3664), .ZN(n3299) );
  NAND2_X1 U4107 ( .A1(n3299), .A2(n3334), .ZN(n3304) );
  NOR2_X1 U4108 ( .A1(STATE_REG_SCAN_IN), .A2(n4040), .ZN(n4693) );
  OAI22_X1 U4109 ( .A1(n3300), .A2(n4653), .B1(n3659), .B2(n4568), .ZN(n3301)
         );
  AOI211_X1 U4110 ( .C1(n3302), .C2(n4656), .A(n4693), .B(n3301), .ZN(n3303)
         );
  OAI211_X1 U4111 ( .C1(n4668), .C2(n3305), .A(n3304), .B(n3303), .ZN(U3214)
         );
  INV_X1 U4112 ( .A(n4423), .ZN(n3306) );
  NOR2_X1 U4113 ( .A1(n4424), .A2(n3306), .ZN(n3710) );
  XNOR2_X1 U4114 ( .A(n4425), .B(n3710), .ZN(n3307) );
  NAND2_X1 U4115 ( .A1(n3307), .A2(n4789), .ZN(n4571) );
  INV_X1 U4116 ( .A(n3710), .ZN(n3309) );
  XNOR2_X1 U4117 ( .A(n3308), .B(n3309), .ZN(n4562) );
  NAND2_X1 U4118 ( .A1(n4562), .A2(n4407), .ZN(n3316) );
  AOI21_X1 U4119 ( .B1(n3311), .B2(n3310), .A(n2194), .ZN(n4636) );
  AOI22_X1 U4120 ( .A1(n4412), .A2(n3829), .B1(n4411), .B2(n4566), .ZN(n3313)
         );
  AOI22_X1 U4121 ( .A1(n4806), .A2(REG2_REG_12__SCAN_IN), .B1(n3552), .B2(
        n4810), .ZN(n3312) );
  OAI211_X1 U4122 ( .C1(n4564), .C2(n4416), .A(n3313), .B(n3312), .ZN(n3314)
         );
  AOI21_X1 U4123 ( .B1(n4636), .B2(n4802), .A(n3314), .ZN(n3315) );
  OAI211_X1 U4124 ( .C1(n4806), .C2(n4571), .A(n3316), .B(n3315), .ZN(U3278)
         );
  NAND2_X1 U4125 ( .A1(n3317), .A2(n4873), .ZN(n3322) );
  NAND2_X1 U4126 ( .A1(n3619), .A2(n4791), .ZN(n3319) );
  NAND2_X1 U4127 ( .A1(n3830), .A2(n4549), .ZN(n3318) );
  OAI211_X1 U4128 ( .C1(n4431), .C2(n4547), .A(n3319), .B(n3318), .ZN(n3320)
         );
  INV_X1 U4129 ( .A(n3320), .ZN(n3321) );
  OAI211_X1 U4130 ( .C1(n3323), .C2(n4551), .A(n3322), .B(n3321), .ZN(n3326)
         );
  MUX2_X1 U4131 ( .A(n3326), .B(REG1_REG_11__SCAN_IN), .S(n4895), .Z(n3324) );
  INV_X1 U4132 ( .A(n3324), .ZN(n3325) );
  OAI21_X1 U4133 ( .B1(n4561), .B2(n3329), .A(n3325), .ZN(U3529) );
  MUX2_X1 U4134 ( .A(n3326), .B(REG0_REG_11__SCAN_IN), .S(n4885), .Z(n3327) );
  INV_X1 U4135 ( .A(n3327), .ZN(n3328) );
  OAI21_X1 U4136 ( .B1(n3329), .B2(n4632), .A(n3328), .ZN(U3489) );
  INV_X1 U4137 ( .A(n3330), .ZN(n3331) );
  NAND2_X1 U4138 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  OAI22_X1 U4139 ( .A1(n4568), .A2(n2984), .B1(n2162), .B2(n3335), .ZN(n3613)
         );
  OAI22_X1 U4140 ( .A1(n4568), .A2(n2162), .B1(n3519), .B2(n3335), .ZN(n3336)
         );
  XNOR2_X1 U4141 ( .A(n3336), .B(n3011), .ZN(n3614) );
  OAI22_X1 U4142 ( .A1(n4431), .A2(n2162), .B1(n3519), .B2(n4564), .ZN(n3337)
         );
  XNOR2_X1 U4143 ( .A(n3337), .B(n3011), .ZN(n3340) );
  OAI22_X1 U4144 ( .A1(n4431), .A2(n2984), .B1(n2162), .B2(n4564), .ZN(n3339)
         );
  AND2_X1 U4145 ( .A1(n3340), .A2(n3339), .ZN(n3545) );
  AOI21_X1 U4146 ( .B1(n3613), .B2(n3614), .A(n3545), .ZN(n3338) );
  NAND2_X1 U4147 ( .A1(n3541), .A2(n3338), .ZN(n3344) );
  NOR2_X1 U4148 ( .A1(n3614), .A2(n3613), .ZN(n3342) );
  INV_X1 U4149 ( .A(n3545), .ZN(n3341) );
  NOR2_X1 U4150 ( .A1(n3340), .A2(n3339), .ZN(n3546) );
  AOI21_X1 U4151 ( .B1(n3342), .B2(n3341), .A(n3546), .ZN(n3343) );
  AOI22_X1 U4152 ( .A1(n4566), .A2(n2176), .B1(n3477), .B2(n4428), .ZN(n3345)
         );
  XNOR2_X1 U4153 ( .A(n3345), .B(n3011), .ZN(n3596) );
  AOI22_X1 U4154 ( .A1(n4566), .A2(n3483), .B1(n2176), .B2(n4428), .ZN(n3597)
         );
  OAI22_X1 U4155 ( .A1(n4542), .A2(n2162), .B1(n3519), .B2(n4546), .ZN(n3346)
         );
  XNOR2_X1 U4156 ( .A(n3346), .B(n3011), .ZN(n3348) );
  OAI22_X1 U4157 ( .A1(n4542), .A2(n2984), .B1(n2162), .B2(n4546), .ZN(n3347)
         );
  OR2_X1 U4158 ( .A1(n3348), .A2(n3347), .ZN(n3368) );
  INV_X1 U4159 ( .A(n3368), .ZN(n3349) );
  AND2_X1 U4160 ( .A1(n3348), .A2(n3347), .ZN(n3369) );
  NOR2_X1 U4161 ( .A1(n3349), .A2(n3369), .ZN(n3350) );
  XNOR2_X1 U4162 ( .A(n3370), .B(n3350), .ZN(n3354) );
  INV_X1 U4163 ( .A(n4653), .ZN(n3630) );
  AOI22_X1 U4164 ( .A1(n3630), .A2(n4566), .B1(n3631), .B2(n4410), .ZN(n3351)
         );
  NAND2_X1 U4165 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4723) );
  OAI211_X1 U4166 ( .C1(n3652), .C2(n4546), .A(n3351), .B(n4723), .ZN(n3352)
         );
  AOI21_X1 U4167 ( .B1(n4413), .B2(n3661), .A(n3352), .ZN(n3353) );
  OAI21_X1 U4168 ( .B1(n3354), .B2(n3664), .A(n3353), .ZN(U3212) );
  MUX2_X1 U4169 ( .A(n3355), .B(REG2_REG_2__SCAN_IN), .S(n4806), .Z(n3367) );
  INV_X1 U4170 ( .A(n4411), .ZN(n3357) );
  OAI22_X1 U4171 ( .A1(n3358), .A2(n3357), .B1(n4441), .B2(n3356), .ZN(n3359)
         );
  AOI21_X1 U4172 ( .B1(n3360), .B2(n4811), .A(n3359), .ZN(n3363) );
  AOI22_X1 U4173 ( .A1(n3361), .A2(n3629), .B1(REG3_REG_2__SCAN_IN), .B2(n4810), .ZN(n3362) );
  OAI211_X1 U4174 ( .C1(n3365), .C2(n3364), .A(n3363), .B(n3362), .ZN(n3366)
         );
  OR2_X1 U4175 ( .A1(n3367), .A2(n3366), .ZN(U3288) );
  OAI22_X1 U4176 ( .A1(n4652), .A2(n2162), .B1(n3519), .B2(n4399), .ZN(n3371)
         );
  XOR2_X1 U4177 ( .A(n3011), .B(n3371), .Z(n3374) );
  NAND2_X1 U4178 ( .A1(n3375), .A2(n3374), .ZN(n3657) );
  NAND2_X1 U4179 ( .A1(n4410), .A2(n3483), .ZN(n3373) );
  NAND2_X1 U4180 ( .A1(n4538), .A2(n2176), .ZN(n3372) );
  NAND2_X1 U4181 ( .A1(n3373), .A2(n3372), .ZN(n4659) );
  NAND2_X1 U4182 ( .A1(n3657), .A2(n4659), .ZN(n3379) );
  OAI22_X1 U4183 ( .A1(n4525), .A2(n2162), .B1(n3519), .B2(n4381), .ZN(n3376)
         );
  XNOR2_X1 U4184 ( .A(n3376), .B(n3011), .ZN(n3378) );
  OAI22_X1 U4185 ( .A1(n4525), .A2(n2984), .B1(n2162), .B2(n4381), .ZN(n3377)
         );
  NOR2_X1 U4186 ( .A1(n3378), .A2(n3377), .ZN(n3380) );
  AOI21_X1 U4187 ( .B1(n3378), .B2(n3377), .A(n3380), .ZN(n4661) );
  NAND3_X1 U4188 ( .A1(n3379), .A2(n4658), .A3(n4661), .ZN(n3442) );
  INV_X1 U4189 ( .A(n3380), .ZN(n3501) );
  OAI22_X1 U4190 ( .A1(n4326), .A2(n2162), .B1(n4312), .B2(n3519), .ZN(n3381)
         );
  XNOR2_X1 U4191 ( .A(n3381), .B(n3011), .ZN(n3385) );
  INV_X1 U4192 ( .A(n3385), .ZN(n3383) );
  OAI22_X1 U4193 ( .A1(n4326), .A2(n2984), .B1(n4312), .B2(n2162), .ZN(n3384)
         );
  INV_X1 U4194 ( .A(n3384), .ZN(n3382) );
  NAND2_X1 U4195 ( .A1(n3383), .A2(n3382), .ZN(n3589) );
  NAND2_X1 U4196 ( .A1(n3385), .A2(n3384), .ZN(n3587) );
  INV_X1 U4197 ( .A(n3587), .ZN(n3397) );
  OAI22_X1 U4198 ( .A1(n4304), .A2(n2162), .B1(n3519), .B2(n4333), .ZN(n3386)
         );
  XNOR2_X1 U4199 ( .A(n3386), .B(n3011), .ZN(n3390) );
  INV_X1 U4200 ( .A(n3390), .ZN(n3388) );
  OAI22_X1 U4201 ( .A1(n4304), .A2(n2984), .B1(n2162), .B2(n4333), .ZN(n3391)
         );
  INV_X1 U4202 ( .A(n3391), .ZN(n3387) );
  NAND2_X1 U4203 ( .A1(n3388), .A2(n3387), .ZN(n3396) );
  OAI22_X1 U4204 ( .A1(n4325), .A2(n2162), .B1(n3519), .B2(n2556), .ZN(n3389)
         );
  XNOR2_X1 U4205 ( .A(n3389), .B(n3011), .ZN(n3394) );
  OAI22_X1 U4206 ( .A1(n4325), .A2(n2984), .B1(n2162), .B2(n2556), .ZN(n3393)
         );
  NAND2_X1 U4207 ( .A1(n3394), .A2(n3393), .ZN(n3637) );
  XOR2_X1 U4208 ( .A(n3391), .B(n3390), .Z(n3508) );
  AND2_X1 U4209 ( .A1(n3637), .A2(n3508), .ZN(n3401) );
  INV_X1 U4210 ( .A(n3401), .ZN(n3395) );
  OAI22_X1 U4211 ( .A1(n4654), .A2(n2162), .B1(n4369), .B2(n3519), .ZN(n3392)
         );
  XNOR2_X1 U4212 ( .A(n3392), .B(n3011), .ZN(n3400) );
  OAI22_X1 U4213 ( .A1(n4654), .A2(n2984), .B1(n4369), .B2(n2162), .ZN(n3399)
         );
  OR2_X1 U4214 ( .A1(n3400), .A2(n3399), .ZN(n3635) );
  OR2_X1 U4215 ( .A1(n3394), .A2(n3393), .ZN(n3638) );
  AND2_X1 U4216 ( .A1(n3635), .A2(n3638), .ZN(n3502) );
  OR2_X1 U4217 ( .A1(n3395), .A2(n3502), .ZN(n3505) );
  AND2_X1 U4218 ( .A1(n3396), .A2(n3505), .ZN(n3584) );
  OR2_X1 U4219 ( .A1(n3397), .A2(n3584), .ZN(n3582) );
  AND2_X1 U4220 ( .A1(n3589), .A2(n3582), .ZN(n3398) );
  AND2_X1 U4221 ( .A1(n3501), .A2(n3398), .ZN(n3435) );
  NAND2_X1 U4222 ( .A1(n3442), .A2(n3435), .ZN(n3403) );
  INV_X1 U4223 ( .A(n3398), .ZN(n3402) );
  NAND2_X1 U4224 ( .A1(n3400), .A2(n3399), .ZN(n3565) );
  AND2_X1 U4225 ( .A1(n3565), .A2(n3401), .ZN(n3504) );
  AND2_X1 U4226 ( .A1(n3504), .A2(n3587), .ZN(n3580) );
  OR2_X1 U4227 ( .A1(n3402), .A2(n3580), .ZN(n3449) );
  AND2_X1 U4228 ( .A1(n3403), .A2(n3449), .ZN(n3406) );
  OAI22_X1 U4229 ( .A1(n4305), .A2(n2162), .B1(n3519), .B2(n4501), .ZN(n3404)
         );
  XNOR2_X1 U4230 ( .A(n3404), .B(n3011), .ZN(n3445) );
  OAI22_X1 U4231 ( .A1(n4305), .A2(n2984), .B1(n2162), .B2(n4501), .ZN(n3444)
         );
  XNOR2_X1 U4232 ( .A(n3445), .B(n3444), .ZN(n3405) );
  XNOR2_X1 U4233 ( .A(n3406), .B(n3405), .ZN(n3411) );
  OAI22_X1 U4234 ( .A1(n4326), .A2(n4653), .B1(n3659), .B2(n4502), .ZN(n3409)
         );
  OAI22_X1 U4235 ( .A1(n3652), .A2(n4501), .B1(STATE_REG_SCAN_IN), .B2(n3407), 
        .ZN(n3408) );
  AOI211_X1 U4236 ( .C1(n4292), .C2(n3661), .A(n3409), .B(n3408), .ZN(n3410)
         );
  OAI21_X1 U4237 ( .B1(n3411), .B2(n3664), .A(n3410), .ZN(U3220) );
  INV_X1 U4238 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n3413) );
  NAND2_X1 U4239 ( .A1(n2858), .A2(U4043), .ZN(n3412) );
  OAI21_X1 U4240 ( .B1(U4043), .B2(n3413), .A(n3412), .ZN(U3550) );
  INV_X1 U4241 ( .A(n3415), .ZN(n3421) );
  AOI22_X1 U4242 ( .A1(n4412), .A2(n4466), .B1(n4411), .B2(n3828), .ZN(n3417)
         );
  AOI22_X1 U4243 ( .A1(n4806), .A2(REG2_REG_28__SCAN_IN), .B1(n3530), .B2(
        n4810), .ZN(n3416) );
  OAI211_X1 U4244 ( .C1(n3527), .C2(n4416), .A(n3417), .B(n3416), .ZN(n3420)
         );
  NOR2_X1 U4245 ( .A1(n3418), .A2(n4806), .ZN(n3419) );
  AOI211_X1 U4246 ( .C1(n4802), .C2(n3421), .A(n3420), .B(n3419), .ZN(n3422)
         );
  OAI21_X1 U4247 ( .B1(n3423), .B2(n4388), .A(n3422), .ZN(U3262) );
  INV_X1 U4248 ( .A(n3424), .ZN(n3427) );
  NAND3_X1 U4249 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n2342), 
        .ZN(n3426) );
  INV_X1 U4250 ( .A(DATAI_31_), .ZN(n3425) );
  OAI22_X1 U4251 ( .A1(n3427), .A2(n3426), .B1(STATE_REG_SCAN_IN), .B2(n3425), 
        .ZN(U3321) );
  INV_X1 U4252 ( .A(n3428), .ZN(n3429) );
  INV_X1 U4253 ( .A(D_REG_0__SCAN_IN), .ZN(n3973) );
  NOR2_X1 U4254 ( .A1(n3431), .A2(n4639), .ZN(n3433) );
  AOI22_X1 U4255 ( .A1(n4835), .A2(n3973), .B1(n3433), .B2(n3432), .ZN(U3458)
         );
  INV_X1 U4256 ( .A(D_REG_1__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U4257 ( .A1(n4835), .A2(n4101), .B1(n2705), .B2(n3433), .ZN(U3459)
         );
  NOR2_X1 U4258 ( .A1(n3445), .A2(n3444), .ZN(n3450) );
  INV_X1 U4259 ( .A(n3450), .ZN(n3434) );
  AND2_X1 U4260 ( .A1(n3435), .A2(n3434), .ZN(n3488) );
  OAI22_X1 U4261 ( .A1(n4502), .A2(n2162), .B1(n3519), .B2(n4283), .ZN(n3436)
         );
  XNOR2_X1 U4262 ( .A(n3436), .B(n3011), .ZN(n3447) );
  OAI22_X1 U4263 ( .A1(n4502), .A2(n2984), .B1(n2162), .B2(n4283), .ZN(n3446)
         );
  NOR2_X1 U4264 ( .A1(n3447), .A2(n3446), .ZN(n3494) );
  NAND2_X1 U4265 ( .A1(n4483), .A2(n2176), .ZN(n3438) );
  NAND2_X1 U4266 ( .A1(n4489), .A2(n3477), .ZN(n3437) );
  NAND2_X1 U4267 ( .A1(n3438), .A2(n3437), .ZN(n3439) );
  XNOR2_X1 U4268 ( .A(n3439), .B(n3480), .ZN(n3457) );
  NOR2_X1 U4269 ( .A1(n2162), .A2(n4268), .ZN(n3440) );
  AOI21_X1 U4270 ( .B1(n4483), .B2(n3483), .A(n3440), .ZN(n3456) );
  XNOR2_X1 U4271 ( .A(n3457), .B(n3456), .ZN(n3493) );
  NOR2_X1 U4272 ( .A1(n3494), .A2(n3493), .ZN(n3443) );
  AND2_X1 U4273 ( .A1(n3488), .A2(n3443), .ZN(n3441) );
  NAND2_X1 U4274 ( .A1(n3442), .A2(n3441), .ZN(n3455) );
  INV_X1 U4275 ( .A(n3443), .ZN(n3453) );
  NAND2_X1 U4276 ( .A1(n3445), .A2(n3444), .ZN(n3491) );
  XNOR2_X1 U4277 ( .A(n3447), .B(n3446), .ZN(n3607) );
  INV_X1 U4278 ( .A(n3607), .ZN(n3448) );
  AND2_X1 U4279 ( .A1(n3491), .A2(n3448), .ZN(n3451) );
  OR2_X1 U4280 ( .A1(n3450), .A2(n3449), .ZN(n3489) );
  AND2_X1 U4281 ( .A1(n3451), .A2(n3489), .ZN(n3452) );
  OR2_X1 U4282 ( .A1(n3453), .A2(n3452), .ZN(n3454) );
  NOR2_X1 U4283 ( .A1(n3457), .A2(n3456), .ZN(n3460) );
  OAI22_X1 U4284 ( .A1(n4476), .A2(n2984), .B1(n2162), .B2(n4480), .ZN(n3462)
         );
  NAND2_X1 U4285 ( .A1(n2319), .A2(n3458), .ZN(n3571) );
  OAI22_X1 U4286 ( .A1(n4476), .A2(n2162), .B1(n3519), .B2(n4480), .ZN(n3459)
         );
  XNOR2_X1 U4287 ( .A(n3459), .B(n3011), .ZN(n3574) );
  NAND2_X1 U4288 ( .A1(n3571), .A2(n3574), .ZN(n3464) );
  INV_X1 U4289 ( .A(n3460), .ZN(n3461) );
  NAND2_X1 U4290 ( .A1(n2319), .A2(n3461), .ZN(n3463) );
  NAND2_X1 U4291 ( .A1(n3463), .A2(n3462), .ZN(n3572) );
  NAND2_X1 U4292 ( .A1(n3464), .A2(n3572), .ZN(n3557) );
  OAI22_X1 U4293 ( .A1(n4481), .A2(n2162), .B1(n4223), .B2(n3519), .ZN(n3465)
         );
  XNOR2_X1 U4294 ( .A(n3465), .B(n3011), .ZN(n3467) );
  OAI22_X1 U4295 ( .A1(n4481), .A2(n2984), .B1(n4223), .B2(n2162), .ZN(n3466)
         );
  OR2_X1 U4296 ( .A1(n3467), .A2(n3466), .ZN(n3556) );
  NAND2_X1 U4297 ( .A1(n3467), .A2(n3466), .ZN(n3555) );
  NAND2_X1 U4298 ( .A1(n4473), .A2(n2176), .ZN(n3470) );
  NAND2_X1 U4299 ( .A1(n3468), .A2(n3477), .ZN(n3469) );
  NAND2_X1 U4300 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  XNOR2_X1 U4301 ( .A(n3471), .B(n3480), .ZN(n3475) );
  NOR2_X1 U4302 ( .A1(n2162), .A2(n4464), .ZN(n3472) );
  AOI21_X1 U4303 ( .B1(n4473), .B2(n3483), .A(n3472), .ZN(n3474) );
  NOR2_X1 U4304 ( .A1(n3475), .A2(n3474), .ZN(n3649) );
  INV_X1 U4305 ( .A(n3649), .ZN(n3473) );
  NAND2_X1 U4306 ( .A1(n3475), .A2(n3474), .ZN(n3647) );
  NAND2_X1 U4307 ( .A1(n3476), .A2(n3647), .ZN(n3518) );
  NAND2_X1 U4308 ( .A1(n4466), .A2(n2176), .ZN(n3479) );
  NAND2_X1 U4309 ( .A1(n3897), .A2(n3477), .ZN(n3478) );
  NAND2_X1 U4310 ( .A1(n3479), .A2(n3478), .ZN(n3481) );
  XNOR2_X1 U4311 ( .A(n3481), .B(n3480), .ZN(n3515) );
  NOR2_X1 U4312 ( .A1(n2162), .A2(n4456), .ZN(n3482) );
  AOI21_X1 U4313 ( .B1(n4466), .B2(n3483), .A(n3482), .ZN(n3514) );
  XNOR2_X1 U4314 ( .A(n3515), .B(n3514), .ZN(n3517) );
  XNOR2_X1 U4315 ( .A(n3518), .B(n3517), .ZN(n3487) );
  INV_X1 U4316 ( .A(n4473), .ZN(n3559) );
  OAI22_X1 U4317 ( .A1(n3521), .A2(n3659), .B1(n4653), .B2(n3559), .ZN(n3485)
         );
  OAI22_X1 U4318 ( .A1(n3652), .A2(n4456), .B1(STATE_REG_SCAN_IN), .B2(n4098), 
        .ZN(n3484) );
  AOI211_X1 U4319 ( .C1(n3900), .C2(n3661), .A(n3485), .B(n3484), .ZN(n3486)
         );
  OAI21_X1 U4320 ( .B1(n3487), .B2(n3664), .A(n3486), .ZN(U3211) );
  NAND2_X1 U4321 ( .A1(n3442), .A2(n3488), .ZN(n3490) );
  AND2_X1 U4322 ( .A1(n3490), .A2(n3489), .ZN(n3492) );
  NAND2_X1 U4323 ( .A1(n3492), .A2(n3491), .ZN(n3606) );
  NOR2_X1 U4324 ( .A1(n3606), .A2(n3607), .ZN(n3605) );
  OAI21_X1 U4325 ( .B1(n3605), .B2(n3494), .A(n3493), .ZN(n3495) );
  NAND3_X1 U4326 ( .A1(n2319), .A2(n3495), .A3(n4663), .ZN(n3499) );
  OAI22_X1 U4327 ( .A1(n4502), .A2(n4653), .B1(n3659), .B2(n4476), .ZN(n3497)
         );
  INV_X1 U4328 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4052) );
  OAI22_X1 U4329 ( .A1(n3652), .A2(n4268), .B1(STATE_REG_SCAN_IN), .B2(n4052), 
        .ZN(n3496) );
  AOI211_X1 U4330 ( .C1(n4265), .C2(n3661), .A(n3497), .B(n3496), .ZN(n3498)
         );
  NAND2_X1 U4331 ( .A1(n3499), .A2(n3498), .ZN(U3213) );
  INV_X1 U4332 ( .A(n3500), .ZN(n4335) );
  NAND2_X1 U4333 ( .A1(n3442), .A2(n3501), .ZN(n3581) );
  NAND2_X1 U4334 ( .A1(n3581), .A2(n3565), .ZN(n3636) );
  NAND2_X1 U4335 ( .A1(n3636), .A2(n3502), .ZN(n3503) );
  AND2_X1 U4336 ( .A1(n3503), .A2(n3637), .ZN(n3507) );
  NAND2_X1 U4337 ( .A1(n3581), .A2(n3504), .ZN(n3585) );
  AND2_X1 U4338 ( .A1(n3585), .A2(n3505), .ZN(n3506) );
  OAI21_X1 U4339 ( .B1(n3508), .B2(n3507), .A(n3506), .ZN(n3509) );
  NAND2_X1 U4340 ( .A1(n3509), .A2(n4663), .ZN(n3513) );
  NAND2_X1 U4341 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3877) );
  INV_X1 U4342 ( .A(n3877), .ZN(n3511) );
  OAI22_X1 U4343 ( .A1(n4325), .A2(n4653), .B1(n3659), .B2(n4326), .ZN(n3510)
         );
  AOI211_X1 U4344 ( .C1(n3719), .C2(n4656), .A(n3511), .B(n3510), .ZN(n3512)
         );
  OAI211_X1 U4345 ( .C1(n4668), .C2(n4335), .A(n3513), .B(n3512), .ZN(U3216)
         );
  OAI22_X1 U4346 ( .A1(n3521), .A2(n2162), .B1(n3519), .B2(n3527), .ZN(n3520)
         );
  XNOR2_X1 U4347 ( .A(n3520), .B(n3011), .ZN(n3523) );
  OAI22_X1 U4348 ( .A1(n3521), .A2(n2984), .B1(n2162), .B2(n3527), .ZN(n3522)
         );
  XNOR2_X1 U4349 ( .A(n3523), .B(n3522), .ZN(n3524) );
  OAI22_X1 U4350 ( .A1(n3803), .A2(n4653), .B1(n3659), .B2(n3525), .ZN(n3529)
         );
  OAI22_X1 U4351 ( .A1(n3652), .A2(n3527), .B1(STATE_REG_SCAN_IN), .B2(n3526), 
        .ZN(n3528) );
  AOI211_X1 U4352 ( .C1(n3530), .C2(n3661), .A(n3529), .B(n3528), .ZN(n3531)
         );
  AOI211_X1 U4353 ( .C1(n3534), .C2(n3533), .A(n3664), .B(n3532), .ZN(n3535)
         );
  INV_X1 U4354 ( .A(n3535), .ZN(n3540) );
  AOI22_X1 U4355 ( .A1(n4656), .A2(n3536), .B1(REG3_REG_1__SCAN_IN), .B2(n3628), .ZN(n3539) );
  AOI22_X1 U4356 ( .A1(n3630), .A2(n2858), .B1(n3631), .B2(n3537), .ZN(n3538)
         );
  NAND3_X1 U4357 ( .A1(n3540), .A2(n3539), .A3(n3538), .ZN(U3219) );
  INV_X1 U4358 ( .A(n3613), .ZN(n3544) );
  INV_X1 U4359 ( .A(n3541), .ZN(n3542) );
  OAI21_X1 U4360 ( .B1(n3542), .B2(n3613), .A(n3614), .ZN(n3543) );
  OAI21_X1 U4361 ( .B1(n3541), .B2(n3544), .A(n3543), .ZN(n3548) );
  NOR2_X1 U4362 ( .A1(n3546), .A2(n3545), .ZN(n3547) );
  XNOR2_X1 U4363 ( .A(n3548), .B(n3547), .ZN(n3554) );
  AOI22_X1 U4364 ( .A1(n3630), .A2(n3829), .B1(n3631), .B2(n4566), .ZN(n3550)
         );
  OAI211_X1 U4365 ( .C1(n3652), .C2(n4564), .A(n3550), .B(n3549), .ZN(n3551)
         );
  AOI21_X1 U4366 ( .B1(n3552), .B2(n3661), .A(n3551), .ZN(n3553) );
  OAI21_X1 U4367 ( .B1(n3554), .B2(n3664), .A(n3553), .ZN(U3221) );
  NAND2_X1 U4368 ( .A1(n3556), .A2(n3555), .ZN(n3558) );
  XOR2_X1 U4369 ( .A(n3558), .B(n3557), .Z(n3564) );
  OAI22_X1 U4370 ( .A1(n4476), .A2(n4653), .B1(n3659), .B2(n3559), .ZN(n3562)
         );
  OAI22_X1 U4371 ( .A1(n3652), .A2(n4223), .B1(STATE_REG_SCAN_IN), .B2(n3560), 
        .ZN(n3561) );
  AOI211_X1 U4372 ( .C1(n4220), .C2(n3661), .A(n3562), .B(n3561), .ZN(n3563)
         );
  OAI21_X1 U4373 ( .B1(n3564), .B2(n3664), .A(n3563), .ZN(U3222) );
  NAND2_X1 U4374 ( .A1(n3635), .A2(n3565), .ZN(n3566) );
  XNOR2_X1 U4375 ( .A(n3581), .B(n3566), .ZN(n3570) );
  AND2_X1 U4376 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4759) );
  OAI22_X1 U4377 ( .A1(n4525), .A2(n4653), .B1(n3659), .B2(n4325), .ZN(n3567)
         );
  AOI211_X1 U4378 ( .C1(n4521), .C2(n4656), .A(n4759), .B(n3567), .ZN(n3569)
         );
  NAND2_X1 U4379 ( .A1(n3661), .A2(n4366), .ZN(n3568) );
  OAI211_X1 U4380 ( .C1(n3570), .C2(n3664), .A(n3569), .B(n3568), .ZN(U3225)
         );
  NAND2_X1 U4381 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  XOR2_X1 U4382 ( .A(n3574), .B(n3573), .Z(n3579) );
  OAI22_X1 U4383 ( .A1(n3608), .A2(n4653), .B1(n3659), .B2(n4481), .ZN(n3577)
         );
  INV_X1 U4384 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3575) );
  OAI22_X1 U4385 ( .A1(n3652), .A2(n4480), .B1(STATE_REG_SCAN_IN), .B2(n3575), 
        .ZN(n3576) );
  AOI211_X1 U4386 ( .C1(n4233), .C2(n3661), .A(n3577), .B(n3576), .ZN(n3578)
         );
  OAI21_X1 U4387 ( .B1(n3579), .B2(n3664), .A(n3578), .ZN(U3226) );
  NAND2_X1 U4388 ( .A1(n3581), .A2(n3580), .ZN(n3583) );
  NAND2_X1 U4389 ( .A1(n3583), .A2(n3582), .ZN(n3590) );
  NAND2_X1 U4390 ( .A1(n3585), .A2(n3584), .ZN(n3586) );
  AOI21_X1 U4391 ( .B1(n3589), .B2(n3587), .A(n3586), .ZN(n3588) );
  AOI21_X1 U4392 ( .B1(n3590), .B2(n3589), .A(n3588), .ZN(n3595) );
  OAI22_X1 U4393 ( .A1(n4305), .A2(n3659), .B1(n4653), .B2(n4304), .ZN(n3593)
         );
  OAI22_X1 U4394 ( .A1(n3652), .A2(n4312), .B1(STATE_REG_SCAN_IN), .B2(n3591), 
        .ZN(n3592) );
  AOI211_X1 U4395 ( .C1(n4314), .C2(n3661), .A(n3593), .B(n3592), .ZN(n3594)
         );
  OAI21_X1 U4396 ( .B1(n3595), .B2(n3664), .A(n3594), .ZN(U3230) );
  XOR2_X1 U4397 ( .A(n3597), .B(n3596), .Z(n3598) );
  XNOR2_X1 U4398 ( .A(n3599), .B(n3598), .ZN(n3600) );
  NAND2_X1 U4399 ( .A1(n3600), .A2(n4663), .ZN(n3603) );
  INV_X1 U4400 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4014) );
  NOR2_X1 U4401 ( .A1(STATE_REG_SCAN_IN), .A2(n4014), .ZN(n4712) );
  OAI22_X1 U4402 ( .A1(n4431), .A2(n4653), .B1(n3659), .B2(n4542), .ZN(n3601)
         );
  AOI211_X1 U4403 ( .C1(n4428), .C2(n4656), .A(n4712), .B(n3601), .ZN(n3602)
         );
  OAI211_X1 U4404 ( .C1(n4668), .C2(n3604), .A(n3603), .B(n3602), .ZN(U3231)
         );
  AOI21_X1 U4405 ( .B1(n3607), .B2(n3606), .A(n3605), .ZN(n3612) );
  OAI22_X1 U4406 ( .A1(n3608), .A2(n3659), .B1(n4653), .B2(n4305), .ZN(n3610)
         );
  OAI22_X1 U4407 ( .A1(n3652), .A2(n4283), .B1(STATE_REG_SCAN_IN), .B2(n4035), 
        .ZN(n3609) );
  AOI211_X1 U4408 ( .C1(n4282), .C2(n3661), .A(n3610), .B(n3609), .ZN(n3611)
         );
  OAI21_X1 U4409 ( .B1(n3612), .B2(n3664), .A(n3611), .ZN(U3232) );
  XNOR2_X1 U4410 ( .A(n3614), .B(n3613), .ZN(n3615) );
  XNOR2_X1 U4411 ( .A(n3541), .B(n3615), .ZN(n3623) );
  NOR2_X1 U4412 ( .A1(STATE_REG_SCAN_IN), .A2(n3616), .ZN(n4701) );
  OAI22_X1 U4413 ( .A1(n4431), .A2(n3659), .B1(n4653), .B2(n3617), .ZN(n3618)
         );
  AOI211_X1 U4414 ( .C1(n3619), .C2(n4656), .A(n4701), .B(n3618), .ZN(n3622)
         );
  NAND2_X1 U4415 ( .A1(n3661), .A2(n3620), .ZN(n3621) );
  OAI211_X1 U4416 ( .C1(n3623), .C2(n3664), .A(n3622), .B(n3621), .ZN(U3233)
         );
  OAI21_X1 U4417 ( .B1(n3626), .B2(n3624), .A(n3625), .ZN(n3627) );
  NAND2_X1 U4418 ( .A1(n3627), .A2(n4663), .ZN(n3634) );
  AOI22_X1 U4419 ( .A1(n4656), .A2(n3629), .B1(REG3_REG_2__SCAN_IN), .B2(n3628), .ZN(n3633) );
  AOI22_X1 U4420 ( .A1(n3631), .A2(n3835), .B1(n3630), .B2(n2872), .ZN(n3632)
         );
  NAND3_X1 U4421 ( .A1(n3634), .A2(n3633), .A3(n3632), .ZN(U3234) );
  NAND2_X1 U4422 ( .A1(n3636), .A2(n3635), .ZN(n3640) );
  NAND2_X1 U4423 ( .A1(n3638), .A2(n3637), .ZN(n3639) );
  XNOR2_X1 U4424 ( .A(n3640), .B(n3639), .ZN(n3645) );
  OAI22_X1 U4425 ( .A1(n4304), .A2(n3659), .B1(n4653), .B2(n4654), .ZN(n3642)
         );
  NAND2_X1 U4426 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4765) );
  OAI21_X1 U4427 ( .B1(n3652), .B2(n2556), .A(n4765), .ZN(n3641) );
  AOI211_X1 U4428 ( .C1(n3643), .C2(n3661), .A(n3642), .B(n3641), .ZN(n3644)
         );
  OAI21_X1 U4429 ( .B1(n3645), .B2(n3664), .A(n3644), .ZN(U3235) );
  INV_X1 U4430 ( .A(n3647), .ZN(n3648) );
  NOR2_X1 U4431 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  XNOR2_X1 U4432 ( .A(n3646), .B(n3650), .ZN(n3656) );
  INV_X1 U4433 ( .A(n3651), .ZN(n4202) );
  OAI22_X1 U4434 ( .A1(n4481), .A2(n4653), .B1(n3659), .B2(n3803), .ZN(n3654)
         );
  OAI22_X1 U4435 ( .A1(n3652), .A2(n4464), .B1(STATE_REG_SCAN_IN), .B2(n3923), 
        .ZN(n3653) );
  AOI211_X1 U4436 ( .C1(n4202), .C2(n3661), .A(n3654), .B(n3653), .ZN(n3655)
         );
  OAI21_X1 U4437 ( .B1(n3656), .B2(n3664), .A(n3655), .ZN(U3237) );
  NAND2_X1 U4438 ( .A1(n4658), .A2(n3657), .ZN(n3658) );
  XOR2_X1 U4439 ( .A(n4659), .B(n3658), .Z(n3665) );
  NOR2_X1 U4440 ( .A1(STATE_REG_SCAN_IN), .A2(n2518), .ZN(n4738) );
  OAI22_X1 U4441 ( .A1(n4542), .A2(n4653), .B1(n3659), .B2(n4525), .ZN(n3660)
         );
  AOI211_X1 U4442 ( .C1(n4538), .C2(n4656), .A(n4738), .B(n3660), .ZN(n3663)
         );
  NAND2_X1 U4443 ( .A1(n3661), .A2(n4396), .ZN(n3662) );
  OAI211_X1 U4444 ( .C1(n3665), .C2(n3664), .A(n3663), .B(n3662), .ZN(U3238)
         );
  NAND2_X1 U4445 ( .A1(n3666), .A2(DATAI_31_), .ZN(n3887) );
  INV_X1 U4446 ( .A(n3887), .ZN(n3884) );
  NAND2_X1 U4447 ( .A1(n3666), .A2(DATAI_30_), .ZN(n4452) );
  AND2_X1 U4448 ( .A1(n3680), .A2(n4452), .ZN(n3723) );
  NOR2_X1 U4449 ( .A1(n3886), .A2(n3887), .ZN(n3722) );
  INV_X1 U4450 ( .A(n4452), .ZN(n4450) );
  INV_X1 U4451 ( .A(n3707), .ZN(n3667) );
  NOR2_X1 U4452 ( .A1(n3667), .A2(n3706), .ZN(n3800) );
  NAND2_X1 U4453 ( .A1(n3668), .A2(n3671), .ZN(n3739) );
  NAND2_X1 U4454 ( .A1(n3670), .A2(n3669), .ZN(n3767) );
  NAND2_X1 U4455 ( .A1(n3767), .A2(n3671), .ZN(n3787) );
  OAI21_X1 U4456 ( .B1(n4404), .B2(n3739), .A(n3787), .ZN(n3673) );
  INV_X1 U4457 ( .A(n3672), .ZN(n3789) );
  AOI21_X1 U4458 ( .B1(n3673), .B2(n3788), .A(n3789), .ZN(n3676) );
  OAI21_X1 U4459 ( .B1(n3676), .B2(n3675), .A(n3674), .ZN(n3677) );
  NAND2_X1 U4460 ( .A1(n3677), .A2(n3799), .ZN(n3681) );
  NAND2_X1 U4461 ( .A1(n3679), .A2(n3678), .ZN(n3688) );
  NAND2_X1 U4462 ( .A1(n3886), .A2(n3887), .ZN(n3810) );
  OR2_X1 U4463 ( .A1(n3680), .A2(n4452), .ZN(n3721) );
  OAI211_X1 U4464 ( .C1(n3828), .C2(n3684), .A(n3810), .B(n3721), .ZN(n3686)
         );
  AOI211_X1 U4465 ( .C1(n3800), .C2(n3681), .A(n3688), .B(n3686), .ZN(n3690)
         );
  INV_X1 U4466 ( .A(n3682), .ZN(n3683) );
  AOI21_X1 U4467 ( .B1(n3684), .B2(n3828), .A(n3683), .ZN(n3687) );
  NAND2_X1 U4468 ( .A1(n3687), .A2(n3700), .ZN(n3804) );
  INV_X1 U4469 ( .A(n3804), .ZN(n3685) );
  NAND2_X1 U4470 ( .A1(n3890), .A2(n3685), .ZN(n3689) );
  AOI21_X1 U4471 ( .B1(n3688), .B2(n3687), .A(n3686), .ZN(n3811) );
  AOI22_X1 U4472 ( .A1(n3690), .A2(n3807), .B1(n3689), .B2(n3811), .ZN(n3691)
         );
  AOI21_X1 U4473 ( .B1(n3692), .B2(n4450), .A(n3691), .ZN(n3693) );
  AOI211_X1 U4474 ( .C1(n3884), .C2(n3723), .A(n3722), .B(n3693), .ZN(n3818)
         );
  NOR4_X1 U4475 ( .A1(n4274), .A2(n4375), .A3(n3695), .A4(n3694), .ZN(n3697)
         );
  NOR2_X1 U4476 ( .A1(n2648), .A2(n4392), .ZN(n3696) );
  NAND4_X1 U4477 ( .A1(n3697), .A2(n4405), .A3(n3107), .A4(n3696), .ZN(n3705)
         );
  INV_X1 U4478 ( .A(n3698), .ZN(n3703) );
  NAND2_X1 U4479 ( .A1(n3700), .A2(n3699), .ZN(n4201) );
  INV_X1 U4480 ( .A(n4201), .ZN(n4207) );
  NAND2_X1 U4481 ( .A1(n4207), .A2(n3701), .ZN(n3702) );
  NOR4_X1 U4482 ( .A1(n3705), .A2(n3704), .A3(n3703), .A4(n3702), .ZN(n3735)
         );
  NAND2_X1 U4483 ( .A1(n2676), .A2(n4205), .ZN(n4217) );
  INV_X1 U4484 ( .A(n4217), .ZN(n3711) );
  NAND2_X1 U4485 ( .A1(n3708), .A2(n3707), .ZN(n4229) );
  INV_X1 U4486 ( .A(n4229), .ZN(n4238) );
  INV_X1 U4487 ( .A(n4320), .ZN(n3709) );
  NAND4_X1 U4488 ( .A1(n3711), .A2(n4238), .A3(n4364), .A4(n3710), .ZN(n3727)
         );
  INV_X1 U4489 ( .A(n3712), .ZN(n3713) );
  NOR2_X1 U4490 ( .A1(n3714), .A2(n3713), .ZN(n4426) );
  INV_X1 U4491 ( .A(n3715), .ZN(n3716) );
  NOR2_X1 U4492 ( .A1(n3717), .A2(n3716), .ZN(n4303) );
  INV_X1 U4493 ( .A(n4254), .ZN(n3718) );
  XNOR2_X1 U4494 ( .A(n4483), .B(n4268), .ZN(n4262) );
  XNOR2_X1 U4495 ( .A(n4304), .B(n3719), .ZN(n4330) );
  NOR4_X1 U4496 ( .A1(n4303), .A2(n4253), .A3(n4262), .A4(n4330), .ZN(n3720)
         );
  NAND3_X1 U4497 ( .A1(n3721), .A2(n3720), .A3(n3810), .ZN(n3726) );
  INV_X1 U4498 ( .A(n3722), .ZN(n3725) );
  INV_X1 U4499 ( .A(n3723), .ZN(n3724) );
  NAND2_X1 U4500 ( .A1(n3725), .A2(n3724), .ZN(n3809) );
  NOR4_X1 U4501 ( .A1(n3727), .A2(n4426), .A3(n3726), .A4(n3809), .ZN(n3734)
         );
  NOR4_X1 U4502 ( .A1(n3730), .A2(n3729), .A3(n4353), .A4(n3728), .ZN(n3733)
         );
  INV_X1 U4503 ( .A(n4788), .ZN(n4784) );
  NOR4_X1 U4504 ( .A1(n2650), .A2(n4784), .A3(n2962), .A4(n3731), .ZN(n3732)
         );
  NAND4_X1 U4505 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3737)
         );
  OAI21_X1 U4506 ( .B1(n3737), .B2(n3892), .A(n3736), .ZN(n3815) );
  INV_X1 U4507 ( .A(n3738), .ZN(n3781) );
  INV_X1 U4508 ( .A(n3739), .ZN(n3740) );
  OAI211_X1 U4509 ( .C1(n3742), .C2(n3781), .A(n3741), .B(n3740), .ZN(n3786)
         );
  INV_X1 U4510 ( .A(n3743), .ZN(n3747) );
  OAI211_X1 U4511 ( .C1(n3747), .C2(n3746), .A(n3745), .B(n3744), .ZN(n3749)
         );
  NAND3_X1 U4512 ( .A1(n3749), .A2(n3748), .A3(n2649), .ZN(n3752) );
  NAND3_X1 U4513 ( .A1(n3752), .A2(n3751), .A3(n3750), .ZN(n3754) );
  NAND3_X1 U4514 ( .A1(n3754), .A2(n2652), .A3(n3753), .ZN(n3757) );
  NAND4_X1 U4515 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3770), .ZN(n3760)
         );
  INV_X1 U4516 ( .A(n3758), .ZN(n3769) );
  AOI21_X1 U4517 ( .B1(n3760), .B2(n3759), .A(n3769), .ZN(n3762) );
  OAI21_X1 U4518 ( .B1(n3762), .B2(n3761), .A(n3771), .ZN(n3765) );
  NAND3_X1 U4519 ( .A1(n3765), .A2(n3764), .A3(n3763), .ZN(n3778) );
  NOR2_X1 U4520 ( .A1(n3767), .A2(n3766), .ZN(n3777) );
  NOR2_X1 U4521 ( .A1(n3769), .A2(n3768), .ZN(n3773) );
  NAND4_X1 U4522 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3775)
         );
  NAND2_X1 U4523 ( .A1(n3775), .A2(n3774), .ZN(n3776) );
  AOI22_X1 U4524 ( .A1(n3778), .A2(n3777), .B1(n3787), .B2(n3776), .ZN(n3784)
         );
  INV_X1 U4525 ( .A(n3779), .ZN(n3783) );
  INV_X1 U4526 ( .A(n3780), .ZN(n3782) );
  NOR4_X1 U4527 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3785)
         );
  AOI21_X1 U4528 ( .B1(n3787), .B2(n3786), .A(n3785), .ZN(n3790) );
  OAI21_X1 U4529 ( .B1(n3790), .B2(n3789), .A(n3788), .ZN(n3794) );
  INV_X1 U4530 ( .A(n3791), .ZN(n3792) );
  AOI21_X1 U4531 ( .B1(n3794), .B2(n3793), .A(n3792), .ZN(n3796) );
  AOI221_X1 U4532 ( .B1(n3798), .B2(n3797), .C1(n3796), .C2(n3797), .A(n3795), 
        .ZN(n3802) );
  INV_X1 U4533 ( .A(n3799), .ZN(n3801) );
  OAI21_X1 U4534 ( .B1(n3802), .B2(n3801), .A(n3800), .ZN(n3806) );
  NOR2_X1 U4535 ( .A1(n3803), .A2(n3897), .ZN(n3805) );
  AOI211_X1 U4536 ( .C1(n3807), .C2(n3806), .A(n3805), .B(n3804), .ZN(n3808)
         );
  INV_X1 U4537 ( .A(n3808), .ZN(n3812) );
  AOI22_X1 U4538 ( .A1(n3812), .A2(n3811), .B1(n3810), .B2(n3809), .ZN(n3814)
         );
  MUX2_X1 U4539 ( .A(n3815), .B(n3814), .S(n3813), .Z(n3816) );
  OAI21_X1 U4540 ( .B1(n3818), .B2(n3817), .A(n3816), .ZN(n3819) );
  XNOR2_X1 U4541 ( .A(n3819), .B(n3878), .ZN(n3827) );
  NAND2_X1 U4542 ( .A1(n3821), .A2(n3820), .ZN(n3822) );
  OAI211_X1 U4543 ( .C1(n3824), .C2(n3823), .A(B_REG_SCAN_IN), .B(n3822), .ZN(
        n3825) );
  OAI21_X1 U4544 ( .B1(n3827), .B2(n3826), .A(n3825), .ZN(U3239) );
  MUX2_X1 U4545 ( .A(n3828), .B(DATAO_REG_29__SCAN_IN), .S(n3836), .Z(U3579)
         );
  MUX2_X1 U4546 ( .A(n4458), .B(DATAO_REG_28__SCAN_IN), .S(n3836), .Z(U3578)
         );
  MUX2_X1 U4547 ( .A(n4473), .B(DATAO_REG_26__SCAN_IN), .S(n3836), .Z(U3576)
         );
  MUX2_X1 U4548 ( .A(n4490), .B(DATAO_REG_24__SCAN_IN), .S(n3836), .Z(U3574)
         );
  MUX2_X1 U4549 ( .A(n4291), .B(DATAO_REG_22__SCAN_IN), .S(n3836), .Z(U3572)
         );
  MUX2_X1 U4550 ( .A(n4504), .B(DATAO_REG_20__SCAN_IN), .S(n3836), .Z(U3570)
         );
  MUX2_X1 U4551 ( .A(n4522), .B(DATAO_REG_18__SCAN_IN), .S(n3836), .Z(U3568)
         );
  MUX2_X1 U4552 ( .A(n4410), .B(DATAO_REG_15__SCAN_IN), .S(n3836), .Z(U3565)
         );
  MUX2_X1 U4553 ( .A(n4566), .B(DATAO_REG_13__SCAN_IN), .S(n3836), .Z(U3563)
         );
  MUX2_X1 U4554 ( .A(n3829), .B(DATAO_REG_11__SCAN_IN), .S(n3836), .Z(U3561)
         );
  MUX2_X1 U4555 ( .A(n3830), .B(DATAO_REG_10__SCAN_IN), .S(n3836), .Z(U3560)
         );
  MUX2_X1 U4556 ( .A(n3831), .B(DATAO_REG_9__SCAN_IN), .S(n3836), .Z(U3559) );
  MUX2_X1 U4557 ( .A(n3832), .B(DATAO_REG_8__SCAN_IN), .S(n3836), .Z(U3558) );
  MUX2_X1 U4558 ( .A(n3833), .B(DATAO_REG_7__SCAN_IN), .S(n3836), .Z(U3557) );
  MUX2_X1 U4559 ( .A(n3834), .B(DATAO_REG_6__SCAN_IN), .S(n3836), .Z(U3556) );
  MUX2_X1 U4560 ( .A(n4793), .B(DATAO_REG_4__SCAN_IN), .S(n3836), .Z(U3554) );
  MUX2_X1 U4561 ( .A(n3835), .B(DATAO_REG_3__SCAN_IN), .S(n3836), .Z(U3553) );
  MUX2_X1 U4562 ( .A(n2872), .B(DATAO_REG_1__SCAN_IN), .S(n3836), .Z(U3551) );
  XNOR2_X1 U4563 ( .A(n4642), .B(REG1_REG_7__SCAN_IN), .ZN(n3838) );
  AOI21_X1 U4564 ( .B1(n3839), .B2(n3838), .A(n4756), .ZN(n3837) );
  OAI21_X1 U4565 ( .B1(n3839), .B2(n3838), .A(n3837), .ZN(n3848) );
  AOI21_X1 U4566 ( .B1(n4767), .B2(ADDR_REG_7__SCAN_IN), .A(n3840), .ZN(n3847)
         );
  OAI211_X1 U4567 ( .C1(n3843), .C2(n3842), .A(n3841), .B(n4762), .ZN(n3846)
         );
  INV_X1 U4568 ( .A(n4775), .ZN(n3844) );
  NAND2_X1 U4569 ( .A1(n3844), .A2(n4642), .ZN(n3845) );
  NAND4_X1 U4570 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(U3247)
         );
  INV_X1 U4571 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3908) );
  INV_X1 U4572 ( .A(n3849), .ZN(n3851) );
  NAND2_X1 U4573 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4709), .ZN(n4708) );
  INV_X1 U4574 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4000) );
  XNOR2_X1 U4575 ( .A(n3853), .B(n3852), .ZN(n4721) );
  NAND2_X1 U4576 ( .A1(n4721), .A2(REG2_REG_14__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U4577 ( .A1(n4719), .A2(n3853), .ZN(n3854) );
  NAND2_X1 U4578 ( .A1(n4720), .A2(n3854), .ZN(n4733) );
  INV_X1 U4579 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3855) );
  INV_X1 U4580 ( .A(n3869), .ZN(n4844) );
  AOI22_X1 U4581 ( .A1(n3869), .A2(REG2_REG_15__SCAN_IN), .B1(n3855), .B2(
        n4844), .ZN(n4734) );
  NAND2_X1 U4582 ( .A1(n4733), .A2(n4734), .ZN(n4732) );
  NAND2_X1 U4583 ( .A1(n3869), .A2(REG2_REG_15__SCAN_IN), .ZN(n3856) );
  XNOR2_X1 U4584 ( .A(n3857), .B(n4740), .ZN(n4744) );
  NOR2_X1 U4585 ( .A1(n4740), .A2(n3857), .ZN(n3858) );
  INV_X1 U4586 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4587 ( .A1(REG2_REG_17__SCAN_IN), .A2(n4840), .B1(n3873), .B2(
        n4001), .ZN(n4753) );
  AOI22_X1 U4588 ( .A1(REG2_REG_18__SCAN_IN), .A2(n3862), .B1(n4839), .B2(
        n3908), .ZN(n4764) );
  OAI21_X1 U4589 ( .B1(n3908), .B2(n4839), .A(n4761), .ZN(n3861) );
  XNOR2_X1 U4590 ( .A(n3878), .B(REG2_REG_19__SCAN_IN), .ZN(n3860) );
  XNOR2_X1 U4591 ( .A(n3861), .B(n3860), .ZN(n3882) );
  INV_X1 U4592 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4593 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3862), .B1(n4839), .B2(
        n3910), .ZN(n4773) );
  INV_X1 U4594 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3949) );
  INV_X1 U4595 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4559) );
  AOI22_X1 U4596 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4709), .B1(n4847), .B2(
        n4559), .ZN(n4716) );
  NAND2_X1 U4597 ( .A1(n3863), .A2(n4641), .ZN(n3864) );
  NAND2_X1 U4598 ( .A1(n4719), .A2(n3866), .ZN(n3867) );
  NAND2_X1 U4599 ( .A1(n3867), .A2(n4725), .ZN(n4730) );
  INV_X1 U4600 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4601 ( .A1(n3869), .A2(REG1_REG_15__SCAN_IN), .B1(n3868), .B2(
        n4844), .ZN(n4731) );
  NAND2_X1 U4602 ( .A1(n3869), .A2(REG1_REG_15__SCAN_IN), .ZN(n3870) );
  NOR2_X1 U4603 ( .A1(n4740), .A2(n3871), .ZN(n3872) );
  XNOR2_X1 U4604 ( .A(n3871), .B(n4740), .ZN(n4742) );
  AOI22_X1 U4605 ( .A1(REG1_REG_17__SCAN_IN), .A2(n4840), .B1(n3873), .B2(
        n3949), .ZN(n4751) );
  NAND2_X1 U4606 ( .A1(n4773), .A2(n4772), .ZN(n4770) );
  OAI21_X1 U4607 ( .B1(n3910), .B2(n4839), .A(n4770), .ZN(n3875) );
  INV_X1 U4608 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3915) );
  MUX2_X1 U4609 ( .A(REG1_REG_19__SCAN_IN), .B(n3915), .S(n3878), .Z(n3874) );
  XNOR2_X1 U4610 ( .A(n3875), .B(n3874), .ZN(n3880) );
  NAND2_X1 U4611 ( .A1(n4767), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3876) );
  OAI211_X1 U4612 ( .C1(n4775), .C2(n3878), .A(n3877), .B(n3876), .ZN(n3879)
         );
  AOI21_X1 U4613 ( .B1(n3880), .B2(n4771), .A(n3879), .ZN(n3881) );
  OAI21_X1 U4614 ( .B1(n3882), .B2(n4754), .A(n3881), .ZN(U3259) );
  NAND2_X1 U4615 ( .A1(n3883), .A2(n4452), .ZN(n4447) );
  XNOR2_X1 U4616 ( .A(n4447), .B(n3884), .ZN(n4580) );
  NAND2_X1 U4617 ( .A1(n3886), .A2(n3885), .ZN(n4451) );
  OAI21_X1 U4618 ( .B1(n3887), .B2(n4563), .A(n4451), .ZN(n4578) );
  NAND2_X1 U4619 ( .A1(n4578), .A2(n4815), .ZN(n3889) );
  NAND2_X1 U4620 ( .A1(n4806), .A2(REG2_REG_31__SCAN_IN), .ZN(n3888) );
  OAI211_X1 U4621 ( .C1(n4580), .C2(n4441), .A(n3889), .B(n3888), .ZN(U3260)
         );
  XNOR2_X1 U4622 ( .A(n3891), .B(n3890), .ZN(n4463) );
  INV_X1 U4623 ( .A(n4463), .ZN(n3906) );
  NAND2_X1 U4624 ( .A1(n3893), .A2(n3892), .ZN(n3894) );
  AOI21_X1 U4625 ( .B1(n3895), .B2(n3894), .A(n4551), .ZN(n4462) );
  NAND2_X1 U4626 ( .A1(n3896), .A2(n3897), .ZN(n3898) );
  NOR2_X1 U4627 ( .A1(n4461), .A2(n4441), .ZN(n3904) );
  AOI22_X1 U4628 ( .A1(n4412), .A2(n4473), .B1(n4458), .B2(n4411), .ZN(n3902)
         );
  AOI22_X1 U4629 ( .A1(n4806), .A2(REG2_REG_27__SCAN_IN), .B1(n3900), .B2(
        n4810), .ZN(n3901) );
  OAI211_X1 U4630 ( .C1(n4456), .C2(n4416), .A(n3902), .B(n3901), .ZN(n3903)
         );
  OAI21_X1 U4631 ( .B1(n3906), .B2(n4388), .A(n3905), .ZN(n4199) );
  AOI22_X1 U4632 ( .A1(n3908), .A2(keyinput84), .B1(U3149), .B2(keyinput35), 
        .ZN(n3907) );
  OAI221_X1 U4633 ( .B1(n3908), .B2(keyinput84), .C1(U3149), .C2(keyinput35), 
        .A(n3907), .ZN(n3993) );
  INV_X1 U4634 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4336) );
  AOI22_X1 U4635 ( .A1(n3910), .A2(keyinput29), .B1(n4336), .B2(keyinput104), 
        .ZN(n3909) );
  OAI221_X1 U4636 ( .B1(n3910), .B2(keyinput29), .C1(n4336), .C2(keyinput104), 
        .A(n3909), .ZN(n3992) );
  INV_X1 U4637 ( .A(keyinput64), .ZN(n4140) );
  INV_X1 U4638 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3913) );
  INV_X1 U4639 ( .A(keyinput68), .ZN(n3912) );
  AOI22_X1 U4640 ( .A1(n3913), .A2(keyinput125), .B1(ADDR_REG_19__SCAN_IN), 
        .B2(n3912), .ZN(n3911) );
  OAI221_X1 U4641 ( .B1(n3913), .B2(keyinput125), .C1(n3912), .C2(
        ADDR_REG_19__SCAN_IN), .A(n3911), .ZN(n3914) );
  AOI221_X1 U4642 ( .B1(REG1_REG_19__SCAN_IN), .B2(n4140), .C1(n3915), .C2(
        keyinput64), .A(n3914), .ZN(n3932) );
  INV_X1 U4643 ( .A(keyinput88), .ZN(n3918) );
  INV_X1 U4644 ( .A(keyinput89), .ZN(n3917) );
  AOI22_X1 U4645 ( .A1(n3918), .A2(DATAO_REG_0__SCAN_IN), .B1(
        DATAO_REG_12__SCAN_IN), .B2(n3917), .ZN(n3916) );
  OAI221_X1 U4646 ( .B1(n3918), .B2(DATAO_REG_0__SCAN_IN), .C1(n3917), .C2(
        DATAO_REG_12__SCAN_IN), .A(n3916), .ZN(n3930) );
  INV_X1 U4647 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3921) );
  INV_X1 U4648 ( .A(keyinput111), .ZN(n3920) );
  AOI22_X1 U4649 ( .A1(n3921), .A2(keyinput124), .B1(ADDR_REG_3__SCAN_IN), 
        .B2(n3920), .ZN(n3919) );
  OAI221_X1 U4650 ( .B1(n3921), .B2(keyinput124), .C1(n3920), .C2(
        ADDR_REG_3__SCAN_IN), .A(n3919), .ZN(n3929) );
  AOI22_X1 U4651 ( .A1(n2746), .A2(keyinput16), .B1(keyinput56), .B2(n3923), 
        .ZN(n3922) );
  OAI221_X1 U4652 ( .B1(n2746), .B2(keyinput16), .C1(n3923), .C2(keyinput56), 
        .A(n3922), .ZN(n3928) );
  INV_X1 U4653 ( .A(keyinput91), .ZN(n3926) );
  INV_X1 U4654 ( .A(keyinput28), .ZN(n3925) );
  AOI22_X1 U4655 ( .A1(n3926), .A2(DATAO_REG_5__SCAN_IN), .B1(
        DATAO_REG_2__SCAN_IN), .B2(n3925), .ZN(n3924) );
  OAI221_X1 U4656 ( .B1(n3926), .B2(DATAO_REG_5__SCAN_IN), .C1(n3925), .C2(
        DATAO_REG_2__SCAN_IN), .A(n3924), .ZN(n3927) );
  NOR4_X1 U4657 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3931)
         );
  OAI211_X1 U4658 ( .C1(keyinput72), .C2(n2448), .A(n3932), .B(n3931), .ZN(
        n3991) );
  INV_X1 U4659 ( .A(keyinput27), .ZN(n3935) );
  INV_X1 U4660 ( .A(keyinput45), .ZN(n3934) );
  AOI22_X1 U4661 ( .A1(n3935), .A2(DATAO_REG_23__SCAN_IN), .B1(
        DATAO_REG_25__SCAN_IN), .B2(n3934), .ZN(n3933) );
  OAI221_X1 U4662 ( .B1(n3935), .B2(DATAO_REG_23__SCAN_IN), .C1(n3934), .C2(
        DATAO_REG_25__SCAN_IN), .A(n3933), .ZN(n3947) );
  INV_X1 U4663 ( .A(keyinput69), .ZN(n3938) );
  INV_X1 U4664 ( .A(keyinput17), .ZN(n3937) );
  AOI22_X1 U4665 ( .A1(n3938), .A2(DATAO_REG_19__SCAN_IN), .B1(
        DATAO_REG_21__SCAN_IN), .B2(n3937), .ZN(n3936) );
  OAI221_X1 U4666 ( .B1(n3938), .B2(DATAO_REG_19__SCAN_IN), .C1(n3937), .C2(
        DATAO_REG_21__SCAN_IN), .A(n3936), .ZN(n3946) );
  INV_X1 U4667 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3941) );
  INV_X1 U4668 ( .A(keyinput108), .ZN(n3940) );
  AOI22_X1 U4669 ( .A1(n3941), .A2(keyinput8), .B1(DATAO_REG_30__SCAN_IN), 
        .B2(n3940), .ZN(n3939) );
  OAI221_X1 U4670 ( .B1(n3941), .B2(keyinput8), .C1(n3940), .C2(
        DATAO_REG_30__SCAN_IN), .A(n3939), .ZN(n3945) );
  INV_X1 U4671 ( .A(keyinput25), .ZN(n3943) );
  AOI22_X1 U4672 ( .A1(n2726), .A2(keyinput18), .B1(DATAO_REG_27__SCAN_IN), 
        .B2(n3943), .ZN(n3942) );
  OAI221_X1 U4673 ( .B1(n2726), .B2(keyinput18), .C1(n3943), .C2(
        DATAO_REG_27__SCAN_IN), .A(n3942), .ZN(n3944) );
  NOR4_X1 U4674 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3989)
         );
  AOI22_X1 U4675 ( .A1(n3227), .A2(keyinput34), .B1(n3949), .B2(keyinput118), 
        .ZN(n3948) );
  OAI221_X1 U4676 ( .B1(n3227), .B2(keyinput34), .C1(n3949), .C2(keyinput118), 
        .A(n3948), .ZN(n3960) );
  AOI22_X1 U4677 ( .A1(n3951), .A2(keyinput61), .B1(keyinput23), .B2(n2794), 
        .ZN(n3950) );
  OAI221_X1 U4678 ( .B1(n3951), .B2(keyinput61), .C1(n2794), .C2(keyinput23), 
        .A(n3950), .ZN(n3959) );
  INV_X1 U4679 ( .A(keyinput47), .ZN(n4152) );
  INV_X1 U4680 ( .A(keyinput78), .ZN(n3953) );
  AOI22_X1 U4681 ( .A1(n4152), .A2(DATAO_REG_16__SCAN_IN), .B1(
        DATAO_REG_17__SCAN_IN), .B2(n3953), .ZN(n3952) );
  OAI221_X1 U4682 ( .B1(n4152), .B2(DATAO_REG_16__SCAN_IN), .C1(n3953), .C2(
        DATAO_REG_17__SCAN_IN), .A(n3952), .ZN(n3958) );
  INV_X1 U4683 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3954) );
  XOR2_X1 U4684 ( .A(n3954), .B(keyinput0), .Z(n3956) );
  XNOR2_X1 U4685 ( .A(IR_REG_31__SCAN_IN), .B(keyinput50), .ZN(n3955) );
  NAND2_X1 U4686 ( .A1(n3956), .A2(n3955), .ZN(n3957) );
  NOR4_X1 U4687 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n3988)
         );
  INV_X1 U4688 ( .A(DATAI_28_), .ZN(n4649) );
  AOI22_X1 U4689 ( .A1(n4649), .A2(keyinput38), .B1(n3962), .B2(keyinput39), 
        .ZN(n3961) );
  OAI221_X1 U4690 ( .B1(n4649), .B2(keyinput38), .C1(n3962), .C2(keyinput39), 
        .A(n3961), .ZN(n3971) );
  INV_X1 U4691 ( .A(IR_REG_29__SCAN_IN), .ZN(n3964) );
  INV_X1 U4692 ( .A(D_REG_14__SCAN_IN), .ZN(n4828) );
  AOI22_X1 U4693 ( .A1(n3964), .A2(keyinput31), .B1(n4828), .B2(keyinput30), 
        .ZN(n3963) );
  OAI221_X1 U4694 ( .B1(n3964), .B2(keyinput31), .C1(n4828), .C2(keyinput30), 
        .A(n3963), .ZN(n3970) );
  INV_X1 U4695 ( .A(DATAI_15_), .ZN(n4843) );
  INV_X1 U4696 ( .A(D_REG_19__SCAN_IN), .ZN(n4825) );
  AOI22_X1 U4697 ( .A1(n4843), .A2(keyinput51), .B1(n4825), .B2(keyinput55), 
        .ZN(n3965) );
  OAI221_X1 U4698 ( .B1(n4843), .B2(keyinput51), .C1(n4825), .C2(keyinput55), 
        .A(n3965), .ZN(n3969) );
  INV_X1 U4699 ( .A(keyinput42), .ZN(n3967) );
  AOI22_X1 U4700 ( .A1(n4651), .A2(keyinput46), .B1(ADDR_REG_18__SCAN_IN), 
        .B2(n3967), .ZN(n3966) );
  OAI221_X1 U4701 ( .B1(n4651), .B2(keyinput46), .C1(n3967), .C2(
        ADDR_REG_18__SCAN_IN), .A(n3966), .ZN(n3968) );
  NOR4_X1 U4702 ( .A1(n3971), .A2(n3970), .A3(n3969), .A4(n3968), .ZN(n3987)
         );
  INV_X1 U4703 ( .A(D_REG_13__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U4704 ( .A1(n3973), .A2(keyinput15), .B1(keyinput19), .B2(n4829), 
        .ZN(n3972) );
  OAI221_X1 U4705 ( .B1(n3973), .B2(keyinput15), .C1(n4829), .C2(keyinput19), 
        .A(n3972), .ZN(n3985) );
  INV_X1 U4706 ( .A(IR_REG_1__SCAN_IN), .ZN(n3976) );
  INV_X1 U4707 ( .A(keyinput106), .ZN(n3975) );
  AOI22_X1 U4708 ( .A1(n3976), .A2(keyinput7), .B1(DATAO_REG_31__SCAN_IN), 
        .B2(n3975), .ZN(n3974) );
  OAI221_X1 U4709 ( .B1(n3976), .B2(keyinput7), .C1(n3975), .C2(
        DATAO_REG_31__SCAN_IN), .A(n3974), .ZN(n3984) );
  INV_X1 U4710 ( .A(IR_REG_10__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4711 ( .A1(n3979), .A2(keyinput10), .B1(keyinput14), .B2(n3978), 
        .ZN(n3977) );
  OAI221_X1 U4712 ( .B1(n3979), .B2(keyinput10), .C1(n3978), .C2(keyinput14), 
        .A(n3977), .ZN(n3983) );
  XNOR2_X1 U4713 ( .A(IR_REG_5__SCAN_IN), .B(keyinput26), .ZN(n3981) );
  XNOR2_X1 U4714 ( .A(DATAI_4_), .B(keyinput22), .ZN(n3980) );
  NAND2_X1 U4715 ( .A1(n3981), .A2(n3980), .ZN(n3982) );
  NOR4_X1 U4716 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3986)
         );
  NAND4_X1 U4717 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3990)
         );
  NOR4_X1 U4718 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n4136)
         );
  AOI22_X1 U4719 ( .A1(n3118), .A2(keyinput6), .B1(n3995), .B2(keyinput13), 
        .ZN(n3994) );
  OAI221_X1 U4720 ( .B1(n3118), .B2(keyinput6), .C1(n3995), .C2(keyinput13), 
        .A(n3994), .ZN(n4008) );
  INV_X1 U4721 ( .A(keyinput113), .ZN(n3997) );
  AOI22_X1 U4722 ( .A1(n3998), .A2(keyinput3), .B1(ADDR_REG_5__SCAN_IN), .B2(
        n3997), .ZN(n3996) );
  OAI221_X1 U4723 ( .B1(n3998), .B2(keyinput3), .C1(n3997), .C2(
        ADDR_REG_5__SCAN_IN), .A(n3996), .ZN(n4007) );
  AOI22_X1 U4724 ( .A1(n4001), .A2(keyinput83), .B1(keyinput63), .B2(n4000), 
        .ZN(n3999) );
  OAI221_X1 U4725 ( .B1(n4001), .B2(keyinput83), .C1(n4000), .C2(keyinput63), 
        .A(n3999), .ZN(n4006) );
  INV_X1 U4726 ( .A(keyinput48), .ZN(n4004) );
  INV_X1 U4727 ( .A(keyinput43), .ZN(n4003) );
  AOI22_X1 U4728 ( .A1(n4004), .A2(ADDR_REG_14__SCAN_IN), .B1(
        ADDR_REG_17__SCAN_IN), .B2(n4003), .ZN(n4002) );
  OAI221_X1 U4729 ( .B1(n4004), .B2(ADDR_REG_14__SCAN_IN), .C1(n4003), .C2(
        ADDR_REG_17__SCAN_IN), .A(n4002), .ZN(n4005) );
  NOR4_X1 U4730 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4135)
         );
  AOI22_X1 U4731 ( .A1(n4010), .A2(keyinput98), .B1(n2518), .B2(keyinput103), 
        .ZN(n4009) );
  OAI221_X1 U4732 ( .B1(n4010), .B2(keyinput98), .C1(n2518), .C2(keyinput103), 
        .A(n4009), .ZN(n4020) );
  INV_X1 U4733 ( .A(D_REG_8__SCAN_IN), .ZN(n4832) );
  INV_X1 U4734 ( .A(D_REG_21__SCAN_IN), .ZN(n4824) );
  AOI22_X1 U4735 ( .A1(n4832), .A2(keyinput102), .B1(n4824), .B2(keyinput107), 
        .ZN(n4011) );
  OAI221_X1 U4736 ( .B1(n4832), .B2(keyinput102), .C1(n4824), .C2(keyinput107), 
        .A(n4011), .ZN(n4019) );
  INV_X1 U4737 ( .A(keyinput110), .ZN(n4013) );
  AOI22_X1 U4738 ( .A1(n4014), .A2(keyinput115), .B1(DATAO_REG_14__SCAN_IN), 
        .B2(n4013), .ZN(n4012) );
  OAI221_X1 U4739 ( .B1(n4014), .B2(keyinput115), .C1(n4013), .C2(
        DATAO_REG_14__SCAN_IN), .A(n4012), .ZN(n4018) );
  INV_X1 U4740 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4016) );
  INV_X1 U4741 ( .A(DATAI_16_), .ZN(n4841) );
  AOI22_X1 U4742 ( .A1(n4016), .A2(keyinput114), .B1(keyinput119), .B2(n4841), 
        .ZN(n4015) );
  OAI221_X1 U4743 ( .B1(n4016), .B2(keyinput114), .C1(n4841), .C2(keyinput119), 
        .A(n4015), .ZN(n4017) );
  NOR4_X1 U4744 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4134)
         );
  INV_X1 U4745 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4022) );
  INV_X1 U4746 ( .A(DATAI_0_), .ZN(n4856) );
  AOI22_X1 U4747 ( .A1(n4022), .A2(keyinput70), .B1(keyinput75), .B2(n4856), 
        .ZN(n4021) );
  OAI221_X1 U4748 ( .B1(n4022), .B2(keyinput70), .C1(n4856), .C2(keyinput75), 
        .A(n4021), .ZN(n4031) );
  INV_X1 U4749 ( .A(DATAI_26_), .ZN(n4024) );
  AOI22_X1 U4750 ( .A1(n4025), .A2(keyinput1), .B1(keyinput5), .B2(n4024), 
        .ZN(n4023) );
  OAI221_X1 U4751 ( .B1(n4025), .B2(keyinput1), .C1(n4024), .C2(keyinput5), 
        .A(n4023), .ZN(n4030) );
  INV_X1 U4752 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4028) );
  INV_X1 U4753 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4754 ( .A1(n4028), .A2(keyinput37), .B1(n4027), .B2(keyinput49), 
        .ZN(n4026) );
  OAI221_X1 U4755 ( .B1(n4028), .B2(keyinput37), .C1(n4027), .C2(keyinput49), 
        .A(n4026), .ZN(n4029) );
  NOR3_X1 U4756 ( .A1(n4031), .A2(n4030), .A3(n4029), .ZN(n4050) );
  AOI22_X1 U4757 ( .A1(n2440), .A2(keyinput100), .B1(keyinput92), .B2(n2377), 
        .ZN(n4032) );
  OAI221_X1 U4758 ( .B1(n2440), .B2(keyinput100), .C1(n2377), .C2(keyinput92), 
        .A(n4032), .ZN(n4037) );
  INV_X1 U4759 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U4760 ( .A1(n4035), .A2(keyinput36), .B1(keyinput44), .B2(n4034), 
        .ZN(n4033) );
  OAI221_X1 U4761 ( .B1(n4035), .B2(keyinput36), .C1(n4034), .C2(keyinput44), 
        .A(n4033), .ZN(n4036) );
  NOR2_X1 U4762 ( .A1(n4037), .A2(n4036), .ZN(n4049) );
  AOI22_X1 U4763 ( .A1(n4626), .A2(keyinput81), .B1(n4823), .B2(keyinput85), 
        .ZN(n4038) );
  OAI221_X1 U4764 ( .B1(n4626), .B2(keyinput81), .C1(n4823), .C2(keyinput85), 
        .A(n4038), .ZN(n4042) );
  AOI22_X1 U4765 ( .A1(n4040), .A2(keyinput74), .B1(keyinput79), .B2(n4604), 
        .ZN(n4039) );
  OAI221_X1 U4766 ( .B1(n4040), .B2(keyinput74), .C1(n4604), .C2(keyinput79), 
        .A(n4039), .ZN(n4041) );
  NOR2_X1 U4767 ( .A1(n4042), .A2(n4041), .ZN(n4048) );
  AOI22_X1 U4768 ( .A1(n2479), .A2(keyinput32), .B1(keyinput60), .B2(n2346), 
        .ZN(n4043) );
  OAI221_X1 U4769 ( .B1(n2479), .B2(keyinput32), .C1(n2346), .C2(keyinput60), 
        .A(n4043), .ZN(n4046) );
  AOI22_X1 U4770 ( .A1(n2342), .A2(keyinput40), .B1(n4830), .B2(keyinput52), 
        .ZN(n4044) );
  OAI221_X1 U4771 ( .B1(n2342), .B2(keyinput40), .C1(n4830), .C2(keyinput52), 
        .A(n4044), .ZN(n4045) );
  NOR2_X1 U4772 ( .A1(n4046), .A2(n4045), .ZN(n4047) );
  NAND4_X1 U4773 ( .A1(n4050), .A2(n4049), .A3(n4048), .A4(n4047), .ZN(n4082)
         );
  INV_X1 U4774 ( .A(D_REG_28__SCAN_IN), .ZN(n4821) );
  AOI22_X1 U4775 ( .A1(n4052), .A2(keyinput4), .B1(n4821), .B2(keyinput12), 
        .ZN(n4051) );
  OAI221_X1 U4776 ( .B1(n4052), .B2(keyinput4), .C1(n4821), .C2(keyinput12), 
        .A(n4051), .ZN(n4056) );
  INV_X1 U4777 ( .A(D_REG_4__SCAN_IN), .ZN(n4833) );
  AOI22_X1 U4778 ( .A1(n4054), .A2(keyinput116), .B1(n4833), .B2(keyinput120), 
        .ZN(n4053) );
  OAI221_X1 U4779 ( .B1(n4054), .B2(keyinput116), .C1(n4833), .C2(keyinput120), 
        .A(n4053), .ZN(n4055) );
  NOR2_X1 U4780 ( .A1(n4056), .A2(n4055), .ZN(n4080) );
  INV_X1 U4781 ( .A(keyinput2), .ZN(n4059) );
  INV_X1 U4782 ( .A(keyinput58), .ZN(n4058) );
  AOI22_X1 U4783 ( .A1(n4059), .A2(ADDR_REG_0__SCAN_IN), .B1(
        ADDR_REG_1__SCAN_IN), .B2(n4058), .ZN(n4057) );
  OAI221_X1 U4784 ( .B1(n4059), .B2(ADDR_REG_0__SCAN_IN), .C1(n4058), .C2(
        ADDR_REG_1__SCAN_IN), .A(n4057), .ZN(n4063) );
  INV_X1 U4785 ( .A(keyinput117), .ZN(n4061) );
  AOI22_X1 U4786 ( .A1(n4892), .A2(keyinput11), .B1(ADDR_REG_4__SCAN_IN), .B2(
        n4061), .ZN(n4060) );
  OAI221_X1 U4787 ( .B1(n4892), .B2(keyinput11), .C1(n4061), .C2(
        ADDR_REG_4__SCAN_IN), .A(n4060), .ZN(n4062) );
  NOR2_X1 U4788 ( .A1(n4063), .A2(n4062), .ZN(n4079) );
  INV_X1 U4789 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4065) );
  INV_X1 U4790 ( .A(D_REG_30__SCAN_IN), .ZN(n4819) );
  AOI22_X1 U4791 ( .A1(n4065), .A2(keyinput123), .B1(n4819), .B2(keyinput126), 
        .ZN(n4064) );
  OAI221_X1 U4792 ( .B1(n4065), .B2(keyinput123), .C1(n4819), .C2(keyinput126), 
        .A(n4064), .ZN(n4069) );
  INV_X1 U4793 ( .A(D_REG_29__SCAN_IN), .ZN(n4820) );
  AOI22_X1 U4794 ( .A1(n4067), .A2(keyinput67), .B1(n4820), .B2(keyinput71), 
        .ZN(n4066) );
  OAI221_X1 U4795 ( .B1(n4067), .B2(keyinput67), .C1(n4820), .C2(keyinput71), 
        .A(n4066), .ZN(n4068) );
  NOR2_X1 U4796 ( .A1(n4069), .A2(n4068), .ZN(n4078) );
  INV_X1 U4797 ( .A(DATAI_1_), .ZN(n4072) );
  INV_X1 U4798 ( .A(IR_REG_16__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4799 ( .A1(n4072), .A2(keyinput95), .B1(n4071), .B2(keyinput99), 
        .ZN(n4070) );
  OAI221_X1 U4800 ( .B1(n4072), .B2(keyinput95), .C1(n4071), .C2(keyinput99), 
        .A(n4070), .ZN(n4076) );
  AOI22_X1 U4801 ( .A1(n4827), .A2(keyinput105), .B1(keyinput97), .B2(n4074), 
        .ZN(n4073) );
  OAI221_X1 U4802 ( .B1(n4827), .B2(keyinput105), .C1(n4074), .C2(keyinput97), 
        .A(n4073), .ZN(n4075) );
  NOR2_X1 U4803 ( .A1(n4076), .A2(n4075), .ZN(n4077) );
  NAND4_X1 U4804 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4081)
         );
  OR2_X1 U4805 ( .A1(n4082), .A2(n4081), .ZN(n4132) );
  INV_X1 U4806 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4672) );
  INV_X1 U4807 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U4808 ( .A1(n4672), .A2(keyinput122), .B1(n4084), .B2(keyinput77), 
        .ZN(n4083) );
  OAI221_X1 U4809 ( .B1(n4672), .B2(keyinput122), .C1(n4084), .C2(keyinput77), 
        .A(n4083), .ZN(n4088) );
  AOI22_X1 U4810 ( .A1(n2429), .A2(keyinput96), .B1(n4086), .B2(keyinput112), 
        .ZN(n4085) );
  OAI221_X1 U4811 ( .B1(n2429), .B2(keyinput96), .C1(n4086), .C2(keyinput112), 
        .A(n4085), .ZN(n4087) );
  NOR2_X1 U4812 ( .A1(n4088), .A2(n4087), .ZN(n4096) );
  INV_X1 U4813 ( .A(DATAI_23_), .ZN(n4837) );
  INV_X1 U4814 ( .A(DATAI_18_), .ZN(n4838) );
  AOI22_X1 U4815 ( .A1(n4837), .A2(keyinput101), .B1(keyinput109), .B2(n4838), 
        .ZN(n4089) );
  OAI221_X1 U4816 ( .B1(n4837), .B2(keyinput101), .C1(n4838), .C2(keyinput109), 
        .A(n4089), .ZN(n4094) );
  INV_X1 U4817 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4092) );
  INV_X1 U4818 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U4819 ( .A1(n4092), .A2(keyinput82), .B1(keyinput86), .B2(n4091), 
        .ZN(n4090) );
  OAI221_X1 U4820 ( .B1(n4092), .B2(keyinput82), .C1(n4091), .C2(keyinput86), 
        .A(n4090), .ZN(n4093) );
  NOR2_X1 U4821 ( .A1(n4094), .A2(n4093), .ZN(n4095) );
  AND2_X1 U4822 ( .A1(n4096), .A2(n4095), .ZN(n4130) );
  AOI22_X1 U4823 ( .A1(n4831), .A2(keyinput73), .B1(keyinput93), .B2(n4098), 
        .ZN(n4097) );
  OAI221_X1 U4824 ( .B1(n4831), .B2(keyinput73), .C1(n4098), .C2(keyinput93), 
        .A(n4097), .ZN(n4112) );
  AOI22_X1 U4825 ( .A1(n4101), .A2(keyinput21), .B1(keyinput33), .B2(n4100), 
        .ZN(n4099) );
  OAI221_X1 U4826 ( .B1(n4101), .B2(keyinput21), .C1(n4100), .C2(keyinput33), 
        .A(n4099), .ZN(n4111) );
  XNOR2_X1 U4827 ( .A(IR_REG_28__SCAN_IN), .B(keyinput41), .ZN(n4105) );
  XNOR2_X1 U4828 ( .A(IR_REG_14__SCAN_IN), .B(keyinput87), .ZN(n4104) );
  XNOR2_X1 U4829 ( .A(IR_REG_26__SCAN_IN), .B(keyinput121), .ZN(n4103) );
  XNOR2_X1 U4830 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput57), .ZN(n4102) );
  AND4_X1 U4831 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4109)
         );
  XNOR2_X1 U4832 ( .A(keyinput54), .B(DATAI_20_), .ZN(n4108) );
  XNOR2_X1 U4833 ( .A(IR_REG_11__SCAN_IN), .B(keyinput62), .ZN(n4107) );
  XNOR2_X1 U4834 ( .A(DATAI_3_), .B(keyinput59), .ZN(n4106) );
  NAND4_X1 U4835 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4110)
         );
  NOR3_X1 U4836 ( .A1(n4112), .A2(n4111), .A3(n4110), .ZN(n4129) );
  XNOR2_X1 U4837 ( .A(REG0_REG_22__SCAN_IN), .B(keyinput9), .ZN(n4116) );
  XNOR2_X1 U4838 ( .A(IR_REG_17__SCAN_IN), .B(keyinput53), .ZN(n4115) );
  XNOR2_X1 U4839 ( .A(IR_REG_9__SCAN_IN), .B(keyinput76), .ZN(n4114) );
  XNOR2_X1 U4840 ( .A(IR_REG_2__SCAN_IN), .B(keyinput20), .ZN(n4113) );
  AND4_X1 U4841 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4122)
         );
  XNOR2_X1 U4842 ( .A(keyinput127), .B(REG3_REG_3__SCAN_IN), .ZN(n4121) );
  XNOR2_X1 U4843 ( .A(keyinput65), .B(n4617), .ZN(n4118) );
  XNOR2_X1 U4844 ( .A(keyinput66), .B(n2639), .ZN(n4117) );
  NOR2_X1 U4845 ( .A1(n4118), .A2(n4117), .ZN(n4120) );
  XNOR2_X1 U4846 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput94), .ZN(n4119) );
  NAND4_X1 U4847 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4124)
         );
  INV_X1 U4848 ( .A(D_REG_31__SCAN_IN), .ZN(n4818) );
  XNOR2_X1 U4849 ( .A(n4818), .B(keyinput80), .ZN(n4123) );
  NOR2_X1 U4850 ( .A1(n4124), .A2(n4123), .ZN(n4128) );
  INV_X1 U4851 ( .A(D_REG_27__SCAN_IN), .ZN(n4822) );
  XNOR2_X1 U4852 ( .A(n4822), .B(keyinput24), .ZN(n4126) );
  INV_X1 U4853 ( .A(D_REG_17__SCAN_IN), .ZN(n4826) );
  XNOR2_X1 U4854 ( .A(n4826), .B(keyinput90), .ZN(n4125) );
  NOR2_X1 U4855 ( .A1(n4126), .A2(n4125), .ZN(n4127) );
  NAND4_X1 U4856 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(n4131)
         );
  NOR2_X1 U4857 ( .A1(n4132), .A2(n4131), .ZN(n4133) );
  AND4_X1 U4858 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4197)
         );
  NOR2_X1 U4859 ( .A1(keyinput77), .A2(keyinput94), .ZN(n4137) );
  NAND3_X1 U4860 ( .A1(keyinput127), .A2(keyinput2), .A3(n4137), .ZN(n4138) );
  NOR3_X1 U4861 ( .A1(keyinput58), .A2(keyinput11), .A3(n4138), .ZN(n4150) );
  INV_X1 U4862 ( .A(keyinput35), .ZN(n4148) );
  NOR4_X1 U4863 ( .A1(keyinput124), .A2(keyinput88), .A3(keyinput89), .A4(
        keyinput91), .ZN(n4139) );
  NAND3_X1 U4864 ( .A1(keyinput28), .A2(keyinput16), .A3(n4139), .ZN(n4147) );
  NOR4_X1 U4865 ( .A1(keyinput125), .A2(keyinput29), .A3(keyinput104), .A4(
        keyinput84), .ZN(n4145) );
  NOR3_X1 U4866 ( .A1(keyinput76), .A2(keyinput68), .A3(n4140), .ZN(n4144) );
  NOR4_X1 U4867 ( .A1(keyinput3), .A2(keyinput6), .A3(keyinput43), .A4(
        keyinput83), .ZN(n4143) );
  NAND3_X1 U4868 ( .A1(keyinput48), .A2(keyinput13), .A3(keyinput113), .ZN(
        n4141) );
  NOR2_X1 U4869 ( .A1(keyinput117), .A2(n4141), .ZN(n4142) );
  NAND4_X1 U4870 ( .A1(n4145), .A2(n4144), .A3(n4143), .A4(n4142), .ZN(n4146)
         );
  NOR4_X1 U4871 ( .A1(keyinput111), .A2(n4148), .A3(n4147), .A4(n4146), .ZN(
        n4149) );
  NAND4_X1 U4872 ( .A1(keyinput56), .A2(keyinput122), .A3(n4150), .A4(n4149), 
        .ZN(n4194) );
  NAND4_X1 U4873 ( .A1(keyinput7), .A2(keyinput10), .A3(keyinput14), .A4(
        keyinput15), .ZN(n4151) );
  NOR3_X1 U4874 ( .A1(keyinput19), .A2(keyinput22), .A3(n4151), .ZN(n4162) );
  NOR4_X1 U4875 ( .A1(keyinput23), .A2(keyinput0), .A3(keyinput50), .A4(n4152), 
        .ZN(n4153) );
  NAND3_X1 U4876 ( .A1(keyinput63), .A2(keyinput34), .A3(n4153), .ZN(n4160) );
  NOR4_X1 U4877 ( .A1(keyinput17), .A2(keyinput27), .A3(keyinput45), .A4(
        keyinput25), .ZN(n4158) );
  AND4_X1 U4878 ( .A1(keyinput78), .A2(keyinput69), .A3(keyinput18), .A4(
        keyinput8), .ZN(n4157) );
  AND4_X1 U4879 ( .A1(keyinput30), .A2(keyinput38), .A3(keyinput46), .A4(
        keyinput51), .ZN(n4156) );
  INV_X1 U4880 ( .A(keyinput39), .ZN(n4154) );
  NOR4_X1 U4881 ( .A1(keyinput26), .A2(keyinput31), .A3(keyinput42), .A4(n4154), .ZN(n4155) );
  NAND4_X1 U4882 ( .A1(n4158), .A2(n4157), .A3(n4156), .A4(n4155), .ZN(n4159)
         );
  NOR4_X1 U4883 ( .A1(keyinput118), .A2(keyinput61), .A3(n4160), .A4(n4159), 
        .ZN(n4161) );
  NAND4_X1 U4884 ( .A1(keyinput108), .A2(keyinput106), .A3(n4162), .A4(n4161), 
        .ZN(n4193) );
  INV_X1 U4885 ( .A(keyinput126), .ZN(n4163) );
  NAND4_X1 U4886 ( .A1(keyinput65), .A2(keyinput109), .A3(keyinput105), .A4(
        n4163), .ZN(n4164) );
  NOR3_X1 U4887 ( .A1(keyinput41), .A2(keyinput101), .A3(n4164), .ZN(n4176) );
  NAND2_X1 U4888 ( .A1(keyinput82), .A2(keyinput74), .ZN(n4165) );
  NOR3_X1 U4889 ( .A1(keyinput75), .A2(keyinput79), .A3(n4165), .ZN(n4166) );
  NAND3_X1 U4890 ( .A1(keyinput86), .A2(keyinput87), .A3(n4166), .ZN(n4174) );
  NAND2_X1 U4891 ( .A1(keyinput70), .A2(keyinput67), .ZN(n4167) );
  NOR3_X1 U4892 ( .A1(keyinput66), .A2(keyinput71), .A3(n4167), .ZN(n4172) );
  NOR4_X1 U4893 ( .A1(keyinput55), .A2(keyinput54), .A3(keyinput59), .A4(
        keyinput62), .ZN(n4171) );
  NAND2_X1 U4894 ( .A1(keyinput114), .A2(keyinput107), .ZN(n4168) );
  NOR3_X1 U4895 ( .A1(keyinput115), .A2(keyinput110), .A3(n4168), .ZN(n4170)
         );
  NOR4_X1 U4896 ( .A1(keyinput99), .A2(keyinput98), .A3(keyinput103), .A4(
        keyinput102), .ZN(n4169) );
  NAND4_X1 U4897 ( .A1(n4172), .A2(n4171), .A3(n4170), .A4(n4169), .ZN(n4173)
         );
  NOR4_X1 U4898 ( .A1(keyinput90), .A2(keyinput95), .A3(n4174), .A4(n4173), 
        .ZN(n4175) );
  NAND4_X1 U4899 ( .A1(keyinput119), .A2(keyinput123), .A3(n4176), .A4(n4175), 
        .ZN(n4192) );
  INV_X1 U4900 ( .A(keyinput21), .ZN(n4177) );
  NAND4_X1 U4901 ( .A1(keyinput5), .A2(keyinput33), .A3(keyinput37), .A4(n4177), .ZN(n4178) );
  NOR3_X1 U4902 ( .A1(keyinput9), .A2(keyinput1), .A3(n4178), .ZN(n4190) );
  NAND2_X1 U4903 ( .A1(keyinput80), .A2(keyinput100), .ZN(n4179) );
  NOR3_X1 U4904 ( .A1(keyinput60), .A2(keyinput92), .A3(n4179), .ZN(n4180) );
  NAND3_X1 U4905 ( .A1(keyinput52), .A2(keyinput32), .A3(n4180), .ZN(n4188) );
  NAND2_X1 U4906 ( .A1(keyinput93), .A2(keyinput73), .ZN(n4181) );
  NOR3_X1 U4907 ( .A1(keyinput85), .A2(keyinput116), .A3(n4181), .ZN(n4186) );
  NOR4_X1 U4908 ( .A1(keyinput49), .A2(keyinput53), .A3(keyinput57), .A4(
        keyinput81), .ZN(n4185) );
  AND4_X1 U4909 ( .A1(keyinput112), .A2(keyinput4), .A3(keyinput12), .A4(
        keyinput24), .ZN(n4184) );
  INV_X1 U4910 ( .A(keyinput96), .ZN(n4182) );
  NOR4_X1 U4911 ( .A1(keyinput120), .A2(keyinput20), .A3(keyinput36), .A4(
        n4182), .ZN(n4183) );
  NAND4_X1 U4912 ( .A1(n4186), .A2(n4185), .A3(n4184), .A4(n4183), .ZN(n4187)
         );
  NOR4_X1 U4913 ( .A1(keyinput44), .A2(keyinput40), .A3(n4188), .A4(n4187), 
        .ZN(n4189) );
  NAND4_X1 U4914 ( .A1(keyinput97), .A2(keyinput121), .A3(n4190), .A4(n4189), 
        .ZN(n4191) );
  NOR4_X1 U4915 ( .A1(n4194), .A2(n4193), .A3(n4192), .A4(n4191), .ZN(n4195)
         );
  OAI21_X1 U4916 ( .B1(keyinput72), .B2(n4195), .A(n2448), .ZN(n4196) );
  NAND2_X1 U4917 ( .A1(n4197), .A2(n4196), .ZN(n4198) );
  XNOR2_X1 U4918 ( .A(n4199), .B(n4198), .ZN(U3263) );
  XOR2_X1 U4919 ( .A(n4201), .B(n4200), .Z(n4469) );
  OAI21_X1 U4920 ( .B1(n4218), .B2(n4464), .A(n3896), .ZN(n4587) );
  INV_X1 U4921 ( .A(n4587), .ZN(n4212) );
  AOI22_X1 U4922 ( .A1(n4412), .A2(n4232), .B1(n4411), .B2(n4466), .ZN(n4204)
         );
  AOI22_X1 U4923 ( .A1(n4806), .A2(REG2_REG_26__SCAN_IN), .B1(n4202), .B2(
        n4810), .ZN(n4203) );
  OAI211_X1 U4924 ( .C1(n4464), .C2(n4416), .A(n4204), .B(n4203), .ZN(n4211)
         );
  NAND2_X1 U4925 ( .A1(n4206), .A2(n4205), .ZN(n4208) );
  XNOR2_X1 U4926 ( .A(n4208), .B(n4207), .ZN(n4209) );
  NAND2_X1 U4927 ( .A1(n4209), .A2(n4789), .ZN(n4467) );
  NOR2_X1 U4928 ( .A1(n4467), .A2(n4806), .ZN(n4210) );
  AOI211_X1 U4929 ( .C1(n4212), .C2(n4802), .A(n4211), .B(n4210), .ZN(n4213)
         );
  OAI21_X1 U4930 ( .B1(n4469), .B2(n4388), .A(n4213), .ZN(U3264) );
  XNOR2_X1 U4931 ( .A(n4214), .B(n4217), .ZN(n4215) );
  NAND2_X1 U4932 ( .A1(n4215), .A2(n4789), .ZN(n4475) );
  XOR2_X1 U4933 ( .A(n4217), .B(n4216), .Z(n4478) );
  NAND2_X1 U4934 ( .A1(n4478), .A2(n4407), .ZN(n4227) );
  INV_X1 U4935 ( .A(n4218), .ZN(n4219) );
  OAI21_X1 U4936 ( .B1(n4230), .B2(n4223), .A(n4219), .ZN(n4591) );
  INV_X1 U4937 ( .A(n4591), .ZN(n4225) );
  AOI22_X1 U4938 ( .A1(n4412), .A2(n4490), .B1(n4411), .B2(n4473), .ZN(n4222)
         );
  AOI22_X1 U4939 ( .A1(n4806), .A2(REG2_REG_25__SCAN_IN), .B1(n4220), .B2(
        n4810), .ZN(n4221) );
  OAI211_X1 U4940 ( .C1(n4223), .C2(n4416), .A(n4222), .B(n4221), .ZN(n4224)
         );
  AOI21_X1 U4941 ( .B1(n4225), .B2(n4802), .A(n4224), .ZN(n4226) );
  OAI211_X1 U4942 ( .C1(n4806), .C2(n4475), .A(n4227), .B(n4226), .ZN(U3265)
         );
  XOR2_X1 U4943 ( .A(n4229), .B(n4228), .Z(n4486) );
  AOI21_X1 U4944 ( .B1(n4231), .B2(n4263), .A(n4230), .ZN(n4594) );
  AOI22_X1 U4945 ( .A1(n4412), .A2(n4483), .B1(n4411), .B2(n4232), .ZN(n4235)
         );
  AOI22_X1 U4946 ( .A1(n4806), .A2(REG2_REG_24__SCAN_IN), .B1(n4233), .B2(
        n4810), .ZN(n4234) );
  OAI211_X1 U4947 ( .C1(n4480), .C2(n4416), .A(n4235), .B(n4234), .ZN(n4242)
         );
  NAND2_X1 U4948 ( .A1(n4237), .A2(n4236), .ZN(n4239) );
  XNOR2_X1 U4949 ( .A(n4239), .B(n4238), .ZN(n4240) );
  NAND2_X1 U4950 ( .A1(n4240), .A2(n4789), .ZN(n4484) );
  NOR2_X1 U4951 ( .A1(n4484), .A2(n4806), .ZN(n4241) );
  AOI211_X1 U4952 ( .C1(n4594), .C2(n4802), .A(n4242), .B(n4241), .ZN(n4243)
         );
  OAI21_X1 U4953 ( .B1(n4486), .B2(n4388), .A(n4243), .ZN(U3266) );
  INV_X1 U4954 ( .A(n4244), .ZN(n4245) );
  OR2_X1 U4955 ( .A1(n4361), .A2(n4245), .ZN(n4248) );
  INV_X1 U4956 ( .A(n4246), .ZN(n4247) );
  NAND2_X1 U4957 ( .A1(n4248), .A2(n4247), .ZN(n4302) );
  NAND2_X1 U4958 ( .A1(n4302), .A2(n4249), .ZN(n4252) );
  INV_X1 U4959 ( .A(n4250), .ZN(n4251) );
  NAND2_X1 U4960 ( .A1(n4252), .A2(n4251), .ZN(n4296) );
  NAND2_X1 U4961 ( .A1(n4296), .A2(n4295), .ZN(n4255) );
  NAND2_X1 U4962 ( .A1(n4255), .A2(n4254), .ZN(n4277) );
  INV_X1 U4963 ( .A(n4274), .ZN(n4276) );
  NAND2_X1 U4964 ( .A1(n4277), .A2(n4276), .ZN(n4257) );
  NAND2_X1 U4965 ( .A1(n4257), .A2(n4256), .ZN(n4259) );
  INV_X1 U4966 ( .A(n4262), .ZN(n4258) );
  XNOR2_X1 U4967 ( .A(n4259), .B(n4258), .ZN(n4260) );
  NAND2_X1 U4968 ( .A1(n4260), .A2(n4789), .ZN(n4492) );
  XOR2_X1 U4969 ( .A(n4262), .B(n4261), .Z(n4494) );
  NAND2_X1 U4970 ( .A1(n4494), .A2(n4407), .ZN(n4272) );
  INV_X1 U4971 ( .A(n4496), .ZN(n4264) );
  OAI21_X1 U4972 ( .B1(n4264), .B2(n4268), .A(n4263), .ZN(n4599) );
  INV_X1 U4973 ( .A(n4599), .ZN(n4270) );
  AOI22_X1 U4974 ( .A1(n4412), .A2(n4291), .B1(n4411), .B2(n4490), .ZN(n4267)
         );
  AOI22_X1 U4975 ( .A1(n4806), .A2(REG2_REG_23__SCAN_IN), .B1(n4265), .B2(
        n4810), .ZN(n4266) );
  OAI211_X1 U4976 ( .C1(n4268), .C2(n4416), .A(n4267), .B(n4266), .ZN(n4269)
         );
  AOI21_X1 U4977 ( .B1(n4270), .B2(n4802), .A(n4269), .ZN(n4271) );
  OAI211_X1 U4978 ( .C1(n4806), .C2(n4492), .A(n4272), .B(n4271), .ZN(U3267)
         );
  OAI21_X1 U4979 ( .B1(n4275), .B2(n4274), .A(n4273), .ZN(n4500) );
  XNOR2_X1 U4980 ( .A(n4277), .B(n4276), .ZN(n4281) );
  NOR2_X1 U4981 ( .A1(n4283), .A2(n4563), .ZN(n4278) );
  AOI21_X1 U4982 ( .B1(n4483), .B2(n4792), .A(n4278), .ZN(n4279) );
  OAI21_X1 U4983 ( .B1(n4305), .B2(n4796), .A(n4279), .ZN(n4280) );
  AOI21_X1 U4984 ( .B1(n4281), .B2(n4789), .A(n4280), .ZN(n4499) );
  AOI22_X1 U4985 ( .A1(n4806), .A2(REG2_REG_22__SCAN_IN), .B1(n4282), .B2(
        n4810), .ZN(n4285) );
  OR2_X1 U4986 ( .A1(n4289), .A2(n4283), .ZN(n4497) );
  NAND3_X1 U4987 ( .A1(n4497), .A2(n4802), .A3(n4496), .ZN(n4284) );
  OAI211_X1 U4988 ( .C1(n4499), .C2(n4806), .A(n4285), .B(n4284), .ZN(n4286)
         );
  INV_X1 U4989 ( .A(n4286), .ZN(n4287) );
  OAI21_X1 U4990 ( .B1(n4500), .B2(n4388), .A(n4287), .ZN(U3268) );
  XNOR2_X1 U4991 ( .A(n4288), .B(n4295), .ZN(n4507) );
  AOI21_X1 U4992 ( .B1(n4290), .B2(n4311), .A(n4289), .ZN(n4601) );
  AOI22_X1 U4993 ( .A1(n4412), .A2(n4504), .B1(n4411), .B2(n4291), .ZN(n4294)
         );
  AOI22_X1 U4994 ( .A1(n4806), .A2(REG2_REG_21__SCAN_IN), .B1(n4292), .B2(
        n4810), .ZN(n4293) );
  OAI211_X1 U4995 ( .C1(n4501), .C2(n4416), .A(n4294), .B(n4293), .ZN(n4299)
         );
  XNOR2_X1 U4996 ( .A(n4296), .B(n4295), .ZN(n4297) );
  NAND2_X1 U4997 ( .A1(n4297), .A2(n4789), .ZN(n4505) );
  NOR2_X1 U4998 ( .A1(n4505), .A2(n4806), .ZN(n4298) );
  AOI211_X1 U4999 ( .C1(n4601), .C2(n4802), .A(n4299), .B(n4298), .ZN(n4300)
         );
  OAI21_X1 U5000 ( .B1(n4507), .B2(n4388), .A(n4300), .ZN(U3269) );
  XNOR2_X1 U5001 ( .A(n4301), .B(n4303), .ZN(n4310) );
  XOR2_X1 U5002 ( .A(n4303), .B(n4302), .Z(n4308) );
  NOR2_X1 U5003 ( .A1(n4304), .A2(n4796), .ZN(n4307) );
  OAI22_X1 U5004 ( .A1(n4305), .A2(n4547), .B1(n4312), .B2(n4563), .ZN(n4306)
         );
  AOI211_X1 U5005 ( .C1(n4308), .C2(n4789), .A(n4307), .B(n4306), .ZN(n4309)
         );
  OAI21_X1 U5006 ( .B1(n4310), .B2(n4435), .A(n4309), .ZN(n4510) );
  INV_X1 U5007 ( .A(n4510), .ZN(n4318) );
  INV_X1 U5008 ( .A(n4310), .ZN(n4511) );
  INV_X1 U5009 ( .A(n4332), .ZN(n4313) );
  OAI21_X1 U5010 ( .B1(n4313), .B2(n4312), .A(n4311), .ZN(n4610) );
  AOI22_X1 U5011 ( .A1(n4806), .A2(REG2_REG_20__SCAN_IN), .B1(n4314), .B2(
        n4810), .ZN(n4315) );
  OAI21_X1 U5012 ( .B1(n4610), .B2(n4441), .A(n4315), .ZN(n4316) );
  AOI21_X1 U5013 ( .B1(n4511), .B2(n4811), .A(n4316), .ZN(n4317) );
  OAI21_X1 U5014 ( .B1(n4318), .B2(n4806), .A(n4317), .ZN(U3270) );
  OAI21_X1 U5015 ( .B1(n4361), .B2(n4320), .A(n4319), .ZN(n4343) );
  INV_X1 U5016 ( .A(n4321), .ZN(n4323) );
  OAI21_X1 U5017 ( .B1(n4343), .B2(n4323), .A(n4322), .ZN(n4324) );
  XNOR2_X1 U5018 ( .A(n4324), .B(n4330), .ZN(n4329) );
  NOR2_X1 U5019 ( .A1(n4325), .A2(n4796), .ZN(n4328) );
  OAI22_X1 U5020 ( .A1(n4326), .A2(n4547), .B1(n4563), .B2(n4333), .ZN(n4327)
         );
  AOI211_X1 U5021 ( .C1(n4329), .C2(n4789), .A(n4328), .B(n4327), .ZN(n4514)
         );
  XNOR2_X1 U5022 ( .A(n4331), .B(n4330), .ZN(n4516) );
  NAND2_X1 U5023 ( .A1(n4516), .A2(n4407), .ZN(n4340) );
  INV_X1 U5024 ( .A(n4342), .ZN(n4334) );
  OAI21_X1 U5025 ( .B1(n4334), .B2(n4333), .A(n4332), .ZN(n4614) );
  INV_X1 U5026 ( .A(n4614), .ZN(n4338) );
  OAI22_X1 U5027 ( .A1(n4815), .A2(n4336), .B1(n4335), .B2(n4350), .ZN(n4337)
         );
  AOI21_X1 U5028 ( .B1(n4338), .B2(n4802), .A(n4337), .ZN(n4339) );
  OAI211_X1 U5029 ( .C1(n4806), .C2(n4514), .A(n4340), .B(n4339), .ZN(U3271)
         );
  OAI211_X1 U5030 ( .C1(n4341), .C2(n2556), .A(n4532), .B(n4342), .ZN(n4518)
         );
  XOR2_X1 U5031 ( .A(n4353), .B(n4343), .Z(n4348) );
  AOI22_X1 U5032 ( .A1(n4345), .A2(n4792), .B1(n4344), .B2(n4791), .ZN(n4346)
         );
  OAI21_X1 U5033 ( .B1(n4654), .B2(n4796), .A(n4346), .ZN(n4347) );
  AOI21_X1 U5034 ( .B1(n4348), .B2(n4789), .A(n4347), .ZN(n4519) );
  OAI21_X1 U5035 ( .B1(n4349), .B2(n4518), .A(n4519), .ZN(n4358) );
  OAI22_X1 U5036 ( .A1(n4815), .A2(n3908), .B1(n4351), .B2(n4350), .ZN(n4357)
         );
  OAI21_X1 U5037 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n4355) );
  INV_X1 U5038 ( .A(n4355), .ZN(n4520) );
  NOR2_X1 U5039 ( .A1(n4520), .A2(n4388), .ZN(n4356) );
  AOI211_X1 U5040 ( .C1(n4815), .C2(n4358), .A(n4357), .B(n4356), .ZN(n4359)
         );
  INV_X1 U5041 ( .A(n4359), .ZN(U3272) );
  INV_X1 U5042 ( .A(n4364), .ZN(n4360) );
  XNOR2_X1 U5043 ( .A(n4361), .B(n4360), .ZN(n4362) );
  NAND2_X1 U5044 ( .A1(n4362), .A2(n4789), .ZN(n4524) );
  XNOR2_X1 U5045 ( .A(n4363), .B(n4364), .ZN(n4527) );
  NAND2_X1 U5046 ( .A1(n4527), .A2(n4407), .ZN(n4373) );
  INV_X1 U5047 ( .A(n4341), .ZN(n4365) );
  OAI21_X1 U5048 ( .B1(n4377), .B2(n4369), .A(n4365), .ZN(n4619) );
  INV_X1 U5049 ( .A(n4619), .ZN(n4371) );
  AOI22_X1 U5050 ( .A1(n4412), .A2(n4539), .B1(n4411), .B2(n4522), .ZN(n4368)
         );
  AOI22_X1 U5051 ( .A1(n4806), .A2(REG2_REG_17__SCAN_IN), .B1(n4366), .B2(
        n4810), .ZN(n4367) );
  OAI211_X1 U5052 ( .C1(n4369), .C2(n4416), .A(n4368), .B(n4367), .ZN(n4370)
         );
  AOI21_X1 U5053 ( .B1(n4371), .B2(n4802), .A(n4370), .ZN(n4372) );
  OAI211_X1 U5054 ( .C1(n4806), .C2(n4524), .A(n4373), .B(n4372), .ZN(U3273)
         );
  OAI21_X1 U5055 ( .B1(n4376), .B2(n4375), .A(n4374), .ZN(n4537) );
  AOI21_X1 U5056 ( .B1(n4657), .B2(n4394), .A(n4377), .ZN(n4533) );
  AOI22_X1 U5057 ( .A1(n4412), .A2(n4410), .B1(n4411), .B2(n4529), .ZN(n4380)
         );
  AOI22_X1 U5058 ( .A1(n4806), .A2(REG2_REG_16__SCAN_IN), .B1(n4378), .B2(
        n4810), .ZN(n4379) );
  OAI211_X1 U5059 ( .C1(n4381), .C2(n4416), .A(n4380), .B(n4379), .ZN(n4386)
         );
  OAI211_X1 U5060 ( .C1(n4384), .C2(n4383), .A(n4382), .B(n4789), .ZN(n4534)
         );
  NOR2_X1 U5061 ( .A1(n4534), .A2(n4806), .ZN(n4385) );
  AOI211_X1 U5062 ( .C1(n4533), .C2(n4802), .A(n4386), .B(n4385), .ZN(n4387)
         );
  OAI21_X1 U5063 ( .B1(n4388), .B2(n4537), .A(n4387), .ZN(U3274) );
  AOI21_X1 U5064 ( .B1(n4389), .B2(n4392), .A(n4551), .ZN(n4391) );
  NAND2_X1 U5065 ( .A1(n4391), .A2(n4390), .ZN(n4541) );
  XNOR2_X1 U5066 ( .A(n4393), .B(n4392), .ZN(n4544) );
  NAND2_X1 U5067 ( .A1(n4544), .A2(n4407), .ZN(n4403) );
  INV_X1 U5068 ( .A(n4409), .ZN(n4395) );
  OAI21_X1 U5069 ( .B1(n4395), .B2(n4399), .A(n4394), .ZN(n4624) );
  INV_X1 U5070 ( .A(n4624), .ZN(n4401) );
  AOI22_X1 U5071 ( .A1(n4412), .A2(n4429), .B1(n4411), .B2(n4539), .ZN(n4398)
         );
  AOI22_X1 U5072 ( .A1(n4806), .A2(REG2_REG_15__SCAN_IN), .B1(n4396), .B2(
        n4810), .ZN(n4397) );
  OAI211_X1 U5073 ( .C1(n4399), .C2(n4416), .A(n4398), .B(n4397), .ZN(n4400)
         );
  AOI21_X1 U5074 ( .B1(n4401), .B2(n4802), .A(n4400), .ZN(n4402) );
  OAI211_X1 U5075 ( .C1(n4806), .C2(n4541), .A(n4403), .B(n4402), .ZN(U3275)
         );
  XOR2_X1 U5076 ( .A(n4404), .B(n4405), .Z(n4552) );
  XNOR2_X1 U5077 ( .A(n4406), .B(n4405), .ZN(n4554) );
  NAND2_X1 U5078 ( .A1(n4554), .A2(n4407), .ZN(n4420) );
  OAI21_X1 U5079 ( .B1(n4408), .B2(n4546), .A(n4409), .ZN(n4628) );
  INV_X1 U5080 ( .A(n4628), .ZN(n4418) );
  AOI22_X1 U5081 ( .A1(n4412), .A2(n4566), .B1(n4411), .B2(n4410), .ZN(n4415)
         );
  AOI22_X1 U5082 ( .A1(n4806), .A2(REG2_REG_14__SCAN_IN), .B1(n4413), .B2(
        n4810), .ZN(n4414) );
  OAI211_X1 U5083 ( .C1(n4546), .C2(n4416), .A(n4415), .B(n4414), .ZN(n4417)
         );
  AOI21_X1 U5084 ( .B1(n4418), .B2(n4802), .A(n4417), .ZN(n4419) );
  OAI211_X1 U5085 ( .C1(n4552), .C2(n4421), .A(n4420), .B(n4419), .ZN(U3276)
         );
  XOR2_X1 U5086 ( .A(n4426), .B(n4422), .Z(n4436) );
  OAI21_X1 U5087 ( .B1(n4425), .B2(n4424), .A(n4423), .ZN(n4427) );
  XNOR2_X1 U5088 ( .A(n4427), .B(n4426), .ZN(n4433) );
  AOI22_X1 U5089 ( .A1(n4429), .A2(n4792), .B1(n4791), .B2(n4428), .ZN(n4430)
         );
  OAI21_X1 U5090 ( .B1(n4431), .B2(n4796), .A(n4430), .ZN(n4432) );
  AOI21_X1 U5091 ( .B1(n4433), .B2(n4789), .A(n4432), .ZN(n4434) );
  OAI21_X1 U5092 ( .B1(n4436), .B2(n4435), .A(n4434), .ZN(n4557) );
  INV_X1 U5093 ( .A(n4557), .ZN(n4444) );
  INV_X1 U5094 ( .A(n4436), .ZN(n4558) );
  NOR2_X1 U5095 ( .A1(n2194), .A2(n4437), .ZN(n4438) );
  AOI22_X1 U5096 ( .A1(n4806), .A2(REG2_REG_13__SCAN_IN), .B1(n4439), .B2(
        n4810), .ZN(n4440) );
  OAI21_X1 U5097 ( .B1(n4633), .B2(n4441), .A(n4440), .ZN(n4442) );
  AOI21_X1 U5098 ( .B1(n4558), .B2(n4811), .A(n4442), .ZN(n4443) );
  OAI21_X1 U5099 ( .B1(n4444), .B2(n4806), .A(n4443), .ZN(U3277) );
  NAND2_X1 U5100 ( .A1(n4578), .A2(n4898), .ZN(n4446) );
  NAND2_X1 U5101 ( .A1(n4895), .A2(REG1_REG_31__SCAN_IN), .ZN(n4445) );
  OAI211_X1 U5102 ( .C1(n4580), .C2(n4561), .A(n4446), .B(n4445), .ZN(U3549)
         );
  INV_X1 U5103 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4455) );
  INV_X1 U5104 ( .A(n3883), .ZN(n4449) );
  INV_X1 U5105 ( .A(n4447), .ZN(n4448) );
  NAND2_X1 U5106 ( .A1(n4670), .A2(n4888), .ZN(n4454) );
  OAI21_X1 U5107 ( .B1(n4452), .B2(n4563), .A(n4451), .ZN(n4669) );
  NAND2_X1 U5108 ( .A1(n4669), .A2(n4898), .ZN(n4453) );
  OAI211_X1 U5109 ( .C1(n4898), .C2(n4455), .A(n4454), .B(n4453), .ZN(U3548)
         );
  NOR2_X1 U5110 ( .A1(n4456), .A2(n4563), .ZN(n4457) );
  AOI21_X1 U5111 ( .B1(n4473), .B2(n4549), .A(n4457), .ZN(n4460) );
  NAND2_X1 U5112 ( .A1(n4458), .A2(n4792), .ZN(n4459) );
  MUX2_X1 U5113 ( .A(REG1_REG_27__SCAN_IN), .B(n4583), .S(n4898), .Z(U3545) );
  OAI22_X1 U5114 ( .A1(n4481), .A2(n4796), .B1(n4464), .B2(n4563), .ZN(n4465)
         );
  AOI21_X1 U5115 ( .B1(n4792), .B2(n4466), .A(n4465), .ZN(n4468) );
  OAI211_X1 U5116 ( .C1(n4469), .C2(n4536), .A(n4468), .B(n4467), .ZN(n4584)
         );
  MUX2_X1 U5117 ( .A(REG1_REG_26__SCAN_IN), .B(n4584), .S(n4898), .Z(n4470) );
  INV_X1 U5118 ( .A(n4470), .ZN(n4471) );
  OAI21_X1 U5119 ( .B1(n4561), .B2(n4587), .A(n4471), .ZN(U3544) );
  AOI22_X1 U5120 ( .A1(n4473), .A2(n4792), .B1(n4791), .B2(n4472), .ZN(n4474)
         );
  OAI211_X1 U5121 ( .C1(n4476), .C2(n4796), .A(n4475), .B(n4474), .ZN(n4477)
         );
  AOI21_X1 U5122 ( .B1(n4478), .B2(n4873), .A(n4477), .ZN(n4588) );
  MUX2_X1 U5123 ( .A(n4034), .B(n4588), .S(n4898), .Z(n4479) );
  OAI21_X1 U5124 ( .B1(n4561), .B2(n4591), .A(n4479), .ZN(U3543) );
  OAI22_X1 U5125 ( .A1(n4481), .A2(n4547), .B1(n4563), .B2(n4480), .ZN(n4482)
         );
  AOI21_X1 U5126 ( .B1(n4549), .B2(n4483), .A(n4482), .ZN(n4485) );
  OAI211_X1 U5127 ( .C1(n4486), .C2(n4536), .A(n4485), .B(n4484), .ZN(n4592)
         );
  MUX2_X1 U5128 ( .A(REG1_REG_24__SCAN_IN), .B(n4592), .S(n4898), .Z(n4487) );
  AOI21_X1 U5129 ( .B1(n4888), .B2(n4594), .A(n4487), .ZN(n4488) );
  INV_X1 U5130 ( .A(n4488), .ZN(U3542) );
  AOI22_X1 U5131 ( .A1(n4490), .A2(n4792), .B1(n4791), .B2(n4489), .ZN(n4491)
         );
  OAI211_X1 U5132 ( .C1(n4502), .C2(n4796), .A(n4492), .B(n4491), .ZN(n4493)
         );
  AOI21_X1 U5133 ( .B1(n4494), .B2(n4873), .A(n4493), .ZN(n4596) );
  MUX2_X1 U5134 ( .A(n4022), .B(n4596), .S(n4898), .Z(n4495) );
  OAI21_X1 U5135 ( .B1(n4561), .B2(n4599), .A(n4495), .ZN(U3541) );
  NAND3_X1 U5136 ( .A1(n4497), .A2(n4532), .A3(n4496), .ZN(n4498) );
  OAI211_X1 U5137 ( .C1(n4500), .C2(n4536), .A(n4499), .B(n4498), .ZN(n4600)
         );
  MUX2_X1 U5138 ( .A(REG1_REG_22__SCAN_IN), .B(n4600), .S(n4898), .Z(U3540) );
  OAI22_X1 U5139 ( .A1(n4502), .A2(n4547), .B1(n4563), .B2(n4501), .ZN(n4503)
         );
  AOI21_X1 U5140 ( .B1(n4549), .B2(n4504), .A(n4503), .ZN(n4506) );
  OAI211_X1 U5141 ( .C1(n4507), .C2(n4536), .A(n4506), .B(n4505), .ZN(n4602)
         );
  MUX2_X1 U5142 ( .A(REG1_REG_21__SCAN_IN), .B(n4602), .S(n4898), .Z(n4508) );
  AOI21_X1 U5143 ( .B1(n4888), .B2(n4601), .A(n4508), .ZN(n4509) );
  INV_X1 U5144 ( .A(n4509), .ZN(U3539) );
  INV_X1 U5145 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4512) );
  AOI21_X1 U5146 ( .B1(n4883), .B2(n4511), .A(n4510), .ZN(n4607) );
  MUX2_X1 U5147 ( .A(n4512), .B(n4607), .S(n4898), .Z(n4513) );
  OAI21_X1 U5148 ( .B1(n4561), .B2(n4610), .A(n4513), .ZN(U3538) );
  INV_X1 U5149 ( .A(n4514), .ZN(n4515) );
  AOI21_X1 U5150 ( .B1(n4516), .B2(n4873), .A(n4515), .ZN(n4611) );
  MUX2_X1 U5151 ( .A(n3915), .B(n4611), .S(n4898), .Z(n4517) );
  OAI21_X1 U5152 ( .B1(n4561), .B2(n4614), .A(n4517), .ZN(U3537) );
  OAI211_X1 U5153 ( .C1(n4520), .C2(n4536), .A(n4519), .B(n4518), .ZN(n4615)
         );
  MUX2_X1 U5154 ( .A(REG1_REG_18__SCAN_IN), .B(n4615), .S(n4898), .Z(U3536) );
  AOI22_X1 U5155 ( .A1(n4522), .A2(n4792), .B1(n4791), .B2(n4521), .ZN(n4523)
         );
  OAI211_X1 U5156 ( .C1(n4525), .C2(n4796), .A(n4524), .B(n4523), .ZN(n4526)
         );
  AOI21_X1 U5157 ( .B1(n4527), .B2(n4873), .A(n4526), .ZN(n4616) );
  MUX2_X1 U5158 ( .A(n3949), .B(n4616), .S(n4898), .Z(n4528) );
  OAI21_X1 U5159 ( .B1(n4561), .B2(n4619), .A(n4528), .ZN(U3535) );
  AOI22_X1 U5160 ( .A1(n4529), .A2(n4792), .B1(n4657), .B2(n4791), .ZN(n4530)
         );
  OAI21_X1 U5161 ( .B1(n4652), .B2(n4796), .A(n4530), .ZN(n4531) );
  AOI21_X1 U5162 ( .B1(n4533), .B2(n4532), .A(n4531), .ZN(n4535) );
  OAI211_X1 U5163 ( .C1(n4537), .C2(n4536), .A(n4535), .B(n4534), .ZN(n4620)
         );
  MUX2_X1 U5164 ( .A(REG1_REG_16__SCAN_IN), .B(n4620), .S(n4898), .Z(U3534) );
  AOI22_X1 U5165 ( .A1(n4539), .A2(n4792), .B1(n4791), .B2(n4538), .ZN(n4540)
         );
  OAI211_X1 U5166 ( .C1(n4542), .C2(n4796), .A(n4541), .B(n4540), .ZN(n4543)
         );
  AOI21_X1 U5167 ( .B1(n4544), .B2(n4873), .A(n4543), .ZN(n4621) );
  MUX2_X1 U5168 ( .A(n3868), .B(n4621), .S(n4898), .Z(n4545) );
  OAI21_X1 U5169 ( .B1(n4561), .B2(n4624), .A(n4545), .ZN(U3533) );
  INV_X1 U5170 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4555) );
  OAI22_X1 U5171 ( .A1(n4652), .A2(n4547), .B1(n4563), .B2(n4546), .ZN(n4548)
         );
  AOI21_X1 U5172 ( .B1(n4549), .B2(n4566), .A(n4548), .ZN(n4550) );
  OAI21_X1 U5173 ( .B1(n4552), .B2(n4551), .A(n4550), .ZN(n4553) );
  AOI21_X1 U5174 ( .B1(n4554), .B2(n4873), .A(n4553), .ZN(n4625) );
  MUX2_X1 U5175 ( .A(n4555), .B(n4625), .S(n4898), .Z(n4556) );
  OAI21_X1 U5176 ( .B1(n4561), .B2(n4628), .A(n4556), .ZN(U3532) );
  AOI21_X1 U5177 ( .B1(n4883), .B2(n4558), .A(n4557), .ZN(n4629) );
  MUX2_X1 U5178 ( .A(n4559), .B(n4629), .S(n4898), .Z(n4560) );
  OAI21_X1 U5179 ( .B1(n4561), .B2(n4633), .A(n4560), .ZN(U3531) );
  NAND2_X1 U5180 ( .A1(n4562), .A2(n4873), .ZN(n4573) );
  NOR2_X1 U5181 ( .A1(n4564), .A2(n4563), .ZN(n4565) );
  AOI21_X1 U5182 ( .B1(n4566), .B2(n4792), .A(n4565), .ZN(n4567) );
  OAI21_X1 U5183 ( .B1(n4568), .B2(n4796), .A(n4567), .ZN(n4569) );
  INV_X1 U5184 ( .A(n4569), .ZN(n4570) );
  AND2_X1 U5185 ( .A1(n4571), .A2(n4570), .ZN(n4572) );
  NAND2_X1 U5186 ( .A1(n4573), .A2(n4572), .ZN(n4634) );
  MUX2_X1 U5187 ( .A(REG1_REG_12__SCAN_IN), .B(n4634), .S(n4898), .Z(n4574) );
  AOI21_X1 U5188 ( .B1(n4888), .B2(n4636), .A(n4574), .ZN(n4575) );
  INV_X1 U5189 ( .A(n4575), .ZN(U3530) );
  NOR2_X1 U5190 ( .A1(n4886), .A2(n4576), .ZN(n4577) );
  AOI21_X1 U5191 ( .B1(n4578), .B2(n4886), .A(n4577), .ZN(n4579) );
  OAI21_X1 U5192 ( .B1(n4580), .B2(n4632), .A(n4579), .ZN(U3517) );
  NAND2_X1 U5193 ( .A1(n4670), .A2(n4865), .ZN(n4582) );
  NAND2_X1 U5194 ( .A1(n4669), .A2(n4886), .ZN(n4581) );
  OAI211_X1 U5195 ( .C1(n4886), .C2(n2691), .A(n4582), .B(n4581), .ZN(U3516)
         );
  MUX2_X1 U5196 ( .A(REG0_REG_27__SCAN_IN), .B(n4583), .S(n4886), .Z(U3513) );
  MUX2_X1 U5197 ( .A(REG0_REG_26__SCAN_IN), .B(n4584), .S(n4886), .Z(n4585) );
  INV_X1 U5198 ( .A(n4585), .ZN(n4586) );
  OAI21_X1 U5199 ( .B1(n4587), .B2(n4632), .A(n4586), .ZN(U3512) );
  MUX2_X1 U5200 ( .A(n4589), .B(n4588), .S(n4886), .Z(n4590) );
  OAI21_X1 U5201 ( .B1(n4591), .B2(n4632), .A(n4590), .ZN(U3511) );
  MUX2_X1 U5202 ( .A(REG0_REG_24__SCAN_IN), .B(n4592), .S(n4886), .Z(n4593) );
  AOI21_X1 U5203 ( .B1(n4594), .B2(n4865), .A(n4593), .ZN(n4595) );
  INV_X1 U5204 ( .A(n4595), .ZN(U3510) );
  MUX2_X1 U5205 ( .A(n4597), .B(n4596), .S(n4886), .Z(n4598) );
  OAI21_X1 U5206 ( .B1(n4599), .B2(n4632), .A(n4598), .ZN(U3509) );
  MUX2_X1 U5207 ( .A(REG0_REG_22__SCAN_IN), .B(n4600), .S(n4886), .Z(U3508) );
  INV_X1 U5208 ( .A(n4601), .ZN(n4606) );
  INV_X1 U5209 ( .A(n4602), .ZN(n4603) );
  MUX2_X1 U5210 ( .A(n4604), .B(n4603), .S(n4886), .Z(n4605) );
  OAI21_X1 U5211 ( .B1(n4606), .B2(n4632), .A(n4605), .ZN(U3507) );
  MUX2_X1 U5212 ( .A(n4608), .B(n4607), .S(n4886), .Z(n4609) );
  OAI21_X1 U5213 ( .B1(n4610), .B2(n4632), .A(n4609), .ZN(U3506) );
  MUX2_X1 U5214 ( .A(n4612), .B(n4611), .S(n4886), .Z(n4613) );
  OAI21_X1 U5215 ( .B1(n4614), .B2(n4632), .A(n4613), .ZN(U3505) );
  MUX2_X1 U5216 ( .A(REG0_REG_18__SCAN_IN), .B(n4615), .S(n4886), .Z(U3503) );
  MUX2_X1 U5217 ( .A(n4617), .B(n4616), .S(n4886), .Z(n4618) );
  OAI21_X1 U5218 ( .B1(n4619), .B2(n4632), .A(n4618), .ZN(U3501) );
  MUX2_X1 U5219 ( .A(REG0_REG_16__SCAN_IN), .B(n4620), .S(n4886), .Z(U3499) );
  MUX2_X1 U5220 ( .A(n4622), .B(n4621), .S(n4886), .Z(n4623) );
  OAI21_X1 U5221 ( .B1(n4624), .B2(n4632), .A(n4623), .ZN(U3497) );
  MUX2_X1 U5222 ( .A(n4626), .B(n4625), .S(n4886), .Z(n4627) );
  OAI21_X1 U5223 ( .B1(n4628), .B2(n4632), .A(n4627), .ZN(U3495) );
  MUX2_X1 U5224 ( .A(n4630), .B(n4629), .S(n4886), .Z(n4631) );
  OAI21_X1 U5225 ( .B1(n4633), .B2(n4632), .A(n4631), .ZN(U3493) );
  MUX2_X1 U5226 ( .A(REG0_REG_12__SCAN_IN), .B(n4634), .S(n4886), .Z(n4635) );
  AOI21_X1 U5227 ( .B1(n4636), .B2(n4865), .A(n4635), .ZN(n4637) );
  INV_X1 U5228 ( .A(n4637), .ZN(U3491) );
  MUX2_X1 U5229 ( .A(n4638), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5230 ( .A(n4639), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5231 ( .A(DATAI_20_), .B(n4640), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5232 ( .A(n4641), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  MUX2_X1 U5233 ( .A(n4642), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5234 ( .A(n4643), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5235 ( .A(n4644), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5236 ( .A(DATAI_4_), .B(n4645), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5237 ( .A(n4646), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5238 ( .A(n2161), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5239 ( .A(n4648), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U5240 ( .A1(STATE_REG_SCAN_IN), .A2(n4650), .B1(n4649), .B2(U3149), 
        .ZN(U3324) );
  NOR2_X1 U5241 ( .A1(STATE_REG_SCAN_IN), .A2(n4651), .ZN(n4748) );
  OAI22_X1 U5242 ( .A1(n4654), .A2(n3659), .B1(n4653), .B2(n4652), .ZN(n4655)
         );
  AOI211_X1 U5243 ( .C1(n4657), .C2(n4656), .A(n4748), .B(n4655), .ZN(n4666)
         );
  INV_X1 U5244 ( .A(n4658), .ZN(n4660) );
  OAI21_X1 U5245 ( .B1(n4660), .B2(n4659), .A(n3657), .ZN(n4662) );
  XNOR2_X1 U5246 ( .A(n4662), .B(n4661), .ZN(n4664) );
  NAND2_X1 U5247 ( .A1(n4664), .A2(n4663), .ZN(n4665) );
  OAI211_X1 U5248 ( .C1(n4668), .C2(n4667), .A(n4666), .B(n4665), .ZN(U3223)
         );
  AOI22_X1 U5249 ( .A1(n4670), .A2(n4802), .B1(n4815), .B2(n4669), .ZN(n4671)
         );
  OAI21_X1 U5250 ( .B1(n4672), .B2(n4815), .A(n4671), .ZN(U3261) );
  AOI211_X1 U5251 ( .C1(n3118), .C2(n4674), .A(n4673), .B(n4754), .ZN(n4676)
         );
  AOI211_X1 U5252 ( .C1(n4767), .C2(ADDR_REG_8__SCAN_IN), .A(n4676), .B(n4675), 
        .ZN(n4680) );
  OAI211_X1 U5253 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4678), .A(n4771), .B(n4677), 
        .ZN(n4679) );
  OAI211_X1 U5254 ( .C1(n4775), .C2(n4855), .A(n4680), .B(n4679), .ZN(U3248)
         );
  AOI211_X1 U5255 ( .C1(n4683), .C2(n4682), .A(n4681), .B(n4754), .ZN(n4685)
         );
  AOI211_X1 U5256 ( .C1(n4767), .C2(ADDR_REG_9__SCAN_IN), .A(n4685), .B(n4684), 
        .ZN(n4690) );
  OAI211_X1 U5257 ( .C1(n4688), .C2(n4687), .A(n4771), .B(n4686), .ZN(n4689)
         );
  OAI211_X1 U5258 ( .C1(n4775), .C2(n4853), .A(n4690), .B(n4689), .ZN(U3249)
         );
  AOI211_X1 U5259 ( .C1(n3250), .C2(n4692), .A(n4691), .B(n4754), .ZN(n4694)
         );
  AOI211_X1 U5260 ( .C1(n4767), .C2(ADDR_REG_10__SCAN_IN), .A(n4694), .B(n4693), .ZN(n4698) );
  OAI211_X1 U5261 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4696), .A(n4771), .B(n4695), .ZN(n4697) );
  OAI211_X1 U5262 ( .C1(n4775), .C2(n4851), .A(n4698), .B(n4697), .ZN(U3250)
         );
  AOI211_X1 U5263 ( .C1(n2193), .C2(n4700), .A(n4699), .B(n4754), .ZN(n4702)
         );
  AOI211_X1 U5264 ( .C1(n4767), .C2(ADDR_REG_11__SCAN_IN), .A(n4702), .B(n4701), .ZN(n4707) );
  OAI211_X1 U5265 ( .C1(n4705), .C2(n4704), .A(n4771), .B(n4703), .ZN(n4706)
         );
  OAI211_X1 U5266 ( .C1(n4775), .C2(n4849), .A(n4707), .B(n4706), .ZN(U3251)
         );
  OAI21_X1 U5267 ( .B1(REG2_REG_13__SCAN_IN), .B2(n4709), .A(n4708), .ZN(n4711) );
  OAI21_X1 U5268 ( .B1(n2171), .B2(n4711), .A(n4762), .ZN(n4710) );
  AOI21_X1 U5269 ( .B1(n2171), .B2(n4711), .A(n4710), .ZN(n4713) );
  AOI211_X1 U5270 ( .C1(n4767), .C2(ADDR_REG_13__SCAN_IN), .A(n4713), .B(n4712), .ZN(n4718) );
  OAI211_X1 U5271 ( .C1(n4716), .C2(n4715), .A(n4771), .B(n4714), .ZN(n4717)
         );
  OAI211_X1 U5272 ( .C1(n4775), .C2(n4847), .A(n4718), .B(n4717), .ZN(U3253)
         );
  OAI211_X1 U5273 ( .C1(REG2_REG_14__SCAN_IN), .C2(n4721), .A(n4762), .B(n4720), .ZN(n4722) );
  NAND2_X1 U5274 ( .A1(n4723), .A2(n4722), .ZN(n4724) );
  AOI21_X1 U5275 ( .B1(ADDR_REG_14__SCAN_IN), .B2(n4767), .A(n4724), .ZN(n4728) );
  OAI211_X1 U5276 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4726), .A(n4771), .B(n4725), .ZN(n4727) );
  OAI211_X1 U5277 ( .C1(n4775), .C2(n3852), .A(n4728), .B(n4727), .ZN(U3254)
         );
  OAI211_X1 U5278 ( .C1(n4731), .C2(n4730), .A(n4771), .B(n4729), .ZN(n4736)
         );
  OAI211_X1 U5279 ( .C1(n4734), .C2(n4733), .A(n4762), .B(n4732), .ZN(n4735)
         );
  OAI211_X1 U5280 ( .C1(n4775), .C2(n4844), .A(n4736), .B(n4735), .ZN(n4737)
         );
  AOI211_X1 U5281 ( .C1(n4767), .C2(ADDR_REG_15__SCAN_IN), .A(n4738), .B(n4737), .ZN(n4739) );
  INV_X1 U5282 ( .A(n4739), .ZN(U3255) );
  INV_X1 U5283 ( .A(n4740), .ZN(n4842) );
  AOI21_X1 U5284 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4742), .A(n4741), .ZN(n4746) );
  AOI21_X1 U5285 ( .B1(REG2_REG_16__SCAN_IN), .B2(n4744), .A(n4743), .ZN(n4745) );
  OAI22_X1 U5286 ( .A1(n4746), .A2(n4756), .B1(n4745), .B2(n4754), .ZN(n4747)
         );
  AOI211_X1 U5287 ( .C1(n4767), .C2(ADDR_REG_16__SCAN_IN), .A(n4748), .B(n4747), .ZN(n4749) );
  OAI21_X1 U5288 ( .B1(n4842), .B2(n4775), .A(n4749), .ZN(U3256) );
  AOI21_X1 U5289 ( .B1(n2184), .B2(n4751), .A(n4750), .ZN(n4757) );
  AOI21_X1 U5290 ( .B1(n2182), .B2(n4753), .A(n4752), .ZN(n4755) );
  OAI22_X1 U5291 ( .A1(n4757), .A2(n4756), .B1(n4755), .B2(n4754), .ZN(n4758)
         );
  OAI21_X1 U5292 ( .B1(n4840), .B2(n4775), .A(n4760), .ZN(U3257) );
  OAI211_X1 U5293 ( .C1(n4764), .C2(n4763), .A(n4762), .B(n4761), .ZN(n4769)
         );
  INV_X1 U5294 ( .A(n4765), .ZN(n4766) );
  OAI211_X1 U5295 ( .C1(n4773), .C2(n4772), .A(n4771), .B(n4770), .ZN(n4774)
         );
  OAI211_X1 U5296 ( .C1(n4775), .C2(n4839), .A(n2310), .B(n4774), .ZN(U3258)
         );
  AOI22_X1 U5297 ( .A1(n4776), .A2(n4810), .B1(REG2_REG_6__SCAN_IN), .B2(n4806), .ZN(n4782) );
  INV_X1 U5298 ( .A(n4777), .ZN(n4780) );
  INV_X1 U5299 ( .A(n4778), .ZN(n4779) );
  AOI22_X1 U5300 ( .A1(n4780), .A2(n4811), .B1(n4802), .B2(n4779), .ZN(n4781)
         );
  OAI211_X1 U5301 ( .C1(n4806), .C2(n4783), .A(n4782), .B(n4781), .ZN(U3284)
         );
  XNOR2_X1 U5302 ( .A(n4785), .B(n4784), .ZN(n4864) );
  OAI21_X1 U5303 ( .B1(n4788), .B2(n4787), .A(n4786), .ZN(n4790) );
  NAND2_X1 U5304 ( .A1(n4790), .A2(n4789), .ZN(n4795) );
  AOI22_X1 U5305 ( .A1(n4793), .A2(n4792), .B1(n4791), .B2(n4801), .ZN(n4794)
         );
  OAI211_X1 U5306 ( .C1(n2374), .C2(n4796), .A(n4795), .B(n4794), .ZN(n4863)
         );
  AOI21_X1 U5307 ( .B1(n4797), .B2(n4864), .A(n4863), .ZN(n4805) );
  AOI22_X1 U5308 ( .A1(n4806), .A2(REG2_REG_3__SCAN_IN), .B1(n4810), .B2(n4798), .ZN(n4804) );
  AOI21_X1 U5309 ( .B1(n4801), .B2(n4800), .A(n4799), .ZN(n4889) );
  AOI22_X1 U5310 ( .A1(n4864), .A2(n4811), .B1(n4802), .B2(n4889), .ZN(n4803)
         );
  OAI211_X1 U5311 ( .C1(n4806), .C2(n4805), .A(n4804), .B(n4803), .ZN(U3287)
         );
  AOI21_X1 U5312 ( .B1(n4809), .B2(n4808), .A(n4807), .ZN(n4816) );
  AOI22_X1 U5313 ( .A1(n4812), .A2(n4811), .B1(REG3_REG_0__SCAN_IN), .B2(n4810), .ZN(n4813) );
  OAI221_X1 U5314 ( .B1(n4806), .B2(n4816), .C1(n4815), .C2(n4814), .A(n4813), 
        .ZN(U3290) );
  NOR2_X1 U5315 ( .A1(n4834), .A2(n4818), .ZN(U3291) );
  NOR2_X1 U5316 ( .A1(n4834), .A2(n4819), .ZN(U3292) );
  NOR2_X1 U5317 ( .A1(n4834), .A2(n4820), .ZN(U3293) );
  NOR2_X1 U5318 ( .A1(n4834), .A2(n4821), .ZN(U3294) );
  NOR2_X1 U5319 ( .A1(n4834), .A2(n4822), .ZN(U3295) );
  AND2_X1 U5320 ( .A1(D_REG_26__SCAN_IN), .A2(n4835), .ZN(U3296) );
  NOR2_X1 U5321 ( .A1(n4834), .A2(n4823), .ZN(U3297) );
  AND2_X1 U5322 ( .A1(D_REG_24__SCAN_IN), .A2(n4835), .ZN(U3298) );
  AND2_X1 U5323 ( .A1(D_REG_23__SCAN_IN), .A2(n4835), .ZN(U3299) );
  AND2_X1 U5324 ( .A1(D_REG_22__SCAN_IN), .A2(n4835), .ZN(U3300) );
  NOR2_X1 U5325 ( .A1(n4834), .A2(n4824), .ZN(U3301) );
  AND2_X1 U5326 ( .A1(D_REG_20__SCAN_IN), .A2(n4835), .ZN(U3302) );
  NOR2_X1 U5327 ( .A1(n4834), .A2(n4825), .ZN(U3303) );
  AND2_X1 U5328 ( .A1(D_REG_18__SCAN_IN), .A2(n4835), .ZN(U3304) );
  NOR2_X1 U5329 ( .A1(n4834), .A2(n4826), .ZN(U3305) );
  NOR2_X1 U5330 ( .A1(n4834), .A2(n4827), .ZN(U3306) );
  AND2_X1 U5331 ( .A1(D_REG_15__SCAN_IN), .A2(n4835), .ZN(U3307) );
  NOR2_X1 U5332 ( .A1(n4834), .A2(n4828), .ZN(U3308) );
  NOR2_X1 U5333 ( .A1(n4834), .A2(n4829), .ZN(U3309) );
  NOR2_X1 U5334 ( .A1(n4834), .A2(n4830), .ZN(U3310) );
  AND2_X1 U5335 ( .A1(D_REG_11__SCAN_IN), .A2(n4835), .ZN(U3311) );
  NOR2_X1 U5336 ( .A1(n4834), .A2(n4831), .ZN(U3312) );
  AND2_X1 U5337 ( .A1(D_REG_9__SCAN_IN), .A2(n4835), .ZN(U3313) );
  NOR2_X1 U5338 ( .A1(n4834), .A2(n4832), .ZN(U3314) );
  AND2_X1 U5339 ( .A1(D_REG_7__SCAN_IN), .A2(n4835), .ZN(U3315) );
  AND2_X1 U5340 ( .A1(D_REG_6__SCAN_IN), .A2(n4835), .ZN(U3316) );
  AND2_X1 U5341 ( .A1(D_REG_5__SCAN_IN), .A2(n4835), .ZN(U3317) );
  NOR2_X1 U5342 ( .A1(n4834), .A2(n4833), .ZN(U3318) );
  AND2_X1 U5343 ( .A1(D_REG_3__SCAN_IN), .A2(n4835), .ZN(U3319) );
  AND2_X1 U5344 ( .A1(D_REG_2__SCAN_IN), .A2(n4835), .ZN(U3320) );
  AOI21_X1 U5345 ( .B1(U3149), .B2(n4837), .A(n4836), .ZN(U3329) );
  AOI22_X1 U5346 ( .A1(STATE_REG_SCAN_IN), .A2(n4839), .B1(n4838), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5347 ( .A1(STATE_REG_SCAN_IN), .A2(n4840), .B1(n2545), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5348 ( .A1(STATE_REG_SCAN_IN), .A2(n4842), .B1(n4841), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5349 ( .A1(STATE_REG_SCAN_IN), .A2(n4844), .B1(n4843), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5350 ( .A(DATAI_14_), .ZN(n4845) );
  AOI22_X1 U5351 ( .A1(STATE_REG_SCAN_IN), .A2(n3852), .B1(n4845), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5352 ( .A(DATAI_13_), .ZN(n4846) );
  AOI22_X1 U5353 ( .A1(STATE_REG_SCAN_IN), .A2(n4847), .B1(n4846), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5354 ( .A(DATAI_11_), .ZN(n4848) );
  AOI22_X1 U5355 ( .A1(STATE_REG_SCAN_IN), .A2(n4849), .B1(n4848), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5356 ( .A(DATAI_10_), .ZN(n4850) );
  AOI22_X1 U5357 ( .A1(STATE_REG_SCAN_IN), .A2(n4851), .B1(n4850), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5358 ( .A(DATAI_9_), .ZN(n4852) );
  AOI22_X1 U5359 ( .A1(STATE_REG_SCAN_IN), .A2(n4853), .B1(n4852), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5360 ( .A1(STATE_REG_SCAN_IN), .A2(n4855), .B1(n4854), .B2(U3149), 
        .ZN(U3344) );
  AOI22_X1 U5361 ( .A1(STATE_REG_SCAN_IN), .A2(n2270), .B1(n4856), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5362 ( .A1(n4886), .A2(n4857), .B1(n2358), .B2(n4885), .ZN(U3467)
         );
  OAI22_X1 U5363 ( .A1(n4860), .A2(n4859), .B1(n4878), .B2(n4858), .ZN(n4861)
         );
  NOR2_X1 U5364 ( .A1(n4862), .A2(n4861), .ZN(n4887) );
  AOI22_X1 U5365 ( .A1(n4886), .A2(n4887), .B1(n2346), .B2(n4885), .ZN(U3469)
         );
  AOI21_X1 U5366 ( .B1(n4873), .B2(n4864), .A(n4863), .ZN(n4891) );
  AOI22_X1 U5367 ( .A1(n4889), .A2(n4865), .B1(REG0_REG_3__SCAN_IN), .B2(n4885), .ZN(n4866) );
  OAI21_X1 U5368 ( .B1(n4891), .B2(n4885), .A(n4866), .ZN(U3473) );
  INV_X1 U5369 ( .A(n4867), .ZN(n4871) );
  INV_X1 U5370 ( .A(n4868), .ZN(n4870) );
  AOI211_X1 U5371 ( .C1(n4871), .C2(n4883), .A(n4870), .B(n4869), .ZN(n4893)
         );
  AOI22_X1 U5372 ( .A1(n4886), .A2(n4893), .B1(n2395), .B2(n4885), .ZN(U3475)
         );
  AND3_X1 U5373 ( .A1(n4874), .A2(n4873), .A3(n4872), .ZN(n4875) );
  NOR3_X1 U5374 ( .A1(n4877), .A2(n4876), .A3(n4875), .ZN(n4894) );
  AOI22_X1 U5375 ( .A1(n4886), .A2(n4894), .B1(n2437), .B2(n4885), .ZN(U3481)
         );
  NOR3_X1 U5376 ( .A1(n4880), .A2(n4879), .A3(n4878), .ZN(n4882) );
  AOI211_X1 U5377 ( .C1(n4884), .C2(n4883), .A(n4882), .B(n4881), .ZN(n4897)
         );
  AOI22_X1 U5378 ( .A1(n4886), .A2(n4897), .B1(n2429), .B2(n4885), .ZN(U3483)
         );
  AOI22_X1 U5379 ( .A1(n4898), .A2(n4887), .B1(n2794), .B2(n4895), .ZN(U3519)
         );
  AOI22_X1 U5380 ( .A1(n4889), .A2(n4888), .B1(REG1_REG_3__SCAN_IN), .B2(n4895), .ZN(n4890) );
  OAI21_X1 U5381 ( .B1(n4891), .B2(n4895), .A(n4890), .ZN(U3521) );
  AOI22_X1 U5382 ( .A1(n4898), .A2(n4893), .B1(n4892), .B2(n4895), .ZN(U3522)
         );
  AOI22_X1 U5383 ( .A1(n4898), .A2(n4894), .B1(n3202), .B2(n4895), .ZN(U3525)
         );
  INV_X1 U5384 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4896) );
  AOI22_X1 U5385 ( .A1(n4898), .A2(n4897), .B1(n4896), .B2(n4895), .ZN(U3526)
         );
  INV_X2 U3008 ( .A(n4815), .ZN(n4806) );
  CLKBUF_X1 U2401 ( .A(n2359), .Z(n2885) );
endmodule

