

module b15_C_SARLock_k_64_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744;

  NAND2_X1 U3438 ( .A1(n3306), .A2(n3305), .ZN(n3307) );
  BUF_X1 U3439 ( .A(n3587), .Z(n3621) );
  CLKBUF_X2 U3440 ( .A(n2997), .Z(n3989) );
  NOR2_X1 U3441 ( .A1(n4280), .A2(n3629), .ZN(n3625) );
  CLKBUF_X2 U3442 ( .A(n4175), .Z(n4144) );
  CLKBUF_X2 U3443 ( .A(n3094), .Z(n3856) );
  CLKBUF_X2 U3444 ( .A(n3207), .Z(n4173) );
  CLKBUF_X2 U34450 ( .A(n3088), .Z(n4151) );
  CLKBUF_X2 U34460 ( .A(n3161), .Z(n4057) );
  CLKBUF_X2 U34470 ( .A(n3294), .Z(n2992) );
  CLKBUF_X2 U34480 ( .A(n3162), .Z(n2999) );
  INV_X2 U3449 ( .A(n3202), .ZN(n4096) );
  CLKBUF_X2 U3450 ( .A(n3149), .Z(n4174) );
  CLKBUF_X2 U34510 ( .A(n3089), .Z(n3988) );
  OR2_X1 U34530 ( .A1(n3085), .A2(n3084), .ZN(n3515) );
  CLKBUF_X1 U3454 ( .A(n3117), .Z(n3510) );
  AND2_X1 U34550 ( .A1(n3025), .A2(n4397), .ZN(n4175) );
  AND2_X2 U34560 ( .A1(n4294), .A2(n4377), .ZN(n3010) );
  AND2_X2 U3457 ( .A1(n4333), .A2(n4397), .ZN(n3149) );
  AND2_X2 U3458 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4397) );
  AND2_X2 U34590 ( .A1(n4286), .A2(n3019), .ZN(n2997) );
  NAND3_X1 U34600 ( .A1(n4256), .A2(n4322), .A3(n3190), .ZN(n4280) );
  NAND2_X1 U34610 ( .A1(n3515), .A2(n3648), .ZN(n3587) );
  NAND2_X2 U34620 ( .A1(n3648), .A2(n6065), .ZN(n4324) );
  OR2_X1 U34630 ( .A1(n5294), .A2(n5334), .ZN(n5427) );
  AND2_X1 U34640 ( .A1(n5987), .A2(n4998), .ZN(n5999) );
  INV_X1 U34650 ( .A(n6001), .ZN(n5955) );
  INV_X1 U3466 ( .A(n5999), .ZN(n6037) );
  XNOR2_X1 U3467 ( .A(n3624), .B(n3623), .ZN(n5355) );
  AND2_X2 U34680 ( .A1(n3642), .A2(n3116), .ZN(n3137) );
  AND2_X1 U34690 ( .A1(n4291), .A2(n4377), .ZN(n2989) );
  AND2_X1 U34700 ( .A1(n4291), .A2(n4377), .ZN(n2990) );
  NAND2_X2 U34720 ( .A1(n4341), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3233) );
  OAI21_X2 U34730 ( .B1(n4942), .B2(n3447), .A(n3182), .ZN(n4341) );
  AND2_X2 U34740 ( .A1(n3016), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4337) );
  NAND2_X2 U3475 ( .A1(n4225), .A2(n4224), .ZN(n4226) );
  NOR2_X2 U3476 ( .A1(n5545), .A2(n3652), .ZN(n5527) );
  AND2_X1 U3477 ( .A1(n5855), .A2(n5856), .ZN(n3419) );
  CLKBUF_X1 U3478 ( .A(n5457), .Z(n5465) );
  OR2_X1 U3479 ( .A1(n5494), .A2(n5487), .ZN(n5488) );
  AND2_X1 U3480 ( .A1(n5486), .A2(n5485), .ZN(n5494) );
  CLKBUF_X1 U3481 ( .A(n5291), .Z(n5332) );
  NAND2_X1 U3482 ( .A1(n5304), .A2(n5303), .ZN(n5484) );
  NAND2_X1 U3483 ( .A1(n3968), .A2(n3967), .ZN(n5293) );
  CLKBUF_X1 U3484 ( .A(n5273), .Z(n5300) );
  NAND2_X1 U3485 ( .A1(n5402), .A2(n3621), .ZN(n5398) );
  CLKBUF_X1 U3486 ( .A(n5068), .Z(n5069) );
  AND2_X1 U3487 ( .A1(n5256), .A2(n3408), .ZN(n5614) );
  INV_X1 U3488 ( .A(n5576), .ZN(n4227) );
  AOI21_X1 U3489 ( .B1(n3725), .B2(n3932), .A(n3724), .ZN(n4442) );
  NAND2_X1 U3490 ( .A1(n3369), .A2(n3368), .ZN(n3391) );
  OR2_X1 U3491 ( .A1(n3701), .A2(n3700), .ZN(n4410) );
  NAND2_X1 U3492 ( .A1(n3682), .A2(n3920), .ZN(n3701) );
  CLKBUF_X1 U3493 ( .A(n4433), .Z(n4736) );
  CLKBUF_X2 U3494 ( .A(n3704), .Z(n6539) );
  OR2_X1 U3495 ( .A1(n3273), .A2(n3272), .ZN(n3274) );
  AND2_X1 U3496 ( .A1(n5138), .A2(n5221), .ZN(n5250) );
  NAND2_X1 U3497 ( .A1(n3302), .A2(n3301), .ZN(n4519) );
  CLKBUF_X1 U3498 ( .A(n3284), .Z(n4389) );
  NAND2_X1 U3499 ( .A1(n3245), .A2(n3244), .ZN(n3284) );
  NAND2_X1 U3500 ( .A1(n3216), .A2(n3215), .ZN(n3267) );
  NAND2_X1 U3501 ( .A1(n3174), .A2(n3175), .ZN(n3178) );
  CLKBUF_X1 U3502 ( .A(n4332), .Z(n5359) );
  AND2_X1 U3503 ( .A1(n3236), .A2(n3238), .ZN(n3201) );
  NAND2_X1 U3504 ( .A1(n3532), .A2(n3007), .ZN(n4419) );
  AND3_X1 U3505 ( .A1(n3136), .A2(n3135), .A3(n3134), .ZN(n3138) );
  NAND2_X1 U3506 ( .A1(n3177), .A2(n3176), .ZN(n3217) );
  AND2_X1 U3507 ( .A1(n3185), .A2(n3184), .ZN(n3502) );
  NAND2_X1 U3508 ( .A1(n3172), .A2(n3171), .ZN(n3176) );
  CLKBUF_X1 U3509 ( .A(n3485), .Z(n4308) );
  AOI21_X1 U3510 ( .B1(n3131), .B2(n3508), .A(n3130), .ZN(n3631) );
  CLKBUF_X1 U3511 ( .A(n3118), .Z(n4360) );
  NAND2_X1 U3512 ( .A1(n3491), .A2(n3132), .ZN(n3508) );
  INV_X1 U3513 ( .A(n4324), .ZN(n4366) );
  BUF_X2 U3514 ( .A(n3587), .Z(n5478) );
  CLKBUF_X1 U3515 ( .A(n3189), .Z(n3190) );
  OR2_X1 U3516 ( .A1(n3168), .A2(n3167), .ZN(n3392) );
  INV_X1 U3517 ( .A(n3112), .ZN(n3189) );
  INV_X1 U3518 ( .A(n6065), .ZN(n3180) );
  BUF_X2 U3519 ( .A(n3112), .Z(n3491) );
  OR2_X2 U3520 ( .A1(n3110), .A2(n3109), .ZN(n3648) );
  OR2_X1 U3521 ( .A1(n3061), .A2(n3060), .ZN(n3635) );
  BUF_X2 U3522 ( .A(n4145), .Z(n4172) );
  BUF_X2 U3523 ( .A(n3995), .Z(n2991) );
  AND2_X1 U3524 ( .A1(n3025), .A2(n4397), .ZN(n2998) );
  BUF_X2 U3525 ( .A(n3208), .Z(n3156) );
  INV_X2 U3526 ( .A(n6570), .ZN(n6556) );
  CLKBUF_X1 U3527 ( .A(n4897), .Z(n6536) );
  AND2_X1 U3528 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4286) );
  AND2_X1 U3529 ( .A1(n5449), .A2(n5547), .ZN(n2993) );
  AND2_X1 U3530 ( .A1(n5458), .A2(n5547), .ZN(n5448) );
  AND2_X1 U3531 ( .A1(n3025), .A2(n3026), .ZN(n2994) );
  AND2_X2 U3532 ( .A1(n3025), .A2(n3026), .ZN(n4145) );
  AND2_X1 U3533 ( .A1(n4333), .A2(n4397), .ZN(n2995) );
  AND2_X2 U3534 ( .A1(n4333), .A2(n3026), .ZN(n3089) );
  AND2_X2 U3535 ( .A1(n3026), .A2(n4377), .ZN(n3208) );
  AND2_X2 U3536 ( .A1(n3026), .A2(n4377), .ZN(n3001) );
  NAND2_X1 U3537 ( .A1(n3273), .A2(n3272), .ZN(n3310) );
  XNOR2_X1 U3538 ( .A(n3266), .B(n3265), .ZN(n3273) );
  NAND2_X1 U3539 ( .A1(n3183), .A2(n4256), .ZN(n3642) );
  NAND2_X1 U3540 ( .A1(n3502), .A2(n4510), .ZN(n4303) );
  NAND2_X1 U3541 ( .A1(n3003), .A2(n3011), .ZN(n3117) );
  AND2_X1 U3542 ( .A1(n4397), .A2(n4377), .ZN(n2996) );
  AND2_X2 U3543 ( .A1(n4397), .A2(n4377), .ZN(n3162) );
  AND2_X4 U3544 ( .A1(n4337), .A2(n3026), .ZN(n3051) );
  AND2_X2 U3545 ( .A1(n4337), .A2(n4291), .ZN(n3088) );
  NAND2_X1 U3546 ( .A1(n3497), .A2(n5503), .ZN(n3688) );
  AND2_X4 U3547 ( .A1(n4294), .A2(n4333), .ZN(n3094) );
  AND2_X2 U3548 ( .A1(n5457), .A2(n4095), .ZN(n5458) );
  NAND2_X2 U3549 ( .A1(n4408), .A2(n4437), .ZN(n4443) );
  NAND2_X2 U3550 ( .A1(n3703), .A2(n3702), .ZN(n4408) );
  INV_X1 U3551 ( .A(n3962), .ZN(n5302) );
  XNOR2_X2 U3552 ( .A(n3962), .B(n5301), .ZN(n5273) );
  AND2_X1 U3553 ( .A1(n3026), .A2(n4377), .ZN(n3000) );
  NAND2_X2 U3554 ( .A1(n3237), .A2(n3143), .ZN(n3690) );
  NAND2_X2 U3555 ( .A1(n3139), .A2(n3140), .ZN(n3237) );
  INV_X1 U3556 ( .A(n3263), .ZN(n3276) );
  INV_X1 U3557 ( .A(n3608), .ZN(n3603) );
  AND2_X1 U3558 ( .A1(n3651), .A2(n3650), .ZN(n4298) );
  NAND2_X1 U3559 ( .A1(n6557), .A2(n4198), .ZN(n5987) );
  OR2_X2 U3560 ( .A1(n3072), .A2(n3071), .ZN(n5503) );
  OR3_X1 U3561 ( .A1(n5731), .A2(READY_N), .A3(n4309), .ZN(n6140) );
  AND2_X1 U3562 ( .A1(n3132), .A2(n3635), .ZN(n3073) );
  AND2_X1 U3563 ( .A1(n3367), .A2(n3366), .ZN(n3370) );
  NAND2_X1 U3564 ( .A1(n3497), .A2(n3112), .ZN(n3118) );
  OR2_X1 U3565 ( .A1(n3259), .A2(n3258), .ZN(n3263) );
  NOR2_X1 U3566 ( .A1(n3220), .A2(n3219), .ZN(n3221) );
  INV_X1 U3567 ( .A(n3217), .ZN(n3220) );
  INV_X1 U3568 ( .A(n3471), .ZN(n3354) );
  OR2_X1 U3569 ( .A1(n3300), .A2(n3299), .ZN(n3304) );
  AOI22_X1 U3570 ( .A1(n3094), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3105) );
  OR2_X1 U3571 ( .A1(n3344), .A2(n3343), .ZN(n3345) );
  OR2_X1 U3572 ( .A1(n4349), .A2(n6562), .ZN(n4162) );
  INV_X1 U3573 ( .A(n3952), .ZN(n4165) );
  INV_X1 U3574 ( .A(n4788), .ZN(n3740) );
  NOR2_X1 U3575 ( .A1(n3681), .A2(n6560), .ZN(n3932) );
  CLKBUF_X1 U3576 ( .A(n3952), .Z(n4188) );
  INV_X1 U3577 ( .A(n3932), .ZN(n3956) );
  NAND2_X1 U3578 ( .A1(n3530), .A2(n3529), .ZN(n4413) );
  NAND2_X1 U3579 ( .A1(n3526), .A2(n3525), .ZN(n3530) );
  NAND2_X1 U3580 ( .A1(n3118), .A2(n3515), .ZN(n3129) );
  AND2_X1 U3581 ( .A1(n3115), .A2(n4281), .ZN(n3116) );
  NAND2_X1 U3582 ( .A1(n3496), .A2(n3014), .ZN(n3115) );
  NAND2_X1 U3583 ( .A1(n3144), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3471) );
  INV_X1 U3584 ( .A(n3289), .ZN(n3144) );
  INV_X1 U3585 ( .A(n6026), .ZN(n6009) );
  INV_X1 U3586 ( .A(n3920), .ZN(n4191) );
  NOR2_X1 U3587 ( .A1(n4140), .A2(n5540), .ZN(n4141) );
  NOR2_X2 U3588 ( .A1(n5411), .A2(n5413), .ZN(n5412) );
  INV_X1 U3589 ( .A(n5460), .ZN(n4095) );
  NAND2_X1 U3590 ( .A1(n3735), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3742)
         );
  NOR2_X2 U3591 ( .A1(n5429), .A2(n4230), .ZN(n5469) );
  NOR2_X2 U3592 ( .A1(n5438), .A2(n5439), .ZN(n5499) );
  AND2_X1 U3593 ( .A1(n3655), .A2(n3647), .ZN(n5215) );
  OR2_X1 U3594 ( .A1(n5708), .A2(n3404), .ZN(n5201) );
  NAND2_X1 U3595 ( .A1(n3549), .A2(n3548), .ZN(n5030) );
  INV_X1 U3596 ( .A(n4498), .ZN(n3549) );
  NOR2_X2 U3597 ( .A1(n4419), .A2(n4420), .ZN(n4500) );
  INV_X1 U3598 ( .A(n6192), .ZN(n5592) );
  XNOR2_X1 U3599 ( .A(n4389), .B(n4936), .ZN(n4279) );
  CLKBUF_X1 U3600 ( .A(n4374), .Z(n4375) );
  OR3_X1 U3601 ( .A1(n4314), .A2(n4358), .A3(n4313), .ZN(n4391) );
  OR2_X1 U3602 ( .A1(n6540), .A2(n5154), .ZN(n4895) );
  INV_X1 U3603 ( .A(n4610), .ZN(n4612) );
  INV_X1 U3604 ( .A(n4523), .ZN(n4893) );
  NOR2_X1 U3605 ( .A1(n4728), .A2(n4518), .ZN(n4455) );
  OR2_X1 U3606 ( .A1(n3441), .A2(n3440), .ZN(n3443) );
  AND2_X1 U3607 ( .A1(n4997), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4998) );
  AND2_X1 U3608 ( .A1(n5987), .A2(n4201), .ZN(n6001) );
  AND2_X1 U3609 ( .A1(n5505), .A2(n5504), .ZN(n6062) );
  OAI21_X1 U3610 ( .B1(n3690), .B2(STATE2_REG_0__SCAN_IN), .A(n3176), .ZN(
        n3174) );
  CLKBUF_X1 U3611 ( .A(n4279), .Z(n6540) );
  INV_X1 U3612 ( .A(n4856), .ZN(n4883) );
  INV_X1 U3613 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3018) );
  NAND2_X1 U3614 ( .A1(n3603), .A2(n3524), .ZN(n3526) );
  NAND2_X1 U3615 ( .A1(n3120), .A2(n3119), .ZN(n3126) );
  AND2_X1 U3616 ( .A1(n3132), .A2(n3392), .ZN(n3173) );
  AND2_X1 U3617 ( .A1(n3129), .A2(n5503), .ZN(n3086) );
  AND2_X1 U3618 ( .A1(n5299), .A2(n3963), .ZN(n3961) );
  AND2_X2 U3619 ( .A1(n4337), .A2(n4397), .ZN(n3294) );
  AND2_X1 U3620 ( .A1(n3958), .A2(n5342), .ZN(n5306) );
  INV_X1 U3621 ( .A(n5227), .ZN(n3820) );
  AND2_X1 U3622 ( .A1(n3719), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3727)
         );
  INV_X1 U3623 ( .A(n5584), .ZN(n4224) );
  INV_X1 U3624 ( .A(n3371), .ZN(n3369) );
  OR2_X1 U3625 ( .A1(n5236), .A2(n3406), .ZN(n5239) );
  OAI22_X1 U3626 ( .A1(n3714), .A2(n3447), .B1(n3328), .B2(n4249), .ZN(n3329)
         );
  INV_X1 U3627 ( .A(n3173), .ZN(n3389) );
  NAND2_X1 U3628 ( .A1(n3271), .A2(n3270), .ZN(n3272) );
  XNOR2_X1 U3629 ( .A(n3267), .B(n3225), .ZN(n4429) );
  NAND2_X1 U3630 ( .A1(n3114), .A2(n3113), .ZN(n4281) );
  INV_X1 U3631 ( .A(n3587), .ZN(n3113) );
  INV_X1 U3632 ( .A(n3508), .ZN(n3114) );
  INV_X1 U3633 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4642) );
  AOI21_X1 U3634 ( .B1(n6450), .B2(n5732), .A(n5387), .ZN(n4453) );
  OR2_X1 U3635 ( .A1(n5731), .A2(n4261), .ZN(n4251) );
  CLKBUF_X1 U3636 ( .A(n3502), .Z(n4259) );
  OAI211_X1 U3637 ( .C1(n3870), .C2(n3734), .A(n3733), .B(n3732), .ZN(n4554)
         );
  AND2_X1 U3638 ( .A1(n5738), .A2(n4188), .ZN(n4137) );
  AND2_X1 U3639 ( .A1(n4120), .A2(n4119), .ZN(n5547) );
  AND2_X1 U3640 ( .A1(n4072), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4073)
         );
  NAND2_X1 U3641 ( .A1(n4073), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4113)
         );
  NOR2_X1 U3642 ( .A1(n4033), .A2(n5579), .ZN(n4034) );
  AND2_X1 U3643 ( .A1(n4034), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4072)
         );
  CLKBUF_X1 U3644 ( .A(n5422), .Z(n5423) );
  INV_X1 U3645 ( .A(n5331), .ZN(n4007) );
  AND2_X1 U3646 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3983), .ZN(n3984)
         );
  NAND2_X1 U3647 ( .A1(n3984), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4033)
         );
  NAND2_X1 U3648 ( .A1(n3854), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3982)
         );
  AND2_X1 U3649 ( .A1(n3918), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3903)
         );
  AND2_X1 U3650 ( .A1(n3949), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3918)
         );
  OR2_X1 U3651 ( .A1(n5576), .A2(n5898), .ZN(n5616) );
  NOR2_X1 U3652 ( .A1(n6621), .A2(n3948), .ZN(n3949) );
  INV_X1 U3653 ( .A(n3742), .ZN(n3743) );
  AOI21_X1 U3654 ( .B1(n3739), .B2(n3932), .A(n3738), .ZN(n4788) );
  NAND2_X1 U3655 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3706) );
  CLKBUF_X1 U3656 ( .A(n5315), .Z(n5316) );
  AND2_X1 U3657 ( .A1(n3572), .A2(n3571), .ZN(n5266) );
  NAND2_X1 U3658 ( .A1(n5250), .A2(n3569), .ZN(n5267) );
  CLKBUF_X1 U3659 ( .A(n5208), .Z(n5209) );
  AND2_X1 U3660 ( .A1(n3558), .A2(n3557), .ZN(n5109) );
  AND2_X1 U3661 ( .A1(n3552), .A2(n3551), .ZN(n5029) );
  AND2_X1 U3662 ( .A1(n3547), .A2(n3546), .ZN(n5013) );
  AND2_X1 U3663 ( .A1(n3537), .A2(n3536), .ZN(n4420) );
  INV_X1 U3664 ( .A(n4412), .ZN(n3532) );
  AND2_X1 U3665 ( .A1(n3649), .A2(n5248), .ZN(n5214) );
  NAND2_X1 U3666 ( .A1(n3655), .A2(n4298), .ZN(n5698) );
  AND2_X1 U3667 ( .A1(n3631), .A2(n3133), .ZN(n3134) );
  INV_X1 U3668 ( .A(n3175), .ZN(n3177) );
  CLKBUF_X1 U3669 ( .A(n4429), .Z(n4735) );
  INV_X1 U3670 ( .A(n5359), .ZN(n4575) );
  INV_X1 U3671 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4347) );
  INV_X1 U3672 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3024) );
  OR2_X1 U3673 ( .A1(n6339), .A2(n4735), .ZN(n4648) );
  AND2_X1 U3674 ( .A1(n5155), .A2(n6540), .ZN(n6341) );
  NAND2_X1 U3675 ( .A1(n6539), .A2(n4736), .ZN(n6339) );
  OR3_X1 U3676 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4453), .A3(n6718), .ZN(n4511) );
  NOR2_X1 U3677 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4453), .ZN(n4523) );
  INV_X1 U3678 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5059) );
  OR2_X1 U3679 ( .A1(n4996), .A2(n4204), .ZN(n6026) );
  OR2_X1 U3680 ( .A1(n4996), .A2(n4995), .ZN(n6004) );
  INV_X1 U3681 ( .A(n6045), .ZN(n5501) );
  AND2_X1 U3682 ( .A1(n6045), .A2(n5376), .ZN(n6040) );
  AND2_X2 U3683 ( .A1(n4327), .A2(n6436), .ZN(n6045) );
  INV_X1 U3684 ( .A(n6040), .ZN(n5817) );
  NAND2_X1 U3685 ( .A1(n4359), .A2(n6140), .ZN(n5505) );
  NOR2_X1 U3687 ( .A1(n6091), .A2(n6103), .ZN(n6102) );
  OR2_X1 U3688 ( .A1(n4199), .A2(n5522), .ZN(n4200) );
  INV_X1 U3689 ( .A(n4192), .ZN(n4193) );
  INV_X1 U3690 ( .A(n5393), .ZN(n5394) );
  INV_X1 U3691 ( .A(n5465), .ZN(n5459) );
  INV_X1 U3692 ( .A(n6200), .ZN(n6186) );
  INV_X1 U3693 ( .A(n5873), .ZN(n6197) );
  AND2_X1 U3694 ( .A1(n5404), .A2(n5403), .ZN(n5628) );
  CLKBUF_X1 U3695 ( .A(n5198), .Z(n5199) );
  INV_X1 U3696 ( .A(n5698), .ZN(n6241) );
  INV_X1 U3697 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6408) );
  INV_X1 U3698 ( .A(n6542), .ZN(n6545) );
  INV_X1 U3699 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4339) );
  INV_X1 U3700 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5389) );
  NOR2_X1 U3701 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5902) );
  INV_X1 U3702 ( .A(n4631), .ZN(n4599) );
  OAI21_X1 U3703 ( .B1(n4899), .B2(n4894), .A(n5166), .ZN(n4927) );
  AND2_X1 U3704 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6299), .ZN(n6327)
         );
  INV_X1 U3705 ( .A(n6300), .ZN(n6328) );
  OR2_X1 U3706 ( .A1(n6294), .A2(n4807), .ZN(n6300) );
  OR2_X1 U3707 ( .A1(n4859), .A2(n4858), .ZN(n4888) );
  NAND2_X1 U3708 ( .A1(n4455), .A2(n4942), .ZN(n4885) );
  AOI21_X1 U3709 ( .B1(n3484), .B2(n3483), .A(n3482), .ZN(n6407) );
  NOR2_X1 U3710 ( .A1(n3481), .A2(n3480), .ZN(n3482) );
  NAND2_X1 U3711 ( .A1(n3473), .A2(n3472), .ZN(n3484) );
  INV_X1 U3712 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6441) );
  NOR2_X1 U3713 ( .A1(n5881), .A2(n3012), .ZN(n4236) );
  XOR2_X1 U3714 ( .A(n5528), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .Z(n3002) );
  AND4_X1 U3715 ( .A1(n3023), .A2(n3022), .A3(n3021), .A4(n3020), .ZN(n3003)
         );
  NOR2_X2 U3716 ( .A1(n5648), .A2(n5647), .ZN(n5451) );
  NAND2_X2 U3717 ( .A1(n3391), .A2(n3390), .ZN(n5576) );
  OR2_X1 U3718 ( .A1(n4318), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3004)
         );
  NAND2_X1 U3719 ( .A1(n5708), .A2(n5112), .ZN(n3005) );
  OR2_X1 U3720 ( .A1(n5576), .A2(n3415), .ZN(n3006) );
  INV_X1 U3721 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5142) );
  AND2_X1 U3722 ( .A1(n3531), .A2(n4413), .ZN(n3007) );
  NAND2_X1 U3723 ( .A1(n5108), .A2(n3560), .ZN(n3561) );
  INV_X1 U3724 ( .A(n3561), .ZN(n5138) );
  NAND2_X1 U3725 ( .A1(n5576), .A2(n5898), .ZN(n3008) );
  NOR2_X1 U3726 ( .A1(n5708), .A2(n5265), .ZN(n3009) );
  NAND2_X1 U3727 ( .A1(n3655), .A2(n3512), .ZN(n5717) );
  AND4_X1 U3728 ( .A1(n3030), .A2(n3029), .A3(n3028), .A4(n3027), .ZN(n3011)
         );
  INV_X1 U3729 ( .A(n3683), .ZN(n3870) );
  NAND2_X1 U3730 ( .A1(n3327), .A2(n3326), .ZN(n3714) );
  AND2_X1 U3731 ( .A1(n4235), .A2(n4234), .ZN(n3012) );
  AND2_X1 U3732 ( .A1(n3679), .A2(n3678), .ZN(n3013) );
  AND2_X1 U3733 ( .A1(n4510), .A2(n6065), .ZN(n3014) );
  INV_X1 U3734 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U3735 ( .A1(n5708), .A2(n3659), .ZN(n3015) );
  AND2_X1 U3737 ( .A1(n5902), .A2(n6443), .ZN(n6238) );
  NAND2_X1 U3738 ( .A1(n4360), .A2(n3510), .ZN(n3119) );
  INV_X1 U3739 ( .A(n3218), .ZN(n3219) );
  AOI22_X1 U3740 ( .A1(n4145), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3020) );
  NOR2_X1 U3741 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3019) );
  AND2_X1 U3742 ( .A1(n3323), .A2(n3322), .ZN(n3324) );
  AOI22_X1 U3743 ( .A1(n3088), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3042) );
  AOI21_X1 U3744 ( .B1(n3285), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3243), 
        .ZN(n3246) );
  NAND2_X1 U3745 ( .A1(n6065), .A2(n3510), .ZN(n3289) );
  INV_X1 U3746 ( .A(EBX_REG_2__SCAN_IN), .ZN(n3524) );
  OR2_X1 U3747 ( .A1(n5747), .A2(n4165), .ZN(n4119) );
  AND2_X1 U3748 ( .A1(n3008), .A2(n5614), .ZN(n3409) );
  INV_X1 U3749 ( .A(n5140), .ZN(n3560) );
  OR2_X1 U3750 ( .A1(n3364), .A2(n3363), .ZN(n3381) );
  OR2_X1 U3751 ( .A1(n3214), .A2(n3213), .ZN(n3226) );
  NAND2_X1 U3752 ( .A1(n3289), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3475) );
  OR2_X1 U3753 ( .A1(n3471), .A2(n4590), .ZN(n3172) );
  OR3_X1 U3754 ( .A1(n3441), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6419), 
        .ZN(n3436) );
  OR2_X1 U3755 ( .A1(n4324), .A2(EBX_REG_1__SCAN_IN), .ZN(n3516) );
  AND2_X1 U3756 ( .A1(n3960), .A2(n5305), .ZN(n3963) );
  OR2_X1 U3757 ( .A1(n3850), .A2(n5284), .ZN(n3948) );
  INV_X1 U3758 ( .A(n5011), .ZN(n3748) );
  OAI211_X1 U3759 ( .C1(n3118), .C2(n3510), .A(n5503), .B(n4321), .ZN(n3630)
         );
  AND2_X1 U3760 ( .A1(n5708), .A2(n6612), .ZN(n3418) );
  INV_X1 U3761 ( .A(n3370), .ZN(n3368) );
  OR2_X1 U3762 ( .A1(n3341), .A2(n3340), .ZN(n3348) );
  OR2_X1 U3763 ( .A1(n3155), .A2(n3154), .ZN(n3227) );
  OR2_X1 U3764 ( .A1(n3199), .A2(n3198), .ZN(n3236) );
  NAND2_X1 U3765 ( .A1(n3142), .A2(n3141), .ZN(n3143) );
  AND2_X1 U3766 ( .A1(n3187), .A2(n3186), .ZN(n3485) );
  NOR2_X1 U3767 ( .A1(n6026), .A2(n5960), .ZN(n5950) );
  AND2_X1 U3768 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3705), .ZN(n3719)
         );
  INV_X1 U3769 ( .A(n3870), .ZN(n4187) );
  NOR2_X1 U3770 ( .A1(n5012), .A2(n5013), .ZN(n3548) );
  INV_X1 U3771 ( .A(n3714), .ZN(n3725) );
  NAND2_X1 U3772 ( .A1(n2993), .A2(n5458), .ZN(n5411) );
  AND2_X1 U3773 ( .A1(n3957), .A2(n5483), .ZN(n5342) );
  OR2_X1 U3774 ( .A1(n5239), .A2(n3009), .ZN(n5613) );
  NAND2_X1 U3775 ( .A1(n3801), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3805)
         );
  XNOR2_X1 U3776 ( .A(n3391), .B(n3379), .ZN(n3747) );
  OR2_X1 U3777 ( .A1(n5576), .A2(n3413), .ZN(n3414) );
  OR2_X1 U3778 ( .A1(n3406), .A2(n5237), .ZN(n5240) );
  OR2_X1 U3779 ( .A1(n5083), .A2(n3399), .ZN(n3401) );
  NAND2_X1 U3780 ( .A1(n4500), .A2(n4499), .ZN(n4498) );
  NAND2_X1 U3781 ( .A1(n3281), .A2(n3280), .ZN(n6182) );
  AND2_X1 U3782 ( .A1(n4643), .A2(n4897), .ZN(n4645) );
  NAND2_X1 U3783 ( .A1(n3288), .A2(n3287), .ZN(n4936) );
  OR2_X1 U3784 ( .A1(n3471), .A2(n3447), .ZN(n3481) );
  NAND2_X1 U3785 ( .A1(n3180), .A2(n3648), .ZN(n3634) );
  AND2_X1 U3786 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n4114), .ZN(n4115)
         );
  INV_X1 U3787 ( .A(n3982), .ZN(n3983) );
  NOR2_X1 U3788 ( .A1(n3805), .A2(n5142), .ZN(n3822) );
  NOR2_X1 U3789 ( .A1(n3777), .A2(n5076), .ZN(n3801) );
  AND2_X1 U3790 ( .A1(n3727), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3735)
         );
  NAND2_X1 U3791 ( .A1(n5987), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4996) );
  OR2_X1 U3792 ( .A1(n4996), .A2(n5354), .ZN(n4216) );
  AND2_X1 U3793 ( .A1(n3959), .A2(n5306), .ZN(n5305) );
  OR2_X1 U3794 ( .A1(n5436), .A2(n5437), .ZN(n5493) );
  OR2_X1 U3795 ( .A1(n3726), .A2(n3956), .ZN(n3733) );
  AND2_X1 U3796 ( .A1(n4414), .A2(n4415), .ZN(n3700) );
  XNOR2_X1 U3797 ( .A(n4200), .B(n4209), .ZN(n4997) );
  NOR2_X1 U3798 ( .A1(n3902), .A2(n3851), .ZN(n3854) );
  OR2_X1 U3799 ( .A1(n3764), .A2(n5059), .ZN(n3777) );
  AOI21_X1 U3800 ( .B1(n3747), .B2(n3932), .A(n3746), .ZN(n5011) );
  NAND2_X1 U3801 ( .A1(n4217), .A2(n6240), .ZN(n3679) );
  BUF_X1 U3802 ( .A(n5517), .Z(n5555) );
  AND2_X1 U3803 ( .A1(n3407), .A2(n5240), .ZN(n5256) );
  OAI21_X1 U3804 ( .B1(n3726), .B2(n3447), .A(n3350), .ZN(n3351) );
  NAND2_X1 U3805 ( .A1(n4363), .A2(n3235), .ZN(n6183) );
  NAND2_X1 U3806 ( .A1(n3491), .A2(n3648), .ZN(n3447) );
  INV_X1 U3807 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3016) );
  INV_X1 U3808 ( .A(n6540), .ZN(n6254) );
  OR3_X1 U3809 ( .A1(n6539), .A2(n4574), .A3(n4735), .ZN(n4610) );
  OR2_X1 U3810 ( .A1(n6539), .A2(n4737), .ZN(n6571) );
  XNOR2_X1 U3811 ( .A(n3310), .B(n4519), .ZN(n3704) );
  OR2_X1 U3812 ( .A1(n6294), .A2(n4735), .ZN(n4943) );
  INV_X1 U3813 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4769) );
  OR2_X1 U3814 ( .A1(n4648), .A2(n4942), .ZN(n5159) );
  OR2_X1 U3815 ( .A1(n4728), .A2(n4735), .ZN(n4778) );
  AND2_X1 U3816 ( .A1(n6441), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3506) );
  NAND2_X1 U3817 ( .A1(n4115), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4140)
         );
  NAND2_X1 U3818 ( .A1(n3903), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3902)
         );
  AND2_X1 U3819 ( .A1(n5987), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U3820 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n3743), .ZN(n3764)
         );
  INV_X1 U3821 ( .A(n5994), .ZN(n6022) );
  INV_X1 U3822 ( .A(n6004), .ZN(n6028) );
  NAND2_X1 U3823 ( .A1(n5467), .A2(n5461), .ZN(n5648) );
  OR2_X1 U3824 ( .A1(n5427), .A2(n5426), .ZN(n5429) );
  NAND2_X1 U3825 ( .A1(n5496), .A2(n5320), .ZN(n5339) );
  OR2_X1 U3826 ( .A1(n5267), .A2(n5266), .ZN(n5438) );
  AND2_X1 U3827 ( .A1(n6045), .A2(n5503), .ZN(n6041) );
  AND2_X1 U3828 ( .A1(n5505), .A2(n5378), .ZN(n6052) );
  INV_X1 U3829 ( .A(n5505), .ZN(n6061) );
  AND2_X1 U3830 ( .A1(n5505), .A2(n4362), .ZN(n5514) );
  INV_X1 U3831 ( .A(n6105), .ZN(n6091) );
  INV_X1 U3832 ( .A(n6115), .ZN(n6178) );
  AND2_X1 U3833 ( .A1(n5411), .A2(n5450), .ZN(n5823) );
  INV_X1 U3834 ( .A(n5806), .ZN(n5862) );
  AND2_X1 U3835 ( .A1(n5489), .A2(n5488), .ZN(n6054) );
  AND2_X1 U3836 ( .A1(n5436), .A2(n5346), .ZN(n5968) );
  INV_X1 U3837 ( .A(n6191), .ZN(n5868) );
  OR2_X1 U3838 ( .A1(n6407), .A2(n6445), .ZN(n5731) );
  MUX2_X1 U3839 ( .A(n5526), .B(n5527), .S(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .Z(n5519) );
  INV_X1 U3840 ( .A(n4226), .ZN(n5583) );
  INV_X1 U3841 ( .A(n5717), .ZN(n6245) );
  AND2_X1 U3842 ( .A1(n3655), .A2(n3627), .ZN(n6240) );
  AND2_X1 U3843 ( .A1(n3507), .A2(n6436), .ZN(n3655) );
  NOR2_X1 U3844 ( .A1(n6407), .A2(n6718), .ZN(n5387) );
  INV_X1 U3845 ( .A(n6571), .ZN(n4932) );
  INV_X1 U3846 ( .A(n4953), .ZN(n4986) );
  INV_X1 U3847 ( .A(n6287), .ZN(n6329) );
  OR2_X1 U3848 ( .A1(n4693), .A2(n4692), .ZN(n4721) );
  INV_X1 U3849 ( .A(n4942), .ZN(n4777) );
  INV_X1 U3850 ( .A(n5159), .ZN(n5192) );
  OR2_X1 U3851 ( .A1(n4812), .A2(n4811), .ZN(n4849) );
  NOR2_X1 U3852 ( .A1(n4778), .A2(n4942), .ZN(n4856) );
  INV_X1 U3853 ( .A(n6259), .ZN(n6290) );
  AND2_X1 U3854 ( .A1(n3506), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6436) );
  INV_X1 U3855 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6562) );
  AND2_X1 U3856 ( .A1(n4251), .A2(n4252), .ZN(n6557) );
  INV_X1 U3857 ( .A(n5993), .ZN(n6018) );
  INV_X1 U3858 ( .A(n6007), .ZN(n6031) );
  INV_X1 U3859 ( .A(n6033), .ZN(n5367) );
  OR2_X1 U3860 ( .A1(n5495), .A2(n5494), .ZN(n6059) );
  INV_X1 U3861 ( .A(n5278), .ZN(n5327) );
  INV_X1 U3862 ( .A(n5514), .ZN(n5329) );
  OR3_X1 U3863 ( .A1(n5731), .A2(n5730), .A3(n6461), .ZN(n6105) );
  INV_X1 U3864 ( .A(n6110), .ZN(n6115) );
  NAND2_X1 U3865 ( .A1(n6193), .A2(n4240), .ZN(n5873) );
  NAND2_X1 U3866 ( .A1(n5873), .A2(n6196), .ZN(n6191) );
  NOR2_X1 U3867 ( .A1(n4232), .A2(n4236), .ZN(n4237) );
  INV_X1 U3868 ( .A(n6238), .ZN(n6192) );
  INV_X1 U3869 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6544) );
  AND2_X1 U3870 ( .A1(n4581), .A2(n4580), .ZN(n4638) );
  NAND2_X1 U3871 ( .A1(n4612), .A2(n4777), .ZN(n4935) );
  OR3_X1 U3872 ( .A1(n6539), .A2(n4518), .A3(n4517), .ZN(n6575) );
  INV_X1 U3873 ( .A(n4952), .ZN(n4989) );
  OR2_X1 U3874 ( .A1(n6294), .A2(n6253), .ZN(n6287) );
  OR2_X1 U3875 ( .A1(n4648), .A2(n4777), .ZN(n4727) );
  AOI21_X1 U3876 ( .B1(n5164), .B2(n6341), .A(n5158), .ZN(n5194) );
  OR2_X1 U3877 ( .A1(n6339), .A2(n6253), .ZN(n6399) );
  OR2_X1 U3878 ( .A1(n6339), .A2(n4807), .ZN(n6388) );
  INV_X1 U3879 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6463) );
  NOR2_X4 U3880 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3026) );
  INV_X1 U3881 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3017) );
  NOR2_X2 U3882 ( .A1(n3017), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4291)
         );
  NOR2_X4 U3883 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4333) );
  AND2_X2 U3884 ( .A1(n4291), .A2(n4333), .ZN(n3161) );
  AOI22_X1 U3885 ( .A1(n3051), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3161), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3023) );
  NOR2_X2 U3886 ( .A1(n3018), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3025)
         );
  AOI22_X1 U3887 ( .A1(n3088), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3022) );
  AOI22_X1 U3888 ( .A1(n3149), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3021) );
  AND2_X4 U3889 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4377) );
  NOR2_X2 U3890 ( .A1(n3024), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4294)
         );
  AND2_X2 U3891 ( .A1(n4291), .A2(n3025), .ZN(n3995) );
  AOI22_X1 U3892 ( .A1(n3094), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3030) );
  AOI22_X1 U3893 ( .A1(n3010), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3029) );
  AOI22_X1 U3894 ( .A1(n3294), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3028) );
  AND2_X2 U3895 ( .A1(n4294), .A2(n4337), .ZN(n3207) );
  AOI22_X1 U3896 ( .A1(n3207), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3027) );
  INV_X2 U3897 ( .A(n3117), .ZN(n3132) );
  AOI22_X1 U3898 ( .A1(n3094), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3010), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3034) );
  AOI22_X1 U3899 ( .A1(n3051), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3033) );
  AOI22_X1 U3900 ( .A1(n3995), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3032) );
  AOI22_X1 U3901 ( .A1(n3253), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3031) );
  NAND4_X1 U3902 ( .A1(n3034), .A2(n3033), .A3(n3032), .A4(n3031), .ZN(n3040)
         );
  AOI22_X1 U3903 ( .A1(n3088), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3038) );
  AOI22_X1 U3904 ( .A1(n3207), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n2995), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3037) );
  AOI22_X1 U3905 ( .A1(n3001), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3036) );
  AOI22_X1 U3906 ( .A1(n3161), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3035) );
  NAND4_X1 U3907 ( .A1(n3038), .A2(n3037), .A3(n3036), .A4(n3035), .ZN(n3039)
         );
  OR2_X2 U3908 ( .A1(n3040), .A2(n3039), .ZN(n3681) );
  AOI22_X1 U3909 ( .A1(n3051), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3044) );
  AOI22_X1 U3910 ( .A1(n3161), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3043) );
  AOI22_X1 U3911 ( .A1(n4145), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3041) );
  NAND4_X1 U3912 ( .A1(n3044), .A2(n3043), .A3(n3042), .A4(n3041), .ZN(n3050)
         );
  AOI22_X1 U3913 ( .A1(n3010), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3048) );
  AOI22_X1 U3914 ( .A1(n3294), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3047) );
  AOI22_X1 U3915 ( .A1(n3207), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3046) );
  AOI22_X1 U3916 ( .A1(n3094), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3045) );
  NAND4_X1 U3917 ( .A1(n3048), .A2(n3047), .A3(n3046), .A4(n3045), .ZN(n3049)
         );
  OR2_X2 U3918 ( .A1(n3050), .A2(n3049), .ZN(n3112) );
  OAI21_X1 U3920 ( .B1(n3132), .B2(n3681), .A(n4321), .ZN(n3062) );
  AOI22_X1 U3921 ( .A1(n3088), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3055) );
  AOI22_X1 U3922 ( .A1(n4145), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3054) );
  AOI22_X1 U3923 ( .A1(n3051), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U3924 ( .A1(n3161), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3052) );
  NAND4_X1 U3925 ( .A1(n3055), .A2(n3054), .A3(n3053), .A4(n3052), .ZN(n3061)
         );
  AOI22_X1 U3926 ( .A1(n3010), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3059) );
  AOI22_X1 U3927 ( .A1(n3294), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3058) );
  AOI22_X1 U3928 ( .A1(n3207), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U3929 ( .A1(n3094), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3056) );
  NAND4_X1 U3930 ( .A1(n3059), .A2(n3058), .A3(n3057), .A4(n3056), .ZN(n3060)
         );
  NAND2_X1 U3931 ( .A1(n3062), .A2(n4454), .ZN(n3075) );
  INV_X2 U3932 ( .A(n3681), .ZN(n3497) );
  AOI22_X1 U3933 ( .A1(n3088), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3066) );
  AOI22_X1 U3934 ( .A1(n4145), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3065) );
  AOI22_X1 U3935 ( .A1(n3051), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U3936 ( .A1(n3161), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3063) );
  NAND4_X1 U3937 ( .A1(n3066), .A2(n3065), .A3(n3064), .A4(n3063), .ZN(n3072)
         );
  AOI22_X1 U3938 ( .A1(n3010), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3070) );
  AOI22_X1 U3939 ( .A1(n3294), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U3940 ( .A1(n3207), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3068) );
  AOI22_X1 U3941 ( .A1(n3094), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3067) );
  NAND4_X1 U3942 ( .A1(n3070), .A2(n3069), .A3(n3068), .A4(n3067), .ZN(n3071)
         );
  NAND3_X1 U3943 ( .A1(n3073), .A2(n3688), .A3(n4321), .ZN(n3074) );
  NAND2_X1 U3944 ( .A1(n3075), .A2(n3074), .ZN(n3087) );
  AOI22_X1 U3945 ( .A1(n3088), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3079) );
  AOI22_X1 U3946 ( .A1(n2994), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3078) );
  AOI22_X1 U3947 ( .A1(n3051), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3077) );
  AOI22_X1 U3948 ( .A1(n3161), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3076) );
  NAND4_X1 U3949 ( .A1(n3079), .A2(n3078), .A3(n3077), .A4(n3076), .ZN(n3085)
         );
  AOI22_X1 U3950 ( .A1(n3010), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3083) );
  AOI22_X1 U3951 ( .A1(n3294), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3082) );
  AOI22_X1 U3952 ( .A1(n3207), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3081) );
  AOI22_X1 U3953 ( .A1(n3094), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3080) );
  NAND4_X1 U3954 ( .A1(n3083), .A2(n3082), .A3(n3081), .A4(n3080), .ZN(n3084)
         );
  NAND2_X1 U3955 ( .A1(n3087), .A2(n3086), .ZN(n3183) );
  AOI22_X1 U3956 ( .A1(n3207), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3051), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3093) );
  AOI22_X1 U3957 ( .A1(n3088), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3092) );
  AOI22_X1 U3958 ( .A1(n3010), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3091) );
  AOI22_X1 U3959 ( .A1(n3161), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3090) );
  NAND4_X1 U3960 ( .A1(n3093), .A2(n3092), .A3(n3091), .A4(n3090), .ZN(n3100)
         );
  AOI22_X1 U3961 ( .A1(n3294), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3098) );
  AOI22_X1 U3962 ( .A1(n3094), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3097) );
  AOI22_X1 U3963 ( .A1(n3995), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3096) );
  AOI22_X1 U3964 ( .A1(n3253), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3095) );
  NAND4_X1 U3965 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3099)
         );
  OR2_X4 U3966 ( .A1(n3100), .A2(n3099), .ZN(n6065) );
  AOI22_X1 U3967 ( .A1(n3088), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3995), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3104) );
  AOI22_X1 U3968 ( .A1(n4145), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4175), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3103) );
  AOI22_X1 U3969 ( .A1(n3051), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3149), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3102) );
  AOI22_X1 U3970 ( .A1(n3161), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3101) );
  NAND4_X1 U3971 ( .A1(n3104), .A2(n3103), .A3(n3102), .A4(n3101), .ZN(n3110)
         );
  AOI22_X1 U3972 ( .A1(n3010), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n2990), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U3973 ( .A1(n3294), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3089), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3107) );
  AOI22_X1 U3974 ( .A1(n3207), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3106) );
  NAND4_X1 U3975 ( .A1(n3108), .A2(n3107), .A3(n3106), .A4(n3105), .ZN(n3109)
         );
  NOR2_X2 U3976 ( .A1(n6065), .A2(n3648), .ZN(n4256) );
  AND2_X1 U3977 ( .A1(n3132), .A2(n5503), .ZN(n3111) );
  NAND2_X1 U3978 ( .A1(n3111), .A2(n4321), .ZN(n3496) );
  INV_X2 U3979 ( .A(n3648), .ZN(n4510) );
  INV_X1 U3980 ( .A(n3630), .ZN(n3120) );
  INV_X1 U3981 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6455) );
  NOR2_X1 U3982 ( .A1(n6463), .A2(n6455), .ZN(n6469) );
  NOR2_X1 U3983 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n3121) );
  NOR2_X1 U3984 ( .A1(n6469), .A2(n3121), .ZN(n3423) );
  NOR2_X1 U3985 ( .A1(n3648), .A2(n3423), .ZN(n3188) );
  INV_X2 U3986 ( .A(n3635), .ZN(n4454) );
  NAND2_X1 U3987 ( .A1(n4454), .A2(n3515), .ZN(n3637) );
  INV_X1 U3988 ( .A(n3637), .ZN(n3228) );
  OAI211_X1 U3989 ( .C1(n3188), .C2(n3491), .A(n3228), .B(n3634), .ZN(n3122)
         );
  NOR2_X1 U3990 ( .A1(n3126), .A2(n3122), .ZN(n3123) );
  NAND2_X1 U3991 ( .A1(n3137), .A2(n3123), .ZN(n3124) );
  NAND2_X1 U3992 ( .A1(n3124), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U3993 ( .A1(n5902), .A2(n6562), .ZN(n4239) );
  MUX2_X1 U3994 ( .A(n4239), .B(n3506), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3125) );
  OAI21_X2 U3995 ( .B1(n3240), .B2(n4347), .A(n3125), .ZN(n3139) );
  INV_X1 U3996 ( .A(n3126), .ZN(n3127) );
  NAND2_X1 U3997 ( .A1(n3127), .A2(n3515), .ZN(n3128) );
  NAND2_X1 U3998 ( .A1(n3128), .A2(n3648), .ZN(n3136) );
  AND2_X1 U3999 ( .A1(n4510), .A2(n6065), .ZN(n3179) );
  NAND2_X1 U4000 ( .A1(n5902), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6444) );
  AOI21_X1 U4001 ( .B1(n3129), .B2(n3179), .A(n6444), .ZN(n3135) );
  INV_X1 U4002 ( .A(n3634), .ZN(n3131) );
  AND2_X1 U4003 ( .A1(n6065), .A2(n3635), .ZN(n3130) );
  NOR2_X1 U4004 ( .A1(n3688), .A2(n3132), .ZN(n3492) );
  NOR2_X2 U4005 ( .A1(n3635), .A2(n3515), .ZN(n4322) );
  NAND2_X1 U4006 ( .A1(n3492), .A2(n4322), .ZN(n3133) );
  NAND2_X1 U4007 ( .A1(n3138), .A2(n3137), .ZN(n3140) );
  INV_X1 U4008 ( .A(n3139), .ZN(n3142) );
  INV_X1 U4009 ( .A(n3140), .ZN(n3141) );
  INV_X1 U4010 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4590) );
  AOI22_X1 U4011 ( .A1(n4173), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4012 ( .A1(n4151), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4013 ( .A1(n4096), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4014 ( .A1(n3051), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3145) );
  NAND4_X1 U4015 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n3155)
         );
  AOI22_X1 U4016 ( .A1(n2991), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4017 ( .A1(n3856), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4018 ( .A1(n4057), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4019 ( .A1(n2992), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3150) );
  NAND4_X1 U4020 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n3154)
         );
  INV_X1 U4021 ( .A(n3227), .ZN(n3169) );
  AOI22_X1 U4022 ( .A1(n4096), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4023 ( .A1(n4151), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4024 ( .A1(n3856), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4025 ( .A1(n3988), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3157) );
  NAND4_X1 U4026 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .ZN(n3168)
         );
  AOI22_X1 U4027 ( .A1(n4173), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4028 ( .A1(n2991), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4029 ( .A1(n3051), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4030 ( .A1(n2998), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3163) );
  NAND4_X1 U4031 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3167)
         );
  OAI211_X1 U4032 ( .C1(n3169), .C2(n6065), .A(n3389), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3170) );
  INV_X1 U4033 ( .A(n3170), .ZN(n3171) );
  NAND2_X1 U4034 ( .A1(n3173), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3218) );
  NOR2_X1 U4035 ( .A1(n3510), .A2(n6562), .ZN(n3260) );
  INV_X1 U4036 ( .A(n3392), .ZN(n3378) );
  NAND2_X1 U4037 ( .A1(n3260), .A2(n3378), .ZN(n3222) );
  MUX2_X1 U4038 ( .A(n3218), .B(n3222), .S(n3227), .Z(n3175) );
  NAND2_X2 U4039 ( .A1(n3178), .A2(n3217), .ZN(n4942) );
  INV_X1 U4040 ( .A(n3179), .ZN(n4249) );
  NAND2_X1 U4041 ( .A1(n3180), .A2(n3515), .ZN(n3277) );
  OAI21_X1 U4042 ( .B1(n4249), .B2(n3227), .A(n3277), .ZN(n3181) );
  INV_X1 U4043 ( .A(n3181), .ZN(n3182) );
  XNOR2_X1 U4044 ( .A(n3233), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4365)
         );
  INV_X1 U4045 ( .A(n3183), .ZN(n3185) );
  NOR2_X1 U4046 ( .A1(n3508), .A2(n6065), .ZN(n3184) );
  INV_X1 U4047 ( .A(n3496), .ZN(n3187) );
  NOR2_X1 U4048 ( .A1(n3637), .A2(n3491), .ZN(n3186) );
  AND2_X2 U4049 ( .A1(n3485), .A2(n6065), .ZN(n4255) );
  INV_X1 U4050 ( .A(n3188), .ZN(n3191) );
  NAND2_X1 U4051 ( .A1(n3681), .A2(n5503), .ZN(n3629) );
  AOI21_X1 U4052 ( .B1(n4255), .B2(n3191), .A(n3625), .ZN(n3192) );
  NAND2_X1 U4053 ( .A1(n4303), .A2(n3192), .ZN(n3193) );
  NAND2_X1 U4054 ( .A1(n3193), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3199) );
  XNOR2_X1 U4055 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5156) );
  INV_X1 U4056 ( .A(n5156), .ZN(n6255) );
  INV_X1 U4057 ( .A(n4239), .ZN(n3196) );
  INV_X1 U4058 ( .A(n3506), .ZN(n3194) );
  AND2_X1 U4059 ( .A1(n3194), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3195)
         );
  AOI21_X1 U4060 ( .B1(n6255), .B2(n3196), .A(n3195), .ZN(n3200) );
  INV_X1 U4061 ( .A(n3200), .ZN(n3197) );
  NOR2_X1 U4062 ( .A1(n3197), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3198)
         );
  OAI211_X1 U4063 ( .C1(n3240), .C2(n4339), .A(n3200), .B(n3199), .ZN(n3238)
         );
  XNOR2_X1 U4064 ( .A(n3237), .B(n3201), .ZN(n4332) );
  NAND2_X1 U4065 ( .A1(n4332), .A2(n6562), .ZN(n3216) );
  INV_X1 U4066 ( .A(n3010), .ZN(n3202) );
  AOI22_X1 U4067 ( .A1(n4096), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4068 ( .A1(n4151), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4069 ( .A1(n3856), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4070 ( .A1(n4057), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3203) );
  NAND4_X1 U4071 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3214)
         );
  AOI22_X1 U4072 ( .A1(n2992), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4073 ( .A1(n4173), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4074 ( .A1(n4145), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4075 ( .A1(n4150), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3209) );
  NAND4_X1 U4076 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3213)
         );
  NAND2_X1 U4077 ( .A1(n3260), .A2(n3226), .ZN(n3215) );
  OAI21_X2 U4078 ( .B1(n3690), .B2(STATE2_REG_0__SCAN_IN), .A(n3221), .ZN(
        n3269) );
  INV_X1 U4079 ( .A(n3226), .ZN(n3224) );
  NAND2_X1 U4080 ( .A1(n3180), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3262) );
  INV_X1 U4081 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6694) );
  OR2_X1 U4082 ( .A1(n3471), .A2(n6694), .ZN(n3223) );
  OAI211_X1 U4083 ( .C1(n3224), .C2(n3262), .A(n3223), .B(n3222), .ZN(n3268)
         );
  XNOR2_X1 U4084 ( .A(n3269), .B(n3268), .ZN(n3225) );
  INV_X1 U4085 ( .A(n3447), .ZN(n3498) );
  NAND2_X1 U4086 ( .A1(n4429), .A2(n3498), .ZN(n3232) );
  NAND2_X1 U4087 ( .A1(n3226), .A2(n3227), .ZN(n3275) );
  OAI21_X1 U4088 ( .B1(n3227), .B2(n3226), .A(n3275), .ZN(n3229) );
  OAI211_X1 U4089 ( .C1(n3229), .C2(n4249), .A(n3228), .B(n3491), .ZN(n3230)
         );
  INV_X1 U4090 ( .A(n3230), .ZN(n3231) );
  NAND2_X1 U4091 ( .A1(n3232), .A2(n3231), .ZN(n4364) );
  NAND2_X1 U4092 ( .A1(n4365), .A2(n4364), .ZN(n4363) );
  INV_X1 U4093 ( .A(n3233), .ZN(n3234) );
  NAND2_X1 U4094 ( .A1(n3234), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3235)
         );
  NAND2_X1 U4095 ( .A1(n3237), .A2(n3236), .ZN(n3239) );
  NAND2_X1 U4096 ( .A1(n3239), .A2(n3238), .ZN(n3247) );
  INV_X1 U4097 ( .A(n3247), .ZN(n3245) );
  INV_X1 U4098 ( .A(n3240), .ZN(n3285) );
  NAND2_X1 U4099 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4100 ( .A1(n3241), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3242) );
  NOR2_X1 U4101 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n4769), .ZN(n5160)
         );
  NAND2_X1 U4102 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5160), .ZN(n4731) );
  AND2_X1 U4103 ( .A1(n3242), .A2(n4731), .ZN(n4526) );
  OAI22_X1 U4104 ( .A1(n4239), .A2(n4526), .B1(n3506), .B2(n4642), .ZN(n3243)
         );
  INV_X1 U4105 ( .A(n3246), .ZN(n3244) );
  NAND2_X1 U4106 ( .A1(n3247), .A2(n3246), .ZN(n3248) );
  NAND2_X1 U4107 ( .A1(n3284), .A2(n3248), .ZN(n4374) );
  AOI22_X1 U4108 ( .A1(n4151), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4109 ( .A1(n2994), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4110 ( .A1(n3051), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4111 ( .A1(n4057), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3249) );
  NAND4_X1 U4112 ( .A1(n3252), .A2(n3251), .A3(n3250), .A4(n3249), .ZN(n3259)
         );
  AOI22_X1 U4113 ( .A1(n4096), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4114 ( .A1(n2992), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4115 ( .A1(n4173), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4116 ( .A1(n3856), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3254) );
  NAND4_X1 U4117 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3258)
         );
  INV_X1 U4118 ( .A(n3260), .ZN(n3261) );
  OAI22_X2 U4119 ( .A1(n4374), .A2(STATE2_REG_0__SCAN_IN), .B1(n3276), .B2(
        n3261), .ZN(n3266) );
  INV_X1 U4120 ( .A(n3262), .ZN(n3264) );
  AOI22_X1 U4121 ( .A1(n3354), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3264), 
        .B2(n3263), .ZN(n3265) );
  OAI21_X1 U4122 ( .B1(n3269), .B2(n3268), .A(n3267), .ZN(n3271) );
  NAND2_X1 U4123 ( .A1(n3269), .A2(n3268), .ZN(n3270) );
  NAND2_X1 U4124 ( .A1(n3310), .A2(n3274), .ZN(n4433) );
  OR2_X1 U4125 ( .A1(n4433), .A2(n3447), .ZN(n3281) );
  NAND2_X1 U4126 ( .A1(n3275), .A2(n3276), .ZN(n3303) );
  OAI21_X1 U4127 ( .B1(n3276), .B2(n3275), .A(n3303), .ZN(n3279) );
  INV_X1 U4128 ( .A(n3277), .ZN(n3278) );
  AOI21_X1 U4129 ( .B1(n3279), .B2(n3179), .A(n3278), .ZN(n3280) );
  OAI21_X1 U4130 ( .B1(n6183), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6182), 
        .ZN(n3283) );
  NAND2_X1 U4131 ( .A1(n6183), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3282)
         );
  NAND2_X1 U4132 ( .A1(n3283), .A2(n3282), .ZN(n5368) );
  NAND2_X1 U4133 ( .A1(n3285), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3288) );
  NOR3_X1 U4134 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4642), .A3(n4769), 
        .ZN(n6299) );
  NAND3_X1 U4135 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4854) );
  INV_X1 U4136 ( .A(n4854), .ZN(n4447) );
  NAND2_X1 U4137 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4447), .ZN(n4512) );
  OAI21_X1 U4138 ( .B1(n6327), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n4512), 
        .ZN(n4691) );
  OAI22_X1 U4139 ( .A1(n4691), .A2(n4239), .B1(n3506), .B2(n6544), .ZN(n3286)
         );
  INV_X1 U4140 ( .A(n3286), .ZN(n3287) );
  NAND2_X1 U4141 ( .A1(n4279), .A2(n6562), .ZN(n3302) );
  INV_X1 U4142 ( .A(n3475), .ZN(n3463) );
  AOI22_X1 U4143 ( .A1(n4151), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4144 ( .A1(n4172), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3292) );
  BUF_X1 U4145 ( .A(n3051), .Z(n3994) );
  AOI22_X1 U4146 ( .A1(n3994), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4147 ( .A1(n4057), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3290) );
  NAND4_X1 U4148 ( .A1(n3293), .A2(n3292), .A3(n3291), .A4(n3290), .ZN(n3300)
         );
  AOI22_X1 U4149 ( .A1(n4096), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4150 ( .A1(n2992), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3297) );
  INV_X1 U4151 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6711) );
  AOI22_X1 U4152 ( .A1(n4173), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4153 ( .A1(n3856), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3295) );
  NAND4_X1 U4154 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3299)
         );
  AOI22_X1 U4155 ( .A1(n3463), .A2(n3304), .B1(n3354), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4156 ( .A1(n3704), .A2(n3498), .ZN(n3306) );
  NAND2_X1 U4157 ( .A1(n3303), .A2(n3304), .ZN(n3347) );
  OAI211_X1 U4158 ( .C1(n3304), .C2(n3303), .A(n3347), .B(n3179), .ZN(n3305)
         );
  INV_X1 U4159 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U4160 ( .A1(n5368), .A2(n5369), .ZN(n3309) );
  NAND2_X1 U4161 ( .A1(n3307), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3308)
         );
  NAND2_X1 U4162 ( .A1(n3309), .A2(n3308), .ZN(n4418) );
  INV_X1 U4163 ( .A(n3310), .ZN(n3311) );
  NAND2_X1 U4164 ( .A1(n3311), .A2(n4519), .ZN(n3325) );
  NAND2_X1 U4165 ( .A1(n3354), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4166 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4173), .B1(n3094), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4167 ( .A1(n4151), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4168 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4144), .B1(n4172), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4169 ( .A1(n2992), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3312) );
  NAND4_X1 U4170 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), .ZN(n3321)
         );
  AOI22_X1 U4171 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4150), .B1(n3994), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4172 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4096), .B1(n3001), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4173 ( .A1(n4057), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4174 ( .A1(n3988), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3316) );
  NAND4_X1 U4175 ( .A1(n3319), .A2(n3318), .A3(n3317), .A4(n3316), .ZN(n3320)
         );
  NOR2_X1 U4176 ( .A1(n3321), .A2(n3320), .ZN(n3346) );
  OR2_X1 U4177 ( .A1(n3475), .A2(n3346), .ZN(n3322) );
  NOR2_X2 U4178 ( .A1(n3325), .A2(n3324), .ZN(n3344) );
  INV_X1 U4179 ( .A(n3344), .ZN(n3327) );
  NAND2_X1 U4180 ( .A1(n3325), .A2(n3324), .ZN(n3326) );
  XNOR2_X1 U4181 ( .A(n3347), .B(n3346), .ZN(n3328) );
  INV_X1 U4182 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4423) );
  XNOR2_X1 U4183 ( .A(n3329), .B(n4423), .ZN(n4417) );
  NAND2_X1 U4184 ( .A1(n4418), .A2(n4417), .ZN(n3331) );
  NAND2_X1 U4185 ( .A1(n3329), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3330)
         );
  NAND2_X1 U4186 ( .A1(n3331), .A2(n3330), .ZN(n4496) );
  INV_X1 U4187 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4598) );
  AOI22_X1 U4188 ( .A1(n4151), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4189 ( .A1(n4172), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4190 ( .A1(n3051), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4191 ( .A1(n4057), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3332) );
  NAND4_X1 U4192 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3341)
         );
  AOI22_X1 U4193 ( .A1(n4096), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4194 ( .A1(n2992), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4195 ( .A1(n4173), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4196 ( .A1(n3856), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3336) );
  NAND4_X1 U4197 ( .A1(n3339), .A2(n3338), .A3(n3337), .A4(n3336), .ZN(n3340)
         );
  INV_X1 U4198 ( .A(n3348), .ZN(n3342) );
  OAI22_X1 U4199 ( .A1(n3471), .A2(n4598), .B1(n3475), .B2(n3342), .ZN(n3343)
         );
  NAND2_X1 U4200 ( .A1(n3344), .A2(n3343), .ZN(n3371) );
  NAND2_X1 U4201 ( .A1(n3371), .A2(n3345), .ZN(n3726) );
  NOR2_X1 U4202 ( .A1(n3347), .A2(n3346), .ZN(n3349) );
  NAND2_X1 U4203 ( .A1(n3349), .A2(n3348), .ZN(n3380) );
  OAI211_X1 U4204 ( .C1(n3349), .C2(n3348), .A(n3380), .B(n3179), .ZN(n3350)
         );
  INV_X1 U4205 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4504) );
  XNOR2_X1 U4206 ( .A(n3351), .B(n4504), .ZN(n4497) );
  NAND2_X1 U4207 ( .A1(n4496), .A2(n4497), .ZN(n3353) );
  NAND2_X1 U4208 ( .A1(n3351), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3352)
         );
  NAND2_X1 U4209 ( .A1(n3353), .A2(n3352), .ZN(n4563) );
  NAND2_X1 U4210 ( .A1(n3354), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4211 ( .A1(n4150), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4212 ( .A1(n4151), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4213 ( .A1(n3856), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4214 ( .A1(n3051), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3355) );
  NAND4_X1 U4215 ( .A1(n3358), .A2(n3357), .A3(n3356), .A4(n3355), .ZN(n3364)
         );
  AOI22_X1 U4216 ( .A1(n2991), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4217 ( .A1(n4096), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4218 ( .A1(n4173), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4219 ( .A1(n4057), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3359) );
  NAND4_X1 U4220 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3363)
         );
  INV_X1 U4221 ( .A(n3381), .ZN(n3365) );
  OR2_X1 U4222 ( .A1(n3475), .A2(n3365), .ZN(n3366) );
  NAND2_X1 U4223 ( .A1(n3371), .A2(n3370), .ZN(n3739) );
  NAND3_X1 U4224 ( .A1(n3391), .A2(n3739), .A3(n3498), .ZN(n3374) );
  XNOR2_X1 U4225 ( .A(n3380), .B(n3381), .ZN(n3372) );
  NAND2_X1 U4226 ( .A1(n3372), .A2(n3179), .ZN(n3373) );
  NAND2_X1 U4227 ( .A1(n3374), .A2(n3373), .ZN(n3375) );
  INV_X1 U4228 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3543) );
  XNOR2_X1 U4229 ( .A(n3375), .B(n3543), .ZN(n4564) );
  NAND2_X1 U4230 ( .A1(n4563), .A2(n4564), .ZN(n3377) );
  NAND2_X1 U4231 ( .A1(n3375), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3376)
         );
  NAND2_X1 U4232 ( .A1(n3377), .A2(n3376), .ZN(n5018) );
  INV_X1 U4233 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4627) );
  OAI22_X1 U4234 ( .A1(n3471), .A2(n4627), .B1(n3475), .B2(n3378), .ZN(n3379)
         );
  NAND2_X1 U4235 ( .A1(n3747), .A2(n3498), .ZN(n3385) );
  INV_X1 U4236 ( .A(n3380), .ZN(n3382) );
  NAND2_X1 U4237 ( .A1(n3382), .A2(n3381), .ZN(n3394) );
  XNOR2_X1 U4238 ( .A(n3394), .B(n3392), .ZN(n3383) );
  NAND2_X1 U4239 ( .A1(n3383), .A2(n3179), .ZN(n3384) );
  NAND2_X1 U4240 ( .A1(n3385), .A2(n3384), .ZN(n3386) );
  INV_X1 U4241 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6225) );
  XNOR2_X1 U4242 ( .A(n3386), .B(n6225), .ZN(n5019) );
  NAND2_X1 U4243 ( .A1(n5018), .A2(n5019), .ZN(n3388) );
  NAND2_X1 U4244 ( .A1(n3386), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3387)
         );
  NAND2_X1 U4245 ( .A1(n3388), .A2(n3387), .ZN(n5024) );
  NOR2_X1 U4246 ( .A1(n3389), .A2(n3447), .ZN(n3390) );
  NAND2_X1 U4247 ( .A1(n3179), .A2(n3392), .ZN(n3393) );
  OR2_X1 U4248 ( .A1(n3394), .A2(n3393), .ZN(n3395) );
  NAND2_X1 U4249 ( .A1(n5576), .A2(n3395), .ZN(n3396) );
  INV_X1 U4250 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5035) );
  XNOR2_X1 U4251 ( .A(n3396), .B(n5035), .ZN(n5025) );
  NAND2_X1 U4252 ( .A1(n5024), .A2(n5025), .ZN(n3398) );
  NAND2_X1 U4253 ( .A1(n3396), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3397)
         );
  NAND2_X1 U4254 ( .A1(n3398), .A2(n3397), .ZN(n5083) );
  INV_X1 U4255 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5113) );
  NOR2_X1 U4256 ( .A1(n5576), .A2(n5113), .ZN(n3399) );
  INV_X4 U4257 ( .A(n4227), .ZN(n5708) );
  NAND2_X1 U4258 ( .A1(n5708), .A2(n5113), .ZN(n3400) );
  NAND2_X1 U4259 ( .A1(n3401), .A2(n3400), .ZN(n5103) );
  INV_X1 U4260 ( .A(n5103), .ZN(n3402) );
  INV_X1 U4261 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U4262 ( .A1(n3402), .A2(n3005), .ZN(n3403) );
  OR2_X1 U4263 ( .A1(n5708), .A2(n5112), .ZN(n5104) );
  NAND2_X1 U4264 ( .A1(n3403), .A2(n5104), .ZN(n5198) );
  INV_X1 U4265 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3404) );
  NAND2_X1 U4266 ( .A1(n5708), .A2(n3404), .ZN(n5200) );
  NAND2_X1 U4267 ( .A1(n5198), .A2(n5200), .ZN(n3405) );
  NAND2_X1 U4268 ( .A1(n3405), .A2(n5201), .ZN(n5208) );
  INV_X1 U4269 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3562) );
  NOR2_X1 U4270 ( .A1(n5576), .A2(n3562), .ZN(n5236) );
  XNOR2_X1 U4271 ( .A(n5576), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5242)
         );
  INV_X1 U4272 ( .A(n5242), .ZN(n3406) );
  INV_X1 U4273 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5265) );
  INV_X1 U4274 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5898) );
  INV_X1 U4275 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3653) );
  NAND2_X1 U4276 ( .A1(n5708), .A2(n3653), .ZN(n3407) );
  NAND2_X1 U4277 ( .A1(n5708), .A2(n3562), .ZN(n5237) );
  NAND2_X1 U4278 ( .A1(n5708), .A2(n5265), .ZN(n3408) );
  OAI21_X1 U4279 ( .B1(n5208), .B2(n5613), .A(n3409), .ZN(n3410) );
  NAND2_X1 U4280 ( .A1(n3410), .A2(n5616), .ZN(n5315) );
  INV_X1 U4281 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U4282 ( .A1(n5576), .A2(n6708), .ZN(n3411) );
  NAND2_X1 U4283 ( .A1(n5315), .A2(n3411), .ZN(n5598) );
  INV_X1 U4284 ( .A(n5598), .ZN(n3412) );
  NAND2_X1 U4285 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3659) );
  NAND2_X1 U4286 ( .A1(n3412), .A2(n3015), .ZN(n5569) );
  NOR2_X1 U4287 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5596) );
  INV_X1 U4288 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5726) );
  AND2_X1 U4289 ( .A1(n5596), .A2(n5726), .ZN(n3413) );
  NAND2_X1 U4290 ( .A1(n5569), .A2(n3414), .ZN(n4221) );
  INV_X1 U4291 ( .A(n4221), .ZN(n3416) );
  NOR2_X1 U4292 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5693) );
  NOR2_X1 U4293 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5680) );
  INV_X1 U4294 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4234) );
  INV_X1 U4295 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5668) );
  AND4_X1 U4296 ( .A1(n5693), .A2(n5680), .A3(n4234), .A4(n5668), .ZN(n3415)
         );
  NAND2_X1 U4297 ( .A1(n3416), .A2(n3006), .ZN(n5536) );
  AND2_X1 U4298 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5694) );
  AND2_X1 U4299 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5679) );
  AND2_X1 U4300 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3664) );
  NAND3_X1 U4301 ( .A1(n5694), .A2(n5679), .A3(n3664), .ZN(n3671) );
  NAND2_X1 U4302 ( .A1(n5576), .A2(n3671), .ZN(n3417) );
  NAND2_X1 U4303 ( .A1(n5536), .A2(n3417), .ZN(n5855) );
  XNOR2_X1 U4304 ( .A(n5708), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5856)
         );
  INV_X1 U4305 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6612) );
  NOR2_X2 U4306 ( .A1(n3419), .A2(n3418), .ZN(n5517) );
  INV_X1 U4307 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5659) );
  NOR2_X1 U4308 ( .A1(n4227), .A2(n5659), .ZN(n5554) );
  NAND2_X1 U4309 ( .A1(n5517), .A2(n5554), .ZN(n5545) );
  NAND2_X1 U4310 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3652) );
  AND2_X1 U4311 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3674) );
  INV_X1 U4312 ( .A(n3419), .ZN(n5854) );
  NOR2_X1 U4313 ( .A1(n5576), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5553)
         );
  INV_X1 U4314 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5640) );
  INV_X1 U4315 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5650) );
  NAND3_X1 U4316 ( .A1(n5553), .A2(n5640), .A3(n5650), .ZN(n5518) );
  NOR4_X1 U4317 ( .A1(n5854), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5518), .ZN(n3420) );
  AOI21_X1 U4318 ( .B1(n5527), .B2(n3674), .A(n3420), .ZN(n3421) );
  INV_X1 U4319 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4336) );
  XNOR2_X1 U4320 ( .A(n3421), .B(n4336), .ZN(n4248) );
  INV_X1 U4321 ( .A(n4248), .ZN(n3513) );
  INV_X1 U4322 ( .A(STATE_REG_0__SCAN_IN), .ZN(n3422) );
  NAND2_X1 U4323 ( .A1(n3423), .A2(n3422), .ZN(n6461) );
  NAND2_X1 U4324 ( .A1(n6461), .A2(n3648), .ZN(n3445) );
  NAND2_X1 U4325 ( .A1(n6408), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3453) );
  INV_X1 U4326 ( .A(n3453), .ZN(n3424) );
  XNOR2_X1 U4327 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3439) );
  NAND2_X1 U4328 ( .A1(n3424), .A2(n3439), .ZN(n3426) );
  NAND2_X1 U4329 ( .A1(n4769), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3425) );
  NAND2_X1 U4330 ( .A1(n3426), .A2(n3425), .ZN(n3438) );
  XNOR2_X1 U4331 ( .A(n5389), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3437)
         );
  INV_X1 U4332 ( .A(n3437), .ZN(n3427) );
  NAND2_X1 U4333 ( .A1(n3438), .A2(n3427), .ZN(n3429) );
  NAND2_X1 U4334 ( .A1(n4642), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3428) );
  NAND2_X1 U4335 ( .A1(n3429), .A2(n3428), .ZN(n3434) );
  XNOR2_X1 U4336 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3432) );
  NAND2_X1 U4337 ( .A1(n3434), .A2(n3432), .ZN(n3431) );
  NAND2_X1 U4338 ( .A1(n6544), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3430) );
  NAND2_X1 U4339 ( .A1(n3431), .A2(n3430), .ZN(n3441) );
  INV_X1 U4340 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6419) );
  INV_X1 U4341 ( .A(n3432), .ZN(n3433) );
  XNOR2_X1 U4342 ( .A(n3434), .B(n3433), .ZN(n3435) );
  NAND2_X1 U4343 ( .A1(n3436), .A2(n3435), .ZN(n3474) );
  XNOR2_X1 U4344 ( .A(n3438), .B(n3437), .ZN(n3466) );
  XNOR2_X1 U4345 ( .A(n3439), .B(n3453), .ZN(n3448) );
  NAND2_X1 U4346 ( .A1(n3466), .A2(n3448), .ZN(n3444) );
  AND2_X1 U4347 ( .A1(n6419), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3440)
         );
  INV_X1 U4348 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U4349 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5905), .ZN(n3442) );
  NAND2_X1 U4350 ( .A1(n3443), .A2(n3442), .ZN(n3480) );
  OAI21_X1 U4351 ( .B1(n3474), .B2(n3444), .A(n3480), .ZN(n4195) );
  NOR2_X1 U4352 ( .A1(READY_N), .A2(n4195), .ZN(n4304) );
  NAND2_X1 U4353 ( .A1(n3445), .A2(n4304), .ZN(n3490) );
  INV_X1 U4354 ( .A(n3448), .ZN(n3450) );
  OR2_X1 U4355 ( .A1(n3475), .A2(n4510), .ZN(n3446) );
  NAND2_X1 U4356 ( .A1(n3446), .A2(n3491), .ZN(n3460) );
  NAND2_X1 U4357 ( .A1(n3448), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3451) );
  NAND2_X1 U4358 ( .A1(n3481), .A2(n3451), .ZN(n3449) );
  OAI21_X1 U4359 ( .B1(n3450), .B2(n3460), .A(n3449), .ZN(n3462) );
  INV_X1 U4360 ( .A(n3451), .ZN(n3459) );
  NAND2_X1 U4361 ( .A1(n4347), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3452) );
  NAND2_X1 U4362 ( .A1(n3453), .A2(n3452), .ZN(n3454) );
  OAI21_X1 U4363 ( .B1(n3475), .B2(n3454), .A(n3481), .ZN(n3458) );
  INV_X1 U4364 ( .A(n3454), .ZN(n3455) );
  AOI21_X1 U4365 ( .B1(n3508), .B2(n3455), .A(n3180), .ZN(n3456) );
  AOI21_X1 U4366 ( .B1(n3190), .B2(n6065), .A(n3648), .ZN(n3464) );
  OR2_X1 U4367 ( .A1(n3456), .A2(n3464), .ZN(n3457) );
  OAI211_X1 U4368 ( .C1(n3460), .C2(n3459), .A(n3458), .B(n3457), .ZN(n3461)
         );
  NAND2_X1 U4369 ( .A1(n3462), .A2(n3461), .ZN(n3468) );
  OAI211_X1 U4370 ( .C1(n3468), .C2(n3464), .A(n3463), .B(n3466), .ZN(n3470)
         );
  INV_X1 U4371 ( .A(n3464), .ZN(n3465) );
  OAI21_X1 U4372 ( .B1(n3471), .B2(n3466), .A(n3465), .ZN(n3467) );
  NAND2_X1 U4373 ( .A1(n3468), .A2(n3467), .ZN(n3469) );
  NAND2_X1 U4374 ( .A1(n3470), .A2(n3469), .ZN(n3473) );
  NAND2_X1 U4375 ( .A1(n3471), .A2(n3474), .ZN(n3472) );
  INV_X1 U4376 ( .A(n3474), .ZN(n3478) );
  NOR2_X1 U4377 ( .A1(n3475), .A2(n3480), .ZN(n3476) );
  AOI21_X1 U4378 ( .B1(n6562), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n3476), 
        .ZN(n3477) );
  OAI21_X1 U4379 ( .B1(n3481), .B2(n3478), .A(n3477), .ZN(n3479) );
  INV_X1 U4380 ( .A(n3479), .ZN(n3483) );
  NAND2_X1 U4381 ( .A1(n4510), .A2(n6461), .ZN(n4203) );
  INV_X1 U4382 ( .A(READY_N), .ZN(n6462) );
  AND2_X1 U4383 ( .A1(n4203), .A2(n6462), .ZN(n3487) );
  NAND2_X1 U4384 ( .A1(n3629), .A2(n6065), .ZN(n3486) );
  AOI21_X1 U4385 ( .B1(n4308), .B2(n3487), .A(n3486), .ZN(n3488) );
  OR2_X1 U4386 ( .A1(n6407), .A2(n3488), .ZN(n3489) );
  MUX2_X1 U4387 ( .A(n3490), .B(n3489), .S(n4454), .Z(n3505) );
  NAND2_X1 U4388 ( .A1(n3492), .A2(n3491), .ZN(n4349) );
  NOR2_X1 U4389 ( .A1(n4349), .A2(n4510), .ZN(n3650) );
  NOR2_X1 U4390 ( .A1(n3630), .A2(n3637), .ZN(n3494) );
  NAND2_X1 U4391 ( .A1(n4349), .A2(n3180), .ZN(n3493) );
  NAND2_X1 U4392 ( .A1(n3494), .A2(n3493), .ZN(n3509) );
  INV_X1 U4393 ( .A(n4360), .ZN(n3495) );
  OR2_X1 U4394 ( .A1(n3496), .A2(n3495), .ZN(n3500) );
  AOI21_X1 U4395 ( .B1(n3498), .B2(n3497), .A(n3180), .ZN(n3499) );
  NAND2_X1 U4396 ( .A1(n3500), .A2(n3499), .ZN(n3640) );
  INV_X1 U4397 ( .A(n3640), .ZN(n3501) );
  NOR2_X1 U4398 ( .A1(n3509), .A2(n3501), .ZN(n3503) );
  NOR2_X1 U4399 ( .A1(n3503), .A2(n4259), .ZN(n4299) );
  AOI21_X1 U4400 ( .B1(n6407), .B2(n3650), .A(n4299), .ZN(n3504) );
  NAND2_X1 U4401 ( .A1(n3505), .A2(n3504), .ZN(n3507) );
  OR2_X1 U4402 ( .A1(n3509), .A2(n3508), .ZN(n6424) );
  INV_X1 U4403 ( .A(n4256), .ZN(n4990) );
  OR2_X1 U4404 ( .A1(n3509), .A2(n4990), .ZN(n4302) );
  AND2_X1 U4405 ( .A1(n6424), .A2(n4302), .ZN(n4262) );
  NAND2_X1 U4406 ( .A1(n4255), .A2(n3648), .ZN(n4309) );
  NAND2_X1 U4407 ( .A1(n3625), .A2(n3510), .ZN(n3511) );
  NAND4_X1 U4408 ( .A1(n4303), .A2(n4262), .A3(n4309), .A4(n3511), .ZN(n3512)
         );
  NAND2_X1 U4409 ( .A1(n3513), .A2(n6245), .ZN(n3680) );
  NOR2_X4 U4410 ( .A1(n5478), .A2(n4324), .ZN(n3608) );
  INV_X1 U4411 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U4412 ( .A1(n3608), .A2(n3514), .ZN(n3519) );
  INV_X1 U4413 ( .A(n3515), .ZN(n4460) );
  NAND2_X2 U4414 ( .A1(n4460), .A2(n6065), .ZN(n3609) );
  INV_X1 U4415 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U4416 ( .A1(n3609), .A2(n4369), .ZN(n3517) );
  NAND3_X1 U4417 ( .A1(n3517), .A2(n5478), .A3(n3516), .ZN(n3518) );
  NAND2_X1 U4418 ( .A1(n3519), .A2(n3518), .ZN(n3522) );
  NAND2_X1 U4419 ( .A1(n3609), .A2(EBX_REG_0__SCAN_IN), .ZN(n3521) );
  INV_X1 U4420 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U4421 ( .A1(n3621), .A2(n5052), .ZN(n3520) );
  NAND2_X1 U4422 ( .A1(n3521), .A2(n3520), .ZN(n4319) );
  XNOR2_X1 U4423 ( .A(n3522), .B(n4319), .ZN(n5363) );
  NAND2_X1 U4424 ( .A1(n5363), .A2(n4366), .ZN(n4368) );
  NAND2_X1 U4425 ( .A1(n4368), .A2(n3522), .ZN(n4412) );
  NAND2_X2 U4426 ( .A1(n3609), .A2(n3621), .ZN(n4318) );
  NAND2_X2 U4427 ( .A1(n4366), .A2(n5478), .ZN(n3606) );
  MUX2_X1 U4428 ( .A(n3606), .B(n3621), .S(EBX_REG_3__SCAN_IN), .Z(n3523) );
  OAI21_X1 U4429 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n4318), .A(n3523), 
        .ZN(n4438) );
  INV_X1 U4430 ( .A(n4438), .ZN(n3531) );
  NAND2_X1 U4431 ( .A1(n3609), .A2(EBX_REG_2__SCAN_IN), .ZN(n3525) );
  INV_X1 U4432 ( .A(n3609), .ZN(n3527) );
  NAND2_X1 U4433 ( .A1(n3527), .A2(n4324), .ZN(n3575) );
  NAND2_X1 U4434 ( .A1(n4324), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3528)
         );
  AND2_X1 U4435 ( .A1(n3575), .A2(n3528), .ZN(n3529) );
  INV_X1 U4436 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U4437 ( .A1(n3608), .A2(n3533), .ZN(n3537) );
  NAND2_X1 U4438 ( .A1(n3609), .A2(n4423), .ZN(n3535) );
  NAND2_X1 U4439 ( .A1(n4366), .A2(n3533), .ZN(n3534) );
  NAND3_X1 U4440 ( .A1(n3535), .A2(n3621), .A3(n3534), .ZN(n3536) );
  MUX2_X1 U4441 ( .A(n3606), .B(n3621), .S(EBX_REG_5__SCAN_IN), .Z(n3538) );
  INV_X1 U4442 ( .A(n3538), .ZN(n3540) );
  NOR2_X1 U4443 ( .A1(n4318), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3539)
         );
  NOR2_X1 U4444 ( .A1(n3540), .A2(n3539), .ZN(n4499) );
  NAND2_X1 U4445 ( .A1(n3621), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3541)
         );
  OAI211_X1 U4446 ( .C1(n4324), .C2(EBX_REG_7__SCAN_IN), .A(n3609), .B(n3541), 
        .ZN(n3542) );
  OAI21_X1 U4447 ( .B1(n3606), .B2(EBX_REG_7__SCAN_IN), .A(n3542), .ZN(n5012)
         );
  INV_X1 U4448 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U4449 ( .A1(n3608), .A2(n6044), .ZN(n3547) );
  NAND2_X1 U4450 ( .A1(n3609), .A2(n3543), .ZN(n3545) );
  NAND2_X1 U4451 ( .A1(n4366), .A2(n6044), .ZN(n3544) );
  NAND3_X1 U4452 ( .A1(n3545), .A2(n5478), .A3(n3544), .ZN(n3546) );
  MUX2_X1 U4453 ( .A(n3603), .B(n3609), .S(EBX_REG_8__SCAN_IN), .Z(n3552) );
  NAND2_X1 U4454 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n4324), .ZN(n3550)
         );
  AND2_X1 U4455 ( .A1(n3575), .A2(n3550), .ZN(n3551) );
  NOR2_X2 U4456 ( .A1(n5030), .A2(n5029), .ZN(n5073) );
  MUX2_X1 U4457 ( .A(n3606), .B(n3621), .S(EBX_REG_9__SCAN_IN), .Z(n3553) );
  INV_X1 U4458 ( .A(n3553), .ZN(n3555) );
  NOR2_X1 U4459 ( .A1(n4318), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3554)
         );
  NOR2_X1 U4460 ( .A1(n3555), .A2(n3554), .ZN(n5072) );
  NAND2_X1 U4461 ( .A1(n5073), .A2(n5072), .ZN(n5071) );
  MUX2_X1 U4462 ( .A(n3603), .B(n3609), .S(EBX_REG_10__SCAN_IN), .Z(n3558) );
  NAND2_X1 U4463 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4324), .ZN(n3556) );
  AND2_X1 U4464 ( .A1(n3575), .A2(n3556), .ZN(n3557) );
  NOR2_X2 U4465 ( .A1(n5071), .A2(n5109), .ZN(n5108) );
  MUX2_X1 U4466 ( .A(n3606), .B(n5478), .S(EBX_REG_11__SCAN_IN), .Z(n3559) );
  NAND2_X1 U4467 ( .A1(n3559), .A2(n3004), .ZN(n5140) );
  INV_X1 U4468 ( .A(EBX_REG_12__SCAN_IN), .ZN(n3563) );
  NAND2_X1 U4469 ( .A1(n3608), .A2(n3563), .ZN(n3567) );
  NAND2_X1 U4470 ( .A1(n3609), .A2(n3562), .ZN(n3565) );
  NAND2_X1 U4471 ( .A1(n4366), .A2(n3563), .ZN(n3564) );
  NAND3_X1 U4472 ( .A1(n3565), .A2(n3621), .A3(n3564), .ZN(n3566) );
  NAND2_X1 U4473 ( .A1(n3567), .A2(n3566), .ZN(n5221) );
  MUX2_X1 U4474 ( .A(n3606), .B(n5478), .S(EBX_REG_13__SCAN_IN), .Z(n3568) );
  OAI21_X1 U4475 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n4318), .A(n3568), 
        .ZN(n5253) );
  INV_X1 U4476 ( .A(n5253), .ZN(n3569) );
  MUX2_X1 U4477 ( .A(n3603), .B(n3609), .S(EBX_REG_14__SCAN_IN), .Z(n3572) );
  NAND2_X1 U4478 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4324), .ZN(n3570) );
  AND2_X1 U4479 ( .A1(n3575), .A2(n3570), .ZN(n3571) );
  MUX2_X1 U4480 ( .A(n3606), .B(n5478), .S(EBX_REG_15__SCAN_IN), .Z(n3573) );
  OAI21_X1 U4481 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n4318), .A(n3573), 
        .ZN(n5439) );
  MUX2_X1 U4482 ( .A(n3603), .B(n3609), .S(EBX_REG_16__SCAN_IN), .Z(n3577) );
  NAND2_X1 U4483 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4324), .ZN(n3574) );
  AND2_X1 U4484 ( .A1(n3575), .A2(n3574), .ZN(n3576) );
  NAND2_X1 U4485 ( .A1(n3577), .A2(n3576), .ZN(n5498) );
  AND2_X2 U4486 ( .A1(n5499), .A2(n5498), .ZN(n5496) );
  MUX2_X1 U4487 ( .A(n3606), .B(n5478), .S(EBX_REG_17__SCAN_IN), .Z(n3578) );
  OAI21_X1 U4488 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n4318), .A(n3578), 
        .ZN(n3579) );
  INV_X1 U4489 ( .A(n3579), .ZN(n5320) );
  INV_X1 U4490 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5312) );
  NAND2_X1 U4491 ( .A1(n3608), .A2(n5312), .ZN(n3583) );
  INV_X1 U4492 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U4493 ( .A1(n3609), .A2(n5713), .ZN(n3581) );
  NAND2_X1 U4494 ( .A1(n4366), .A2(n5312), .ZN(n3580) );
  NAND3_X1 U4495 ( .A1(n3581), .A2(n3621), .A3(n3580), .ZN(n3582) );
  AND2_X1 U4496 ( .A1(n3583), .A2(n3582), .ZN(n5310) );
  OR2_X2 U4497 ( .A1(n5339), .A2(n5310), .ZN(n5477) );
  INV_X1 U4498 ( .A(n4318), .ZN(n3636) );
  INV_X1 U4499 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4223) );
  NOR2_X1 U4500 ( .A1(n4324), .A2(EBX_REG_20__SCAN_IN), .ZN(n3584) );
  AOI21_X1 U4501 ( .B1(n3636), .B2(n4223), .A(n3584), .ZN(n5481) );
  OR2_X1 U4502 ( .A1(n4318), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3586)
         );
  INV_X1 U4503 ( .A(EBX_REG_18__SCAN_IN), .ZN(n3585) );
  NAND2_X1 U4504 ( .A1(n4366), .A2(n3585), .ZN(n5309) );
  NAND2_X1 U4505 ( .A1(n3586), .A2(n5309), .ZN(n5479) );
  INV_X1 U4506 ( .A(n3587), .ZN(n5399) );
  NAND2_X1 U4507 ( .A1(n5399), .A2(EBX_REG_20__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4508 ( .A1(n5479), .A2(n3621), .ZN(n3588) );
  OAI211_X1 U4509 ( .C1(n5481), .C2(n5479), .A(n3589), .B(n3588), .ZN(n3590)
         );
  NOR2_X2 U4510 ( .A1(n5477), .A2(n3590), .ZN(n5296) );
  MUX2_X1 U4511 ( .A(n3606), .B(n3621), .S(EBX_REG_21__SCAN_IN), .Z(n3591) );
  OAI21_X1 U4512 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4318), .A(n3591), 
        .ZN(n3592) );
  INV_X1 U4513 ( .A(n3592), .ZN(n5295) );
  NAND2_X1 U4514 ( .A1(n5296), .A2(n5295), .ZN(n5294) );
  INV_X1 U4515 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6721) );
  NAND2_X1 U4516 ( .A1(n3608), .A2(n6721), .ZN(n3597) );
  INV_X1 U4517 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3593) );
  NAND2_X1 U4518 ( .A1(n3609), .A2(n3593), .ZN(n3595) );
  NAND2_X1 U4519 ( .A1(n4366), .A2(n6721), .ZN(n3594) );
  NAND3_X1 U4520 ( .A1(n3595), .A2(n5478), .A3(n3594), .ZN(n3596) );
  AND2_X1 U4521 ( .A1(n3597), .A2(n3596), .ZN(n5334) );
  MUX2_X1 U4522 ( .A(n3606), .B(n3621), .S(EBX_REG_23__SCAN_IN), .Z(n3598) );
  OAI21_X1 U4523 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n4318), .A(n3598), 
        .ZN(n5426) );
  MUX2_X1 U4524 ( .A(n3603), .B(n3609), .S(EBX_REG_24__SCAN_IN), .Z(n3600) );
  NAND2_X1 U4525 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n4324), .ZN(n3599) );
  AND2_X1 U4526 ( .A1(n3600), .A2(n3599), .ZN(n4230) );
  MUX2_X1 U4527 ( .A(n3606), .B(n5478), .S(EBX_REG_25__SCAN_IN), .Z(n3601) );
  OAI21_X1 U4528 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4318), .A(n3601), 
        .ZN(n3602) );
  INV_X1 U4529 ( .A(n3602), .ZN(n5470) );
  AND2_X2 U4530 ( .A1(n5469), .A2(n5470), .ZN(n5467) );
  MUX2_X1 U4531 ( .A(n3603), .B(n3609), .S(EBX_REG_26__SCAN_IN), .Z(n3605) );
  NAND2_X1 U4532 ( .A1(n4324), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3604) );
  NAND2_X1 U4533 ( .A1(n3605), .A2(n3604), .ZN(n5461) );
  MUX2_X1 U4534 ( .A(n3606), .B(n3621), .S(EBX_REG_27__SCAN_IN), .Z(n3607) );
  OAI21_X1 U4535 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4318), .A(n3607), 
        .ZN(n5647) );
  INV_X1 U4536 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U4537 ( .A1(n3608), .A2(n5734), .ZN(n3613) );
  NAND2_X1 U4538 ( .A1(n3609), .A2(n5640), .ZN(n3611) );
  NAND2_X1 U4539 ( .A1(n4366), .A2(n5734), .ZN(n3610) );
  NAND3_X1 U4540 ( .A1(n3611), .A2(n5478), .A3(n3610), .ZN(n3612) );
  NAND2_X1 U4541 ( .A1(n3613), .A2(n3612), .ZN(n5452) );
  NAND2_X2 U4542 ( .A1(n5451), .A2(n5452), .ZN(n5454) );
  INV_X1 U4543 ( .A(EBX_REG_29__SCAN_IN), .ZN(n3617) );
  OR2_X1 U4544 ( .A1(n4318), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3615)
         );
  NAND2_X1 U4545 ( .A1(n4366), .A2(n3617), .ZN(n3614) );
  NAND2_X1 U4546 ( .A1(n3615), .A2(n3614), .ZN(n3620) );
  INV_X1 U4547 ( .A(n3620), .ZN(n3616) );
  MUX2_X1 U4548 ( .A(n3617), .B(n3616), .S(n3621), .Z(n5414) );
  NAND2_X1 U4549 ( .A1(n4318), .A2(EBX_REG_30__SCAN_IN), .ZN(n3619) );
  NAND2_X1 U4550 ( .A1(n4324), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3618) );
  AND2_X1 U4551 ( .A1(n3619), .A2(n3618), .ZN(n5401) );
  NAND2_X1 U4552 ( .A1(n5414), .A2(n5401), .ZN(n3622) );
  OR2_X2 U4553 ( .A1(n5454), .A2(n3620), .ZN(n5402) );
  OAI21_X1 U4554 ( .B1(n5454), .B2(n3622), .A(n5398), .ZN(n3624) );
  OAI22_X1 U4555 ( .A1(n4318), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4324), .ZN(n3623) );
  NAND2_X1 U4556 ( .A1(n3625), .A2(n3132), .ZN(n3626) );
  NAND2_X1 U4557 ( .A1(n4308), .A2(n3179), .ZN(n6402) );
  NAND2_X1 U4558 ( .A1(n3626), .A2(n6402), .ZN(n3627) );
  INV_X1 U4559 ( .A(n6240), .ZN(n3628) );
  INV_X1 U4560 ( .A(n3674), .ZN(n3668) );
  INV_X1 U4561 ( .A(n3629), .ZN(n5378) );
  NAND2_X1 U4562 ( .A1(n3630), .A2(n5399), .ZN(n3632) );
  OAI211_X1 U4563 ( .C1(n4454), .C2(n5378), .A(n3632), .B(n3631), .ZN(n3633)
         );
  INV_X1 U4564 ( .A(n3633), .ZN(n3641) );
  OR2_X1 U4565 ( .A1(n3634), .A2(n3635), .ZN(n4300) );
  NAND2_X1 U4566 ( .A1(n3636), .A2(n4300), .ZN(n3638) );
  NAND2_X1 U4567 ( .A1(n3638), .A2(n3637), .ZN(n3639) );
  NAND4_X1 U4568 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n4284)
         );
  OAI22_X1 U4569 ( .A1(n4280), .A2(n3688), .B1(n4281), .B2(n6065), .ZN(n3643)
         );
  INV_X1 U4570 ( .A(n3643), .ZN(n3645) );
  INV_X1 U4571 ( .A(n4322), .ZN(n3644) );
  OR3_X1 U4572 ( .A1(n4349), .A2(n6065), .A3(n3644), .ZN(n4380) );
  NAND2_X1 U4573 ( .A1(n3645), .A2(n4380), .ZN(n3646) );
  NOR2_X1 U4574 ( .A1(n4284), .A2(n3646), .ZN(n3651) );
  INV_X1 U4575 ( .A(n3651), .ZN(n3647) );
  INV_X1 U4576 ( .A(n5215), .ZN(n3649) );
  AND2_X1 U4577 ( .A1(n4259), .A2(n3648), .ZN(n5729) );
  NAND2_X1 U4578 ( .A1(n3655), .A2(n5729), .ZN(n5248) );
  NAND2_X1 U4579 ( .A1(n5214), .A2(n5698), .ZN(n5883) );
  INV_X1 U4580 ( .A(n3652), .ZN(n3673) );
  INV_X1 U4581 ( .A(n5883), .ZN(n5107) );
  NAND2_X1 U4582 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U4583 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5249) );
  NOR2_X1 U4584 ( .A1(n3653), .A2(n5249), .ZN(n5263) );
  NAND2_X1 U4585 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5263), .ZN(n5887) );
  NAND2_X1 U4586 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5888) );
  NOR2_X1 U4587 ( .A1(n5887), .A2(n5888), .ZN(n3657) );
  NOR2_X1 U4588 ( .A1(n6225), .A2(n5035), .ZN(n5111) );
  NAND3_X1 U4589 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5111), .ZN(n3656) );
  AOI21_X1 U4590 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6243) );
  NOR2_X1 U4591 ( .A1(n6235), .A2(n4423), .ZN(n4502) );
  INV_X1 U4592 ( .A(n4502), .ZN(n3654) );
  NOR2_X1 U4593 ( .A1(n6243), .A2(n3654), .ZN(n4503) );
  NAND4_X1 U4594 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6241), .A4(n4503), .ZN(n5032) );
  NOR2_X1 U4595 ( .A1(n3656), .A2(n5032), .ZN(n5216) );
  NAND2_X1 U4596 ( .A1(n3657), .A2(n5216), .ZN(n3670) );
  NOR2_X1 U4597 ( .A1(n6241), .A2(n5215), .ZN(n5245) );
  NOR2_X1 U4598 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5245), .ZN(n4343)
         );
  INV_X2 U4599 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U4600 ( .A1(n6562), .A2(n6560), .ZN(n6449) );
  INV_X1 U4601 ( .A(n6449), .ZN(n6443) );
  NOR2_X1 U4602 ( .A1(n6238), .A2(n3655), .ZN(n4344) );
  NOR2_X1 U4603 ( .A1(n4343), .A2(n4344), .ZN(n4422) );
  NAND2_X1 U4604 ( .A1(n4422), .A2(n5698), .ZN(n5212) );
  INV_X1 U4605 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6247) );
  NOR2_X1 U4606 ( .A1(n6247), .A2(n4369), .ZN(n6242) );
  NAND4_X1 U4607 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6242), .A4(n4502), .ZN(n5033) );
  NOR2_X1 U4608 ( .A1(n5033), .A2(n3656), .ZN(n5219) );
  AND2_X1 U4609 ( .A1(n5219), .A2(n3657), .ZN(n3669) );
  NOR2_X1 U4610 ( .A1(n5214), .A2(n3669), .ZN(n3658) );
  AOI21_X1 U4611 ( .B1(n3670), .B2(n5212), .A(n3658), .ZN(n5702) );
  INV_X1 U4612 ( .A(n5694), .ZN(n4233) );
  OAI21_X1 U4613 ( .B1(n4233), .B2(n3659), .A(n5883), .ZN(n3660) );
  AND2_X1 U4614 ( .A1(n5702), .A2(n3660), .ZN(n5676) );
  INV_X1 U4615 ( .A(n5679), .ZN(n3661) );
  NAND2_X1 U4616 ( .A1(n5883), .A2(n3661), .ZN(n3662) );
  AND2_X1 U4617 ( .A1(n5676), .A2(n3662), .ZN(n5667) );
  INV_X1 U4618 ( .A(n5248), .ZN(n5220) );
  NOR2_X1 U4619 ( .A1(n5220), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4371)
         );
  NOR2_X1 U4620 ( .A1(n5214), .A2(n4371), .ZN(n6248) );
  INV_X1 U4621 ( .A(n6248), .ZN(n3663) );
  NAND2_X1 U4622 ( .A1(n5698), .A2(n3663), .ZN(n3666) );
  INV_X1 U4623 ( .A(n3664), .ZN(n3665) );
  NAND2_X1 U4624 ( .A1(n3666), .A2(n3665), .ZN(n3667) );
  NAND2_X1 U4625 ( .A1(n5667), .A2(n3667), .ZN(n5874) );
  AOI21_X1 U4626 ( .B1(n5883), .B2(n5661), .A(n5874), .ZN(n5639) );
  OAI21_X1 U4627 ( .B1(n3673), .B2(n5107), .A(n5639), .ZN(n5632) );
  AOI21_X1 U4628 ( .B1(n3668), .B2(n5883), .A(n5632), .ZN(n5626) );
  NAND2_X1 U4629 ( .A1(n3669), .A2(n6248), .ZN(n5699) );
  NAND2_X1 U4630 ( .A1(n3670), .A2(n5699), .ZN(n5322) );
  NAND3_X1 U4631 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5322), .ZN(n5714) );
  NOR2_X1 U4632 ( .A1(n5714), .A2(n3671), .ZN(n5875) );
  INV_X1 U4633 ( .A(n5661), .ZN(n3672) );
  AND2_X1 U4634 ( .A1(n5875), .A2(n3672), .ZN(n5651) );
  AND2_X1 U4635 ( .A1(n5651), .A2(n3673), .ZN(n5631) );
  NAND3_X1 U4636 ( .A1(n5631), .A2(n3674), .A3(n4336), .ZN(n3676) );
  INV_X1 U4637 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6524) );
  NOR2_X1 U4638 ( .A1(n6192), .A2(n6524), .ZN(n4243) );
  INV_X1 U4639 ( .A(n4243), .ZN(n3675) );
  OAI211_X1 U4640 ( .C1(n5626), .C2(n4336), .A(n3676), .B(n3675), .ZN(n3677)
         );
  INV_X1 U4641 ( .A(n3677), .ZN(n3678) );
  NAND2_X1 U4642 ( .A1(n3680), .A2(n3013), .ZN(U2987) );
  INV_X1 U4643 ( .A(n4433), .ZN(n4574) );
  NAND2_X1 U4644 ( .A1(n4574), .A2(n3932), .ZN(n3682) );
  NAND2_X1 U4645 ( .A1(n6560), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3920) );
  NAND2_X1 U4646 ( .A1(n4429), .A2(n3932), .ZN(n3687) );
  AND2_X1 U4647 ( .A1(n5378), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3697) );
  NAND2_X1 U4648 ( .A1(n3697), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3685) );
  NOR2_X1 U4649 ( .A1(n5503), .A2(n6560), .ZN(n3683) );
  AOI22_X1 U4650 ( .A1(n3683), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6560), .ZN(n3684) );
  AND2_X1 U4651 ( .A1(n3685), .A2(n3684), .ZN(n3686) );
  NAND2_X1 U4652 ( .A1(n3687), .A2(n3686), .ZN(n4414) );
  INV_X1 U4653 ( .A(n3688), .ZN(n3689) );
  AOI21_X1 U4654 ( .B1(n4942), .B2(n3689), .A(n6560), .ZN(n4330) );
  OR2_X1 U4655 ( .A1(n3690), .A2(n3956), .ZN(n3694) );
  NAND2_X1 U4656 ( .A1(n3697), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4657 ( .A1(n3683), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6560), .ZN(n3691) );
  AND2_X1 U4658 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  NAND2_X1 U4659 ( .A1(n3694), .A2(n3693), .ZN(n4329) );
  NAND2_X1 U4660 ( .A1(n4330), .A2(n4329), .ZN(n4328) );
  INV_X1 U4661 ( .A(n4329), .ZN(n3695) );
  NOR2_X1 U4662 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3952) );
  NAND2_X1 U4663 ( .A1(n3695), .A2(n4188), .ZN(n3696) );
  NAND2_X1 U4664 ( .A1(n4328), .A2(n3696), .ZN(n4415) );
  INV_X1 U4665 ( .A(n3697), .ZN(n3717) );
  OAI21_X1 U4666 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3706), .ZN(n6190) );
  AOI22_X1 U4667 ( .A1(n4191), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4188), 
        .B2(n6190), .ZN(n3699) );
  NAND2_X1 U4668 ( .A1(n4187), .A2(EAX_REG_2__SCAN_IN), .ZN(n3698) );
  OAI211_X1 U4669 ( .C1(n3717), .C2(n5389), .A(n3699), .B(n3698), .ZN(n4409)
         );
  NAND2_X1 U4670 ( .A1(n4410), .A2(n4409), .ZN(n3703) );
  NAND2_X1 U4671 ( .A1(n3700), .A2(n3701), .ZN(n3702) );
  NAND2_X1 U4672 ( .A1(n6539), .A2(n3932), .ZN(n3713) );
  INV_X1 U4673 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4290) );
  INV_X1 U4674 ( .A(n3706), .ZN(n3705) );
  INV_X1 U4675 ( .A(n3719), .ZN(n3720) );
  INV_X1 U4676 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3707) );
  NAND2_X1 U4677 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  NAND2_X1 U4678 ( .A1(n3720), .A2(n3708), .ZN(n5370) );
  AOI22_X1 U4679 ( .A1(n5370), .A2(n4188), .B1(n4191), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3710) );
  NAND2_X1 U4680 ( .A1(n4187), .A2(EAX_REG_3__SCAN_IN), .ZN(n3709) );
  OAI211_X1 U4681 ( .C1(n3717), .C2(n4290), .A(n3710), .B(n3709), .ZN(n3711)
         );
  INV_X1 U4682 ( .A(n3711), .ZN(n3712) );
  NAND2_X1 U4683 ( .A1(n3713), .A2(n3712), .ZN(n4437) );
  NAND2_X1 U4684 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3716)
         );
  NAND2_X1 U4685 ( .A1(n4187), .A2(EAX_REG_4__SCAN_IN), .ZN(n3715) );
  OAI211_X1 U4686 ( .C1(n3717), .C2(n5905), .A(n3716), .B(n3715), .ZN(n3718)
         );
  NAND2_X1 U4687 ( .A1(n3718), .A2(n4165), .ZN(n3723) );
  INV_X1 U4688 ( .A(n3727), .ZN(n3729) );
  INV_X1 U4689 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U4690 ( .A1(n3720), .A2(n6019), .ZN(n3721) );
  NAND2_X1 U4691 ( .A1(n3729), .A2(n3721), .ZN(n6038) );
  NAND2_X1 U4692 ( .A1(n6038), .A2(n3952), .ZN(n3722) );
  NAND2_X1 U4693 ( .A1(n3723), .A2(n3722), .ZN(n3724) );
  NOR2_X2 U4694 ( .A1(n4443), .A2(n4442), .ZN(n4441) );
  INV_X1 U4695 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3734) );
  INV_X1 U4696 ( .A(n3735), .ZN(n3731) );
  INV_X1 U4697 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U4698 ( .A1(n3729), .A2(n3728), .ZN(n3730) );
  NAND2_X1 U4699 ( .A1(n3731), .A2(n3730), .ZN(n6017) );
  AOI22_X1 U4700 ( .A1(n6017), .A2(n3952), .B1(n4191), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U4701 ( .A1(n4441), .A2(n4554), .ZN(n4553) );
  INV_X1 U4702 ( .A(n4553), .ZN(n3741) );
  OAI21_X1 U4703 ( .B1(n3735), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3742), 
        .ZN(n5998) );
  INV_X1 U4704 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4790) );
  INV_X1 U4705 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3736) );
  OAI22_X1 U4706 ( .A1(n3870), .A2(n4790), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3736), .ZN(n3737) );
  MUX2_X1 U4707 ( .A(n5998), .B(n3737), .S(n4165), .Z(n3738) );
  NAND2_X1 U4708 ( .A1(n3741), .A2(n3740), .ZN(n4787) );
  INV_X1 U4709 ( .A(n4787), .ZN(n3749) );
  OAI21_X1 U4710 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3743), .A(n3764), 
        .ZN(n5992) );
  NAND2_X1 U4711 ( .A1(n5992), .A2(n4188), .ZN(n3745) );
  AOI22_X1 U4712 ( .A1(n4187), .A2(EAX_REG_7__SCAN_IN), .B1(n4191), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4713 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  NAND2_X1 U4714 ( .A1(n3749), .A2(n3748), .ZN(n5009) );
  XOR2_X1 U4715 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3764), .Z(n5062) );
  AOI22_X1 U4716 ( .A1(n4151), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4717 ( .A1(n4173), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4718 ( .A1(n3994), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4719 ( .A1(n4150), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3750) );
  NAND4_X1 U4720 ( .A1(n3753), .A2(n3752), .A3(n3751), .A4(n3750), .ZN(n3759)
         );
  AOI22_X1 U4721 ( .A1(n3856), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4722 ( .A1(n4096), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4723 ( .A1(n2992), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4724 ( .A1(n4172), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4725 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3758)
         );
  NOR2_X1 U4726 ( .A1(n3759), .A2(n3758), .ZN(n3762) );
  NAND2_X1 U4727 ( .A1(n4187), .A2(EAX_REG_8__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U4728 ( .A1(n4191), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3760)
         );
  OAI211_X1 U4729 ( .C1(n3956), .C2(n3762), .A(n3761), .B(n3760), .ZN(n3763)
         );
  AOI21_X1 U4730 ( .B1(n5062), .B2(n3952), .A(n3763), .ZN(n5041) );
  NOR2_X2 U4731 ( .A1(n5009), .A2(n5041), .ZN(n5040) );
  XNOR2_X1 U4732 ( .A(n3777), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5087) );
  AOI22_X1 U4733 ( .A1(n3683), .A2(EAX_REG_9__SCAN_IN), .B1(n4191), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4734 ( .A1(n4173), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4735 ( .A1(n2991), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4736 ( .A1(n4057), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4737 ( .A1(n3156), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3765) );
  NAND4_X1 U4738 ( .A1(n3768), .A2(n3767), .A3(n3766), .A4(n3765), .ZN(n3774)
         );
  AOI22_X1 U4739 ( .A1(n3856), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4740 ( .A1(n4151), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4741 ( .A1(n4150), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4742 ( .A1(n2992), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3769) );
  NAND4_X1 U4743 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3773)
         );
  OAI21_X1 U4744 ( .B1(n3774), .B2(n3773), .A(n3932), .ZN(n3775) );
  OAI211_X1 U4745 ( .C1(n5087), .C2(n4165), .A(n3776), .B(n3775), .ZN(n5070)
         );
  NAND2_X1 U4746 ( .A1(n5040), .A2(n5070), .ZN(n5068) );
  XOR2_X1 U4747 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3801), .Z(n5131) );
  AOI22_X1 U4748 ( .A1(n4096), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4749 ( .A1(n3994), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4750 ( .A1(n3856), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4751 ( .A1(n4172), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4752 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3787)
         );
  AOI22_X1 U4753 ( .A1(n4151), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4754 ( .A1(n4057), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4755 ( .A1(n3988), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4756 ( .A1(n4173), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3782) );
  NAND4_X1 U4757 ( .A1(n3785), .A2(n3784), .A3(n3783), .A4(n3782), .ZN(n3786)
         );
  OR2_X1 U4758 ( .A1(n3787), .A2(n3786), .ZN(n3788) );
  AOI22_X1 U4759 ( .A1(n3932), .A2(n3788), .B1(n4191), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3790) );
  NAND2_X1 U4760 ( .A1(n3683), .A2(EAX_REG_10__SCAN_IN), .ZN(n3789) );
  OAI211_X1 U4761 ( .C1(n5131), .C2(n4165), .A(n3790), .B(n3789), .ZN(n5118)
         );
  NOR2_X2 U4762 ( .A1(n5068), .A2(n5119), .ZN(n5136) );
  AOI22_X1 U4763 ( .A1(n3994), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4764 ( .A1(n4151), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4765 ( .A1(n4172), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4766 ( .A1(n2992), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4767 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3800)
         );
  AOI22_X1 U4768 ( .A1(n3856), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4769 ( .A1(n4173), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4770 ( .A1(n4174), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4771 ( .A1(n4057), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4772 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3799)
         );
  NOR2_X1 U4773 ( .A1(n3800), .A2(n3799), .ZN(n3804) );
  XNOR2_X1 U4774 ( .A(n3805), .B(n5142), .ZN(n5203) );
  NAND2_X1 U4775 ( .A1(n5203), .A2(n3952), .ZN(n3803) );
  AOI22_X1 U4776 ( .A1(n3683), .A2(EAX_REG_11__SCAN_IN), .B1(n4191), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3802) );
  OAI211_X1 U4777 ( .C1(n3804), .C2(n3956), .A(n3803), .B(n3802), .ZN(n5135)
         );
  NAND2_X1 U4778 ( .A1(n5136), .A2(n5135), .ZN(n5134) );
  INV_X1 U4779 ( .A(n5134), .ZN(n3821) );
  XOR2_X1 U4780 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3822), .Z(n5976) );
  INV_X1 U4781 ( .A(n5976), .ZN(n5232) );
  AOI22_X1 U4782 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3856), .B1(n3994), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4783 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n2992), .B1(n4144), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4784 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n2991), .B1(n4174), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4785 ( .A1(n4150), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4786 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3815)
         );
  AOI22_X1 U4787 ( .A1(n4151), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4788 ( .A1(n4172), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4789 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4096), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4790 ( .A1(n4173), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3810) );
  NAND4_X1 U4791 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3814)
         );
  NOR2_X1 U4792 ( .A1(n3815), .A2(n3814), .ZN(n3818) );
  NAND2_X1 U4793 ( .A1(n3683), .A2(EAX_REG_12__SCAN_IN), .ZN(n3817) );
  NAND2_X1 U4794 ( .A1(n4191), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3816)
         );
  OAI211_X1 U4795 ( .C1(n3956), .C2(n3818), .A(n3817), .B(n3816), .ZN(n3819)
         );
  AOI21_X1 U4796 ( .B1(n5232), .B2(n3952), .A(n3819), .ZN(n5227) );
  NAND2_X1 U4797 ( .A1(n3821), .A2(n3820), .ZN(n3962) );
  NAND2_X1 U4798 ( .A1(n3822), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3850)
         );
  INV_X1 U4799 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5284) );
  XNOR2_X1 U4800 ( .A(n3850), .B(n5284), .ZN(n5286) );
  NAND2_X1 U4801 ( .A1(n5286), .A2(n3952), .ZN(n3825) );
  NOR2_X1 U4802 ( .A1(n3920), .A2(n5284), .ZN(n3823) );
  AOI21_X1 U4803 ( .B1(n4187), .B2(EAX_REG_13__SCAN_IN), .A(n3823), .ZN(n3824)
         );
  NAND2_X1 U4804 ( .A1(n3825), .A2(n3824), .ZN(n5301) );
  AOI22_X1 U4805 ( .A1(n4151), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4806 ( .A1(n4172), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4807 ( .A1(n3994), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4808 ( .A1(n4057), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3826) );
  NAND4_X1 U4809 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3835)
         );
  AOI22_X1 U4810 ( .A1(n4096), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4811 ( .A1(n2992), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4812 ( .A1(n4173), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4813 ( .A1(n3856), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4814 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3834)
         );
  OR2_X1 U4815 ( .A1(n3835), .A2(n3834), .ZN(n3836) );
  AND2_X1 U4816 ( .A1(n3932), .A2(n3836), .ZN(n5299) );
  AOI22_X1 U4817 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4151), .B1(n2991), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4818 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4144), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4819 ( .A1(n3994), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4820 ( .A1(n4057), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4821 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3846)
         );
  AOI22_X1 U4822 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4096), .B1(n4150), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4823 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n2992), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4824 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4173), .B1(n3156), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4825 ( .A1(n3856), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3841) );
  NAND4_X1 U4826 ( .A1(n3844), .A2(n3843), .A3(n3842), .A4(n3841), .ZN(n3845)
         );
  NOR2_X1 U4827 ( .A1(n3846), .A2(n3845), .ZN(n3849) );
  INV_X1 U4828 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5796) );
  AOI21_X1 U4829 ( .B1(n5796), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3847) );
  AOI21_X1 U4830 ( .B1(n4187), .B2(EAX_REG_20__SCAN_IN), .A(n3847), .ZN(n3848)
         );
  OAI21_X1 U4831 ( .B1(n4162), .B2(n3849), .A(n3848), .ZN(n3853) );
  INV_X1 U4832 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6621) );
  INV_X1 U4833 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3851) );
  XNOR2_X1 U4834 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3982), .ZN(n5800)
         );
  NAND2_X1 U4835 ( .A1(n4188), .A2(n5800), .ZN(n3852) );
  NAND2_X1 U4836 ( .A1(n3853), .A2(n3852), .ZN(n5475) );
  INV_X1 U4837 ( .A(n5475), .ZN(n3960) );
  OR2_X1 U4838 ( .A1(n3854), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3855)
         );
  NAND2_X1 U4839 ( .A1(n3855), .A2(n3982), .ZN(n5866) );
  AOI22_X1 U4840 ( .A1(n3856), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4841 ( .A1(n4096), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4842 ( .A1(n4151), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4843 ( .A1(n4144), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4844 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3866)
         );
  AOI22_X1 U4845 ( .A1(n2991), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4846 ( .A1(n3988), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4847 ( .A1(n4173), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4848 ( .A1(n4150), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4849 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3865)
         );
  NOR2_X1 U4850 ( .A1(n3866), .A2(n3865), .ZN(n3867) );
  NOR2_X1 U4851 ( .A1(n4162), .A2(n3867), .ZN(n3872) );
  INV_X1 U4852 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4853 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3868)
         );
  OAI211_X1 U4854 ( .C1(n3870), .C2(n3869), .A(n4165), .B(n3868), .ZN(n3871)
         );
  OAI22_X1 U4855 ( .A1(n5866), .A2(n4165), .B1(n3872), .B2(n3871), .ZN(n5307)
         );
  INV_X1 U4856 ( .A(n5307), .ZN(n3959) );
  AOI22_X1 U4857 ( .A1(n4057), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4858 ( .A1(n2991), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4859 ( .A1(n3856), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4860 ( .A1(n4173), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4861 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3882)
         );
  AOI22_X1 U4862 ( .A1(n4096), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4863 ( .A1(n3994), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4864 ( .A1(n4150), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4865 ( .A1(n4151), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4866 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3881)
         );
  NOR2_X1 U4867 ( .A1(n3882), .A2(n3881), .ZN(n3886) );
  NAND2_X1 U4868 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3883)
         );
  NAND2_X1 U4869 ( .A1(n4165), .A2(n3883), .ZN(n3884) );
  AOI21_X1 U4870 ( .B1(n4187), .B2(EAX_REG_18__SCAN_IN), .A(n3884), .ZN(n3885)
         );
  OAI21_X1 U4871 ( .B1(n4162), .B2(n3886), .A(n3885), .ZN(n3888) );
  XNOR2_X1 U4872 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3902), .ZN(n5603)
         );
  NAND2_X1 U4873 ( .A1(n3952), .A2(n5603), .ZN(n3887) );
  NAND2_X1 U4874 ( .A1(n3888), .A2(n3887), .ZN(n5343) );
  INV_X1 U4875 ( .A(n5343), .ZN(n3958) );
  AOI22_X1 U4876 ( .A1(n4173), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4877 ( .A1(n3994), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4878 ( .A1(n2991), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4879 ( .A1(n4057), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4880 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3898)
         );
  AOI22_X1 U4881 ( .A1(n4096), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4882 ( .A1(n4151), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4883 ( .A1(n3856), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4884 ( .A1(n3988), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4885 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  NOR2_X1 U4886 ( .A1(n3898), .A2(n3897), .ZN(n3899) );
  OR2_X1 U4887 ( .A1(n4162), .A2(n3899), .ZN(n3906) );
  NAND2_X1 U4888 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3900)
         );
  NAND2_X1 U4889 ( .A1(n4165), .A2(n3900), .ZN(n3901) );
  AOI21_X1 U4890 ( .B1(n4187), .B2(EAX_REG_17__SCAN_IN), .A(n3901), .ZN(n3905)
         );
  OAI21_X1 U4891 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3903), .A(n3902), 
        .ZN(n5947) );
  NOR2_X1 U4892 ( .A1(n5947), .A2(n4165), .ZN(n3904) );
  AOI21_X1 U4893 ( .B1(n3906), .B2(n3905), .A(n3904), .ZN(n5487) );
  AOI22_X1 U4894 ( .A1(n4151), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4895 ( .A1(n4173), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4896 ( .A1(n4096), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4897 ( .A1(n4057), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3907) );
  NAND4_X1 U4898 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3916)
         );
  AOI22_X1 U4899 ( .A1(n4172), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4900 ( .A1(n3856), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4901 ( .A1(n3994), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4902 ( .A1(n2992), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3911) );
  NAND4_X1 U4903 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3915)
         );
  NOR2_X1 U4904 ( .A1(n3916), .A2(n3915), .ZN(n3917) );
  OR2_X1 U4905 ( .A1(n4162), .A2(n3917), .ZN(n3923) );
  INV_X1 U4906 ( .A(n3918), .ZN(n3919) );
  XNOR2_X1 U4907 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3919), .ZN(n5953)
         );
  INV_X1 U4908 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5609) );
  OAI22_X1 U4909 ( .A1(n5953), .A2(n4165), .B1(n3920), .B2(n5609), .ZN(n3921)
         );
  AOI21_X1 U4910 ( .B1(n4187), .B2(EAX_REG_16__SCAN_IN), .A(n3921), .ZN(n3922)
         );
  AND2_X1 U4911 ( .A1(n3923), .A2(n3922), .ZN(n5492) );
  AOI22_X1 U4912 ( .A1(n4173), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4913 ( .A1(n3994), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4914 ( .A1(n4150), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4915 ( .A1(n4151), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3924) );
  NAND4_X1 U4916 ( .A1(n3927), .A2(n3926), .A3(n3925), .A4(n3924), .ZN(n3934)
         );
  AOI22_X1 U4917 ( .A1(n3856), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4918 ( .A1(n4172), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4919 ( .A1(n4096), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4920 ( .A1(n2992), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U4921 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3933)
         );
  OAI21_X1 U4922 ( .B1(n3934), .B2(n3933), .A(n3932), .ZN(n3937) );
  XNOR2_X1 U4923 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3949), .ZN(n5620)
         );
  AOI22_X1 U4924 ( .A1(n4191), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n3952), 
        .B2(n5620), .ZN(n3936) );
  NAND2_X1 U4925 ( .A1(n4187), .A2(EAX_REG_15__SCAN_IN), .ZN(n3935) );
  AND3_X1 U4926 ( .A1(n3937), .A2(n3936), .A3(n3935), .ZN(n5437) );
  NOR2_X1 U4927 ( .A1(n5492), .A2(n5437), .ZN(n5485) );
  AND2_X1 U4928 ( .A1(n5487), .A2(n5485), .ZN(n3957) );
  AOI22_X1 U4929 ( .A1(n4096), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4930 ( .A1(n4151), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4931 ( .A1(n4057), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4932 ( .A1(n4150), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3938) );
  NAND4_X1 U4933 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3947)
         );
  AOI22_X1 U4934 ( .A1(n3994), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4935 ( .A1(n3856), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4936 ( .A1(n4173), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4937 ( .A1(n3988), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4938 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3946)
         );
  NOR2_X1 U4939 ( .A1(n3947), .A2(n3946), .ZN(n3955) );
  INV_X1 U4940 ( .A(n3948), .ZN(n3951) );
  INV_X1 U4941 ( .A(n3949), .ZN(n3950) );
  OAI21_X1 U4942 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n3951), .A(n3950), 
        .ZN(n5966) );
  AOI22_X1 U4943 ( .A1(n3952), .A2(n5966), .B1(n4191), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3954) );
  NAND2_X1 U4944 ( .A1(n4187), .A2(EAX_REG_14__SCAN_IN), .ZN(n3953) );
  OAI211_X1 U4945 ( .C1(n3956), .C2(n3955), .A(n3954), .B(n3953), .ZN(n5483)
         );
  NAND2_X1 U4946 ( .A1(n5273), .A2(n3961), .ZN(n3968) );
  INV_X1 U4947 ( .A(n3963), .ZN(n3965) );
  INV_X1 U4948 ( .A(n5301), .ZN(n3964) );
  NOR2_X1 U4949 ( .A1(n3965), .A2(n3964), .ZN(n3966) );
  NAND2_X1 U4950 ( .A1(n5302), .A2(n3966), .ZN(n3967) );
  AOI22_X1 U4951 ( .A1(n4151), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4952 ( .A1(n4096), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4953 ( .A1(n3994), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4954 ( .A1(n4172), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3969) );
  NAND4_X1 U4955 ( .A1(n3972), .A2(n3971), .A3(n3970), .A4(n3969), .ZN(n3978)
         );
  AOI22_X1 U4956 ( .A1(n3856), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4957 ( .A1(n4057), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4958 ( .A1(n3988), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4959 ( .A1(n4173), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3973) );
  NAND4_X1 U4960 ( .A1(n3976), .A2(n3975), .A3(n3974), .A4(n3973), .ZN(n3977)
         );
  NOR2_X1 U4961 ( .A1(n3978), .A2(n3977), .ZN(n3979) );
  OR2_X1 U4962 ( .A1(n4162), .A2(n3979), .ZN(n3987) );
  INV_X1 U4963 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6561) );
  OAI21_X1 U4964 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6561), .A(n6560), 
        .ZN(n3980) );
  INV_X1 U4965 ( .A(n3980), .ZN(n3981) );
  AOI21_X1 U4966 ( .B1(n4187), .B2(EAX_REG_21__SCAN_IN), .A(n3981), .ZN(n3986)
         );
  OAI21_X1 U4967 ( .B1(n3984), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4033), 
        .ZN(n5794) );
  NOR2_X1 U4968 ( .A1(n5794), .A2(n4165), .ZN(n3985) );
  AOI21_X1 U4969 ( .B1(n3987), .B2(n3986), .A(n3985), .ZN(n5292) );
  NAND2_X1 U4970 ( .A1(n5293), .A2(n5292), .ZN(n5291) );
  INV_X1 U4971 ( .A(n5291), .ZN(n4008) );
  AOI22_X1 U4972 ( .A1(n4096), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4973 ( .A1(n4151), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4974 ( .A1(n4057), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4975 ( .A1(n3856), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3990) );
  NAND4_X1 U4976 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n4001)
         );
  AOI22_X1 U4977 ( .A1(n3994), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4978 ( .A1(n2991), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4979 ( .A1(n4172), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4980 ( .A1(n4174), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3996) );
  NAND4_X1 U4981 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n4000)
         );
  NOR2_X1 U4982 ( .A1(n4001), .A2(n4000), .ZN(n4004) );
  INV_X1 U4983 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5579) );
  OAI21_X1 U4984 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5579), .A(n4165), .ZN(
        n4002) );
  AOI21_X1 U4985 ( .B1(n4187), .B2(EAX_REG_22__SCAN_IN), .A(n4002), .ZN(n4003)
         );
  OAI21_X1 U4986 ( .B1(n4162), .B2(n4004), .A(n4003), .ZN(n4006) );
  XNOR2_X1 U4987 ( .A(n4033), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5780)
         );
  NAND2_X1 U4988 ( .A1(n5780), .A2(n4188), .ZN(n4005) );
  NAND2_X1 U4989 ( .A1(n4006), .A2(n4005), .ZN(n5331) );
  NAND2_X1 U4990 ( .A1(n4008), .A2(n4007), .ZN(n5330) );
  AOI22_X1 U4991 ( .A1(n2991), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4992 ( .A1(n4096), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4993 ( .A1(n4174), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4994 ( .A1(n4144), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4009) );
  NAND4_X1 U4995 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(n4018)
         );
  AOI22_X1 U4996 ( .A1(n3094), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4997 ( .A1(n4173), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4998 ( .A1(n4151), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4999 ( .A1(n4150), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4013) );
  NAND4_X1 U5000 ( .A1(n4016), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(n4017)
         );
  NOR2_X1 U5001 ( .A1(n4018), .A2(n4017), .ZN(n4039) );
  AOI22_X1 U5002 ( .A1(n3094), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4096), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U5003 ( .A1(n4173), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3994), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U5004 ( .A1(n4150), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U5005 ( .A1(n4144), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4019) );
  NAND4_X1 U5006 ( .A1(n4022), .A2(n4021), .A3(n4020), .A4(n4019), .ZN(n4028)
         );
  AOI22_X1 U5007 ( .A1(n4151), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U5008 ( .A1(n4057), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5009 ( .A1(n3156), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5010 ( .A1(n2992), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U5011 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4027)
         );
  NOR2_X1 U5012 ( .A1(n4028), .A2(n4027), .ZN(n4040) );
  XNOR2_X1 U5013 ( .A(n4039), .B(n4040), .ZN(n4032) );
  NAND2_X1 U5014 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4029)
         );
  NAND2_X1 U5015 ( .A1(n4165), .A2(n4029), .ZN(n4030) );
  AOI21_X1 U5016 ( .B1(n4187), .B2(EAX_REG_23__SCAN_IN), .A(n4030), .ZN(n4031)
         );
  OAI21_X1 U5017 ( .B1(n4162), .B2(n4032), .A(n4031), .ZN(n4038) );
  NOR2_X1 U5018 ( .A1(n4034), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4035)
         );
  OR2_X1 U5019 ( .A1(n4072), .A2(n4035), .ZN(n5572) );
  INV_X1 U5020 ( .A(n5572), .ZN(n4036) );
  NAND2_X1 U5021 ( .A1(n4036), .A2(n4188), .ZN(n4037) );
  NAND2_X1 U5022 ( .A1(n4038), .A2(n4037), .ZN(n5424) );
  NOR2_X2 U5023 ( .A1(n5330), .A2(n5424), .ZN(n5422) );
  INV_X1 U5024 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5562) );
  XNOR2_X1 U5025 ( .A(n4072), .B(n5562), .ZN(n5770) );
  NOR2_X1 U5026 ( .A1(n4040), .A2(n4039), .ZN(n4056) );
  AOI22_X1 U5027 ( .A1(n4151), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5028 ( .A1(n4172), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5029 ( .A1(n3994), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5030 ( .A1(n4057), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U5031 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4050)
         );
  AOI22_X1 U5032 ( .A1(n4096), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5033 ( .A1(n2992), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5034 ( .A1(n4173), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5035 ( .A1(n3094), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U5036 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4049)
         );
  OR2_X1 U5037 ( .A1(n4050), .A2(n4049), .ZN(n4055) );
  INV_X1 U5038 ( .A(n4055), .ZN(n4051) );
  XNOR2_X1 U5039 ( .A(n4056), .B(n4051), .ZN(n4052) );
  INV_X1 U5040 ( .A(n4162), .ZN(n4184) );
  NAND2_X1 U5041 ( .A1(n4052), .A2(n4184), .ZN(n4054) );
  AOI22_X1 U5042 ( .A1(n3683), .A2(EAX_REG_24__SCAN_IN), .B1(n4191), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4053) );
  OAI211_X1 U5043 ( .C1(n5770), .C2(n4165), .A(n4054), .B(n4053), .ZN(n5472)
         );
  NAND2_X1 U5044 ( .A1(n5422), .A2(n5472), .ZN(n5464) );
  NAND2_X1 U5045 ( .A1(n4056), .A2(n4055), .ZN(n4078) );
  AOI22_X1 U5046 ( .A1(n4096), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5047 ( .A1(n4173), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5048 ( .A1(n4172), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5049 ( .A1(n4150), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U5050 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4067)
         );
  AOI22_X1 U5051 ( .A1(n4151), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5052 ( .A1(n3094), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5053 ( .A1(n3994), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5054 ( .A1(n4174), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5055 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4066)
         );
  NOR2_X1 U5056 ( .A1(n4067), .A2(n4066), .ZN(n4079) );
  XNOR2_X1 U5057 ( .A(n4078), .B(n4079), .ZN(n4071) );
  NAND2_X1 U5058 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4068)
         );
  NAND2_X1 U5059 ( .A1(n4165), .A2(n4068), .ZN(n4069) );
  AOI21_X1 U5060 ( .B1(n4187), .B2(EAX_REG_25__SCAN_IN), .A(n4069), .ZN(n4070)
         );
  OAI21_X1 U5061 ( .B1(n4071), .B2(n4162), .A(n4070), .ZN(n4077) );
  OR2_X1 U5062 ( .A1(n4073), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4074)
         );
  NAND2_X1 U5063 ( .A1(n4074), .A2(n4113), .ZN(n5860) );
  INV_X1 U5064 ( .A(n5860), .ZN(n4075) );
  NAND2_X1 U5065 ( .A1(n4075), .A2(n4188), .ZN(n4076) );
  NAND2_X1 U5066 ( .A1(n4077), .A2(n4076), .ZN(n5466) );
  NOR2_X2 U5067 ( .A1(n5464), .A2(n5466), .ZN(n5457) );
  NOR2_X1 U5068 ( .A1(n4079), .A2(n4078), .ZN(n4108) );
  AOI22_X1 U5069 ( .A1(n4151), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5070 ( .A1(n4172), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5071 ( .A1(n3994), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5072 ( .A1(n4057), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4080) );
  NAND4_X1 U5073 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4089)
         );
  AOI22_X1 U5074 ( .A1(n4096), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5075 ( .A1(n2992), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5076 ( .A1(n4173), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5077 ( .A1(n3094), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4084) );
  NAND4_X1 U5078 ( .A1(n4087), .A2(n4086), .A3(n4085), .A4(n4084), .ZN(n4088)
         );
  OR2_X1 U5079 ( .A1(n4089), .A2(n4088), .ZN(n4107) );
  XNOR2_X1 U5080 ( .A(n4108), .B(n4107), .ZN(n4092) );
  INV_X1 U5081 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5757) );
  AOI21_X1 U5082 ( .B1(n5757), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4090) );
  AOI21_X1 U5083 ( .B1(n4187), .B2(EAX_REG_26__SCAN_IN), .A(n4090), .ZN(n4091)
         );
  OAI21_X1 U5084 ( .B1(n4092), .B2(n4162), .A(n4091), .ZN(n4094) );
  XNOR2_X1 U5085 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4113), .ZN(n5748)
         );
  NAND2_X1 U5086 ( .A1(n5748), .A2(n4188), .ZN(n4093) );
  NAND2_X1 U5087 ( .A1(n4094), .A2(n4093), .ZN(n5460) );
  AOI22_X1 U5088 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4173), .B1(n4096), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5089 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n2991), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5090 ( .A1(n4150), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5091 ( .A1(n4144), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4097) );
  NAND4_X1 U5092 ( .A1(n4100), .A2(n4099), .A3(n4098), .A4(n4097), .ZN(n4106)
         );
  AOI22_X1 U5093 ( .A1(n4151), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5094 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3856), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5095 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n2992), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5096 ( .A1(n3994), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4101) );
  NAND4_X1 U5097 ( .A1(n4104), .A2(n4103), .A3(n4102), .A4(n4101), .ZN(n4105)
         );
  NOR2_X1 U5098 ( .A1(n4106), .A2(n4105), .ZN(n4122) );
  NAND2_X1 U5099 ( .A1(n4108), .A2(n4107), .ZN(n4121) );
  XNOR2_X1 U5100 ( .A(n4122), .B(n4121), .ZN(n4112) );
  NAND2_X1 U5101 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4109)
         );
  NAND2_X1 U5102 ( .A1(n4165), .A2(n4109), .ZN(n4110) );
  AOI21_X1 U5103 ( .B1(n4187), .B2(EAX_REG_27__SCAN_IN), .A(n4110), .ZN(n4111)
         );
  OAI21_X1 U5104 ( .B1(n4112), .B2(n4162), .A(n4111), .ZN(n4120) );
  INV_X1 U5105 ( .A(n4113), .ZN(n4114) );
  INV_X1 U5106 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4117) );
  INV_X1 U5107 ( .A(n4115), .ZN(n4116) );
  NAND2_X1 U5108 ( .A1(n4117), .A2(n4116), .ZN(n4118) );
  NAND2_X1 U5109 ( .A1(n4140), .A2(n4118), .ZN(n5747) );
  NOR2_X1 U5110 ( .A1(n4122), .A2(n4121), .ZN(n4159) );
  AOI22_X1 U5111 ( .A1(n4151), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5112 ( .A1(n4172), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5113 ( .A1(n3051), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5114 ( .A1(n4057), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U5115 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4132)
         );
  AOI22_X1 U5116 ( .A1(n4096), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5117 ( .A1(n2992), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5118 ( .A1(n4173), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5119 ( .A1(n3094), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4127) );
  NAND4_X1 U5120 ( .A1(n4130), .A2(n4129), .A3(n4128), .A4(n4127), .ZN(n4131)
         );
  OR2_X1 U5121 ( .A1(n4132), .A2(n4131), .ZN(n4158) );
  INV_X1 U5122 ( .A(n4158), .ZN(n4133) );
  XNOR2_X1 U5123 ( .A(n4159), .B(n4133), .ZN(n4134) );
  NAND2_X1 U5124 ( .A1(n4134), .A2(n4184), .ZN(n4139) );
  NAND2_X1 U5125 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4135)
         );
  NAND2_X1 U5126 ( .A1(n4165), .A2(n4135), .ZN(n4136) );
  AOI21_X1 U5127 ( .B1(n4187), .B2(EAX_REG_28__SCAN_IN), .A(n4136), .ZN(n4138)
         );
  XNOR2_X1 U5128 ( .A(n4140), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5738)
         );
  AOI21_X1 U5129 ( .B1(n4139), .B2(n4138), .A(n4137), .ZN(n5449) );
  INV_X1 U5130 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U5131 ( .A1(n4141), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4199)
         );
  INV_X1 U5132 ( .A(n4141), .ZN(n4142) );
  INV_X1 U5133 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U5134 ( .A1(n4142), .A2(n5530), .ZN(n4143) );
  NAND2_X1 U5135 ( .A1(n4199), .A2(n4143), .ZN(n5529) );
  AOI22_X1 U5136 ( .A1(n4172), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5137 ( .A1(n3094), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5138 ( .A1(n3988), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5139 ( .A1(n3051), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4146) );
  NAND4_X1 U5140 ( .A1(n4149), .A2(n4148), .A3(n4147), .A4(n4146), .ZN(n4157)
         );
  AOI22_X1 U5141 ( .A1(n4096), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5142 ( .A1(n4151), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5143 ( .A1(n4173), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5144 ( .A1(n4057), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U5145 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4156)
         );
  NOR2_X1 U5146 ( .A1(n4157), .A2(n4156), .ZN(n4167) );
  NAND2_X1 U5147 ( .A1(n4159), .A2(n4158), .ZN(n4166) );
  XNOR2_X1 U5148 ( .A(n4167), .B(n4166), .ZN(n4163) );
  AOI21_X1 U5149 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6560), .A(n4188), 
        .ZN(n4161) );
  NAND2_X1 U5150 ( .A1(n4187), .A2(EAX_REG_29__SCAN_IN), .ZN(n4160) );
  OAI211_X1 U5151 ( .C1(n4163), .C2(n4162), .A(n4161), .B(n4160), .ZN(n4164)
         );
  OAI21_X1 U5152 ( .B1(n4165), .B2(n5529), .A(n4164), .ZN(n5413) );
  NOR2_X1 U5153 ( .A1(n4167), .A2(n4166), .ZN(n4183) );
  AOI22_X1 U5154 ( .A1(n4096), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5155 ( .A1(n2991), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4057), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5156 ( .A1(n3094), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3989), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5157 ( .A1(n4150), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4168) );
  NAND4_X1 U5158 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4181)
         );
  AOI22_X1 U5159 ( .A1(n4151), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5160 ( .A1(n4173), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3988), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5161 ( .A1(n3051), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5162 ( .A1(n4144), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4176) );
  NAND4_X1 U5163 ( .A1(n4179), .A2(n4178), .A3(n4177), .A4(n4176), .ZN(n4180)
         );
  NOR2_X1 U5164 ( .A1(n4181), .A2(n4180), .ZN(n4182) );
  XNOR2_X1 U5165 ( .A(n4183), .B(n4182), .ZN(n4185) );
  NAND2_X1 U5166 ( .A1(n4185), .A2(n4184), .ZN(n4190) );
  INV_X1 U5167 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5522) );
  NOR2_X1 U5168 ( .A1(n5522), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4186) );
  AOI211_X1 U5169 ( .C1(n4187), .C2(EAX_REG_30__SCAN_IN), .A(n4186), .B(n4188), 
        .ZN(n4189) );
  XNOR2_X1 U5170 ( .A(n4199), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5520)
         );
  AOI22_X1 U5171 ( .A1(n4190), .A2(n4189), .B1(n5520), .B2(n4188), .ZN(n5393)
         );
  NAND2_X1 U5172 ( .A1(n5412), .A2(n5393), .ZN(n4194) );
  AOI22_X1 U5173 ( .A1(n3683), .A2(EAX_REG_31__SCAN_IN), .B1(n4191), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4192) );
  XNOR2_X2 U5174 ( .A(n4194), .B(n4193), .ZN(n5377) );
  INV_X1 U5175 ( .A(n6436), .ZN(n6445) );
  INV_X1 U5176 ( .A(n4255), .ZN(n4261) );
  INV_X1 U5177 ( .A(n4195), .ZN(n4267) );
  AND2_X1 U5178 ( .A1(n4259), .A2(n4267), .ZN(n4254) );
  NAND2_X1 U5179 ( .A1(n4254), .A2(n6436), .ZN(n4252) );
  NOR2_X1 U5180 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6566) );
  NAND2_X1 U5181 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6566), .ZN(n6434) );
  NOR3_X1 U5182 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6449), .A3(n6441), .ZN(
        n6448) );
  NOR2_X1 U5183 ( .A1(n5592), .A2(n6448), .ZN(n4196) );
  OAI21_X1 U5184 ( .B1(n6434), .B2(n6562), .A(n4196), .ZN(n4197) );
  INV_X1 U5185 ( .A(n4197), .ZN(n4198) );
  INV_X1 U5186 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4209) );
  NOR2_X1 U5187 ( .A1(n4997), .A2(n6441), .ZN(n4201) );
  NAND2_X1 U5188 ( .A1(n5377), .A2(n6001), .ZN(n4220) );
  NAND2_X1 U5189 ( .A1(n6462), .A2(n6561), .ZN(n4992) );
  INV_X1 U5190 ( .A(n4992), .ZN(n4202) );
  NAND3_X1 U5191 ( .A1(n4203), .A2(n4202), .A3(n6065), .ZN(n4204) );
  INV_X1 U5192 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6520) );
  INV_X1 U5193 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6703) );
  INV_X1 U5194 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6513) );
  INV_X1 U5195 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6511) );
  NOR3_X1 U5196 ( .A1(n6703), .A2(n6513), .A3(n6511), .ZN(n4211) );
  NAND3_X1 U5197 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4206) );
  INV_X1 U5198 ( .A(n5987), .ZN(n5441) );
  INV_X1 U5199 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6484) );
  INV_X1 U5200 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6478) );
  NAND3_X1 U5201 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6025) );
  NOR2_X1 U5202 ( .A1(n6478), .A2(n6025), .ZN(n6008) );
  NAND2_X1 U5203 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6008), .ZN(n5986) );
  NAND2_X1 U5204 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5057) );
  NOR3_X1 U5205 ( .A1(n6484), .A2(n5986), .A3(n5057), .ZN(n5127) );
  NAND4_X1 U5206 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n5127), .ZN(n5974) );
  NAND2_X1 U5207 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n5281) );
  NOR2_X1 U5208 ( .A1(n5974), .A2(n5281), .ZN(n5962) );
  NAND2_X1 U5209 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5962), .ZN(n5960) );
  NAND3_X1 U5210 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n4205) );
  NOR3_X1 U5211 ( .A1(n5441), .A2(n5960), .A3(n4205), .ZN(n5810) );
  NAND4_X1 U5212 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5810), .ZN(n5774) );
  NOR2_X1 U5213 ( .A1(n4206), .A2(n5774), .ZN(n5425) );
  NOR2_X1 U5214 ( .A1(n5441), .A2(n6009), .ZN(n5811) );
  AOI21_X1 U5215 ( .B1(n4211), .B2(n5425), .A(n5811), .ZN(n5754) );
  AND2_X1 U5216 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4207) );
  NOR2_X1 U5217 ( .A1(n6026), .A2(n4207), .ZN(n4208) );
  OR2_X1 U5218 ( .A1(n5754), .A2(n4208), .ZN(n5415) );
  AOI21_X1 U5219 ( .B1(n6009), .B2(n6520), .A(n5415), .ZN(n5407) );
  OAI21_X1 U5220 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6026), .A(n5407), .ZN(n4214) );
  INV_X1 U5221 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5354) );
  OR2_X1 U5222 ( .A1(n6461), .A2(n4992), .ZN(n6401) );
  NAND2_X1 U5223 ( .A1(n3179), .A2(n6401), .ZN(n4994) );
  OAI22_X1 U5224 ( .A1(n6018), .A2(n4209), .B1(n4216), .B2(n4994), .ZN(n4213)
         );
  NAND4_X1 U5225 ( .A1(n5950), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(REIP_REG_15__SCAN_IN), .ZN(n5931) );
  NAND3_X1 U5226 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4210) );
  NOR2_X1 U5227 ( .A1(n5931), .A2(n4210), .ZN(n5776) );
  NAND4_X1 U5228 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5776), .ZN(n5763) );
  INV_X1 U5229 ( .A(n5763), .ZN(n5749) );
  NAND2_X1 U5230 ( .A1(n5749), .A2(n4211), .ZN(n5733) );
  INV_X1 U5231 ( .A(n5733), .ZN(n5743) );
  NAND3_X1 U5232 ( .A1(n5743), .A2(REIP_REG_27__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n5419) );
  INV_X1 U5233 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6522) );
  NOR4_X1 U5234 ( .A1(n5419), .A2(REIP_REG_31__SCAN_IN), .A3(n6522), .A4(n6520), .ZN(n4212) );
  AOI211_X1 U5235 ( .C1(REIP_REG_31__SCAN_IN), .C2(n4214), .A(n4213), .B(n4212), .ZN(n4219) );
  INV_X1 U5236 ( .A(n5355), .ZN(n4217) );
  NAND2_X1 U5237 ( .A1(n4366), .A2(n4992), .ZN(n4215) );
  NOR2_X2 U5238 ( .A1(n4216), .A2(n4215), .ZN(n6007) );
  NAND2_X1 U5239 ( .A1(n4217), .A2(n6007), .ZN(n4218) );
  NAND3_X1 U5240 ( .A1(n4220), .A2(n4219), .A3(n4218), .ZN(U2796) );
  BUF_X1 U5241 ( .A(n4221), .Z(n5710) );
  NAND2_X1 U5242 ( .A1(n5708), .A2(n5713), .ZN(n4222) );
  AOI22_X2 U5243 ( .A1(n5710), .A2(n4222), .B1(n4227), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5590) );
  XNOR2_X1 U5244 ( .A(n5708), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5591)
         );
  AOI22_X1 U5245 ( .A1(n5590), .A2(n5591), .B1(n5708), .B2(n4223), .ZN(n5585)
         );
  INV_X1 U5246 ( .A(n5585), .ZN(n4225) );
  XNOR2_X1 U5247 ( .A(n4227), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5584)
         );
  NOR2_X1 U5248 ( .A1(n5576), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5575)
         );
  NAND2_X1 U5249 ( .A1(n5583), .A2(n5575), .ZN(n5567) );
  NAND3_X1 U5250 ( .A1(n5576), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4228) );
  OAI21_X1 U5251 ( .B1(n4227), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n4226), 
        .ZN(n5578) );
  OAI22_X2 U5252 ( .A1(n5567), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n4228), .B2(n5578), .ZN(n4229) );
  XNOR2_X1 U5253 ( .A(n4229), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5566)
         );
  AND2_X1 U5254 ( .A1(n5429), .A2(n4230), .ZN(n4231) );
  OR2_X1 U5255 ( .A1(n4231), .A2(n5469), .ZN(n5773) );
  NAND2_X1 U5256 ( .A1(n5592), .A2(REIP_REG_24__SCAN_IN), .ZN(n5561) );
  OAI21_X1 U5257 ( .B1(n5773), .B2(n3628), .A(n5561), .ZN(n4232) );
  NOR2_X1 U5258 ( .A1(n5714), .A2(n4233), .ZN(n5678) );
  NAND3_X1 U5259 ( .A1(n5678), .A2(n5679), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4235) );
  OAI21_X1 U5260 ( .B1(n5566), .B2(n5717), .A(n4237), .ZN(U2994) );
  OR2_X2 U5261 ( .A1(n5731), .A2(n6424), .ZN(n6193) );
  NAND3_X1 U5262 ( .A1(n6562), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6453) );
  INV_X1 U5263 ( .A(n6453), .ZN(n4238) );
  NOR2_X1 U5264 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n4897) );
  NAND2_X1 U5265 ( .A1(n4238), .A2(n6536), .ZN(n6200) );
  NAND2_X1 U5266 ( .A1(n5377), .A2(n6186), .ZN(n4247) );
  INV_X1 U5267 ( .A(n4897), .ZN(n6343) );
  AND2_X1 U5268 ( .A1(n6343), .A2(n4239), .ZN(n6558) );
  OR2_X1 U5269 ( .A1(n6558), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4240) );
  NAND2_X1 U5270 ( .A1(n6562), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4242) );
  NAND2_X1 U5271 ( .A1(n6561), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4241) );
  NAND2_X1 U5272 ( .A1(n4242), .A2(n4241), .ZN(n6196) );
  AOI21_X1 U5273 ( .B1(n6197), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4243), 
        .ZN(n4244) );
  OAI21_X1 U5274 ( .B1(n6191), .B2(n4997), .A(n4244), .ZN(n4245) );
  INV_X1 U5275 ( .A(n4245), .ZN(n4246) );
  OAI211_X1 U5276 ( .C1(n4248), .C2(n6193), .A(n4247), .B(n4246), .ZN(U2955)
         );
  NAND2_X1 U5277 ( .A1(n4249), .A2(n3634), .ZN(n4258) );
  NOR2_X1 U5278 ( .A1(n6343), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5060) );
  OAI21_X1 U5279 ( .B1(n5060), .B2(READREQUEST_REG_SCAN_IN), .A(n6557), .ZN(
        n4250) );
  OAI21_X1 U5280 ( .B1(n6557), .B2(n4258), .A(n4250), .ZN(U3474) );
  INV_X1 U5281 ( .A(n4251), .ZN(n4270) );
  AOI211_X1 U5282 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4252), .A(n5060), .B(
        n4270), .ZN(n4253) );
  INV_X1 U5283 ( .A(n4253), .ZN(U2788) );
  INV_X1 U5284 ( .A(n6407), .ZN(n4257) );
  OAI22_X1 U5285 ( .A1(n4257), .A2(n4256), .B1(n4255), .B2(n4254), .ZN(n5908)
         );
  AOI21_X1 U5286 ( .B1(n4258), .B2(n6461), .A(READY_N), .ZN(n6564) );
  NOR2_X1 U5287 ( .A1(n5908), .A2(n6564), .ZN(n6427) );
  NOR2_X1 U5288 ( .A1(n6427), .A2(n6445), .ZN(n5914) );
  INV_X1 U5289 ( .A(MORE_REG_SCAN_IN), .ZN(n4269) );
  INV_X1 U5290 ( .A(n4259), .ZN(n4266) );
  INV_X1 U5291 ( .A(n4298), .ZN(n4260) );
  OR2_X1 U5292 ( .A1(n4260), .A2(n6407), .ZN(n4265) );
  NAND2_X1 U5293 ( .A1(n4262), .A2(n4261), .ZN(n4263) );
  NAND2_X1 U5294 ( .A1(n6407), .A2(n4263), .ZN(n4264) );
  OAI211_X1 U5295 ( .C1(n4267), .C2(n4266), .A(n4265), .B(n4264), .ZN(n6426)
         );
  NAND2_X1 U5296 ( .A1(n5914), .A2(n6426), .ZN(n4268) );
  OAI21_X1 U5297 ( .B1(n5914), .B2(n4269), .A(n4268), .ZN(U3471) );
  OAI21_X1 U5298 ( .B1(n3179), .B2(n6462), .A(n4270), .ZN(n6110) );
  INV_X1 U5299 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6724) );
  INV_X1 U5300 ( .A(n5731), .ZN(n4271) );
  INV_X1 U5301 ( .A(n6402), .ZN(n5728) );
  NAND2_X2 U5302 ( .A1(n4271), .A2(n5728), .ZN(n6180) );
  INV_X1 U5303 ( .A(n6180), .ZN(n4277) );
  NAND2_X1 U5304 ( .A1(n4277), .A2(EAX_REG_7__SCAN_IN), .ZN(n4272) );
  INV_X1 U5305 ( .A(n6140), .ZN(n6177) );
  NAND2_X1 U5306 ( .A1(n6177), .A2(DATAI_7_), .ZN(n4273) );
  OAI211_X1 U5307 ( .C1(n6115), .C2(n6724), .A(n4272), .B(n4273), .ZN(U2946)
         );
  INV_X1 U5308 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U5309 ( .A1(n4277), .A2(EAX_REG_23__SCAN_IN), .ZN(n4274) );
  OAI211_X1 U5310 ( .C1(n6115), .C2(n6742), .A(n4274), .B(n4273), .ZN(U2931)
         );
  INV_X1 U5311 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6675) );
  INV_X1 U5312 ( .A(DATAI_12_), .ZN(n4275) );
  NOR2_X1 U5313 ( .A1(n6140), .A2(n4275), .ZN(n6134) );
  AOI21_X1 U5314 ( .B1(EAX_REG_12__SCAN_IN), .B2(n4277), .A(n6134), .ZN(n4276)
         );
  OAI21_X1 U5315 ( .B1(n6115), .B2(n6675), .A(n4276), .ZN(U2951) );
  INV_X1 U5316 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6659) );
  AND2_X1 U5317 ( .A1(n6177), .A2(DATAI_3_), .ZN(n6113) );
  AOI21_X1 U5318 ( .B1(EAX_REG_3__SCAN_IN), .B2(n4277), .A(n6113), .ZN(n4278)
         );
  OAI21_X1 U5319 ( .B1(n6115), .B2(n6659), .A(n4278), .ZN(U2942) );
  INV_X1 U5320 ( .A(n4308), .ZN(n4282) );
  NAND3_X1 U5321 ( .A1(n4282), .A2(n4281), .A3(n4280), .ZN(n4283) );
  NOR2_X1 U5322 ( .A1(n4284), .A2(n4283), .ZN(n4285) );
  AND2_X1 U5323 ( .A1(n4285), .A2(n4303), .ZN(n4376) );
  XNOR2_X1 U5324 ( .A(n4286), .B(n4290), .ZN(n4289) );
  INV_X1 U5325 ( .A(n4380), .ZN(n4288) );
  INV_X1 U5326 ( .A(n4377), .ZN(n5388) );
  OAI21_X1 U5327 ( .B1(n5388), .B2(n5389), .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .ZN(n4287) );
  NAND2_X1 U5328 ( .A1(n3202), .A2(n4287), .ZN(n4297) );
  AOI22_X1 U5329 ( .A1(n5729), .A2(n4289), .B1(n4288), .B2(n4297), .ZN(n4296)
         );
  MUX2_X1 U5330 ( .A(n4291), .B(n4290), .S(n4377), .Z(n4293) );
  INV_X1 U5331 ( .A(n4302), .ZN(n4292) );
  OR2_X1 U5332 ( .A1(n4298), .A2(n4292), .ZN(n4383) );
  OAI21_X1 U5333 ( .B1(n4294), .B2(n4293), .A(n4383), .ZN(n4295) );
  OAI211_X1 U5334 ( .C1(n6254), .C2(n4376), .A(n4296), .B(n4295), .ZN(n4388)
         );
  INV_X1 U5335 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6718) );
  AOI22_X1 U5336 ( .A1(n4388), .A2(n5902), .B1(n5387), .B2(n4297), .ZN(n4317)
         );
  NAND2_X1 U5337 ( .A1(n6407), .A2(n4298), .ZN(n4326) );
  INV_X1 U5338 ( .A(n4299), .ZN(n4301) );
  NAND3_X1 U5339 ( .A1(n4326), .A2(n4301), .A3(n4300), .ZN(n4314) );
  OR2_X1 U5340 ( .A1(n6407), .A2(n4302), .ZN(n4306) );
  INV_X1 U5341 ( .A(n4303), .ZN(n5903) );
  NAND2_X1 U5342 ( .A1(n5903), .A2(n4304), .ZN(n4305) );
  NAND2_X1 U5343 ( .A1(n4306), .A2(n4305), .ZN(n4358) );
  INV_X1 U5344 ( .A(n6461), .ZN(n4307) );
  OAI21_X1 U5345 ( .B1(n5729), .B2(n4308), .A(n4307), .ZN(n4310) );
  NAND2_X1 U5346 ( .A1(n4310), .A2(n4309), .ZN(n4311) );
  NAND2_X1 U5347 ( .A1(n4311), .A2(n6462), .ZN(n4312) );
  NOR2_X1 U5348 ( .A1(n4312), .A2(n6407), .ZN(n4313) );
  INV_X1 U5349 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5913) );
  NAND2_X1 U5350 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n5732) );
  INV_X1 U5351 ( .A(n5732), .ZN(n4403) );
  NAND2_X1 U5352 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4403), .ZN(n6532) );
  NOR2_X1 U5353 ( .A1(n5913), .A2(n6532), .ZN(n4315) );
  AOI21_X1 U5354 ( .B1(n4391), .B2(n6436), .A(n4315), .ZN(n5900) );
  OAI21_X1 U5355 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6718), .A(n5900), .ZN(
        n5906) );
  INV_X1 U5356 ( .A(n5906), .ZN(n5391) );
  NAND2_X1 U5357 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n5391), .ZN(n4316) );
  OAI21_X1 U5358 ( .B1(n4317), .B2(n5391), .A(n4316), .ZN(U3456) );
  OR2_X1 U5359 ( .A1(n4318), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4320)
         );
  AND2_X1 U5360 ( .A1(n4320), .A2(n4319), .ZN(n5055) );
  INV_X1 U5361 ( .A(n5055), .ZN(n4331) );
  INV_X1 U5362 ( .A(n4321), .ZN(n4323) );
  INV_X1 U5363 ( .A(n5503), .ZN(n5376) );
  NAND4_X1 U5364 ( .A1(n4323), .A2(n3132), .A3(n5376), .A4(n4322), .ZN(n4356)
         );
  OR2_X1 U5365 ( .A1(n4356), .A2(n4324), .ZN(n4325) );
  NAND2_X1 U5366 ( .A1(n4326), .A2(n4325), .ZN(n4327) );
  OAI21_X1 U5367 ( .B1(n4330), .B2(n4329), .A(n4328), .ZN(n6201) );
  INV_X2 U5368 ( .A(n6041), .ZN(n5819) );
  OAI222_X1 U5369 ( .A1(n4331), .A2(n5817), .B1(n5052), .B2(n6045), .C1(n6201), 
        .C2(n5819), .ZN(U2859) );
  NOR3_X1 U5370 ( .A1(n4349), .A2(n4333), .A3(n4377), .ZN(n4334) );
  AOI21_X1 U5371 ( .B1(n5729), .B2(n4339), .A(n4334), .ZN(n4335) );
  OAI21_X1 U5372 ( .B1(n4575), .B2(n4376), .A(n4335), .ZN(n6411) );
  AOI22_X1 U5373 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4336), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4369), .ZN(n5381) );
  INV_X1 U5374 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5382) );
  NOR2_X1 U5375 ( .A1(n6441), .A2(n5382), .ZN(n4338) );
  AOI222_X1 U5376 ( .A1(n6411), .A2(n5902), .B1(n5381), .B2(n4338), .C1(n4337), 
        .C2(n5387), .ZN(n4340) );
  AOI21_X1 U5377 ( .B1(n4347), .B2(n5387), .A(n5391), .ZN(n4350) );
  OAI22_X1 U5378 ( .A1(n4340), .A2(n5391), .B1(n4350), .B2(n4339), .ZN(U3460)
         );
  OAI21_X1 U5379 ( .B1(n4341), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n3233), 
        .ZN(n6194) );
  INV_X1 U5380 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6552) );
  NOR2_X1 U5381 ( .A1(n6192), .A2(n6552), .ZN(n4342) );
  AOI211_X1 U5382 ( .C1(n6240), .C2(n5055), .A(n4343), .B(n4342), .ZN(n4346)
         );
  OAI21_X1 U5383 ( .B1(n5220), .B2(n4344), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4345) );
  OAI211_X1 U5384 ( .C1(n6194), .C2(n5717), .A(n4346), .B(n4345), .ZN(U3018)
         );
  INV_X1 U5385 ( .A(n5729), .ZN(n4348) );
  NOR2_X1 U5386 ( .A1(n4348), .A2(n4347), .ZN(n6409) );
  INV_X1 U5387 ( .A(n6409), .ZN(n4355) );
  INV_X1 U5388 ( .A(n5902), .ZN(n4354) );
  OAI22_X1 U5389 ( .A1(n3690), .A2(n4376), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4349), .ZN(n6410) );
  NAND2_X1 U5390 ( .A1(n6410), .A2(n5902), .ZN(n4351) );
  OAI211_X1 U5391 ( .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n6441), .A(n4351), 
        .B(n4350), .ZN(n4352) );
  OAI21_X1 U5392 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5906), .A(n4352), 
        .ZN(n4353) );
  OAI21_X1 U5393 ( .B1(n4355), .B2(n4354), .A(n4353), .ZN(U3461) );
  NOR2_X1 U5394 ( .A1(n4356), .A2(n4990), .ZN(n4357) );
  OAI21_X1 U5395 ( .B1(n4358), .B2(n4357), .A(n6436), .ZN(n4359) );
  NAND2_X1 U5396 ( .A1(n4360), .A2(n5503), .ZN(n4361) );
  NAND2_X2 U5397 ( .A1(n5505), .A2(n4361), .ZN(n6047) );
  INV_X1 U5398 ( .A(n4361), .ZN(n4362) );
  INV_X1 U5399 ( .A(DATAI_0_), .ZN(n4465) );
  INV_X1 U5400 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6145) );
  OAI222_X1 U5401 ( .A1(n6201), .A2(n6047), .B1(n5329), .B2(n4465), .C1(n5505), 
        .C2(n6145), .ZN(U2891) );
  OAI21_X1 U5402 ( .B1(n4365), .B2(n4364), .A(n4363), .ZN(n4480) );
  OR2_X1 U5403 ( .A1(n5363), .A2(n4366), .ZN(n4367) );
  NAND2_X1 U5404 ( .A1(n4368), .A2(n4367), .ZN(n5356) );
  AND2_X1 U5405 ( .A1(n6238), .A2(REIP_REG_1__SCAN_IN), .ZN(n4477) );
  NOR2_X1 U5406 ( .A1(n4369), .A2(n4422), .ZN(n4370) );
  AOI211_X1 U5407 ( .C1(n6240), .C2(n5356), .A(n4477), .B(n4370), .ZN(n4373)
         );
  OR3_X1 U5408 ( .A1(n5107), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4371), 
        .ZN(n4372) );
  OAI211_X1 U5409 ( .C1(n4480), .C2(n5717), .A(n4373), .B(n4372), .ZN(U3017)
         );
  INV_X1 U5410 ( .A(n6566), .ZN(n6450) );
  OR2_X1 U5411 ( .A1(n4375), .A2(n4376), .ZN(n4385) );
  XNOR2_X1 U5412 ( .A(n4377), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4382)
         );
  XNOR2_X1 U5413 ( .A(n5389), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4378)
         );
  NAND2_X1 U5414 ( .A1(n5729), .A2(n4378), .ZN(n4379) );
  OAI21_X1 U5415 ( .B1(n4382), .B2(n4380), .A(n4379), .ZN(n4381) );
  AOI21_X1 U5416 ( .B1(n4383), .B2(n4382), .A(n4381), .ZN(n4384) );
  NAND2_X1 U5417 ( .A1(n4385), .A2(n4384), .ZN(n5386) );
  NAND2_X1 U5418 ( .A1(n5386), .A2(n4391), .ZN(n4387) );
  INV_X1 U5419 ( .A(n4391), .ZN(n6412) );
  NAND2_X1 U5420 ( .A1(n6412), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4386) );
  AND2_X1 U5421 ( .A1(n4387), .A2(n4386), .ZN(n6418) );
  MUX2_X1 U5422 ( .A(n4388), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6412), 
        .Z(n6422) );
  NAND2_X1 U5423 ( .A1(n6441), .A2(n6422), .ZN(n4399) );
  INV_X1 U5424 ( .A(n4936), .ZN(n4520) );
  NOR2_X1 U5425 ( .A1(n4389), .A2(n4520), .ZN(n4390) );
  XNOR2_X1 U5426 ( .A(n4390), .B(n5905), .ZN(n6024) );
  NAND3_X1 U5427 ( .A1(n6024), .A2(n5903), .A3(n6441), .ZN(n4394) );
  NAND2_X1 U5428 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5913), .ZN(n4395) );
  OAI21_X1 U5429 ( .B1(n4391), .B2(STATE2_REG_1__SCAN_IN), .A(n4395), .ZN(
        n4392) );
  NAND2_X1 U5430 ( .A1(n4392), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4393) );
  AND2_X1 U5431 ( .A1(n4394), .A2(n4393), .ZN(n4400) );
  INV_X1 U5432 ( .A(n4395), .ZN(n4396) );
  NAND2_X1 U5433 ( .A1(n4397), .A2(n4396), .ZN(n4398) );
  OAI211_X1 U5434 ( .C1(n6418), .C2(n4399), .A(n4400), .B(n4398), .ZN(n6423)
         );
  NAND2_X1 U5435 ( .A1(n4400), .A2(n4333), .ZN(n4401) );
  NAND2_X1 U5436 ( .A1(n6423), .A2(n4401), .ZN(n4404) );
  AOI21_X1 U5437 ( .B1(n4404), .B2(n5913), .A(n6532), .ZN(n4402) );
  OR2_X1 U5438 ( .A1(n4523), .A2(n4402), .ZN(n6542) );
  NAND2_X1 U5439 ( .A1(n4404), .A2(n4403), .ZN(n6433) );
  INV_X1 U5440 ( .A(n6433), .ZN(n4406) );
  NOR2_X1 U5441 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6441), .ZN(n4428) );
  OAI22_X1 U5442 ( .A1(n4942), .A2(n6343), .B1(n4428), .B2(n3690), .ZN(n4405)
         );
  OAI21_X1 U5443 ( .B1(n4406), .B2(n4405), .A(n6542), .ZN(n4407) );
  OAI21_X1 U5444 ( .B1(n6542), .B2(n6408), .A(n4407), .ZN(U3465) );
  NOR2_X1 U5445 ( .A1(n4410), .A2(n4409), .ZN(n4411) );
  NOR2_X1 U5446 ( .A1(n4408), .A2(n4411), .ZN(n6187) );
  INV_X1 U5447 ( .A(n6187), .ZN(n5008) );
  INV_X1 U5448 ( .A(n4413), .ZN(n4439) );
  XNOR2_X1 U5449 ( .A(n4412), .B(n4439), .ZN(n6237) );
  OAI222_X1 U5450 ( .A1(n5819), .A2(n5008), .B1(n3524), .B2(n6045), .C1(n5817), 
        .C2(n6237), .ZN(U2857) );
  INV_X1 U5451 ( .A(DATAI_2_), .ZN(n6707) );
  INV_X1 U5452 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6151) );
  OAI222_X1 U5453 ( .A1(n5008), .A2(n6047), .B1(n5329), .B2(n6707), .C1(n5505), 
        .C2(n6151), .ZN(U2889) );
  NOR2_X1 U5454 ( .A1(n4414), .A2(n4415), .ZN(n4416) );
  OR2_X1 U5455 ( .A1(n3700), .A2(n4416), .ZN(n5366) );
  INV_X1 U5456 ( .A(DATAI_1_), .ZN(n6633) );
  INV_X1 U5457 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6148) );
  OAI222_X1 U5458 ( .A1(n5366), .A2(n6047), .B1(n5329), .B2(n6633), .C1(n5505), 
        .C2(n6148), .ZN(U2890) );
  XNOR2_X1 U5459 ( .A(n4418), .B(n4417), .ZN(n4609) );
  AOI21_X1 U5460 ( .B1(n6235), .B2(n4423), .A(n4502), .ZN(n4426) );
  AOI21_X1 U5461 ( .B1(n6242), .B2(n6248), .A(n6241), .ZN(n4566) );
  NOR2_X1 U5462 ( .A1(n6243), .A2(n4566), .ZN(n6228) );
  AND2_X1 U5463 ( .A1(n4419), .A2(n4420), .ZN(n4421) );
  OR2_X1 U5464 ( .A1(n4421), .A2(n4500), .ZN(n6030) );
  NAND2_X1 U5465 ( .A1(n5592), .A2(REIP_REG_4__SCAN_IN), .ZN(n4605) );
  OAI21_X1 U5466 ( .B1(n3628), .B2(n6030), .A(n4605), .ZN(n4425) );
  OAI22_X1 U5467 ( .A1(n5214), .A2(n6242), .B1(n6241), .B2(n4422), .ZN(n6246)
         );
  AOI21_X1 U5468 ( .B1(n6241), .B2(n6243), .A(n6246), .ZN(n6236) );
  NOR2_X1 U5469 ( .A1(n6236), .A2(n4423), .ZN(n4424) );
  AOI211_X1 U5470 ( .C1(n4426), .C2(n6228), .A(n4425), .B(n4424), .ZN(n4427)
         );
  OAI21_X1 U5471 ( .B1(n5717), .B2(n4609), .A(n4427), .ZN(U3014) );
  INV_X1 U5472 ( .A(n4428), .ZN(n6541) );
  INV_X1 U5473 ( .A(n4735), .ZN(n4518) );
  AND2_X1 U5474 ( .A1(n4735), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6293) );
  AOI211_X1 U5475 ( .C1(n4518), .C2(n6561), .A(n6343), .B(n6293), .ZN(n4430)
         );
  AOI21_X1 U5476 ( .B1(n6541), .B2(n5359), .A(n4430), .ZN(n4432) );
  NAND2_X1 U5477 ( .A1(n6545), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4431) );
  OAI21_X1 U5478 ( .B1(n4432), .B2(n6545), .A(n4431), .ZN(U3464) );
  XNOR2_X1 U5479 ( .A(n6293), .B(n4736), .ZN(n4434) );
  INV_X1 U5480 ( .A(n4375), .ZN(n5006) );
  AOI22_X1 U5481 ( .A1(n4434), .A2(n6536), .B1(n5006), .B2(n6541), .ZN(n4436)
         );
  NAND2_X1 U5482 ( .A1(n6545), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4435) );
  OAI21_X1 U5483 ( .B1(n6545), .B2(n4436), .A(n4435), .ZN(U3463) );
  OAI21_X1 U5484 ( .B1(n4408), .B2(n4437), .A(n4443), .ZN(n5375) );
  INV_X1 U5485 ( .A(DATAI_3_), .ZN(n4459) );
  INV_X1 U5486 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6098) );
  OAI222_X1 U5487 ( .A1(n5375), .A2(n6047), .B1(n5329), .B2(n4459), .C1(n5505), 
        .C2(n6098), .ZN(U2888) );
  INV_X1 U5488 ( .A(EBX_REG_3__SCAN_IN), .ZN(n5096) );
  OAI21_X1 U5489 ( .B1(n4412), .B2(n4439), .A(n4438), .ZN(n4440) );
  NAND2_X1 U5490 ( .A1(n4440), .A2(n4419), .ZN(n6227) );
  OAI222_X1 U5491 ( .A1(n5375), .A2(n5819), .B1(n5096), .B2(n6045), .C1(n6227), 
        .C2(n5817), .ZN(U2856) );
  AND2_X1 U5492 ( .A1(n4443), .A2(n4442), .ZN(n4444) );
  OR2_X1 U5493 ( .A1(n4441), .A2(n4444), .ZN(n4604) );
  INV_X1 U5494 ( .A(n6030), .ZN(n4445) );
  AOI22_X1 U5495 ( .A1(n6040), .A2(n4445), .B1(n5501), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4446) );
  OAI21_X1 U5496 ( .B1(n4604), .B2(n5819), .A(n4446), .ZN(U2855) );
  NOR2_X1 U5497 ( .A1(n6254), .A2(n3690), .ZN(n4771) );
  OR2_X1 U5498 ( .A1(n4375), .A2(n4575), .ZN(n6259) );
  INV_X1 U5499 ( .A(n4512), .ZN(n4484) );
  AOI21_X1 U5500 ( .B1(n4771), .B2(n6290), .A(n4484), .ZN(n4451) );
  INV_X1 U5501 ( .A(n4451), .ZN(n4448) );
  AOI22_X1 U5502 ( .A1(n4448), .A2(n4897), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4447), .ZN(n4508) );
  NOR2_X1 U5503 ( .A1(n6707), .A2(n4893), .ZN(n6360) );
  INV_X1 U5504 ( .A(n6360), .ZN(n6310) );
  OAI21_X1 U5505 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6718), .A(n4523), 
        .ZN(n6342) );
  INV_X1 U5506 ( .A(n6342), .ZN(n6297) );
  INV_X1 U5507 ( .A(n4519), .ZN(n4449) );
  OR2_X1 U5508 ( .A1(n4736), .A2(n4449), .ZN(n4728) );
  NAND2_X1 U5509 ( .A1(n6536), .A2(n6561), .ZN(n5152) );
  OAI21_X1 U5510 ( .B1(n4455), .B2(n6200), .A(n5152), .ZN(n4450) );
  AOI22_X1 U5511 ( .A1(n4451), .A2(n4450), .B1(n4854), .B2(n6343), .ZN(n4452)
         );
  NAND2_X1 U5512 ( .A1(n6297), .A2(n4452), .ZN(n4515) );
  NAND2_X1 U5513 ( .A1(n4515), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4458)
         );
  NOR2_X1 U5514 ( .A1(n4511), .A2(n4454), .ZN(n6358) );
  INV_X1 U5515 ( .A(DATAI_26_), .ZN(n6642) );
  OR2_X1 U5516 ( .A1(n6200), .A2(n6642), .ZN(n4968) );
  NAND2_X1 U5517 ( .A1(n4455), .A2(n4777), .ZN(n4631) );
  INV_X1 U5518 ( .A(DATAI_18_), .ZN(n6046) );
  OR2_X1 U5519 ( .A1(n6200), .A2(n6046), .ZN(n6363) );
  OAI22_X1 U5520 ( .A1(n4968), .A2(n4885), .B1(n4631), .B2(n6363), .ZN(n4456)
         );
  AOI21_X1 U5521 ( .B1(n4484), .B2(n6358), .A(n4456), .ZN(n4457) );
  OAI211_X1 U5522 ( .C1(n4508), .C2(n6310), .A(n4458), .B(n4457), .ZN(U3142)
         );
  NOR2_X1 U5523 ( .A1(n4459), .A2(n4893), .ZN(n6366) );
  INV_X1 U5524 ( .A(n6366), .ZN(n6314) );
  NAND2_X1 U5525 ( .A1(n4515), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4464)
         );
  NOR2_X1 U5526 ( .A1(n4511), .A2(n4460), .ZN(n6364) );
  INV_X1 U5527 ( .A(DATAI_27_), .ZN(n5826) );
  OR2_X1 U5528 ( .A1(n6200), .A2(n5826), .ZN(n4973) );
  INV_X1 U5529 ( .A(DATAI_19_), .ZN(n4461) );
  OR2_X1 U5530 ( .A1(n6200), .A2(n4461), .ZN(n6369) );
  OAI22_X1 U5531 ( .A1(n4973), .A2(n4885), .B1(n4631), .B2(n6369), .ZN(n4462)
         );
  AOI21_X1 U5532 ( .B1(n4484), .B2(n6364), .A(n4462), .ZN(n4463) );
  OAI211_X1 U5533 ( .C1(n4508), .C2(n6314), .A(n4464), .B(n4463), .ZN(U3143)
         );
  NOR2_X1 U5534 ( .A1(n4465), .A2(n4893), .ZN(n6349) );
  INV_X1 U5535 ( .A(n6349), .ZN(n6303) );
  NAND2_X1 U5536 ( .A1(n4515), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4469)
         );
  NOR2_X1 U5537 ( .A1(n4511), .A2(n3180), .ZN(n6336) );
  INV_X1 U5538 ( .A(DATAI_24_), .ZN(n4466) );
  OR2_X1 U5539 ( .A1(n6200), .A2(n4466), .ZN(n6352) );
  INV_X1 U5540 ( .A(DATAI_16_), .ZN(n6057) );
  OR2_X1 U5541 ( .A1(n6200), .A2(n6057), .ZN(n6267) );
  OAI22_X1 U5542 ( .A1(n6352), .A2(n4885), .B1(n4631), .B2(n6267), .ZN(n4467)
         );
  AOI21_X1 U5543 ( .B1(n4484), .B2(n6336), .A(n4467), .ZN(n4468) );
  OAI211_X1 U5544 ( .C1(n4508), .C2(n6303), .A(n4469), .B(n4468), .ZN(U3140)
         );
  INV_X1 U5545 ( .A(DATAI_4_), .ZN(n4474) );
  NOR2_X1 U5546 ( .A1(n4474), .A2(n4893), .ZN(n6372) );
  INV_X1 U5547 ( .A(n6372), .ZN(n6318) );
  NAND2_X1 U5548 ( .A1(n4515), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4473)
         );
  NOR2_X1 U5549 ( .A1(n4511), .A2(n3132), .ZN(n6370) );
  INV_X1 U5550 ( .A(DATAI_28_), .ZN(n4470) );
  OR2_X1 U5551 ( .A1(n6200), .A2(n4470), .ZN(n4978) );
  INV_X1 U5552 ( .A(DATAI_20_), .ZN(n5847) );
  OR2_X1 U5553 ( .A1(n6200), .A2(n5847), .ZN(n6375) );
  OAI22_X1 U5554 ( .A1(n4978), .A2(n4885), .B1(n4631), .B2(n6375), .ZN(n4471)
         );
  AOI21_X1 U5555 ( .B1(n4484), .B2(n6370), .A(n4471), .ZN(n4472) );
  OAI211_X1 U5556 ( .C1(n4508), .C2(n6318), .A(n4473), .B(n4472), .ZN(U3144)
         );
  INV_X1 U5557 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6154) );
  OAI222_X1 U5558 ( .A1(n4604), .A2(n6047), .B1(n5329), .B2(n4474), .C1(n5505), 
        .C2(n6154), .ZN(U2887) );
  INV_X1 U5559 ( .A(n5366), .ZN(n4475) );
  NAND2_X1 U5560 ( .A1(n4475), .A2(n6186), .ZN(n4479) );
  NOR2_X1 U5561 ( .A1(n6191), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4476)
         );
  AOI211_X1 U5562 ( .C1(n6197), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4477), 
        .B(n4476), .ZN(n4478) );
  OAI211_X1 U5563 ( .C1(n6193), .C2(n4480), .A(n4479), .B(n4478), .ZN(U2985)
         );
  INV_X1 U5564 ( .A(DATAI_5_), .ZN(n4556) );
  NOR2_X1 U5565 ( .A1(n4556), .A2(n4893), .ZN(n6378) );
  INV_X1 U5566 ( .A(n6378), .ZN(n6322) );
  NAND2_X1 U5567 ( .A1(n4515), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4486)
         );
  NOR2_X1 U5568 ( .A1(n4511), .A2(n3190), .ZN(n6376) );
  INV_X1 U5569 ( .A(DATAI_29_), .ZN(n4481) );
  OR2_X1 U5570 ( .A1(n6200), .A2(n4481), .ZN(n6381) );
  INV_X1 U5571 ( .A(DATAI_21_), .ZN(n4482) );
  OR2_X1 U5572 ( .A1(n6200), .A2(n4482), .ZN(n6278) );
  OAI22_X1 U5573 ( .A1(n6381), .A2(n4885), .B1(n4631), .B2(n6278), .ZN(n4483)
         );
  AOI21_X1 U5574 ( .B1(n4484), .B2(n6376), .A(n4483), .ZN(n4485) );
  OAI211_X1 U5575 ( .C1(n4508), .C2(n6322), .A(n4486), .B(n4485), .ZN(U3145)
         );
  NAND2_X1 U5576 ( .A1(DATAI_7_), .A2(n4523), .ZN(n6334) );
  INV_X1 U5577 ( .A(DATAI_23_), .ZN(n4487) );
  OR2_X1 U5578 ( .A1(n6200), .A2(n4487), .ZN(n6288) );
  OAI22_X1 U5579 ( .A1(n6334), .A2(n4508), .B1(n4631), .B2(n6288), .ZN(n4490)
         );
  INV_X1 U5580 ( .A(DATAI_31_), .ZN(n4488) );
  OR2_X1 U5581 ( .A1(n6200), .A2(n4488), .ZN(n6400) );
  NOR2_X1 U5582 ( .A1(n4511), .A2(n5376), .ZN(n6391) );
  INV_X1 U5583 ( .A(n6391), .ZN(n4915) );
  OAI22_X1 U5584 ( .A1(n4885), .A2(n6400), .B1(n4915), .B2(n4512), .ZN(n4489)
         );
  AOI211_X1 U5585 ( .C1(n4515), .C2(INSTQUEUE_REG_15__7__SCAN_IN), .A(n4490), 
        .B(n4489), .ZN(n4491) );
  INV_X1 U5586 ( .A(n4491), .ZN(U3147) );
  NAND2_X1 U5587 ( .A1(DATAI_6_), .A2(n4523), .ZN(n6326) );
  INV_X1 U5588 ( .A(DATAI_22_), .ZN(n5839) );
  OR2_X1 U5589 ( .A1(n6200), .A2(n5839), .ZN(n6389) );
  OAI22_X1 U5590 ( .A1(n6326), .A2(n4508), .B1(n4631), .B2(n6389), .ZN(n4494)
         );
  INV_X1 U5591 ( .A(DATAI_30_), .ZN(n4492) );
  OR2_X1 U5592 ( .A1(n6200), .A2(n4492), .ZN(n4963) );
  NOR2_X1 U5593 ( .A1(n4511), .A2(n3497), .ZN(n6382) );
  INV_X1 U5594 ( .A(n6382), .ZN(n4904) );
  OAI22_X1 U5595 ( .A1(n4885), .A2(n4963), .B1(n4904), .B2(n4512), .ZN(n4493)
         );
  AOI211_X1 U5596 ( .C1(n4515), .C2(INSTQUEUE_REG_15__6__SCAN_IN), .A(n4494), 
        .B(n4493), .ZN(n4495) );
  INV_X1 U5597 ( .A(n4495), .ZN(U3146) );
  XNOR2_X1 U5598 ( .A(n4496), .B(n4497), .ZN(n4768) );
  OR2_X1 U5599 ( .A1(n4500), .A2(n4499), .ZN(n4501) );
  AND2_X1 U5600 ( .A1(n4498), .A2(n4501), .ZN(n6006) );
  AND2_X1 U5601 ( .A1(n6238), .A2(REIP_REG_5__SCAN_IN), .ZN(n4764) );
  NAND2_X1 U5602 ( .A1(n4502), .A2(n6228), .ZN(n5027) );
  NAND2_X1 U5603 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4503), .ZN(n4565)
         );
  AOI21_X1 U5604 ( .B1(n5883), .B2(n4565), .A(n6246), .ZN(n4567) );
  AOI21_X1 U5605 ( .B1(n4504), .B2(n5027), .A(n4567), .ZN(n4505) );
  AOI211_X1 U5606 ( .C1(n6240), .C2(n6006), .A(n4764), .B(n4505), .ZN(n4506)
         );
  OAI21_X1 U5607 ( .B1(n5717), .B2(n4768), .A(n4506), .ZN(U3013) );
  NAND2_X1 U5608 ( .A1(DATAI_1_), .A2(n4523), .ZN(n6577) );
  INV_X1 U5609 ( .A(DATAI_17_), .ZN(n4507) );
  OR2_X1 U5610 ( .A1(n6200), .A2(n4507), .ZN(n6576) );
  OAI22_X1 U5611 ( .A1(n4508), .A2(n6577), .B1(n4631), .B2(n6576), .ZN(n4514)
         );
  INV_X1 U5612 ( .A(DATAI_25_), .ZN(n4509) );
  OR2_X1 U5613 ( .A1(n6200), .A2(n4509), .ZN(n6572) );
  NOR2_X1 U5614 ( .A1(n4511), .A2(n4510), .ZN(n6353) );
  INV_X1 U5615 ( .A(n6353), .ZN(n6574) );
  OAI22_X1 U5616 ( .A1(n4885), .A2(n6572), .B1(n6574), .B2(n4512), .ZN(n4513)
         );
  AOI211_X1 U5617 ( .C1(n4515), .C2(INSTQUEUE_REG_15__1__SCAN_IN), .A(n4514), 
        .B(n4513), .ZN(n4516) );
  INV_X1 U5618 ( .A(n4516), .ZN(U3141) );
  NAND2_X1 U5619 ( .A1(n4736), .A2(n4777), .ZN(n4517) );
  INV_X1 U5620 ( .A(n5152), .ZN(n6538) );
  NOR2_X1 U5621 ( .A1(n4375), .A2(n5359), .ZN(n4937) );
  OR2_X1 U5622 ( .A1(n4736), .A2(n4519), .ZN(n6294) );
  OAI21_X1 U5623 ( .B1(n4943), .B2(n6561), .A(n4897), .ZN(n4949) );
  AOI21_X1 U5624 ( .B1(n4520), .B2(n4937), .A(n4949), .ZN(n4521) );
  OAI21_X1 U5625 ( .B1(n6538), .B2(n6575), .A(n4521), .ZN(n4525) );
  NAND3_X1 U5626 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6544), .A3(n4769), .ZN(n4946) );
  OR2_X1 U5627 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4946), .ZN(n4558)
         );
  AND2_X1 U5628 ( .A1(n4526), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4855) );
  INV_X1 U5629 ( .A(n4691), .ZN(n4522) );
  NOR2_X1 U5630 ( .A1(n4522), .A2(n6255), .ZN(n4582) );
  OAI21_X1 U5631 ( .B1(n4582), .B2(n6560), .A(n4523), .ZN(n4578) );
  AOI211_X1 U5632 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4558), .A(n4855), .B(
        n4578), .ZN(n4524) );
  NAND2_X1 U5633 ( .A1(n4525), .A2(n4524), .ZN(n4557) );
  NAND2_X1 U5634 ( .A1(n4557), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4532) );
  INV_X1 U5635 ( .A(n4582), .ZN(n4528) );
  NOR2_X1 U5636 ( .A1(n4526), .A2(n6560), .ZN(n6256) );
  INV_X1 U5637 ( .A(n6256), .ZN(n4851) );
  NAND3_X1 U5638 ( .A1(n6254), .A2(n6536), .A3(n4937), .ZN(n4527) );
  OAI21_X1 U5639 ( .B1(n4528), .B2(n4851), .A(n4527), .ZN(n4560) );
  INV_X1 U5640 ( .A(n4943), .ZN(n4529) );
  NAND2_X1 U5641 ( .A1(n4529), .A2(n4942), .ZN(n4984) );
  INV_X1 U5642 ( .A(n6364), .ZN(n4900) );
  OAI22_X1 U5643 ( .A1(n4984), .A2(n6369), .B1(n4900), .B2(n4558), .ZN(n4530)
         );
  AOI21_X1 U5644 ( .B1(n6366), .B2(n4560), .A(n4530), .ZN(n4531) );
  OAI211_X1 U5645 ( .C1(n6575), .C2(n4973), .A(n4532), .B(n4531), .ZN(U3055)
         );
  NAND2_X1 U5646 ( .A1(n4557), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4535) );
  INV_X1 U5647 ( .A(n6288), .ZN(n6392) );
  INV_X1 U5648 ( .A(n4984), .ZN(n4550) );
  INV_X1 U5649 ( .A(n4560), .ZN(n4548) );
  OAI22_X1 U5650 ( .A1(n6334), .A2(n4548), .B1(n4915), .B2(n4558), .ZN(n4533)
         );
  AOI21_X1 U5651 ( .B1(n6392), .B2(n4550), .A(n4533), .ZN(n4534) );
  OAI211_X1 U5652 ( .C1(n6575), .C2(n6400), .A(n4535), .B(n4534), .ZN(U3059)
         );
  NAND2_X1 U5653 ( .A1(n4557), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4538) );
  INV_X1 U5654 ( .A(n6336), .ZN(n4929) );
  OAI22_X1 U5655 ( .A1(n6267), .A2(n4984), .B1(n4929), .B2(n4558), .ZN(n4536)
         );
  AOI21_X1 U5656 ( .B1(n6349), .B2(n4560), .A(n4536), .ZN(n4537) );
  OAI211_X1 U5657 ( .C1(n6575), .C2(n6352), .A(n4538), .B(n4537), .ZN(U3052)
         );
  NAND2_X1 U5658 ( .A1(n4557), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4541) );
  INV_X1 U5659 ( .A(n6370), .ZN(n4911) );
  OAI22_X1 U5660 ( .A1(n4984), .A2(n6375), .B1(n4911), .B2(n4558), .ZN(n4539)
         );
  AOI21_X1 U5661 ( .B1(n6372), .B2(n4560), .A(n4539), .ZN(n4540) );
  OAI211_X1 U5662 ( .C1(n6575), .C2(n4978), .A(n4541), .B(n4540), .ZN(U3056)
         );
  NAND2_X1 U5663 ( .A1(n4557), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4544) );
  INV_X1 U5664 ( .A(n6358), .ZN(n4919) );
  OAI22_X1 U5665 ( .A1(n4984), .A2(n6363), .B1(n4919), .B2(n4558), .ZN(n4542)
         );
  AOI21_X1 U5666 ( .B1(n6360), .B2(n4560), .A(n4542), .ZN(n4543) );
  OAI211_X1 U5667 ( .C1(n6575), .C2(n4968), .A(n4544), .B(n4543), .ZN(U3054)
         );
  NAND2_X1 U5668 ( .A1(n4557), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4547) );
  INV_X1 U5669 ( .A(n6576), .ZN(n6354) );
  OAI22_X1 U5670 ( .A1(n6574), .A2(n4558), .B1(n4548), .B2(n6577), .ZN(n4545)
         );
  AOI21_X1 U5671 ( .B1(n6354), .B2(n4550), .A(n4545), .ZN(n4546) );
  OAI211_X1 U5672 ( .C1(n6575), .C2(n6572), .A(n4547), .B(n4546), .ZN(U3053)
         );
  NAND2_X1 U5673 ( .A1(n4557), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4552) );
  INV_X1 U5674 ( .A(n6389), .ZN(n6323) );
  OAI22_X1 U5675 ( .A1(n6326), .A2(n4548), .B1(n4904), .B2(n4558), .ZN(n4549)
         );
  AOI21_X1 U5676 ( .B1(n6323), .B2(n4550), .A(n4549), .ZN(n4551) );
  OAI211_X1 U5677 ( .C1(n6575), .C2(n4963), .A(n4552), .B(n4551), .ZN(U3058)
         );
  OAI21_X1 U5678 ( .B1(n4441), .B2(n4554), .A(n4553), .ZN(n4763) );
  INV_X1 U5679 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6691) );
  INV_X1 U5680 ( .A(n6006), .ZN(n4555) );
  OAI222_X1 U5681 ( .A1(n4763), .A2(n5819), .B1(n6045), .B2(n6691), .C1(n4555), 
        .C2(n5817), .ZN(U2854) );
  OAI222_X1 U5682 ( .A1(n4763), .A2(n6047), .B1(n5329), .B2(n4556), .C1(n5505), 
        .C2(n3734), .ZN(U2886) );
  NAND2_X1 U5683 ( .A1(n4557), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4562) );
  INV_X1 U5684 ( .A(n6376), .ZN(n4923) );
  OAI22_X1 U5685 ( .A1(n4984), .A2(n6278), .B1(n4923), .B2(n4558), .ZN(n4559)
         );
  AOI21_X1 U5686 ( .B1(n6378), .B2(n4560), .A(n4559), .ZN(n4561) );
  OAI211_X1 U5687 ( .C1(n6575), .C2(n6381), .A(n4562), .B(n4561), .ZN(U3057)
         );
  XNOR2_X1 U5688 ( .A(n4563), .B(n4564), .ZN(n4806) );
  NOR2_X1 U5689 ( .A1(n4566), .A2(n4565), .ZN(n4569) );
  INV_X1 U5690 ( .A(n4567), .ZN(n4568) );
  MUX2_X1 U5691 ( .A(n4569), .B(n4568), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4570) );
  INV_X1 U5692 ( .A(n4570), .ZN(n4573) );
  INV_X1 U5693 ( .A(n5013), .ZN(n4571) );
  XNOR2_X1 U5694 ( .A(n4498), .B(n4571), .ZN(n6039) );
  AOI22_X1 U5695 ( .A1(n6240), .A2(n6039), .B1(n6238), .B2(REIP_REG_6__SCAN_IN), .ZN(n4572) );
  OAI211_X1 U5696 ( .C1(n4806), .C2(n5717), .A(n4573), .B(n4572), .ZN(U3012)
         );
  NOR2_X2 U5697 ( .A1(n4610), .A2(n4777), .ZN(n4686) );
  NOR3_X1 U5698 ( .A1(n4599), .A2(n4686), .A3(n6343), .ZN(n4577) );
  NAND2_X1 U5699 ( .A1(n4375), .A2(n4575), .ZN(n4641) );
  NOR2_X1 U5700 ( .A1(n6540), .A2(n4641), .ZN(n4611) );
  INV_X1 U5701 ( .A(n4611), .ZN(n4576) );
  OAI21_X1 U5702 ( .B1(n4577), .B2(n6538), .A(n4576), .ZN(n4581) );
  NAND3_X1 U5703 ( .A1(n6544), .A2(n4642), .A3(n4769), .ZN(n4615) );
  NOR2_X1 U5704 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4615), .ZN(n4634)
         );
  INV_X1 U5705 ( .A(n4634), .ZN(n4579) );
  AOI211_X1 U5706 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4579), .A(n6256), .B(
        n4578), .ZN(n4580) );
  INV_X1 U5707 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4586) );
  INV_X1 U5708 ( .A(n6369), .ZN(n6311) );
  AOI22_X1 U5709 ( .A1(n4611), .A2(n4897), .B1(n4855), .B2(n4582), .ZN(n4632)
         );
  INV_X1 U5710 ( .A(n4973), .ZN(n6365) );
  AOI22_X1 U5711 ( .A1(n4599), .A2(n6365), .B1(n6364), .B2(n4634), .ZN(n4583)
         );
  OAI21_X1 U5712 ( .B1(n6314), .B2(n4632), .A(n4583), .ZN(n4584) );
  AOI21_X1 U5713 ( .B1(n6311), .B2(n4686), .A(n4584), .ZN(n4585) );
  OAI21_X1 U5714 ( .B1(n4638), .B2(n4586), .A(n4585), .ZN(U3023) );
  INV_X1 U5715 ( .A(n6267), .ZN(n6337) );
  INV_X1 U5716 ( .A(n6352), .ZN(n6292) );
  AOI22_X1 U5717 ( .A1(n4599), .A2(n6292), .B1(n6336), .B2(n4634), .ZN(n4587)
         );
  OAI21_X1 U5718 ( .B1(n6303), .B2(n4632), .A(n4587), .ZN(n4588) );
  AOI21_X1 U5719 ( .B1(n6337), .B2(n4686), .A(n4588), .ZN(n4589) );
  OAI21_X1 U5720 ( .B1(n4638), .B2(n4590), .A(n4589), .ZN(U3020) );
  INV_X1 U5721 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4594) );
  INV_X1 U5722 ( .A(n6363), .ZN(n6307) );
  INV_X1 U5723 ( .A(n4968), .ZN(n6359) );
  AOI22_X1 U5724 ( .A1(n4599), .A2(n6359), .B1(n6358), .B2(n4634), .ZN(n4591)
         );
  OAI21_X1 U5725 ( .B1(n6310), .B2(n4632), .A(n4591), .ZN(n4592) );
  AOI21_X1 U5726 ( .B1(n6307), .B2(n4686), .A(n4592), .ZN(n4593) );
  OAI21_X1 U5727 ( .B1(n4638), .B2(n4594), .A(n4593), .ZN(U3022) );
  INV_X1 U5728 ( .A(n6278), .ZN(n6377) );
  INV_X1 U5729 ( .A(n6381), .ZN(n6319) );
  AOI22_X1 U5730 ( .A1(n4599), .A2(n6319), .B1(n6376), .B2(n4634), .ZN(n4595)
         );
  OAI21_X1 U5731 ( .B1(n6322), .B2(n4632), .A(n4595), .ZN(n4596) );
  AOI21_X1 U5732 ( .B1(n6377), .B2(n4686), .A(n4596), .ZN(n4597) );
  OAI21_X1 U5733 ( .B1(n4638), .B2(n4598), .A(n4597), .ZN(U3025) );
  INV_X1 U5734 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4603) );
  INV_X1 U5735 ( .A(n6375), .ZN(n6315) );
  INV_X1 U5736 ( .A(n4978), .ZN(n6371) );
  AOI22_X1 U5737 ( .A1(n4599), .A2(n6371), .B1(n6370), .B2(n4634), .ZN(n4600)
         );
  OAI21_X1 U5738 ( .B1(n6318), .B2(n4632), .A(n4600), .ZN(n4601) );
  AOI21_X1 U5739 ( .B1(n6315), .B2(n4686), .A(n4601), .ZN(n4602) );
  OAI21_X1 U5740 ( .B1(n4638), .B2(n4603), .A(n4602), .ZN(U3024) );
  INV_X1 U5741 ( .A(n4604), .ZN(n6034) );
  NOR2_X1 U5742 ( .A1(n6191), .A2(n6038), .ZN(n4607) );
  OAI21_X1 U5743 ( .B1(n5873), .B2(n6019), .A(n4605), .ZN(n4606) );
  AOI211_X1 U5744 ( .C1(n6034), .C2(n6186), .A(n4607), .B(n4606), .ZN(n4608)
         );
  OAI21_X1 U5745 ( .B1(n6193), .B2(n4609), .A(n4608), .ZN(U2982) );
  INV_X1 U5746 ( .A(n3690), .ZN(n6340) );
  NOR2_X1 U5747 ( .A1(n6408), .A2(n4615), .ZN(n4685) );
  AOI21_X1 U5748 ( .B1(n4611), .B2(n6340), .A(n4685), .ZN(n4616) );
  AOI21_X1 U5749 ( .B1(n4612), .B2(STATEBS16_REG_SCAN_IN), .A(n6343), .ZN(
        n4614) );
  AOI22_X1 U5750 ( .A1(n4616), .A2(n4614), .B1(n6343), .B2(n4615), .ZN(n4613)
         );
  NAND2_X1 U5751 ( .A1(n6297), .A2(n4613), .ZN(n4684) );
  INV_X1 U5752 ( .A(n6326), .ZN(n6385) );
  INV_X1 U5753 ( .A(n4614), .ZN(n4617) );
  OAI22_X1 U5754 ( .A1(n4617), .A2(n4616), .B1(n6560), .B2(n4615), .ZN(n4683)
         );
  AOI22_X1 U5755 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4684), .B1(n6385), 
        .B2(n4683), .ZN(n4619) );
  INV_X1 U5756 ( .A(n4963), .ZN(n6383) );
  AOI22_X1 U5757 ( .A1(n4686), .A2(n6383), .B1(n6382), .B2(n4685), .ZN(n4618)
         );
  OAI211_X1 U5758 ( .C1(n6389), .C2(n4935), .A(n4619), .B(n4618), .ZN(U3034)
         );
  INV_X1 U5759 ( .A(n6577), .ZN(n6355) );
  AOI22_X1 U5760 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4684), .B1(n6355), 
        .B2(n4683), .ZN(n4621) );
  INV_X1 U5761 ( .A(n6572), .ZN(n6304) );
  AOI22_X1 U5762 ( .A1(n4686), .A2(n6304), .B1(n6353), .B2(n4685), .ZN(n4620)
         );
  OAI211_X1 U5763 ( .C1(n6576), .C2(n4935), .A(n4621), .B(n4620), .ZN(U3029)
         );
  INV_X1 U5764 ( .A(n6334), .ZN(n6395) );
  AOI22_X1 U5765 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4684), .B1(n6395), 
        .B2(n4683), .ZN(n4623) );
  INV_X1 U5766 ( .A(n6400), .ZN(n6330) );
  AOI22_X1 U5767 ( .A1(n4686), .A2(n6330), .B1(n6391), .B2(n4685), .ZN(n4622)
         );
  OAI211_X1 U5768 ( .C1(n6288), .C2(n4935), .A(n4623), .B(n4622), .ZN(U3035)
         );
  OAI22_X1 U5769 ( .A1(n6334), .A2(n4632), .B1(n4631), .B2(n6400), .ZN(n4624)
         );
  AOI21_X1 U5770 ( .B1(n6391), .B2(n4634), .A(n4624), .ZN(n4626) );
  NAND2_X1 U5771 ( .A1(n4686), .A2(n6392), .ZN(n4625) );
  OAI211_X1 U5772 ( .C1(n4638), .C2(n4627), .A(n4626), .B(n4625), .ZN(U3027)
         );
  OAI22_X1 U5773 ( .A1(n4631), .A2(n6572), .B1(n4632), .B2(n6577), .ZN(n4628)
         );
  AOI21_X1 U5774 ( .B1(n6353), .B2(n4634), .A(n4628), .ZN(n4630) );
  NAND2_X1 U5775 ( .A1(n4686), .A2(n6354), .ZN(n4629) );
  OAI211_X1 U5776 ( .C1(n4638), .C2(n6694), .A(n4630), .B(n4629), .ZN(U3021)
         );
  INV_X1 U5777 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4637) );
  OAI22_X1 U5778 ( .A1(n6326), .A2(n4632), .B1(n4631), .B2(n4963), .ZN(n4633)
         );
  AOI21_X1 U5779 ( .B1(n6382), .B2(n4634), .A(n4633), .ZN(n4636) );
  NAND2_X1 U5780 ( .A1(n4686), .A2(n6323), .ZN(n4635) );
  OAI211_X1 U5781 ( .C1(n4638), .C2(n4637), .A(n4636), .B(n4635), .ZN(U3026)
         );
  AOI22_X1 U5782 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4684), .B1(n6349), 
        .B2(n4683), .ZN(n4640) );
  AOI22_X1 U5783 ( .A1(n4686), .A2(n6292), .B1(n6336), .B2(n4685), .ZN(n4639)
         );
  OAI211_X1 U5784 ( .C1(n6267), .C2(n4935), .A(n4640), .B(n4639), .ZN(U3028)
         );
  INV_X1 U5785 ( .A(n4641), .ZN(n4694) );
  NAND3_X1 U5786 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4642), .A3(n4769), .ZN(n4690) );
  NOR2_X1 U5787 ( .A1(n6408), .A2(n4690), .ZN(n4649) );
  AOI21_X1 U5788 ( .B1(n4771), .B2(n4694), .A(n4649), .ZN(n4647) );
  OR3_X1 U5789 ( .A1(n6339), .A2(n4735), .A3(n6561), .ZN(n4643) );
  AOI22_X1 U5790 ( .A1(n4647), .A2(n4645), .B1(n6343), .B2(n4690), .ZN(n4644)
         );
  NAND2_X1 U5791 ( .A1(n6297), .A2(n4644), .ZN(n4672) );
  INV_X1 U5792 ( .A(n4645), .ZN(n4646) );
  OAI22_X1 U5793 ( .A1(n4647), .A2(n4646), .B1(n6560), .B2(n4690), .ZN(n4671)
         );
  AOI22_X1 U5794 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4672), .B1(n6385), 
        .B2(n4671), .ZN(n4652) );
  INV_X1 U5795 ( .A(n4649), .ZN(n4673) );
  OAI22_X1 U5796 ( .A1(n5159), .A2(n6389), .B1(n4673), .B2(n4904), .ZN(n4650)
         );
  INV_X1 U5797 ( .A(n4650), .ZN(n4651) );
  OAI211_X1 U5798 ( .C1(n4727), .C2(n4963), .A(n4652), .B(n4651), .ZN(U3098)
         );
  AOI22_X1 U5799 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4672), .B1(n6360), 
        .B2(n4671), .ZN(n4655) );
  OAI22_X1 U5800 ( .A1(n5159), .A2(n6363), .B1(n4673), .B2(n4919), .ZN(n4653)
         );
  INV_X1 U5801 ( .A(n4653), .ZN(n4654) );
  OAI211_X1 U5802 ( .C1(n4727), .C2(n4968), .A(n4655), .B(n4654), .ZN(U3094)
         );
  AOI22_X1 U5803 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4672), .B1(n6366), 
        .B2(n4671), .ZN(n4658) );
  OAI22_X1 U5804 ( .A1(n5159), .A2(n6369), .B1(n4673), .B2(n4900), .ZN(n4656)
         );
  INV_X1 U5805 ( .A(n4656), .ZN(n4657) );
  OAI211_X1 U5806 ( .C1(n4727), .C2(n4973), .A(n4658), .B(n4657), .ZN(U3095)
         );
  AOI22_X1 U5807 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4672), .B1(n6355), 
        .B2(n4671), .ZN(n4661) );
  OAI22_X1 U5808 ( .A1(n5159), .A2(n6576), .B1(n4673), .B2(n6574), .ZN(n4659)
         );
  INV_X1 U5809 ( .A(n4659), .ZN(n4660) );
  OAI211_X1 U5810 ( .C1(n4727), .C2(n6572), .A(n4661), .B(n4660), .ZN(U3093)
         );
  AOI22_X1 U5811 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4672), .B1(n6372), 
        .B2(n4671), .ZN(n4664) );
  OAI22_X1 U5812 ( .A1(n5159), .A2(n6375), .B1(n4673), .B2(n4911), .ZN(n4662)
         );
  INV_X1 U5813 ( .A(n4662), .ZN(n4663) );
  OAI211_X1 U5814 ( .C1(n4727), .C2(n4978), .A(n4664), .B(n4663), .ZN(U3096)
         );
  AOI22_X1 U5815 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4672), .B1(n6395), 
        .B2(n4671), .ZN(n4667) );
  OAI22_X1 U5816 ( .A1(n5159), .A2(n6288), .B1(n4673), .B2(n4915), .ZN(n4665)
         );
  INV_X1 U5817 ( .A(n4665), .ZN(n4666) );
  OAI211_X1 U5818 ( .C1(n4727), .C2(n6400), .A(n4667), .B(n4666), .ZN(U3099)
         );
  AOI22_X1 U5819 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4672), .B1(n6349), 
        .B2(n4671), .ZN(n4670) );
  OAI22_X1 U5820 ( .A1(n5159), .A2(n6267), .B1(n4929), .B2(n4673), .ZN(n4668)
         );
  INV_X1 U5821 ( .A(n4668), .ZN(n4669) );
  OAI211_X1 U5822 ( .C1(n4727), .C2(n6352), .A(n4670), .B(n4669), .ZN(U3092)
         );
  AOI22_X1 U5823 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4672), .B1(n6378), 
        .B2(n4671), .ZN(n4676) );
  OAI22_X1 U5824 ( .A1(n5159), .A2(n6278), .B1(n4673), .B2(n4923), .ZN(n4674)
         );
  INV_X1 U5825 ( .A(n4674), .ZN(n4675) );
  OAI211_X1 U5826 ( .C1(n4727), .C2(n6381), .A(n4676), .B(n4675), .ZN(U3097)
         );
  AOI22_X1 U5827 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4684), .B1(n6360), 
        .B2(n4683), .ZN(n4678) );
  AOI22_X1 U5828 ( .A1(n4686), .A2(n6359), .B1(n6358), .B2(n4685), .ZN(n4677)
         );
  OAI211_X1 U5829 ( .C1(n6363), .C2(n4935), .A(n4678), .B(n4677), .ZN(U3030)
         );
  AOI22_X1 U5830 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4684), .B1(n6366), 
        .B2(n4683), .ZN(n4680) );
  AOI22_X1 U5831 ( .A1(n4686), .A2(n6365), .B1(n6364), .B2(n4685), .ZN(n4679)
         );
  OAI211_X1 U5832 ( .C1(n6369), .C2(n4935), .A(n4680), .B(n4679), .ZN(U3031)
         );
  AOI22_X1 U5833 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4684), .B1(n6372), 
        .B2(n4683), .ZN(n4682) );
  AOI22_X1 U5834 ( .A1(n4686), .A2(n6371), .B1(n6370), .B2(n4685), .ZN(n4681)
         );
  OAI211_X1 U5835 ( .C1(n6375), .C2(n4935), .A(n4682), .B(n4681), .ZN(U3032)
         );
  AOI22_X1 U5836 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4684), .B1(n6378), 
        .B2(n4683), .ZN(n4688) );
  AOI22_X1 U5837 ( .A1(n4686), .A2(n6319), .B1(n6376), .B2(n4685), .ZN(n4687)
         );
  OAI211_X1 U5838 ( .C1(n6278), .C2(n4935), .A(n4688), .B(n4687), .ZN(U3033)
         );
  NAND2_X1 U5839 ( .A1(n4735), .A2(n4777), .ZN(n4807) );
  NAND3_X1 U5840 ( .A1(n4727), .A2(n6536), .A3(n6300), .ZN(n4689) );
  AOI22_X1 U5841 ( .A1(n4689), .A2(n5152), .B1(n4694), .B2(n6540), .ZN(n4693)
         );
  NOR2_X1 U5842 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4690), .ZN(n4718)
         );
  OR2_X1 U5843 ( .A1(n6255), .A2(n4691), .ZN(n4695) );
  AOI21_X1 U5844 ( .B1(n4695), .B2(STATE2_REG_2__SCAN_IN), .A(n4893), .ZN(
        n4810) );
  OAI211_X1 U5845 ( .C1(n6718), .C2(n4718), .A(n4851), .B(n4810), .ZN(n4692)
         );
  NAND2_X1 U5846 ( .A1(n4721), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4700) );
  AND2_X1 U5847 ( .A1(n6540), .A2(n4897), .ZN(n4853) );
  NAND2_X1 U5848 ( .A1(n4853), .A2(n4694), .ZN(n4697) );
  INV_X1 U5849 ( .A(n4695), .ZN(n4813) );
  NAND2_X1 U5850 ( .A1(n4813), .A2(n4855), .ZN(n4696) );
  NAND2_X1 U5851 ( .A1(n4697), .A2(n4696), .ZN(n4724) );
  INV_X1 U5852 ( .A(n4718), .ZN(n4722) );
  OAI22_X1 U5853 ( .A1(n4900), .A2(n4722), .B1(n4973), .B2(n6300), .ZN(n4698)
         );
  AOI21_X1 U5854 ( .B1(n6366), .B2(n4724), .A(n4698), .ZN(n4699) );
  OAI211_X1 U5855 ( .C1(n6369), .C2(n4727), .A(n4700), .B(n4699), .ZN(U3087)
         );
  NAND2_X1 U5856 ( .A1(n4721), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4703) );
  OAI22_X1 U5857 ( .A1(n4929), .A2(n4722), .B1(n6352), .B2(n6300), .ZN(n4701)
         );
  AOI21_X1 U5858 ( .B1(n6349), .B2(n4724), .A(n4701), .ZN(n4702) );
  OAI211_X1 U5859 ( .C1(n6267), .C2(n4727), .A(n4703), .B(n4702), .ZN(U3084)
         );
  NAND2_X1 U5860 ( .A1(n4721), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4706) );
  OAI22_X1 U5861 ( .A1(n4923), .A2(n4722), .B1(n6381), .B2(n6300), .ZN(n4704)
         );
  AOI21_X1 U5862 ( .B1(n6378), .B2(n4724), .A(n4704), .ZN(n4705) );
  OAI211_X1 U5863 ( .C1(n6278), .C2(n4727), .A(n4706), .B(n4705), .ZN(U3089)
         );
  NAND2_X1 U5864 ( .A1(n4721), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4709) );
  OAI22_X1 U5865 ( .A1(n4911), .A2(n4722), .B1(n4978), .B2(n6300), .ZN(n4707)
         );
  AOI21_X1 U5866 ( .B1(n6372), .B2(n4724), .A(n4707), .ZN(n4708) );
  OAI211_X1 U5867 ( .C1(n6375), .C2(n4727), .A(n4709), .B(n4708), .ZN(U3088)
         );
  NAND2_X1 U5868 ( .A1(n4721), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4712) );
  INV_X1 U5869 ( .A(n4724), .ZN(n4716) );
  OAI22_X1 U5870 ( .A1(n6300), .A2(n6572), .B1(n4716), .B2(n6577), .ZN(n4710)
         );
  AOI21_X1 U5871 ( .B1(n6353), .B2(n4718), .A(n4710), .ZN(n4711) );
  OAI211_X1 U5872 ( .C1(n6576), .C2(n4727), .A(n4712), .B(n4711), .ZN(U3085)
         );
  NAND2_X1 U5873 ( .A1(n4721), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4715) );
  OAI22_X1 U5874 ( .A1(n6334), .A2(n4716), .B1(n6400), .B2(n6300), .ZN(n4713)
         );
  AOI21_X1 U5875 ( .B1(n6391), .B2(n4718), .A(n4713), .ZN(n4714) );
  OAI211_X1 U5876 ( .C1(n6288), .C2(n4727), .A(n4715), .B(n4714), .ZN(U3091)
         );
  NAND2_X1 U5877 ( .A1(n4721), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4720) );
  OAI22_X1 U5878 ( .A1(n6326), .A2(n4716), .B1(n4963), .B2(n6300), .ZN(n4717)
         );
  AOI21_X1 U5879 ( .B1(n6382), .B2(n4718), .A(n4717), .ZN(n4719) );
  OAI211_X1 U5880 ( .C1(n6389), .C2(n4727), .A(n4720), .B(n4719), .ZN(U3090)
         );
  NAND2_X1 U5881 ( .A1(n4721), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4726) );
  OAI22_X1 U5882 ( .A1(n4919), .A2(n4722), .B1(n4968), .B2(n6300), .ZN(n4723)
         );
  AOI21_X1 U5883 ( .B1(n6360), .B2(n4724), .A(n4723), .ZN(n4725) );
  OAI211_X1 U5884 ( .C1(n6363), .C2(n4727), .A(n4726), .B(n4725), .ZN(U3086)
         );
  INV_X1 U5885 ( .A(n4778), .ZN(n4729) );
  NAND2_X1 U5886 ( .A1(n4729), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4774) );
  NAND2_X1 U5887 ( .A1(n4774), .A2(n6339), .ZN(n6535) );
  NAND2_X1 U5888 ( .A1(n6293), .A2(n4736), .ZN(n4730) );
  OAI21_X1 U5889 ( .B1(n6535), .B2(n4730), .A(n6536), .ZN(n4741) );
  INV_X1 U5890 ( .A(n4741), .ZN(n4734) );
  NAND2_X1 U5891 ( .A1(n4375), .A2(n5359), .ZN(n5154) );
  INV_X1 U5892 ( .A(n4731), .ZN(n4732) );
  NAND2_X1 U5893 ( .A1(n4732), .A2(n6544), .ZN(n6573) );
  OAI21_X1 U5894 ( .B1(n4895), .B2(n3690), .A(n6573), .ZN(n4740) );
  NAND2_X1 U5895 ( .A1(n5160), .A2(n6544), .ZN(n4890) );
  INV_X1 U5896 ( .A(n4890), .ZN(n4733) );
  AOI22_X1 U5897 ( .A1(n4734), .A2(n4740), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4733), .ZN(n6578) );
  INV_X1 U5898 ( .A(n6575), .ZN(n4760) );
  AND2_X1 U5899 ( .A1(n4735), .A2(n4942), .ZN(n5151) );
  NAND2_X1 U5900 ( .A1(n5151), .A2(n4736), .ZN(n4737) );
  OAI22_X1 U5901 ( .A1(n4911), .A2(n6573), .B1(n4978), .B2(n6571), .ZN(n4738)
         );
  AOI21_X1 U5902 ( .B1(n6315), .B2(n4760), .A(n4738), .ZN(n4743) );
  AOI21_X1 U5903 ( .B1(n6343), .B2(n4890), .A(n6342), .ZN(n4739) );
  OAI21_X1 U5904 ( .B1(n4741), .B2(n4740), .A(n4739), .ZN(n6581) );
  NAND2_X1 U5905 ( .A1(n6581), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4742) );
  OAI211_X1 U5906 ( .C1(n6578), .C2(n6318), .A(n4743), .B(n4742), .ZN(U3048)
         );
  OAI22_X1 U5907 ( .A1(n4900), .A2(n6573), .B1(n4973), .B2(n6571), .ZN(n4744)
         );
  AOI21_X1 U5908 ( .B1(n6311), .B2(n4760), .A(n4744), .ZN(n4746) );
  NAND2_X1 U5909 ( .A1(n6581), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4745) );
  OAI211_X1 U5910 ( .C1(n6578), .C2(n6314), .A(n4746), .B(n4745), .ZN(U3047)
         );
  OAI22_X1 U5911 ( .A1(n4919), .A2(n6573), .B1(n4968), .B2(n6571), .ZN(n4747)
         );
  AOI21_X1 U5912 ( .B1(n6307), .B2(n4760), .A(n4747), .ZN(n4749) );
  NAND2_X1 U5913 ( .A1(n6581), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4748) );
  OAI211_X1 U5914 ( .C1(n6578), .C2(n6310), .A(n4749), .B(n4748), .ZN(U3046)
         );
  OAI22_X1 U5915 ( .A1(n4929), .A2(n6573), .B1(n6352), .B2(n6571), .ZN(n4750)
         );
  AOI21_X1 U5916 ( .B1(n6337), .B2(n4760), .A(n4750), .ZN(n4752) );
  NAND2_X1 U5917 ( .A1(n6581), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4751) );
  OAI211_X1 U5918 ( .C1(n6578), .C2(n6303), .A(n4752), .B(n4751), .ZN(U3044)
         );
  OAI22_X1 U5919 ( .A1(n4904), .A2(n6573), .B1(n4963), .B2(n6571), .ZN(n4753)
         );
  AOI21_X1 U5920 ( .B1(n6323), .B2(n4760), .A(n4753), .ZN(n4755) );
  NAND2_X1 U5921 ( .A1(n6581), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4754) );
  OAI211_X1 U5922 ( .C1(n6578), .C2(n6326), .A(n4755), .B(n4754), .ZN(U3050)
         );
  OAI22_X1 U5923 ( .A1(n4923), .A2(n6573), .B1(n6381), .B2(n6571), .ZN(n4756)
         );
  AOI21_X1 U5924 ( .B1(n6377), .B2(n4760), .A(n4756), .ZN(n4758) );
  NAND2_X1 U5925 ( .A1(n6581), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4757) );
  OAI211_X1 U5926 ( .C1(n6578), .C2(n6322), .A(n4758), .B(n4757), .ZN(U3049)
         );
  OAI22_X1 U5927 ( .A1(n4915), .A2(n6573), .B1(n6400), .B2(n6571), .ZN(n4759)
         );
  AOI21_X1 U5928 ( .B1(n6392), .B2(n4760), .A(n4759), .ZN(n4762) );
  NAND2_X1 U5929 ( .A1(n6581), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4761) );
  OAI211_X1 U5930 ( .C1(n6578), .C2(n6334), .A(n4762), .B(n4761), .ZN(U3051)
         );
  INV_X1 U5931 ( .A(n4763), .ZN(n6014) );
  AOI21_X1 U5932 ( .B1(n6197), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4764), 
        .ZN(n4765) );
  OAI21_X1 U5933 ( .B1(n6017), .B2(n6191), .A(n4765), .ZN(n4766) );
  AOI21_X1 U5934 ( .B1(n6014), .B2(n6186), .A(n4766), .ZN(n4767) );
  OAI21_X1 U5935 ( .B1(n6193), .B2(n4768), .A(n4767), .ZN(U2981) );
  NAND3_X1 U5936 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n4769), .ZN(n4809) );
  NOR2_X1 U5937 ( .A1(n6408), .A2(n4809), .ZN(n4770) );
  INV_X1 U5938 ( .A(n4770), .ZN(n4802) );
  INV_X1 U5939 ( .A(n4809), .ZN(n4773) );
  AOI21_X1 U5940 ( .B1(n4771), .B2(n4937), .A(n4770), .ZN(n4776) );
  NAND3_X1 U5941 ( .A1(n6536), .A2(n4776), .A3(n4774), .ZN(n4772) );
  OAI211_X1 U5942 ( .C1(n6536), .C2(n4773), .A(n6297), .B(n4772), .ZN(n4799)
         );
  NAND2_X1 U5943 ( .A1(n4897), .A2(n4774), .ZN(n4775) );
  OAI22_X1 U5944 ( .A1(n4776), .A2(n4775), .B1(n6560), .B2(n4809), .ZN(n4798)
         );
  AOI22_X1 U5945 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4799), .B1(n6355), 
        .B2(n4798), .ZN(n4780) );
  NOR2_X2 U5946 ( .A1(n4778), .A2(n4777), .ZN(n4845) );
  AOI22_X1 U5947 ( .A1(n6304), .A2(n4845), .B1(n4856), .B2(n6354), .ZN(n4779)
         );
  OAI211_X1 U5948 ( .C1(n6574), .C2(n4802), .A(n4780), .B(n4779), .ZN(U3125)
         );
  AOI22_X1 U5949 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4799), .B1(n6385), 
        .B2(n4798), .ZN(n4782) );
  AOI22_X1 U5950 ( .A1(n6383), .A2(n4845), .B1(n4856), .B2(n6323), .ZN(n4781)
         );
  OAI211_X1 U5951 ( .C1(n4904), .C2(n4802), .A(n4782), .B(n4781), .ZN(U3130)
         );
  AOI22_X1 U5952 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4799), .B1(n6395), 
        .B2(n4798), .ZN(n4784) );
  AOI22_X1 U5953 ( .A1(n6330), .A2(n4845), .B1(n4856), .B2(n6392), .ZN(n4783)
         );
  OAI211_X1 U5954 ( .C1(n4915), .C2(n4802), .A(n4784), .B(n4783), .ZN(U3131)
         );
  AOI22_X1 U5955 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4799), .B1(n6349), 
        .B2(n4798), .ZN(n4786) );
  AOI22_X1 U5956 ( .A1(n6292), .A2(n4845), .B1(n4856), .B2(n6337), .ZN(n4785)
         );
  OAI211_X1 U5957 ( .C1(n4929), .C2(n4802), .A(n4786), .B(n4785), .ZN(U3124)
         );
  NAND2_X1 U5958 ( .A1(n4553), .A2(n4788), .ZN(n4789) );
  AND2_X1 U5959 ( .A1(n4787), .A2(n4789), .ZN(n6042) );
  INV_X1 U5960 ( .A(n6042), .ZN(n4791) );
  INV_X1 U5961 ( .A(DATAI_6_), .ZN(n6120) );
  OAI222_X1 U5962 ( .A1(n4791), .A2(n6047), .B1(n5505), .B2(n4790), .C1(n5329), 
        .C2(n6120), .ZN(U2885) );
  AOI22_X1 U5963 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4799), .B1(n6360), 
        .B2(n4798), .ZN(n4793) );
  AOI22_X1 U5964 ( .A1(n6359), .A2(n4845), .B1(n4856), .B2(n6307), .ZN(n4792)
         );
  OAI211_X1 U5965 ( .C1(n4919), .C2(n4802), .A(n4793), .B(n4792), .ZN(U3126)
         );
  AOI22_X1 U5966 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4799), .B1(n6366), 
        .B2(n4798), .ZN(n4795) );
  AOI22_X1 U5967 ( .A1(n6365), .A2(n4845), .B1(n4856), .B2(n6311), .ZN(n4794)
         );
  OAI211_X1 U5968 ( .C1(n4900), .C2(n4802), .A(n4795), .B(n4794), .ZN(U3127)
         );
  AOI22_X1 U5969 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4799), .B1(n6372), 
        .B2(n4798), .ZN(n4797) );
  AOI22_X1 U5970 ( .A1(n6371), .A2(n4845), .B1(n4856), .B2(n6315), .ZN(n4796)
         );
  OAI211_X1 U5971 ( .C1(n4911), .C2(n4802), .A(n4797), .B(n4796), .ZN(U3128)
         );
  AOI22_X1 U5972 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4799), .B1(n6378), 
        .B2(n4798), .ZN(n4801) );
  AOI22_X1 U5973 ( .A1(n6319), .A2(n4845), .B1(n4856), .B2(n6377), .ZN(n4800)
         );
  OAI211_X1 U5974 ( .C1(n4923), .C2(n4802), .A(n4801), .B(n4800), .ZN(U3129)
         );
  AOI22_X1 U5975 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6238), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n4803) );
  OAI21_X1 U5976 ( .B1(n5998), .B2(n6191), .A(n4803), .ZN(n4804) );
  AOI21_X1 U5977 ( .B1(n6042), .B2(n6186), .A(n4804), .ZN(n4805) );
  OAI21_X1 U5978 ( .B1(n4806), .B2(n6193), .A(n4805), .ZN(U2980) );
  INV_X1 U5979 ( .A(n4845), .ZN(n4822) );
  AOI21_X1 U5980 ( .B1(n4822), .B2(n6388), .A(n6561), .ZN(n4808) );
  AOI211_X1 U5981 ( .C1(n4937), .C2(n4936), .A(n6343), .B(n4808), .ZN(n4812)
         );
  NOR2_X1 U5982 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4809), .ZN(n4844)
         );
  INV_X1 U5983 ( .A(n4855), .ZN(n5157) );
  OAI211_X1 U5984 ( .C1(n6718), .C2(n4844), .A(n5157), .B(n4810), .ZN(n4811)
         );
  NAND2_X1 U5985 ( .A1(n4849), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4818)
         );
  NAND2_X1 U5986 ( .A1(n4853), .A2(n4937), .ZN(n4815) );
  NAND2_X1 U5987 ( .A1(n4813), .A2(n6256), .ZN(n4814) );
  AND2_X1 U5988 ( .A1(n4815), .A2(n4814), .ZN(n4826) );
  OAI22_X1 U5989 ( .A1(n4822), .A2(n6576), .B1(n4826), .B2(n6577), .ZN(n4816)
         );
  AOI21_X1 U5990 ( .B1(n6353), .B2(n4844), .A(n4816), .ZN(n4817) );
  OAI211_X1 U5991 ( .C1(n6388), .C2(n6572), .A(n4818), .B(n4817), .ZN(U3117)
         );
  NAND2_X1 U5992 ( .A1(n4849), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4821)
         );
  OAI22_X1 U5993 ( .A1(n4822), .A2(n6288), .B1(n6334), .B2(n4826), .ZN(n4819)
         );
  AOI21_X1 U5994 ( .B1(n6391), .B2(n4844), .A(n4819), .ZN(n4820) );
  OAI211_X1 U5995 ( .C1(n6388), .C2(n6400), .A(n4821), .B(n4820), .ZN(U3123)
         );
  NAND2_X1 U5996 ( .A1(n4849), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4825)
         );
  OAI22_X1 U5997 ( .A1(n4822), .A2(n6389), .B1(n6326), .B2(n4826), .ZN(n4823)
         );
  AOI21_X1 U5998 ( .B1(n6382), .B2(n4844), .A(n4823), .ZN(n4824) );
  OAI211_X1 U5999 ( .C1(n6388), .C2(n4963), .A(n4825), .B(n4824), .ZN(U3122)
         );
  INV_X1 U6000 ( .A(n4826), .ZN(n4843) );
  NAND2_X1 U6001 ( .A1(n6366), .A2(n4843), .ZN(n4828) );
  AOI22_X1 U6002 ( .A1(n4845), .A2(n6311), .B1(n6364), .B2(n4844), .ZN(n4827)
         );
  OAI211_X1 U6003 ( .C1(n6388), .C2(n4973), .A(n4828), .B(n4827), .ZN(n4829)
         );
  AOI21_X1 U6004 ( .B1(n4849), .B2(INSTQUEUE_REG_12__3__SCAN_IN), .A(n4829), 
        .ZN(n4830) );
  INV_X1 U6005 ( .A(n4830), .ZN(U3119) );
  NAND2_X1 U6006 ( .A1(n6360), .A2(n4843), .ZN(n4832) );
  AOI22_X1 U6007 ( .A1(n4845), .A2(n6307), .B1(n6358), .B2(n4844), .ZN(n4831)
         );
  OAI211_X1 U6008 ( .C1(n6388), .C2(n4968), .A(n4832), .B(n4831), .ZN(n4833)
         );
  AOI21_X1 U6009 ( .B1(n4849), .B2(INSTQUEUE_REG_12__2__SCAN_IN), .A(n4833), 
        .ZN(n4834) );
  INV_X1 U6010 ( .A(n4834), .ZN(U3118) );
  NAND2_X1 U6011 ( .A1(n6349), .A2(n4843), .ZN(n4836) );
  AOI22_X1 U6012 ( .A1(n4845), .A2(n6337), .B1(n6336), .B2(n4844), .ZN(n4835)
         );
  OAI211_X1 U6013 ( .C1(n6388), .C2(n6352), .A(n4836), .B(n4835), .ZN(n4837)
         );
  AOI21_X1 U6014 ( .B1(n4849), .B2(INSTQUEUE_REG_12__0__SCAN_IN), .A(n4837), 
        .ZN(n4838) );
  INV_X1 U6015 ( .A(n4838), .ZN(U3116) );
  NAND2_X1 U6016 ( .A1(n6378), .A2(n4843), .ZN(n4840) );
  AOI22_X1 U6017 ( .A1(n4845), .A2(n6377), .B1(n6376), .B2(n4844), .ZN(n4839)
         );
  OAI211_X1 U6018 ( .C1(n6388), .C2(n6381), .A(n4840), .B(n4839), .ZN(n4841)
         );
  AOI21_X1 U6019 ( .B1(n4849), .B2(INSTQUEUE_REG_12__5__SCAN_IN), .A(n4841), 
        .ZN(n4842) );
  INV_X1 U6020 ( .A(n4842), .ZN(U3121) );
  NAND2_X1 U6021 ( .A1(n6372), .A2(n4843), .ZN(n4847) );
  AOI22_X1 U6022 ( .A1(n4845), .A2(n6315), .B1(n6370), .B2(n4844), .ZN(n4846)
         );
  OAI211_X1 U6023 ( .C1(n6388), .C2(n4978), .A(n4847), .B(n4846), .ZN(n4848)
         );
  AOI21_X1 U6024 ( .B1(n4849), .B2(INSTQUEUE_REG_12__4__SCAN_IN), .A(n4848), 
        .ZN(n4850) );
  INV_X1 U6025 ( .A(n4850), .ZN(U3120) );
  NOR3_X1 U6026 ( .A1(n4851), .A2(n5156), .A3(n6544), .ZN(n4852) );
  AOI21_X1 U6027 ( .B1(n4853), .B2(n6290), .A(n4852), .ZN(n4882) );
  NOR2_X1 U6028 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4854), .ZN(n4875)
         );
  AOI211_X1 U6029 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n5156), .A(n4855), .B(
        n4893), .ZN(n6263) );
  NAND2_X1 U6030 ( .A1(n6544), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5161) );
  OAI211_X1 U6031 ( .C1(n4875), .C2(n6718), .A(n6263), .B(n5161), .ZN(n4859)
         );
  NAND3_X1 U6032 ( .A1(n4883), .A2(n6536), .A3(n4885), .ZN(n4857) );
  AOI22_X1 U6033 ( .A1(n4857), .A2(n5152), .B1(n6290), .B2(n6540), .ZN(n4858)
         );
  NAND2_X1 U6034 ( .A1(n4888), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4862)
         );
  OAI22_X1 U6035 ( .A1(n4883), .A2(n4978), .B1(n6375), .B2(n4885), .ZN(n4860)
         );
  AOI21_X1 U6036 ( .B1(n6370), .B2(n4875), .A(n4860), .ZN(n4861) );
  OAI211_X1 U6037 ( .C1(n4882), .C2(n6318), .A(n4862), .B(n4861), .ZN(U3136)
         );
  NAND2_X1 U6038 ( .A1(n4888), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4865)
         );
  OAI22_X1 U6039 ( .A1(n4883), .A2(n4968), .B1(n6363), .B2(n4885), .ZN(n4863)
         );
  AOI21_X1 U6040 ( .B1(n6358), .B2(n4875), .A(n4863), .ZN(n4864) );
  OAI211_X1 U6041 ( .C1(n4882), .C2(n6310), .A(n4865), .B(n4864), .ZN(U3134)
         );
  NAND2_X1 U6042 ( .A1(n4888), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4868)
         );
  OAI22_X1 U6043 ( .A1(n4883), .A2(n6381), .B1(n6278), .B2(n4885), .ZN(n4866)
         );
  AOI21_X1 U6044 ( .B1(n6376), .B2(n4875), .A(n4866), .ZN(n4867) );
  OAI211_X1 U6045 ( .C1(n4882), .C2(n6322), .A(n4868), .B(n4867), .ZN(U3137)
         );
  NAND2_X1 U6046 ( .A1(n4888), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4871)
         );
  OAI22_X1 U6047 ( .A1(n4883), .A2(n4973), .B1(n6369), .B2(n4885), .ZN(n4869)
         );
  AOI21_X1 U6048 ( .B1(n6364), .B2(n4875), .A(n4869), .ZN(n4870) );
  OAI211_X1 U6049 ( .C1(n4882), .C2(n6314), .A(n4871), .B(n4870), .ZN(U3135)
         );
  NAND2_X1 U6050 ( .A1(n4888), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4874)
         );
  OAI22_X1 U6051 ( .A1(n4883), .A2(n6352), .B1(n6267), .B2(n4885), .ZN(n4872)
         );
  AOI21_X1 U6052 ( .B1(n6336), .B2(n4875), .A(n4872), .ZN(n4873) );
  OAI211_X1 U6053 ( .C1(n4882), .C2(n6303), .A(n4874), .B(n4873), .ZN(U3132)
         );
  OAI22_X1 U6054 ( .A1(n4883), .A2(n6400), .B1(n6334), .B2(n4882), .ZN(n4877)
         );
  INV_X1 U6055 ( .A(n4875), .ZN(n4884) );
  OAI22_X1 U6056 ( .A1(n4885), .A2(n6288), .B1(n4915), .B2(n4884), .ZN(n4876)
         );
  AOI211_X1 U6057 ( .C1(n4888), .C2(INSTQUEUE_REG_14__7__SCAN_IN), .A(n4877), 
        .B(n4876), .ZN(n4878) );
  INV_X1 U6058 ( .A(n4878), .ZN(U3139) );
  OAI22_X1 U6059 ( .A1(n4883), .A2(n6572), .B1(n4882), .B2(n6577), .ZN(n4880)
         );
  OAI22_X1 U6060 ( .A1(n4885), .A2(n6576), .B1(n6574), .B2(n4884), .ZN(n4879)
         );
  AOI211_X1 U6061 ( .C1(n4888), .C2(INSTQUEUE_REG_14__1__SCAN_IN), .A(n4880), 
        .B(n4879), .ZN(n4881) );
  INV_X1 U6062 ( .A(n4881), .ZN(U3133) );
  OAI22_X1 U6063 ( .A1(n4883), .A2(n4963), .B1(n6326), .B2(n4882), .ZN(n4887)
         );
  OAI22_X1 U6064 ( .A1(n4885), .A2(n6389), .B1(n4904), .B2(n4884), .ZN(n4886)
         );
  AOI211_X1 U6065 ( .C1(n4888), .C2(INSTQUEUE_REG_14__6__SCAN_IN), .A(n4887), 
        .B(n4886), .ZN(n4889) );
  INV_X1 U6066 ( .A(n4889), .ZN(U3138) );
  NOR2_X1 U6067 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4890), .ZN(n4899)
         );
  INV_X1 U6068 ( .A(n4935), .ZN(n4891) );
  OAI21_X1 U6069 ( .B1(n4891), .B2(n4932), .A(n5152), .ZN(n4892) );
  AOI21_X1 U6070 ( .B1(n4892), .B2(n4895), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4894) );
  AOI211_X1 U6071 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n5156), .A(n6256), .B(
        n4893), .ZN(n5166) );
  NAND2_X1 U6072 ( .A1(n4927), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4903) );
  INV_X1 U6073 ( .A(n4895), .ZN(n4898) );
  NOR3_X1 U6074 ( .A1(n5157), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5156), 
        .ZN(n4896) );
  AOI21_X1 U6075 ( .B1(n4898), .B2(n4897), .A(n4896), .ZN(n4930) );
  INV_X1 U6076 ( .A(n4899), .ZN(n4928) );
  OAI22_X1 U6077 ( .A1(n6314), .A2(n4930), .B1(n4900), .B2(n4928), .ZN(n4901)
         );
  AOI21_X1 U6078 ( .B1(n6311), .B2(n4932), .A(n4901), .ZN(n4902) );
  OAI211_X1 U6079 ( .C1(n4935), .C2(n4973), .A(n4903), .B(n4902), .ZN(U3039)
         );
  NAND2_X1 U6080 ( .A1(n4927), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4907) );
  OAI22_X1 U6081 ( .A1(n6326), .A2(n4930), .B1(n4904), .B2(n4928), .ZN(n4905)
         );
  AOI21_X1 U6082 ( .B1(n6323), .B2(n4932), .A(n4905), .ZN(n4906) );
  OAI211_X1 U6083 ( .C1(n4935), .C2(n4963), .A(n4907), .B(n4906), .ZN(U3042)
         );
  NAND2_X1 U6084 ( .A1(n4927), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4910) );
  OAI22_X1 U6085 ( .A1(n6574), .A2(n4928), .B1(n4930), .B2(n6577), .ZN(n4908)
         );
  AOI21_X1 U6086 ( .B1(n6354), .B2(n4932), .A(n4908), .ZN(n4909) );
  OAI211_X1 U6087 ( .C1(n4935), .C2(n6572), .A(n4910), .B(n4909), .ZN(U3037)
         );
  NAND2_X1 U6088 ( .A1(n4927), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4914) );
  OAI22_X1 U6089 ( .A1(n6318), .A2(n4930), .B1(n4911), .B2(n4928), .ZN(n4912)
         );
  AOI21_X1 U6090 ( .B1(n6315), .B2(n4932), .A(n4912), .ZN(n4913) );
  OAI211_X1 U6091 ( .C1(n4935), .C2(n4978), .A(n4914), .B(n4913), .ZN(U3040)
         );
  NAND2_X1 U6092 ( .A1(n4927), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4918) );
  OAI22_X1 U6093 ( .A1(n6334), .A2(n4930), .B1(n4915), .B2(n4928), .ZN(n4916)
         );
  AOI21_X1 U6094 ( .B1(n6392), .B2(n4932), .A(n4916), .ZN(n4917) );
  OAI211_X1 U6095 ( .C1(n4935), .C2(n6400), .A(n4918), .B(n4917), .ZN(U3043)
         );
  NAND2_X1 U6096 ( .A1(n4927), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4922) );
  OAI22_X1 U6097 ( .A1(n6310), .A2(n4930), .B1(n4919), .B2(n4928), .ZN(n4920)
         );
  AOI21_X1 U6098 ( .B1(n6307), .B2(n4932), .A(n4920), .ZN(n4921) );
  OAI211_X1 U6099 ( .C1(n4935), .C2(n4968), .A(n4922), .B(n4921), .ZN(U3038)
         );
  NAND2_X1 U6100 ( .A1(n4927), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4926) );
  OAI22_X1 U6101 ( .A1(n6322), .A2(n4930), .B1(n4923), .B2(n4928), .ZN(n4924)
         );
  AOI21_X1 U6102 ( .B1(n6377), .B2(n4932), .A(n4924), .ZN(n4925) );
  OAI211_X1 U6103 ( .C1(n4935), .C2(n6381), .A(n4926), .B(n4925), .ZN(U3041)
         );
  NAND2_X1 U6104 ( .A1(n4927), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4934) );
  OAI22_X1 U6105 ( .A1(n6303), .A2(n4930), .B1(n4929), .B2(n4928), .ZN(n4931)
         );
  AOI21_X1 U6106 ( .B1(n6337), .B2(n4932), .A(n4931), .ZN(n4933) );
  OAI211_X1 U6107 ( .C1(n4935), .C2(n6352), .A(n4934), .B(n4933), .ZN(U3036)
         );
  INV_X1 U6108 ( .A(n4949), .ZN(n4941) );
  NOR2_X1 U6109 ( .A1(n3690), .A2(n4936), .ZN(n6289) );
  NAND2_X1 U6110 ( .A1(n4937), .A2(n6289), .ZN(n4939) );
  NOR2_X1 U6111 ( .A1(n6408), .A2(n4946), .ZN(n4982) );
  INV_X1 U6112 ( .A(n4982), .ZN(n4938) );
  NAND2_X1 U6113 ( .A1(n4939), .A2(n4938), .ZN(n4948) );
  INV_X1 U6114 ( .A(n4946), .ZN(n4940) );
  AOI22_X1 U6115 ( .A1(n4941), .A2(n4948), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4940), .ZN(n4953) );
  NOR2_X2 U6116 ( .A1(n4943), .A2(n4942), .ZN(n6283) );
  INV_X1 U6117 ( .A(n6283), .ZN(n4944) );
  OAI22_X1 U6118 ( .A1(n4944), .A2(n6267), .B1(n6352), .B2(n4984), .ZN(n4945)
         );
  AOI21_X1 U6119 ( .B1(n6336), .B2(n4982), .A(n4945), .ZN(n4951) );
  AOI21_X1 U6120 ( .B1(n6343), .B2(n4946), .A(n6342), .ZN(n4947) );
  OAI21_X1 U6121 ( .B1(n4949), .B2(n4948), .A(n4947), .ZN(n4952) );
  NAND2_X1 U6122 ( .A1(n4952), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4950) );
  OAI211_X1 U6123 ( .C1(n4953), .C2(n6303), .A(n4951), .B(n4950), .ZN(U3060)
         );
  INV_X1 U6124 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U6125 ( .A1(n6283), .A2(n6392), .B1(n6391), .B2(n4982), .ZN(n4954)
         );
  OAI21_X1 U6126 ( .B1(n6400), .B2(n4984), .A(n4954), .ZN(n4955) );
  AOI21_X1 U6127 ( .B1(n4986), .B2(n6395), .A(n4955), .ZN(n4956) );
  OAI21_X1 U6128 ( .B1(n4989), .B2(n4957), .A(n4956), .ZN(U3067) );
  INV_X1 U6129 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U6130 ( .A1(n6283), .A2(n6354), .B1(n6353), .B2(n4982), .ZN(n4958)
         );
  OAI21_X1 U6131 ( .B1(n6572), .B2(n4984), .A(n4958), .ZN(n4959) );
  AOI21_X1 U6132 ( .B1(n4986), .B2(n6355), .A(n4959), .ZN(n4960) );
  OAI21_X1 U6133 ( .B1(n4989), .B2(n4961), .A(n4960), .ZN(U3061) );
  INV_X1 U6134 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4966) );
  AOI22_X1 U6135 ( .A1(n6283), .A2(n6323), .B1(n6382), .B2(n4982), .ZN(n4962)
         );
  OAI21_X1 U6136 ( .B1(n4963), .B2(n4984), .A(n4962), .ZN(n4964) );
  AOI21_X1 U6137 ( .B1(n4986), .B2(n6385), .A(n4964), .ZN(n4965) );
  OAI21_X1 U6138 ( .B1(n4989), .B2(n4966), .A(n4965), .ZN(U3066) );
  INV_X1 U6139 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4971) );
  AOI22_X1 U6140 ( .A1(n6283), .A2(n6307), .B1(n6358), .B2(n4982), .ZN(n4967)
         );
  OAI21_X1 U6141 ( .B1(n4968), .B2(n4984), .A(n4967), .ZN(n4969) );
  AOI21_X1 U6142 ( .B1(n4986), .B2(n6360), .A(n4969), .ZN(n4970) );
  OAI21_X1 U6143 ( .B1(n4989), .B2(n4971), .A(n4970), .ZN(U3062) );
  INV_X1 U6144 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4976) );
  AOI22_X1 U6145 ( .A1(n6283), .A2(n6311), .B1(n6364), .B2(n4982), .ZN(n4972)
         );
  OAI21_X1 U6146 ( .B1(n4973), .B2(n4984), .A(n4972), .ZN(n4974) );
  AOI21_X1 U6147 ( .B1(n4986), .B2(n6366), .A(n4974), .ZN(n4975) );
  OAI21_X1 U6148 ( .B1(n4989), .B2(n4976), .A(n4975), .ZN(U3063) );
  INV_X1 U6149 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4981) );
  AOI22_X1 U6150 ( .A1(n6283), .A2(n6315), .B1(n6370), .B2(n4982), .ZN(n4977)
         );
  OAI21_X1 U6151 ( .B1(n4978), .B2(n4984), .A(n4977), .ZN(n4979) );
  AOI21_X1 U6152 ( .B1(n4986), .B2(n6372), .A(n4979), .ZN(n4980) );
  OAI21_X1 U6153 ( .B1(n4989), .B2(n4981), .A(n4980), .ZN(U3064) );
  INV_X1 U6154 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4988) );
  AOI22_X1 U6155 ( .A1(n6283), .A2(n6377), .B1(n6376), .B2(n4982), .ZN(n4983)
         );
  OAI21_X1 U6156 ( .B1(n6381), .B2(n4984), .A(n4983), .ZN(n4985) );
  AOI21_X1 U6157 ( .B1(n4986), .B2(n6378), .A(n4985), .ZN(n4987) );
  OAI21_X1 U6158 ( .B1(n4989), .B2(n4988), .A(n4987), .ZN(U3065) );
  NOR2_X1 U6159 ( .A1(n4996), .A2(n4990), .ZN(n4991) );
  OR2_X1 U6160 ( .A1(n4991), .A2(n6001), .ZN(n6033) );
  NOR2_X1 U6161 ( .A1(n4996), .A2(n3634), .ZN(n6023) );
  NAND3_X1 U6162 ( .A1(n6065), .A2(n5354), .A3(n4992), .ZN(n4993) );
  AND2_X1 U6163 ( .A1(n4994), .A2(n4993), .ZN(n4995) );
  INV_X1 U6164 ( .A(n6190), .ZN(n4999) );
  NAND2_X1 U6165 ( .A1(n5999), .A2(n4999), .ZN(n5001) );
  NAND2_X1 U6166 ( .A1(n5993), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5000)
         );
  OAI211_X1 U6167 ( .C1(n6004), .C2(n3524), .A(n5001), .B(n5000), .ZN(n5005)
         );
  AOI21_X1 U6168 ( .B1(n6009), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5003) );
  OAI211_X1 U6169 ( .C1(REIP_REG_1__SCAN_IN), .C2(n6026), .A(
        REIP_REG_2__SCAN_IN), .B(n5987), .ZN(n5091) );
  INV_X1 U6170 ( .A(n5091), .ZN(n5002) );
  OAI22_X1 U6171 ( .A1(n6031), .A2(n6237), .B1(n5003), .B2(n5002), .ZN(n5004)
         );
  AOI211_X1 U6172 ( .C1(n5006), .C2(n6023), .A(n5005), .B(n5004), .ZN(n5007)
         );
  OAI21_X1 U6173 ( .B1(n5008), .B2(n5367), .A(n5007), .ZN(U2825) );
  INV_X1 U6174 ( .A(n5009), .ZN(n5010) );
  AOI21_X1 U6175 ( .B1(n5011), .B2(n4787), .A(n5010), .ZN(n5985) );
  INV_X1 U6176 ( .A(n5985), .ZN(n5017) );
  OAI21_X1 U6177 ( .B1(n4498), .B2(n5013), .A(n5012), .ZN(n5014) );
  AND2_X1 U6178 ( .A1(n5014), .A2(n5030), .ZN(n6218) );
  AOI22_X1 U6179 ( .A1(n6040), .A2(n6218), .B1(n5501), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5015) );
  OAI21_X1 U6180 ( .B1(n5017), .B2(n5819), .A(n5015), .ZN(U2852) );
  AOI22_X1 U6181 ( .A1(n5514), .A2(DATAI_7_), .B1(n6061), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n5016) );
  OAI21_X1 U6182 ( .B1(n5017), .B2(n6047), .A(n5016), .ZN(U2884) );
  XOR2_X1 U6183 ( .A(n5019), .B(n5018), .Z(n6223) );
  INV_X1 U6184 ( .A(n6223), .ZN(n5023) );
  NAND2_X1 U6185 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5020)
         );
  NAND2_X1 U6186 ( .A1(n6238), .A2(REIP_REG_7__SCAN_IN), .ZN(n6219) );
  OAI211_X1 U6187 ( .C1(n6191), .C2(n5992), .A(n5020), .B(n6219), .ZN(n5021)
         );
  AOI21_X1 U6188 ( .B1(n5985), .B2(n6186), .A(n5021), .ZN(n5022) );
  OAI21_X1 U6189 ( .B1(n5023), .B2(n6193), .A(n5022), .ZN(U2979) );
  CLKBUF_X1 U6190 ( .A(n5024), .Z(n5026) );
  XNOR2_X1 U6191 ( .A(n5026), .B(n5025), .ZN(n5046) );
  NAND2_X1 U6192 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5028) );
  NOR2_X1 U6193 ( .A1(n5028), .A2(n5027), .ZN(n6217) );
  AOI21_X1 U6194 ( .B1(n6225), .B2(n5035), .A(n5111), .ZN(n5038) );
  AND2_X1 U6195 ( .A1(n5030), .A2(n5029), .ZN(n5031) );
  OR2_X1 U6196 ( .A1(n5031), .A2(n5073), .ZN(n5058) );
  NAND2_X1 U6197 ( .A1(n5592), .A2(REIP_REG_8__SCAN_IN), .ZN(n5043) );
  OAI21_X1 U6198 ( .B1(n3628), .B2(n5058), .A(n5043), .ZN(n5037) );
  INV_X1 U6199 ( .A(n5214), .ZN(n5034) );
  AOI22_X1 U6200 ( .A1(n5034), .A2(n5033), .B1(n5212), .B2(n5032), .ZN(n6226)
         );
  NOR2_X1 U6201 ( .A1(n6226), .A2(n5035), .ZN(n5036) );
  AOI211_X1 U6202 ( .C1(n6217), .C2(n5038), .A(n5037), .B(n5036), .ZN(n5039)
         );
  OAI21_X1 U6203 ( .B1(n5717), .B2(n5046), .A(n5039), .ZN(U3010) );
  AOI21_X1 U6204 ( .B1(n5041), .B2(n5009), .A(n5040), .ZN(n5047) );
  NAND2_X1 U6205 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5042)
         );
  OAI211_X1 U6206 ( .C1(n6191), .C2(n5062), .A(n5043), .B(n5042), .ZN(n5044)
         );
  AOI21_X1 U6207 ( .B1(n5047), .B2(n6186), .A(n5044), .ZN(n5045) );
  OAI21_X1 U6208 ( .B1(n6193), .B2(n5046), .A(n5045), .ZN(U2978) );
  INV_X1 U6209 ( .A(n5047), .ZN(n5067) );
  AOI22_X1 U6210 ( .A1(n5514), .A2(DATAI_8_), .B1(n6061), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5048) );
  OAI21_X1 U6211 ( .B1(n5067), .B2(n6047), .A(n5048), .ZN(U2883) );
  INV_X1 U6212 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5049) );
  OAI222_X1 U6213 ( .A1(n5067), .A2(n5819), .B1(n6045), .B2(n5049), .C1(n5058), 
        .C2(n5817), .ZN(U2851) );
  OAI21_X1 U6214 ( .B1(n5993), .B2(n5999), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5050) );
  OAI21_X1 U6215 ( .B1(n5811), .B2(n6552), .A(n5050), .ZN(n5054) );
  NAND2_X1 U6216 ( .A1(n6023), .A2(n6340), .ZN(n5051) );
  OAI21_X1 U6217 ( .B1(n5052), .B2(n6004), .A(n5051), .ZN(n5053) );
  AOI211_X1 U6218 ( .C1(n6007), .C2(n5055), .A(n5054), .B(n5053), .ZN(n5056)
         );
  OAI21_X1 U6219 ( .B1(n5367), .B2(n6201), .A(n5056), .ZN(U2827) );
  NAND3_X1 U6220 ( .A1(n6009), .A2(REIP_REG_5__SCAN_IN), .A3(n6008), .ZN(n5989) );
  AOI221_X1 U6221 ( .B1(n5057), .B2(n6484), .C1(n5989), .C2(n6484), .A(n5811), 
        .ZN(n5065) );
  NAND2_X1 U6222 ( .A1(n5127), .A2(n5987), .ZN(n5077) );
  OAI22_X1 U6223 ( .A1(n5059), .A2(n6018), .B1(n6031), .B2(n5058), .ZN(n5064)
         );
  NAND2_X1 U6224 ( .A1(n6028), .A2(EBX_REG_8__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U6225 ( .A1(n5987), .A2(n5060), .ZN(n5994) );
  OAI211_X1 U6226 ( .C1(n6037), .C2(n5062), .A(n5061), .B(n5994), .ZN(n5063)
         );
  AOI211_X1 U6227 ( .C1(n5065), .C2(n5077), .A(n5064), .B(n5063), .ZN(n5066)
         );
  OAI21_X1 U6228 ( .B1(n5067), .B2(n5955), .A(n5066), .ZN(U2819) );
  OAI21_X1 U6229 ( .B1(n5040), .B2(n5070), .A(n5069), .ZN(n5117) );
  OR2_X1 U6230 ( .A1(n5073), .A2(n5072), .ZN(n5074) );
  AND2_X1 U6231 ( .A1(n5071), .A2(n5074), .ZN(n6211) );
  AOI22_X1 U6232 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6028), .B1(n6007), .B2(n6211), 
        .ZN(n5075) );
  OAI211_X1 U6233 ( .C1(n6018), .C2(n5076), .A(n5075), .B(n5994), .ZN(n5080)
         );
  INV_X1 U6234 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U6235 ( .A1(n6009), .A2(n5127), .ZN(n5078) );
  INV_X1 U6236 ( .A(n5811), .ZN(n5775) );
  OAI21_X1 U6237 ( .B1(n6486), .B2(n5077), .A(n5775), .ZN(n5128) );
  AOI21_X1 U6238 ( .B1(n6486), .B2(n5078), .A(n5128), .ZN(n5079) );
  AOI211_X1 U6239 ( .C1(n5999), .C2(n5087), .A(n5080), .B(n5079), .ZN(n5081)
         );
  OAI21_X1 U6240 ( .B1(n5117), .B2(n5955), .A(n5081), .ZN(U2818) );
  AOI22_X1 U6241 ( .A1(n6211), .A2(n6040), .B1(EBX_REG_9__SCAN_IN), .B2(n5501), 
        .ZN(n5082) );
  OAI21_X1 U6242 ( .B1(n5117), .B2(n5819), .A(n5082), .ZN(U2850) );
  CLKBUF_X1 U6243 ( .A(n5083), .Z(n5084) );
  XNOR2_X1 U6244 ( .A(n5708), .B(n5113), .ZN(n5085) );
  XNOR2_X1 U6245 ( .A(n5084), .B(n5085), .ZN(n6213) );
  INV_X1 U6246 ( .A(n6193), .ZN(n6185) );
  NAND2_X1 U6247 ( .A1(n6213), .A2(n6185), .ZN(n5089) );
  NAND2_X1 U6248 ( .A1(n6238), .A2(REIP_REG_9__SCAN_IN), .ZN(n6209) );
  OAI21_X1 U6249 ( .B1(n5873), .B2(n5076), .A(n6209), .ZN(n5086) );
  AOI21_X1 U6250 ( .B1(n5868), .B2(n5087), .A(n5086), .ZN(n5088) );
  OAI211_X1 U6251 ( .C1(n6200), .C2(n5117), .A(n5089), .B(n5088), .ZN(U2977)
         );
  AOI21_X1 U6252 ( .B1(n6009), .B2(n6025), .A(n5441), .ZN(n6020) );
  INV_X1 U6253 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6475) );
  INV_X1 U6254 ( .A(n6227), .ZN(n5098) );
  NAND2_X1 U6255 ( .A1(n6009), .A2(n6025), .ZN(n5090) );
  NOR2_X1 U6256 ( .A1(n5091), .A2(n5090), .ZN(n5092) );
  AOI21_X1 U6257 ( .B1(n5993), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5092), 
        .ZN(n5095) );
  INV_X1 U6258 ( .A(n5370), .ZN(n5093) );
  NAND2_X1 U6259 ( .A1(n5999), .A2(n5093), .ZN(n5094) );
  OAI211_X1 U6260 ( .C1(n6004), .C2(n5096), .A(n5095), .B(n5094), .ZN(n5097)
         );
  AOI21_X1 U6261 ( .B1(n6007), .B2(n5098), .A(n5097), .ZN(n5099) );
  OAI21_X1 U6262 ( .B1(n6020), .B2(n6475), .A(n5099), .ZN(n5101) );
  NOR2_X1 U6263 ( .A1(n5375), .A2(n5367), .ZN(n5100) );
  AOI211_X1 U6264 ( .C1(n6023), .C2(n6540), .A(n5101), .B(n5100), .ZN(n5102)
         );
  INV_X1 U6265 ( .A(n5102), .ZN(U2824) );
  CLKBUF_X1 U6266 ( .A(n5103), .Z(n5106) );
  NAND2_X1 U6267 ( .A1(n3005), .A2(n5104), .ZN(n5105) );
  XNOR2_X1 U6268 ( .A(n5106), .B(n5105), .ZN(n5124) );
  OAI21_X1 U6269 ( .B1(n5107), .B2(n5111), .A(n6226), .ZN(n6212) );
  INV_X1 U6270 ( .A(n5108), .ZN(n5139) );
  NAND2_X1 U6271 ( .A1(n5071), .A2(n5109), .ZN(n5110) );
  NAND2_X1 U6272 ( .A1(n5139), .A2(n5110), .ZN(n5197) );
  INV_X1 U6273 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6488) );
  OAI22_X1 U6274 ( .A1(n5197), .A2(n3628), .B1(n6488), .B2(n6192), .ZN(n5115)
         );
  NAND2_X1 U6275 ( .A1(n5111), .A2(n6217), .ZN(n6216) );
  AOI221_X1 U6276 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5113), .C2(n5112), .A(n6216), 
        .ZN(n5114) );
  AOI211_X1 U6277 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6212), .A(n5115), .B(n5114), .ZN(n5116) );
  OAI21_X1 U6278 ( .B1(n5717), .B2(n5124), .A(n5116), .ZN(U3008) );
  INV_X1 U6279 ( .A(DATAI_9_), .ZN(n6631) );
  INV_X1 U6280 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6164) );
  OAI222_X1 U6281 ( .A1(n5117), .A2(n6047), .B1(n5329), .B2(n6631), .C1(n5505), 
        .C2(n6164), .ZN(U2882) );
  INV_X1 U6282 ( .A(n5118), .ZN(n5119) );
  AOI21_X1 U6283 ( .B1(n5119), .B2(n5069), .A(n5136), .ZN(n5125) );
  INV_X1 U6284 ( .A(n5131), .ZN(n5121) );
  AOI22_X1 U6285 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6238), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5120) );
  OAI21_X1 U6286 ( .B1(n6191), .B2(n5121), .A(n5120), .ZN(n5122) );
  AOI21_X1 U6287 ( .B1(n5125), .B2(n6186), .A(n5122), .ZN(n5123) );
  OAI21_X1 U6288 ( .B1(n6193), .B2(n5124), .A(n5123), .ZN(U2976) );
  INV_X1 U6289 ( .A(n5125), .ZN(n5195) );
  AOI22_X1 U6290 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6028), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n5993), .ZN(n5126) );
  OAI211_X1 U6291 ( .C1(n6031), .C2(n5197), .A(n5126), .B(n5994), .ZN(n5130)
         );
  NAND3_X1 U6292 ( .A1(n6009), .A2(REIP_REG_9__SCAN_IN), .A3(n5127), .ZN(n5143) );
  AOI22_X1 U6293 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5128), .B1(n5143), .B2(
        n6488), .ZN(n5129) );
  AOI211_X1 U6294 ( .C1(n5131), .C2(n5999), .A(n5130), .B(n5129), .ZN(n5132)
         );
  OAI21_X1 U6295 ( .B1(n5195), .B2(n5955), .A(n5132), .ZN(U2817) );
  AOI22_X1 U6296 ( .A1(n5514), .A2(DATAI_10_), .B1(n6061), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5133) );
  OAI21_X1 U6297 ( .B1(n5195), .B2(n6047), .A(n5133), .ZN(U2881) );
  OAI21_X1 U6298 ( .B1(n5136), .B2(n5135), .A(n5134), .ZN(n5207) );
  AOI22_X1 U6299 ( .A1(n5514), .A2(DATAI_11_), .B1(n6061), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5137) );
  OAI21_X1 U6300 ( .B1(n5207), .B2(n6047), .A(n5137), .ZN(U2880) );
  INV_X1 U6301 ( .A(n5203), .ZN(n5148) );
  AOI21_X1 U6302 ( .B1(n5140), .B2(n5139), .A(n5138), .ZN(n6203) );
  AOI22_X1 U6303 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6028), .B1(n6007), .B2(n6203), .ZN(n5141) );
  OAI211_X1 U6304 ( .C1(n6018), .C2(n5142), .A(n5141), .B(n5994), .ZN(n5147)
         );
  NOR2_X1 U6305 ( .A1(n6488), .A2(n5143), .ZN(n5145) );
  AOI21_X1 U6306 ( .B1(n5974), .B2(n6009), .A(n5441), .ZN(n5144) );
  INV_X1 U6307 ( .A(n5144), .ZN(n5972) );
  MUX2_X1 U6308 ( .A(n5145), .B(n5972), .S(REIP_REG_11__SCAN_IN), .Z(n5146) );
  AOI211_X1 U6309 ( .C1(n5999), .C2(n5148), .A(n5147), .B(n5146), .ZN(n5149)
         );
  OAI21_X1 U6310 ( .B1(n5207), .B2(n5955), .A(n5149), .ZN(U2816) );
  AOI22_X1 U6311 ( .A1(n6203), .A2(n6040), .B1(EBX_REG_11__SCAN_IN), .B2(n5501), .ZN(n5150) );
  OAI21_X1 U6312 ( .B1(n5207), .B2(n5819), .A(n5150), .ZN(U2848) );
  INV_X1 U6313 ( .A(n5151), .ZN(n6253) );
  NAND3_X1 U6314 ( .A1(n5159), .A2(n6536), .A3(n6399), .ZN(n5153) );
  NAND2_X1 U6315 ( .A1(n5153), .A2(n5152), .ZN(n5164) );
  INV_X1 U6316 ( .A(n5154), .ZN(n5155) );
  NOR3_X1 U6317 ( .A1(n5157), .A2(n5156), .A3(n6544), .ZN(n5158) );
  NAND2_X1 U6318 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5160), .ZN(n6346) );
  NOR2_X1 U6319 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6346), .ZN(n5189)
         );
  INV_X1 U6320 ( .A(n6341), .ZN(n5163) );
  INV_X1 U6321 ( .A(n5161), .ZN(n5162) );
  AOI21_X1 U6322 ( .B1(n5164), .B2(n5163), .A(n5162), .ZN(n5165) );
  OAI211_X1 U6323 ( .C1(n5189), .C2(n6718), .A(n5166), .B(n5165), .ZN(n5188)
         );
  AOI22_X1 U6324 ( .A1(n6353), .A2(n5189), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5188), .ZN(n5167) );
  OAI21_X1 U6325 ( .B1(n6576), .B2(n6399), .A(n5167), .ZN(n5168) );
  AOI21_X1 U6326 ( .B1(n5192), .B2(n6304), .A(n5168), .ZN(n5169) );
  OAI21_X1 U6327 ( .B1(n5194), .B2(n6577), .A(n5169), .ZN(U3101) );
  AOI22_X1 U6328 ( .A1(n6336), .A2(n5189), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5188), .ZN(n5170) );
  OAI21_X1 U6329 ( .B1(n6267), .B2(n6399), .A(n5170), .ZN(n5171) );
  AOI21_X1 U6330 ( .B1(n6292), .B2(n5192), .A(n5171), .ZN(n5172) );
  OAI21_X1 U6331 ( .B1(n5194), .B2(n6303), .A(n5172), .ZN(U3100) );
  AOI22_X1 U6332 ( .A1(n6391), .A2(n5189), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5188), .ZN(n5173) );
  OAI21_X1 U6333 ( .B1(n6288), .B2(n6399), .A(n5173), .ZN(n5174) );
  AOI21_X1 U6334 ( .B1(n5192), .B2(n6330), .A(n5174), .ZN(n5175) );
  OAI21_X1 U6335 ( .B1(n5194), .B2(n6334), .A(n5175), .ZN(U3107) );
  AOI22_X1 U6336 ( .A1(n6370), .A2(n5189), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5188), .ZN(n5176) );
  OAI21_X1 U6337 ( .B1(n6375), .B2(n6399), .A(n5176), .ZN(n5177) );
  AOI21_X1 U6338 ( .B1(n5192), .B2(n6371), .A(n5177), .ZN(n5178) );
  OAI21_X1 U6339 ( .B1(n5194), .B2(n6318), .A(n5178), .ZN(U3104) );
  AOI22_X1 U6340 ( .A1(n6358), .A2(n5189), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5188), .ZN(n5179) );
  OAI21_X1 U6341 ( .B1(n6363), .B2(n6399), .A(n5179), .ZN(n5180) );
  AOI21_X1 U6342 ( .B1(n5192), .B2(n6359), .A(n5180), .ZN(n5181) );
  OAI21_X1 U6343 ( .B1(n5194), .B2(n6310), .A(n5181), .ZN(U3102) );
  AOI22_X1 U6344 ( .A1(n6382), .A2(n5189), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5188), .ZN(n5182) );
  OAI21_X1 U6345 ( .B1(n6389), .B2(n6399), .A(n5182), .ZN(n5183) );
  AOI21_X1 U6346 ( .B1(n5192), .B2(n6383), .A(n5183), .ZN(n5184) );
  OAI21_X1 U6347 ( .B1(n5194), .B2(n6326), .A(n5184), .ZN(U3106) );
  AOI22_X1 U6348 ( .A1(n6376), .A2(n5189), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5188), .ZN(n5185) );
  OAI21_X1 U6349 ( .B1(n6278), .B2(n6399), .A(n5185), .ZN(n5186) );
  AOI21_X1 U6350 ( .B1(n5192), .B2(n6319), .A(n5186), .ZN(n5187) );
  OAI21_X1 U6351 ( .B1(n5194), .B2(n6322), .A(n5187), .ZN(U3105) );
  AOI22_X1 U6352 ( .A1(n6364), .A2(n5189), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5188), .ZN(n5190) );
  OAI21_X1 U6353 ( .B1(n6369), .B2(n6399), .A(n5190), .ZN(n5191) );
  AOI21_X1 U6354 ( .B1(n5192), .B2(n6365), .A(n5191), .ZN(n5193) );
  OAI21_X1 U6355 ( .B1(n5194), .B2(n6314), .A(n5193), .ZN(U3103) );
  INV_X1 U6356 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5196) );
  OAI222_X1 U6357 ( .A1(n5197), .A2(n5817), .B1(n6045), .B2(n5196), .C1(n5195), 
        .C2(n5819), .ZN(U2849) );
  NAND2_X1 U6358 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  XNOR2_X1 U6359 ( .A(n5199), .B(n5202), .ZN(n6205) );
  NAND2_X1 U6360 ( .A1(n6205), .A2(n6185), .ZN(n5206) );
  AND2_X1 U6361 ( .A1(n6238), .A2(REIP_REG_11__SCAN_IN), .ZN(n6202) );
  NOR2_X1 U6362 ( .A1(n6191), .A2(n5203), .ZN(n5204) );
  AOI211_X1 U6363 ( .C1(n6197), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6202), 
        .B(n5204), .ZN(n5205) );
  OAI211_X1 U6364 ( .C1(n6200), .C2(n5207), .A(n5206), .B(n5205), .ZN(U2975)
         );
  INV_X1 U6365 ( .A(n5237), .ZN(n5210) );
  NOR2_X1 U6366 ( .A1(n5236), .A2(n5210), .ZN(n5211) );
  XNOR2_X1 U6367 ( .A(n5209), .B(n5211), .ZN(n5235) );
  INV_X1 U6368 ( .A(n5212), .ZN(n5213) );
  OAI22_X1 U6369 ( .A1(n5214), .A2(n5219), .B1(n5213), .B2(n5216), .ZN(n6204)
         );
  INV_X1 U6370 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6705) );
  NAND3_X1 U6371 ( .A1(n5215), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n5219), 
        .ZN(n5218) );
  INV_X1 U6372 ( .A(n5216), .ZN(n5217) );
  NAND2_X1 U6373 ( .A1(n5218), .A2(n5217), .ZN(n5260) );
  AOI21_X1 U6374 ( .B1(n5220), .B2(n5219), .A(n5260), .ZN(n6208) );
  INV_X1 U6375 ( .A(n6208), .ZN(n5264) );
  OAI211_X1 U6376 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5264), .B(n5249), .ZN(n5224) );
  INV_X1 U6377 ( .A(n5221), .ZN(n5222) );
  AOI21_X1 U6378 ( .B1(n5222), .B2(n3561), .A(n5250), .ZN(n5973) );
  NAND2_X1 U6379 ( .A1(n5973), .A2(n6240), .ZN(n5223) );
  OAI211_X1 U6380 ( .C1(n6705), .C2(n6192), .A(n5224), .B(n5223), .ZN(n5225)
         );
  AOI21_X1 U6381 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6204), .A(n5225), 
        .ZN(n5226) );
  OAI21_X1 U6382 ( .B1(n5235), .B2(n5717), .A(n5226), .ZN(U3006) );
  AOI21_X1 U6383 ( .B1(n5227), .B2(n5134), .A(n5302), .ZN(n5977) );
  INV_X1 U6384 ( .A(n5977), .ZN(n5230) );
  AOI22_X1 U6385 ( .A1(n5973), .A2(n6040), .B1(EBX_REG_12__SCAN_IN), .B2(n5501), .ZN(n5228) );
  OAI21_X1 U6386 ( .B1(n5230), .B2(n5819), .A(n5228), .ZN(U2847) );
  AOI22_X1 U6387 ( .A1(n5514), .A2(DATAI_12_), .B1(n6061), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5229) );
  OAI21_X1 U6388 ( .B1(n5230), .B2(n6047), .A(n5229), .ZN(U2879) );
  AOI22_X1 U6389 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6238), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5231) );
  OAI21_X1 U6390 ( .B1(n6191), .B2(n5232), .A(n5231), .ZN(n5233) );
  AOI21_X1 U6391 ( .B1(n5977), .B2(n6186), .A(n5233), .ZN(n5234) );
  OAI21_X1 U6392 ( .B1(n5235), .B2(n6193), .A(n5234), .ZN(U2974) );
  OR2_X1 U6393 ( .A1(n5209), .A2(n5236), .ZN(n5238) );
  NAND2_X1 U6394 ( .A1(n5238), .A2(n5237), .ZN(n5243) );
  OR2_X1 U6395 ( .A1(n5209), .A2(n5239), .ZN(n5257) );
  AND2_X1 U6396 ( .A1(n5257), .A2(n5240), .ZN(n5241) );
  OAI21_X1 U6397 ( .B1(n5243), .B2(n5242), .A(n5241), .ZN(n5244) );
  INV_X1 U6398 ( .A(n5244), .ZN(n5280) );
  INV_X1 U6399 ( .A(n5245), .ZN(n5246) );
  AOI21_X1 U6400 ( .B1(n5249), .B2(n5246), .A(n6204), .ZN(n5247) );
  OAI21_X1 U6401 ( .B1(n5263), .B2(n5248), .A(n5247), .ZN(n5262) );
  NOR2_X1 U6402 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5249), .ZN(n5261)
         );
  AOI22_X1 U6403 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5262), .B1(n5261), .B2(n5264), .ZN(n5255) );
  INV_X1 U6404 ( .A(n5250), .ZN(n5252) );
  INV_X1 U6405 ( .A(n5267), .ZN(n5251) );
  AOI21_X1 U6406 ( .B1(n5253), .B2(n5252), .A(n5251), .ZN(n5288) );
  NOR2_X1 U6407 ( .A1(n6192), .A2(n6492), .ZN(n5275) );
  AOI21_X1 U6408 ( .B1(n5288), .B2(n6240), .A(n5275), .ZN(n5254) );
  OAI211_X1 U6409 ( .C1(n5280), .C2(n5717), .A(n5255), .B(n5254), .ZN(U3005)
         );
  NAND2_X1 U6410 ( .A1(n5257), .A2(n5256), .ZN(n5259) );
  XNOR2_X1 U6411 ( .A(n5708), .B(n5265), .ZN(n5258) );
  XNOR2_X1 U6412 ( .A(n5259), .B(n5258), .ZN(n5351) );
  OAI221_X1 U6413 ( .B1(n5262), .B2(n5261), .C1(n5262), .C2(n5260), .A(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5272) );
  AND3_X1 U6414 ( .A1(n5265), .A2(n5264), .A3(n5263), .ZN(n5270) );
  NAND2_X1 U6415 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  NAND2_X1 U6416 ( .A1(n5438), .A2(n5268), .ZN(n5971) );
  INV_X1 U6417 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6494) );
  OAI22_X1 U6418 ( .A1(n5971), .A2(n3628), .B1(n6494), .B2(n6192), .ZN(n5269)
         );
  NOR2_X1 U6419 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  OAI211_X1 U6420 ( .C1(n5351), .C2(n5717), .A(n5272), .B(n5271), .ZN(U3004)
         );
  XOR2_X1 U6421 ( .A(n5299), .B(n5300), .Z(n5278) );
  AOI22_X1 U6422 ( .A1(n5288), .A2(n6040), .B1(EBX_REG_13__SCAN_IN), .B2(n5501), .ZN(n5274) );
  OAI21_X1 U6423 ( .B1(n5327), .B2(n5819), .A(n5274), .ZN(U2846) );
  AOI21_X1 U6424 ( .B1(n6197), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5275), 
        .ZN(n5276) );
  OAI21_X1 U6425 ( .B1(n5286), .B2(n6191), .A(n5276), .ZN(n5277) );
  AOI21_X1 U6426 ( .B1(n5278), .B2(n6186), .A(n5277), .ZN(n5279) );
  OAI21_X1 U6427 ( .B1(n5280), .B2(n6193), .A(n5279), .ZN(U2973) );
  INV_X1 U6428 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6492) );
  AOI211_X1 U6429 ( .C1(n6705), .C2(n6492), .A(n5974), .B(n6026), .ZN(n5282)
         );
  AOI22_X1 U6430 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6028), .B1(n5282), .B2(n5281), .ZN(n5283) );
  OAI211_X1 U6431 ( .C1(n6018), .C2(n5284), .A(n5283), .B(n5994), .ZN(n5285)
         );
  AOI21_X1 U6432 ( .B1(REIP_REG_13__SCAN_IN), .B2(n5972), .A(n5285), .ZN(n5290) );
  INV_X1 U6433 ( .A(n5286), .ZN(n5287) );
  AOI22_X1 U6434 ( .A1(n5288), .A2(n6007), .B1(n5999), .B2(n5287), .ZN(n5289)
         );
  OAI211_X1 U6435 ( .C1(n5327), .C2(n5955), .A(n5290), .B(n5289), .ZN(U2814)
         );
  OAI21_X1 U6436 ( .B1(n5293), .B2(n5292), .A(n5332), .ZN(n5586) );
  INV_X1 U6437 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5298) );
  OR2_X1 U6438 ( .A1(n5296), .A2(n5295), .ZN(n5297) );
  NAND2_X1 U6439 ( .A1(n5294), .A2(n5297), .ZN(n5790) );
  OAI222_X1 U6440 ( .A1(n5586), .A2(n5819), .B1(n5298), .B2(n6045), .C1(n5817), 
        .C2(n5790), .ZN(U2838) );
  NAND2_X1 U6441 ( .A1(n5300), .A2(n5299), .ZN(n5304) );
  NAND2_X1 U6442 ( .A1(n5302), .A2(n5301), .ZN(n5303) );
  NAND2_X1 U6443 ( .A1(n5484), .A2(n5305), .ZN(n5476) );
  NAND2_X1 U6444 ( .A1(n5484), .A2(n5306), .ZN(n5345) );
  NAND2_X1 U6445 ( .A1(n5345), .A2(n5307), .ZN(n5308) );
  NAND2_X1 U6446 ( .A1(n5476), .A2(n5308), .ZN(n5806) );
  MUX2_X1 U6447 ( .A(n5479), .B(n5309), .S(n5399), .Z(n5338) );
  OR2_X1 U6448 ( .A1(n5339), .A2(n5338), .ZN(n5341) );
  INV_X1 U6449 ( .A(n5310), .ZN(n5311) );
  XNOR2_X1 U6450 ( .A(n5341), .B(n5311), .ZN(n5807) );
  NOR2_X1 U6451 ( .A1(n6045), .A2(n5312), .ZN(n5313) );
  AOI21_X1 U6452 ( .B1(n5807), .B2(n6040), .A(n5313), .ZN(n5314) );
  OAI21_X1 U6453 ( .B1(n5806), .B2(n5819), .A(n5314), .ZN(U2840) );
  NAND2_X1 U6454 ( .A1(n4227), .A2(n6708), .ZN(n5318) );
  NAND3_X1 U6455 ( .A1(n5316), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5576), .ZN(n5317) );
  OAI21_X1 U6456 ( .B1(n5316), .B2(n5318), .A(n5317), .ZN(n5319) );
  XNOR2_X1 U6457 ( .A(n5319), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5867)
         );
  INV_X1 U6458 ( .A(n5702), .ZN(n5325) );
  OR2_X1 U6459 ( .A1(n5496), .A2(n5320), .ZN(n5321) );
  NAND2_X1 U6460 ( .A1(n5339), .A2(n5321), .ZN(n5943) );
  NAND2_X1 U6461 ( .A1(n6238), .A2(REIP_REG_17__SCAN_IN), .ZN(n5871) );
  OAI21_X1 U6462 ( .B1(n5943), .B2(n3628), .A(n5871), .ZN(n5324) );
  INV_X1 U6463 ( .A(n5322), .ZN(n5720) );
  NOR2_X1 U6464 ( .A1(n5720), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5323)
         );
  AOI211_X1 U6465 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5325), .A(n5324), .B(n5323), .ZN(n5326) );
  OAI21_X1 U6466 ( .B1(n5867), .B2(n5717), .A(n5326), .ZN(U3001) );
  INV_X1 U6467 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6173) );
  INV_X1 U6468 ( .A(DATAI_13_), .ZN(n5328) );
  OAI222_X1 U6469 ( .A1(n5505), .A2(n6173), .B1(n5329), .B2(n5328), .C1(n6047), 
        .C2(n5327), .ZN(U2878) );
  NAND2_X1 U6470 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  NAND2_X1 U6471 ( .A1(n5330), .A2(n5333), .ZN(n5840) );
  NAND2_X1 U6472 ( .A1(n5294), .A2(n5334), .ZN(n5335) );
  NAND2_X1 U6473 ( .A1(n5427), .A2(n5335), .ZN(n5785) );
  OAI22_X1 U6474 ( .A1(n5785), .A2(n5817), .B1(n6721), .B2(n6045), .ZN(n5336)
         );
  INV_X1 U6475 ( .A(n5336), .ZN(n5337) );
  OAI21_X1 U6476 ( .B1(n5840), .B2(n5819), .A(n5337), .ZN(U2837) );
  NAND2_X1 U6477 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  NAND2_X1 U6478 ( .A1(n5341), .A2(n5340), .ZN(n5937) );
  NAND2_X1 U6479 ( .A1(n5484), .A2(n5342), .ZN(n5489) );
  NAND2_X1 U6480 ( .A1(n5489), .A2(n5343), .ZN(n5344) );
  NAND2_X1 U6481 ( .A1(n5345), .A2(n5344), .ZN(n6048) );
  OAI222_X1 U6482 ( .A1(n5937), .A2(n5817), .B1(n6045), .B2(n3585), .C1(n6048), 
        .C2(n5819), .ZN(U2841) );
  NAND2_X1 U6483 ( .A1(n5484), .A2(n5483), .ZN(n5436) );
  OR2_X1 U6484 ( .A1(n5484), .A2(n5483), .ZN(n5346) );
  INV_X1 U6485 ( .A(n5968), .ZN(n5352) );
  AOI22_X1 U6486 ( .A1(n5514), .A2(DATAI_14_), .B1(n6061), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5347) );
  OAI21_X1 U6487 ( .B1(n5352), .B2(n6047), .A(n5347), .ZN(U2877) );
  AOI22_X1 U6488 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6238), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5348) );
  OAI21_X1 U6489 ( .B1(n5966), .B2(n6191), .A(n5348), .ZN(n5349) );
  AOI21_X1 U6490 ( .B1(n5968), .B2(n6186), .A(n5349), .ZN(n5350) );
  OAI21_X1 U6491 ( .B1(n5351), .B2(n6193), .A(n5350), .ZN(U2972) );
  INV_X1 U6492 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5353) );
  OAI222_X1 U6493 ( .A1(n5971), .A2(n5817), .B1(n6045), .B2(n5353), .C1(n5352), 
        .C2(n5819), .ZN(U2845) );
  OAI22_X1 U6494 ( .A1(n5355), .A2(n5817), .B1(n6045), .B2(n5354), .ZN(U2828)
         );
  AOI22_X1 U6495 ( .A1(n6040), .A2(n5356), .B1(n5501), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5357) );
  OAI21_X1 U6496 ( .B1(n5366), .B2(n5819), .A(n5357), .ZN(U2858) );
  AOI22_X1 U6497 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6028), .B1(n5441), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n5365) );
  INV_X1 U6498 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5358) );
  AOI22_X1 U6499 ( .A1(n5993), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5999), 
        .B2(n5358), .ZN(n5361) );
  NAND2_X1 U6500 ( .A1(n6023), .A2(n5359), .ZN(n5360) );
  OAI211_X1 U6501 ( .C1(REIP_REG_1__SCAN_IN), .C2(n6026), .A(n5361), .B(n5360), 
        .ZN(n5362) );
  AOI21_X1 U6502 ( .B1(n6007), .B2(n5363), .A(n5362), .ZN(n5364) );
  OAI211_X1 U6503 ( .C1(n5367), .C2(n5366), .A(n5365), .B(n5364), .ZN(U2826)
         );
  XOR2_X1 U6504 ( .A(n5369), .B(n5368), .Z(n6233) );
  NAND2_X1 U6505 ( .A1(n6233), .A2(n6185), .ZN(n5374) );
  NAND2_X1 U6506 ( .A1(n6238), .A2(REIP_REG_3__SCAN_IN), .ZN(n6229) );
  INV_X1 U6507 ( .A(n6229), .ZN(n5372) );
  NOR2_X1 U6508 ( .A1(n6191), .A2(n5370), .ZN(n5371) );
  AOI211_X1 U6509 ( .C1(n6197), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5372), 
        .B(n5371), .ZN(n5373) );
  OAI211_X1 U6510 ( .C1(n6200), .C2(n5375), .A(n5374), .B(n5373), .ZN(U2983)
         );
  NAND3_X1 U6511 ( .A1(n5377), .A2(n5376), .A3(n5505), .ZN(n5380) );
  AOI22_X1 U6512 ( .A1(n6052), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6061), .ZN(n5379) );
  NAND2_X1 U6513 ( .A1(n5380), .A2(n5379), .ZN(U2860) );
  NOR3_X1 U6514 ( .A1(n6441), .A2(n5382), .A3(n5381), .ZN(n5385) );
  INV_X1 U6515 ( .A(n5387), .ZN(n5383) );
  NOR3_X1 U6516 ( .A1(n5388), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5383), 
        .ZN(n5384) );
  AOI211_X1 U6517 ( .C1(n5386), .C2(n5902), .A(n5385), .B(n5384), .ZN(n5392)
         );
  AOI21_X1 U6518 ( .B1(n5388), .B2(n5387), .A(n5391), .ZN(n5390) );
  OAI22_X1 U6519 ( .A1(n5392), .A2(n5391), .B1(n5390), .B2(n5389), .ZN(U3459)
         );
  XNOR2_X1 U6520 ( .A(n5412), .B(n5394), .ZN(n5524) );
  INV_X1 U6521 ( .A(n5524), .ZN(n5508) );
  INV_X1 U6522 ( .A(n5401), .ZN(n5397) );
  INV_X1 U6523 ( .A(n5454), .ZN(n5395) );
  NAND2_X1 U6524 ( .A1(n5402), .A2(n5395), .ZN(n5396) );
  NAND3_X1 U6525 ( .A1(n5398), .A2(n5397), .A3(n5396), .ZN(n5404) );
  NAND2_X1 U6526 ( .A1(n5454), .A2(n5399), .ZN(n5400) );
  NAND3_X1 U6527 ( .A1(n5402), .A2(n5401), .A3(n5400), .ZN(n5403) );
  NOR3_X1 U6528 ( .A1(n5419), .A2(REIP_REG_30__SCAN_IN), .A3(n6520), .ZN(n5409) );
  AOI22_X1 U6529 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5993), .B1(n5999), 
        .B2(n5520), .ZN(n5406) );
  NAND2_X1 U6530 ( .A1(n6028), .A2(EBX_REG_30__SCAN_IN), .ZN(n5405) );
  OAI211_X1 U6531 ( .C1(n5407), .C2(n6522), .A(n5406), .B(n5405), .ZN(n5408)
         );
  AOI211_X1 U6532 ( .C1(n5628), .C2(n6007), .A(n5409), .B(n5408), .ZN(n5410)
         );
  OAI21_X1 U6533 ( .B1(n5508), .B2(n5955), .A(n5410), .ZN(U2797) );
  AOI21_X1 U6534 ( .B1(n5413), .B2(n5411), .A(n5412), .ZN(n5533) );
  INV_X1 U6535 ( .A(n5533), .ZN(n5511) );
  XNOR2_X1 U6536 ( .A(n5454), .B(n5414), .ZN(n5637) );
  OAI22_X1 U6537 ( .A1(n5530), .A2(n6018), .B1(n6037), .B2(n5529), .ZN(n5417)
         );
  INV_X1 U6538 ( .A(n5415), .ZN(n5735) );
  NOR2_X1 U6539 ( .A1(n5735), .A2(n6520), .ZN(n5416) );
  AOI211_X1 U6540 ( .C1(EBX_REG_29__SCAN_IN), .C2(n6028), .A(n5417), .B(n5416), 
        .ZN(n5418) );
  OAI21_X1 U6541 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5419), .A(n5418), .ZN(n5420) );
  AOI21_X1 U6542 ( .B1(n6007), .B2(n5637), .A(n5420), .ZN(n5421) );
  OAI21_X1 U6543 ( .B1(n5511), .B2(n5955), .A(n5421), .ZN(U2798) );
  AOI21_X1 U6544 ( .B1(n5424), .B2(n5330), .A(n5423), .ZN(n5836) );
  INV_X1 U6545 ( .A(n5836), .ZN(n5474) );
  INV_X1 U6546 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U6547 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5776), .ZN(n5777) );
  INV_X1 U6548 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6648) );
  OAI21_X1 U6549 ( .B1(n6507), .B2(n5777), .A(n6648), .ZN(n5433) );
  NOR2_X1 U6550 ( .A1(n5811), .A2(n5425), .ZN(n5768) );
  NAND2_X1 U6551 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  NAND2_X1 U6552 ( .A1(n5429), .A2(n5428), .ZN(n5671) );
  INV_X1 U6553 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5473) );
  OAI22_X1 U6554 ( .A1(n5671), .A2(n6031), .B1(n6004), .B2(n5473), .ZN(n5432)
         );
  INV_X1 U6555 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5430) );
  OAI22_X1 U6556 ( .A1(n5430), .A2(n6018), .B1(n5572), .B2(n6037), .ZN(n5431)
         );
  AOI211_X1 U6557 ( .C1(n5433), .C2(n5768), .A(n5432), .B(n5431), .ZN(n5434)
         );
  OAI21_X1 U6558 ( .B1(n5474), .B2(n5955), .A(n5434), .ZN(U2804) );
  INV_X1 U6559 ( .A(n5493), .ZN(n5435) );
  AOI21_X1 U6560 ( .B1(n5437), .B2(n5436), .A(n5435), .ZN(n5622) );
  INV_X1 U6561 ( .A(n5622), .ZN(n5516) );
  AOI21_X1 U6562 ( .B1(n5439), .B2(n5438), .A(n5499), .ZN(n5894) );
  AOI21_X1 U6563 ( .B1(n5993), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6022), 
        .ZN(n5440) );
  OAI21_X1 U6564 ( .B1(n6037), .B2(n5620), .A(n5440), .ZN(n5444) );
  AOI21_X1 U6565 ( .B1(n6009), .B2(n5960), .A(n5441), .ZN(n5964) );
  INV_X1 U6566 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6497) );
  AOI22_X1 U6567 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6028), .B1(n5950), .B2(n6497), .ZN(n5442) );
  OAI21_X1 U6568 ( .B1(n5964), .B2(n6497), .A(n5442), .ZN(n5443) );
  AOI211_X1 U6569 ( .C1(n5894), .C2(n6007), .A(n5444), .B(n5443), .ZN(n5445)
         );
  OAI21_X1 U6570 ( .B1(n5516), .B2(n5955), .A(n5445), .ZN(U2812) );
  AOI22_X1 U6571 ( .A1(n5628), .A2(n6040), .B1(EBX_REG_30__SCAN_IN), .B2(n5501), .ZN(n5446) );
  OAI21_X1 U6572 ( .B1(n5508), .B2(n5819), .A(n5446), .ZN(U2829) );
  AOI22_X1 U6573 ( .A1(n5637), .A2(n6040), .B1(EBX_REG_29__SCAN_IN), .B2(n5501), .ZN(n5447) );
  OAI21_X1 U6574 ( .B1(n5511), .B2(n5819), .A(n5447), .ZN(U2830) );
  OR2_X1 U6575 ( .A1(n5448), .A2(n5449), .ZN(n5450) );
  OR2_X1 U6576 ( .A1(n5451), .A2(n5452), .ZN(n5453) );
  NAND2_X1 U6577 ( .A1(n5454), .A2(n5453), .ZN(n5741) );
  OAI22_X1 U6578 ( .A1(n5741), .A2(n5817), .B1(n5734), .B2(n6045), .ZN(n5455)
         );
  AOI21_X1 U6579 ( .B1(n5823), .B2(n6041), .A(n5455), .ZN(n5456) );
  INV_X1 U6580 ( .A(n5456), .ZN(U2831) );
  AOI21_X1 U6581 ( .B1(n5460), .B2(n5459), .A(n5458), .ZN(n5559) );
  INV_X1 U6582 ( .A(n5559), .ZN(n5751) );
  INV_X1 U6583 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5463) );
  OR2_X1 U6584 ( .A1(n5467), .A2(n5461), .ZN(n5462) );
  NAND2_X1 U6585 ( .A1(n5648), .A2(n5462), .ZN(n5750) );
  OAI222_X1 U6586 ( .A1(n5819), .A2(n5751), .B1(n6045), .B2(n5463), .C1(n5750), 
        .C2(n5817), .ZN(U2833) );
  AOI21_X1 U6587 ( .B1(n5466), .B2(n5464), .A(n5465), .ZN(n5857) );
  INV_X1 U6588 ( .A(n5857), .ZN(n5760) );
  INV_X1 U6589 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5471) );
  INV_X1 U6590 ( .A(n5467), .ZN(n5468) );
  OAI21_X1 U6591 ( .B1(n5470), .B2(n5469), .A(n5468), .ZN(n5876) );
  OAI222_X1 U6592 ( .A1(n5760), .A2(n5819), .B1(n5471), .B2(n6045), .C1(n5817), 
        .C2(n5876), .ZN(U2834) );
  OAI21_X1 U6593 ( .B1(n5423), .B2(n5472), .A(n5464), .ZN(n5769) );
  INV_X1 U6594 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6671) );
  OAI222_X1 U6595 ( .A1(n5819), .A2(n5769), .B1(n6045), .B2(n6671), .C1(n5773), 
        .C2(n5817), .ZN(U2835) );
  OAI222_X1 U6596 ( .A1(n5819), .A2(n5474), .B1(n5473), .B2(n6045), .C1(n5671), 
        .C2(n5817), .ZN(U2836) );
  XNOR2_X1 U6597 ( .A(n5476), .B(n5475), .ZN(n5848) );
  INV_X1 U6598 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5482) );
  MUX2_X1 U6599 ( .A(n5479), .B(n5478), .S(n5477), .Z(n5480) );
  XOR2_X1 U6600 ( .A(n5481), .B(n5480), .Z(n5805) );
  OAI222_X1 U6601 ( .A1(n5848), .A2(n5819), .B1(n5482), .B2(n6045), .C1(n5817), 
        .C2(n5805), .ZN(U2839) );
  AND2_X1 U6602 ( .A1(n5484), .A2(n5483), .ZN(n5486) );
  INV_X1 U6603 ( .A(n6054), .ZN(n5491) );
  INV_X1 U6604 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5490) );
  OAI222_X1 U6605 ( .A1(n5491), .A2(n5819), .B1(n5490), .B2(n6045), .C1(n5817), 
        .C2(n5943), .ZN(U2842) );
  AND2_X1 U6606 ( .A1(n5493), .A2(n5492), .ZN(n5495) );
  INV_X1 U6607 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5500) );
  INV_X1 U6608 ( .A(n5496), .ZN(n5497) );
  OAI21_X1 U6609 ( .B1(n5499), .B2(n5498), .A(n5497), .ZN(n5959) );
  OAI222_X1 U6610 ( .A1(n6059), .A2(n5819), .B1(n6045), .B2(n5500), .C1(n5959), 
        .C2(n5817), .ZN(U2843) );
  AOI22_X1 U6611 ( .A1(n5894), .A2(n6040), .B1(EBX_REG_15__SCAN_IN), .B2(n5501), .ZN(n5502) );
  OAI21_X1 U6612 ( .B1(n5516), .B2(n5819), .A(n5502), .ZN(U2844) );
  AOI22_X1 U6613 ( .A1(n6052), .A2(DATAI_30_), .B1(n6061), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5507) );
  AND2_X1 U6614 ( .A1(n3190), .A2(n5503), .ZN(n5504) );
  NAND2_X1 U6615 ( .A1(n6062), .A2(DATAI_14_), .ZN(n5506) );
  OAI211_X1 U6616 ( .C1(n5508), .C2(n6047), .A(n5507), .B(n5506), .ZN(U2861)
         );
  AOI22_X1 U6617 ( .A1(n6052), .A2(DATAI_29_), .B1(n6061), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U6618 ( .A1(n6062), .A2(DATAI_13_), .ZN(n5509) );
  OAI211_X1 U6619 ( .C1(n5511), .C2(n6047), .A(n5510), .B(n5509), .ZN(U2862)
         );
  AOI22_X1 U6620 ( .A1(n6062), .A2(DATAI_10_), .B1(n6061), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U6621 ( .A1(n6052), .A2(DATAI_26_), .ZN(n5512) );
  OAI211_X1 U6622 ( .C1(n5751), .C2(n6047), .A(n5513), .B(n5512), .ZN(U2865)
         );
  AOI22_X1 U6623 ( .A1(n5514), .A2(DATAI_15_), .B1(n6061), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5515) );
  OAI21_X1 U6624 ( .B1(n5516), .B2(n6047), .A(n5515), .ZN(U2876) );
  NOR2_X1 U6625 ( .A1(n5555), .A2(n5518), .ZN(n5526) );
  XNOR2_X1 U6626 ( .A(n5519), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5630)
         );
  NAND2_X1 U6627 ( .A1(n5868), .A2(n5520), .ZN(n5521) );
  NAND2_X1 U6628 ( .A1(n6238), .A2(REIP_REG_30__SCAN_IN), .ZN(n5624) );
  OAI211_X1 U6629 ( .C1(n5522), .C2(n5873), .A(n5521), .B(n5624), .ZN(n5523)
         );
  AOI21_X1 U6630 ( .B1(n5524), .B2(n6186), .A(n5523), .ZN(n5525) );
  OAI21_X1 U6631 ( .B1(n5630), .B2(n6193), .A(n5525), .ZN(U2956) );
  NOR2_X1 U6632 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  NOR2_X1 U6633 ( .A1(n6191), .A2(n5529), .ZN(n5532) );
  NAND2_X1 U6634 ( .A1(n5592), .A2(REIP_REG_29__SCAN_IN), .ZN(n5633) );
  OAI21_X1 U6635 ( .B1(n5873), .B2(n5530), .A(n5633), .ZN(n5531) );
  AOI211_X1 U6636 ( .C1(n5533), .C2(n6186), .A(n5532), .B(n5531), .ZN(n5534)
         );
  OAI21_X1 U6637 ( .B1(n3002), .B2(n6193), .A(n5534), .ZN(U2957) );
  AND3_X1 U6638 ( .A1(n5555), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5576), 
        .ZN(n5537) );
  NAND2_X1 U6639 ( .A1(n5553), .A2(n6612), .ZN(n5535) );
  NOR2_X1 U6640 ( .A1(n5536), .A2(n5535), .ZN(n5543) );
  OAI22_X1 U6641 ( .A1(n5537), .A2(n5543), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5650), .ZN(n5538) );
  XNOR2_X1 U6642 ( .A(n5538), .B(n5640), .ZN(n5646) );
  NAND2_X1 U6643 ( .A1(n5868), .A2(n5738), .ZN(n5539) );
  NAND2_X1 U6644 ( .A1(n5592), .A2(REIP_REG_28__SCAN_IN), .ZN(n5643) );
  OAI211_X1 U6645 ( .C1(n5873), .C2(n5540), .A(n5539), .B(n5643), .ZN(n5541)
         );
  AOI21_X1 U6646 ( .B1(n5823), .B2(n6186), .A(n5541), .ZN(n5542) );
  OAI21_X1 U6647 ( .B1(n6193), .B2(n5646), .A(n5542), .ZN(U2958) );
  INV_X1 U6648 ( .A(n5543), .ZN(n5544) );
  NAND2_X1 U6649 ( .A1(n5545), .A2(n5544), .ZN(n5546) );
  XNOR2_X1 U6650 ( .A(n5546), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5657)
         );
  NOR2_X1 U6651 ( .A1(n5458), .A2(n5547), .ZN(n5548) );
  OR2_X1 U6652 ( .A1(n5448), .A2(n5548), .ZN(n5827) );
  INV_X1 U6653 ( .A(n5827), .ZN(n5551) );
  NAND2_X1 U6654 ( .A1(n5592), .A2(REIP_REG_27__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U6655 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5549)
         );
  OAI211_X1 U6656 ( .C1(n6191), .C2(n5747), .A(n5653), .B(n5549), .ZN(n5550)
         );
  AOI21_X1 U6657 ( .B1(n5551), .B2(n6186), .A(n5550), .ZN(n5552) );
  OAI21_X1 U6658 ( .B1(n5657), .B2(n6193), .A(n5552), .ZN(U2959) );
  NOR2_X1 U6659 ( .A1(n5554), .A2(n5553), .ZN(n5556) );
  XOR2_X1 U6660 ( .A(n5556), .B(n5555), .Z(n5666) );
  NAND2_X1 U6661 ( .A1(n5868), .A2(n5748), .ZN(n5557) );
  NAND2_X1 U6662 ( .A1(n5592), .A2(REIP_REG_26__SCAN_IN), .ZN(n5663) );
  OAI211_X1 U6663 ( .C1(n5873), .C2(n5757), .A(n5557), .B(n5663), .ZN(n5558)
         );
  AOI21_X1 U6664 ( .B1(n5559), .B2(n6186), .A(n5558), .ZN(n5560) );
  OAI21_X1 U6665 ( .B1(n5666), .B2(n6193), .A(n5560), .ZN(U2960) );
  OAI21_X1 U6666 ( .B1(n5873), .B2(n5562), .A(n5561), .ZN(n5564) );
  NOR2_X1 U6667 ( .A1(n5769), .A2(n6200), .ZN(n5563) );
  AOI211_X1 U6668 ( .C1(n5868), .C2(n5770), .A(n5564), .B(n5563), .ZN(n5565)
         );
  OAI21_X1 U6669 ( .B1(n5566), .B2(n6193), .A(n5565), .ZN(U2962) );
  NAND3_X1 U6670 ( .A1(n5576), .A2(n5694), .A3(n5679), .ZN(n5568) );
  OAI21_X1 U6671 ( .B1(n5569), .B2(n5568), .A(n5567), .ZN(n5570) );
  XNOR2_X1 U6672 ( .A(n5570), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5675)
         );
  NAND2_X1 U6673 ( .A1(n5592), .A2(REIP_REG_23__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U6674 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5571)
         );
  OAI211_X1 U6675 ( .C1(n6191), .C2(n5572), .A(n5670), .B(n5571), .ZN(n5573)
         );
  AOI21_X1 U6676 ( .B1(n5836), .B2(n6186), .A(n5573), .ZN(n5574) );
  OAI21_X1 U6677 ( .B1(n5675), .B2(n6193), .A(n5574), .ZN(U2963) );
  AOI21_X1 U6678 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5576), .A(n5575), 
        .ZN(n5577) );
  XNOR2_X1 U6679 ( .A(n5578), .B(n5577), .ZN(n5684) );
  NAND2_X1 U6680 ( .A1(n5592), .A2(REIP_REG_22__SCAN_IN), .ZN(n5677) );
  OAI21_X1 U6681 ( .B1(n5873), .B2(n5579), .A(n5677), .ZN(n5581) );
  NOR2_X1 U6682 ( .A1(n5840), .A2(n6200), .ZN(n5580) );
  AOI211_X1 U6683 ( .C1(n5868), .C2(n5780), .A(n5581), .B(n5580), .ZN(n5582)
         );
  OAI21_X1 U6684 ( .B1(n5684), .B2(n6193), .A(n5582), .ZN(U2964) );
  AOI21_X1 U6685 ( .B1(n5585), .B2(n5584), .A(n5583), .ZN(n5691) );
  INV_X1 U6686 ( .A(n5586), .ZN(n5844) );
  NAND2_X1 U6687 ( .A1(n5592), .A2(REIP_REG_21__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U6688 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5587)
         );
  OAI211_X1 U6689 ( .C1(n6191), .C2(n5794), .A(n5685), .B(n5587), .ZN(n5588)
         );
  AOI21_X1 U6690 ( .B1(n5844), .B2(n6186), .A(n5588), .ZN(n5589) );
  OAI21_X1 U6691 ( .B1(n5691), .B2(n6193), .A(n5589), .ZN(U2965) );
  XOR2_X1 U6692 ( .A(n5591), .B(n5590), .Z(n5707) );
  NAND2_X1 U6693 ( .A1(n5592), .A2(REIP_REG_20__SCAN_IN), .ZN(n5692) );
  OAI21_X1 U6694 ( .B1(n5873), .B2(n5796), .A(n5692), .ZN(n5594) );
  NOR2_X1 U6695 ( .A1(n5848), .A2(n6200), .ZN(n5593) );
  AOI211_X1 U6696 ( .C1(n5868), .C2(n5800), .A(n5594), .B(n5593), .ZN(n5595)
         );
  OAI21_X1 U6697 ( .B1(n5707), .B2(n6193), .A(n5595), .ZN(U2966) );
  INV_X1 U6698 ( .A(n5596), .ZN(n5597) );
  NOR2_X1 U6699 ( .A1(n5316), .A2(n5597), .ZN(n5600) );
  INV_X1 U6700 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5719) );
  NOR2_X1 U6701 ( .A1(n5598), .A2(n5719), .ZN(n5599) );
  MUX2_X1 U6702 ( .A(n5600), .B(n5599), .S(n5708), .Z(n5601) );
  XNOR2_X1 U6703 ( .A(n5601), .B(n5726), .ZN(n5718) );
  NAND2_X1 U6704 ( .A1(n5718), .A2(n6185), .ZN(n5606) );
  INV_X1 U6705 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5602) );
  NOR2_X1 U6706 ( .A1(n6192), .A2(n5602), .ZN(n5722) );
  INV_X1 U6707 ( .A(n5603), .ZN(n5933) );
  NOR2_X1 U6708 ( .A1(n6191), .A2(n5933), .ZN(n5604) );
  AOI211_X1 U6709 ( .C1(n6197), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5722), 
        .B(n5604), .ZN(n5605) );
  OAI211_X1 U6710 ( .C1(n6200), .C2(n6048), .A(n5606), .B(n5605), .ZN(U2968)
         );
  XNOR2_X1 U6711 ( .A(n5708), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5607)
         );
  XNOR2_X1 U6712 ( .A(n5316), .B(n5607), .ZN(n5882) );
  INV_X1 U6713 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5608) );
  OAI22_X1 U6714 ( .A1(n5873), .A2(n5609), .B1(n6192), .B2(n5608), .ZN(n5611)
         );
  NOR2_X1 U6715 ( .A1(n6059), .A2(n6200), .ZN(n5610) );
  AOI211_X1 U6716 ( .C1(n5868), .C2(n5953), .A(n5611), .B(n5610), .ZN(n5612)
         );
  OAI21_X1 U6717 ( .B1(n5882), .B2(n6193), .A(n5612), .ZN(U2970) );
  OR2_X1 U6718 ( .A1(n5209), .A2(n5613), .ZN(n5615) );
  NAND2_X1 U6719 ( .A1(n5615), .A2(n5614), .ZN(n5618) );
  NAND2_X1 U6720 ( .A1(n3008), .A2(n5616), .ZN(n5617) );
  XNOR2_X1 U6721 ( .A(n5618), .B(n5617), .ZN(n5893) );
  AOI22_X1 U6722 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6238), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5619) );
  OAI21_X1 U6723 ( .B1(n6191), .B2(n5620), .A(n5619), .ZN(n5621) );
  AOI21_X1 U6724 ( .B1(n5622), .B2(n6186), .A(n5621), .ZN(n5623) );
  OAI21_X1 U6725 ( .B1(n6193), .B2(n5893), .A(n5623), .ZN(U2971) );
  AOI21_X1 U6726 ( .B1(n5631), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5625) );
  OAI21_X1 U6727 ( .B1(n5626), .B2(n5625), .A(n5624), .ZN(n5627) );
  AOI21_X1 U6728 ( .B1(n5628), .B2(n6240), .A(n5627), .ZN(n5629) );
  OAI21_X1 U6729 ( .B1(n5630), .B2(n5717), .A(n5629), .ZN(U2988) );
  INV_X1 U6730 ( .A(n5631), .ZN(n5635) );
  NAND2_X1 U6731 ( .A1(n5632), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5634) );
  OAI211_X1 U6732 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n5635), .A(n5634), .B(n5633), .ZN(n5636) );
  AOI21_X1 U6733 ( .B1(n5637), .B2(n6240), .A(n5636), .ZN(n5638) );
  OAI21_X1 U6734 ( .B1(n3002), .B2(n5717), .A(n5638), .ZN(U2989) );
  INV_X1 U6735 ( .A(n5639), .ZN(n5655) );
  XNOR2_X1 U6736 ( .A(n5640), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5641)
         );
  NAND2_X1 U6737 ( .A1(n5651), .A2(n5641), .ZN(n5642) );
  OAI211_X1 U6738 ( .C1(n5741), .C2(n3628), .A(n5643), .B(n5642), .ZN(n5644)
         );
  AOI21_X1 U6739 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5655), .A(n5644), 
        .ZN(n5645) );
  OAI21_X1 U6740 ( .B1(n5646), .B2(n5717), .A(n5645), .ZN(U2990) );
  AND2_X1 U6741 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  OR2_X1 U6742 ( .A1(n5451), .A2(n5649), .ZN(n5818) );
  NAND2_X1 U6743 ( .A1(n5651), .A2(n5650), .ZN(n5652) );
  OAI211_X1 U6744 ( .C1(n5818), .C2(n3628), .A(n5653), .B(n5652), .ZN(n5654)
         );
  AOI21_X1 U6745 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5655), .A(n5654), 
        .ZN(n5656) );
  OAI21_X1 U6746 ( .B1(n5657), .B2(n5717), .A(n5656), .ZN(U2991) );
  INV_X1 U6747 ( .A(n5875), .ZN(n5658) );
  AOI21_X1 U6748 ( .B1(n5659), .B2(n6612), .A(n5658), .ZN(n5660) );
  NAND2_X1 U6749 ( .A1(n5661), .A2(n5660), .ZN(n5662) );
  OAI211_X1 U6750 ( .C1(n5750), .C2(n3628), .A(n5663), .B(n5662), .ZN(n5664)
         );
  AOI21_X1 U6751 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5874), .A(n5664), 
        .ZN(n5665) );
  OAI21_X1 U6752 ( .B1(n5666), .B2(n5717), .A(n5665), .ZN(U2992) );
  INV_X1 U6753 ( .A(n5667), .ZN(n5673) );
  NAND3_X1 U6754 ( .A1(n5678), .A2(n5679), .A3(n5668), .ZN(n5669) );
  OAI211_X1 U6755 ( .C1(n5671), .C2(n3628), .A(n5670), .B(n5669), .ZN(n5672)
         );
  AOI21_X1 U6756 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5673), .A(n5672), 
        .ZN(n5674) );
  OAI21_X1 U6757 ( .B1(n5675), .B2(n5717), .A(n5674), .ZN(U2995) );
  INV_X1 U6758 ( .A(n5676), .ZN(n5689) );
  OAI21_X1 U6759 ( .B1(n5785), .B2(n3628), .A(n5677), .ZN(n5682) );
  INV_X1 U6760 ( .A(n5678), .ZN(n5686) );
  NOR3_X1 U6761 ( .A1(n5686), .A2(n5680), .A3(n5679), .ZN(n5681) );
  AOI211_X1 U6762 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5689), .A(n5682), .B(n5681), .ZN(n5683) );
  OAI21_X1 U6763 ( .B1(n5684), .B2(n5717), .A(n5683), .ZN(U2996) );
  OAI21_X1 U6764 ( .B1(n5790), .B2(n3628), .A(n5685), .ZN(n5688) );
  NOR2_X1 U6765 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5687)
         );
  AOI211_X1 U6766 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5689), .A(n5688), .B(n5687), .ZN(n5690) );
  OAI21_X1 U6767 ( .B1(n5691), .B2(n5717), .A(n5690), .ZN(U2997) );
  INV_X1 U6768 ( .A(n5805), .ZN(n5697) );
  INV_X1 U6769 ( .A(n5692), .ZN(n5696) );
  NOR3_X1 U6770 ( .A1(n5694), .A2(n5693), .A3(n5714), .ZN(n5695) );
  AOI211_X1 U6771 ( .C1(n5697), .C2(n6240), .A(n5696), .B(n5695), .ZN(n5706)
         );
  NAND2_X1 U6772 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  NAND2_X1 U6773 ( .A1(n5700), .A2(n5719), .ZN(n5701) );
  AND2_X1 U6774 ( .A1(n5702), .A2(n5701), .ZN(n5727) );
  NAND2_X1 U6775 ( .A1(n5883), .A2(n5726), .ZN(n5703) );
  AND2_X1 U6776 ( .A1(n5727), .A2(n5703), .ZN(n5712) );
  INV_X1 U6777 ( .A(n5712), .ZN(n5704) );
  NAND2_X1 U6778 ( .A1(n5704), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5705) );
  OAI211_X1 U6779 ( .C1(n5707), .C2(n5717), .A(n5706), .B(n5705), .ZN(U2998)
         );
  XNOR2_X1 U6780 ( .A(n5708), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5709)
         );
  XNOR2_X1 U6781 ( .A(n5710), .B(n5709), .ZN(n5861) );
  NAND2_X1 U6782 ( .A1(n6238), .A2(REIP_REG_19__SCAN_IN), .ZN(n5711) );
  OAI221_X1 U6783 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5714), .C1(
        n5713), .C2(n5712), .A(n5711), .ZN(n5715) );
  AOI21_X1 U6784 ( .B1(n6240), .B2(n5807), .A(n5715), .ZN(n5716) );
  OAI21_X1 U6785 ( .B1(n5861), .B2(n5717), .A(n5716), .ZN(U2999) );
  NAND2_X1 U6786 ( .A1(n5718), .A2(n6245), .ZN(n5725) );
  INV_X1 U6787 ( .A(n5937), .ZN(n5723) );
  NOR3_X1 U6788 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5720), .A3(n5719), 
        .ZN(n5721) );
  AOI211_X1 U6789 ( .C1(n5723), .C2(n6240), .A(n5722), .B(n5721), .ZN(n5724)
         );
  OAI211_X1 U6790 ( .C1(n5727), .C2(n5726), .A(n5725), .B(n5724), .ZN(U3000)
         );
  NOR2_X1 U6791 ( .A1(n5729), .A2(n5728), .ZN(n5730) );
  NOR2_X1 U6792 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5732), .ZN(n6096) );
  INV_X1 U6793 ( .A(n6096), .ZN(n6559) );
  INV_X1 U6794 ( .A(n6559), .ZN(n6103) );
  AND2_X1 U6795 ( .A1(n6102), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6796 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6628) );
  NOR3_X1 U6797 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6628), .A3(n5733), .ZN(n5737) );
  INV_X1 U6798 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6514) );
  OAI22_X1 U6799 ( .A1(n5735), .A2(n6514), .B1(n5734), .B2(n6004), .ZN(n5736)
         );
  AOI211_X1 U6800 ( .C1(n5993), .C2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5737), 
        .B(n5736), .ZN(n5740) );
  AOI22_X1 U6801 ( .A1(n5823), .A2(n6001), .B1(n5738), .B2(n5999), .ZN(n5739)
         );
  OAI211_X1 U6802 ( .C1(n5741), .C2(n6031), .A(n5740), .B(n5739), .ZN(U2799)
         );
  INV_X1 U6803 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5822) );
  OAI22_X1 U6804 ( .A1(n5822), .A2(n6004), .B1(n4117), .B2(n6018), .ZN(n5742)
         );
  AOI221_X1 U6805 ( .B1(n5754), .B2(REIP_REG_27__SCAN_IN), .C1(n5743), .C2(
        n6628), .A(n5742), .ZN(n5746) );
  OAI22_X1 U6806 ( .A1(n5827), .A2(n5955), .B1(n5818), .B2(n6031), .ZN(n5744)
         );
  INV_X1 U6807 ( .A(n5744), .ZN(n5745) );
  OAI211_X1 U6808 ( .C1(n5747), .C2(n6037), .A(n5746), .B(n5745), .ZN(U2800)
         );
  AOI22_X1 U6809 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6028), .B1(n5748), .B2(n5999), .ZN(n5756) );
  NAND2_X1 U6810 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5749), .ZN(n5759) );
  OAI21_X1 U6811 ( .B1(n6511), .B2(n5759), .A(n6513), .ZN(n5753) );
  OAI22_X1 U6812 ( .A1(n5751), .A2(n5955), .B1(n6031), .B2(n5750), .ZN(n5752)
         );
  AOI21_X1 U6813 ( .B1(n5754), .B2(n5753), .A(n5752), .ZN(n5755) );
  OAI211_X1 U6814 ( .C1(n5757), .C2(n6018), .A(n5756), .B(n5755), .ZN(U2801)
         );
  INV_X1 U6815 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5758) );
  OAI22_X1 U6816 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5759), .B1(n5758), .B2(
        n6018), .ZN(n5762) );
  OAI22_X1 U6817 ( .A1(n5760), .A2(n5955), .B1(n6031), .B2(n5876), .ZN(n5761)
         );
  AOI211_X1 U6818 ( .C1(EBX_REG_25__SCAN_IN), .C2(n6028), .A(n5762), .B(n5761), 
        .ZN(n5765) );
  NOR2_X1 U6819 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5763), .ZN(n5767) );
  OAI21_X1 U6820 ( .B1(n5768), .B2(n5767), .A(REIP_REG_25__SCAN_IN), .ZN(n5764) );
  OAI211_X1 U6821 ( .C1(n6037), .C2(n5860), .A(n5765), .B(n5764), .ZN(U2802)
         );
  OAI22_X1 U6822 ( .A1(n6671), .A2(n6004), .B1(n5562), .B2(n6018), .ZN(n5766)
         );
  AOI211_X1 U6823 ( .C1(n5768), .C2(REIP_REG_24__SCAN_IN), .A(n5767), .B(n5766), .ZN(n5772) );
  INV_X1 U6824 ( .A(n5769), .ZN(n5833) );
  AOI22_X1 U6825 ( .A1(n5833), .A2(n6001), .B1(n5770), .B2(n5999), .ZN(n5771)
         );
  OAI211_X1 U6826 ( .C1(n5773), .C2(n6031), .A(n5772), .B(n5771), .ZN(U2803)
         );
  NAND2_X1 U6827 ( .A1(n5775), .A2(n5774), .ZN(n5797) );
  INV_X1 U6828 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U6829 ( .A1(n5776), .A2(n6505), .ZN(n5786) );
  AOI21_X1 U6830 ( .B1(n5797), .B2(n5786), .A(n6507), .ZN(n5779) );
  OAI22_X1 U6831 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5777), .B1(n6721), .B2(
        n6004), .ZN(n5778) );
  AOI211_X1 U6832 ( .C1(n5993), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5779), 
        .B(n5778), .ZN(n5784) );
  INV_X1 U6833 ( .A(n5780), .ZN(n5781) );
  OAI22_X1 U6834 ( .A1(n5840), .A2(n5955), .B1(n5781), .B2(n6037), .ZN(n5782)
         );
  INV_X1 U6835 ( .A(n5782), .ZN(n5783) );
  OAI211_X1 U6836 ( .C1(n5785), .C2(n6031), .A(n5784), .B(n5783), .ZN(U2805)
         );
  INV_X1 U6837 ( .A(n5786), .ZN(n5789) );
  INV_X1 U6838 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5787) );
  OAI22_X1 U6839 ( .A1(n5787), .A2(n6018), .B1(n6505), .B2(n5797), .ZN(n5788)
         );
  AOI211_X1 U6840 ( .C1(n6028), .C2(EBX_REG_21__SCAN_IN), .A(n5789), .B(n5788), 
        .ZN(n5793) );
  INV_X1 U6841 ( .A(n5790), .ZN(n5791) );
  AOI22_X1 U6842 ( .A1(n5844), .A2(n6001), .B1(n6007), .B2(n5791), .ZN(n5792)
         );
  OAI211_X1 U6843 ( .C1(n5794), .C2(n6037), .A(n5793), .B(n5792), .ZN(U2806)
         );
  INV_X1 U6844 ( .A(n5931), .ZN(n5795) );
  INV_X1 U6845 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6502) );
  NOR2_X1 U6846 ( .A1(n6502), .A2(n5602), .ZN(n5808) );
  AOI21_X1 U6847 ( .B1(n5795), .B2(n5808), .A(REIP_REG_20__SCAN_IN), .ZN(n5798) );
  OAI22_X1 U6848 ( .A1(n5798), .A2(n5797), .B1(n5796), .B2(n6018), .ZN(n5799)
         );
  AOI21_X1 U6849 ( .B1(EBX_REG_20__SCAN_IN), .B2(n6028), .A(n5799), .ZN(n5804)
         );
  INV_X1 U6850 ( .A(n5800), .ZN(n5801) );
  OAI22_X1 U6851 ( .A1(n5848), .A2(n5955), .B1(n5801), .B2(n6037), .ZN(n5802)
         );
  INV_X1 U6852 ( .A(n5802), .ZN(n5803) );
  OAI211_X1 U6853 ( .C1(n5805), .C2(n6031), .A(n5804), .B(n5803), .ZN(U2807)
         );
  INV_X1 U6854 ( .A(n5807), .ZN(n5814) );
  AOI211_X1 U6855 ( .C1(n6502), .C2(n5602), .A(n5808), .B(n5931), .ZN(n5809)
         );
  AOI211_X1 U6856 ( .C1(n5993), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5809), 
        .B(n6022), .ZN(n5813) );
  NOR2_X1 U6857 ( .A1(n5811), .A2(n5810), .ZN(n5938) );
  AOI22_X1 U6858 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6028), .B1(
        REIP_REG_19__SCAN_IN), .B2(n5938), .ZN(n5812) );
  OAI211_X1 U6859 ( .C1(n5814), .C2(n6031), .A(n5813), .B(n5812), .ZN(n5815)
         );
  AOI21_X1 U6860 ( .B1(n5862), .B2(n6001), .A(n5815), .ZN(n5816) );
  OAI21_X1 U6861 ( .B1(n5866), .B2(n6037), .A(n5816), .ZN(U2808) );
  OAI22_X1 U6862 ( .A1(n5827), .A2(n5819), .B1(n5818), .B2(n5817), .ZN(n5820)
         );
  INV_X1 U6863 ( .A(n5820), .ZN(n5821) );
  OAI21_X1 U6864 ( .B1(n6045), .B2(n5822), .A(n5821), .ZN(U2832) );
  INV_X1 U6865 ( .A(n6047), .ZN(n6053) );
  AOI22_X1 U6866 ( .A1(n5823), .A2(n6053), .B1(n6052), .B2(DATAI_28_), .ZN(
        n5825) );
  AOI22_X1 U6867 ( .A1(n6062), .A2(DATAI_12_), .B1(n6061), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U6868 ( .A1(n5825), .A2(n5824), .ZN(U2863) );
  INV_X1 U6869 ( .A(n6052), .ZN(n6058) );
  OAI22_X1 U6870 ( .A1(n5827), .A2(n6047), .B1(n6058), .B2(n5826), .ZN(n5828)
         );
  INV_X1 U6871 ( .A(n5828), .ZN(n5830) );
  AOI22_X1 U6872 ( .A1(n6062), .A2(DATAI_11_), .B1(n6061), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U6873 ( .A1(n5830), .A2(n5829), .ZN(U2864) );
  AOI22_X1 U6874 ( .A1(n5857), .A2(n6053), .B1(n6052), .B2(DATAI_25_), .ZN(
        n5832) );
  AOI22_X1 U6875 ( .A1(n6062), .A2(DATAI_9_), .B1(n6061), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U6876 ( .A1(n5832), .A2(n5831), .ZN(U2866) );
  AOI22_X1 U6877 ( .A1(n5833), .A2(n6053), .B1(n6052), .B2(DATAI_24_), .ZN(
        n5835) );
  AOI22_X1 U6878 ( .A1(n6062), .A2(DATAI_8_), .B1(n6061), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U6879 ( .A1(n5835), .A2(n5834), .ZN(U2867) );
  AOI22_X1 U6880 ( .A1(n5836), .A2(n6053), .B1(n6052), .B2(DATAI_23_), .ZN(
        n5838) );
  AOI22_X1 U6881 ( .A1(n6062), .A2(DATAI_7_), .B1(n6061), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U6882 ( .A1(n5838), .A2(n5837), .ZN(U2868) );
  OAI22_X1 U6883 ( .A1(n5840), .A2(n6047), .B1(n6058), .B2(n5839), .ZN(n5841)
         );
  INV_X1 U6884 ( .A(n5841), .ZN(n5843) );
  AOI22_X1 U6885 ( .A1(n6062), .A2(DATAI_6_), .B1(n6061), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U6886 ( .A1(n5843), .A2(n5842), .ZN(U2869) );
  AOI22_X1 U6887 ( .A1(n5844), .A2(n6053), .B1(n6052), .B2(DATAI_21_), .ZN(
        n5846) );
  AOI22_X1 U6888 ( .A1(n6062), .A2(DATAI_5_), .B1(n6061), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U6889 ( .A1(n5846), .A2(n5845), .ZN(U2870) );
  OAI22_X1 U6890 ( .A1(n5848), .A2(n6047), .B1(n6058), .B2(n5847), .ZN(n5849)
         );
  INV_X1 U6891 ( .A(n5849), .ZN(n5851) );
  AOI22_X1 U6892 ( .A1(n6062), .A2(DATAI_4_), .B1(n6061), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U6893 ( .A1(n5851), .A2(n5850), .ZN(U2871) );
  AOI22_X1 U6894 ( .A1(n5862), .A2(n6053), .B1(n6052), .B2(DATAI_19_), .ZN(
        n5853) );
  AOI22_X1 U6895 ( .A1(n6062), .A2(DATAI_3_), .B1(n6061), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U6896 ( .A1(n5853), .A2(n5852), .ZN(U2872) );
  AOI22_X1 U6897 ( .A1(n6238), .A2(REIP_REG_25__SCAN_IN), .B1(n6197), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5859) );
  OAI21_X1 U6898 ( .B1(n5856), .B2(n5855), .A(n5854), .ZN(n5878) );
  AOI22_X1 U6899 ( .A1(n5857), .A2(n6186), .B1(n6185), .B2(n5878), .ZN(n5858)
         );
  OAI211_X1 U6900 ( .C1(n6191), .C2(n5860), .A(n5859), .B(n5858), .ZN(U2961)
         );
  AOI22_X1 U6901 ( .A1(n6238), .A2(REIP_REG_19__SCAN_IN), .B1(n6197), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5865) );
  INV_X1 U6902 ( .A(n5861), .ZN(n5863) );
  AOI22_X1 U6903 ( .A1(n5863), .A2(n6185), .B1(n6186), .B2(n5862), .ZN(n5864)
         );
  OAI211_X1 U6904 ( .C1(n6191), .C2(n5866), .A(n5865), .B(n5864), .ZN(U2967)
         );
  INV_X1 U6905 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5939) );
  INV_X1 U6906 ( .A(n5867), .ZN(n5870) );
  INV_X1 U6907 ( .A(n5947), .ZN(n5869) );
  AOI222_X1 U6908 ( .A1(n5870), .A2(n6185), .B1(n5869), .B2(n5868), .C1(n6186), 
        .C2(n6054), .ZN(n5872) );
  OAI211_X1 U6909 ( .C1(n5939), .C2(n5873), .A(n5872), .B(n5871), .ZN(U2969)
         );
  INV_X1 U6910 ( .A(n5874), .ZN(n5881) );
  AOI22_X1 U6911 ( .A1(n6238), .A2(REIP_REG_25__SCAN_IN), .B1(n5875), .B2(
        n6612), .ZN(n5880) );
  INV_X1 U6912 ( .A(n5876), .ZN(n5877) );
  AOI22_X1 U6913 ( .A1(n5878), .A2(n6245), .B1(n6240), .B2(n5877), .ZN(n5879)
         );
  OAI211_X1 U6914 ( .C1(n5881), .C2(n6612), .A(n5880), .B(n5879), .ZN(U2993)
         );
  INV_X1 U6915 ( .A(n5882), .ZN(n5886) );
  INV_X1 U6916 ( .A(n5959), .ZN(n5885) );
  AND2_X1 U6917 ( .A1(n5883), .A2(n5887), .ZN(n5884) );
  OR2_X1 U6918 ( .A1(n6204), .A2(n5884), .ZN(n5891) );
  AOI222_X1 U6919 ( .A1(n5886), .A2(n6245), .B1(n6240), .B2(n5885), .C1(n5891), 
        .C2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5890) );
  NOR2_X1 U6920 ( .A1(n6208), .A2(n5887), .ZN(n5892) );
  OAI211_X1 U6921 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5892), .B(n5888), .ZN(n5889) );
  OAI211_X1 U6922 ( .C1(n5608), .C2(n6192), .A(n5890), .B(n5889), .ZN(U3002)
         );
  INV_X1 U6923 ( .A(n5891), .ZN(n5899) );
  AOI22_X1 U6924 ( .A1(n6238), .A2(REIP_REG_15__SCAN_IN), .B1(n5892), .B2(
        n5898), .ZN(n5897) );
  INV_X1 U6925 ( .A(n5893), .ZN(n5895) );
  AOI22_X1 U6926 ( .A1(n5895), .A2(n6245), .B1(n6240), .B2(n5894), .ZN(n5896)
         );
  OAI211_X1 U6927 ( .C1(n5899), .C2(n5898), .A(n5897), .B(n5896), .ZN(U3003)
         );
  INV_X1 U6928 ( .A(n5900), .ZN(n5901) );
  NAND4_X1 U6929 ( .A1(n6024), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(n5904)
         );
  OAI21_X1 U6930 ( .B1(n5906), .B2(n5905), .A(n5904), .ZN(U3455) );
  AOI21_X1 U6931 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6455), .A(n3422), .ZN(n5911) );
  INV_X1 U6932 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5907) );
  NOR2_X2 U6933 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6463), .ZN(n6570) );
  AOI21_X1 U6934 ( .B1(n5911), .B2(n5907), .A(n6570), .ZN(U2789) );
  OAI21_X1 U6935 ( .B1(n5908), .B2(n6445), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5909) );
  OAI21_X1 U6936 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6444), .A(n5909), .ZN(
        U2790) );
  NOR2_X1 U6937 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5912) );
  OAI21_X1 U6938 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5912), .A(n6556), .ZN(n5910)
         );
  OAI21_X1 U6939 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6556), .A(n5910), .ZN(
        U2791) );
  NOR2_X1 U6940 ( .A1(n6570), .A2(n5911), .ZN(n6530) );
  OAI21_X1 U6941 ( .B1(BS16_N), .B2(n5912), .A(n6530), .ZN(n6528) );
  OAI21_X1 U6942 ( .B1(n6530), .B2(n6561), .A(n6528), .ZN(U2792) );
  OAI21_X1 U6943 ( .B1(n5914), .B2(n5913), .A(n6193), .ZN(U2793) );
  NOR4_X1 U6944 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5918) );
  NOR4_X1 U6945 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5917) );
  NOR4_X1 U6946 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5916) );
  NOR4_X1 U6947 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5915) );
  NAND4_X1 U6948 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n5924)
         );
  NOR4_X1 U6949 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n5922) );
  AOI211_X1 U6950 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_12__SCAN_IN), .B(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n5921) );
  NOR4_X1 U6951 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5920) );
  NOR4_X1 U6952 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n5919) );
  NAND4_X1 U6953 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(n5923)
         );
  NOR2_X1 U6954 ( .A1(n5924), .A2(n5923), .ZN(n6550) );
  INV_X1 U6955 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5926) );
  NOR3_X1 U6956 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5927) );
  OAI21_X1 U6957 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5927), .A(n6550), .ZN(n5925)
         );
  OAI21_X1 U6958 ( .B1(n6550), .B2(n5926), .A(n5925), .ZN(U2794) );
  INV_X1 U6959 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6546) );
  INV_X1 U6960 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6529) );
  AOI21_X1 U6961 ( .B1(n6546), .B2(n6529), .A(n5927), .ZN(n5929) );
  INV_X1 U6962 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5928) );
  INV_X1 U6963 ( .A(n6550), .ZN(n6553) );
  AOI22_X1 U6964 ( .A1(n6550), .A2(n5929), .B1(n5928), .B2(n6553), .ZN(U2795)
         );
  AOI22_X1 U6965 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6028), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5938), .ZN(n5930) );
  OAI21_X1 U6966 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5931), .A(n5930), .ZN(n5932) );
  AOI211_X1 U6967 ( .C1(n5993), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6022), 
        .B(n5932), .ZN(n5936) );
  OAI22_X1 U6968 ( .A1(n6048), .A2(n5955), .B1(n5933), .B2(n6037), .ZN(n5934)
         );
  INV_X1 U6969 ( .A(n5934), .ZN(n5935) );
  OAI211_X1 U6970 ( .C1(n6031), .C2(n5937), .A(n5936), .B(n5935), .ZN(U2809)
         );
  NOR2_X1 U6971 ( .A1(n5608), .A2(n6497), .ZN(n5948) );
  AOI21_X1 U6972 ( .B1(n5950), .B2(n5948), .A(REIP_REG_17__SCAN_IN), .ZN(n5941) );
  INV_X1 U6973 ( .A(n5938), .ZN(n5940) );
  OAI22_X1 U6974 ( .A1(n5941), .A2(n5940), .B1(n5939), .B2(n6018), .ZN(n5942)
         );
  AOI211_X1 U6975 ( .C1(n6028), .C2(EBX_REG_17__SCAN_IN), .A(n6022), .B(n5942), 
        .ZN(n5946) );
  NOR2_X1 U6976 ( .A1(n5943), .A2(n6031), .ZN(n5944) );
  AOI21_X1 U6977 ( .B1(n6054), .B2(n6001), .A(n5944), .ZN(n5945) );
  OAI211_X1 U6978 ( .C1(n5947), .C2(n6037), .A(n5946), .B(n5945), .ZN(U2810)
         );
  AOI21_X1 U6979 ( .B1(n5608), .B2(n6497), .A(n5948), .ZN(n5949) );
  AOI22_X1 U6980 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6028), .B1(n5950), .B2(n5949), .ZN(n5951) );
  OAI21_X1 U6981 ( .B1(n5964), .B2(n5608), .A(n5951), .ZN(n5952) );
  AOI211_X1 U6982 ( .C1(n5993), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6022), 
        .B(n5952), .ZN(n5958) );
  INV_X1 U6983 ( .A(n5953), .ZN(n5954) );
  OAI22_X1 U6984 ( .A1(n6059), .A2(n5955), .B1(n5954), .B2(n6037), .ZN(n5956)
         );
  INV_X1 U6985 ( .A(n5956), .ZN(n5957) );
  OAI211_X1 U6986 ( .C1(n6031), .C2(n5959), .A(n5958), .B(n5957), .ZN(U2811)
         );
  AND2_X1 U6987 ( .A1(n5960), .A2(n6009), .ZN(n5961) );
  AOI22_X1 U6988 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6028), .B1(n5962), .B2(n5961), .ZN(n5963) );
  OAI21_X1 U6989 ( .B1(n5964), .B2(n6494), .A(n5963), .ZN(n5965) );
  AOI211_X1 U6990 ( .C1(n5993), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6022), 
        .B(n5965), .ZN(n5970) );
  INV_X1 U6991 ( .A(n5966), .ZN(n5967) );
  AOI22_X1 U6992 ( .A1(n5968), .A2(n6001), .B1(n5967), .B2(n5999), .ZN(n5969)
         );
  OAI211_X1 U6993 ( .C1(n6031), .C2(n5971), .A(n5970), .B(n5969), .ZN(U2813)
         );
  AOI22_X1 U6994 ( .A1(n6007), .A2(n5973), .B1(REIP_REG_12__SCAN_IN), .B2(
        n5972), .ZN(n5981) );
  AOI22_X1 U6995 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6028), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5993), .ZN(n5980) );
  NOR2_X1 U6996 ( .A1(n6026), .A2(n5974), .ZN(n5975) );
  AOI21_X1 U6997 ( .B1(n5975), .B2(n6705), .A(n6022), .ZN(n5979) );
  AOI22_X1 U6998 ( .A1(n5977), .A2(n6001), .B1(n5999), .B2(n5976), .ZN(n5978)
         );
  NAND4_X1 U6999 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(U2815)
         );
  INV_X1 U7000 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6480) );
  NOR3_X1 U7001 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6480), .A3(n5989), .ZN(n5984)
         );
  INV_X1 U7002 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6645) );
  AOI22_X1 U7003 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6028), .B1(n6007), .B2(n6218), 
        .ZN(n5982) );
  OAI211_X1 U7004 ( .C1(n6018), .C2(n6645), .A(n5994), .B(n5982), .ZN(n5983)
         );
  AOI211_X1 U7005 ( .C1(n5985), .C2(n6001), .A(n5984), .B(n5983), .ZN(n5991)
         );
  INV_X1 U7006 ( .A(n5986), .ZN(n5988) );
  OAI21_X1 U7007 ( .B1(n6026), .B2(n5988), .A(n5987), .ZN(n6012) );
  NOR2_X1 U7008 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5989), .ZN(n5997) );
  OAI21_X1 U7009 ( .B1(n6012), .B2(n5997), .A(REIP_REG_7__SCAN_IN), .ZN(n5990)
         );
  OAI211_X1 U7010 ( .C1(n6037), .C2(n5992), .A(n5991), .B(n5990), .ZN(U2820)
         );
  AOI22_X1 U7011 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n5993), .B1(n6007), 
        .B2(n6039), .ZN(n5995) );
  OAI211_X1 U7012 ( .C1(n6004), .C2(n6044), .A(n5995), .B(n5994), .ZN(n5996)
         );
  AOI211_X1 U7013 ( .C1(n6012), .C2(REIP_REG_6__SCAN_IN), .A(n5997), .B(n5996), 
        .ZN(n6003) );
  INV_X1 U7014 ( .A(n5998), .ZN(n6000) );
  AOI22_X1 U7015 ( .A1(n6042), .A2(n6001), .B1(n6000), .B2(n5999), .ZN(n6002)
         );
  NAND2_X1 U7016 ( .A1(n6003), .A2(n6002), .ZN(U2821) );
  OAI22_X1 U7017 ( .A1(n6691), .A2(n6004), .B1(n3728), .B2(n6018), .ZN(n6005)
         );
  AOI211_X1 U7018 ( .C1(n6007), .C2(n6006), .A(n6022), .B(n6005), .ZN(n6016)
         );
  INV_X1 U7019 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7020 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  NAND2_X1 U7021 ( .A1(n6011), .A2(n6010), .ZN(n6013) );
  AOI22_X1 U7022 ( .A1(n6014), .A2(n6033), .B1(n6013), .B2(n6012), .ZN(n6015)
         );
  OAI211_X1 U7023 ( .C1(n6017), .C2(n6037), .A(n6016), .B(n6015), .ZN(U2822)
         );
  OAI22_X1 U7024 ( .A1(n6020), .A2(n6478), .B1(n6019), .B2(n6018), .ZN(n6021)
         );
  AOI211_X1 U7025 ( .C1(n6024), .C2(n6023), .A(n6022), .B(n6021), .ZN(n6036)
         );
  NOR3_X1 U7026 ( .A1(n6026), .A2(REIP_REG_4__SCAN_IN), .A3(n6025), .ZN(n6027)
         );
  AOI21_X1 U7027 ( .B1(n6028), .B2(EBX_REG_4__SCAN_IN), .A(n6027), .ZN(n6029)
         );
  OAI21_X1 U7028 ( .B1(n6031), .B2(n6030), .A(n6029), .ZN(n6032) );
  AOI21_X1 U7029 ( .B1(n6034), .B2(n6033), .A(n6032), .ZN(n6035) );
  OAI211_X1 U7030 ( .C1(n6038), .C2(n6037), .A(n6036), .B(n6035), .ZN(U2823)
         );
  AOI22_X1 U7031 ( .A1(n6042), .A2(n6041), .B1(n6040), .B2(n6039), .ZN(n6043)
         );
  OAI21_X1 U7032 ( .B1(n6045), .B2(n6044), .A(n6043), .ZN(U2853) );
  OAI22_X1 U7033 ( .A1(n6048), .A2(n6047), .B1(n6058), .B2(n6046), .ZN(n6049)
         );
  INV_X1 U7034 ( .A(n6049), .ZN(n6051) );
  AOI22_X1 U7035 ( .A1(n6062), .A2(DATAI_2_), .B1(n6061), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7036 ( .A1(n6051), .A2(n6050), .ZN(U2873) );
  AOI22_X1 U7037 ( .A1(n6054), .A2(n6053), .B1(n6052), .B2(DATAI_17_), .ZN(
        n6056) );
  AOI22_X1 U7038 ( .A1(n6062), .A2(DATAI_1_), .B1(n6061), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7039 ( .A1(n6056), .A2(n6055), .ZN(U2874) );
  OAI22_X1 U7040 ( .A1(n6059), .A2(n6047), .B1(n6058), .B2(n6057), .ZN(n6060)
         );
  INV_X1 U7041 ( .A(n6060), .ZN(n6064) );
  AOI22_X1 U7042 ( .A1(n6062), .A2(DATAI_0_), .B1(n6061), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7043 ( .A1(n6064), .A2(n6063), .ZN(U2875) );
  INV_X1 U7044 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7045 ( .A1(n6091), .A2(n6065), .ZN(n6082) );
  AOI22_X1 U7046 ( .A1(n6103), .A2(UWORD_REG_14__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n6066) );
  OAI21_X1 U7047 ( .B1(n6142), .B2(n6082), .A(n6066), .ZN(U2893) );
  INV_X1 U7048 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6138) );
  AOI22_X1 U7049 ( .A1(DATAO_REG_29__SCAN_IN), .A2(n6100), .B1(n6096), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n6067) );
  OAI21_X1 U7050 ( .B1(n6138), .B2(n6082), .A(n6067), .ZN(U2894) );
  INV_X1 U7051 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6136) );
  AOI22_X1 U7052 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6096), .B1(
        DATAO_REG_28__SCAN_IN), .B2(n6100), .ZN(n6068) );
  OAI21_X1 U7053 ( .B1(n6136), .B2(n6082), .A(n6068), .ZN(U2895) );
  INV_X1 U7054 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6133) );
  AOI22_X1 U7055 ( .A1(n6096), .A2(UWORD_REG_11__SCAN_IN), .B1(n6102), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n6069) );
  OAI21_X1 U7056 ( .B1(n6133), .B2(n6082), .A(n6069), .ZN(U2896) );
  INV_X1 U7057 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6130) );
  AOI22_X1 U7058 ( .A1(n6103), .A2(UWORD_REG_10__SCAN_IN), .B1(n6102), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n6070) );
  OAI21_X1 U7059 ( .B1(n6130), .B2(n6082), .A(n6070), .ZN(U2897) );
  INV_X1 U7060 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6127) );
  AOI22_X1 U7061 ( .A1(n6103), .A2(UWORD_REG_9__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n6071) );
  OAI21_X1 U7062 ( .B1(n6127), .B2(n6082), .A(n6071), .ZN(U2898) );
  INV_X1 U7063 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6125) );
  AOI22_X1 U7064 ( .A1(n6103), .A2(UWORD_REG_8__SCAN_IN), .B1(n6102), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n6072) );
  OAI21_X1 U7065 ( .B1(n6125), .B2(n6082), .A(n6072), .ZN(U2899) );
  INV_X1 U7066 ( .A(n6082), .ZN(n6073) );
  AOI22_X1 U7067 ( .A1(EAX_REG_23__SCAN_IN), .A2(n6073), .B1(n6102), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n6074) );
  OAI21_X1 U7068 ( .B1(n6742), .B2(n6559), .A(n6074), .ZN(U2900) );
  INV_X1 U7069 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6122) );
  AOI22_X1 U7070 ( .A1(DATAO_REG_22__SCAN_IN), .A2(n6100), .B1(
        UWORD_REG_6__SCAN_IN), .B2(n6103), .ZN(n6075) );
  OAI21_X1 U7071 ( .B1(n6122), .B2(n6082), .A(n6075), .ZN(U2901) );
  INV_X1 U7072 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6119) );
  AOI22_X1 U7073 ( .A1(n6103), .A2(UWORD_REG_5__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n6076) );
  OAI21_X1 U7074 ( .B1(n6119), .B2(n6082), .A(n6076), .ZN(U2902) );
  INV_X1 U7075 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6117) );
  AOI22_X1 U7076 ( .A1(DATAO_REG_20__SCAN_IN), .A2(n6100), .B1(n6096), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n6077) );
  OAI21_X1 U7077 ( .B1(n6117), .B2(n6082), .A(n6077), .ZN(U2903) );
  AOI22_X1 U7078 ( .A1(n6103), .A2(UWORD_REG_3__SCAN_IN), .B1(n6102), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n6078) );
  OAI21_X1 U7079 ( .B1(n3869), .B2(n6082), .A(n6078), .ZN(U2904) );
  INV_X1 U7080 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6112) );
  AOI22_X1 U7081 ( .A1(n6103), .A2(UWORD_REG_2__SCAN_IN), .B1(n6102), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n6079) );
  OAI21_X1 U7082 ( .B1(n6112), .B2(n6082), .A(n6079), .ZN(U2905) );
  INV_X1 U7083 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6109) );
  AOI22_X1 U7084 ( .A1(DATAO_REG_17__SCAN_IN), .A2(n6100), .B1(n6096), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n6080) );
  OAI21_X1 U7085 ( .B1(n6109), .B2(n6082), .A(n6080), .ZN(U2906) );
  INV_X1 U7086 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6107) );
  AOI22_X1 U7087 ( .A1(n6103), .A2(UWORD_REG_0__SCAN_IN), .B1(n6102), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n6081) );
  OAI21_X1 U7088 ( .B1(n6107), .B2(n6082), .A(n6081), .ZN(U2907) );
  INV_X1 U7089 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6181) );
  AOI22_X1 U7090 ( .A1(DATAO_REG_15__SCAN_IN), .A2(n6100), .B1(n6096), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6083) );
  OAI21_X1 U7091 ( .B1(n6181), .B2(n6105), .A(n6083), .ZN(U2908) );
  INV_X1 U7092 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6176) );
  AOI22_X1 U7093 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6096), .B1(n6100), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6084) );
  OAI21_X1 U7094 ( .B1(n6176), .B2(n6105), .A(n6084), .ZN(U2909) );
  AOI22_X1 U7095 ( .A1(DATAO_REG_13__SCAN_IN), .A2(n6100), .B1(n6096), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6085) );
  OAI21_X1 U7096 ( .B1(n6173), .B2(n6105), .A(n6085), .ZN(U2910) );
  AOI22_X1 U7097 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6091), .B1(n6102), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6086) );
  OAI21_X1 U7098 ( .B1(n6675), .B2(n6559), .A(n6086), .ZN(U2911) );
  INV_X1 U7099 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6170) );
  AOI22_X1 U7100 ( .A1(n6103), .A2(LWORD_REG_11__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6087) );
  OAI21_X1 U7101 ( .B1(n6170), .B2(n6105), .A(n6087), .ZN(U2912) );
  INV_X1 U7102 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6167) );
  AOI22_X1 U7103 ( .A1(n6103), .A2(LWORD_REG_10__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6088) );
  OAI21_X1 U7104 ( .B1(n6167), .B2(n6105), .A(n6088), .ZN(U2913) );
  AOI22_X1 U7105 ( .A1(n6103), .A2(LWORD_REG_9__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6089) );
  OAI21_X1 U7106 ( .B1(n6164), .B2(n6105), .A(n6089), .ZN(U2914) );
  INV_X1 U7107 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6161) );
  AOI22_X1 U7108 ( .A1(n6103), .A2(LWORD_REG_8__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6090) );
  OAI21_X1 U7109 ( .B1(n6161), .B2(n6105), .A(n6090), .ZN(U2915) );
  AOI22_X1 U7110 ( .A1(EAX_REG_7__SCAN_IN), .A2(n6091), .B1(n6102), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6092) );
  OAI21_X1 U7111 ( .B1(n6724), .B2(n6559), .A(n6092), .ZN(U2916) );
  AOI22_X1 U7112 ( .A1(DATAO_REG_6__SCAN_IN), .A2(n6100), .B1(n6096), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n6093) );
  OAI21_X1 U7113 ( .B1(n4790), .B2(n6105), .A(n6093), .ZN(U2917) );
  AOI22_X1 U7114 ( .A1(n6103), .A2(LWORD_REG_5__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6094) );
  OAI21_X1 U7115 ( .B1(n3734), .B2(n6105), .A(n6094), .ZN(U2918) );
  AOI22_X1 U7116 ( .A1(n6103), .A2(LWORD_REG_4__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6095) );
  OAI21_X1 U7117 ( .B1(n6154), .B2(n6105), .A(n6095), .ZN(U2919) );
  AOI22_X1 U7118 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6096), .B1(n6100), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6097) );
  OAI21_X1 U7119 ( .B1(n6098), .B2(n6105), .A(n6097), .ZN(U2920) );
  AOI22_X1 U7120 ( .A1(n6103), .A2(LWORD_REG_2__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6099) );
  OAI21_X1 U7121 ( .B1(n6151), .B2(n6105), .A(n6099), .ZN(U2921) );
  AOI22_X1 U7122 ( .A1(n6103), .A2(LWORD_REG_1__SCAN_IN), .B1(n6100), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6101) );
  OAI21_X1 U7123 ( .B1(n6148), .B2(n6105), .A(n6101), .ZN(U2922) );
  AOI22_X1 U7124 ( .A1(n6103), .A2(LWORD_REG_0__SCAN_IN), .B1(n6102), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6104) );
  OAI21_X1 U7125 ( .B1(n6145), .B2(n6105), .A(n6104), .ZN(U2923) );
  AND2_X1 U7126 ( .A1(n6177), .A2(DATAI_0_), .ZN(n6143) );
  AOI21_X1 U7127 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6110), .A(n6143), .ZN(n6106) );
  OAI21_X1 U7128 ( .B1(n6107), .B2(n6180), .A(n6106), .ZN(U2924) );
  AND2_X1 U7129 ( .A1(n6177), .A2(DATAI_1_), .ZN(n6146) );
  AOI21_X1 U7130 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6110), .A(n6146), .ZN(n6108) );
  OAI21_X1 U7131 ( .B1(n6109), .B2(n6180), .A(n6108), .ZN(U2925) );
  AND2_X1 U7132 ( .A1(n6177), .A2(DATAI_2_), .ZN(n6149) );
  AOI21_X1 U7133 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6110), .A(n6149), .ZN(n6111) );
  OAI21_X1 U7134 ( .B1(n6112), .B2(n6180), .A(n6111), .ZN(U2926) );
  AOI21_X1 U7135 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6178), .A(n6113), .ZN(n6114) );
  OAI21_X1 U7136 ( .B1(n3869), .B2(n6180), .A(n6114), .ZN(U2927) );
  AND2_X1 U7137 ( .A1(n6177), .A2(DATAI_4_), .ZN(n6152) );
  AOI21_X1 U7138 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6110), .A(n6152), .ZN(n6116) );
  OAI21_X1 U7139 ( .B1(n6117), .B2(n6180), .A(n6116), .ZN(U2928) );
  AND2_X1 U7140 ( .A1(n6177), .A2(DATAI_5_), .ZN(n6155) );
  AOI21_X1 U7141 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6178), .A(n6155), .ZN(n6118) );
  OAI21_X1 U7142 ( .B1(n6119), .B2(n6180), .A(n6118), .ZN(U2929) );
  NOR2_X1 U7143 ( .A1(n6140), .A2(n6120), .ZN(n6157) );
  AOI21_X1 U7144 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6178), .A(n6157), .ZN(n6121) );
  OAI21_X1 U7145 ( .B1(n6122), .B2(n6180), .A(n6121), .ZN(U2930) );
  INV_X1 U7146 ( .A(DATAI_8_), .ZN(n6123) );
  NOR2_X1 U7147 ( .A1(n6140), .A2(n6123), .ZN(n6159) );
  AOI21_X1 U7148 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6110), .A(n6159), .ZN(n6124) );
  OAI21_X1 U7149 ( .B1(n6125), .B2(n6180), .A(n6124), .ZN(U2932) );
  AND2_X1 U7150 ( .A1(n6177), .A2(DATAI_9_), .ZN(n6162) );
  AOI21_X1 U7151 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6110), .A(n6162), .ZN(n6126) );
  OAI21_X1 U7152 ( .B1(n6127), .B2(n6180), .A(n6126), .ZN(U2933) );
  INV_X1 U7153 ( .A(DATAI_10_), .ZN(n6128) );
  NOR2_X1 U7154 ( .A1(n6140), .A2(n6128), .ZN(n6165) );
  AOI21_X1 U7155 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6110), .A(n6165), .ZN(
        n6129) );
  OAI21_X1 U7156 ( .B1(n6130), .B2(n6180), .A(n6129), .ZN(U2934) );
  INV_X1 U7157 ( .A(DATAI_11_), .ZN(n6131) );
  NOR2_X1 U7158 ( .A1(n6140), .A2(n6131), .ZN(n6168) );
  AOI21_X1 U7159 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6110), .A(n6168), .ZN(
        n6132) );
  OAI21_X1 U7160 ( .B1(n6133), .B2(n6180), .A(n6132), .ZN(U2935) );
  AOI21_X1 U7161 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6110), .A(n6134), .ZN(
        n6135) );
  OAI21_X1 U7162 ( .B1(n6136), .B2(n6180), .A(n6135), .ZN(U2936) );
  AND2_X1 U7163 ( .A1(n6177), .A2(DATAI_13_), .ZN(n6171) );
  AOI21_X1 U7164 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6178), .A(n6171), .ZN(
        n6137) );
  OAI21_X1 U7165 ( .B1(n6138), .B2(n6180), .A(n6137), .ZN(U2937) );
  INV_X1 U7166 ( .A(DATAI_14_), .ZN(n6139) );
  NOR2_X1 U7167 ( .A1(n6140), .A2(n6139), .ZN(n6174) );
  AOI21_X1 U7168 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6110), .A(n6174), .ZN(
        n6141) );
  OAI21_X1 U7169 ( .B1(n6142), .B2(n6180), .A(n6141), .ZN(U2938) );
  AOI21_X1 U7170 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6178), .A(n6143), .ZN(n6144) );
  OAI21_X1 U7171 ( .B1(n6145), .B2(n6180), .A(n6144), .ZN(U2939) );
  AOI21_X1 U7172 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6178), .A(n6146), .ZN(n6147) );
  OAI21_X1 U7173 ( .B1(n6148), .B2(n6180), .A(n6147), .ZN(U2940) );
  AOI21_X1 U7174 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6178), .A(n6149), .ZN(n6150) );
  OAI21_X1 U7175 ( .B1(n6151), .B2(n6180), .A(n6150), .ZN(U2941) );
  AOI21_X1 U7176 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6178), .A(n6152), .ZN(n6153) );
  OAI21_X1 U7177 ( .B1(n6154), .B2(n6180), .A(n6153), .ZN(U2943) );
  AOI21_X1 U7178 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6178), .A(n6155), .ZN(n6156) );
  OAI21_X1 U7179 ( .B1(n3734), .B2(n6180), .A(n6156), .ZN(U2944) );
  AOI21_X1 U7180 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6178), .A(n6157), .ZN(n6158) );
  OAI21_X1 U7181 ( .B1(n4790), .B2(n6180), .A(n6158), .ZN(U2945) );
  AOI21_X1 U7182 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6178), .A(n6159), .ZN(n6160) );
  OAI21_X1 U7183 ( .B1(n6161), .B2(n6180), .A(n6160), .ZN(U2947) );
  AOI21_X1 U7184 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6178), .A(n6162), .ZN(n6163) );
  OAI21_X1 U7185 ( .B1(n6164), .B2(n6180), .A(n6163), .ZN(U2948) );
  AOI21_X1 U7186 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6178), .A(n6165), .ZN(
        n6166) );
  OAI21_X1 U7187 ( .B1(n6167), .B2(n6180), .A(n6166), .ZN(U2949) );
  AOI21_X1 U7188 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6178), .A(n6168), .ZN(
        n6169) );
  OAI21_X1 U7189 ( .B1(n6170), .B2(n6180), .A(n6169), .ZN(U2950) );
  AOI21_X1 U7190 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6178), .A(n6171), .ZN(
        n6172) );
  OAI21_X1 U7191 ( .B1(n6173), .B2(n6180), .A(n6172), .ZN(U2952) );
  AOI21_X1 U7192 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6178), .A(n6174), .ZN(
        n6175) );
  OAI21_X1 U7193 ( .B1(n6176), .B2(n6180), .A(n6175), .ZN(U2953) );
  AOI22_X1 U7194 ( .A1(n6178), .A2(LWORD_REG_15__SCAN_IN), .B1(n6177), .B2(
        DATAI_15_), .ZN(n6179) );
  OAI21_X1 U7195 ( .B1(n6181), .B2(n6180), .A(n6179), .ZN(U2954) );
  AOI22_X1 U7196 ( .A1(n6238), .A2(REIP_REG_2__SCAN_IN), .B1(n6197), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6189) );
  XNOR2_X1 U7197 ( .A(n6182), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6184)
         );
  XNOR2_X1 U7198 ( .A(n6184), .B(n6183), .ZN(n6244) );
  AOI22_X1 U7199 ( .A1(n6187), .A2(n6186), .B1(n6185), .B2(n6244), .ZN(n6188)
         );
  OAI211_X1 U7200 ( .C1(n6191), .C2(n6190), .A(n6189), .B(n6188), .ZN(U2984)
         );
  OAI22_X1 U7201 ( .A1(n6194), .A2(n6193), .B1(n6192), .B2(n6552), .ZN(n6195)
         );
  INV_X1 U7202 ( .A(n6195), .ZN(n6199) );
  OAI21_X1 U7203 ( .B1(n6197), .B2(n6196), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6198) );
  OAI211_X1 U7204 ( .C1(n6201), .C2(n6200), .A(n6199), .B(n6198), .ZN(U2986)
         );
  AOI21_X1 U7205 ( .B1(n6203), .B2(n6240), .A(n6202), .ZN(n6207) );
  AOI22_X1 U7206 ( .A1(n6205), .A2(n6245), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6204), .ZN(n6206) );
  OAI211_X1 U7207 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6208), .A(n6207), .B(n6206), .ZN(U3007) );
  INV_X1 U7208 ( .A(n6209), .ZN(n6210) );
  AOI21_X1 U7209 ( .B1(n6211), .B2(n6240), .A(n6210), .ZN(n6215) );
  AOI22_X1 U7210 ( .A1(n6213), .A2(n6245), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6212), .ZN(n6214) );
  OAI211_X1 U7211 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6216), .A(n6215), 
        .B(n6214), .ZN(U3009) );
  INV_X1 U7212 ( .A(n6217), .ZN(n6221) );
  NAND2_X1 U7213 ( .A1(n6240), .A2(n6218), .ZN(n6220) );
  OAI211_X1 U7214 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6221), .A(n6220), 
        .B(n6219), .ZN(n6222) );
  AOI21_X1 U7215 ( .B1(n6223), .B2(n6245), .A(n6222), .ZN(n6224) );
  OAI21_X1 U7216 ( .B1(n6226), .B2(n6225), .A(n6224), .ZN(U3011) );
  NOR2_X1 U7217 ( .A1(n3628), .A2(n6227), .ZN(n6232) );
  INV_X1 U7218 ( .A(n6228), .ZN(n6230) );
  OAI21_X1 U7219 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6230), .A(n6229), 
        .ZN(n6231) );
  AOI211_X1 U7220 ( .C1(n6233), .C2(n6245), .A(n6232), .B(n6231), .ZN(n6234)
         );
  OAI21_X1 U7221 ( .B1(n6236), .B2(n6235), .A(n6234), .ZN(U3015) );
  INV_X1 U7222 ( .A(n6237), .ZN(n6239) );
  AOI22_X1 U7223 ( .A1(n6240), .A2(n6239), .B1(n6238), .B2(REIP_REG_2__SCAN_IN), .ZN(n6252) );
  OAI221_X1 U7224 ( .B1(n6243), .B2(n6242), .C1(n6243), .C2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6241), .ZN(n6251) );
  AOI22_X1 U7225 ( .A1(n6246), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6245), 
        .B2(n6244), .ZN(n6250) );
  NAND3_X1 U7226 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6248), .A3(n6247), 
        .ZN(n6249) );
  NAND4_X1 U7227 ( .A1(n6252), .A2(n6251), .A3(n6250), .A4(n6249), .ZN(U3016)
         );
  NOR2_X1 U7228 ( .A1(n6419), .A2(n6542), .ZN(U3019) );
  NAND2_X1 U7229 ( .A1(n6408), .A2(n6299), .ZN(n6261) );
  INV_X1 U7230 ( .A(n6261), .ZN(n6281) );
  NAND3_X1 U7231 ( .A1(n6254), .A2(n6536), .A3(n6290), .ZN(n6258) );
  NAND3_X1 U7232 ( .A1(n6256), .A2(n6255), .A3(n6544), .ZN(n6257) );
  NAND2_X1 U7233 ( .A1(n6258), .A2(n6257), .ZN(n6282) );
  AOI22_X1 U7234 ( .A1(n6336), .A2(n6281), .B1(n6349), .B2(n6282), .ZN(n6266)
         );
  NOR3_X1 U7235 ( .A1(n6283), .A2(n6329), .A3(n6343), .ZN(n6260) );
  OAI21_X1 U7236 ( .B1(n6260), .B2(n6538), .A(n6259), .ZN(n6264) );
  AOI21_X1 U7237 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6261), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6262) );
  NAND3_X1 U7238 ( .A1(n6264), .A2(n6263), .A3(n6262), .ZN(n6284) );
  AOI22_X1 U7239 ( .A1(n6284), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6292), 
        .B2(n6283), .ZN(n6265) );
  OAI211_X1 U7240 ( .C1(n6267), .C2(n6287), .A(n6266), .B(n6265), .ZN(U3068)
         );
  AOI22_X1 U7241 ( .A1(n6353), .A2(n6281), .B1(n6355), .B2(n6282), .ZN(n6269)
         );
  AOI22_X1 U7242 ( .A1(n6284), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6304), 
        .B2(n6283), .ZN(n6268) );
  OAI211_X1 U7243 ( .C1(n6576), .C2(n6287), .A(n6269), .B(n6268), .ZN(U3069)
         );
  AOI22_X1 U7244 ( .A1(n6360), .A2(n6282), .B1(n6358), .B2(n6281), .ZN(n6271)
         );
  AOI22_X1 U7245 ( .A1(n6284), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6359), 
        .B2(n6283), .ZN(n6270) );
  OAI211_X1 U7246 ( .C1(n6363), .C2(n6287), .A(n6271), .B(n6270), .ZN(U3070)
         );
  AOI22_X1 U7247 ( .A1(n6366), .A2(n6282), .B1(n6364), .B2(n6281), .ZN(n6273)
         );
  AOI22_X1 U7248 ( .A1(n6284), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6365), 
        .B2(n6283), .ZN(n6272) );
  OAI211_X1 U7249 ( .C1(n6369), .C2(n6287), .A(n6273), .B(n6272), .ZN(U3071)
         );
  AOI22_X1 U7250 ( .A1(n6372), .A2(n6282), .B1(n6370), .B2(n6281), .ZN(n6275)
         );
  AOI22_X1 U7251 ( .A1(n6284), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6371), 
        .B2(n6283), .ZN(n6274) );
  OAI211_X1 U7252 ( .C1(n6375), .C2(n6287), .A(n6275), .B(n6274), .ZN(U3072)
         );
  AOI22_X1 U7253 ( .A1(n6378), .A2(n6282), .B1(n6376), .B2(n6281), .ZN(n6277)
         );
  AOI22_X1 U7254 ( .A1(n6284), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6319), 
        .B2(n6283), .ZN(n6276) );
  OAI211_X1 U7255 ( .C1(n6278), .C2(n6287), .A(n6277), .B(n6276), .ZN(U3073)
         );
  AOI22_X1 U7256 ( .A1(n6385), .A2(n6282), .B1(n6382), .B2(n6281), .ZN(n6280)
         );
  AOI22_X1 U7257 ( .A1(n6284), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6383), 
        .B2(n6283), .ZN(n6279) );
  OAI211_X1 U7258 ( .C1(n6389), .C2(n6287), .A(n6280), .B(n6279), .ZN(U3074)
         );
  AOI22_X1 U7259 ( .A1(n6395), .A2(n6282), .B1(n6391), .B2(n6281), .ZN(n6286)
         );
  AOI22_X1 U7260 ( .A1(n6284), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6330), 
        .B2(n6283), .ZN(n6285) );
  OAI211_X1 U7261 ( .C1(n6288), .C2(n6287), .A(n6286), .B(n6285), .ZN(U3075)
         );
  AOI21_X1 U7262 ( .B1(n6290), .B2(n6289), .A(n6327), .ZN(n6295) );
  NOR2_X1 U7263 ( .A1(n6295), .A2(n6343), .ZN(n6291) );
  AOI21_X1 U7264 ( .B1(n6299), .B2(STATE2_REG_2__SCAN_IN), .A(n6291), .ZN(
        n6335) );
  AOI22_X1 U7265 ( .A1(n6327), .A2(n6336), .B1(n6292), .B2(n6329), .ZN(n6302)
         );
  INV_X1 U7266 ( .A(n6293), .ZN(n6338) );
  NOR2_X1 U7267 ( .A1(n6338), .A2(n6294), .ZN(n6534) );
  INV_X1 U7268 ( .A(n6534), .ZN(n6296) );
  NAND3_X1 U7269 ( .A1(n6296), .A2(n6536), .A3(n6295), .ZN(n6298) );
  OAI211_X1 U7270 ( .C1(n6299), .C2(n6536), .A(n6298), .B(n6297), .ZN(n6331)
         );
  AOI22_X1 U7271 ( .A1(n6331), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n6337), 
        .B2(n6328), .ZN(n6301) );
  OAI211_X1 U7272 ( .C1(n6335), .C2(n6303), .A(n6302), .B(n6301), .ZN(U3076)
         );
  AOI22_X1 U7273 ( .A1(n6329), .A2(n6304), .B1(n6327), .B2(n6353), .ZN(n6306)
         );
  AOI22_X1 U7274 ( .A1(n6331), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n6354), 
        .B2(n6328), .ZN(n6305) );
  OAI211_X1 U7275 ( .C1(n6335), .C2(n6577), .A(n6306), .B(n6305), .ZN(U3077)
         );
  AOI22_X1 U7276 ( .A1(n6329), .A2(n6359), .B1(n6327), .B2(n6358), .ZN(n6309)
         );
  AOI22_X1 U7277 ( .A1(n6331), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n6307), 
        .B2(n6328), .ZN(n6308) );
  OAI211_X1 U7278 ( .C1(n6335), .C2(n6310), .A(n6309), .B(n6308), .ZN(U3078)
         );
  AOI22_X1 U7279 ( .A1(n6328), .A2(n6311), .B1(n6364), .B2(n6327), .ZN(n6313)
         );
  AOI22_X1 U7280 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6331), .B1(n6365), 
        .B2(n6329), .ZN(n6312) );
  OAI211_X1 U7281 ( .C1(n6335), .C2(n6314), .A(n6313), .B(n6312), .ZN(U3079)
         );
  AOI22_X1 U7282 ( .A1(n6329), .A2(n6371), .B1(n6327), .B2(n6370), .ZN(n6317)
         );
  AOI22_X1 U7283 ( .A1(n6331), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n6315), 
        .B2(n6328), .ZN(n6316) );
  OAI211_X1 U7284 ( .C1(n6335), .C2(n6318), .A(n6317), .B(n6316), .ZN(U3080)
         );
  AOI22_X1 U7285 ( .A1(n6329), .A2(n6319), .B1(n6327), .B2(n6376), .ZN(n6321)
         );
  AOI22_X1 U7286 ( .A1(n6331), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n6377), 
        .B2(n6328), .ZN(n6320) );
  OAI211_X1 U7287 ( .C1(n6335), .C2(n6322), .A(n6321), .B(n6320), .ZN(U3081)
         );
  AOI22_X1 U7288 ( .A1(n6329), .A2(n6383), .B1(n6327), .B2(n6382), .ZN(n6325)
         );
  AOI22_X1 U7289 ( .A1(n6331), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n6323), 
        .B2(n6328), .ZN(n6324) );
  OAI211_X1 U7290 ( .C1(n6335), .C2(n6326), .A(n6325), .B(n6324), .ZN(U3082)
         );
  AOI22_X1 U7291 ( .A1(n6328), .A2(n6392), .B1(n6391), .B2(n6327), .ZN(n6333)
         );
  AOI22_X1 U7292 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6331), .B1(n6330), 
        .B2(n6329), .ZN(n6332) );
  OAI211_X1 U7293 ( .C1(n6335), .C2(n6334), .A(n6333), .B(n6332), .ZN(U3083)
         );
  INV_X1 U7294 ( .A(n6388), .ZN(n6393) );
  NOR2_X1 U7295 ( .A1(n6408), .A2(n6346), .ZN(n6390) );
  AOI22_X1 U7296 ( .A1(n6337), .A2(n6393), .B1(n6336), .B2(n6390), .ZN(n6351)
         );
  OAI21_X1 U7297 ( .B1(n6339), .B2(n6338), .A(n6536), .ZN(n6348) );
  AOI21_X1 U7298 ( .B1(n6341), .B2(n6340), .A(n6390), .ZN(n6347) );
  INV_X1 U7299 ( .A(n6347), .ZN(n6345) );
  AOI21_X1 U7300 ( .B1(n6343), .B2(n6346), .A(n6342), .ZN(n6344) );
  OAI21_X1 U7301 ( .B1(n6348), .B2(n6345), .A(n6344), .ZN(n6396) );
  OAI22_X1 U7302 ( .A1(n6348), .A2(n6347), .B1(n6346), .B2(n6560), .ZN(n6394)
         );
  AOI22_X1 U7303 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6396), .B1(n6349), 
        .B2(n6394), .ZN(n6350) );
  OAI211_X1 U7304 ( .C1(n6352), .C2(n6399), .A(n6351), .B(n6350), .ZN(U3108)
         );
  AOI22_X1 U7305 ( .A1(n6393), .A2(n6354), .B1(n6353), .B2(n6390), .ZN(n6357)
         );
  AOI22_X1 U7306 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6396), .B1(n6355), 
        .B2(n6394), .ZN(n6356) );
  OAI211_X1 U7307 ( .C1(n6572), .C2(n6399), .A(n6357), .B(n6356), .ZN(U3109)
         );
  INV_X1 U7308 ( .A(n6399), .ZN(n6384) );
  AOI22_X1 U7309 ( .A1(n6384), .A2(n6359), .B1(n6358), .B2(n6390), .ZN(n6362)
         );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6396), .B1(n6360), 
        .B2(n6394), .ZN(n6361) );
  OAI211_X1 U7311 ( .C1(n6363), .C2(n6388), .A(n6362), .B(n6361), .ZN(U3110)
         );
  AOI22_X1 U7312 ( .A1(n6384), .A2(n6365), .B1(n6364), .B2(n6390), .ZN(n6368)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6396), .B1(n6366), 
        .B2(n6394), .ZN(n6367) );
  OAI211_X1 U7314 ( .C1(n6369), .C2(n6388), .A(n6368), .B(n6367), .ZN(U3111)
         );
  AOI22_X1 U7315 ( .A1(n6384), .A2(n6371), .B1(n6370), .B2(n6390), .ZN(n6374)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6396), .B1(n6372), 
        .B2(n6394), .ZN(n6373) );
  OAI211_X1 U7317 ( .C1(n6375), .C2(n6388), .A(n6374), .B(n6373), .ZN(U3112)
         );
  AOI22_X1 U7318 ( .A1(n6393), .A2(n6377), .B1(n6376), .B2(n6390), .ZN(n6380)
         );
  AOI22_X1 U7319 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6396), .B1(n6378), 
        .B2(n6394), .ZN(n6379) );
  OAI211_X1 U7320 ( .C1(n6381), .C2(n6399), .A(n6380), .B(n6379), .ZN(U3113)
         );
  AOI22_X1 U7321 ( .A1(n6384), .A2(n6383), .B1(n6382), .B2(n6390), .ZN(n6387)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6396), .B1(n6385), 
        .B2(n6394), .ZN(n6386) );
  OAI211_X1 U7323 ( .C1(n6389), .C2(n6388), .A(n6387), .B(n6386), .ZN(U3114)
         );
  AOI22_X1 U7324 ( .A1(n6393), .A2(n6392), .B1(n6391), .B2(n6390), .ZN(n6398)
         );
  AOI22_X1 U7325 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6396), .B1(n6395), 
        .B2(n6394), .ZN(n6397) );
  OAI211_X1 U7326 ( .C1(n6400), .C2(n6399), .A(n6398), .B(n6397), .ZN(U3115)
         );
  OR2_X1 U7327 ( .A1(n6402), .A2(n6401), .ZN(n6406) );
  AOI21_X1 U7328 ( .B1(STATE2_REG_1__SCAN_IN), .B2(READY_N), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6403) );
  INV_X1 U7329 ( .A(n6403), .ZN(n6404) );
  AND2_X1 U7330 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6404), .ZN(n6405) );
  AND2_X1 U7331 ( .A1(n6406), .A2(n6405), .ZN(n6440) );
  OAI21_X1 U7332 ( .B1(n6407), .B2(n6434), .A(n6562), .ZN(n6439) );
  NOR3_X1 U7333 ( .A1(n6410), .A2(n6409), .A3(n6408), .ZN(n6414) );
  NAND2_X1 U7334 ( .A1(n6414), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6416) );
  INV_X1 U7335 ( .A(n6411), .ZN(n6413) );
  OAI22_X1 U7336 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6414), .B1(n6413), .B2(n6412), .ZN(n6415) );
  NAND2_X1 U7337 ( .A1(n6416), .A2(n6415), .ZN(n6417) );
  AOI222_X1 U7338 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6418), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6417), .C1(n6418), .C2(n6417), 
        .ZN(n6421) );
  AND2_X1 U7339 ( .A1(n6422), .A2(n6544), .ZN(n6420) );
  OAI221_X1 U7340 ( .B1(n6422), .B2(n6544), .C1(n6421), .C2(n6420), .A(n6419), 
        .ZN(n6431) );
  INV_X1 U7341 ( .A(n6423), .ZN(n6430) );
  INV_X1 U7342 ( .A(n6424), .ZN(n6425) );
  NOR2_X1 U7343 ( .A1(n6426), .A2(n6425), .ZN(n6429) );
  OAI21_X1 U7344 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6427), 
        .ZN(n6428) );
  NAND4_X1 U7345 ( .A1(n6431), .A2(n6430), .A3(n6429), .A4(n6428), .ZN(n6435)
         );
  INV_X1 U7346 ( .A(n6440), .ZN(n6432) );
  AOI221_X1 U7347 ( .B1(STATE2_REG_1__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(n6435), .C2(STATE2_REG_0__SCAN_IN), .A(n6432), .ZN(n6531) );
  AOI21_X1 U7348 ( .B1(READY_N), .B2(n6560), .A(n6531), .ZN(n6442) );
  NAND3_X1 U7349 ( .A1(n6442), .A2(n6434), .A3(n6433), .ZN(n6437) );
  AOI22_X1 U7350 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6437), .B1(n6436), .B2(
        n6435), .ZN(n6438) );
  OAI21_X1 U7351 ( .B1(n6440), .B2(n6439), .A(n6438), .ZN(U3148) );
  NOR3_X1 U7352 ( .A1(n6443), .A2(n6442), .A3(n6441), .ZN(n6447) );
  AOI221_X1 U7353 ( .B1(READY_N), .B2(n6445), .C1(n6444), .C2(n6445), .A(n6531), .ZN(n6446) );
  OR3_X1 U7354 ( .A1(n6448), .A2(n6447), .A3(n6446), .ZN(U3149) );
  OAI211_X1 U7355 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6462), .A(n6450), .B(
        n6449), .ZN(n6452) );
  INV_X1 U7356 ( .A(n6532), .ZN(n6451) );
  AOI21_X1 U7357 ( .B1(n6453), .B2(n6452), .A(n6451), .ZN(U3150) );
  INV_X1 U7358 ( .A(n6530), .ZN(n6527) );
  AND2_X1 U7359 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6527), .ZN(U3151) );
  AND2_X1 U7360 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6527), .ZN(U3152) );
  AND2_X1 U7361 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6527), .ZN(U3153) );
  AND2_X1 U7362 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6527), .ZN(U3154) );
  AND2_X1 U7363 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6527), .ZN(U3155) );
  AND2_X1 U7364 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6527), .ZN(U3156) );
  AND2_X1 U7365 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6527), .ZN(U3157) );
  AND2_X1 U7366 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6527), .ZN(U3158) );
  AND2_X1 U7367 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6527), .ZN(U3159) );
  AND2_X1 U7368 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6527), .ZN(U3160) );
  AND2_X1 U7369 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6527), .ZN(U3161) );
  AND2_X1 U7370 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6527), .ZN(U3162) );
  AND2_X1 U7371 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6527), .ZN(U3163) );
  AND2_X1 U7372 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6527), .ZN(U3164) );
  AND2_X1 U7373 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6527), .ZN(U3165) );
  AND2_X1 U7374 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6527), .ZN(U3166) );
  AND2_X1 U7375 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6527), .ZN(U3167) );
  AND2_X1 U7376 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6527), .ZN(U3168) );
  AND2_X1 U7377 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6527), .ZN(U3169) );
  AND2_X1 U7378 ( .A1(n6527), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U7379 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6527), .ZN(U3171) );
  AND2_X1 U7380 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6527), .ZN(U3172) );
  AND2_X1 U7381 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6527), .ZN(U3173) );
  AND2_X1 U7382 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6527), .ZN(U3174) );
  AND2_X1 U7383 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6527), .ZN(U3175) );
  AND2_X1 U7384 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6527), .ZN(U3176) );
  AND2_X1 U7385 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6527), .ZN(U3177) );
  AND2_X1 U7386 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6527), .ZN(U3178) );
  AND2_X1 U7387 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6527), .ZN(U3179) );
  AND2_X1 U7388 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6527), .ZN(U3180) );
  NAND2_X1 U7389 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6464) );
  OAI21_X1 U7390 ( .B1(n6463), .B2(n6462), .A(n6464), .ZN(n6468) );
  INV_X1 U7391 ( .A(n6468), .ZN(n6457) );
  AND2_X1 U7392 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6458) );
  INV_X1 U7393 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6568) );
  OAI21_X1 U7394 ( .B1(n6458), .B2(n6568), .A(n6556), .ZN(n6456) );
  INV_X1 U7395 ( .A(n6469), .ZN(n6454) );
  OAI211_X1 U7396 ( .C1(NA_N), .C2(n6455), .A(n3422), .B(n6454), .ZN(n6467) );
  OAI211_X1 U7397 ( .C1(n6469), .C2(n6457), .A(n6456), .B(n6467), .ZN(U3181)
         );
  NOR2_X1 U7398 ( .A1(n3422), .A2(n6568), .ZN(n6459) );
  OAI21_X1 U7399 ( .B1(n6459), .B2(n6458), .A(n6464), .ZN(n6460) );
  OAI211_X1 U7400 ( .C1(n6463), .C2(n6462), .A(n6461), .B(n6460), .ZN(U3182)
         );
  NOR2_X1 U7401 ( .A1(NA_N), .A2(n6462), .ZN(n6470) );
  OAI211_X1 U7402 ( .C1(n6470), .C2(n6463), .A(HOLD), .B(n6568), .ZN(n6465) );
  NAND3_X1 U7403 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6465), .A3(n6464), .ZN(
        n6466) );
  AOI22_X1 U7404 ( .A1(n6469), .A2(n6468), .B1(n6467), .B2(n6466), .ZN(n6472)
         );
  NAND4_X1 U7405 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .A3(
        REQUESTPENDING_REG_SCAN_IN), .A4(n6470), .ZN(n6471) );
  NAND2_X1 U7406 ( .A1(n6472), .A2(n6471), .ZN(U3183) );
  NAND2_X1 U7407 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6570), .ZN(n6521) );
  NOR2_X2 U7408 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6556), .ZN(n6518) );
  AOI22_X1 U7409 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6556), .ZN(n6473) );
  OAI21_X1 U7410 ( .B1(n6546), .B2(n6521), .A(n6473), .ZN(U3184) );
  INV_X1 U7411 ( .A(n6518), .ZN(n6525) );
  INV_X1 U7412 ( .A(n6521), .ZN(n6516) );
  AOI22_X1 U7413 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6516), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6556), .ZN(n6474) );
  OAI21_X1 U7414 ( .B1(n6475), .B2(n6525), .A(n6474), .ZN(U3185) );
  AOI22_X1 U7415 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6516), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6556), .ZN(n6476) );
  OAI21_X1 U7416 ( .B1(n6478), .B2(n6525), .A(n6476), .ZN(U3186) );
  AOI22_X1 U7417 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6556), .ZN(n6477) );
  OAI21_X1 U7418 ( .B1(n6478), .B2(n6521), .A(n6477), .ZN(U3187) );
  AOI22_X1 U7419 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6516), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6556), .ZN(n6479) );
  OAI21_X1 U7420 ( .B1(n6480), .B2(n6525), .A(n6479), .ZN(U3188) );
  AOI222_X1 U7421 ( .A1(n6516), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6556), .C1(REIP_REG_7__SCAN_IN), .C2(
        n6518), .ZN(n6481) );
  INV_X1 U7422 ( .A(n6481), .ZN(U3189) );
  AOI22_X1 U7423 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6516), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6556), .ZN(n6482) );
  OAI21_X1 U7424 ( .B1(n6484), .B2(n6525), .A(n6482), .ZN(U3190) );
  AOI22_X1 U7425 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6556), .ZN(n6483) );
  OAI21_X1 U7426 ( .B1(n6484), .B2(n6521), .A(n6483), .ZN(U3191) );
  AOI22_X1 U7427 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6556), .ZN(n6485) );
  OAI21_X1 U7428 ( .B1(n6486), .B2(n6521), .A(n6485), .ZN(U3192) );
  AOI22_X1 U7429 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6556), .ZN(n6487) );
  OAI21_X1 U7430 ( .B1(n6488), .B2(n6521), .A(n6487), .ZN(U3193) );
  INV_X1 U7431 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6490) );
  AOI22_X1 U7432 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6556), .ZN(n6489) );
  OAI21_X1 U7433 ( .B1(n6490), .B2(n6521), .A(n6489), .ZN(U3194) );
  AOI22_X1 U7434 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6516), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6556), .ZN(n6491) );
  OAI21_X1 U7435 ( .B1(n6492), .B2(n6525), .A(n6491), .ZN(U3195) );
  AOI22_X1 U7436 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6516), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6556), .ZN(n6493) );
  OAI21_X1 U7437 ( .B1(n6494), .B2(n6525), .A(n6493), .ZN(U3196) );
  AOI22_X1 U7438 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6516), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6556), .ZN(n6495) );
  OAI21_X1 U7439 ( .B1(n6497), .B2(n6525), .A(n6495), .ZN(U3197) );
  INV_X1 U7440 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6496) );
  OAI222_X1 U7441 ( .A1(n6521), .A2(n6497), .B1(n6496), .B2(n6570), .C1(n5608), 
        .C2(n6525), .ZN(U3198) );
  INV_X1 U7442 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6498) );
  INV_X1 U7443 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6681) );
  OAI222_X1 U7444 ( .A1(n6521), .A2(n5608), .B1(n6498), .B2(n6570), .C1(n6681), 
        .C2(n6525), .ZN(U3199) );
  AOI22_X1 U7445 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6556), .ZN(n6499) );
  OAI21_X1 U7446 ( .B1(n6681), .B2(n6521), .A(n6499), .ZN(U3200) );
  AOI22_X1 U7447 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6556), .ZN(n6500) );
  OAI21_X1 U7448 ( .B1(n5602), .B2(n6521), .A(n6500), .ZN(U3201) );
  AOI22_X1 U7449 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6556), .ZN(n6501) );
  OAI21_X1 U7450 ( .B1(n6502), .B2(n6521), .A(n6501), .ZN(U3202) );
  AOI22_X1 U7451 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6516), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6556), .ZN(n6503) );
  OAI21_X1 U7452 ( .B1(n6505), .B2(n6525), .A(n6503), .ZN(U3203) );
  AOI22_X1 U7453 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6556), .ZN(n6504) );
  OAI21_X1 U7454 ( .B1(n6505), .B2(n6521), .A(n6504), .ZN(U3204) );
  AOI22_X1 U7455 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6556), .ZN(n6506) );
  OAI21_X1 U7456 ( .B1(n6507), .B2(n6521), .A(n6506), .ZN(U3205) );
  AOI22_X1 U7457 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6556), .ZN(n6508) );
  OAI21_X1 U7458 ( .B1(n6648), .B2(n6521), .A(n6508), .ZN(U3206) );
  AOI22_X1 U7459 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6556), .ZN(n6509) );
  OAI21_X1 U7460 ( .B1(n6703), .B2(n6521), .A(n6509), .ZN(U3207) );
  INV_X1 U7461 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6510) );
  OAI222_X1 U7462 ( .A1(n6521), .A2(n6511), .B1(n6510), .B2(n6570), .C1(n6513), 
        .C2(n6525), .ZN(U3208) );
  AOI22_X1 U7463 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6556), .ZN(n6512) );
  OAI21_X1 U7464 ( .B1(n6513), .B2(n6521), .A(n6512), .ZN(U3209) );
  INV_X1 U7465 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6515) );
  OAI222_X1 U7466 ( .A1(n6521), .A2(n6628), .B1(n6515), .B2(n6570), .C1(n6514), 
        .C2(n6525), .ZN(U3210) );
  AOI22_X1 U7467 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6516), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6556), .ZN(n6517) );
  OAI21_X1 U7468 ( .B1(n6520), .B2(n6525), .A(n6517), .ZN(U3211) );
  AOI22_X1 U7469 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6518), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6556), .ZN(n6519) );
  OAI21_X1 U7470 ( .B1(n6520), .B2(n6521), .A(n6519), .ZN(U3212) );
  INV_X1 U7471 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6523) );
  OAI222_X1 U7472 ( .A1(n6525), .A2(n6524), .B1(n6523), .B2(n6570), .C1(n6522), 
        .C2(n6521), .ZN(U3213) );
  MUX2_X1 U7473 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6570), .Z(U3445) );
  MUX2_X1 U7474 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6570), .Z(U3446) );
  MUX2_X1 U7475 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6570), .Z(U3447) );
  MUX2_X1 U7476 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6570), .Z(U3448) );
  INV_X1 U7477 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6727) );
  INV_X1 U7478 ( .A(n6528), .ZN(n6526) );
  AOI21_X1 U7479 ( .B1(n6727), .B2(n6527), .A(n6526), .ZN(U3451) );
  OAI21_X1 U7480 ( .B1(n6530), .B2(n6529), .A(n6528), .ZN(U3452) );
  INV_X1 U7481 ( .A(n6531), .ZN(n6533) );
  OAI221_X1 U7482 ( .B1(n6718), .B2(STATE2_REG_0__SCAN_IN), .C1(n6718), .C2(
        n6533), .A(n6532), .ZN(U3453) );
  OR2_X1 U7483 ( .A1(n6535), .A2(n6534), .ZN(n6537) );
  AOI222_X1 U7484 ( .A1(n6541), .A2(n6540), .B1(n6539), .B2(n6538), .C1(n6537), 
        .C2(n6536), .ZN(n6543) );
  AOI22_X1 U7485 ( .A1(n6545), .A2(n6544), .B1(n6543), .B2(n6542), .ZN(U3462)
         );
  AOI21_X1 U7486 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6547) );
  AOI22_X1 U7487 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6547), .B2(n6546), .ZN(n6549) );
  INV_X1 U7488 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6548) );
  AOI22_X1 U7489 ( .A1(n6550), .A2(n6549), .B1(n6548), .B2(n6553), .ZN(U3468)
         );
  INV_X1 U7490 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6554) );
  NOR2_X1 U7491 ( .A1(n6553), .A2(REIP_REG_1__SCAN_IN), .ZN(n6551) );
  AOI22_X1 U7492 ( .A1(n6554), .A2(n6553), .B1(n6552), .B2(n6551), .ZN(U3469)
         );
  NAND2_X1 U7493 ( .A1(n6556), .A2(W_R_N_REG_SCAN_IN), .ZN(n6555) );
  OAI21_X1 U7494 ( .B1(n6556), .B2(READREQUEST_REG_SCAN_IN), .A(n6555), .ZN(
        U3470) );
  OAI211_X1 U7495 ( .C1(READY_N), .C2(n6559), .A(n6558), .B(n6557), .ZN(n6569)
         );
  AOI21_X1 U7496 ( .B1(n3179), .B2(n6561), .A(n6560), .ZN(n6563) );
  AOI21_X1 U7497 ( .B1(n6564), .B2(n6563), .A(n6562), .ZN(n6565) );
  OAI21_X1 U7498 ( .B1(n6566), .B2(n6565), .A(n6569), .ZN(n6567) );
  OAI21_X1 U7499 ( .B1(n6569), .B2(n6568), .A(n6567), .ZN(U3472) );
  MUX2_X1 U7500 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6570), .Z(U3473) );
  OAI22_X1 U7501 ( .A1(n6574), .A2(n6573), .B1(n6572), .B2(n6571), .ZN(n6580)
         );
  OAI22_X1 U7502 ( .A1(n6578), .A2(n6577), .B1(n6576), .B2(n6575), .ZN(n6579)
         );
  AOI211_X1 U7503 ( .C1(INSTQUEUE_REG_3__1__SCAN_IN), .C2(n6581), .A(n6580), 
        .B(n6579), .ZN(n6744) );
  NAND2_X1 U7504 ( .A1(keyinput50), .A2(keyinput57), .ZN(n6586) );
  NOR2_X1 U7505 ( .A1(keyinput36), .A2(keyinput23), .ZN(n6584) );
  INV_X1 U7506 ( .A(keyinput35), .ZN(n6582) );
  NOR4_X1 U7507 ( .A1(keyinput62), .A2(keyinput13), .A3(keyinput12), .A4(n6582), .ZN(n6583) );
  NAND4_X1 U7508 ( .A1(keyinput45), .A2(keyinput0), .A3(n6584), .A4(n6583), 
        .ZN(n6585) );
  NOR4_X1 U7509 ( .A1(keyinput18), .A2(keyinput25), .A3(n6586), .A4(n6585), 
        .ZN(n6588) );
  INV_X1 U7510 ( .A(keyinput46), .ZN(n6587) );
  NAND4_X1 U7511 ( .A1(keyinput24), .A2(keyinput2), .A3(n6588), .A4(n6587), 
        .ZN(n6609) );
  INV_X1 U7512 ( .A(keyinput10), .ZN(n6614) );
  INV_X1 U7513 ( .A(keyinput6), .ZN(n6617) );
  AND3_X1 U7514 ( .A1(n6614), .A2(n6617), .A3(keyinput11), .ZN(n6593) );
  NOR4_X1 U7515 ( .A1(keyinput44), .A2(keyinput48), .A3(keyinput15), .A4(
        keyinput29), .ZN(n6592) );
  NAND4_X1 U7516 ( .A1(keyinput63), .A2(keyinput19), .A3(keyinput47), .A4(
        keyinput26), .ZN(n6590) );
  NAND2_X1 U7517 ( .A1(keyinput33), .A2(keyinput61), .ZN(n6589) );
  NOR4_X1 U7518 ( .A1(keyinput52), .A2(keyinput7), .A3(n6590), .A4(n6589), 
        .ZN(n6591) );
  NAND4_X1 U7519 ( .A1(keyinput16), .A2(n6593), .A3(n6592), .A4(n6591), .ZN(
        n6608) );
  NOR2_X1 U7520 ( .A1(keyinput60), .A2(keyinput14), .ZN(n6599) );
  NAND2_X1 U7521 ( .A1(keyinput38), .A2(keyinput28), .ZN(n6597) );
  NOR3_X1 U7522 ( .A1(keyinput54), .A2(keyinput4), .A3(keyinput53), .ZN(n6595)
         );
  NOR3_X1 U7523 ( .A1(keyinput41), .A2(keyinput43), .A3(keyinput58), .ZN(n6594) );
  NAND4_X1 U7524 ( .A1(keyinput59), .A2(n6595), .A3(keyinput27), .A4(n6594), 
        .ZN(n6596) );
  NOR4_X1 U7525 ( .A1(keyinput49), .A2(keyinput1), .A3(n6597), .A4(n6596), 
        .ZN(n6598) );
  NAND4_X1 U7526 ( .A1(keyinput21), .A2(keyinput31), .A3(n6599), .A4(n6598), 
        .ZN(n6607) );
  NAND2_X1 U7527 ( .A1(keyinput17), .A2(keyinput3), .ZN(n6600) );
  NOR3_X1 U7528 ( .A1(keyinput5), .A2(keyinput56), .A3(n6600), .ZN(n6605) );
  NOR3_X1 U7529 ( .A1(keyinput22), .A2(keyinput37), .A3(keyinput9), .ZN(n6604)
         );
  NAND4_X1 U7530 ( .A1(keyinput34), .A2(keyinput40), .A3(keyinput8), .A4(
        keyinput32), .ZN(n6602) );
  NAND2_X1 U7531 ( .A1(keyinput30), .A2(keyinput20), .ZN(n6601) );
  NOR4_X1 U7532 ( .A1(keyinput51), .A2(keyinput42), .A3(n6602), .A4(n6601), 
        .ZN(n6603) );
  NAND4_X1 U7533 ( .A1(n6605), .A2(keyinput55), .A3(n6604), .A4(n6603), .ZN(
        n6606) );
  NOR4_X1 U7534 ( .A1(n6609), .A2(n6608), .A3(n6607), .A4(n6606), .ZN(n6741)
         );
  INV_X1 U7535 ( .A(keyinput19), .ZN(n6611) );
  AOI22_X1 U7536 ( .A1(n6612), .A2(keyinput47), .B1(ADDRESS_REG_14__SCAN_IN), 
        .B2(n6611), .ZN(n6610) );
  OAI221_X1 U7537 ( .B1(n6612), .B2(keyinput47), .C1(n6611), .C2(
        ADDRESS_REG_14__SCAN_IN), .A(n6610), .ZN(n6625) );
  INV_X1 U7538 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6615) );
  AOI22_X1 U7539 ( .A1(n6615), .A2(keyinput26), .B1(ADDRESS_REG_5__SCAN_IN), 
        .B2(n6614), .ZN(n6613) );
  OAI221_X1 U7540 ( .B1(n6615), .B2(keyinput26), .C1(n6614), .C2(
        ADDRESS_REG_5__SCAN_IN), .A(n6613), .ZN(n6624) );
  INV_X1 U7541 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6618) );
  AOI22_X1 U7542 ( .A1(n6618), .A2(keyinput16), .B1(DATAO_REG_6__SCAN_IN), 
        .B2(n6617), .ZN(n6616) );
  OAI221_X1 U7543 ( .B1(n6618), .B2(keyinput16), .C1(n6617), .C2(
        DATAO_REG_6__SCAN_IN), .A(n6616), .ZN(n6623) );
  INV_X1 U7544 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U7545 ( .A1(n6621), .A2(keyinput11), .B1(n6620), .B2(keyinput33), 
        .ZN(n6619) );
  OAI221_X1 U7546 ( .B1(n6621), .B2(keyinput11), .C1(n6620), .C2(keyinput33), 
        .A(n6619), .ZN(n6622) );
  NOR4_X1 U7547 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6739)
         );
  INV_X1 U7548 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U7549 ( .A1(n6628), .A2(keyinput7), .B1(n6627), .B2(keyinput52), 
        .ZN(n6626) );
  OAI221_X1 U7550 ( .B1(n6628), .B2(keyinput7), .C1(n6627), .C2(keyinput52), 
        .A(n6626), .ZN(n6639) );
  INV_X1 U7551 ( .A(keyinput61), .ZN(n6630) );
  AOI22_X1 U7552 ( .A1(n6631), .A2(keyinput44), .B1(DATAO_REG_20__SCAN_IN), 
        .B2(n6630), .ZN(n6629) );
  OAI221_X1 U7553 ( .B1(n6631), .B2(keyinput44), .C1(n6630), .C2(
        DATAO_REG_20__SCAN_IN), .A(n6629), .ZN(n6638) );
  AOI22_X1 U7554 ( .A1(n4590), .A2(keyinput48), .B1(keyinput15), .B2(n6633), 
        .ZN(n6632) );
  OAI221_X1 U7555 ( .B1(n4590), .B2(keyinput48), .C1(n6633), .C2(keyinput15), 
        .A(n6632), .ZN(n6637) );
  INV_X1 U7556 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6635) );
  AOI22_X1 U7557 ( .A1(n5358), .A2(keyinput29), .B1(n6635), .B2(keyinput54), 
        .ZN(n6634) );
  OAI221_X1 U7558 ( .B1(n5358), .B2(keyinput29), .C1(n6635), .C2(keyinput54), 
        .A(n6634), .ZN(n6636) );
  NOR4_X1 U7559 ( .A1(n6639), .A2(n6638), .A3(n6637), .A4(n6636), .ZN(n6738)
         );
  INV_X1 U7560 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U7561 ( .A1(n6642), .A2(keyinput46), .B1(n6641), .B2(keyinput50), 
        .ZN(n6640) );
  OAI221_X1 U7562 ( .B1(n6642), .B2(keyinput46), .C1(n6641), .C2(keyinput50), 
        .A(n6640), .ZN(n6669) );
  INV_X1 U7563 ( .A(keyinput25), .ZN(n6644) );
  AOI22_X1 U7564 ( .A1(n6645), .A2(keyinput18), .B1(LWORD_REG_14__SCAN_IN), 
        .B2(n6644), .ZN(n6643) );
  OAI221_X1 U7565 ( .B1(n6645), .B2(keyinput18), .C1(n6644), .C2(
        LWORD_REG_14__SCAN_IN), .A(n6643), .ZN(n6668) );
  INV_X1 U7566 ( .A(DATAI_15_), .ZN(n6647) );
  OAI22_X1 U7567 ( .A1(n6648), .A2(keyinput57), .B1(n6647), .B2(keyinput36), 
        .ZN(n6646) );
  AOI221_X1 U7568 ( .B1(n6648), .B2(keyinput57), .C1(keyinput36), .C2(n6647), 
        .A(n6646), .ZN(n6650) );
  XNOR2_X1 U7569 ( .A(keyinput24), .B(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6649)
         );
  OAI211_X1 U7570 ( .C1(keyinput39), .C2(n6742), .A(n6650), .B(n6649), .ZN(
        n6667) );
  INV_X1 U7571 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6653) );
  INV_X1 U7572 ( .A(keyinput23), .ZN(n6652) );
  OAI22_X1 U7573 ( .A1(n6653), .A2(keyinput45), .B1(n6652), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n6651) );
  AOI221_X1 U7574 ( .B1(n6653), .B2(keyinput45), .C1(DATAO_REG_22__SCAN_IN), 
        .C2(n6652), .A(n6651), .ZN(n6665) );
  INV_X1 U7575 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6656) );
  INV_X1 U7576 ( .A(keyinput0), .ZN(n6655) );
  OAI22_X1 U7577 ( .A1(n6656), .A2(keyinput62), .B1(n6655), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n6654) );
  AOI221_X1 U7578 ( .B1(n6656), .B2(keyinput62), .C1(DATAO_REG_29__SCAN_IN), 
        .C2(n6655), .A(n6654), .ZN(n6664) );
  INV_X1 U7579 ( .A(keyinput13), .ZN(n6658) );
  OAI22_X1 U7580 ( .A1(keyinput35), .A2(n6659), .B1(n6658), .B2(
        ADDRESS_REG_26__SCAN_IN), .ZN(n6657) );
  AOI221_X1 U7581 ( .B1(n6659), .B2(keyinput35), .C1(n6658), .C2(
        ADDRESS_REG_26__SCAN_IN), .A(n6657), .ZN(n6663) );
  INV_X1 U7582 ( .A(keyinput63), .ZN(n6661) );
  OAI22_X1 U7583 ( .A1(n5473), .A2(keyinput12), .B1(n6661), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n6660) );
  AOI221_X1 U7584 ( .B1(n5473), .B2(keyinput12), .C1(UWORD_REG_6__SCAN_IN), 
        .C2(n6661), .A(n6660), .ZN(n6662) );
  NAND4_X1 U7585 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6666)
         );
  NOR4_X1 U7586 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6737)
         );
  INV_X1 U7587 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6672) );
  OAI22_X1 U7588 ( .A1(n6672), .A2(keyinput43), .B1(n6671), .B2(keyinput58), 
        .ZN(n6670) );
  AOI221_X1 U7589 ( .B1(n6672), .B2(keyinput43), .C1(keyinput58), .C2(n6671), 
        .A(n6670), .ZN(n6685) );
  INV_X1 U7590 ( .A(keyinput49), .ZN(n6674) );
  OAI22_X1 U7591 ( .A1(keyinput27), .A2(n6675), .B1(n6674), .B2(
        MEMORYFETCH_REG_SCAN_IN), .ZN(n6673) );
  AOI221_X1 U7592 ( .B1(n6675), .B2(keyinput27), .C1(n6674), .C2(
        MEMORYFETCH_REG_SCAN_IN), .A(n6673), .ZN(n6684) );
  INV_X1 U7593 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6678) );
  INV_X1 U7594 ( .A(keyinput28), .ZN(n6677) );
  OAI22_X1 U7595 ( .A1(n6678), .A2(keyinput17), .B1(n6677), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n6676) );
  AOI221_X1 U7596 ( .B1(n6678), .B2(keyinput17), .C1(DATAO_REG_28__SCAN_IN), 
        .C2(n6677), .A(n6676), .ZN(n6683) );
  INV_X1 U7597 ( .A(keyinput1), .ZN(n6680) );
  OAI22_X1 U7598 ( .A1(n6681), .A2(keyinput38), .B1(n6680), .B2(
        ADDRESS_REG_29__SCAN_IN), .ZN(n6679) );
  AOI221_X1 U7599 ( .B1(n6681), .B2(keyinput38), .C1(ADDRESS_REG_29__SCAN_IN), 
        .C2(n6680), .A(n6679), .ZN(n6682) );
  NAND4_X1 U7600 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .ZN(n6735)
         );
  INV_X1 U7601 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6688) );
  INV_X1 U7602 ( .A(keyinput4), .ZN(n6687) );
  OAI22_X1 U7603 ( .A1(n6688), .A2(keyinput21), .B1(n6687), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6686) );
  AOI221_X1 U7604 ( .B1(n6688), .B2(keyinput21), .C1(UWORD_REG_12__SCAN_IN), 
        .C2(n6687), .A(n6686), .ZN(n6700) );
  INV_X1 U7605 ( .A(keyinput59), .ZN(n6690) );
  OAI22_X1 U7606 ( .A1(n6691), .A2(keyinput53), .B1(n6690), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6689) );
  AOI221_X1 U7607 ( .B1(n6691), .B2(keyinput53), .C1(DATAO_REG_15__SCAN_IN), 
        .C2(n6690), .A(n6689), .ZN(n6699) );
  INV_X1 U7608 ( .A(keyinput41), .ZN(n6693) );
  OAI22_X1 U7609 ( .A1(n6694), .A2(keyinput14), .B1(n6693), .B2(
        D_C_N_REG_SCAN_IN), .ZN(n6692) );
  AOI221_X1 U7610 ( .B1(n6694), .B2(keyinput14), .C1(D_C_N_REG_SCAN_IN), .C2(
        n6693), .A(n6692), .ZN(n6698) );
  INV_X1 U7611 ( .A(keyinput60), .ZN(n6696) );
  OAI22_X1 U7612 ( .A1(n4981), .A2(keyinput31), .B1(n6696), .B2(
        ADDRESS_REG_24__SCAN_IN), .ZN(n6695) );
  AOI221_X1 U7613 ( .B1(n4981), .B2(keyinput31), .C1(ADDRESS_REG_24__SCAN_IN), 
        .C2(n6696), .A(n6695), .ZN(n6697) );
  NAND4_X1 U7614 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n6734)
         );
  INV_X1 U7615 ( .A(keyinput42), .ZN(n6702) );
  OAI22_X1 U7616 ( .A1(n6703), .A2(keyinput9), .B1(n6702), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6701) );
  AOI221_X1 U7617 ( .B1(n6703), .B2(keyinput9), .C1(DATAO_REG_13__SCAN_IN), 
        .C2(n6702), .A(n6701), .ZN(n6715) );
  OAI22_X1 U7618 ( .A1(n6705), .A2(keyinput37), .B1(n4482), .B2(keyinput55), 
        .ZN(n6704) );
  AOI221_X1 U7619 ( .B1(n6705), .B2(keyinput37), .C1(keyinput55), .C2(n4482), 
        .A(n6704), .ZN(n6714) );
  OAI22_X1 U7620 ( .A1(n6708), .A2(keyinput2), .B1(n6707), .B2(keyinput20), 
        .ZN(n6706) );
  AOI221_X1 U7621 ( .B1(n6708), .B2(keyinput2), .C1(keyinput20), .C2(n6707), 
        .A(n6706), .ZN(n6713) );
  INV_X1 U7622 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6710) );
  OAI22_X1 U7623 ( .A1(n6711), .A2(keyinput30), .B1(n6710), .B2(keyinput51), 
        .ZN(n6709) );
  AOI221_X1 U7624 ( .B1(n6711), .B2(keyinput30), .C1(keyinput51), .C2(n6710), 
        .A(n6709), .ZN(n6712) );
  NAND4_X1 U7625 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6733)
         );
  INV_X1 U7626 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6717) );
  OAI22_X1 U7627 ( .A1(n6718), .A2(keyinput56), .B1(n6717), .B2(keyinput34), 
        .ZN(n6716) );
  AOI221_X1 U7628 ( .B1(n6718), .B2(keyinput56), .C1(keyinput34), .C2(n6717), 
        .A(n6716), .ZN(n6731) );
  INV_X1 U7629 ( .A(keyinput5), .ZN(n6720) );
  OAI22_X1 U7630 ( .A1(n6721), .A2(keyinput3), .B1(n6720), .B2(
        CODEFETCH_REG_SCAN_IN), .ZN(n6719) );
  AOI221_X1 U7631 ( .B1(n6721), .B2(keyinput3), .C1(CODEFETCH_REG_SCAN_IN), 
        .C2(n6720), .A(n6719), .ZN(n6730) );
  INV_X1 U7632 ( .A(keyinput22), .ZN(n6723) );
  OAI22_X1 U7633 ( .A1(keyinput8), .A2(n6724), .B1(n6723), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n6722) );
  AOI221_X1 U7634 ( .B1(n6724), .B2(keyinput8), .C1(n6723), .C2(
        DATAO_REG_17__SCAN_IN), .A(n6722), .ZN(n6729) );
  INV_X1 U7635 ( .A(keyinput32), .ZN(n6726) );
  OAI22_X1 U7636 ( .A1(keyinput40), .A2(n6727), .B1(n6726), .B2(
        ADDRESS_REG_15__SCAN_IN), .ZN(n6725) );
  AOI221_X1 U7637 ( .B1(n6727), .B2(keyinput40), .C1(n6726), .C2(
        ADDRESS_REG_15__SCAN_IN), .A(n6725), .ZN(n6728) );
  NAND4_X1 U7638 ( .A1(n6731), .A2(n6730), .A3(n6729), .A4(n6728), .ZN(n6732)
         );
  NOR4_X1 U7639 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n6736)
         );
  NAND4_X1 U7640 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6740)
         );
  AOI221_X1 U7641 ( .B1(keyinput39), .B2(n6742), .C1(n6741), .C2(n6742), .A(
        n6740), .ZN(n6743) );
  XNOR2_X1 U7642 ( .A(n6744), .B(n6743), .ZN(U3045) );
  AND2_X1 U3736 ( .A1(n4291), .A2(n4377), .ZN(n3253) );
  NAND2_X1 U3919 ( .A1(n3189), .A2(n3681), .ZN(n4321) );
  CLKBUF_X2 U34520 ( .A(n3253), .Z(n4150) );
  XNOR2_X1 U34710 ( .A(n3307), .B(n6235), .ZN(n5369) );
  CLKBUF_X1 U3686 ( .A(n6102), .Z(n6100) );
endmodule

