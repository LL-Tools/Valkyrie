

module b15_C_SARLock_k_64_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2953, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545;

  INV_X2 U3402 ( .A(n5692), .ZN(n5702) );
  INV_X1 U3403 ( .A(n5386), .ZN(n5340) );
  CLKBUF_X2 U3404 ( .A(n3981), .Z(n4869) );
  CLKBUF_X2 U3405 ( .A(n3283), .Z(n4636) );
  CLKBUF_X2 U3407 ( .A(n3078), .Z(n3672) );
  CLKBUF_X2 U3408 ( .A(n3237), .Z(n4140) );
  CLKBUF_X2 U3409 ( .A(n3119), .Z(n3281) );
  CLKBUF_X2 U3410 ( .A(n3066), .Z(n4125) );
  CLKBUF_X2 U3411 ( .A(n3199), .Z(n3844) );
  CLKBUF_X2 U3412 ( .A(n4637), .Z(n4120) );
  CLKBUF_X2 U3413 ( .A(n3103), .Z(n4635) );
  INV_X1 U3414 ( .A(n3175), .ZN(n5684) );
  AND4_X1 U3415 ( .A1(n3102), .A2(n3101), .A3(n3100), .A4(n3099), .ZN(n3109)
         );
  AND2_X1 U3417 ( .A1(n4183), .A2(n4268), .ZN(n3103) );
  AND2_X2 U3418 ( .A1(n3029), .A2(n4184), .ZN(n3117) );
  NOR2_X1 U3419 ( .A1(n3158), .A2(n4072), .ZN(n3183) );
  CLKBUF_X2 U3420 ( .A(n3282), .Z(n3912) );
  NOR2_X1 U3421 ( .A1(n3181), .A2(n3180), .ZN(n4082) );
  AND4_X1 U3422 ( .A1(n3107), .A2(n3106), .A3(n3105), .A4(n3104), .ZN(n3108)
         );
  INV_X1 U3423 ( .A(n4438), .ZN(n3983) );
  NAND2_X1 U3424 ( .A1(n3982), .A2(n2957), .ZN(n4027) );
  AND2_X1 U3425 ( .A1(n4220), .A2(n3989), .ZN(n4246) );
  INV_X2 U3426 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3023) );
  OR3_X2 U3427 ( .A1(n4868), .A2(n4038), .A3(n4037), .ZN(n2974) );
  AND2_X2 U3428 ( .A1(n3159), .A2(n3160), .ZN(n6364) );
  AND2_X1 U3429 ( .A1(n4457), .A2(n4456), .ZN(n4453) );
  OAI21_X1 U3431 ( .B1(n4975), .B2(n5027), .A(n5203), .ZN(n3436) );
  OAI22_X2 U3432 ( .A1(n4946), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n4957), .B2(n4939), .ZN(n4940) );
  NAND2_X2 U3433 ( .A1(n4965), .A2(n4966), .ZN(n4964) );
  AND2_X1 U3434 ( .A1(n4184), .A2(n4269), .ZN(n2953) );
  AND2_X1 U3435 ( .A1(n4184), .A2(n4269), .ZN(n3283) );
  INV_X1 U3437 ( .A(n2956), .ZN(n2955) );
  NAND4_X4 U3438 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n3159)
         );
  AND2_X4 U3439 ( .A1(n3030), .A2(n4269), .ZN(n3077) );
  AND2_X2 U3440 ( .A1(n3024), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3030)
         );
  OAI21_X1 U3441 ( .B1(n4935), .B2(n3437), .A(n3436), .ZN(n3440) );
  NAND2_X1 U3442 ( .A1(n4372), .A2(n3400), .ZN(n4405) );
  AND2_X1 U3443 ( .A1(n4360), .A2(n4411), .ZN(n4392) );
  BUF_X2 U3444 ( .A(n3156), .Z(n4092) );
  AND2_X2 U34450 ( .A1(n3156), .A2(n3155), .ZN(n3444) );
  BUF_X2 U34460 ( .A(n3117), .Z(n4272) );
  BUF_X2 U34470 ( .A(n3118), .Z(n4147) );
  INV_X2 U34480 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n3558) );
  NOR2_X4 U3449 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4268) );
  XNOR2_X1 U3450 ( .A(n2999), .B(n5002), .ZN(n4996) );
  NOR2_X1 U34510 ( .A1(n4111), .A2(n5002), .ZN(n4677) );
  AOI22_X1 U34520 ( .A1(n4912), .A2(n4911), .B1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5026), .ZN(n4913) );
  OR2_X1 U34530 ( .A1(n4900), .A2(n5692), .ZN(n4161) );
  NAND2_X1 U3454 ( .A1(n3937), .A2(n5003), .ZN(n4111) );
  AND2_X1 U34550 ( .A1(n3943), .A2(n3942), .ZN(n3944) );
  AND2_X1 U34560 ( .A1(n3934), .A2(n3933), .ZN(n3935) );
  OR2_X1 U3457 ( .A1(n4906), .A2(n5692), .ZN(n3934) );
  CLKBUF_X1 U3458 ( .A(n3938), .Z(n3939) );
  NAND2_X1 U34590 ( .A1(n3938), .A2(n3439), .ZN(n4676) );
  OAI21_X1 U34600 ( .B1(n3923), .B2(n3924), .A(n4136), .ZN(n4906) );
  AND2_X1 U34610 ( .A1(n4936), .A2(n4935), .ZN(n4971) );
  NAND2_X1 U34620 ( .A1(n3440), .A2(n4931), .ZN(n3938) );
  CLKBUF_X1 U34630 ( .A(n4624), .Z(n2964) );
  AOI21_X1 U34640 ( .B1(n4692), .B2(n4691), .A(n4690), .ZN(n4693) );
  NAND2_X1 U34650 ( .A1(n4687), .A2(n4686), .ZN(n4823) );
  XNOR2_X1 U3466 ( .A(n2987), .B(n4071), .ZN(n4820) );
  NAND2_X1 U3467 ( .A1(n4558), .A2(n4559), .ZN(n5512) );
  AND2_X2 U34680 ( .A1(n4681), .A2(n4740), .ZN(n4685) );
  NAND2_X1 U34690 ( .A1(n2995), .A2(n2996), .ZN(n4558) );
  NAND2_X1 U34700 ( .A1(n4468), .A2(n2972), .ZN(n2995) );
  NAND2_X1 U34710 ( .A1(n4403), .A2(n3413), .ZN(n4468) );
  NAND2_X1 U34720 ( .A1(n3518), .A2(n3517), .ZN(n4361) );
  NOR2_X2 U34730 ( .A1(n4317), .A2(n4318), .ZN(n4360) );
  XNOR2_X1 U34740 ( .A(n3364), .B(n3372), .ZN(n3513) );
  XNOR2_X1 U3475 ( .A(n3351), .B(n3373), .ZN(n2989) );
  NAND2_X1 U3476 ( .A1(n3331), .A2(n4338), .ZN(n3351) );
  NAND2_X1 U3477 ( .A1(n3325), .A2(n3324), .ZN(n5538) );
  NAND2_X1 U3478 ( .A1(n3266), .A2(n3022), .ZN(n3297) );
  OAI21_X1 U3479 ( .B1(n5855), .B2(STATE2_REG_0__SCAN_IN), .A(n3225), .ZN(
        n3307) );
  NAND2_X1 U3480 ( .A1(n4362), .A2(n4363), .ZN(n4376) );
  INV_X1 U3481 ( .A(n4320), .ZN(n4362) );
  NAND2_X1 U3482 ( .A1(n4246), .A2(n4247), .ZN(n4336) );
  AOI21_X1 U3483 ( .B1(n3268), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3193), 
        .ZN(n3194) );
  NAND2_X1 U3484 ( .A1(n3186), .A2(n3185), .ZN(n3538) );
  NAND2_X1 U3485 ( .A1(n3260), .A2(n3259), .ZN(n3305) );
  MUX2_X1 U3486 ( .A(n3317), .B(n3316), .S(n3315), .Z(n6344) );
  NAND2_X1 U3487 ( .A1(n3986), .A2(n3985), .ZN(n3989) );
  AND2_X1 U3488 ( .A1(n3182), .A2(n4082), .ZN(n3186) );
  OAI211_X1 U3489 ( .C1(n3484), .C2(n3264), .A(n3263), .B(n3262), .ZN(n3304)
         );
  NOR2_X1 U3490 ( .A1(n3317), .A2(n3254), .ZN(n3316) );
  NOR2_X1 U3491 ( .A1(n3151), .A2(n3502), .ZN(n3162) );
  AOI22_X1 U3492 ( .A1(n3445), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3261), 
        .B2(n3300), .ZN(n3210) );
  INV_X1 U3493 ( .A(n3484), .ZN(n3445) );
  AOI22_X1 U3494 ( .A1(n3183), .A2(n3175), .B1(n6364), .B2(n3161), .ZN(n3179)
         );
  AND2_X1 U3495 ( .A1(n4438), .A2(n4869), .ZN(n4057) );
  INV_X1 U3496 ( .A(n4438), .ZN(n2957) );
  AND2_X1 U3497 ( .A1(n3250), .A2(n3408), .ZN(n3414) );
  INV_X1 U3498 ( .A(n3981), .ZN(n4785) );
  NAND2_X1 U3499 ( .A1(n3131), .A2(n3157), .ZN(n3128) );
  OR2_X1 U3500 ( .A1(n3248), .A2(n3247), .ZN(n3319) );
  NAND2_X1 U3501 ( .A1(n3131), .A2(n3155), .ZN(n3148) );
  OR2_X1 U3502 ( .A1(n3236), .A2(n3235), .ZN(n3408) );
  CLKBUF_X1 U3504 ( .A(n3135), .Z(n3505) );
  INV_X1 U3505 ( .A(n3156), .ZN(n3160) );
  AND4_X1 U3506 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3111)
         );
  NAND2_X1 U3507 ( .A1(n2973), .A2(n2970), .ZN(n3156) );
  AND2_X1 U3508 ( .A1(n3076), .A2(n3075), .ZN(n3157) );
  AND4_X1 U3509 ( .A1(n3050), .A2(n3049), .A3(n3048), .A4(n3047), .ZN(n3016)
         );
  AND4_X1 U3510 ( .A1(n3083), .A2(n3082), .A3(n3081), .A4(n3080), .ZN(n3089)
         );
  AND4_X1 U3511 ( .A1(n3070), .A2(n3069), .A3(n3068), .A4(n3067), .ZN(n3076)
         );
  AND4_X1 U3512 ( .A1(n3074), .A2(n3073), .A3(n3072), .A4(n3071), .ZN(n3075)
         );
  AND4_X1 U3513 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3110)
         );
  BUF_X2 U3514 ( .A(n3077), .Z(n4146) );
  BUF_X2 U3515 ( .A(n3197), .Z(n4145) );
  AND2_X2 U3516 ( .A1(n3029), .A2(n4183), .ZN(n2968) );
  AND2_X2 U3517 ( .A1(n4178), .A2(n3031), .ZN(n4637) );
  AND2_X2 U3518 ( .A1(n3032), .A2(n4273), .ZN(n3198) );
  AND2_X2 U3519 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n3023), .ZN(n3029)
         );
  AND2_X1 U3520 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4273) );
  INV_X2 U3521 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6366) );
  NOR2_X1 U3522 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4419) );
  NAND2_X1 U3523 ( .A1(n2988), .A2(n2981), .ZN(n4842) );
  OR2_X2 U3524 ( .A1(n3195), .A2(n3194), .ZN(n2958) );
  CLKBUF_X1 U3525 ( .A(n3654), .Z(n2959) );
  AND2_X1 U3526 ( .A1(n3003), .A2(n3667), .ZN(n2960) );
  INV_X1 U3527 ( .A(n3132), .ZN(n2961) );
  OR2_X1 U3528 ( .A1(n3195), .A2(n3194), .ZN(n3267) );
  OR2_X2 U3529 ( .A1(n3065), .A2(n3064), .ZN(n3153) );
  OAI21_X1 U3530 ( .B1(n4745), .B2(n4682), .A(n4679), .ZN(n2987) );
  AND2_X4 U3531 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4184) );
  OR2_X1 U3532 ( .A1(n3168), .A2(n3024), .ZN(n3539) );
  NAND2_X2 U3533 ( .A1(n3923), .A2(n3924), .ZN(n4136) );
  NAND2_X1 U3534 ( .A1(n3187), .A2(n3538), .ZN(n2962) );
  NOR2_X1 U3535 ( .A1(n4111), .A2(n5002), .ZN(n2963) );
  NAND2_X1 U3536 ( .A1(n2958), .A2(n3196), .ZN(n2965) );
  NAND2_X1 U3537 ( .A1(n3187), .A2(n3538), .ZN(n3212) );
  NAND2_X1 U3538 ( .A1(n3267), .A2(n3196), .ZN(n4282) );
  INV_X2 U3539 ( .A(n3155), .ZN(n3146) );
  NAND2_X4 U3540 ( .A1(n3016), .A2(n3055), .ZN(n3155) );
  NOR2_X1 U3541 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3032) );
  AND2_X1 U3542 ( .A1(n3032), .A2(n4273), .ZN(n2966) );
  NAND2_X2 U3543 ( .A1(n3451), .A2(n3128), .ZN(n3170) );
  AND2_X4 U3544 ( .A1(n3030), .A2(n4268), .ZN(n3118) );
  AND2_X2 U3545 ( .A1(n3134), .A2(n3133), .ZN(n3017) );
  XNOR2_X1 U3546 ( .A(n3328), .B(n5628), .ZN(n4324) );
  NAND2_X1 U3547 ( .A1(n3296), .A2(n3295), .ZN(n3328) );
  XNOR2_X1 U3548 ( .A(n2962), .B(n3214), .ZN(n5855) );
  NAND2_X2 U3549 ( .A1(n3948), .A2(n3160), .ZN(n3970) );
  INV_X2 U3550 ( .A(n3135), .ZN(n3131) );
  NAND2_X2 U3551 ( .A1(n3089), .A2(n3088), .ZN(n3135) );
  OR2_X1 U3552 ( .A1(n4681), .A2(n4757), .ZN(n5008) );
  AND2_X4 U3553 ( .A1(n4768), .A2(n4756), .ZN(n4681) );
  AND2_X1 U3554 ( .A1(n3032), .A2(n4273), .ZN(n2967) );
  AND3_X4 U3555 ( .A1(n3017), .A2(n3136), .A3(n2955), .ZN(n3948) );
  NOR2_X4 U3556 ( .A1(n2974), .A2(n5068), .ZN(n5067) );
  XNOR2_X2 U3557 ( .A(n3404), .B(n3403), .ZN(n3512) );
  NAND2_X2 U3558 ( .A1(n3388), .A2(n3387), .ZN(n3404) );
  OAI21_X2 U3559 ( .B1(n5512), .B2(n3426), .A(n3425), .ZN(n4581) );
  NAND2_X2 U3560 ( .A1(n5321), .A2(n4536), .ZN(n5255) );
  NOR2_X4 U3561 ( .A1(n5323), .A2(n5322), .ZN(n5321) );
  AND2_X2 U3562 ( .A1(n4829), .A2(n4830), .ZN(n3923) );
  NOR2_X2 U3563 ( .A1(n4836), .A2(n4837), .ZN(n4829) );
  AND2_X2 U3564 ( .A1(n3164), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4178)
         );
  NAND2_X2 U3565 ( .A1(n4780), .A2(n4783), .ZN(n4781) );
  NOR2_X4 U3566 ( .A1(n4880), .A2(n4879), .ZN(n4780) );
  INV_X1 U3567 ( .A(n4731), .ZN(n4897) );
  NOR2_X2 U3568 ( .A1(n4417), .A2(n4519), .ZN(n4518) );
  AND2_X2 U3569 ( .A1(n4866), .A2(n2980), .ZN(n4845) );
  NOR2_X4 U3570 ( .A1(n4781), .A2(n4867), .ZN(n4866) );
  AND2_X1 U3571 ( .A1(n4183), .A2(n4268), .ZN(n2969) );
  NAND2_X1 U3572 ( .A1(n3445), .A2(n3444), .ZN(n3494) );
  AOI21_X1 U3573 ( .B1(n3143), .B2(n3142), .A(n4092), .ZN(n3144) );
  INV_X1 U3574 ( .A(n3351), .ZN(n3374) );
  NAND2_X1 U3575 ( .A1(n5662), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3275) );
  INV_X1 U3576 ( .A(n3250), .ZN(n3276) );
  NAND2_X1 U3577 ( .A1(n3493), .A2(n3492), .ZN(n3957) );
  OR2_X1 U3578 ( .A1(n3491), .A2(n3490), .ZN(n3493) );
  NOR2_X1 U3579 ( .A1(n4185), .A2(n6366), .ZN(n4154) );
  INV_X1 U3580 ( .A(n4419), .ZN(n4649) );
  INV_X1 U3581 ( .A(n4649), .ZN(n4655) );
  NAND2_X1 U3582 ( .A1(n3276), .A2(n3275), .ZN(n3498) );
  OR3_X1 U3583 ( .A1(n4240), .A2(n3964), .A3(n4239), .ZN(n5463) );
  NAND2_X1 U3584 ( .A1(n4160), .A2(n3013), .ZN(n3012) );
  INV_X1 U3585 ( .A(n4755), .ZN(n3013) );
  NAND2_X1 U3586 ( .A1(n3968), .A2(n3967), .ZN(n4093) );
  OR3_X1 U3587 ( .A1(n4240), .A2(n3966), .A3(n3142), .ZN(n3967) );
  CLKBUF_X1 U3588 ( .A(n3963), .Z(n3964) );
  AND2_X1 U3589 ( .A1(n3449), .A2(n3450), .ZN(n3468) );
  OR2_X1 U3590 ( .A1(n3463), .A2(n3462), .ZN(n3472) );
  INV_X1 U3591 ( .A(n3330), .ZN(n3331) );
  AND2_X1 U3592 ( .A1(n3386), .A2(n3385), .ZN(n3389) );
  AND2_X1 U3593 ( .A1(n2956), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3453) );
  INV_X1 U3594 ( .A(n3300), .ZN(n3292) );
  AND3_X1 U3595 ( .A1(n5684), .A2(n3150), .A3(n3146), .ZN(n4210) );
  INV_X1 U3596 ( .A(n4854), .ZN(n3008) );
  AND2_X1 U3597 ( .A1(n4861), .A2(n3798), .ZN(n3009) );
  INV_X1 U3598 ( .A(n4154), .ZN(n4652) );
  OR2_X1 U3599 ( .A1(n3007), .A2(n3698), .ZN(n3006) );
  INV_X1 U3600 ( .A(n4567), .ZN(n3666) );
  NOR2_X2 U3601 ( .A1(n3505), .A2(n3558), .ZN(n3693) );
  NAND2_X1 U3602 ( .A1(n5067), .A2(n4049), .ZN(n4839) );
  OR2_X1 U3603 ( .A1(n4989), .A2(n3433), .ZN(n2994) );
  NAND2_X1 U3604 ( .A1(n3453), .A2(n4072), .ZN(n3484) );
  OR2_X1 U3605 ( .A1(n3289), .A2(n3288), .ZN(n3344) );
  AND2_X1 U3606 ( .A1(n6010), .A2(n3192), .ZN(n5665) );
  NOR2_X1 U3607 ( .A1(n4086), .A2(n4084), .ZN(n4267) );
  NAND2_X1 U3608 ( .A1(n3500), .A2(n3499), .ZN(n4199) );
  NAND2_X1 U3609 ( .A1(n3498), .A2(n3497), .ZN(n3499) );
  NAND2_X1 U3610 ( .A1(n3496), .A2(n3495), .ZN(n3500) );
  XNOR2_X1 U3611 ( .A(n2958), .B(n5826), .ZN(n4263) );
  INV_X1 U3612 ( .A(n4618), .ZN(n5357) );
  INV_X1 U3613 ( .A(n4496), .ZN(n4709) );
  AND2_X1 U3614 ( .A1(n6368), .A2(n4422), .ZN(n5371) );
  AND2_X1 U3615 ( .A1(n4421), .A2(n5612), .ZN(n4422) );
  OR2_X1 U3616 ( .A1(n5371), .A2(n3558), .ZN(n4496) );
  AOI22_X1 U3617 ( .A1(n3922), .A2(n3921), .B1(n4419), .B2(n4769), .ZN(n3924)
         );
  INV_X1 U3618 ( .A(n3550), .ZN(n4658) );
  AOI22_X1 U3619 ( .A1(n4158), .A2(n4157), .B1(n4419), .B2(n4746), .ZN(n4160)
         );
  NAND2_X1 U3620 ( .A1(n3650), .A2(n3651), .ZN(n3667) );
  INV_X1 U3621 ( .A(n3003), .ZN(n3002) );
  INV_X1 U3622 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3630) );
  AND2_X1 U3623 ( .A1(n3519), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3578)
         );
  OR2_X1 U3624 ( .A1(n4199), .A2(n6236), .ZN(n4240) );
  NAND2_X1 U3625 ( .A1(n5203), .A2(n3438), .ZN(n3439) );
  OR2_X1 U3626 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4920)
         );
  INV_X1 U3627 ( .A(n2991), .ZN(n2990) );
  AOI21_X1 U3628 ( .B1(n2992), .B2(n3433), .A(n2978), .ZN(n2991) );
  NOR2_X1 U3629 ( .A1(n5203), .A2(n3422), .ZN(n3423) );
  AND2_X1 U3630 ( .A1(n6425), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3501) );
  CLKBUF_X1 U3631 ( .A(n4263), .Z(n4264) );
  AND2_X1 U3632 ( .A1(n4894), .A2(n4893), .ZN(n5409) );
  INV_X2 U3633 ( .A(n4894), .ZN(n5408) );
  AND2_X1 U3634 ( .A1(n4894), .A2(n4244), .ZN(n4606) );
  AND2_X1 U3635 ( .A1(n4093), .A2(n4073), .ZN(n5649) );
  INV_X1 U3636 ( .A(n4264), .ZN(n6103) );
  INV_X1 U3637 ( .A(n5947), .ZN(n5918) );
  NOR2_X1 U3638 ( .A1(n4092), .A2(n3952), .ZN(n3147) );
  OR2_X1 U3639 ( .A1(n3361), .A2(n3360), .ZN(n3391) );
  OR2_X1 U3640 ( .A1(n3384), .A2(n3383), .ZN(n3406) );
  NOR2_X1 U3641 ( .A1(n3152), .A2(n3124), .ZN(n3154) );
  AND2_X1 U3642 ( .A1(n3270), .A2(n6144), .ZN(n5913) );
  AOI22_X1 U3643 ( .A1(n3066), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U3644 ( .A1(n3118), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U3645 ( .A1(n3118), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U3646 ( .A1(n3119), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3086) );
  AOI22_X1 U3647 ( .A1(n2968), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3080) );
  INV_X1 U3648 ( .A(n3502), .ZN(n4079) );
  AND2_X1 U3649 ( .A1(n3484), .A2(n3485), .ZN(n3488) );
  AOI21_X1 U3650 ( .B1(n3472), .B2(n3471), .A(n3470), .ZN(n3489) );
  OR2_X1 U3651 ( .A1(n3494), .A2(n3957), .ZN(n3495) );
  AOI22_X1 U3652 ( .A1(n3066), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3060) );
  OR2_X1 U3653 ( .A1(n5133), .A2(n4649), .ZN(n3858) );
  OAI21_X1 U3654 ( .B1(n3402), .B2(n3484), .A(n3401), .ZN(n3403) );
  OR2_X1 U3655 ( .A1(n3209), .A2(n3208), .ZN(n3300) );
  AND2_X1 U3656 ( .A1(n3125), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3547) );
  NOR2_X1 U3657 ( .A1(n2977), .A2(n2993), .ZN(n2992) );
  INV_X1 U3658 ( .A(n3432), .ZN(n2993) );
  OR2_X1 U3659 ( .A1(n4182), .A2(n4083), .ZN(n4086) );
  NAND2_X1 U3660 ( .A1(n2989), .A2(n3444), .ZN(n3348) );
  OR2_X1 U3661 ( .A1(n3305), .A2(n3304), .ZN(n3265) );
  NAND2_X1 U3662 ( .A1(n4210), .A2(n3448), .ZN(n4180) );
  OAI21_X1 U3663 ( .B1(n5270), .B2(n6243), .A(n6333), .ZN(n5661) );
  INV_X1 U3664 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6213) );
  INV_X1 U3665 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6218) );
  OR2_X1 U3666 ( .A1(n4240), .A2(n4164), .ZN(n5113) );
  AND2_X1 U3667 ( .A1(n3959), .A2(n3958), .ZN(n4168) );
  NOR2_X1 U3668 ( .A1(n6303), .A2(n5296), .ZN(n5169) );
  AND2_X1 U3669 ( .A1(n3174), .A2(n3173), .ZN(n3182) );
  AND2_X1 U3670 ( .A1(n3815), .A2(n3814), .ZN(n4861) );
  OR2_X1 U3671 ( .A1(n3006), .A2(n3005), .ZN(n3004) );
  INV_X1 U3672 ( .A(n4796), .ZN(n3005) );
  AND2_X1 U3673 ( .A1(n4023), .A2(n4022), .ZN(n4608) );
  INV_X1 U3674 ( .A(n4579), .ZN(n2984) );
  AND2_X1 U3675 ( .A1(n3146), .A2(n3153), .ZN(n4893) );
  AND2_X1 U3676 ( .A1(n4225), .A2(n4431), .ZN(n5412) );
  OR2_X1 U3677 ( .A1(n4240), .A2(n4223), .ZN(n4224) );
  AND2_X1 U3678 ( .A1(n4113), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4115)
         );
  NAND2_X1 U3679 ( .A1(n4115), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4423)
         );
  AND2_X1 U3680 ( .A1(n3881), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3900)
         );
  NOR2_X1 U3681 ( .A1(n3856), .A2(n4950), .ZN(n3881) );
  INV_X1 U3682 ( .A(n4848), .ZN(n3862) );
  NAND2_X1 U3683 ( .A1(n3813), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3856)
         );
  INV_X1 U3684 ( .A(n3793), .ZN(n3794) );
  AND2_X1 U3685 ( .A1(n3760), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3761)
         );
  NAND2_X1 U3686 ( .A1(n3761), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3793)
         );
  NOR2_X1 U3687 ( .A1(n3728), .A2(n4803), .ZN(n3729) );
  AND2_X1 U3688 ( .A1(n3729), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3760)
         );
  NAND2_X1 U3689 ( .A1(n3713), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3728)
         );
  NOR2_X1 U3690 ( .A1(n3700), .A2(n3699), .ZN(n3713) );
  AND2_X1 U3691 ( .A1(n3646), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3647)
         );
  NAND2_X1 U3692 ( .A1(n3647), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3684)
         );
  NAND2_X1 U3693 ( .A1(n3645), .A2(n3644), .ZN(n4535) );
  NAND2_X1 U3694 ( .A1(n3614), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3631)
         );
  NOR2_X1 U3695 ( .A1(n3598), .A2(n3597), .ZN(n3614) );
  INV_X1 U3696 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3597) );
  CLKBUF_X1 U3697 ( .A(n4417), .Z(n4520) );
  NAND2_X1 U3698 ( .A1(n3583), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3598)
         );
  AND2_X1 U3699 ( .A1(n3578), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3583)
         );
  AOI21_X1 U3700 ( .B1(n3523), .B2(n3693), .A(n3522), .ZN(n4399) );
  NOR2_X1 U3701 ( .A1(n3563), .A2(n6431), .ZN(n3519) );
  INV_X1 U3702 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6431) );
  AND2_X1 U3703 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3507), .ZN(n3564)
         );
  INV_X1 U3704 ( .A(n3548), .ZN(n3507) );
  NAND2_X1 U3705 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3548) );
  INV_X1 U3706 ( .A(n4741), .ZN(n2983) );
  INV_X1 U3707 ( .A(n4839), .ZN(n2988) );
  AOI21_X1 U3708 ( .B1(n4971), .B2(n4970), .A(n4937), .ZN(n4965) );
  OR2_X1 U3709 ( .A1(n5203), .A2(n4625), .ZN(n3430) );
  NOR2_X1 U3710 ( .A1(n5570), .A2(n4091), .ZN(n4593) );
  NOR2_X1 U3711 ( .A1(n5255), .A2(n5256), .ZN(n5258) );
  AND2_X1 U3712 ( .A1(n3414), .A2(n3444), .ZN(n3415) );
  INV_X1 U3713 ( .A(n2997), .ZN(n2996) );
  OAI21_X1 U3714 ( .B1(n3420), .B2(n2998), .A(n4542), .ZN(n2997) );
  AND3_X1 U3715 ( .A1(n4010), .A2(n4027), .A3(n4009), .ZN(n4440) );
  AND2_X1 U3716 ( .A1(n4453), .A2(n4454), .ZN(n5332) );
  AND2_X1 U3717 ( .A1(n4008), .A2(n4007), .ZN(n5331) );
  NAND2_X1 U3718 ( .A1(n5332), .A2(n5331), .ZN(n5334) );
  NAND2_X1 U3719 ( .A1(n4468), .A2(n4470), .ZN(n4469) );
  AND3_X1 U3720 ( .A1(n3999), .A2(n4027), .A3(n3998), .ZN(n4375) );
  AOI21_X1 U3721 ( .B1(n5539), .B2(n3327), .A(n3326), .ZN(n4327) );
  NOR2_X1 U3722 ( .A1(n5538), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3326)
         );
  INV_X1 U3723 ( .A(n5103), .ZN(n5572) );
  NAND2_X1 U3724 ( .A1(n4221), .A2(n4438), .ZN(n4220) );
  NAND2_X1 U3725 ( .A1(n3249), .A2(n3319), .ZN(n3253) );
  INV_X1 U3726 ( .A(n3319), .ZN(n3251) );
  NAND2_X1 U3727 ( .A1(n4263), .A2(n6366), .ZN(n3291) );
  OR2_X1 U3728 ( .A1(n3148), .A2(n3503), .ZN(n4185) );
  AND3_X1 U3729 ( .A1(n4201), .A2(n4200), .A3(n4212), .ZN(n6211) );
  NOR2_X1 U3730 ( .A1(n5762), .A2(n5917), .ZN(n5712) );
  OR2_X1 U3731 ( .A1(n3526), .A2(n5663), .ZN(n5762) );
  INV_X1 U3732 ( .A(n2956), .ZN(n5662) );
  INV_X1 U3733 ( .A(n6344), .ZN(n6071) );
  NAND3_X1 U3734 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6366), .A3(n5661), .ZN(
        n5704) );
  INV_X1 U3735 ( .A(n4199), .ZN(n4177) );
  INV_X1 U3736 ( .A(n6251), .ZN(n6236) );
  NAND2_X1 U3737 ( .A1(n4709), .A2(n4429), .ZN(n4618) );
  INV_X1 U3738 ( .A(n5377), .ZN(n5367) );
  INV_X1 U3739 ( .A(n5374), .ZN(n5364) );
  OR2_X1 U3740 ( .A1(n5371), .A2(n6331), .ZN(n5374) );
  AND2_X1 U3741 ( .A1(n4488), .A2(n5164), .ZN(n5382) );
  AND2_X1 U3742 ( .A1(n4884), .A2(n4883), .ZN(n5298) );
  INV_X1 U3743 ( .A(n5178), .ZN(n5393) );
  AND2_X2 U3744 ( .A1(n4213), .A2(n6251), .ZN(n5398) );
  INV_X1 U3745 ( .A(n5182), .ZN(n5406) );
  NAND2_X1 U3746 ( .A1(n4241), .A2(n5463), .ZN(n4894) );
  OAI21_X1 U3747 ( .B1(n4238), .B2(n4237), .A(n6251), .ZN(n4241) );
  INV_X1 U3748 ( .A(n4606), .ZN(n4402) );
  CLKBUF_X1 U3749 ( .A(n5496), .Z(n5506) );
  XNOR2_X1 U3750 ( .A(n4424), .B(n4711), .ZN(n4704) );
  OR2_X1 U3751 ( .A1(n4654), .A2(n4698), .ZN(n4424) );
  XNOR2_X1 U3752 ( .A(n3014), .B(n4660), .ZN(n4708) );
  NOR2_X1 U3753 ( .A1(n4136), .A2(n3011), .ZN(n3014) );
  OR2_X1 U3754 ( .A1(n3012), .A2(n4695), .ZN(n3011) );
  OAI21_X1 U3755 ( .B1(n4159), .B2(n4160), .A(n4694), .ZN(n4900) );
  INV_X1 U3756 ( .A(n4923), .ZN(n5183) );
  NAND2_X1 U3757 ( .A1(n3002), .A2(n3667), .ZN(n4569) );
  INV_X1 U3758 ( .A(n5546), .ZN(n5517) );
  INV_X1 U3759 ( .A(n5550), .ZN(n5536) );
  INV_X1 U3760 ( .A(n5555), .ZN(n5541) );
  OR2_X1 U3761 ( .A1(n4240), .A2(n6226), .ZN(n5555) );
  OR2_X1 U3762 ( .A1(n5651), .A2(n5244), .ZN(n5103) );
  INV_X1 U3763 ( .A(n4922), .ZN(n3001) );
  NOR2_X1 U3764 ( .A1(n5264), .A2(n4107), .ZN(n5229) );
  INV_X1 U3765 ( .A(n5654), .ZN(n5636) );
  INV_X1 U3766 ( .A(n5077), .ZN(n5632) );
  INV_X1 U3767 ( .A(n4310), .ZN(n4339) );
  INV_X1 U3768 ( .A(n5764), .ZN(n5663) );
  INV_X1 U3769 ( .A(n6348), .ZN(n6352) );
  INV_X1 U3770 ( .A(n6345), .ZN(n6370) );
  OAI21_X1 U3771 ( .B1(n5669), .B2(n5711), .A(n5668), .ZN(n5708) );
  OAI221_X1 U3772 ( .B1(n5756), .B2(n6331), .C1(n5756), .C2(n5741), .A(n5984), 
        .ZN(n5758) );
  INV_X1 U3773 ( .A(n5854), .ZN(n5844) );
  OAI21_X1 U3774 ( .B1(n5927), .B2(n5926), .A(n5925), .ZN(n5944) );
  INV_X1 U3775 ( .A(n6008), .ZN(n5980) );
  INV_X1 U3776 ( .A(n6070), .ZN(n6043) );
  INV_X1 U3777 ( .A(n6101), .ZN(n6089) );
  OAI211_X1 U3778 ( .C1(n6138), .C2(n6331), .A(n6111), .B(n6110), .ZN(n6140)
         );
  INV_X1 U3779 ( .A(n6209), .ZN(n6188) );
  AND2_X1 U3780 ( .A1(n5702), .A2(DATAI_22_), .ZN(n6196) );
  AND2_X1 U3781 ( .A1(DATAI_6_), .A2(n5921), .ZN(n6194) );
  NAND2_X1 U3782 ( .A1(n4177), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6333) );
  AND2_X1 U3783 ( .A1(n3501), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6251) );
  INV_X1 U3784 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6425) );
  INV_X1 U3785 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6523) );
  AND2_X1 U3786 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6523), .ZN(n6376) );
  AOI21_X1 U3787 ( .B1(n4820), .B2(n5649), .A(n2985), .ZN(n4109) );
  NAND2_X1 U3788 ( .A1(n4108), .A2(n2986), .ZN(n2985) );
  NOR2_X1 U3789 ( .A1(n4106), .A2(n4702), .ZN(n2986) );
  INV_X1 U3790 ( .A(n3148), .ZN(n3152) );
  AND4_X1 U3791 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n2970)
         );
  NOR2_X1 U3792 ( .A1(n4136), .A2(n4755), .ZN(n4159) );
  NOR2_X1 U3793 ( .A1(n4572), .A2(n3006), .ZN(n2971) );
  NAND2_X1 U3794 ( .A1(n4866), .A2(n3009), .ZN(n4852) );
  AND2_X1 U3795 ( .A1(n4470), .A2(n4541), .ZN(n2972) );
  OR2_X2 U3796 ( .A1(n3046), .A2(n3045), .ZN(n3175) );
  INV_X1 U3797 ( .A(n3975), .ZN(n3982) );
  NAND2_X2 U3798 ( .A1(n5684), .A2(n3159), .ZN(n3975) );
  NAND2_X1 U3799 ( .A1(n2994), .A2(n3432), .ZN(n4983) );
  AND4_X1 U3800 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n2973)
         );
  AND2_X1 U3801 ( .A1(n3124), .A2(n3160), .ZN(n3448) );
  NAND2_X1 U3802 ( .A1(n4845), .A2(n3862), .ZN(n4836) );
  AND2_X1 U3803 ( .A1(n4866), .A2(n3798), .ZN(n4860) );
  OR2_X1 U3804 ( .A1(n4206), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n2975)
         );
  INV_X1 U3805 ( .A(n3010), .ZN(n4694) );
  INV_X1 U3806 ( .A(n4541), .ZN(n2998) );
  NAND2_X1 U3807 ( .A1(n2994), .A2(n2992), .ZN(n4934) );
  INV_X1 U3808 ( .A(n3506), .ZN(n3877) );
  INV_X1 U3809 ( .A(n3877), .ZN(n4659) );
  INV_X1 U3810 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2982) );
  INV_X1 U3811 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3164) );
  OR2_X1 U3812 ( .A1(n4572), .A2(n3698), .ZN(n2976) );
  OAI21_X1 U3813 ( .B1(n4581), .B2(n4584), .A(n4582), .ZN(n5217) );
  NAND2_X1 U3814 ( .A1(n4469), .A2(n3420), .ZN(n4540) );
  AND2_X1 U3815 ( .A1(n5203), .A2(n3434), .ZN(n2977) );
  NAND2_X1 U3816 ( .A1(n3667), .A2(n2959), .ZN(n4566) );
  NAND2_X1 U3817 ( .A1(n3291), .A2(n3290), .ZN(n4338) );
  NOR2_X1 U3818 ( .A1(n5203), .A2(n3435), .ZN(n2978) );
  AND2_X1 U3819 ( .A1(n3613), .A2(n4393), .ZN(n2979) );
  NAND2_X1 U3820 ( .A1(n3003), .A2(n3667), .ZN(n4573) );
  AND2_X1 U3821 ( .A1(n3009), .A2(n3008), .ZN(n2980) );
  AOI21_X1 U3822 ( .B1(n3512), .B2(n3693), .A(n3511), .ZN(n4398) );
  NAND2_X1 U3823 ( .A1(n3557), .A2(n3556), .ZN(n4317) );
  AOI21_X1 U3824 ( .B1(n3526), .B2(n3693), .A(n3531), .ZN(n4328) );
  AND2_X1 U3825 ( .A1(n4054), .A2(n4849), .ZN(n2981) );
  NOR2_X2 U3826 ( .A1(n5692), .A2(n5674), .ZN(n6116) );
  AND2_X2 U3827 ( .A1(n2982), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3031)
         );
  INV_X1 U3828 ( .A(n4681), .ZN(n4680) );
  AND2_X1 U3829 ( .A1(n4681), .A2(n2983), .ZN(n4066) );
  AND2_X2 U3830 ( .A1(n4833), .A2(n4766), .ZN(n4768) );
  NOR3_X4 U3831 ( .A1(n5255), .A2(n5256), .A3(n2984), .ZN(n4609) );
  NOR2_X2 U3832 ( .A1(n4810), .A2(n4030), .ZN(n4784) );
  NAND2_X2 U3833 ( .A1(n4609), .A2(n4608), .ZN(n4810) );
  NOR2_X2 U3834 ( .A1(n4336), .A2(n4335), .ZN(n4334) );
  OR2_X2 U3835 ( .A1(n5334), .A2(n4440), .ZN(n5323) );
  AOI21_X1 U3836 ( .B1(n2989), .B2(n3693), .A(n3567), .ZN(n4318) );
  INV_X1 U3837 ( .A(n3168), .ZN(n3268) );
  AND2_X2 U3838 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4269) );
  AOI22_X1 U3839 ( .A1(n3066), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3067) );
  AND2_X2 U3840 ( .A1(n3031), .A2(n4184), .ZN(n3066) );
  AOI21_X2 U3841 ( .B1(n4989), .B2(n2992), .A(n2990), .ZN(n4975) );
  INV_X1 U3842 ( .A(n4996), .ZN(n5006) );
  NAND2_X1 U3843 ( .A1(n4111), .A2(n3000), .ZN(n2999) );
  NAND2_X1 U3844 ( .A1(n3001), .A2(n4110), .ZN(n3000) );
  NOR2_X4 U3845 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4183) );
  NAND2_X1 U3846 ( .A1(n3654), .A2(n3666), .ZN(n3003) );
  OR2_X2 U3847 ( .A1(n4572), .A2(n3004), .ZN(n4880) );
  INV_X1 U3848 ( .A(n4808), .ZN(n3007) );
  NOR2_X2 U3849 ( .A1(n4136), .A2(n3012), .ZN(n3010) );
  NAND3_X1 U3850 ( .A1(n4391), .A2(n4392), .A3(n4393), .ZN(n4390) );
  NAND3_X1 U3851 ( .A1(n4391), .A2(n4392), .A3(n2979), .ZN(n4417) );
  NOR2_X1 U3852 ( .A1(n3937), .A2(n3442), .ZN(n3443) );
  AOI21_X1 U3853 ( .B1(n4731), .B2(n5702), .A(n4699), .ZN(n4700) );
  XOR2_X1 U3854 ( .A(n4695), .B(n4694), .Z(n4731) );
  XNOR2_X1 U3855 ( .A(n4678), .B(n4691), .ZN(n4701) );
  AND2_X2 U3856 ( .A1(n3029), .A2(n4178), .ZN(n3119) );
  NOR2_X1 U3857 ( .A1(n2963), .A2(n3020), .ZN(n4678) );
  INV_X1 U3858 ( .A(n4309), .ZN(n5764) );
  INV_X1 U3859 ( .A(n5703), .ZN(n5921) );
  AND4_X1 U3860 ( .A1(n3036), .A2(n3035), .A3(n3034), .A4(n3033), .ZN(n3015)
         );
  INV_X1 U3861 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3438) );
  INV_X1 U3862 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3945) );
  INV_X1 U3863 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4299) );
  INV_X1 U3864 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3699) );
  AND4_X1 U3865 ( .A1(n3028), .A2(n3027), .A3(n3026), .A4(n3025), .ZN(n3018)
         );
  INV_X1 U3866 ( .A(n4416), .ZN(n3613) );
  INV_X1 U3867 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3479) );
  OR2_X1 U3868 ( .A1(n3140), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3019)
         );
  INV_X1 U3869 ( .A(n5203), .ZN(n5204) );
  AND2_X1 U3870 ( .A1(n4676), .A2(n4675), .ZN(n3020) );
  AOI21_X2 U3871 ( .B1(n3152), .B2(n5690), .A(n3149), .ZN(n3169) );
  AND2_X1 U3872 ( .A1(n3373), .A2(n3372), .ZN(n3021) );
  NAND2_X1 U3873 ( .A1(n3305), .A2(n3304), .ZN(n3022) );
  INV_X1 U3874 ( .A(n5639), .ZN(n4380) );
  NAND2_X1 U3875 ( .A1(n4894), .A2(n4243), .ZN(n5182) );
  AND2_X1 U3876 ( .A1(n5398), .A2(n2961), .ZN(n5394) );
  NAND2_X1 U3877 ( .A1(n5398), .A2(n3132), .ZN(n5178) );
  INV_X1 U3878 ( .A(n4846), .ZN(n4853) );
  AND2_X1 U3879 ( .A1(n6349), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3465)
         );
  AOI21_X1 U3880 ( .B1(n3148), .B2(n3175), .A(n3132), .ZN(n3133) );
  AND2_X1 U3881 ( .A1(n6252), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3173) );
  OR2_X1 U3882 ( .A1(n3341), .A2(n3340), .ZN(n3392) );
  NAND2_X1 U3883 ( .A1(n3169), .A2(n3150), .ZN(n3502) );
  INV_X1 U3884 ( .A(n3414), .ZN(n3259) );
  AND2_X1 U3886 ( .A1(n3150), .A2(n3175), .ZN(n3090) );
  INV_X1 U3887 ( .A(n4604), .ZN(n3698) );
  INV_X1 U3888 ( .A(n5513), .ZN(n3424) );
  OR2_X1 U3889 ( .A1(n3224), .A2(n3223), .ZN(n3308) );
  AOI22_X1 U3890 ( .A1(n3077), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3074) );
  NOR2_X1 U3891 ( .A1(n4072), .A2(n6366), .ZN(n3250) );
  INV_X1 U3892 ( .A(n4962), .ZN(n3798) );
  OR2_X1 U3893 ( .A1(n4423), .A2(n4748), .ZN(n4654) );
  OAI21_X1 U3894 ( .B1(n3489), .B2(n3488), .A(n3487), .ZN(n3496) );
  NOR2_X1 U3895 ( .A1(n3424), .A2(n3423), .ZN(n3425) );
  NAND2_X1 U3896 ( .A1(n3274), .A2(n3273), .ZN(n5826) );
  NOR2_X1 U3897 ( .A1(n6300), .A2(n4816), .ZN(n4802) );
  INV_X1 U3898 ( .A(n4964), .ZN(n4938) );
  INV_X1 U3899 ( .A(n3157), .ZN(n4072) );
  AND2_X1 U3900 ( .A1(n5952), .A2(n6345), .ZN(n5954) );
  INV_X1 U3901 ( .A(n6109), .ZN(n6145) );
  AND2_X1 U3902 ( .A1(n3900), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3901)
         );
  INV_X1 U3903 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5304) );
  AND2_X1 U3904 ( .A1(n4618), .A2(n4617), .ZN(n4723) );
  NAND2_X1 U3905 ( .A1(n3975), .A2(n4869), .ZN(n4206) );
  AND2_X1 U3906 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3794), .ZN(n3813)
         );
  OR2_X1 U3907 ( .A1(n3684), .A2(n5304), .ZN(n3700) );
  NOR2_X1 U3908 ( .A1(n3631), .A2(n3630), .ZN(n3646) );
  INV_X1 U3909 ( .A(n5649), .ZN(n5585) );
  OR2_X1 U3910 ( .A1(n5115), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5612) );
  INV_X1 U3911 ( .A(n4338), .ZN(n4342) );
  AND2_X1 U3912 ( .A1(n5982), .A2(n4264), .ZN(n6013) );
  INV_X1 U3913 ( .A(n4339), .ZN(n5917) );
  NAND2_X1 U3914 ( .A1(n6366), .A2(n5661), .ZN(n5703) );
  INV_X1 U3915 ( .A(n6364), .ZN(n4434) );
  AND2_X1 U3916 ( .A1(n4764), .A2(REIP_REG_28__SCAN_IN), .ZN(n4753) );
  NAND2_X1 U3917 ( .A1(n3901), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4112)
         );
  INV_X1 U3918 ( .A(n5164), .ZN(n5351) );
  INV_X1 U3919 ( .A(n4866), .ZN(n4963) );
  INV_X1 U3920 ( .A(n5207), .ZN(n5399) );
  INV_X1 U3921 ( .A(n4572), .ZN(n4605) );
  NAND2_X1 U3922 ( .A1(n3564), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3563)
         );
  NAND2_X1 U3923 ( .A1(n5555), .A2(n3926), .ZN(n5550) );
  NOR2_X1 U3924 ( .A1(n4594), .A2(n4380), .ZN(n5222) );
  OR2_X1 U3925 ( .A1(n5651), .A2(n4094), .ZN(n5569) );
  AND2_X1 U3926 ( .A1(n4100), .A2(n5569), .ZN(n5639) );
  AND2_X1 U3927 ( .A1(n4093), .A2(n6216), .ZN(n5651) );
  NOR2_X1 U3928 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6252) );
  INV_X1 U3929 ( .A(n5761), .ZN(n5739) );
  INV_X1 U3930 ( .A(n5732), .ZN(n5734) );
  INV_X1 U3931 ( .A(n5790), .ZN(n5791) );
  OAI21_X1 U3932 ( .B1(n5819), .B2(n6331), .A(n5804), .ZN(n5821) );
  INV_X1 U3933 ( .A(n5880), .ZN(n5856) );
  OR2_X1 U3934 ( .A1(n5882), .A2(n5917), .ZN(n5825) );
  INV_X1 U3935 ( .A(n5904), .ZN(n5906) );
  INV_X1 U3936 ( .A(n5978), .ZN(n5968) );
  OR2_X1 U3937 ( .A1(n6012), .A2(n5917), .ZN(n5951) );
  INV_X1 U3938 ( .A(n6040), .ZN(n6030) );
  NAND2_X1 U3939 ( .A1(n5764), .A2(n3526), .ZN(n6012) );
  INV_X1 U3940 ( .A(n6143), .ZN(n6107) );
  AND2_X1 U3941 ( .A1(n5113), .A2(n5114), .ZN(n6368) );
  INV_X1 U3942 ( .A(n5368), .ZN(n5361) );
  OR2_X1 U3943 ( .A1(n5371), .A2(n4426), .ZN(n5164) );
  OR2_X1 U3944 ( .A1(n5371), .A2(n4443), .ZN(n5386) );
  OR2_X1 U3945 ( .A1(n3923), .A2(n4831), .ZN(n4923) );
  INV_X1 U3946 ( .A(n5412), .ZN(n5430) );
  OR2_X2 U3947 ( .A1(n4240), .A2(n6239), .ZN(n5511) );
  NAND2_X1 U3948 ( .A1(n5550), .A2(n3929), .ZN(n5546) );
  NOR2_X1 U3949 ( .A1(n4593), .A2(n5222), .ZN(n5264) );
  NAND2_X1 U3950 ( .A1(n4093), .A2(n3974), .ZN(n5654) );
  INV_X1 U3951 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U3952 ( .A1(n5712), .A2(n6344), .ZN(n5761) );
  OR2_X1 U3953 ( .A1(n5762), .A2(n5979), .ZN(n5790) );
  OR2_X1 U3954 ( .A1(n5762), .A2(n6009), .ZN(n5824) );
  OR2_X1 U3955 ( .A1(n5825), .A2(n6344), .ZN(n5854) );
  OR2_X1 U3956 ( .A1(n5825), .A2(n6071), .ZN(n5880) );
  OR2_X1 U3957 ( .A1(n5882), .A2(n5979), .ZN(n5904) );
  OR2_X1 U3958 ( .A1(n5882), .A2(n6009), .ZN(n5947) );
  OR2_X1 U3959 ( .A1(n5951), .A2(n6344), .ZN(n5978) );
  OR2_X1 U3960 ( .A1(n5951), .A2(n6071), .ZN(n6008) );
  OR2_X1 U3961 ( .A1(n6012), .A2(n5979), .ZN(n6040) );
  OR2_X1 U3962 ( .A1(n6012), .A2(n6009), .ZN(n6070) );
  OR2_X1 U3963 ( .A1(n6072), .A2(n6344), .ZN(n6101) );
  OR2_X1 U3964 ( .A1(n6072), .A2(n6071), .ZN(n6143) );
  OR2_X1 U3965 ( .A1(n6150), .A2(n6071), .ZN(n6192) );
  INV_X1 U3966 ( .A(n6328), .ZN(n6324) );
  INV_X1 U3967 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6267) );
  INV_X1 U3968 ( .A(n6542), .ZN(n6319) );
  NAND2_X1 U3969 ( .A1(n3936), .A2(n3935), .ZN(U2959) );
  AOI22_X1 U3970 ( .A1(n3117), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3028) );
  AND2_X2 U3971 ( .A1(n3031), .A2(n4183), .ZN(n3237) );
  AOI22_X1 U3972 ( .A1(n4637), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3027) );
  INV_X1 U3973 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3024) );
  AND2_X2 U3974 ( .A1(n3030), .A2(n3031), .ZN(n3078) );
  AOI22_X1 U3975 ( .A1(n3077), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3078), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3026) );
  AOI22_X1 U3976 ( .A1(n3119), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3025) );
  AND2_X2 U3977 ( .A1(n4178), .A2(n4269), .ZN(n3282) );
  AND2_X2 U3978 ( .A1(n4183), .A2(n4269), .ZN(n3199) );
  AOI22_X1 U3979 ( .A1(n3282), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3036) );
  AND2_X4 U3980 ( .A1(n3029), .A2(n4183), .ZN(n3079) );
  AND2_X2 U3981 ( .A1(n4268), .A2(n4184), .ZN(n3242) );
  AOI22_X1 U3982 ( .A1(n2968), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3035) );
  AOI22_X1 U3983 ( .A1(n3118), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3066), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3034) );
  AND2_X2 U3984 ( .A1(n4178), .A2(n4268), .ZN(n3197) );
  AOI22_X1 U3985 ( .A1(n3197), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3033) );
  NAND2_X1 U3986 ( .A1(n3018), .A2(n3015), .ZN(n3142) );
  INV_X2 U3987 ( .A(n3142), .ZN(n3150) );
  AOI22_X1 U3988 ( .A1(n2968), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3040) );
  AOI22_X1 U3989 ( .A1(n3077), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3039) );
  AOI22_X1 U3990 ( .A1(n4637), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3038) );
  AOI22_X1 U3991 ( .A1(n3078), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3037) );
  NAND4_X1 U3992 ( .A1(n3040), .A2(n3039), .A3(n3038), .A4(n3037), .ZN(n3046)
         );
  AOI22_X1 U3993 ( .A1(n3118), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3044) );
  AOI22_X1 U3994 ( .A1(n3119), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3043) );
  AOI22_X1 U3995 ( .A1(n3282), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3042) );
  AOI22_X1 U3996 ( .A1(n3066), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3041) );
  NAND4_X1 U3997 ( .A1(n3044), .A2(n3043), .A3(n3042), .A4(n3041), .ZN(n3045)
         );
  AOI22_X1 U3998 ( .A1(n3117), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4637), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3050) );
  AOI22_X1 U3999 ( .A1(n3237), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3066), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3049) );
  AOI22_X1 U4000 ( .A1(n2968), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3048) );
  AOI22_X1 U4001 ( .A1(n3077), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3047) );
  AOI22_X1 U4002 ( .A1(n3078), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3054) );
  AOI22_X1 U4003 ( .A1(n3197), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U4004 ( .A1(n3119), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        INSTQUEUE_REG_2__5__SCAN_IN), .B2(n3118), .ZN(n3052) );
  AOI22_X1 U4005 ( .A1(n3242), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3051) );
  AND4_X2 U4006 ( .A1(n3054), .A2(n3053), .A3(n3052), .A4(n3051), .ZN(n3055)
         );
  AOI22_X1 U4007 ( .A1(n2968), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3059) );
  AOI22_X1 U4008 ( .A1(n3077), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3058) );
  AOI22_X1 U4009 ( .A1(n4637), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U4010 ( .A1(n3078), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3056) );
  NAND4_X1 U4011 ( .A1(n3059), .A2(n3058), .A3(n3057), .A4(n3056), .ZN(n3065)
         );
  AOI22_X1 U4012 ( .A1(n3119), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3063) );
  AOI22_X1 U4013 ( .A1(n3118), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3062) );
  AOI22_X1 U4014 ( .A1(n3282), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3061) );
  NAND4_X1 U4015 ( .A1(n3063), .A2(n3062), .A3(n3061), .A4(n3060), .ZN(n3064)
         );
  AOI22_X1 U4016 ( .A1(n3119), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3070) );
  AOI22_X1 U4017 ( .A1(n3282), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3068) );
  AOI22_X1 U4018 ( .A1(n2968), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3073) );
  AOI22_X1 U4019 ( .A1(n4637), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3072) );
  AOI22_X1 U4020 ( .A1(n3078), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3071) );
  NAND2_X1 U4021 ( .A1(n3157), .A2(n3155), .ZN(n3451) );
  AOI22_X1 U4022 ( .A1(n3077), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3083) );
  AOI22_X1 U4023 ( .A1(n4637), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3082) );
  AOI22_X1 U4024 ( .A1(n3078), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3081) );
  AOI22_X1 U4025 ( .A1(n3117), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        INSTQUEUE_REG_2__6__SCAN_IN), .B2(n3118), .ZN(n3087) );
  AOI22_X1 U4026 ( .A1(n3282), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3085) );
  AOI22_X1 U4027 ( .A1(n3066), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3084) );
  NAND3_X1 U4028 ( .A1(n3090), .A2(n4893), .A3(n3170), .ZN(n3963) );
  INV_X1 U4029 ( .A(n3963), .ZN(n3112) );
  NAND2_X1 U4030 ( .A1(n3077), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3094)
         );
  NAND2_X1 U4031 ( .A1(n4637), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3093) );
  NAND2_X1 U4032 ( .A1(n3066), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3092)
         );
  NAND2_X1 U4033 ( .A1(n3198), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U4034 ( .A1(n3078), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3098)
         );
  NAND2_X1 U4035 ( .A1(n3117), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U4036 ( .A1(n3119), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U4037 ( .A1(n3282), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3095)
         );
  NAND2_X1 U4038 ( .A1(n3237), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3102) );
  NAND2_X1 U4039 ( .A1(n3079), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3101) );
  NAND2_X1 U4040 ( .A1(n3197), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3100) );
  NAND2_X1 U4041 ( .A1(n3199), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3099)
         );
  NAND2_X1 U4042 ( .A1(n3118), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U4043 ( .A1(n2969), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U4044 ( .A1(n3230), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U4045 ( .A1(n2953), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3104)
         );
  NAND2_X1 U4046 ( .A1(n3112), .A2(n2956), .ZN(n4164) );
  AOI22_X1 U4047 ( .A1(n2968), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U4048 ( .A1(n3077), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4049 ( .A1(n4637), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4050 ( .A1(n3078), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4051 ( .A1(n3119), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n2969), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3122) );
  AOI22_X1 U4052 ( .A1(n3282), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3121) );
  XNOR2_X1 U4053 ( .A(n6267), .B(STATE_REG_2__SCAN_IN), .ZN(n3952) );
  INV_X1 U4054 ( .A(n3159), .ZN(n3124) );
  INV_X1 U4055 ( .A(n4180), .ZN(n3126) );
  NAND2_X1 U4056 ( .A1(n3135), .A2(n3153), .ZN(n4661) );
  INV_X1 U4057 ( .A(n4661), .ZN(n3125) );
  NAND2_X1 U4058 ( .A1(n3126), .A2(n3125), .ZN(n3971) );
  OAI21_X1 U4059 ( .B1(n4164), .B2(n3147), .A(n3971), .ZN(n3127) );
  INV_X1 U4060 ( .A(n3127), .ZN(n3137) );
  NAND2_X1 U4061 ( .A1(n3135), .A2(n3155), .ZN(n3129) );
  NAND2_X1 U4062 ( .A1(n3129), .A2(n3128), .ZN(n3130) );
  NAND2_X1 U4063 ( .A1(n3130), .A2(n3150), .ZN(n3134) );
  INV_X1 U4064 ( .A(n3153), .ZN(n3132) );
  NAND2_X1 U4065 ( .A1(n3131), .A2(n3153), .ZN(n3176) );
  NAND2_X1 U4066 ( .A1(n3170), .A2(n3176), .ZN(n3143) );
  INV_X1 U4067 ( .A(n3143), .ZN(n3136) );
  NAND2_X1 U4068 ( .A1(n3137), .A2(n3970), .ZN(n3138) );
  NAND2_X1 U4069 ( .A1(n3138), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3165) );
  INV_X1 U4070 ( .A(n3165), .ZN(n3141) );
  NAND2_X1 U4071 ( .A1(n6252), .A2(n6366), .ZN(n6369) );
  INV_X1 U4072 ( .A(n6369), .ZN(n3272) );
  XNOR2_X1 U4073 ( .A(n6349), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5914)
         );
  INV_X1 U4074 ( .A(n3501), .ZN(n3271) );
  AND2_X1 U4075 ( .A1(n3271), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3139)
         );
  AOI21_X1 U4076 ( .B1(n3272), .B2(n5914), .A(n3139), .ZN(n3166) );
  INV_X1 U4077 ( .A(n3166), .ZN(n3140) );
  NAND2_X1 U4078 ( .A1(n3141), .A2(n3019), .ZN(n3167) );
  NAND2_X1 U4079 ( .A1(n3144), .A2(n3017), .ZN(n3145) );
  NAND2_X1 U4080 ( .A1(n3145), .A2(n2955), .ZN(n3184) );
  INV_X1 U4081 ( .A(n3146), .ZN(n3310) );
  NOR2_X1 U4082 ( .A1(n3147), .A2(n3310), .ZN(n3151) );
  NAND2_X1 U4083 ( .A1(n3153), .A2(n3175), .ZN(n3149) );
  NAND2_X1 U4084 ( .A1(n3170), .A2(n3153), .ZN(n3161) );
  NAND2_X1 U4085 ( .A1(n3154), .A2(n3161), .ZN(n4076) );
  INV_X1 U4086 ( .A(n3444), .ZN(n3158) );
  NAND4_X1 U4087 ( .A1(n3184), .A2(n3162), .A3(n4076), .A4(n3179), .ZN(n3163)
         );
  NAND2_X1 U4088 ( .A1(n3163), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3168) );
  OAI211_X1 U4089 ( .C1(n3168), .C2(n3164), .A(n3166), .B(n3165), .ZN(n3188)
         );
  AND2_X2 U4090 ( .A1(n3167), .A2(n3188), .ZN(n3213) );
  MUX2_X1 U4091 ( .A(n3501), .B(n6369), .S(n6349), .Z(n3540) );
  NAND2_X1 U4092 ( .A1(n3539), .A2(n3540), .ZN(n3187) );
  INV_X1 U4093 ( .A(n3169), .ZN(n3172) );
  NOR2_X1 U4094 ( .A1(n3170), .A2(n3152), .ZN(n3171) );
  OAI21_X1 U4095 ( .B1(n3172), .B2(n3171), .A(n4092), .ZN(n3174) );
  NAND2_X1 U4096 ( .A1(n3152), .A2(n6364), .ZN(n4074) );
  AND3_X1 U4097 ( .A1(n3150), .A2(n5684), .A3(n4072), .ZN(n3177) );
  INV_X1 U4098 ( .A(n3176), .ZN(n3537) );
  NAND2_X1 U4099 ( .A1(n3177), .A2(n3537), .ZN(n4286) );
  NAND3_X1 U4100 ( .A1(n4074), .A2(n4286), .A3(n3975), .ZN(n3181) );
  INV_X1 U4101 ( .A(n3179), .ZN(n3180) );
  OAI22_X1 U4102 ( .A1(n3184), .A2(n3183), .B1(n5662), .B2(n3150), .ZN(n4081)
         );
  INV_X1 U4103 ( .A(n4081), .ZN(n3185) );
  NAND2_X1 U4104 ( .A1(n3213), .A2(n3212), .ZN(n3189) );
  NAND2_X1 U4105 ( .A1(n3189), .A2(n3188), .ZN(n3195) );
  AND2_X1 U4106 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U4107 ( .A1(n3190), .A2(n6213), .ZN(n6010) );
  INV_X1 U4108 ( .A(n3190), .ZN(n3191) );
  NAND2_X1 U4109 ( .A1(n3191), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3192) );
  OAI22_X1 U4110 ( .A1(n5665), .A2(n6369), .B1(n3501), .B2(n6213), .ZN(n3193)
         );
  NAND2_X1 U4111 ( .A1(n3195), .A2(n3194), .ZN(n3196) );
  AOI22_X1 U4112 ( .A1(n3079), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3203) );
  AOI22_X1 U4113 ( .A1(n4146), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U4114 ( .A1(n4120), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4115 ( .A1(n3672), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3200) );
  NAND4_X1 U4116 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3209)
         );
  AOI22_X1 U4117 ( .A1(n3118), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3207) );
  INV_X1 U4118 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6491) );
  AOI22_X1 U4119 ( .A1(n3281), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4120 ( .A1(n3282), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4121 ( .A1(n4125), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3204) );
  NAND4_X1 U4122 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3208)
         );
  OAI22_X2 U4123 ( .A1(n4282), .A2(STATE2_REG_0__SCAN_IN), .B1(n3292), .B2(
        n3276), .ZN(n3211) );
  INV_X1 U4124 ( .A(n3275), .ZN(n3261) );
  XNOR2_X2 U4125 ( .A(n3211), .B(n3210), .ZN(n3299) );
  INV_X1 U4126 ( .A(n3213), .ZN(n3214) );
  AOI22_X1 U4127 ( .A1(n3281), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4128 ( .A1(n4145), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U4129 ( .A1(n4140), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4131 ( .A1(n3079), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3215) );
  NAND4_X1 U4132 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n3224)
         );
  AOI22_X1 U4133 ( .A1(n4146), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U4134 ( .A1(n4147), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4135 ( .A1(n4120), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4136 ( .A1(n4125), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3219) );
  NAND4_X1 U4137 ( .A1(n3222), .A2(n3221), .A3(n3220), .A4(n3219), .ZN(n3223)
         );
  NAND2_X1 U4138 ( .A1(n3250), .A2(n3308), .ZN(n3225) );
  AOI22_X1 U4139 ( .A1(n3079), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3229) );
  AOI22_X1 U4140 ( .A1(n4272), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4141 ( .A1(n4120), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4142 ( .A1(n3077), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3283), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3226) );
  NAND4_X1 U4143 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3236)
         );
  AOI22_X1 U4144 ( .A1(n3281), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4145 ( .A1(n4140), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4146 ( .A1(n4147), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U4147 ( .A1(n4125), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3231) );
  NAND4_X1 U4148 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n3235)
         );
  INV_X1 U4149 ( .A(n3408), .ZN(n3416) );
  NAND2_X1 U4150 ( .A1(n3250), .A2(n3416), .ZN(n3263) );
  INV_X1 U4151 ( .A(n3263), .ZN(n3249) );
  AOI22_X1 U4152 ( .A1(n3079), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4153 ( .A1(n4145), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4154 ( .A1(n3077), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4155 ( .A1(n4147), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3238) );
  NAND4_X1 U4156 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3248)
         );
  AOI22_X1 U4157 ( .A1(n3281), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4158 ( .A1(n3117), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4159 ( .A1(n4139), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4160 ( .A1(n3844), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n2953), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3243) );
  NAND4_X1 U4161 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3247)
         );
  NAND2_X1 U4162 ( .A1(n3251), .A2(n3414), .ZN(n3252) );
  NAND2_X1 U4163 ( .A1(n3253), .A2(n3252), .ZN(n3317) );
  AND2_X1 U4164 ( .A1(n3540), .A2(n6366), .ZN(n3254) );
  INV_X1 U4165 ( .A(n3316), .ZN(n3258) );
  INV_X1 U4166 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3257) );
  AOI21_X1 U4167 ( .B1(n5690), .B2(n3408), .A(n6366), .ZN(n3256) );
  NAND2_X1 U4168 ( .A1(n5662), .A2(n3319), .ZN(n3255) );
  OAI211_X1 U4169 ( .C1(n3484), .C2(n3257), .A(n3256), .B(n3255), .ZN(n3315)
         );
  NAND2_X1 U4170 ( .A1(n3258), .A2(n3315), .ZN(n3260) );
  INV_X1 U4171 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3264) );
  NAND2_X1 U4172 ( .A1(n3261), .A2(n3308), .ZN(n3262) );
  NAND2_X1 U4173 ( .A1(n3307), .A2(n3265), .ZN(n3266) );
  NAND2_X2 U4174 ( .A1(n3299), .A2(n3297), .ZN(n3330) );
  NAND2_X1 U4175 ( .A1(n3268), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3274) );
  NAND3_X1 U4176 ( .A1(n3479), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5887) );
  INV_X1 U4177 ( .A(n5887), .ZN(n3269) );
  NAND2_X1 U4178 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3269), .ZN(n5881) );
  NAND2_X1 U4179 ( .A1(n3479), .A2(n5881), .ZN(n3270) );
  NAND3_X1 U4180 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6147) );
  INV_X1 U4181 ( .A(n6147), .ZN(n6157) );
  NAND2_X1 U4182 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6157), .ZN(n6144) );
  AOI22_X1 U4183 ( .A1(n3272), .A2(n5913), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3271), .ZN(n3273) );
  AOI22_X1 U4184 ( .A1(n4146), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4185 ( .A1(n3079), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3279) );
  INV_X1 U4186 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n6520) );
  AOI22_X1 U4187 ( .A1(n3672), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4188 ( .A1(n4140), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3277) );
  NAND4_X1 U4189 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3289)
         );
  AOI22_X1 U4190 ( .A1(n3281), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4191 ( .A1(n4147), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4192 ( .A1(n3282), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4193 ( .A1(n4145), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3284) );
  NAND4_X1 U4194 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3288)
         );
  AOI22_X1 U4195 ( .A1(n3498), .A2(n3344), .B1(n3445), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3290) );
  XNOR2_X2 U4196 ( .A(n3330), .B(n4338), .ZN(n3526) );
  NAND2_X1 U4197 ( .A1(n3526), .A2(n3444), .ZN(n3296) );
  NAND2_X1 U4198 ( .A1(n3319), .A2(n3308), .ZN(n3301) );
  NAND2_X1 U4199 ( .A1(n3301), .A2(n3292), .ZN(n3345) );
  INV_X1 U4200 ( .A(n3344), .ZN(n3293) );
  XNOR2_X1 U4201 ( .A(n3345), .B(n3293), .ZN(n3294) );
  NAND2_X1 U4202 ( .A1(n3294), .A2(n6364), .ZN(n3295) );
  INV_X1 U4203 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5628) );
  INV_X1 U4204 ( .A(n3297), .ZN(n3298) );
  XNOR2_X1 U4205 ( .A(n3299), .B(n3298), .ZN(n4309) );
  XNOR2_X1 U4206 ( .A(n3301), .B(n3300), .ZN(n3302) );
  NAND2_X1 U4207 ( .A1(n5662), .A2(n3175), .ZN(n3318) );
  OAI21_X1 U4208 ( .B1(n3302), .B2(n4434), .A(n3318), .ZN(n3303) );
  AOI21_X1 U4209 ( .B1(n4309), .B2(n3444), .A(n3303), .ZN(n5539) );
  XNOR2_X1 U4210 ( .A(n3305), .B(n3304), .ZN(n3306) );
  XNOR2_X1 U4211 ( .A(n3307), .B(n3306), .ZN(n4310) );
  NAND2_X1 U4212 ( .A1(n4310), .A2(n3444), .ZN(n3314) );
  INV_X1 U4213 ( .A(n3308), .ZN(n3309) );
  XNOR2_X1 U4214 ( .A(n3309), .B(n3319), .ZN(n3312) );
  NAND3_X1 U4215 ( .A1(n3150), .A2(n3310), .A3(n3175), .ZN(n3311) );
  AOI21_X1 U4216 ( .B1(n6364), .B2(n3312), .A(n3311), .ZN(n3313) );
  NAND2_X1 U4217 ( .A1(n3314), .A2(n3313), .ZN(n4231) );
  NAND2_X1 U4218 ( .A1(n6344), .A2(n3444), .ZN(n3322) );
  OAI21_X1 U4219 ( .B1(n4434), .B2(n3319), .A(n3318), .ZN(n3320) );
  INV_X1 U4220 ( .A(n3320), .ZN(n3321) );
  NAND2_X1 U4221 ( .A1(n3322), .A2(n3321), .ZN(n5548) );
  NAND2_X1 U4222 ( .A1(n5548), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5547)
         );
  INV_X1 U4223 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4179) );
  OR2_X1 U4224 ( .A1(n5547), .A2(n4179), .ZN(n3324) );
  NAND2_X1 U4225 ( .A1(n5547), .A2(n4179), .ZN(n3323) );
  AND2_X1 U4226 ( .A1(n3324), .A2(n3323), .ZN(n4230) );
  NAND2_X1 U4227 ( .A1(n4231), .A2(n4230), .ZN(n3325) );
  NAND2_X1 U4228 ( .A1(n5538), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3327)
         );
  NAND2_X1 U4229 ( .A1(n4324), .A2(n4327), .ZN(n4325) );
  NAND2_X1 U4230 ( .A1(n3328), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3329)
         );
  NAND2_X1 U4231 ( .A1(n4325), .A2(n3329), .ZN(n5529) );
  AOI22_X1 U4232 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4272), .B1(n4120), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4233 ( .A1(n3672), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4234 ( .A1(n4146), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4235 ( .A1(n3079), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3332) );
  NAND4_X1 U4236 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3341)
         );
  AOI22_X1 U4237 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3281), .B1(n4147), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4238 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4125), .B1(n4635), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4239 ( .A1(n4139), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4240 ( .A1(n4140), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3336) );
  NAND4_X1 U4241 ( .A1(n3339), .A2(n3338), .A3(n3337), .A4(n3336), .ZN(n3340)
         );
  NAND2_X1 U4242 ( .A1(n3498), .A2(n3392), .ZN(n3343) );
  NAND2_X1 U4243 ( .A1(n3445), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3342) );
  NAND2_X1 U4244 ( .A1(n3343), .A2(n3342), .ZN(n3373) );
  NAND2_X1 U4245 ( .A1(n3345), .A2(n3344), .ZN(n3394) );
  XNOR2_X1 U4246 ( .A(n3394), .B(n3392), .ZN(n3346) );
  NAND2_X1 U4247 ( .A1(n3346), .A2(n6364), .ZN(n3347) );
  NAND2_X1 U4248 ( .A1(n3348), .A2(n3347), .ZN(n3349) );
  INV_X1 U4249 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5620) );
  XNOR2_X1 U4250 ( .A(n3349), .B(n5620), .ZN(n5528) );
  NAND2_X1 U4251 ( .A1(n5529), .A2(n5528), .ZN(n5527) );
  NAND2_X1 U4252 ( .A1(n3349), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3350)
         );
  NAND2_X1 U4253 ( .A1(n5527), .A2(n3350), .ZN(n4367) );
  NAND2_X1 U4254 ( .A1(n3374), .A2(n3373), .ZN(n3364) );
  AOI22_X1 U4255 ( .A1(n3079), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4256 ( .A1(n4146), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4257 ( .A1(n4120), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n2966), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4258 ( .A1(n3672), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3352) );
  NAND4_X1 U4259 ( .A1(n3355), .A2(n3354), .A3(n3353), .A4(n3352), .ZN(n3361)
         );
  INV_X1 U4260 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6454) );
  AOI22_X1 U4261 ( .A1(n4147), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4262 ( .A1(n3281), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4263 ( .A1(n3912), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4264 ( .A1(n4125), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3356) );
  NAND4_X1 U4265 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3360)
         );
  NAND2_X1 U4266 ( .A1(n3498), .A2(n3391), .ZN(n3363) );
  NAND2_X1 U4267 ( .A1(n3445), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3362) );
  NAND2_X1 U4268 ( .A1(n3363), .A2(n3362), .ZN(n3372) );
  NAND2_X1 U4269 ( .A1(n3513), .A2(n3444), .ZN(n3369) );
  INV_X1 U4270 ( .A(n3392), .ZN(n3365) );
  OR2_X1 U4271 ( .A1(n3394), .A2(n3365), .ZN(n3366) );
  XNOR2_X1 U4272 ( .A(n3366), .B(n3391), .ZN(n3367) );
  NAND2_X1 U4273 ( .A1(n3367), .A2(n6364), .ZN(n3368) );
  NAND2_X1 U4274 ( .A1(n3369), .A2(n3368), .ZN(n3370) );
  INV_X1 U4275 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6456) );
  XNOR2_X1 U4276 ( .A(n3370), .B(n6456), .ZN(n4366) );
  NAND2_X1 U4277 ( .A1(n4367), .A2(n4366), .ZN(n4365) );
  NAND2_X1 U4278 ( .A1(n3370), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3371)
         );
  NAND2_X1 U4279 ( .A1(n4365), .A2(n3371), .ZN(n4374) );
  NAND2_X1 U4280 ( .A1(n3374), .A2(n3021), .ZN(n3390) );
  INV_X1 U4281 ( .A(n3390), .ZN(n3388) );
  AOI22_X1 U4282 ( .A1(n3079), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4283 ( .A1(n4146), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4284 ( .A1(n4120), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4285 ( .A1(n3672), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3375) );
  NAND4_X1 U4286 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3384)
         );
  AOI22_X1 U4287 ( .A1(n3118), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4288 ( .A1(n3281), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4289 ( .A1(n3912), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4290 ( .A1(n4125), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3379) );
  NAND4_X1 U4291 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3383)
         );
  NAND2_X1 U4292 ( .A1(n3498), .A2(n3406), .ZN(n3386) );
  NAND2_X1 U4293 ( .A1(n3445), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3385) );
  INV_X1 U4294 ( .A(n3389), .ZN(n3387) );
  NAND2_X1 U4295 ( .A1(n3390), .A2(n3389), .ZN(n3523) );
  NAND3_X1 U4296 ( .A1(n3404), .A2(n3444), .A3(n3523), .ZN(n3397) );
  NAND2_X1 U4297 ( .A1(n3392), .A2(n3391), .ZN(n3393) );
  OR2_X1 U4298 ( .A1(n3394), .A2(n3393), .ZN(n3405) );
  XNOR2_X1 U4299 ( .A(n3405), .B(n3406), .ZN(n3395) );
  NAND2_X1 U4300 ( .A1(n3395), .A2(n6364), .ZN(n3396) );
  NAND2_X1 U4301 ( .A1(n3397), .A2(n3396), .ZN(n3399) );
  INV_X1 U4302 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3398) );
  XNOR2_X1 U4303 ( .A(n3399), .B(n3398), .ZN(n4373) );
  NAND2_X1 U4304 ( .A1(n4374), .A2(n4373), .ZN(n4372) );
  NAND2_X1 U4305 ( .A1(n3399), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3400)
         );
  INV_X1 U4306 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4307 ( .A1(n3498), .A2(n3408), .ZN(n3401) );
  NAND2_X1 U4308 ( .A1(n3512), .A2(n3444), .ZN(n3411) );
  INV_X1 U4309 ( .A(n3405), .ZN(n3407) );
  NAND2_X1 U4310 ( .A1(n3407), .A2(n3406), .ZN(n3417) );
  XNOR2_X1 U4311 ( .A(n3417), .B(n3408), .ZN(n3409) );
  NAND2_X1 U4312 ( .A1(n3409), .A2(n6364), .ZN(n3410) );
  NAND2_X1 U4313 ( .A1(n3411), .A2(n3410), .ZN(n3412) );
  INV_X1 U4314 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6482) );
  XNOR2_X1 U4315 ( .A(n3412), .B(n6482), .ZN(n4404) );
  NAND2_X1 U4316 ( .A1(n4405), .A2(n4404), .ZN(n4403) );
  NAND2_X1 U4317 ( .A1(n3412), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3413)
         );
  NAND2_X4 U4318 ( .A1(n3404), .A2(n3415), .ZN(n5203) );
  OR3_X1 U4319 ( .A1(n3417), .A2(n3416), .A3(n4434), .ZN(n3418) );
  NAND2_X1 U4320 ( .A1(n5203), .A2(n3418), .ZN(n3419) );
  INV_X1 U4321 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5592) );
  XNOR2_X1 U4322 ( .A(n3419), .B(n5592), .ZN(n4470) );
  NAND2_X1 U4323 ( .A1(n3419), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3420)
         );
  INV_X1 U4324 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U4325 ( .A1(n5203), .A2(n5565), .ZN(n4541) );
  OR2_X1 U4326 ( .A1(n5203), .A2(n5565), .ZN(n4542) );
  INV_X1 U4327 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3421) );
  NAND2_X1 U4328 ( .A1(n5203), .A2(n3421), .ZN(n4559) );
  INV_X1 U4329 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3422) );
  AND2_X1 U4330 ( .A1(n5203), .A2(n3422), .ZN(n3426) );
  OR2_X1 U4331 ( .A1(n5203), .A2(n3421), .ZN(n5513) );
  INV_X1 U4332 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4011) );
  NOR2_X1 U4333 ( .A1(n5203), .A2(n4011), .ZN(n4584) );
  NAND2_X1 U4334 ( .A1(n5203), .A2(n4011), .ZN(n4582) );
  XNOR2_X1 U4335 ( .A(n5203), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5218)
         );
  NAND2_X1 U4336 ( .A1(n5217), .A2(n5218), .ZN(n3429) );
  INV_X1 U4337 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3427) );
  NAND2_X1 U4338 ( .A1(n5203), .A2(n3427), .ZN(n3428) );
  NAND2_X1 U4339 ( .A1(n3429), .A2(n3428), .ZN(n4624) );
  INV_X1 U4340 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4625) );
  AND2_X1 U4341 ( .A1(n5203), .A2(n4625), .ZN(n3431) );
  OAI21_X2 U4342 ( .B1(n4624), .B2(n3431), .A(n3430), .ZN(n4989) );
  INV_X1 U4343 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5240) );
  NOR2_X1 U4344 ( .A1(n5203), .A2(n5240), .ZN(n3433) );
  NAND2_X1 U4345 ( .A1(n5203), .A2(n5240), .ZN(n3432) );
  AND2_X1 U4346 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U4347 ( .A1(n5078), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3434) );
  INV_X1 U4348 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5228) );
  INV_X1 U4349 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5223) );
  INV_X1 U4350 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6497) );
  AND3_X1 U4351 ( .A1(n5228), .A2(n5223), .A3(n6497), .ZN(n3435) );
  NAND2_X1 U4352 ( .A1(n4975), .A2(n6476), .ZN(n4935) );
  NOR2_X1 U4353 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5061) );
  INV_X1 U4354 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5044) );
  INV_X1 U4355 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5086) );
  INV_X1 U4356 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5053) );
  NAND4_X1 U4357 ( .A1(n5061), .A2(n5044), .A3(n5086), .A4(n5053), .ZN(n3437)
         );
  NAND2_X1 U4358 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U4359 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5042) );
  NOR2_X1 U4360 ( .A1(n5091), .A2(n5042), .ZN(n4945) );
  AND2_X1 U4361 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4101) );
  NAND2_X1 U4362 ( .A1(n4945), .A2(n4101), .ZN(n5027) );
  XNOR2_X1 U4363 ( .A(n5203), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4931)
         );
  NAND2_X1 U4364 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4919) );
  NOR2_X2 U4365 ( .A1(n4676), .A2(n4919), .ZN(n3937) );
  INV_X1 U4366 ( .A(n4920), .ZN(n3441) );
  NAND3_X1 U4367 ( .A1(n3440), .A2(n3441), .A3(n3438), .ZN(n4911) );
  INV_X1 U4368 ( .A(n4911), .ZN(n3442) );
  XNOR2_X1 U4369 ( .A(n3443), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5017)
         );
  AND2_X1 U4370 ( .A1(n3024), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3446)
         );
  NOR2_X1 U4371 ( .A1(n3465), .A2(n3446), .ZN(n3452) );
  NAND2_X1 U4372 ( .A1(n3498), .A2(n3452), .ZN(n3447) );
  NAND2_X1 U4373 ( .A1(n3494), .A2(n3447), .ZN(n3457) );
  INV_X1 U4374 ( .A(n3448), .ZN(n3449) );
  NAND2_X1 U4375 ( .A1(n3160), .A2(n3310), .ZN(n3450) );
  NAND2_X1 U4376 ( .A1(n3451), .A2(n3452), .ZN(n3454) );
  NAND2_X1 U4377 ( .A1(n3454), .A2(n3453), .ZN(n3455) );
  NAND2_X1 U4378 ( .A1(n3468), .A2(n3455), .ZN(n3456) );
  NAND2_X1 U4379 ( .A1(n3457), .A2(n3456), .ZN(n3461) );
  AOI21_X1 U4380 ( .B1(n3498), .B2(n4092), .A(n3146), .ZN(n3460) );
  XNOR2_X1 U4381 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3464) );
  INV_X1 U4382 ( .A(n3464), .ZN(n3458) );
  XNOR2_X1 U4383 ( .A(n3458), .B(n3465), .ZN(n3955) );
  OAI22_X1 U4384 ( .A1(n3461), .A2(n3460), .B1(n3494), .B2(n3955), .ZN(n3463)
         );
  NAND2_X1 U4385 ( .A1(n3955), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3459) );
  AOI21_X1 U4386 ( .B1(n3461), .B2(n3460), .A(n3459), .ZN(n3462) );
  NAND2_X1 U4387 ( .A1(n3465), .A2(n3464), .ZN(n3467) );
  NAND2_X1 U4388 ( .A1(n6218), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3466) );
  NAND2_X1 U4389 ( .A1(n3467), .A2(n3466), .ZN(n3475) );
  XNOR2_X1 U4390 ( .A(n2982), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3473)
         );
  XNOR2_X1 U4391 ( .A(n3475), .B(n3473), .ZN(n3954) );
  NAND2_X1 U4392 ( .A1(n3498), .A2(n3954), .ZN(n3469) );
  OAI211_X1 U4393 ( .C1(n3954), .C2(n3484), .A(n3469), .B(n3468), .ZN(n3471)
         );
  NOR2_X1 U4394 ( .A1(n3469), .A2(n3468), .ZN(n3470) );
  INV_X1 U4395 ( .A(n3473), .ZN(n3474) );
  NAND2_X1 U4396 ( .A1(n3475), .A2(n3474), .ZN(n3477) );
  NAND2_X1 U4397 ( .A1(n6213), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3476) );
  NAND2_X1 U4398 ( .A1(n3477), .A2(n3476), .ZN(n3483) );
  MUX2_X1 U4399 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n3479), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n3482) );
  INV_X1 U4400 ( .A(n3482), .ZN(n3478) );
  NAND2_X1 U4401 ( .A1(n3483), .A2(n3478), .ZN(n3481) );
  NAND2_X1 U4402 ( .A1(n3479), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U4403 ( .A1(n3481), .A2(n3480), .ZN(n3491) );
  NAND2_X1 U4404 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4299), .ZN(n3492) );
  OR2_X1 U4405 ( .A1(n3491), .A2(n3492), .ZN(n3958) );
  XNOR2_X1 U4406 ( .A(n3483), .B(n3482), .ZN(n3953) );
  NAND2_X1 U4407 ( .A1(n3958), .A2(n3953), .ZN(n3485) );
  INV_X1 U4408 ( .A(n3494), .ZN(n3486) );
  AOI22_X1 U4409 ( .A1(n3486), .A2(n3485), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6366), .ZN(n3487) );
  INV_X1 U4410 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n5656) );
  AND2_X1 U4411 ( .A1(n5656), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3490)
         );
  INV_X1 U4412 ( .A(n3957), .ZN(n3497) );
  NAND2_X1 U4413 ( .A1(n4072), .A2(n2961), .ZN(n3503) );
  NAND2_X1 U4414 ( .A1(n4185), .A2(n5662), .ZN(n3504) );
  NAND2_X1 U4415 ( .A1(n4079), .A2(n3504), .ZN(n3969) );
  OR2_X1 U4416 ( .A1(n3969), .A2(n3451), .ZN(n6226) );
  NAND2_X1 U4417 ( .A1(n5017), .A2(n5541), .ZN(n3936) );
  NOR2_X2 U4418 ( .A1(n2961), .A2(n3558), .ZN(n3506) );
  INV_X1 U4419 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3510) );
  XNOR2_X1 U4420 ( .A(n3578), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4478) );
  NAND2_X1 U4421 ( .A1(n4478), .A2(n4655), .ZN(n3509) );
  NAND2_X1 U4422 ( .A1(n3558), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3550) );
  NAND2_X1 U4423 ( .A1(n4658), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3508)
         );
  OAI211_X1 U4424 ( .C1(n3877), .C2(n3510), .A(n3509), .B(n3508), .ZN(n3511)
         );
  NAND2_X1 U4425 ( .A1(n3513), .A2(n3693), .ZN(n3518) );
  AND2_X1 U4426 ( .A1(n3563), .A2(n6431), .ZN(n3514) );
  OR2_X1 U4427 ( .A1(n3514), .A2(n3519), .ZN(n4527) );
  NAND2_X1 U4428 ( .A1(n4527), .A2(n4655), .ZN(n3515) );
  OAI21_X1 U4429 ( .B1(n6431), .B2(n3550), .A(n3515), .ZN(n3516) );
  AOI21_X1 U4430 ( .B1(n3506), .B2(EAX_REG_5__SCAN_IN), .A(n3516), .ZN(n3517)
         );
  INV_X1 U4431 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4389) );
  NOR2_X1 U4432 ( .A1(n3519), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3520)
         );
  OR2_X1 U4433 ( .A1(n3578), .A2(n3520), .ZN(n5526) );
  AOI22_X1 U4434 ( .A1(n5526), .A2(n4655), .B1(n4658), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3521) );
  OAI21_X1 U4435 ( .B1(n3877), .B2(n4389), .A(n3521), .ZN(n3522) );
  INV_X1 U4436 ( .A(n4399), .ZN(n3524) );
  NAND2_X1 U4437 ( .A1(n4361), .A2(n3524), .ZN(n3525) );
  NOR2_X2 U4438 ( .A1(n4398), .A2(n3525), .ZN(n4391) );
  INV_X1 U4439 ( .A(n3547), .ZN(n3561) );
  INV_X1 U4440 ( .A(n3564), .ZN(n3528) );
  INV_X1 U4441 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U4442 ( .A1(n4501), .A2(n3548), .ZN(n3527) );
  NAND2_X1 U4443 ( .A1(n3528), .A2(n3527), .ZN(n4500) );
  AOI22_X1 U4444 ( .A1(n4500), .A2(n4655), .B1(n4658), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3530) );
  NAND2_X1 U4445 ( .A1(n4659), .A2(EAX_REG_3__SCAN_IN), .ZN(n3529) );
  OAI211_X1 U4446 ( .C1(n3561), .C2(n3023), .A(n3530), .B(n3529), .ZN(n3531)
         );
  INV_X1 U4447 ( .A(n4328), .ZN(n3557) );
  NAND2_X1 U4448 ( .A1(n4309), .A2(n3693), .ZN(n3532) );
  NAND2_X1 U4449 ( .A1(n3532), .A2(n3550), .ZN(n4252) );
  NAND2_X1 U4450 ( .A1(n4310), .A2(n3693), .ZN(n3536) );
  AOI22_X1 U4451 ( .A1(n4659), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n3558), .ZN(n3534) );
  NAND2_X1 U4452 ( .A1(n3547), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3533) );
  AND2_X1 U4453 ( .A1(n3534), .A2(n3533), .ZN(n3535) );
  NAND2_X1 U4454 ( .A1(n3536), .A2(n3535), .ZN(n4217) );
  AOI21_X1 U4455 ( .B1(n6071), .B2(n3537), .A(n3558), .ZN(n4215) );
  INV_X1 U4456 ( .A(n3538), .ZN(n3541) );
  NAND3_X1 U4457 ( .A1(n3541), .A2(n3540), .A3(n3539), .ZN(n3542) );
  NAND2_X1 U4458 ( .A1(n2962), .A2(n3542), .ZN(n5948) );
  INV_X1 U4459 ( .A(n3693), .ZN(n3683) );
  OR2_X1 U4460 ( .A1(n5948), .A2(n3683), .ZN(n3546) );
  AOI22_X1 U4461 ( .A1(n4659), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n3558), .ZN(n3544) );
  NAND2_X1 U4462 ( .A1(n3547), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3543) );
  AND2_X1 U4463 ( .A1(n3544), .A2(n3543), .ZN(n3545) );
  NAND2_X1 U4464 ( .A1(n3546), .A2(n3545), .ZN(n4214) );
  MUX2_X1 U4465 ( .A(n4419), .B(n4215), .S(n4214), .Z(n4216) );
  NAND2_X1 U4466 ( .A1(n4217), .A2(n4216), .ZN(n4219) );
  NAND2_X1 U4467 ( .A1(n3547), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3553) );
  INV_X1 U4468 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4492) );
  OAI21_X1 U4469 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3548), .ZN(n5545) );
  NAND2_X1 U4470 ( .A1(n4419), .A2(n5545), .ZN(n3549) );
  OAI21_X1 U4471 ( .B1(n3550), .B2(n4492), .A(n3549), .ZN(n3551) );
  AOI21_X1 U4472 ( .B1(n4659), .B2(EAX_REG_2__SCAN_IN), .A(n3551), .ZN(n3552)
         );
  AND2_X1 U4473 ( .A1(n3553), .A2(n3552), .ZN(n3554) );
  NOR2_X1 U4474 ( .A1(n4219), .A2(n3554), .ZN(n3555) );
  NAND2_X1 U4475 ( .A1(n4219), .A2(n3554), .ZN(n4253) );
  OAI21_X1 U4476 ( .B1(n4252), .B2(n3555), .A(n4253), .ZN(n4251) );
  INV_X1 U4477 ( .A(n4251), .ZN(n3556) );
  NAND2_X1 U4478 ( .A1(n3558), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3560)
         );
  NAND2_X1 U4479 ( .A1(n3506), .A2(EAX_REG_4__SCAN_IN), .ZN(n3559) );
  OAI211_X1 U4480 ( .C1(n3561), .C2(n4299), .A(n3560), .B(n3559), .ZN(n3562)
         );
  NAND2_X1 U4481 ( .A1(n3562), .A2(n4649), .ZN(n3566) );
  OAI21_X1 U4482 ( .B1(n3564), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3563), 
        .ZN(n5535) );
  NAND2_X1 U4483 ( .A1(n5535), .A2(n4655), .ZN(n3565) );
  NAND2_X1 U4484 ( .A1(n3566), .A2(n3565), .ZN(n3567) );
  AOI22_X1 U4485 ( .A1(n3672), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4486 ( .A1(n3118), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4487 ( .A1(n4140), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4488 ( .A1(n3281), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3568) );
  NAND4_X1 U4489 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(n3577)
         );
  AOI22_X1 U4490 ( .A1(n4272), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4491 ( .A1(n4145), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4492 ( .A1(n3079), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4493 ( .A1(n4146), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3572) );
  NAND4_X1 U4494 ( .A1(n3575), .A2(n3574), .A3(n3573), .A4(n3572), .ZN(n3576)
         );
  OAI21_X1 U4495 ( .B1(n3577), .B2(n3576), .A(n3693), .ZN(n3582) );
  NAND2_X1 U4496 ( .A1(n3506), .A2(EAX_REG_8__SCAN_IN), .ZN(n3581) );
  XNOR2_X1 U4497 ( .A(n3583), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4472) );
  NAND2_X1 U4498 ( .A1(n4472), .A2(n4655), .ZN(n3580) );
  NAND2_X1 U4499 ( .A1(n4658), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3579)
         );
  NAND4_X1 U4500 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n4411)
         );
  XNOR2_X1 U4501 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3598), .ZN(n5339) );
  AOI22_X1 U4502 ( .A1(n4147), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4503 ( .A1(n4120), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4504 ( .A1(n3912), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4505 ( .A1(n3079), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3584) );
  NAND4_X1 U4506 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(n3593)
         );
  AOI22_X1 U4507 ( .A1(n4146), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4508 ( .A1(n3672), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4509 ( .A1(n3281), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4510 ( .A1(n4145), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3588) );
  NAND4_X1 U4511 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3592)
         );
  OR2_X1 U4512 ( .A1(n3593), .A2(n3592), .ZN(n3594) );
  AOI22_X1 U4513 ( .A1(n3693), .A2(n3594), .B1(n4658), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4514 ( .A1(n3506), .A2(EAX_REG_9__SCAN_IN), .ZN(n3595) );
  OAI211_X1 U4515 ( .C1(n5339), .C2(n4649), .A(n3596), .B(n3595), .ZN(n4393)
         );
  XNOR2_X1 U4516 ( .A(n3614), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4561)
         );
  AOI22_X1 U4517 ( .A1(n3079), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4518 ( .A1(n3672), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4519 ( .A1(n4146), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4520 ( .A1(n4120), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4521 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3608)
         );
  AOI22_X1 U4522 ( .A1(n4147), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3606) );
  AOI22_X1 U4523 ( .A1(n3281), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4524 ( .A1(n3844), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4525 ( .A1(n4125), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3603) );
  NAND4_X1 U4526 ( .A1(n3606), .A2(n3605), .A3(n3604), .A4(n3603), .ZN(n3607)
         );
  OAI21_X1 U4527 ( .B1(n3608), .B2(n3607), .A(n3693), .ZN(n3611) );
  NAND2_X1 U4528 ( .A1(n3506), .A2(EAX_REG_10__SCAN_IN), .ZN(n3610) );
  NAND2_X1 U4529 ( .A1(n4658), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3609)
         );
  NAND3_X1 U4530 ( .A1(n3611), .A2(n3610), .A3(n3609), .ZN(n3612) );
  AOI21_X1 U4531 ( .B1(n4561), .B2(n4655), .A(n3612), .ZN(n4416) );
  XNOR2_X1 U4532 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3631), .ZN(n5516)
         );
  INV_X1 U4533 ( .A(n5516), .ZN(n3629) );
  AOI22_X1 U4534 ( .A1(n3079), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4535 ( .A1(n3281), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4536 ( .A1(n4145), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4537 ( .A1(n4147), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3615) );
  NAND4_X1 U4538 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3624)
         );
  AOI22_X1 U4539 ( .A1(n3672), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4540 ( .A1(n4146), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4541 ( .A1(n4140), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4542 ( .A1(n3912), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4543 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3623)
         );
  OAI21_X1 U4544 ( .B1(n3624), .B2(n3623), .A(n3693), .ZN(n3627) );
  NAND2_X1 U4545 ( .A1(n3506), .A2(EAX_REG_11__SCAN_IN), .ZN(n3626) );
  NAND2_X1 U4546 ( .A1(n4658), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3625)
         );
  NAND3_X1 U4547 ( .A1(n3627), .A2(n3626), .A3(n3625), .ZN(n3628) );
  AOI21_X1 U4548 ( .B1(n3629), .B2(n4655), .A(n3628), .ZN(n4519) );
  XNOR2_X1 U4549 ( .A(n3646), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4588)
         );
  INV_X1 U4550 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4551) );
  AOI21_X1 U4551 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n4551), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3633) );
  AND2_X1 U4552 ( .A1(n3506), .A2(EAX_REG_12__SCAN_IN), .ZN(n3632) );
  OAI22_X1 U4553 ( .A1(n4588), .A2(n4649), .B1(n3633), .B2(n3632), .ZN(n3645)
         );
  AOI22_X1 U4554 ( .A1(n4146), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4555 ( .A1(n4120), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4556 ( .A1(n4145), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4557 ( .A1(n4140), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4558 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3643)
         );
  AOI22_X1 U4559 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3079), .B1(n3672), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4560 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4272), .B1(n4147), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4561 ( .A1(n3912), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4562 ( .A1(n3281), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4563 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3642)
         );
  OAI21_X1 U4564 ( .B1(n3643), .B2(n3642), .A(n3693), .ZN(n3644) );
  NAND2_X1 U4565 ( .A1(n4518), .A2(n4535), .ZN(n3653) );
  INV_X1 U4566 ( .A(n3653), .ZN(n3650) );
  NAND2_X1 U4567 ( .A1(n4659), .A2(EAX_REG_13__SCAN_IN), .ZN(n3649) );
  OAI21_X1 U4568 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3647), .A(n3684), 
        .ZN(n5320) );
  AOI22_X1 U4569 ( .A1(n4419), .A2(n5320), .B1(n4658), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3648) );
  NAND2_X1 U4570 ( .A1(n3649), .A2(n3648), .ZN(n3651) );
  INV_X1 U4571 ( .A(n3651), .ZN(n3652) );
  NAND2_X1 U4572 ( .A1(n3653), .A2(n3652), .ZN(n3654) );
  AOI22_X1 U4573 ( .A1(n3281), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4574 ( .A1(n4147), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4575 ( .A1(n3079), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4576 ( .A1(n4140), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3655) );
  NAND4_X1 U4577 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(n3664)
         );
  AOI22_X1 U4578 ( .A1(n3672), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4579 ( .A1(n4125), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4580 ( .A1(n3912), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4581 ( .A1(n4146), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3659) );
  NAND4_X1 U4582 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3663)
         );
  OR2_X1 U4583 ( .A1(n3664), .A2(n3663), .ZN(n3665) );
  NAND2_X1 U4584 ( .A1(n3693), .A2(n3665), .ZN(n4567) );
  AOI22_X1 U4585 ( .A1(n3079), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4586 ( .A1(n4147), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4587 ( .A1(n4120), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4588 ( .A1(n3844), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3668) );
  NAND4_X1 U4589 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(n3678)
         );
  AOI22_X1 U4590 ( .A1(n4146), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3672), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4591 ( .A1(n3281), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3675) );
  AOI22_X1 U4592 ( .A1(n4272), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4593 ( .A1(n4140), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3673) );
  NAND4_X1 U4594 ( .A1(n3676), .A2(n3675), .A3(n3674), .A4(n3673), .ZN(n3677)
         );
  NOR2_X1 U4595 ( .A1(n3678), .A2(n3677), .ZN(n3682) );
  XNOR2_X1 U4596 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3684), .ZN(n5307)
         );
  INV_X1 U4597 ( .A(n5307), .ZN(n3679) );
  AOI22_X1 U4598 ( .A1(n4658), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n4419), 
        .B2(n3679), .ZN(n3681) );
  NAND2_X1 U4599 ( .A1(n4659), .A2(EAX_REG_14__SCAN_IN), .ZN(n3680) );
  OAI211_X1 U4600 ( .C1(n3683), .C2(n3682), .A(n3681), .B(n3680), .ZN(n4574)
         );
  NAND2_X1 U4601 ( .A1(n4573), .A2(n4574), .ZN(n4572) );
  XNOR2_X1 U4602 ( .A(n3700), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4992)
         );
  AOI22_X1 U4603 ( .A1(n4659), .A2(EAX_REG_15__SCAN_IN), .B1(n4658), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4604 ( .A1(n3281), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4147), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4605 ( .A1(n3672), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4606 ( .A1(n4145), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4607 ( .A1(n3844), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3685) );
  NAND4_X1 U4608 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3695)
         );
  AOI22_X1 U4609 ( .A1(n3079), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4610 ( .A1(n3912), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4611 ( .A1(n4272), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4612 ( .A1(n4146), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3689) );
  NAND4_X1 U4613 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3694)
         );
  OAI21_X1 U4614 ( .B1(n3695), .B2(n3694), .A(n3693), .ZN(n3696) );
  OAI211_X1 U4615 ( .C1(n4992), .C2(n4649), .A(n3697), .B(n3696), .ZN(n4604)
         );
  XOR2_X1 U4616 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3713), .Z(n4986) );
  AOI22_X1 U4617 ( .A1(n4659), .A2(EAX_REG_16__SCAN_IN), .B1(n4658), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4618 ( .A1(n3281), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4619 ( .A1(n4147), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4620 ( .A1(n4120), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4621 ( .A1(n3079), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3701) );
  NAND4_X1 U4622 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3710)
         );
  AOI22_X1 U4623 ( .A1(n3672), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4624 ( .A1(n4272), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4625 ( .A1(n4145), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4626 ( .A1(n4146), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3705) );
  NAND4_X1 U4627 ( .A1(n3708), .A2(n3707), .A3(n3706), .A4(n3705), .ZN(n3709)
         );
  OAI21_X1 U4628 ( .B1(n3710), .B2(n3709), .A(n4154), .ZN(n3711) );
  OAI211_X1 U4629 ( .C1(n4986), .C2(n4649), .A(n3712), .B(n3711), .ZN(n4808)
         );
  XNOR2_X1 U4630 ( .A(n3728), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5214)
         );
  AOI22_X1 U4631 ( .A1(n4659), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3558), .ZN(n3727) );
  AOI22_X1 U4632 ( .A1(n3672), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4633 ( .A1(n3281), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4634 ( .A1(n4272), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4635 ( .A1(n4140), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3714) );
  NAND4_X1 U4636 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3725)
         );
  AOI22_X1 U4637 ( .A1(n4146), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4638 ( .A1(n3079), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3722) );
  NAND2_X1 U4639 ( .A1(n4147), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3719) );
  AOI21_X1 U4640 ( .B1(n2967), .B2(INSTQUEUE_REG_9__1__SCAN_IN), .A(n4655), 
        .ZN(n3718) );
  AND2_X1 U4641 ( .A1(n3719), .A2(n3718), .ZN(n3721) );
  AOI22_X1 U4642 ( .A1(n4145), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3720) );
  NAND4_X1 U4643 ( .A1(n3723), .A2(n3722), .A3(n3721), .A4(n3720), .ZN(n3724)
         );
  NAND2_X1 U4644 ( .A1(n4652), .A2(n4649), .ZN(n3788) );
  OAI21_X1 U4645 ( .B1(n3725), .B2(n3724), .A(n3788), .ZN(n3726) );
  AOI22_X1 U4646 ( .A1(n5214), .A2(n4655), .B1(n3727), .B2(n3726), .ZN(n4796)
         );
  INV_X1 U4647 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4803) );
  INV_X1 U4648 ( .A(n3760), .ZN(n3731) );
  OR2_X1 U4649 ( .A1(n3729), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3730)
         );
  NAND2_X1 U4650 ( .A1(n3731), .A2(n3730), .ZN(n5301) );
  AOI22_X1 U4651 ( .A1(n4147), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4652 ( .A1(n3079), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4653 ( .A1(n3672), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4654 ( .A1(n4140), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4655 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3741)
         );
  AOI22_X1 U4656 ( .A1(n4120), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4657 ( .A1(n4146), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4658 ( .A1(n3912), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4659 ( .A1(n3281), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4660 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  NOR2_X1 U4661 ( .A1(n3741), .A2(n3740), .ZN(n3744) );
  INV_X1 U4662 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6363) );
  OAI21_X1 U4663 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6363), .A(n3558), 
        .ZN(n3743) );
  NAND2_X1 U4664 ( .A1(n4659), .A2(EAX_REG_18__SCAN_IN), .ZN(n3742) );
  OAI211_X1 U4665 ( .C1(n4652), .C2(n3744), .A(n3743), .B(n3742), .ZN(n3745)
         );
  OAI21_X1 U4666 ( .B1(n5301), .B2(n4649), .A(n3745), .ZN(n4879) );
  INV_X1 U4667 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4977) );
  XNOR2_X1 U4668 ( .A(n3760), .B(n4977), .ZN(n4981) );
  AOI22_X1 U4669 ( .A1(n4659), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3558), .ZN(n3759) );
  AOI22_X1 U4670 ( .A1(n3079), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4671 ( .A1(n3281), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4147), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4672 ( .A1(n4145), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4673 ( .A1(n4125), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3746) );
  NAND4_X1 U4674 ( .A1(n3749), .A2(n3748), .A3(n3747), .A4(n3746), .ZN(n3757)
         );
  AOI22_X1 U4675 ( .A1(n4146), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4676 ( .A1(n3912), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4677 ( .A1(n3672), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3753) );
  NAND2_X1 U4678 ( .A1(n4272), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3751)
         );
  AOI21_X1 U4679 ( .B1(n2967), .B2(INSTQUEUE_REG_9__3__SCAN_IN), .A(n4655), 
        .ZN(n3750) );
  AND2_X1 U4680 ( .A1(n3751), .A2(n3750), .ZN(n3752) );
  NAND4_X1 U4681 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3756)
         );
  OAI21_X1 U4682 ( .B1(n3757), .B2(n3756), .A(n3788), .ZN(n3758) );
  AOI22_X1 U4683 ( .A1(n4981), .A2(n4655), .B1(n3759), .B2(n3758), .ZN(n4783)
         );
  OR2_X1 U4684 ( .A1(n3761), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3762)
         );
  NAND2_X1 U4685 ( .A1(n3762), .A2(n3793), .ZN(n5176) );
  AOI22_X1 U4686 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4146), .B1(n4125), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4687 ( .A1(n3672), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4688 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3281), .B1(n4635), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4689 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4272), .B1(n3230), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3763) );
  NAND4_X1 U4690 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3772)
         );
  AOI22_X1 U4691 ( .A1(n3079), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4692 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4147), .B1(n3844), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4693 ( .A1(n4120), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4694 ( .A1(n4140), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3767) );
  NAND4_X1 U4695 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3771)
         );
  NOR2_X1 U4696 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  NOR2_X1 U4697 ( .A1(n4652), .A2(n3773), .ZN(n3777) );
  INV_X1 U4698 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U4699 ( .A1(n3558), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3774)
         );
  OAI211_X1 U4700 ( .C1(n3877), .C2(n3775), .A(n4649), .B(n3774), .ZN(n3776)
         );
  OAI22_X1 U4701 ( .A1(n5176), .A2(n4649), .B1(n3777), .B2(n3776), .ZN(n4867)
         );
  AOI22_X1 U4702 ( .A1(n3079), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4703 ( .A1(n3281), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4147), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4704 ( .A1(n3672), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4705 ( .A1(n4145), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4706 ( .A1(n3781), .A2(n3780), .A3(n3779), .A4(n3778), .ZN(n3790)
         );
  AOI22_X1 U4707 ( .A1(n4146), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4708 ( .A1(n4120), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4709 ( .A1(n4635), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3785) );
  NAND2_X1 U4710 ( .A1(n4272), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3783)
         );
  AOI21_X1 U4711 ( .B1(n2967), .B2(INSTQUEUE_REG_9__5__SCAN_IN), .A(n4655), 
        .ZN(n3782) );
  AND2_X1 U4712 ( .A1(n3783), .A2(n3782), .ZN(n3784) );
  NAND4_X1 U4713 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3789)
         );
  OAI21_X1 U4714 ( .B1(n3790), .B2(n3789), .A(n3788), .ZN(n3792) );
  AOI22_X1 U4715 ( .A1(n4659), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n3558), .ZN(n3791) );
  NAND2_X1 U4716 ( .A1(n3792), .A2(n3791), .ZN(n3797) );
  NOR2_X1 U4717 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3794), .ZN(n3795)
         );
  NOR2_X1 U4718 ( .A1(n3813), .A2(n3795), .ZN(n5163) );
  NAND2_X1 U4719 ( .A1(n5163), .A2(n4655), .ZN(n3796) );
  NAND2_X1 U4720 ( .A1(n3797), .A2(n3796), .ZN(n4962) );
  AOI22_X1 U4721 ( .A1(n4147), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4722 ( .A1(n4146), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4723 ( .A1(n3672), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4724 ( .A1(n4125), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3799) );
  NAND4_X1 U4725 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n3808)
         );
  AOI22_X1 U4726 ( .A1(n3281), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4727 ( .A1(n3079), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4728 ( .A1(n4140), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4729 ( .A1(n4145), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4730 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3807)
         );
  NOR2_X1 U4731 ( .A1(n3808), .A2(n3807), .ZN(n3812) );
  NAND2_X1 U4732 ( .A1(n3558), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3809)
         );
  NAND2_X1 U4733 ( .A1(n4649), .A2(n3809), .ZN(n3810) );
  AOI21_X1 U4734 ( .B1(n3506), .B2(EAX_REG_22__SCAN_IN), .A(n3810), .ZN(n3811)
         );
  OAI21_X1 U4735 ( .B1(n4652), .B2(n3812), .A(n3811), .ZN(n3815) );
  OAI21_X1 U4736 ( .B1(n3813), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n3856), 
        .ZN(n5150) );
  OR2_X1 U4737 ( .A1(n5150), .A2(n4649), .ZN(n3814) );
  AOI22_X1 U4738 ( .A1(n3079), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4739 ( .A1(n4272), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4740 ( .A1(n4140), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4741 ( .A1(n3844), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3816) );
  NAND4_X1 U4742 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3825)
         );
  AOI22_X1 U4743 ( .A1(n4120), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4744 ( .A1(n3281), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4147), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4745 ( .A1(n3672), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4746 ( .A1(n4146), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4747 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3824)
         );
  NOR2_X1 U4748 ( .A1(n3825), .A2(n3824), .ZN(n3843) );
  AOI22_X1 U4749 ( .A1(n3079), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4750 ( .A1(n3672), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4751 ( .A1(n4147), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4752 ( .A1(n4146), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3826) );
  NAND4_X1 U4753 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3835)
         );
  AOI22_X1 U4754 ( .A1(n4272), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4755 ( .A1(n3281), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4756 ( .A1(n4140), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4757 ( .A1(n4120), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4758 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3834)
         );
  NOR2_X1 U4759 ( .A1(n3835), .A2(n3834), .ZN(n3842) );
  XOR2_X1 U4760 ( .A(n3843), .B(n3842), .Z(n3836) );
  NAND2_X1 U4761 ( .A1(n3836), .A2(n4154), .ZN(n3839) );
  INV_X1 U4762 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4950) );
  AOI21_X1 U4763 ( .B1(n4950), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3837) );
  AOI21_X1 U4764 ( .B1(n3506), .B2(EAX_REG_23__SCAN_IN), .A(n3837), .ZN(n3838)
         );
  NAND2_X1 U4765 ( .A1(n3839), .A2(n3838), .ZN(n3841) );
  XNOR2_X1 U4766 ( .A(n3856), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5140)
         );
  NAND2_X1 U4767 ( .A1(n5140), .A2(n4655), .ZN(n3840) );
  NAND2_X1 U4768 ( .A1(n3841), .A2(n3840), .ZN(n4854) );
  NOR2_X1 U4769 ( .A1(n3843), .A2(n3842), .ZN(n3874) );
  AOI22_X1 U4770 ( .A1(n3079), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4771 ( .A1(n3077), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4772 ( .A1(n4120), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4773 ( .A1(n3672), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3845) );
  NAND4_X1 U4774 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3854)
         );
  AOI22_X1 U4775 ( .A1(n4147), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4776 ( .A1(n3281), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4777 ( .A1(n3912), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4778 ( .A1(n4125), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4779 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3853)
         );
  OR2_X1 U4780 ( .A1(n3854), .A2(n3853), .ZN(n3873) );
  INV_X1 U4781 ( .A(n3873), .ZN(n3855) );
  XNOR2_X1 U4782 ( .A(n3874), .B(n3855), .ZN(n3861) );
  INV_X1 U4783 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U4784 ( .A1(n4658), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3859)
         );
  INV_X1 U4785 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3857) );
  XNOR2_X1 U4786 ( .A(n3881), .B(n3857), .ZN(n5133) );
  OAI211_X1 U4787 ( .C1(n3877), .C2(n6453), .A(n3859), .B(n3858), .ZN(n3860)
         );
  AOI21_X1 U4788 ( .B1(n3861), .B2(n4154), .A(n3860), .ZN(n4848) );
  AOI22_X1 U4789 ( .A1(n3079), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4790 ( .A1(n4145), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4791 ( .A1(n4146), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4792 ( .A1(n3672), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3863) );
  NAND4_X1 U4793 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3872)
         );
  AOI22_X1 U4794 ( .A1(n4147), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4795 ( .A1(n3281), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4796 ( .A1(n3912), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4797 ( .A1(n4125), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4798 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3871)
         );
  NOR2_X1 U4799 ( .A1(n3872), .A2(n3871), .ZN(n3885) );
  NAND2_X1 U4800 ( .A1(n3874), .A2(n3873), .ZN(n3884) );
  XOR2_X1 U4801 ( .A(n3885), .B(n3884), .Z(n3879) );
  INV_X1 U4802 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3876) );
  NAND2_X1 U4803 ( .A1(n3558), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3875)
         );
  OAI211_X1 U4804 ( .C1(n3877), .C2(n3876), .A(n4649), .B(n3875), .ZN(n3878)
         );
  AOI21_X1 U4805 ( .B1(n3879), .B2(n4154), .A(n3878), .ZN(n3880) );
  INV_X1 U4806 ( .A(n3880), .ZN(n3883) );
  INV_X1 U4807 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4929) );
  XNOR2_X1 U4808 ( .A(n3900), .B(n4929), .ZN(n5125) );
  NAND2_X1 U4809 ( .A1(n5125), .A2(n4655), .ZN(n3882) );
  NAND2_X1 U4810 ( .A1(n3883), .A2(n3882), .ZN(n4837) );
  NOR2_X1 U4811 ( .A1(n3885), .A2(n3884), .ZN(n3907) );
  AOI22_X1 U4812 ( .A1(n3079), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4813 ( .A1(n3077), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4814 ( .A1(n4120), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4815 ( .A1(n3672), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3886) );
  NAND4_X1 U4816 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n3895)
         );
  AOI22_X1 U4817 ( .A1(n4147), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4818 ( .A1(n3281), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4819 ( .A1(n3912), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4820 ( .A1(n4125), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4821 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3894)
         );
  OR2_X1 U4822 ( .A1(n3895), .A2(n3894), .ZN(n3906) );
  INV_X1 U4823 ( .A(n3906), .ZN(n3896) );
  XNOR2_X1 U4824 ( .A(n3907), .B(n3896), .ZN(n3897) );
  NAND2_X1 U4825 ( .A1(n3897), .A2(n4154), .ZN(n3905) );
  NAND2_X1 U4826 ( .A1(n3558), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3898)
         );
  NAND2_X1 U4827 ( .A1(n4649), .A2(n3898), .ZN(n3899) );
  AOI21_X1 U4828 ( .B1(n3506), .B2(EAX_REG_26__SCAN_IN), .A(n3899), .ZN(n3904)
         );
  OR2_X1 U4829 ( .A1(n3901), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3902)
         );
  NAND2_X1 U4830 ( .A1(n4112), .A2(n3902), .ZN(n5123) );
  NOR2_X1 U4831 ( .A1(n5123), .A2(n4649), .ZN(n3903) );
  AOI21_X1 U4832 ( .B1(n3905), .B2(n3904), .A(n3903), .ZN(n4830) );
  NAND2_X1 U4833 ( .A1(n3907), .A2(n3906), .ZN(n4118) );
  AOI22_X1 U4834 ( .A1(n3079), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4835 ( .A1(n4145), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4836 ( .A1(n3077), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4837 ( .A1(n4272), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3908) );
  NAND4_X1 U4838 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3918)
         );
  AOI22_X1 U4839 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3281), .B1(n4125), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4840 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4147), .B1(n4635), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4841 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3912), .B1(n4139), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4842 ( .A1(n3672), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4843 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3917)
         );
  NOR2_X1 U4844 ( .A1(n3918), .A2(n3917), .ZN(n4119) );
  XOR2_X1 U4845 ( .A(n4118), .B(n4119), .Z(n3919) );
  NAND2_X1 U4846 ( .A1(n3919), .A2(n4154), .ZN(n3922) );
  INV_X1 U4847 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3931) );
  NOR2_X1 U4848 ( .A1(n3931), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3920) );
  AOI211_X1 U4849 ( .C1(n3506), .C2(EAX_REG_27__SCAN_IN), .A(n4655), .B(n3920), 
        .ZN(n3921) );
  XNOR2_X1 U4850 ( .A(n4112), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4769)
         );
  AND2_X1 U4851 ( .A1(n6366), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4420) );
  NAND2_X1 U4852 ( .A1(n4420), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6260) );
  NOR2_X2 U4853 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6345) );
  OR2_X2 U4854 ( .A1(n6260), .A2(n6370), .ZN(n5692) );
  NAND2_X1 U4855 ( .A1(n6370), .A2(n6369), .ZN(n3925) );
  NAND2_X1 U4856 ( .A1(n3925), .A2(n6366), .ZN(n3926) );
  NAND2_X1 U4857 ( .A1(n6366), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3928) );
  NAND2_X1 U4858 ( .A1(n6363), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3927) );
  AND2_X1 U4859 ( .A1(n3928), .A2(n3927), .ZN(n5551) );
  INV_X1 U4860 ( .A(n5551), .ZN(n3929) );
  NAND2_X1 U4861 ( .A1(n6345), .A2(n6425), .ZN(n5115) );
  INV_X1 U4862 ( .A(REIP_REG_27__SCAN_IN), .ZN(n3930) );
  NOR2_X1 U4863 ( .A1(n5612), .A2(n3930), .ZN(n5020) );
  NOR2_X1 U4864 ( .A1(n5550), .A2(n3931), .ZN(n3932) );
  AOI211_X1 U4865 ( .C1(n5517), .C2(n4769), .A(n5020), .B(n3932), .ZN(n3933)
         );
  AND2_X1 U4866 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5003) );
  INV_X1 U4867 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5002) );
  INV_X1 U4868 ( .A(n3939), .ZN(n3943) );
  INV_X1 U4869 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3941) );
  INV_X1 U4870 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3940) );
  NAND2_X1 U4871 ( .A1(n3941), .A2(n3940), .ZN(n5012) );
  NOR2_X1 U4872 ( .A1(n4920), .A2(n5012), .ZN(n4110) );
  NAND2_X1 U4873 ( .A1(n4110), .A2(n5002), .ZN(n4674) );
  NOR2_X1 U4874 ( .A1(n4674), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3942)
         );
  AOI21_X1 U4875 ( .B1(n4677), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n3944), 
        .ZN(n3946) );
  XNOR2_X1 U4876 ( .A(n3946), .B(n3945), .ZN(n4707) );
  INV_X1 U4877 ( .A(n4185), .ZN(n6214) );
  NAND2_X1 U4878 ( .A1(n6214), .A2(n4092), .ZN(n4084) );
  INV_X1 U4879 ( .A(n4084), .ZN(n3947) );
  NAND2_X1 U4880 ( .A1(n4199), .A2(n3947), .ZN(n3961) );
  INV_X1 U4881 ( .A(n3948), .ZN(n3951) );
  NAND2_X1 U4882 ( .A1(n4076), .A2(n4074), .ZN(n3949) );
  OR2_X1 U4883 ( .A1(n3969), .A2(n3949), .ZN(n3950) );
  NAND2_X1 U4884 ( .A1(n3951), .A2(n3950), .ZN(n4195) );
  NAND2_X1 U4885 ( .A1(n3952), .A2(n6523), .ZN(n6266) );
  NAND2_X1 U4886 ( .A1(n4092), .A2(n6266), .ZN(n4167) );
  NAND3_X1 U4887 ( .A1(n3955), .A2(n3954), .A3(n3953), .ZN(n3956) );
  NAND2_X1 U4888 ( .A1(n3957), .A2(n3956), .ZN(n3959) );
  NOR2_X1 U4889 ( .A1(n4168), .A2(READY_N), .ZN(n4190) );
  NAND3_X1 U4890 ( .A1(n4167), .A2(n4190), .A3(n3142), .ZN(n3960) );
  NAND3_X1 U4891 ( .A1(n3961), .A2(n4195), .A3(n3960), .ZN(n3962) );
  NAND2_X1 U4892 ( .A1(n3962), .A2(n6251), .ZN(n3968) );
  INV_X1 U4893 ( .A(n6266), .ZN(n4431) );
  INV_X1 U4894 ( .A(READY_N), .ZN(n6271) );
  OAI21_X1 U4895 ( .B1(n4092), .B2(n4431), .A(n6271), .ZN(n4428) );
  OAI211_X1 U4896 ( .C1(n3964), .C2(n4428), .A(n3178), .B(n4661), .ZN(n3965)
         );
  INV_X1 U4897 ( .A(n3965), .ZN(n3966) );
  OR2_X1 U4898 ( .A1(n3969), .A2(n3449), .ZN(n4265) );
  AND2_X4 U4899 ( .A1(n4092), .A2(n3159), .ZN(n4438) );
  OAI22_X1 U4900 ( .A1(n3971), .A2(n5690), .B1(n3964), .B2(n3983), .ZN(n3972)
         );
  INV_X1 U4901 ( .A(n3972), .ZN(n3973) );
  NAND4_X1 U4902 ( .A1(n4265), .A2(n6226), .A3(n3970), .A4(n3973), .ZN(n3974)
         );
  NAND2_X1 U4903 ( .A1(n3175), .A2(n4092), .ZN(n3981) );
  INV_X1 U4904 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U4905 ( .A1(n4057), .A2(n5392), .ZN(n3979) );
  NAND2_X1 U4906 ( .A1(n4438), .A2(n5392), .ZN(n3977) );
  NAND2_X1 U4907 ( .A1(n4869), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3976) );
  NAND3_X1 U4908 ( .A1(n3977), .A2(n3975), .A3(n3976), .ZN(n3978) );
  NAND2_X1 U4909 ( .A1(n3979), .A2(n3978), .ZN(n5322) );
  INV_X1 U4910 ( .A(n4057), .ZN(n4050) );
  MUX2_X1 U4911 ( .A(n4050), .B(n4869), .S(EBX_REG_3__SCAN_IN), .Z(n3980) );
  NAND2_X1 U4912 ( .A1(n3980), .A2(n2975), .ZN(n4335) );
  NAND2_X2 U4913 ( .A1(n4785), .A2(n4438), .ZN(n4061) );
  MUX2_X1 U4914 ( .A(n4061), .B(n3975), .S(EBX_REG_1__SCAN_IN), .Z(n3986) );
  NAND2_X1 U4915 ( .A1(n2957), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3984)
         );
  AND2_X1 U4916 ( .A1(n4027), .A2(n3984), .ZN(n3985) );
  NAND2_X1 U4917 ( .A1(n3975), .A2(EBX_REG_0__SCAN_IN), .ZN(n3988) );
  INV_X1 U4918 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U4919 ( .A1(n4869), .A2(n4512), .ZN(n3987) );
  NAND2_X1 U4920 ( .A1(n3988), .A2(n3987), .ZN(n4207) );
  XNOR2_X1 U4921 ( .A(n3989), .B(n4207), .ZN(n4221) );
  MUX2_X1 U4922 ( .A(n4061), .B(n3975), .S(EBX_REG_2__SCAN_IN), .Z(n3992) );
  NAND3_X1 U4923 ( .A1(n3983), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n4869), 
        .ZN(n3990) );
  AND2_X1 U4924 ( .A1(n4027), .A2(n3990), .ZN(n3991) );
  NAND2_X1 U4925 ( .A1(n3992), .A2(n3991), .ZN(n4247) );
  NAND2_X1 U4926 ( .A1(n3975), .A2(n5620), .ZN(n3994) );
  INV_X1 U4927 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U4928 ( .A1(n4438), .A2(n5360), .ZN(n3993) );
  NAND3_X1 U4929 ( .A1(n3994), .A2(n4869), .A3(n3993), .ZN(n3995) );
  OAI21_X1 U4930 ( .B1(n4061), .B2(EBX_REG_4__SCAN_IN), .A(n3995), .ZN(n4319)
         );
  NAND2_X1 U4931 ( .A1(n4334), .A2(n4319), .ZN(n4320) );
  MUX2_X1 U4932 ( .A(n4057), .B(n4785), .S(EBX_REG_5__SCAN_IN), .Z(n3997) );
  NOR2_X1 U4933 ( .A1(n4206), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3996)
         );
  NOR2_X1 U4934 ( .A1(n3997), .A2(n3996), .ZN(n4363) );
  MUX2_X1 U4935 ( .A(n4061), .B(n3975), .S(EBX_REG_6__SCAN_IN), .Z(n3999) );
  NAND2_X1 U4936 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n3983), .ZN(n3998)
         );
  NOR2_X2 U4937 ( .A1(n4376), .A2(n4375), .ZN(n4457) );
  MUX2_X1 U4938 ( .A(n4057), .B(n4785), .S(EBX_REG_7__SCAN_IN), .Z(n4001) );
  NOR2_X1 U4939 ( .A1(n4206), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4000)
         );
  NOR2_X1 U4940 ( .A1(n4001), .A2(n4000), .ZN(n4456) );
  MUX2_X1 U4941 ( .A(n4061), .B(n3975), .S(EBX_REG_8__SCAN_IN), .Z(n4004) );
  NAND2_X1 U4942 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n3983), .ZN(n4002)
         );
  AND2_X1 U4943 ( .A1(n4027), .A2(n4002), .ZN(n4003) );
  NAND2_X1 U4944 ( .A1(n4004), .A2(n4003), .ZN(n4454) );
  INV_X1 U4945 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U4946 ( .A1(n4057), .A2(n5397), .ZN(n4008) );
  NAND2_X1 U4947 ( .A1(n4438), .A2(n5397), .ZN(n4006) );
  NAND2_X1 U4948 ( .A1(n4869), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4005)
         );
  NAND3_X1 U4949 ( .A1(n4006), .A2(n3975), .A3(n4005), .ZN(n4007) );
  MUX2_X1 U4950 ( .A(n4061), .B(n3975), .S(EBX_REG_10__SCAN_IN), .Z(n4010) );
  NAND2_X1 U4951 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n3983), .ZN(n4009) );
  NAND2_X1 U4952 ( .A1(n3975), .A2(n4011), .ZN(n4013) );
  INV_X1 U4953 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U4954 ( .A1(n4438), .A2(n6413), .ZN(n4012) );
  NAND3_X1 U4955 ( .A1(n4013), .A2(n4869), .A3(n4012), .ZN(n4014) );
  OAI21_X1 U4956 ( .B1(n4061), .B2(EBX_REG_12__SCAN_IN), .A(n4014), .ZN(n4536)
         );
  INV_X1 U4957 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U4958 ( .A1(n4057), .A2(n5390), .ZN(n4017) );
  NAND2_X1 U4959 ( .A1(n4869), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4015) );
  OAI211_X1 U4960 ( .C1(n3983), .C2(EBX_REG_13__SCAN_IN), .A(n3975), .B(n4015), 
        .ZN(n4016) );
  NAND2_X1 U4961 ( .A1(n4017), .A2(n4016), .ZN(n5256) );
  MUX2_X1 U4962 ( .A(n4061), .B(n3975), .S(EBX_REG_14__SCAN_IN), .Z(n4020) );
  NAND2_X1 U4963 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n3983), .ZN(n4018) );
  AND2_X1 U4964 ( .A1(n4027), .A2(n4018), .ZN(n4019) );
  NAND2_X1 U4965 ( .A1(n4020), .A2(n4019), .ZN(n4579) );
  INV_X1 U4966 ( .A(EBX_REG_15__SCAN_IN), .ZN(n4610) );
  NAND2_X1 U4967 ( .A1(n4057), .A2(n4610), .ZN(n4023) );
  NAND2_X1 U4968 ( .A1(n4869), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4021) );
  OAI211_X1 U4969 ( .C1(n3983), .C2(EBX_REG_15__SCAN_IN), .A(n3975), .B(n4021), 
        .ZN(n4022) );
  MUX2_X1 U4970 ( .A(n4050), .B(n4869), .S(EBX_REG_17__SCAN_IN), .Z(n4024) );
  OAI21_X1 U4971 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n4206), .A(n4024), 
        .ZN(n4025) );
  INV_X1 U4972 ( .A(n4025), .ZN(n4797) );
  MUX2_X1 U4973 ( .A(n4061), .B(n3975), .S(EBX_REG_16__SCAN_IN), .Z(n4029) );
  NAND2_X1 U4974 ( .A1(n3983), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4026) );
  AND2_X1 U4975 ( .A1(n4027), .A2(n4026), .ZN(n4028) );
  NAND2_X1 U4976 ( .A1(n4029), .A2(n4028), .ZN(n4809) );
  NAND2_X1 U4977 ( .A1(n4797), .A2(n4809), .ZN(n4030) );
  INV_X1 U4978 ( .A(n4061), .ZN(n4065) );
  INV_X1 U4979 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U4980 ( .A1(n4065), .A2(n4875), .ZN(n4034) );
  INV_X1 U4981 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U4982 ( .A1(n3975), .A2(n6476), .ZN(n4032) );
  NAND2_X1 U4983 ( .A1(n4438), .A2(n4875), .ZN(n4031) );
  NAND3_X1 U4984 ( .A1(n4032), .A2(n4869), .A3(n4031), .ZN(n4033) );
  NAND2_X1 U4985 ( .A1(n4034), .A2(n4033), .ZN(n4788) );
  NAND2_X1 U4986 ( .A1(n4784), .A2(n4788), .ZN(n4868) );
  OR2_X1 U4987 ( .A1(n4206), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4035)
         );
  INV_X1 U4988 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4886) );
  NAND2_X1 U4989 ( .A1(n4438), .A2(n4886), .ZN(n4786) );
  NAND2_X1 U4990 ( .A1(n4035), .A2(n4786), .ZN(n4870) );
  AND2_X1 U4991 ( .A1(n4870), .A2(n4869), .ZN(n4038) );
  INV_X1 U4992 ( .A(n4206), .ZN(n4078) );
  NOR2_X1 U4993 ( .A1(n3983), .A2(EBX_REG_20__SCAN_IN), .ZN(n4036) );
  AOI21_X1 U4994 ( .B1(n4078), .B2(n5086), .A(n4036), .ZN(n4871) );
  INV_X1 U4995 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4873) );
  OAI22_X1 U4996 ( .A1(n4871), .A2(n4870), .B1(n4869), .B2(n4873), .ZN(n4037)
         );
  NAND2_X1 U4997 ( .A1(n4869), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4039) );
  OAI211_X1 U4998 ( .C1(n3983), .C2(EBX_REG_21__SCAN_IN), .A(n3975), .B(n4039), 
        .ZN(n4040) );
  OAI21_X1 U4999 ( .B1(n4050), .B2(EBX_REG_21__SCAN_IN), .A(n4040), .ZN(n5068)
         );
  INV_X1 U5000 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U5001 ( .A1(n4057), .A2(n5149), .ZN(n4043) );
  NAND2_X1 U5002 ( .A1(n4869), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4041) );
  OAI211_X1 U5003 ( .C1(n3983), .C2(EBX_REG_23__SCAN_IN), .A(n3975), .B(n4041), 
        .ZN(n4042) );
  AND2_X1 U5004 ( .A1(n4043), .A2(n4042), .ZN(n4855) );
  INV_X1 U5005 ( .A(EBX_REG_22__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5006 ( .A1(n4065), .A2(n4863), .ZN(n4048) );
  INV_X1 U5007 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4044) );
  NAND2_X1 U5008 ( .A1(n3975), .A2(n4044), .ZN(n4046) );
  NAND2_X1 U5009 ( .A1(n4438), .A2(n4863), .ZN(n4045) );
  NAND3_X1 U5010 ( .A1(n4046), .A2(n4869), .A3(n4045), .ZN(n4047) );
  NAND2_X1 U5011 ( .A1(n4048), .A2(n4047), .ZN(n4862) );
  AND2_X1 U5012 ( .A1(n4855), .A2(n4862), .ZN(n4049) );
  MUX2_X1 U5013 ( .A(n4050), .B(n4869), .S(EBX_REG_25__SCAN_IN), .Z(n4051) );
  OAI21_X1 U5014 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4206), .A(n4051), 
        .ZN(n4840) );
  INV_X1 U5015 ( .A(n4840), .ZN(n4054) );
  MUX2_X1 U5016 ( .A(n4061), .B(n3975), .S(EBX_REG_24__SCAN_IN), .Z(n4053) );
  NAND2_X1 U5017 ( .A1(n3983), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4052) );
  NAND2_X1 U5018 ( .A1(n4053), .A2(n4052), .ZN(n4849) );
  MUX2_X1 U5019 ( .A(n4061), .B(n3975), .S(EBX_REG_26__SCAN_IN), .Z(n4056) );
  NAND2_X1 U5020 ( .A1(n3983), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4055) );
  AND2_X1 U5021 ( .A1(n4056), .A2(n4055), .ZN(n4832) );
  NOR2_X2 U5022 ( .A1(n4842), .A2(n4832), .ZN(n4833) );
  INV_X1 U5023 ( .A(EBX_REG_27__SCAN_IN), .ZN(n4771) );
  NAND2_X1 U5024 ( .A1(n4057), .A2(n4771), .ZN(n4060) );
  NAND2_X1 U5025 ( .A1(n4869), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4058) );
  OAI211_X1 U5026 ( .C1(n3983), .C2(EBX_REG_27__SCAN_IN), .A(n3975), .B(n4058), 
        .ZN(n4059) );
  AND2_X1 U5027 ( .A1(n4060), .A2(n4059), .ZN(n4766) );
  MUX2_X1 U5028 ( .A(n4061), .B(n3975), .S(EBX_REG_28__SCAN_IN), .Z(n4063) );
  NAND2_X1 U5029 ( .A1(n3983), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U5030 ( .A1(n4063), .A2(n4062), .ZN(n4756) );
  NOR2_X1 U5031 ( .A1(n3983), .A2(EBX_REG_29__SCAN_IN), .ZN(n4064) );
  AOI21_X1 U5032 ( .B1(n4078), .B2(n5002), .A(n4064), .ZN(n4740) );
  INV_X1 U5033 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4825) );
  NAND2_X1 U5034 ( .A1(n4065), .A2(n4825), .ZN(n4741) );
  AOI21_X1 U5035 ( .B1(n4685), .B2(n4869), .A(n4066), .ZN(n4745) );
  NAND2_X1 U5036 ( .A1(n4206), .A2(EBX_REG_30__SCAN_IN), .ZN(n4068) );
  NAND2_X1 U5037 ( .A1(n3983), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4067) );
  NAND2_X1 U5038 ( .A1(n4068), .A2(n4067), .ZN(n4682) );
  INV_X1 U5039 ( .A(n4685), .ZN(n4069) );
  NAND2_X1 U5040 ( .A1(n4069), .A2(n4869), .ZN(n4679) );
  OAI22_X1 U5041 ( .A1(n4206), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3983), .ZN(n4070) );
  INV_X1 U5042 ( .A(n4070), .ZN(n4071) );
  OR2_X1 U5043 ( .A1(n3964), .A2(n4434), .ZN(n6239) );
  OAI21_X1 U5044 ( .B1(n3971), .B2(n4072), .A(n6239), .ZN(n4073) );
  INV_X1 U5045 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6322) );
  NOR2_X1 U5046 ( .A1(n5612), .A2(n6322), .ZN(n4702) );
  NAND2_X1 U5047 ( .A1(n5662), .A2(n4092), .ZN(n4495) );
  OR2_X1 U5048 ( .A1(n4495), .A2(n3142), .ZN(n4196) );
  OAI211_X1 U5049 ( .C1(n3150), .C2(n3125), .A(n4074), .B(n4196), .ZN(n4075)
         );
  INV_X1 U5050 ( .A(n4075), .ZN(n4077) );
  OAI211_X1 U5051 ( .C1(n4079), .C2(n4078), .A(n4077), .B(n4076), .ZN(n4080)
         );
  OR2_X1 U5052 ( .A1(n4081), .A2(n4080), .ZN(n4182) );
  NOR2_X1 U5053 ( .A1(n3178), .A2(n4082), .ZN(n4083) );
  NAND2_X1 U5054 ( .A1(n4093), .A2(n4267), .ZN(n5077) );
  AOI21_X1 U5055 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n5634) );
  NOR2_X1 U5056 ( .A1(n5628), .A2(n5620), .ZN(n5610) );
  NAND3_X1 U5057 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n5610), .ZN(n4090) );
  NOR2_X1 U5058 ( .A1(n5634), .A2(n4090), .ZN(n5562) );
  NAND2_X1 U5059 ( .A1(n5632), .A2(n5562), .ZN(n5570) );
  NOR2_X1 U5060 ( .A1(n6482), .A2(n5592), .ZN(n5588) );
  NAND3_X1 U5061 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5588), .ZN(n4091) );
  NAND2_X1 U5062 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5254) );
  NOR2_X1 U5063 ( .A1(n3427), .A2(n5254), .ZN(n5247) );
  NAND2_X1 U5064 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5247), .ZN(n5104) );
  NAND2_X1 U5065 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5105) );
  NOR2_X1 U5066 ( .A1(n5104), .A2(n5105), .ZN(n4089) );
  NAND2_X1 U5067 ( .A1(n4593), .A2(n4089), .ZN(n5082) );
  INV_X1 U5068 ( .A(n5091), .ZN(n4085) );
  AND2_X1 U5069 ( .A1(n4085), .A2(n5078), .ZN(n4095) );
  INV_X1 U5070 ( .A(n4095), .ZN(n4088) );
  INV_X2 U5071 ( .A(n5612), .ZN(n5630) );
  NOR2_X1 U5072 ( .A1(n4093), .A2(n5630), .ZN(n5650) );
  NAND2_X1 U5073 ( .A1(n4093), .A2(n4086), .ZN(n5242) );
  NAND2_X1 U5074 ( .A1(n5077), .A2(n5242), .ZN(n5244) );
  INV_X1 U5075 ( .A(n5244), .ZN(n4087) );
  NOR2_X1 U5076 ( .A1(n4087), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5645)
         );
  NOR2_X1 U5077 ( .A1(n5650), .A2(n5645), .ZN(n4381) );
  NAND2_X1 U5078 ( .A1(n5077), .A2(n4381), .ZN(n5571) );
  OAI21_X1 U5079 ( .B1(n5082), .B2(n4088), .A(n5571), .ZN(n4098) );
  INV_X1 U5080 ( .A(n4089), .ZN(n4107) );
  NAND2_X1 U5081 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4378) );
  OR2_X1 U5082 ( .A1(n4090), .A2(n4378), .ZN(n5568) );
  OR2_X1 U5083 ( .A1(n4091), .A2(n5568), .ZN(n4594) );
  NOR2_X1 U5084 ( .A1(n4107), .A2(n4594), .ZN(n5080) );
  AND2_X1 U5085 ( .A1(n4092), .A2(n3948), .ZN(n6216) );
  INV_X1 U5086 ( .A(n5242), .ZN(n4094) );
  INV_X1 U5087 ( .A(n5569), .ZN(n5079) );
  AOI21_X1 U5088 ( .B1(n4095), .B2(n5080), .A(n5079), .ZN(n4096) );
  INV_X1 U5089 ( .A(n4096), .ZN(n4097) );
  AND2_X1 U5090 ( .A1(n4098), .A2(n4097), .ZN(n5057) );
  NAND2_X1 U5091 ( .A1(n5103), .A2(n5042), .ZN(n4099) );
  AND2_X1 U5092 ( .A1(n5057), .A2(n4099), .ZN(n5050) );
  NOR2_X1 U5093 ( .A1(n5651), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4256)
         );
  INV_X1 U5094 ( .A(n4256), .ZN(n4100) );
  INV_X1 U5095 ( .A(n4101), .ZN(n4102) );
  OAI21_X1 U5096 ( .B1(n5639), .B2(n5632), .A(n4102), .ZN(n4103) );
  NAND2_X1 U5097 ( .A1(n5050), .A2(n4103), .ZN(n5037) );
  AND2_X1 U5098 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5007) );
  AOI21_X1 U5099 ( .B1(n5007), .B2(n5003), .A(n5572), .ZN(n4104) );
  NOR2_X1 U5100 ( .A1(n5037), .A2(n4104), .ZN(n4997) );
  INV_X1 U5101 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4691) );
  OAI21_X1 U5102 ( .B1(n4691), .B2(n5002), .A(n5103), .ZN(n4105) );
  AOI21_X1 U5103 ( .B1(n4997), .B2(n4105), .A(n3945), .ZN(n4106) );
  NAND2_X1 U5104 ( .A1(n5229), .A2(n5078), .ZN(n5090) );
  NOR2_X1 U5105 ( .A1(n5090), .A2(n5027), .ZN(n5025) );
  NAND2_X1 U5106 ( .A1(n5025), .A2(n5007), .ZN(n5024) );
  INV_X1 U5107 ( .A(n5003), .ZN(n5011) );
  NOR3_X1 U5108 ( .A1(n5024), .A2(n5011), .A3(n5002), .ZN(n4692) );
  NAND3_X1 U5109 ( .A1(n4692), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n3945), .ZN(n4108) );
  OAI21_X1 U5110 ( .B1(n4707), .B2(n5654), .A(n4109), .ZN(U2987) );
  INV_X1 U5111 ( .A(n4676), .ZN(n4922) );
  NAND2_X1 U5112 ( .A1(n4996), .A2(n5541), .ZN(n4163) );
  INV_X1 U5113 ( .A(n4112), .ZN(n4113) );
  XNOR2_X1 U5114 ( .A(n4423), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4746)
         );
  INV_X1 U5115 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6421) );
  NOR2_X1 U5116 ( .A1(n5612), .A2(n6421), .ZN(n5000) );
  INV_X1 U5117 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4748) );
  NOR2_X1 U5118 ( .A1(n5550), .A2(n4748), .ZN(n4114) );
  AOI211_X1 U5119 ( .C1(n5517), .C2(n4746), .A(n5000), .B(n4114), .ZN(n4162)
         );
  INV_X1 U5120 ( .A(n4115), .ZN(n4116) );
  INV_X1 U5121 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U5122 ( .A1(n4116), .A2(n4759), .ZN(n4117) );
  NAND2_X1 U5123 ( .A1(n4423), .A2(n4117), .ZN(n4915) );
  NOR2_X1 U5124 ( .A1(n4119), .A2(n4118), .ZN(n4138) );
  AOI22_X1 U5125 ( .A1(n3079), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5126 ( .A1(n3077), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5127 ( .A1(n4120), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5128 ( .A1(n3672), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4121) );
  NAND4_X1 U5129 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), .ZN(n4131)
         );
  AOI22_X1 U5130 ( .A1(n4147), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5131 ( .A1(n3281), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5132 ( .A1(n3912), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3230), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5133 ( .A1(n4125), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4126) );
  NAND4_X1 U5134 ( .A1(n4129), .A2(n4128), .A3(n4127), .A4(n4126), .ZN(n4130)
         );
  OR2_X1 U5135 ( .A1(n4131), .A2(n4130), .ZN(n4137) );
  XNOR2_X1 U5136 ( .A(n4138), .B(n4137), .ZN(n4134) );
  AOI21_X1 U5137 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n3558), .A(n4419), 
        .ZN(n4133) );
  NAND2_X1 U5138 ( .A1(n4659), .A2(EAX_REG_28__SCAN_IN), .ZN(n4132) );
  OAI211_X1 U5139 ( .C1(n4134), .C2(n4652), .A(n4133), .B(n4132), .ZN(n4135)
         );
  OAI21_X1 U5140 ( .B1(n4649), .B2(n4915), .A(n4135), .ZN(n4755) );
  NAND2_X1 U5141 ( .A1(n4138), .A2(n4137), .ZN(n4644) );
  AOI22_X1 U5142 ( .A1(n3079), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5143 ( .A1(n4272), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4635), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5144 ( .A1(n4140), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5145 ( .A1(n4637), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4141) );
  NAND4_X1 U5146 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4141), .ZN(n4153)
         );
  AOI22_X1 U5147 ( .A1(n4146), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5148 ( .A1(n3281), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4147), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5149 ( .A1(n3672), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5150 ( .A1(n3912), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4148) );
  NAND4_X1 U5151 ( .A1(n4151), .A2(n4150), .A3(n4149), .A4(n4148), .ZN(n4152)
         );
  NOR2_X1 U5152 ( .A1(n4153), .A2(n4152), .ZN(n4645) );
  XOR2_X1 U5153 ( .A(n4644), .B(n4645), .Z(n4155) );
  NAND2_X1 U5154 ( .A1(n4155), .A2(n4154), .ZN(n4158) );
  AOI21_X1 U5155 ( .B1(n4748), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4156) );
  AOI21_X1 U5156 ( .B1(n3506), .B2(EAX_REG_29__SCAN_IN), .A(n4156), .ZN(n4157)
         );
  NAND3_X1 U5157 ( .A1(n4163), .A2(n4162), .A3(n4161), .ZN(U2957) );
  INV_X1 U5158 ( .A(n4168), .ZN(n4173) );
  NAND2_X1 U5159 ( .A1(n3948), .A2(n4173), .ZN(n4165) );
  AOI22_X1 U5160 ( .A1(n4199), .A2(n3449), .B1(n4164), .B2(n4165), .ZN(n5271)
         );
  NAND2_X1 U5161 ( .A1(n6364), .A2(n6266), .ZN(n4166) );
  OAI211_X1 U5162 ( .C1(n3178), .C2(n4167), .A(n4166), .B(n6271), .ZN(n6362)
         );
  NAND2_X1 U5163 ( .A1(n5271), .A2(n6362), .ZN(n6227) );
  AND2_X1 U5164 ( .A1(n6227), .A2(n6251), .ZN(n5278) );
  INV_X1 U5165 ( .A(MORE_REG_SCAN_IN), .ZN(n6228) );
  NAND3_X1 U5166 ( .A1(n4265), .A2(n6226), .A3(n4164), .ZN(n4169) );
  AOI22_X1 U5167 ( .A1(n4199), .A2(n4169), .B1(n3948), .B2(n4168), .ZN(n4171)
         );
  NAND2_X1 U5168 ( .A1(n4177), .A2(n4267), .ZN(n4170) );
  NAND2_X1 U5169 ( .A1(n4171), .A2(n4170), .ZN(n6230) );
  NAND2_X1 U5170 ( .A1(n5278), .A2(n6230), .ZN(n4172) );
  OAI21_X1 U5171 ( .B1(n5278), .B2(n6228), .A(n4172), .ZN(U3471) );
  NAND3_X1 U5172 ( .A1(n3948), .A2(n6251), .A3(n4173), .ZN(n5114) );
  NAND2_X1 U5173 ( .A1(n4434), .A2(n4495), .ZN(n4176) );
  INV_X1 U5174 ( .A(n5115), .ZN(n4174) );
  OAI21_X1 U5175 ( .B1(n4174), .B2(READREQUEST_REG_SCAN_IN), .A(n6368), .ZN(
        n4175) );
  OAI21_X1 U5176 ( .B1(n6368), .B2(n4176), .A(n4175), .ZN(U3474) );
  INV_X1 U5177 ( .A(n4178), .ZN(n4189) );
  AOI22_X1 U5178 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n3945), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4179), .ZN(n4664) );
  INV_X1 U5179 ( .A(n4664), .ZN(n4188) );
  NAND2_X1 U5180 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4665) );
  INV_X1 U5181 ( .A(n6252), .ZN(n6342) );
  INV_X1 U5182 ( .A(n5855), .ZN(n5797) );
  NAND3_X1 U5183 ( .A1(n3970), .A2(n4180), .A3(n3964), .ZN(n4181) );
  OR2_X1 U5184 ( .A1(n4182), .A2(n4181), .ZN(n6215) );
  INV_X1 U5185 ( .A(n6216), .ZN(n4223) );
  NOR2_X1 U5186 ( .A1(n4223), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4187)
         );
  NOR3_X1 U5187 ( .A1(n4185), .A2(n4183), .A3(n4184), .ZN(n4186) );
  AOI211_X1 U5188 ( .C1(n5797), .C2(n6215), .A(n4187), .B(n4186), .ZN(n6212)
         );
  OAI222_X1 U5189 ( .A1(n6333), .A2(n4189), .B1(n4188), .B2(n4665), .C1(n6342), 
        .C2(n6212), .ZN(n4204) );
  INV_X1 U5190 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6331) );
  OR2_X1 U5191 ( .A1(n4199), .A2(n4265), .ZN(n4193) );
  INV_X1 U5192 ( .A(n4190), .ZN(n4191) );
  OR2_X1 U5193 ( .A1(n3970), .A2(n4191), .ZN(n4192) );
  NAND2_X1 U5194 ( .A1(n4193), .A2(n4192), .ZN(n4238) );
  INV_X1 U5195 ( .A(n4238), .ZN(n4201) );
  AOI21_X1 U5196 ( .B1(n3983), .B2(n6266), .A(READY_N), .ZN(n4194) );
  OAI21_X1 U5197 ( .B1(n6216), .B2(n3112), .A(n4194), .ZN(n4197) );
  OAI211_X1 U5198 ( .C1(n4199), .C2(n4197), .A(n4196), .B(n4195), .ZN(n4198)
         );
  INV_X1 U5199 ( .A(n4198), .ZN(n4200) );
  NAND2_X1 U5200 ( .A1(n4267), .A2(n4199), .ZN(n4212) );
  OR2_X1 U5201 ( .A1(n6211), .A2(n6236), .ZN(n4203) );
  INV_X1 U5202 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6229) );
  NOR2_X1 U5203 ( .A1(n6425), .A2(n3558), .ZN(n6243) );
  NAND2_X1 U5204 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6243), .ZN(n6329) );
  OR2_X1 U5205 ( .A1(n6229), .A2(n6329), .ZN(n4202) );
  AND2_X1 U5206 ( .A1(n4203), .A2(n4202), .ZN(n5265) );
  OAI21_X1 U5207 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6331), .A(n5265), .ZN(
        n6340) );
  OAI21_X1 U5208 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6333), .A(n6340), 
        .ZN(n6338) );
  AOI22_X1 U5209 ( .A1(n4204), .A2(n6340), .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n6338), .ZN(n4205) );
  INV_X1 U5210 ( .A(n4205), .ZN(U3460) );
  OR2_X1 U5211 ( .A1(n4206), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4208)
         );
  NAND2_X1 U5212 ( .A1(n4208), .A2(n4207), .ZN(n5644) );
  AND3_X1 U5213 ( .A1(n5690), .A2(n3132), .A3(n3505), .ZN(n4209) );
  NAND2_X1 U5214 ( .A1(n4210), .A2(n4209), .ZN(n4236) );
  OR2_X1 U5215 ( .A1(n4236), .A2(n3983), .ZN(n4211) );
  NAND2_X1 U5216 ( .A1(n4212), .A2(n4211), .ZN(n4213) );
  INV_X2 U5217 ( .A(n5394), .ZN(n4891) );
  XOR2_X1 U5218 ( .A(n4215), .B(n4214), .Z(n5553) );
  INV_X1 U5219 ( .A(n5553), .ZN(n4245) );
  OAI222_X1 U5220 ( .A1(n5644), .A2(n5178), .B1(n5398), .B2(n4512), .C1(n4891), 
        .C2(n4245), .ZN(U2859) );
  OR2_X1 U5221 ( .A1(n4217), .A2(n4216), .ZN(n4218) );
  NAND2_X1 U5222 ( .A1(n4219), .A2(n4218), .ZN(n5381) );
  OAI21_X1 U5223 ( .B1(n4221), .B2(n4438), .A(n4220), .ZN(n5376) );
  INV_X1 U5224 ( .A(n5398), .ZN(n4889) );
  AOI22_X1 U5225 ( .A1(n5393), .A2(n5376), .B1(EBX_REG_1__SCAN_IN), .B2(n4889), 
        .ZN(n4222) );
  OAI21_X1 U5226 ( .B1(n5381), .B2(n4891), .A(n4222), .ZN(U2858) );
  INV_X1 U5227 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U5228 ( .A1(n5511), .A2(n4224), .ZN(n4225) );
  NAND2_X1 U5229 ( .A1(n5412), .A2(n3178), .ZN(n4359) );
  AND2_X2 U5230 ( .A1(n6243), .A2(n6366), .ZN(n6237) );
  INV_X1 U5231 ( .A(n6237), .ZN(n6371) );
  NOR2_X4 U5232 ( .A1(n6237), .A2(n5412), .ZN(n5423) );
  AOI22_X1 U5233 ( .A1(n6237), .A2(UWORD_REG_10__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4226) );
  OAI21_X1 U5234 ( .B1(n5453), .B2(n4359), .A(n4226), .ZN(U2897) );
  INV_X1 U5235 ( .A(EAX_REG_29__SCAN_IN), .ZN(n5461) );
  AOI22_X1 U5236 ( .A1(n6237), .A2(UWORD_REG_13__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4227) );
  OAI21_X1 U5237 ( .B1(n5461), .B2(n4359), .A(n4227), .ZN(U2894) );
  INV_X1 U5238 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6526) );
  AOI22_X1 U5239 ( .A1(n6237), .A2(UWORD_REG_12__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4228) );
  OAI21_X1 U5240 ( .B1(n6526), .B2(n4359), .A(n4228), .ZN(U2895) );
  AOI22_X1 U5241 ( .A1(n6237), .A2(UWORD_REG_8__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4229) );
  OAI21_X1 U5242 ( .B1(n6453), .B2(n4359), .A(n4229), .ZN(U2899) );
  XNOR2_X1 U5243 ( .A(n4231), .B(n4230), .ZN(n4262) );
  INV_X1 U5244 ( .A(n5381), .ZN(n4234) );
  AOI22_X1 U5245 ( .A1(n5536), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5630), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4232) );
  OAI21_X1 U5246 ( .B1(n5546), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4232), 
        .ZN(n4233) );
  AOI21_X1 U5247 ( .B1(n4234), .B2(n5702), .A(n4233), .ZN(n4235) );
  OAI21_X1 U5248 ( .B1(n4262), .B2(n5555), .A(n4235), .ZN(U2985) );
  NOR2_X1 U5249 ( .A1(n4236), .A2(n3449), .ZN(n4237) );
  NAND2_X1 U5250 ( .A1(n4438), .A2(n6271), .ZN(n4239) );
  INV_X1 U5251 ( .A(n4893), .ZN(n4242) );
  AND2_X1 U5252 ( .A1(n4242), .A2(n4661), .ZN(n4243) );
  INV_X1 U5253 ( .A(n4243), .ZN(n4244) );
  INV_X1 U5254 ( .A(DATAI_0_), .ZN(n5659) );
  INV_X1 U5255 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5468) );
  OAI222_X1 U5256 ( .A1(n5182), .A2(n4245), .B1(n4402), .B2(n5659), .C1(n4894), 
        .C2(n5468), .ZN(U2891) );
  INV_X1 U5257 ( .A(n4246), .ZN(n4249) );
  INV_X1 U5258 ( .A(n4247), .ZN(n4248) );
  NAND2_X1 U5259 ( .A1(n4249), .A2(n4248), .ZN(n4250) );
  AND2_X1 U5260 ( .A1(n4250), .A2(n4336), .ZN(n5631) );
  INV_X1 U5261 ( .A(n5631), .ZN(n4255) );
  INV_X1 U5262 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4254) );
  OAI21_X1 U5263 ( .B1(n4253), .B2(n4252), .A(n4251), .ZN(n5537) );
  OAI222_X1 U5264 ( .A1(n4255), .A2(n5178), .B1(n5398), .B2(n4254), .C1(n5537), 
        .C2(n4891), .ZN(U2857) );
  INV_X1 U5265 ( .A(DATAI_1_), .ZN(n6474) );
  INV_X1 U5266 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5471) );
  OAI222_X1 U5267 ( .A1(n5381), .A2(n5182), .B1(n4402), .B2(n6474), .C1(n4894), 
        .C2(n5471), .ZN(U2890) );
  NOR2_X1 U5268 ( .A1(n5572), .A2(n4256), .ZN(n4258) );
  INV_X1 U5269 ( .A(n4381), .ZN(n4257) );
  MUX2_X1 U5270 ( .A(n4258), .B(n4257), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4260) );
  INV_X1 U5271 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6353) );
  NOR2_X1 U5272 ( .A1(n5612), .A2(n6353), .ZN(n4259) );
  AOI211_X1 U5273 ( .C1(n5649), .C2(n5376), .A(n4260), .B(n4259), .ZN(n4261)
         );
  OAI21_X1 U5274 ( .B1(n4262), .B2(n5654), .A(n4261), .ZN(U3017) );
  NAND2_X1 U5275 ( .A1(n6425), .A2(n3558), .ZN(n6365) );
  INV_X1 U5276 ( .A(n6365), .ZN(n5270) );
  NAND2_X1 U5277 ( .A1(n4264), .A2(n6215), .ZN(n4279) );
  INV_X1 U5278 ( .A(n4265), .ZN(n4266) );
  OR2_X1 U5279 ( .A1(n4267), .A2(n4266), .ZN(n4289) );
  MUX2_X1 U5280 ( .A(n4268), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4184), 
        .Z(n4270) );
  NOR2_X1 U5281 ( .A1(n4270), .A2(n4269), .ZN(n4277) );
  AOI21_X1 U5282 ( .B1(n4184), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3023), 
        .ZN(n4271) );
  NOR2_X1 U5283 ( .A1(n4272), .A2(n4271), .ZN(n6334) );
  XNOR2_X1 U5284 ( .A(n4273), .B(n3023), .ZN(n4274) );
  NAND2_X1 U5285 ( .A1(n6216), .A2(n4274), .ZN(n4275) );
  OAI21_X1 U5286 ( .B1(n6334), .B2(n4286), .A(n4275), .ZN(n4276) );
  AOI21_X1 U5287 ( .B1(n4289), .B2(n4277), .A(n4276), .ZN(n4278) );
  NAND2_X1 U5288 ( .A1(n4279), .A2(n4278), .ZN(n6332) );
  INV_X1 U5289 ( .A(n6211), .ZN(n4292) );
  NAND2_X1 U5290 ( .A1(n6332), .A2(n4292), .ZN(n4281) );
  NAND2_X1 U5291 ( .A1(n6211), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4280) );
  NAND2_X1 U5292 ( .A1(n4281), .A2(n4280), .ZN(n6225) );
  INV_X1 U5293 ( .A(n6215), .ZN(n4283) );
  OR2_X1 U5294 ( .A1(n2965), .A2(n4283), .ZN(n4291) );
  XNOR2_X1 U5295 ( .A(n4184), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4288)
         );
  XNOR2_X1 U5296 ( .A(n3164), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4284)
         );
  NAND2_X1 U5297 ( .A1(n6216), .A2(n4284), .ZN(n4285) );
  OAI21_X1 U5298 ( .B1(n4288), .B2(n4286), .A(n4285), .ZN(n4287) );
  AOI21_X1 U5299 ( .B1(n4289), .B2(n4288), .A(n4287), .ZN(n4290) );
  NAND2_X1 U5300 ( .A1(n4291), .A2(n4290), .ZN(n4668) );
  NAND2_X1 U5301 ( .A1(n4292), .A2(n4668), .ZN(n4294) );
  NAND2_X1 U5302 ( .A1(n6211), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4293) );
  NAND2_X1 U5303 ( .A1(n4294), .A2(n4293), .ZN(n6220) );
  NAND3_X1 U5304 ( .A1(n6225), .A2(n6425), .A3(n6220), .ZN(n4297) );
  NAND2_X1 U5305 ( .A1(n6229), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4303) );
  INV_X1 U5306 ( .A(n4303), .ZN(n4295) );
  NAND2_X1 U5307 ( .A1(n4269), .A2(n4295), .ZN(n4296) );
  NAND2_X1 U5308 ( .A1(n4297), .A2(n4296), .ZN(n6233) );
  INV_X1 U5309 ( .A(n4183), .ZN(n4298) );
  NAND2_X1 U5310 ( .A1(n6233), .A2(n4298), .ZN(n6245) );
  INV_X1 U5311 ( .A(n5826), .ZN(n5801) );
  NOR2_X1 U5312 ( .A1(n2958), .A2(n5801), .ZN(n4300) );
  XNOR2_X1 U5313 ( .A(n4300), .B(n4299), .ZN(n5354) );
  INV_X1 U5314 ( .A(n3970), .ZN(n5266) );
  NAND2_X1 U5315 ( .A1(n5354), .A2(n5266), .ZN(n4302) );
  NAND2_X1 U5316 ( .A1(n6211), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4301) );
  AOI21_X1 U5317 ( .B1(n4302), .B2(n4301), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n4305) );
  NOR2_X1 U5318 ( .A1(n4303), .A2(n4299), .ZN(n4304) );
  NOR2_X1 U5319 ( .A1(n4305), .A2(n4304), .ZN(n6244) );
  NAND3_X1 U5320 ( .A1(n6245), .A2(n6244), .A3(n6229), .ZN(n4307) );
  INV_X1 U5321 ( .A(n6329), .ZN(n4306) );
  NAND2_X1 U5322 ( .A1(n4307), .A2(n4306), .ZN(n4308) );
  NAND2_X1 U5323 ( .A1(n5703), .A2(n4308), .ZN(n6348) );
  NAND2_X1 U5324 ( .A1(n5917), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6011) );
  XNOR2_X1 U5325 ( .A(n5663), .B(n6011), .ZN(n4311) );
  INV_X1 U5326 ( .A(n2965), .ZN(n4497) );
  NOR2_X1 U5327 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6425), .ZN(n4343) );
  INV_X1 U5328 ( .A(n4343), .ZN(n6346) );
  AOI22_X1 U5329 ( .A1(n4311), .A2(n6345), .B1(n4497), .B2(n6346), .ZN(n4313)
         );
  NAND2_X1 U5330 ( .A1(n6352), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4312) );
  OAI21_X1 U5331 ( .B1(n6352), .B2(n4313), .A(n4312), .ZN(U3463) );
  AOI21_X1 U5332 ( .B1(n4339), .B2(n6363), .A(n6370), .ZN(n4314) );
  AOI22_X1 U5333 ( .A1(n4314), .A2(n6011), .B1(n5797), .B2(n6346), .ZN(n4316)
         );
  NAND2_X1 U5334 ( .A1(n6352), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4315) );
  OAI21_X1 U5335 ( .B1(n6352), .B2(n4316), .A(n4315), .ZN(U3464) );
  XNOR2_X1 U5336 ( .A(n4317), .B(n4318), .ZN(n5531) );
  OR2_X1 U5337 ( .A1(n4319), .A2(n4334), .ZN(n4321) );
  NAND2_X1 U5338 ( .A1(n4321), .A2(n4320), .ZN(n5611) );
  OAI22_X1 U5339 ( .A1(n5178), .A2(n5611), .B1(n5398), .B2(n5360), .ZN(n4322)
         );
  INV_X1 U5340 ( .A(n4322), .ZN(n4323) );
  OAI21_X1 U5341 ( .B1(n5531), .B2(n4891), .A(n4323), .ZN(U2855) );
  CLKBUF_X1 U5342 ( .A(n4325), .Z(n4326) );
  OAI21_X1 U5343 ( .B1(n4324), .B2(n4327), .A(n4326), .ZN(n5623) );
  INV_X1 U5344 ( .A(n4317), .ZN(n4329) );
  AOI21_X1 U5345 ( .B1(n4328), .B2(n4251), .A(n4329), .ZN(n4333) );
  NOR2_X1 U5346 ( .A1(n5612), .A2(n6281), .ZN(n5621) );
  AOI21_X1 U5347 ( .B1(n5536), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5621), 
        .ZN(n4330) );
  OAI21_X1 U5348 ( .B1(n4500), .B2(n5546), .A(n4330), .ZN(n4331) );
  AOI21_X1 U5349 ( .B1(n4333), .B2(n5702), .A(n4331), .ZN(n4332) );
  OAI21_X1 U5350 ( .B1(n5555), .B2(n5623), .A(n4332), .ZN(U2983) );
  INV_X1 U5351 ( .A(n4333), .ZN(n4510) );
  AOI21_X1 U5352 ( .B1(n4336), .B2(n4335), .A(n4334), .ZN(n5622) );
  AOI22_X1 U5353 ( .A1(n5393), .A2(n5622), .B1(EBX_REG_3__SCAN_IN), .B2(n4889), 
        .ZN(n4337) );
  OAI21_X1 U5354 ( .B1(n4510), .B2(n4891), .A(n4337), .ZN(U2856) );
  AND2_X1 U5355 ( .A1(n6345), .A2(n6363), .ZN(n5919) );
  INV_X1 U5356 ( .A(n5919), .ZN(n6151) );
  INV_X1 U5357 ( .A(n3526), .ZN(n4345) );
  AND2_X1 U5358 ( .A1(n4338), .A2(n4339), .ZN(n4340) );
  NAND2_X1 U5359 ( .A1(n5663), .A2(n4340), .ZN(n6072) );
  INV_X1 U5360 ( .A(n6072), .ZN(n4341) );
  NAND2_X1 U5361 ( .A1(n4341), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6076) );
  NAND2_X1 U5362 ( .A1(n6076), .A2(n6012), .ZN(n5766) );
  NAND2_X1 U5363 ( .A1(n5663), .A2(n4342), .ZN(n5882) );
  NOR2_X1 U5364 ( .A1(n5882), .A2(n6011), .ZN(n5883) );
  NOR2_X1 U5365 ( .A1(n5766), .A2(n5883), .ZN(n4344) );
  OAI222_X1 U5366 ( .A1(n6151), .A2(n4345), .B1(n6370), .B2(n4344), .C1(n4343), 
        .C2(n6103), .ZN(n4346) );
  NAND2_X1 U5367 ( .A1(n4346), .A2(n6348), .ZN(n4347) );
  OAI21_X1 U5368 ( .B1(n3479), .B2(n6348), .A(n4347), .ZN(U3462) );
  INV_X1 U5369 ( .A(DATAI_4_), .ZN(n5689) );
  INV_X1 U5370 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5479) );
  OAI222_X1 U5371 ( .A1(n5182), .A2(n5531), .B1(n4402), .B2(n5689), .C1(n4894), 
        .C2(n5479), .ZN(U2887) );
  INV_X1 U5372 ( .A(DATAI_2_), .ZN(n5678) );
  INV_X1 U5373 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5474) );
  OAI222_X1 U5374 ( .A1(n5537), .A2(n5182), .B1(n4402), .B2(n5678), .C1(n4894), 
        .C2(n5474), .ZN(U2889) );
  INV_X1 U5375 ( .A(DATAI_3_), .ZN(n5683) );
  INV_X1 U5376 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6489) );
  OAI222_X1 U5377 ( .A1(n4510), .A2(n5182), .B1(n4402), .B2(n5683), .C1(n4894), 
        .C2(n6489), .ZN(U2888) );
  INV_X1 U5378 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5465) );
  AOI22_X1 U5379 ( .A1(n6237), .A2(UWORD_REG_14__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4348) );
  OAI21_X1 U5380 ( .B1(n5465), .B2(n4359), .A(n4348), .ZN(U2893) );
  INV_X1 U5381 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5444) );
  AOI22_X1 U5382 ( .A1(n6237), .A2(UWORD_REG_6__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4349) );
  OAI21_X1 U5383 ( .B1(n5444), .B2(n4359), .A(n4349), .ZN(U2901) );
  INV_X1 U5384 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5446) );
  AOI22_X1 U5385 ( .A1(n6237), .A2(UWORD_REG_7__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4350) );
  OAI21_X1 U5386 ( .B1(n5446), .B2(n4359), .A(n4350), .ZN(U2900) );
  AOI22_X1 U5387 ( .A1(n6237), .A2(UWORD_REG_9__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4351) );
  OAI21_X1 U5388 ( .B1(n3876), .B2(n4359), .A(n4351), .ZN(U2898) );
  INV_X1 U5389 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5456) );
  AOI22_X1 U5390 ( .A1(n6237), .A2(UWORD_REG_11__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4352) );
  OAI21_X1 U5391 ( .B1(n5456), .B2(n4359), .A(n4352), .ZN(U2896) );
  INV_X1 U5392 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6441) );
  AOI22_X1 U5393 ( .A1(n6237), .A2(UWORD_REG_5__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4353) );
  OAI21_X1 U5394 ( .B1(n6441), .B2(n4359), .A(n4353), .ZN(U2902) );
  INV_X1 U5395 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5433) );
  AOI22_X1 U5396 ( .A1(n6237), .A2(UWORD_REG_0__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4354) );
  OAI21_X1 U5397 ( .B1(n5433), .B2(n4359), .A(n4354), .ZN(U2907) );
  INV_X1 U5398 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5435) );
  AOI22_X1 U5399 ( .A1(n6237), .A2(UWORD_REG_1__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4355) );
  OAI21_X1 U5400 ( .B1(n5435), .B2(n4359), .A(n4355), .ZN(U2906) );
  INV_X1 U5401 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5437) );
  AOI22_X1 U5402 ( .A1(n6237), .A2(UWORD_REG_2__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4356) );
  OAI21_X1 U5403 ( .B1(n5437), .B2(n4359), .A(n4356), .ZN(U2905) );
  INV_X1 U5404 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5439) );
  AOI22_X1 U5405 ( .A1(n6237), .A2(UWORD_REG_3__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4357) );
  OAI21_X1 U5406 ( .B1(n5439), .B2(n4359), .A(n4357), .ZN(U2904) );
  AOI22_X1 U5407 ( .A1(n6237), .A2(UWORD_REG_4__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4358) );
  OAI21_X1 U5408 ( .B1(n3775), .B2(n4359), .A(n4358), .ZN(U2903) );
  NAND2_X1 U5409 ( .A1(n4360), .A2(n4361), .ZN(n4400) );
  OAI21_X1 U5410 ( .B1(n4360), .B2(n4361), .A(n4400), .ZN(n4534) );
  INV_X1 U5411 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4364) );
  OAI21_X1 U5412 ( .B1(n4363), .B2(n4362), .A(n4376), .ZN(n5602) );
  OAI222_X1 U5413 ( .A1(n4534), .A2(n4891), .B1(n5398), .B2(n4364), .C1(n5602), 
        .C2(n5178), .ZN(U2854) );
  INV_X1 U5414 ( .A(DATAI_5_), .ZN(n5696) );
  INV_X1 U5415 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5482) );
  OAI222_X1 U5416 ( .A1(n4534), .A2(n5182), .B1(n4402), .B2(n5696), .C1(n4894), 
        .C2(n5482), .ZN(U2886) );
  OAI21_X1 U5417 ( .B1(n4367), .B2(n4366), .A(n4365), .ZN(n5601) );
  INV_X1 U5418 ( .A(n4534), .ZN(n4370) );
  AOI22_X1 U5419 ( .A1(n5536), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n5630), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4368) );
  OAI21_X1 U5420 ( .B1(n4527), .B2(n5546), .A(n4368), .ZN(n4369) );
  AOI21_X1 U5421 ( .B1(n4370), .B2(n5702), .A(n4369), .ZN(n4371) );
  OAI21_X1 U5422 ( .B1(n5601), .B2(n5555), .A(n4371), .ZN(U2981) );
  OAI21_X1 U5423 ( .B1(n4374), .B2(n4373), .A(n4372), .ZN(n5521) );
  AND2_X1 U5424 ( .A1(n4376), .A2(n4375), .ZN(n4377) );
  OR2_X1 U5425 ( .A1(n4377), .A2(n4457), .ZN(n5348) );
  NOR2_X1 U5426 ( .A1(n5585), .A2(n5348), .ZN(n4387) );
  NAND2_X1 U5427 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5610), .ZN(n4379)
         );
  INV_X1 U5428 ( .A(n4378), .ZN(n5633) );
  AOI21_X1 U5429 ( .B1(n5633), .B2(n5639), .A(n5632), .ZN(n5563) );
  NOR2_X1 U5430 ( .A1(n5634), .A2(n5563), .ZN(n5625) );
  INV_X1 U5431 ( .A(n5625), .ZN(n5609) );
  NOR2_X1 U5432 ( .A1(n4379), .A2(n5609), .ZN(n4385) );
  OAI22_X1 U5433 ( .A1(n5079), .A2(n5633), .B1(n5632), .B2(n4381), .ZN(n5635)
         );
  OAI21_X1 U5434 ( .B1(n5634), .B2(n6456), .A(n5632), .ZN(n4382) );
  OAI21_X1 U5435 ( .B1(n5572), .B2(n5610), .A(n4382), .ZN(n4383) );
  AOI211_X1 U5436 ( .C1(n5639), .C2(n6456), .A(n5635), .B(n4383), .ZN(n5608)
         );
  INV_X1 U5437 ( .A(n5608), .ZN(n4384) );
  MUX2_X1 U5438 ( .A(n4385), .B(n4384), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4386) );
  AOI211_X1 U5439 ( .C1(n5630), .C2(REIP_REG_6__SCAN_IN), .A(n4387), .B(n4386), 
        .ZN(n4388) );
  OAI21_X1 U5440 ( .B1(n5654), .B2(n5521), .A(n4388), .ZN(U3012) );
  INV_X1 U5441 ( .A(DATAI_6_), .ZN(n5442) );
  XOR2_X1 U5442 ( .A(n4399), .B(n4400), .Z(n5522) );
  INV_X1 U5443 ( .A(n5522), .ZN(n4396) );
  OAI222_X1 U5444 ( .A1(n5442), .A2(n4402), .B1(n5182), .B2(n4396), .C1(n4389), 
        .C2(n4894), .ZN(U2885) );
  AND2_X1 U5445 ( .A1(n4391), .A2(n4392), .ZN(n4412) );
  OR2_X1 U5446 ( .A1(n4412), .A2(n4393), .ZN(n4394) );
  NAND2_X1 U5447 ( .A1(n4390), .A2(n4394), .ZN(n5338) );
  AOI22_X1 U5448 ( .A1(n4606), .A2(DATAI_9_), .B1(n5408), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4395) );
  OAI21_X1 U5449 ( .B1(n5338), .B2(n5182), .A(n4395), .ZN(U2882) );
  INV_X1 U5450 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4397) );
  OAI222_X1 U5451 ( .A1(n5348), .A2(n5178), .B1(n4397), .B2(n5398), .C1(n4891), 
        .C2(n4396), .ZN(U2853) );
  OR2_X1 U5452 ( .A1(n4400), .A2(n4399), .ZN(n4401) );
  XOR2_X1 U5453 ( .A(n4398), .B(n4401), .Z(n4409) );
  INV_X1 U5454 ( .A(n4409), .ZN(n4487) );
  INV_X1 U5455 ( .A(DATAI_7_), .ZN(n6479) );
  OAI222_X1 U5456 ( .A1(n5182), .A2(n4487), .B1(n4402), .B2(n6479), .C1(n4894), 
        .C2(n3510), .ZN(U2884) );
  OAI21_X1 U5457 ( .B1(n4405), .B2(n4404), .A(n4403), .ZN(n5595) );
  INV_X1 U5458 ( .A(REIP_REG_7__SCAN_IN), .ZN(n4406) );
  NOR2_X1 U5459 ( .A1(n5612), .A2(n4406), .ZN(n5593) );
  AOI21_X1 U5460 ( .B1(n5536), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5593), 
        .ZN(n4407) );
  OAI21_X1 U5461 ( .B1(n4478), .B2(n5546), .A(n4407), .ZN(n4408) );
  AOI21_X1 U5462 ( .B1(n4409), .B2(n5702), .A(n4408), .ZN(n4410) );
  OAI21_X1 U5463 ( .B1(n5595), .B2(n5555), .A(n4410), .ZN(U2979) );
  INV_X1 U5464 ( .A(n4411), .ZN(n4414) );
  NAND2_X1 U5465 ( .A1(n4360), .A2(n4391), .ZN(n4413) );
  AOI21_X1 U5466 ( .B1(n4414), .B2(n4413), .A(n4412), .ZN(n4474) );
  INV_X1 U5467 ( .A(n4474), .ZN(n4467) );
  AOI22_X1 U5468 ( .A1(n4606), .A2(DATAI_8_), .B1(n5408), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4415) );
  OAI21_X1 U5469 ( .B1(n4467), .B2(n5182), .A(n4415), .ZN(U2883) );
  INV_X1 U5470 ( .A(n4390), .ZN(n4418) );
  OAI21_X1 U5471 ( .B1(n4418), .B2(n3613), .A(n4520), .ZN(n4565) );
  AND2_X1 U5472 ( .A1(n4420), .A2(n4419), .ZN(n6257) );
  NOR3_X1 U5473 ( .A1(n6366), .A2(n6331), .A3(n6365), .ZN(n6246) );
  NOR2_X1 U5474 ( .A1(n6257), .A2(n6246), .ZN(n4421) );
  INV_X1 U5475 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4698) );
  INV_X1 U5476 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4711) );
  INV_X1 U5477 ( .A(n4704), .ZN(n4425) );
  NAND2_X1 U5478 ( .A1(n4425), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4426) );
  INV_X1 U5479 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6292) );
  INV_X1 U5480 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6288) );
  INV_X1 U5481 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4525) );
  INV_X1 U5482 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6281) );
  INV_X1 U5483 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6279) );
  NOR3_X1 U5484 ( .A1(n6353), .A2(n6281), .A3(n6279), .ZN(n5356) );
  NAND2_X1 U5485 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5356), .ZN(n4526) );
  NOR2_X1 U5486 ( .A1(n4525), .A2(n4526), .ZN(n5345) );
  NAND2_X1 U5487 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5345), .ZN(n4444) );
  NOR3_X1 U5488 ( .A1(n6288), .A2(n4406), .A3(n4444), .ZN(n4548) );
  INV_X1 U5489 ( .A(n4548), .ZN(n4430) );
  NAND2_X1 U5490 ( .A1(n3178), .A2(n6363), .ZN(n4427) );
  NOR2_X1 U5491 ( .A1(n4428), .A2(n4427), .ZN(n4429) );
  INV_X1 U5492 ( .A(n5371), .ZN(n4617) );
  INV_X1 U5493 ( .A(n4723), .ZN(n4812) );
  OAI21_X1 U5494 ( .B1(n5371), .B2(n4430), .A(n4812), .ZN(n5336) );
  NOR2_X2 U5495 ( .A1(n5371), .A2(n5115), .ZN(n5344) );
  AOI21_X1 U5496 ( .B1(n5364), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5344), 
        .ZN(n4442) );
  NAND3_X1 U5497 ( .A1(n6271), .A2(n6363), .A3(n4431), .ZN(n6238) );
  INV_X1 U5498 ( .A(n6238), .ZN(n4433) );
  INV_X1 U5499 ( .A(EBX_REG_31__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U5500 ( .A1(n6271), .A2(n6363), .ZN(n4437) );
  NAND3_X1 U5501 ( .A1(n3178), .A2(n4821), .A3(n4437), .ZN(n4432) );
  OAI21_X1 U5502 ( .B1(n4434), .B2(n4433), .A(n4432), .ZN(n4435) );
  INV_X1 U5503 ( .A(n4435), .ZN(n4436) );
  NOR2_X2 U5504 ( .A1(n4496), .A2(n4436), .ZN(n5368) );
  NAND3_X1 U5505 ( .A1(n4438), .A2(EBX_REG_31__SCAN_IN), .A3(n4437), .ZN(n4439) );
  NOR2_X2 U5506 ( .A1(n4496), .A2(n4439), .ZN(n5377) );
  XOR2_X1 U5507 ( .A(n5334), .B(n4440), .Z(n5567) );
  AOI22_X1 U5508 ( .A1(EBX_REG_10__SCAN_IN), .A2(n5368), .B1(n5377), .B2(n5567), .ZN(n4441) );
  OAI211_X1 U5509 ( .C1(n6292), .C2(n5336), .A(n4442), .B(n4441), .ZN(n4449)
         );
  NAND2_X1 U5510 ( .A1(n4704), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4443) );
  NOR2_X1 U5511 ( .A1(n4618), .A2(n4444), .ZN(n4477) );
  NOR2_X1 U5512 ( .A1(n6288), .A2(n4406), .ZN(n4445) );
  AND2_X1 U5513 ( .A1(n4477), .A2(n4445), .ZN(n5330) );
  NAND2_X1 U5514 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n4446) );
  OAI211_X1 U5515 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n5330), .B(n4446), .ZN(n4447) );
  OAI21_X1 U5516 ( .B1(n5386), .B2(n4561), .A(n4447), .ZN(n4448) );
  NOR2_X1 U5517 ( .A1(n4449), .A2(n4448), .ZN(n4450) );
  OAI21_X1 U5518 ( .B1(n4565), .B2(n5164), .A(n4450), .ZN(U2817) );
  AOI22_X1 U5519 ( .A1(n5393), .A2(n5567), .B1(EBX_REG_10__SCAN_IN), .B2(n4889), .ZN(n4451) );
  OAI21_X1 U5520 ( .B1(n4565), .B2(n4891), .A(n4451), .ZN(U2849) );
  AOI22_X1 U5521 ( .A1(n4606), .A2(DATAI_10_), .B1(n5408), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4452) );
  OAI21_X1 U5522 ( .B1(n4565), .B2(n5182), .A(n4452), .ZN(U2881) );
  INV_X1 U5523 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6527) );
  NOR2_X1 U5524 ( .A1(n4453), .A2(n4454), .ZN(n4455) );
  OR2_X1 U5525 ( .A1(n5332), .A2(n4455), .ZN(n5586) );
  OAI222_X1 U5526 ( .A1(n4467), .A2(n4891), .B1(n5398), .B2(n6527), .C1(n5586), 
        .C2(n5178), .ZN(U2851) );
  NOR2_X1 U5527 ( .A1(n4457), .A2(n4456), .ZN(n4458) );
  OR2_X1 U5528 ( .A1(n4453), .A2(n4458), .ZN(n4480) );
  INV_X1 U5529 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4459) );
  OAI222_X1 U5530 ( .A1(n4480), .A2(n5178), .B1(n4459), .B2(n5398), .C1(n4891), 
        .C2(n4487), .ZN(U2852) );
  INV_X1 U5531 ( .A(n4472), .ZN(n4462) );
  AOI22_X1 U5532 ( .A1(EBX_REG_8__SCAN_IN), .A2(n5368), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n5364), .ZN(n4460) );
  INV_X1 U5533 ( .A(n5344), .ZN(n5359) );
  OAI211_X1 U5534 ( .C1(n5367), .C2(n5586), .A(n4460), .B(n5359), .ZN(n4461)
         );
  AOI21_X1 U5535 ( .B1(n5340), .B2(n4462), .A(n4461), .ZN(n4466) );
  NAND2_X1 U5536 ( .A1(REIP_REG_7__SCAN_IN), .A2(n4477), .ZN(n4463) );
  AOI21_X1 U5537 ( .B1(n6288), .B2(n4463), .A(n5336), .ZN(n4464) );
  INV_X1 U5538 ( .A(n4464), .ZN(n4465) );
  OAI211_X1 U5539 ( .C1(n4467), .C2(n5164), .A(n4466), .B(n4465), .ZN(U2819)
         );
  OAI21_X1 U5540 ( .B1(n4468), .B2(n4470), .A(n4469), .ZN(n5584) );
  AOI22_X1 U5541 ( .A1(n5536), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n5630), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4471) );
  OAI21_X1 U5542 ( .B1(n4472), .B2(n5546), .A(n4471), .ZN(n4473) );
  AOI21_X1 U5543 ( .B1(n4474), .B2(n5702), .A(n4473), .ZN(n4475) );
  OAI21_X1 U5544 ( .B1(n5584), .B2(n5555), .A(n4475), .ZN(U2978) );
  INV_X1 U5545 ( .A(n5345), .ZN(n4476) );
  AOI21_X1 U5546 ( .B1(n5357), .B2(n4476), .A(n5371), .ZN(n4524) );
  OAI21_X1 U5547 ( .B1(REIP_REG_6__SCAN_IN), .B2(n4618), .A(n4524), .ZN(n4485)
         );
  INV_X1 U5548 ( .A(n4477), .ZN(n4479) );
  OAI22_X1 U5549 ( .A1(n4479), .A2(REIP_REG_7__SCAN_IN), .B1(n4478), .B2(n5386), .ZN(n4484) );
  INV_X1 U5550 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4482) );
  INV_X1 U5551 ( .A(n4480), .ZN(n5594) );
  AOI22_X1 U5552 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5368), .B1(n5377), .B2(n5594), 
        .ZN(n4481) );
  OAI211_X1 U5553 ( .C1(n5374), .C2(n4482), .A(n4481), .B(n5359), .ZN(n4483)
         );
  AOI211_X1 U5554 ( .C1(REIP_REG_7__SCAN_IN), .C2(n4485), .A(n4484), .B(n4483), 
        .ZN(n4486) );
  OAI21_X1 U5555 ( .B1(n4487), .B2(n5164), .A(n4486), .ZN(U2820) );
  NAND2_X1 U5556 ( .A1(n4709), .A2(n3448), .ZN(n4488) );
  OR2_X1 U5557 ( .A1(n4618), .A2(REIP_REG_1__SCAN_IN), .ZN(n5370) );
  NOR2_X1 U5558 ( .A1(n5371), .A2(n6279), .ZN(n4489) );
  AND2_X1 U5559 ( .A1(n5370), .A2(n4489), .ZN(n4491) );
  AOI21_X1 U5560 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5357), .A(
        REIP_REG_2__SCAN_IN), .ZN(n4490) );
  OAI22_X1 U5561 ( .A1(n4491), .A2(n4490), .B1(n5545), .B2(n5386), .ZN(n4494)
         );
  NOR2_X1 U5562 ( .A1(n5374), .A2(n4492), .ZN(n4493) );
  AOI211_X1 U5563 ( .C1(EBX_REG_2__SCAN_IN), .C2(n5368), .A(n4494), .B(n4493), 
        .ZN(n4499) );
  NOR2_X1 U5564 ( .A1(n4496), .A2(n4495), .ZN(n5378) );
  AOI22_X1 U5565 ( .A1(n4497), .A2(n5378), .B1(n5377), .B2(n5631), .ZN(n4498)
         );
  OAI211_X1 U5566 ( .C1(n5537), .C2(n5382), .A(n4499), .B(n4498), .ZN(U2825)
         );
  OAI21_X1 U5567 ( .B1(n4618), .B2(n5356), .A(n4617), .ZN(n5355) );
  AOI22_X1 U5568 ( .A1(n5377), .A2(n5622), .B1(n5368), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4507) );
  OAI22_X1 U5569 ( .A1(n4501), .A2(n5374), .B1(n5386), .B2(n4500), .ZN(n4502)
         );
  INV_X1 U5570 ( .A(n4502), .ZN(n4506) );
  INV_X1 U5571 ( .A(n5356), .ZN(n4503) );
  NAND4_X1 U5572 ( .A1(n5357), .A2(REIP_REG_2__SCAN_IN), .A3(n4503), .A4(
        REIP_REG_1__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5573 ( .A1(n5378), .A2(n4264), .ZN(n4504) );
  NAND4_X1 U5574 ( .A1(n4507), .A2(n4506), .A3(n4505), .A4(n4504), .ZN(n4508)
         );
  AOI21_X1 U5575 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5355), .A(n4508), .ZN(n4509)
         );
  OAI21_X1 U5576 ( .B1(n4510), .B2(n5382), .A(n4509), .ZN(U2824) );
  INV_X1 U5577 ( .A(n5378), .ZN(n4517) );
  INV_X1 U5578 ( .A(n5382), .ZN(n4511) );
  AOI22_X1 U5579 ( .A1(n4812), .A2(REIP_REG_0__SCAN_IN), .B1(n4511), .B2(n5553), .ZN(n4516) );
  NAND2_X1 U5580 ( .A1(n5374), .A2(n5386), .ZN(n4514) );
  OAI22_X1 U5581 ( .A1(n4512), .A2(n5361), .B1(n5367), .B2(n5644), .ZN(n4513)
         );
  AOI21_X1 U5582 ( .B1(n4514), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n4513), 
        .ZN(n4515) );
  OAI211_X1 U5583 ( .C1(n5948), .C2(n4517), .A(n4516), .B(n4515), .ZN(U2827)
         );
  AND2_X1 U5584 ( .A1(n4520), .A2(n4519), .ZN(n4521) );
  NOR2_X1 U5585 ( .A1(n4518), .A2(n4521), .ZN(n5518) );
  INV_X1 U5586 ( .A(n5518), .ZN(n4523) );
  AOI22_X1 U5587 ( .A1(n4606), .A2(DATAI_11_), .B1(n5408), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4522) );
  OAI21_X1 U5588 ( .B1(n4523), .B2(n5182), .A(n4522), .ZN(U2880) );
  INV_X1 U5589 ( .A(n4524), .ZN(n5350) );
  OAI21_X1 U5590 ( .B1(n4618), .B2(n4526), .A(n4525), .ZN(n4532) );
  INV_X1 U5591 ( .A(n4527), .ZN(n4529) );
  OAI22_X1 U5592 ( .A1(n6431), .A2(n5374), .B1(n5367), .B2(n5602), .ZN(n4528)
         );
  AOI211_X1 U5593 ( .C1(n5340), .C2(n4529), .A(n5344), .B(n4528), .ZN(n4530)
         );
  OAI21_X1 U5594 ( .B1(n5361), .B2(n4364), .A(n4530), .ZN(n4531) );
  AOI21_X1 U5595 ( .B1(n5350), .B2(n4532), .A(n4531), .ZN(n4533) );
  OAI21_X1 U5596 ( .B1(n4534), .B2(n5382), .A(n4533), .ZN(U2822) );
  XOR2_X1 U5597 ( .A(n4535), .B(n4518), .Z(n4590) );
  OR2_X1 U5598 ( .A1(n4536), .A2(n5321), .ZN(n4537) );
  NAND2_X1 U5599 ( .A1(n4537), .A2(n5255), .ZN(n4592) );
  OAI22_X1 U5600 ( .A1(n5178), .A2(n4592), .B1(n5398), .B2(n6413), .ZN(n4538)
         );
  AOI21_X1 U5601 ( .B1(n4590), .B2(n5394), .A(n4538), .ZN(n4539) );
  INV_X1 U5602 ( .A(n4539), .ZN(U2847) );
  NAND2_X1 U5603 ( .A1(n4542), .A2(n4541), .ZN(n4543) );
  XNOR2_X1 U5604 ( .A(n4540), .B(n4543), .ZN(n5580) );
  NAND2_X1 U5605 ( .A1(n5580), .A2(n5541), .ZN(n4546) );
  NOR2_X1 U5606 ( .A1(n5612), .A2(n6290), .ZN(n5577) );
  AND2_X1 U5607 ( .A1(n5536), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4544)
         );
  AOI211_X1 U5608 ( .C1(n5339), .C2(n5517), .A(n5577), .B(n4544), .ZN(n4545)
         );
  OAI211_X1 U5609 ( .C1(n5692), .C2(n5338), .A(n4546), .B(n4545), .ZN(U2977)
         );
  INV_X1 U5610 ( .A(n4590), .ZN(n4557) );
  AOI22_X1 U5611 ( .A1(n4606), .A2(DATAI_12_), .B1(n5408), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4547) );
  OAI21_X1 U5612 ( .B1(n4557), .B2(n5182), .A(n4547), .ZN(U2879) );
  NAND4_X1 U5613 ( .A1(REIP_REG_11__SCAN_IN), .A2(n4548), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n4615) );
  INV_X1 U5614 ( .A(n4615), .ZN(n4549) );
  OR2_X1 U5615 ( .A1(n4618), .A2(n4549), .ZN(n4550) );
  NAND2_X1 U5616 ( .A1(n4550), .A2(n4617), .ZN(n5324) );
  OAI22_X1 U5617 ( .A1(n4551), .A2(n5374), .B1(n5367), .B2(n4592), .ZN(n4553)
         );
  NOR2_X1 U5618 ( .A1(n6413), .A2(n5361), .ZN(n4552) );
  NOR3_X1 U5619 ( .A1(n5344), .A2(n4553), .A3(n4552), .ZN(n4554) );
  OAI21_X1 U5620 ( .B1(n5386), .B2(n4588), .A(n4554), .ZN(n4555) );
  NOR3_X1 U5621 ( .A1(n4618), .A2(REIP_REG_12__SCAN_IN), .A3(n4615), .ZN(n5317) );
  AOI211_X1 U5622 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5324), .A(n4555), .B(n5317), .ZN(n4556) );
  OAI21_X1 U5623 ( .B1(n4557), .B2(n5164), .A(n4556), .ZN(U2815) );
  NAND2_X1 U5624 ( .A1(n5513), .A2(n4559), .ZN(n4560) );
  XNOR2_X1 U5625 ( .A(n4558), .B(n4560), .ZN(n5573) );
  NAND2_X1 U5626 ( .A1(n5573), .A2(n5541), .ZN(n4564) );
  NOR2_X1 U5627 ( .A1(n5612), .A2(n6292), .ZN(n5566) );
  NOR2_X1 U5628 ( .A1(n5546), .A2(n4561), .ZN(n4562) );
  AOI211_X1 U5629 ( .C1(n5536), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5566), 
        .B(n4562), .ZN(n4563) );
  OAI211_X1 U5630 ( .C1(n5692), .C2(n4565), .A(n4564), .B(n4563), .ZN(U2976)
         );
  NAND2_X1 U5631 ( .A1(n4566), .A2(n4567), .ZN(n4568) );
  AND2_X1 U5632 ( .A1(n4569), .A2(n4568), .ZN(n5388) );
  INV_X1 U5633 ( .A(n5388), .ZN(n4571) );
  AOI22_X1 U5634 ( .A1(n4606), .A2(DATAI_13_), .B1(n5408), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n4570) );
  OAI21_X1 U5635 ( .B1(n4571), .B2(n5182), .A(n4570), .ZN(U2878) );
  INV_X1 U5636 ( .A(n4574), .ZN(n4575) );
  NAND2_X1 U5637 ( .A1(n2960), .A2(n4575), .ZN(n4576) );
  NAND2_X1 U5638 ( .A1(n4572), .A2(n4576), .ZN(n5306) );
  AOI22_X1 U5639 ( .A1(n4606), .A2(DATAI_14_), .B1(n5408), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n4577) );
  OAI21_X1 U5640 ( .B1(n5306), .B2(n5182), .A(n4577), .ZN(U2877) );
  INV_X1 U5641 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4580) );
  INV_X1 U5642 ( .A(n4609), .ZN(n4578) );
  OAI21_X1 U5643 ( .B1(n5258), .B2(n4579), .A(n4578), .ZN(n5303) );
  OAI222_X1 U5644 ( .A1(n5306), .A2(n4891), .B1(n4580), .B2(n5398), .C1(n5178), 
        .C2(n5303), .ZN(U2845) );
  INV_X1 U5645 ( .A(n4582), .ZN(n4583) );
  NOR2_X1 U5646 ( .A1(n4584), .A2(n4583), .ZN(n4585) );
  XNOR2_X1 U5647 ( .A(n4581), .B(n4585), .ZN(n4603) );
  INV_X1 U5648 ( .A(REIP_REG_12__SCAN_IN), .ZN(n4586) );
  NOR2_X1 U5649 ( .A1(n5612), .A2(n4586), .ZN(n4600) );
  AOI21_X1 U5650 ( .B1(n5536), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n4600), 
        .ZN(n4587) );
  OAI21_X1 U5651 ( .B1(n4588), .B2(n5546), .A(n4587), .ZN(n4589) );
  AOI21_X1 U5652 ( .B1(n4590), .B2(n5702), .A(n4589), .ZN(n4591) );
  OAI21_X1 U5653 ( .B1(n4603), .B2(n5555), .A(n4591), .ZN(U2974) );
  INV_X1 U5654 ( .A(n4592), .ZN(n4601) );
  NOR2_X1 U5655 ( .A1(n5264), .A2(n3422), .ZN(n4598) );
  INV_X1 U5656 ( .A(n4593), .ZN(n5243) );
  AOI22_X1 U5657 ( .A1(n5571), .A2(n5243), .B1(n5569), .B2(n4594), .ZN(n4595)
         );
  INV_X1 U5658 ( .A(n4595), .ZN(n5558) );
  AOI221_X1 U5659 ( .B1(n5632), .B2(n3422), .C1(n5222), .C2(n3422), .A(n5558), 
        .ZN(n4596) );
  INV_X1 U5660 ( .A(n4596), .ZN(n4597) );
  MUX2_X1 U5661 ( .A(n4598), .B(n4597), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n4599) );
  AOI211_X1 U5662 ( .C1(n5649), .C2(n4601), .A(n4600), .B(n4599), .ZN(n4602)
         );
  OAI21_X1 U5663 ( .B1(n4603), .B2(n5654), .A(n4602), .ZN(U3006) );
  OAI21_X1 U5664 ( .B1(n4605), .B2(n4604), .A(n2976), .ZN(n4995) );
  AOI22_X1 U5665 ( .A1(n4606), .A2(DATAI_15_), .B1(n5408), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n4607) );
  OAI21_X1 U5666 ( .B1(n4995), .B2(n5182), .A(n4607), .ZN(U2876) );
  OAI21_X1 U5667 ( .B1(n4609), .B2(n4608), .A(n4810), .ZN(n4613) );
  OAI22_X1 U5668 ( .A1(n5178), .A2(n4613), .B1(n4610), .B2(n5398), .ZN(n4611)
         );
  INV_X1 U5669 ( .A(n4611), .ZN(n4612) );
  OAI21_X1 U5670 ( .B1(n4995), .B2(n4891), .A(n4612), .ZN(U2844) );
  INV_X1 U5671 ( .A(n4613), .ZN(n5236) );
  INV_X1 U5672 ( .A(n4992), .ZN(n4614) );
  OAI22_X1 U5673 ( .A1(n5361), .A2(n4610), .B1(n4614), .B2(n5386), .ZN(n4622)
         );
  NOR2_X1 U5674 ( .A1(n4586), .A2(n4615), .ZN(n5302) );
  NAND3_X1 U5675 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        n5302), .ZN(n4712) );
  INV_X1 U5676 ( .A(n4712), .ZN(n4616) );
  NAND2_X1 U5677 ( .A1(n4617), .A2(n4616), .ZN(n4813) );
  NAND2_X1 U5678 ( .A1(n4812), .A2(n4813), .ZN(n5312) );
  INV_X1 U5679 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6440) );
  NOR3_X1 U5680 ( .A1(n4618), .A2(REIP_REG_15__SCAN_IN), .A3(n4712), .ZN(n4619) );
  AOI211_X1 U5681 ( .C1(n5364), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5344), 
        .B(n4619), .ZN(n4620) );
  OAI21_X1 U5682 ( .B1(n5312), .B2(n6440), .A(n4620), .ZN(n4621) );
  AOI211_X1 U5683 ( .C1(n5236), .C2(n5377), .A(n4622), .B(n4621), .ZN(n4623)
         );
  OAI21_X1 U5684 ( .B1(n4995), .B2(n5164), .A(n4623), .ZN(U2812) );
  XNOR2_X1 U5685 ( .A(n5203), .B(n4625), .ZN(n4626) );
  XNOR2_X1 U5686 ( .A(n2964), .B(n4626), .ZN(n5248) );
  INV_X1 U5687 ( .A(REIP_REG_14__SCAN_IN), .ZN(n4627) );
  OAI22_X1 U5688 ( .A1(n5550), .A2(n5304), .B1(n5612), .B2(n4627), .ZN(n4628)
         );
  AOI21_X1 U5689 ( .B1(n5517), .B2(n5307), .A(n4628), .ZN(n4630) );
  OR2_X1 U5690 ( .A1(n5306), .A2(n5692), .ZN(n4629) );
  OAI211_X1 U5691 ( .C1(n5248), .C2(n5555), .A(n4630), .B(n4629), .ZN(U2972)
         );
  AOI22_X1 U5692 ( .A1(n3079), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4634) );
  AOI22_X1 U5693 ( .A1(n3672), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5694 ( .A1(n3281), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3912), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4632) );
  AOI22_X1 U5695 ( .A1(n4146), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4139), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4631) );
  NAND4_X1 U5696 ( .A1(n4634), .A2(n4633), .A3(n4632), .A4(n4631), .ZN(n4643)
         );
  AOI22_X1 U5697 ( .A1(n3118), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4641) );
  AOI22_X1 U5698 ( .A1(n4145), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n2967), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5699 ( .A1(n4635), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3844), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5700 ( .A1(n4637), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4636), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4638) );
  NAND4_X1 U5701 ( .A1(n4641), .A2(n4640), .A3(n4639), .A4(n4638), .ZN(n4642)
         );
  NOR2_X1 U5702 ( .A1(n4643), .A2(n4642), .ZN(n4647) );
  NOR2_X1 U5703 ( .A1(n4645), .A2(n4644), .ZN(n4646) );
  XOR2_X1 U5704 ( .A(n4647), .B(n4646), .Z(n4653) );
  NAND2_X1 U5705 ( .A1(n3558), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4648)
         );
  NAND2_X1 U5706 ( .A1(n4649), .A2(n4648), .ZN(n4650) );
  AOI21_X1 U5707 ( .B1(n3506), .B2(EAX_REG_30__SCAN_IN), .A(n4650), .ZN(n4651)
         );
  OAI21_X1 U5708 ( .B1(n4653), .B2(n4652), .A(n4651), .ZN(n4657) );
  XNOR2_X1 U5709 ( .A(n4654), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4732)
         );
  NAND2_X1 U5710 ( .A1(n4732), .A2(n4655), .ZN(n4656) );
  NAND2_X1 U5711 ( .A1(n4657), .A2(n4656), .ZN(n4695) );
  AOI22_X1 U5712 ( .A1(n4659), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4658), .ZN(n4660) );
  NAND3_X1 U5713 ( .A1(n4708), .A2(n3132), .A3(n4894), .ZN(n4663) );
  NOR2_X2 U5714 ( .A1(n5408), .A2(n4661), .ZN(n5405) );
  AOI22_X1 U5715 ( .A1(n5405), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5408), .ZN(n4662) );
  NAND2_X1 U5716 ( .A1(n4663), .A2(n4662), .ZN(U2860) );
  NAND2_X1 U5717 ( .A1(n4184), .A2(n2982), .ZN(n4666) );
  OAI22_X1 U5718 ( .A1(n6333), .A2(n4666), .B1(n4665), .B2(n4664), .ZN(n4667)
         );
  AOI21_X1 U5719 ( .B1(n4668), .B2(n6252), .A(n4667), .ZN(n4673) );
  INV_X1 U5720 ( .A(n6340), .ZN(n4672) );
  INV_X1 U5721 ( .A(n6333), .ZN(n4670) );
  INV_X1 U5722 ( .A(n4184), .ZN(n4669) );
  AOI21_X1 U5723 ( .B1(n4670), .B2(n4669), .A(n4672), .ZN(n4671) );
  OAI22_X1 U5724 ( .A1(n4673), .A2(n4672), .B1(n4671), .B2(n2982), .ZN(U3459)
         );
  INV_X1 U5725 ( .A(n4674), .ZN(n4675) );
  OAI211_X1 U5726 ( .C1(n4685), .C2(n4680), .A(n4679), .B(n4682), .ZN(n4687)
         );
  INV_X1 U5727 ( .A(n4682), .ZN(n4683) );
  OAI21_X1 U5728 ( .B1(n4681), .B2(n4869), .A(n4683), .ZN(n4684) );
  OR2_X1 U5729 ( .A1(n4685), .A2(n4684), .ZN(n4686) );
  NAND2_X1 U5730 ( .A1(n4997), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4688) );
  OAI211_X1 U5731 ( .C1(n5103), .C2(n5037), .A(n4688), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4689) );
  NAND2_X1 U5732 ( .A1(n5630), .A2(REIP_REG_30__SCAN_IN), .ZN(n4696) );
  OAI211_X1 U5733 ( .C1(n5585), .C2(n4823), .A(n4689), .B(n4696), .ZN(n4690)
         );
  OAI21_X1 U5734 ( .B1(n4701), .B2(n5654), .A(n4693), .ZN(U2988) );
  NAND2_X1 U5735 ( .A1(n5517), .A2(n4732), .ZN(n4697) );
  OAI211_X1 U5736 ( .C1(n5550), .C2(n4698), .A(n4697), .B(n4696), .ZN(n4699)
         );
  OAI21_X1 U5737 ( .B1(n4701), .B2(n5555), .A(n4700), .ZN(U2956) );
  AOI21_X1 U5738 ( .B1(n5536), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4702), 
        .ZN(n4703) );
  OAI21_X1 U5739 ( .B1(n5546), .B2(n4704), .A(n4703), .ZN(n4705) );
  AOI21_X1 U5740 ( .B1(n4708), .B2(n5702), .A(n4705), .ZN(n4706) );
  OAI21_X1 U5741 ( .B1(n4707), .B2(n5555), .A(n4706), .ZN(U2955) );
  INV_X1 U5742 ( .A(n4708), .ZN(n4730) );
  NAND4_X1 U5743 ( .A1(n4709), .A2(n6364), .A3(EBX_REG_31__SCAN_IN), .A4(n6238), .ZN(n4710) );
  OAI21_X1 U5744 ( .B1(n5374), .B2(n4711), .A(n4710), .ZN(n4725) );
  INV_X1 U5745 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U5746 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5155) );
  INV_X1 U5747 ( .A(n5155), .ZN(n4718) );
  NOR2_X1 U5748 ( .A1(n6440), .A2(n4712), .ZN(n4726) );
  NAND3_X1 U5749 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        n4726), .ZN(n4713) );
  NOR2_X1 U5750 ( .A1(n5371), .A2(n4713), .ZN(n4714) );
  OR2_X1 U5751 ( .A1(n4723), .A2(n4714), .ZN(n5295) );
  INV_X1 U5752 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6307) );
  INV_X1 U5753 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6305) );
  NOR2_X1 U5754 ( .A1(n6307), .A2(n6305), .ZN(n4715) );
  NAND2_X1 U5755 ( .A1(n4715), .A2(REIP_REG_18__SCAN_IN), .ZN(n4716) );
  NAND2_X1 U5756 ( .A1(n5357), .A2(n4716), .ZN(n4717) );
  NAND2_X1 U5757 ( .A1(n5295), .A2(n4717), .ZN(n5160) );
  INV_X1 U5758 ( .A(n5160), .ZN(n5171) );
  OAI221_X1 U5759 ( .B1(REIP_REG_23__SCAN_IN), .B2(n4723), .C1(n4718), .C2(
        n4723), .A(n5171), .ZN(n5146) );
  AND3_X1 U5760 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4776) );
  NOR2_X1 U5761 ( .A1(n4723), .A2(n4776), .ZN(n4719) );
  NOR2_X1 U5762 ( .A1(n5146), .A2(n4719), .ZN(n5118) );
  NAND2_X1 U5763 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4720) );
  NAND2_X1 U5764 ( .A1(n5357), .A2(n4720), .ZN(n4721) );
  NAND2_X1 U5765 ( .A1(n5118), .A2(n4721), .ZN(n4758) );
  AOI211_X1 U5766 ( .C1(n5357), .C2(n6421), .A(n4722), .B(n4758), .ZN(n4735)
         );
  NOR3_X1 U5767 ( .A1(n4735), .A2(n4723), .A3(n6322), .ZN(n4724) );
  AOI211_X1 U5768 ( .C1(n4820), .C2(n5377), .A(n4725), .B(n4724), .ZN(n4729)
         );
  INV_X1 U5769 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6303) );
  INV_X1 U5770 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U5771 ( .A1(n5357), .A2(n4726), .ZN(n4816) );
  NAND2_X1 U5772 ( .A1(REIP_REG_17__SCAN_IN), .A2(n4802), .ZN(n5296) );
  NAND3_X1 U5773 ( .A1(n5169), .A2(REIP_REG_20__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n5168) );
  NOR2_X1 U5774 ( .A1(n5168), .A2(n5155), .ZN(n5145) );
  NAND2_X1 U5775 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5145), .ZN(n5128) );
  NAND2_X1 U5776 ( .A1(REIP_REG_27__SCAN_IN), .A2(n4776), .ZN(n4727) );
  NOR2_X1 U5777 ( .A1(n5128), .A2(n4727), .ZN(n4764) );
  NAND4_X1 U5778 ( .A1(n4753), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n6322), .ZN(n4728) );
  OAI211_X1 U5779 ( .C1(n4730), .C2(n5164), .A(n4729), .B(n4728), .ZN(U2796)
         );
  INV_X1 U5780 ( .A(n4823), .ZN(n4738) );
  INV_X1 U5781 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4824) );
  AOI22_X1 U5782 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5364), .B1(n5340), 
        .B2(n4732), .ZN(n4733) );
  OAI21_X1 U5783 ( .B1(n5361), .B2(n4824), .A(n4733), .ZN(n4737) );
  AOI21_X1 U5784 ( .B1(n4753), .B2(REIP_REG_29__SCAN_IN), .A(
        REIP_REG_30__SCAN_IN), .ZN(n4734) );
  NOR2_X1 U5785 ( .A1(n4735), .A2(n4734), .ZN(n4736) );
  AOI211_X1 U5786 ( .C1(n5377), .C2(n4738), .A(n4737), .B(n4736), .ZN(n4739)
         );
  OAI21_X1 U5787 ( .B1(n4897), .B2(n5164), .A(n4739), .ZN(U2797) );
  NAND2_X1 U5788 ( .A1(n4740), .A2(n4869), .ZN(n4742) );
  NAND2_X1 U5789 ( .A1(n4742), .A2(n4741), .ZN(n4743) );
  OR2_X1 U5790 ( .A1(n4681), .A2(n4743), .ZN(n4744) );
  NAND2_X1 U5791 ( .A1(n4745), .A2(n4744), .ZN(n4998) );
  NAND2_X1 U5792 ( .A1(n4758), .A2(REIP_REG_29__SCAN_IN), .ZN(n4751) );
  INV_X1 U5793 ( .A(n4746), .ZN(n4747) );
  OAI22_X1 U5794 ( .A1(n4748), .A2(n5374), .B1(n5386), .B2(n4747), .ZN(n4749)
         );
  AOI21_X1 U5795 ( .B1(n5368), .B2(EBX_REG_29__SCAN_IN), .A(n4749), .ZN(n4750)
         );
  OAI211_X1 U5796 ( .C1(n5367), .C2(n4998), .A(n4751), .B(n4750), .ZN(n4752)
         );
  AOI21_X1 U5797 ( .B1(n4753), .B2(n6421), .A(n4752), .ZN(n4754) );
  OAI21_X1 U5798 ( .B1(n4900), .B2(n5164), .A(n4754), .ZN(U2798) );
  AOI21_X1 U5799 ( .B1(n4755), .B2(n4136), .A(n4159), .ZN(n4917) );
  INV_X1 U5800 ( .A(n4917), .ZN(n4903) );
  INV_X1 U5801 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6447) );
  NOR2_X1 U5802 ( .A1(n4768), .A2(n4756), .ZN(n4757) );
  NAND2_X1 U5803 ( .A1(n4758), .A2(REIP_REG_28__SCAN_IN), .ZN(n4762) );
  OAI22_X1 U5804 ( .A1(n4759), .A2(n5374), .B1(n5386), .B2(n4915), .ZN(n4760)
         );
  AOI21_X1 U5805 ( .B1(n5368), .B2(EBX_REG_28__SCAN_IN), .A(n4760), .ZN(n4761)
         );
  OAI211_X1 U5806 ( .C1(n5367), .C2(n5008), .A(n4762), .B(n4761), .ZN(n4763)
         );
  AOI21_X1 U5807 ( .B1(n4764), .B2(n6447), .A(n4763), .ZN(n4765) );
  OAI21_X1 U5808 ( .B1(n4903), .B2(n5164), .A(n4765), .ZN(U2799) );
  INV_X1 U5809 ( .A(n5118), .ZN(n4775) );
  NOR2_X1 U5810 ( .A1(n4833), .A2(n4766), .ZN(n4767) );
  OR2_X1 U5811 ( .A1(n4768), .A2(n4767), .ZN(n5018) );
  AOI22_X1 U5812 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n5364), .B1(n4769), 
        .B2(n5340), .ZN(n4770) );
  OAI21_X1 U5813 ( .B1(n4771), .B2(n5361), .A(n4770), .ZN(n4772) );
  INV_X1 U5814 ( .A(n4772), .ZN(n4773) );
  OAI21_X1 U5815 ( .B1(n5367), .B2(n5018), .A(n4773), .ZN(n4774) );
  AOI21_X1 U5816 ( .B1(n4775), .B2(REIP_REG_27__SCAN_IN), .A(n4774), .ZN(n4779) );
  INV_X1 U5817 ( .A(n5128), .ZN(n4777) );
  NAND3_X1 U5818 ( .A1(n4777), .A2(n3930), .A3(n4776), .ZN(n4778) );
  OAI211_X1 U5819 ( .C1(n4906), .C2(n5164), .A(n4779), .B(n4778), .ZN(U2800)
         );
  BUF_X1 U5820 ( .A(n4781), .Z(n4782) );
  OAI21_X1 U5821 ( .B1(n4780), .B2(n4783), .A(n4782), .ZN(n4978) );
  OAI21_X1 U5822 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5296), .A(n5295), .ZN(n4794) );
  INV_X1 U5823 ( .A(n4981), .ZN(n4790) );
  MUX2_X1 U5824 ( .A(n4870), .B(n4786), .S(n4785), .Z(n4787) );
  INV_X1 U5825 ( .A(n4787), .ZN(n4882) );
  NAND2_X1 U5826 ( .A1(n4784), .A2(n4882), .ZN(n4884) );
  XNOR2_X1 U5827 ( .A(n4884), .B(n4788), .ZN(n5095) );
  AOI21_X1 U5828 ( .B1(n5377), .B2(n5095), .A(n5344), .ZN(n4789) );
  OAI21_X1 U5829 ( .B1(n4790), .B2(n5386), .A(n4789), .ZN(n4793) );
  AOI22_X1 U5830 ( .A1(EBX_REG_19__SCAN_IN), .A2(n5368), .B1(n5169), .B2(n6305), .ZN(n4791) );
  OAI21_X1 U5831 ( .B1(n4977), .B2(n5374), .A(n4791), .ZN(n4792) );
  AOI211_X1 U5832 ( .C1(REIP_REG_19__SCAN_IN), .C2(n4794), .A(n4793), .B(n4792), .ZN(n4795) );
  OAI21_X1 U5833 ( .B1(n4978), .B2(n5164), .A(n4795), .ZN(U2808) );
  XOR2_X1 U5834 ( .A(n4796), .B(n2971), .Z(n5402) );
  INV_X1 U5835 ( .A(n5402), .ZN(n4888) );
  INV_X1 U5836 ( .A(n4810), .ZN(n4798) );
  AOI21_X1 U5837 ( .B1(n4798), .B2(n4809), .A(n4797), .ZN(n4799) );
  NOR2_X1 U5838 ( .A1(n4799), .A2(n4784), .ZN(n5230) );
  INV_X1 U5839 ( .A(n5214), .ZN(n4801) );
  NAND2_X1 U5840 ( .A1(n5368), .A2(EBX_REG_17__SCAN_IN), .ZN(n4800) );
  OAI211_X1 U5841 ( .C1(n4801), .C2(n5386), .A(n4800), .B(n5359), .ZN(n4806)
         );
  NOR2_X1 U5842 ( .A1(REIP_REG_17__SCAN_IN), .A2(n4802), .ZN(n4804) );
  OAI22_X1 U5843 ( .A1(n4804), .A2(n5295), .B1(n4803), .B2(n5374), .ZN(n4805)
         );
  AOI211_X1 U5844 ( .C1(n5377), .C2(n5230), .A(n4806), .B(n4805), .ZN(n4807)
         );
  OAI21_X1 U5845 ( .B1(n4888), .B2(n5164), .A(n4807), .ZN(U2810) );
  AOI21_X1 U5846 ( .B1(n3007), .B2(n2976), .A(n2971), .ZN(n5407) );
  INV_X1 U5847 ( .A(n5407), .ZN(n4892) );
  XNOR2_X1 U5848 ( .A(n4810), .B(n4809), .ZN(n5109) );
  AOI22_X1 U5849 ( .A1(n5368), .A2(EBX_REG_16__SCAN_IN), .B1(n5340), .B2(n4986), .ZN(n4811) );
  INV_X1 U5850 ( .A(n4811), .ZN(n4818) );
  OAI21_X1 U5851 ( .B1(n6440), .B2(n4813), .A(n4812), .ZN(n4815) );
  AOI21_X1 U5852 ( .B1(n5364), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5344), 
        .ZN(n4814) );
  OAI221_X1 U5853 ( .B1(REIP_REG_16__SCAN_IN), .B2(n4816), .C1(n6300), .C2(
        n4815), .A(n4814), .ZN(n4817) );
  AOI211_X1 U5854 ( .C1(n5377), .C2(n5109), .A(n4818), .B(n4817), .ZN(n4819)
         );
  OAI21_X1 U5855 ( .B1(n4892), .B2(n5164), .A(n4819), .ZN(U2811) );
  INV_X1 U5856 ( .A(n4820), .ZN(n4822) );
  OAI22_X1 U5857 ( .A1(n4822), .A2(n5178), .B1(n5398), .B2(n4821), .ZN(U2828)
         );
  OAI222_X1 U5858 ( .A1(n4891), .A2(n4897), .B1(n4824), .B2(n5398), .C1(n4823), 
        .C2(n5178), .ZN(U2829) );
  OAI222_X1 U5859 ( .A1(n4891), .A2(n4900), .B1(n4825), .B2(n5398), .C1(n4998), 
        .C2(n5178), .ZN(U2830) );
  INV_X1 U5860 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4826) );
  OAI222_X1 U5861 ( .A1(n4891), .A2(n4903), .B1(n4826), .B2(n5398), .C1(n5008), 
        .C2(n5178), .ZN(U2831) );
  INV_X1 U5862 ( .A(n5018), .ZN(n4827) );
  AOI22_X1 U5863 ( .A1(n4827), .A2(n5393), .B1(EBX_REG_27__SCAN_IN), .B2(n4889), .ZN(n4828) );
  OAI21_X1 U5864 ( .B1(n4906), .B2(n4891), .A(n4828), .ZN(U2832) );
  NOR2_X1 U5865 ( .A1(n4829), .A2(n4830), .ZN(n4831) );
  INV_X1 U5866 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4835) );
  AND2_X1 U5867 ( .A1(n4842), .A2(n4832), .ZN(n4834) );
  OR2_X1 U5868 ( .A1(n4834), .A2(n4833), .ZN(n5117) );
  OAI222_X1 U5869 ( .A1(n4891), .A2(n4923), .B1(n4835), .B2(n5398), .C1(n5117), 
        .C2(n5178), .ZN(U2833) );
  AND2_X1 U5870 ( .A1(n4836), .A2(n4837), .ZN(n4838) );
  OR2_X1 U5871 ( .A1(n4838), .A2(n4829), .ZN(n5186) );
  INV_X1 U5872 ( .A(EBX_REG_25__SCAN_IN), .ZN(n4844) );
  INV_X1 U5873 ( .A(n4849), .ZN(n4841) );
  OAI21_X1 U5874 ( .B1(n4839), .B2(n4841), .A(n4840), .ZN(n4843) );
  NAND2_X1 U5875 ( .A1(n4843), .A2(n4842), .ZN(n5126) );
  OAI222_X1 U5876 ( .A1(n5186), .A2(n4891), .B1(n4844), .B2(n5398), .C1(n5178), 
        .C2(n5126), .ZN(U2834) );
  INV_X1 U5878 ( .A(n4836), .ZN(n4847) );
  AOI21_X1 U5879 ( .B1(n4848), .B2(n4853), .A(n4847), .ZN(n5190) );
  INV_X1 U5880 ( .A(n5190), .ZN(n4851) );
  XNOR2_X1 U5881 ( .A(n4839), .B(n4849), .ZN(n5134) );
  AOI22_X1 U5882 ( .A1(n5393), .A2(n5134), .B1(EBX_REG_24__SCAN_IN), .B2(n4889), .ZN(n4850) );
  OAI21_X1 U5883 ( .B1(n4851), .B2(n4891), .A(n4850), .ZN(U2835) );
  AOI21_X1 U5884 ( .B1(n4854), .B2(n4852), .A(n4846), .ZN(n4952) );
  INV_X1 U5885 ( .A(n4952), .ZN(n5143) );
  NAND2_X1 U5886 ( .A1(n5067), .A2(n4862), .ZN(n4857) );
  INV_X1 U5887 ( .A(n4855), .ZN(n4856) );
  NAND2_X1 U5888 ( .A1(n4857), .A2(n4856), .ZN(n4858) );
  AND2_X1 U5889 ( .A1(n4858), .A2(n4839), .ZN(n5141) );
  AOI22_X1 U5890 ( .A1(n5393), .A2(n5141), .B1(EBX_REG_23__SCAN_IN), .B2(n4889), .ZN(n4859) );
  OAI21_X1 U5891 ( .B1(n5143), .B2(n4891), .A(n4859), .ZN(U2836) );
  OAI21_X1 U5892 ( .B1(n4860), .B2(n4861), .A(n4852), .ZN(n4958) );
  XNOR2_X1 U5893 ( .A(n5067), .B(n4862), .ZN(n5159) );
  OAI22_X1 U5894 ( .A1(n5159), .A2(n5178), .B1(n4863), .B2(n5398), .ZN(n4864)
         );
  INV_X1 U5895 ( .A(n4864), .ZN(n4865) );
  OAI21_X1 U5896 ( .B1(n4958), .B2(n4891), .A(n4865), .ZN(U2837) );
  AOI21_X1 U5897 ( .B1(n4867), .B2(n4782), .A(n4866), .ZN(n5200) );
  INV_X1 U5898 ( .A(n5200), .ZN(n4874) );
  MUX2_X1 U5899 ( .A(n4870), .B(n4869), .S(n4868), .Z(n4872) );
  XNOR2_X1 U5900 ( .A(n4872), .B(n4871), .ZN(n5089) );
  INV_X1 U5901 ( .A(n5089), .ZN(n5170) );
  OAI222_X1 U5902 ( .A1(n4891), .A2(n4874), .B1(n4873), .B2(n5398), .C1(n5170), 
        .C2(n5178), .ZN(U2839) );
  INV_X1 U5903 ( .A(n5095), .ZN(n4876) );
  OAI22_X1 U5904 ( .A1(n5178), .A2(n4876), .B1(n4875), .B2(n5398), .ZN(n4877)
         );
  INV_X1 U5905 ( .A(n4877), .ZN(n4878) );
  OAI21_X1 U5906 ( .B1(n4978), .B2(n4891), .A(n4878), .ZN(U2840) );
  AND2_X1 U5907 ( .A1(n4880), .A2(n4879), .ZN(n4881) );
  OR2_X1 U5908 ( .A1(n4881), .A2(n4780), .ZN(n5207) );
  OR2_X1 U5909 ( .A1(n4784), .A2(n4882), .ZN(n4883) );
  INV_X1 U5910 ( .A(n5298), .ZN(n4885) );
  OAI222_X1 U5911 ( .A1(n5207), .A2(n4891), .B1(n4886), .B2(n5398), .C1(n5178), 
        .C2(n4885), .ZN(U2841) );
  AOI22_X1 U5912 ( .A1(n5393), .A2(n5230), .B1(EBX_REG_17__SCAN_IN), .B2(n4889), .ZN(n4887) );
  OAI21_X1 U5913 ( .B1(n4888), .B2(n4891), .A(n4887), .ZN(U2842) );
  AOI22_X1 U5914 ( .A1(n5393), .A2(n5109), .B1(EBX_REG_16__SCAN_IN), .B2(n4889), .ZN(n4890) );
  OAI21_X1 U5915 ( .B1(n4892), .B2(n4891), .A(n4890), .ZN(U2843) );
  AOI22_X1 U5916 ( .A1(n5405), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5408), .ZN(n4896) );
  NAND2_X1 U5917 ( .A1(n5409), .A2(DATAI_14_), .ZN(n4895) );
  OAI211_X1 U5918 ( .C1(n4897), .C2(n5182), .A(n4896), .B(n4895), .ZN(U2861)
         );
  AOI22_X1 U5919 ( .A1(n5405), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5408), .ZN(n4899) );
  NAND2_X1 U5920 ( .A1(n5409), .A2(DATAI_13_), .ZN(n4898) );
  OAI211_X1 U5921 ( .C1(n4900), .C2(n5182), .A(n4899), .B(n4898), .ZN(U2862)
         );
  AOI22_X1 U5922 ( .A1(n5405), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5408), .ZN(n4902) );
  NAND2_X1 U5923 ( .A1(n5409), .A2(DATAI_12_), .ZN(n4901) );
  OAI211_X1 U5924 ( .C1(n4903), .C2(n5182), .A(n4902), .B(n4901), .ZN(U2863)
         );
  AOI22_X1 U5925 ( .A1(n5405), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5408), .ZN(n4905) );
  NAND2_X1 U5926 ( .A1(n5409), .A2(DATAI_11_), .ZN(n4904) );
  OAI211_X1 U5927 ( .C1(n4906), .C2(n5182), .A(n4905), .B(n4904), .ZN(U2864)
         );
  AOI22_X1 U5928 ( .A1(n5409), .A2(DATAI_7_), .B1(n5408), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n4908) );
  NAND2_X1 U5929 ( .A1(n5405), .A2(DATAI_23_), .ZN(n4907) );
  OAI211_X1 U5930 ( .C1(n5143), .C2(n5182), .A(n4908), .B(n4907), .ZN(U2868)
         );
  AOI22_X1 U5931 ( .A1(n5405), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5408), .ZN(n4910) );
  NAND2_X1 U5932 ( .A1(n5409), .A2(DATAI_3_), .ZN(n4909) );
  OAI211_X1 U5933 ( .C1(n4978), .C2(n5182), .A(n4910), .B(n4909), .ZN(U2872)
         );
  NAND3_X1 U5934 ( .A1(n4922), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5203), .ZN(n4912) );
  INV_X1 U5935 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5026) );
  XNOR2_X1 U5936 ( .A(n4913), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5016)
         );
  NOR2_X1 U5937 ( .A1(n5612), .A2(n6447), .ZN(n5010) );
  AOI21_X1 U5938 ( .B1(n5536), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5010), 
        .ZN(n4914) );
  OAI21_X1 U5939 ( .B1(n4915), .B2(n5546), .A(n4914), .ZN(n4916) );
  AOI21_X1 U5940 ( .B1(n4917), .B2(n5702), .A(n4916), .ZN(n4918) );
  OAI21_X1 U5941 ( .B1(n5555), .B2(n5016), .A(n4918), .ZN(U2958) );
  NAND2_X1 U5942 ( .A1(n4920), .A2(n4919), .ZN(n4921) );
  XNOR2_X1 U5943 ( .A(n4922), .B(n4921), .ZN(n5033) );
  NOR2_X1 U5944 ( .A1(n5546), .A2(n5123), .ZN(n4927) );
  INV_X1 U5945 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4925) );
  INV_X1 U5946 ( .A(REIP_REG_26__SCAN_IN), .ZN(n4924) );
  OR2_X1 U5947 ( .A1(n5612), .A2(n4924), .ZN(n5028) );
  OAI21_X1 U5948 ( .B1(n5550), .B2(n4925), .A(n5028), .ZN(n4926) );
  AOI211_X1 U5949 ( .C1(n5183), .C2(n5702), .A(n4927), .B(n4926), .ZN(n4928)
         );
  OAI21_X1 U5950 ( .B1(n5033), .B2(n5555), .A(n4928), .ZN(U2960) );
  NAND2_X1 U5951 ( .A1(n5630), .A2(REIP_REG_25__SCAN_IN), .ZN(n5035) );
  OAI21_X1 U5952 ( .B1(n5550), .B2(n4929), .A(n5035), .ZN(n4930) );
  AOI21_X1 U5953 ( .B1(n5517), .B2(n5125), .A(n4930), .ZN(n4933) );
  OAI21_X1 U5954 ( .B1(n3440), .B2(n4931), .A(n3939), .ZN(n5034) );
  NAND2_X1 U5955 ( .A1(n5034), .A2(n5541), .ZN(n4932) );
  OAI211_X1 U5956 ( .C1(n5186), .C2(n5692), .A(n4933), .B(n4932), .ZN(U2961)
         );
  OAI21_X1 U5957 ( .B1(n4934), .B2(n6476), .A(n5203), .ZN(n4936) );
  XNOR2_X1 U5958 ( .A(n5203), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4970)
         );
  NOR2_X1 U5959 ( .A1(n5203), .A2(n5086), .ZN(n4937) );
  XNOR2_X1 U5960 ( .A(n5203), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4966)
         );
  NOR2_X1 U5961 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4955)
         );
  NAND2_X1 U5962 ( .A1(n4938), .A2(n4955), .ZN(n4946) );
  OAI21_X1 U5963 ( .B1(n5204), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n4964), 
        .ZN(n4957) );
  NAND3_X1 U5964 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4939) );
  XNOR2_X1 U5965 ( .A(n4940), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5049)
         );
  INV_X1 U5966 ( .A(n5133), .ZN(n4942) );
  NAND2_X1 U5967 ( .A1(n5630), .A2(REIP_REG_24__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U5968 ( .A1(n5536), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4941)
         );
  OAI211_X1 U5969 ( .C1(n5546), .C2(n4942), .A(n5041), .B(n4941), .ZN(n4943)
         );
  AOI21_X1 U5970 ( .B1(n5190), .B2(n5702), .A(n4943), .ZN(n4944) );
  OAI21_X1 U5971 ( .B1(n5049), .B2(n5555), .A(n4944), .ZN(U2962) );
  NAND2_X1 U5972 ( .A1(n5203), .A2(n4945), .ZN(n4947) );
  OAI21_X1 U5973 ( .B1(n4934), .B2(n4947), .A(n4946), .ZN(n4948) );
  XNOR2_X1 U5974 ( .A(n4948), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5056)
         );
  INV_X1 U5975 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4949) );
  NOR2_X1 U5976 ( .A1(n5612), .A2(n4949), .ZN(n5052) );
  NOR2_X1 U5977 ( .A1(n5550), .A2(n4950), .ZN(n4951) );
  AOI211_X1 U5978 ( .C1(n5517), .C2(n5140), .A(n5052), .B(n4951), .ZN(n4954)
         );
  NAND2_X1 U5979 ( .A1(n4952), .A2(n5702), .ZN(n4953) );
  OAI211_X1 U5980 ( .C1(n5056), .C2(n5555), .A(n4954), .B(n4953), .ZN(U2963)
         );
  AOI21_X1 U5981 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5203), .A(n4955), 
        .ZN(n4956) );
  XNOR2_X1 U5982 ( .A(n4957), .B(n4956), .ZN(n5065) );
  INV_X1 U5983 ( .A(n4958), .ZN(n5193) );
  NAND2_X1 U5984 ( .A1(n5630), .A2(REIP_REG_22__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U5985 ( .A1(n5536), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4959)
         );
  OAI211_X1 U5986 ( .C1(n5546), .C2(n5150), .A(n5058), .B(n4959), .ZN(n4960)
         );
  AOI21_X1 U5987 ( .B1(n5193), .B2(n5702), .A(n4960), .ZN(n4961) );
  OAI21_X1 U5988 ( .B1(n5065), .B2(n5555), .A(n4961), .ZN(U2964) );
  XNOR2_X1 U5989 ( .A(n4963), .B(n4962), .ZN(n5196) );
  OAI21_X1 U5990 ( .B1(n4966), .B2(n4965), .A(n4964), .ZN(n5066) );
  NAND2_X1 U5991 ( .A1(n5066), .A2(n5541), .ZN(n4969) );
  INV_X1 U5992 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U5993 ( .A1(n5630), .A2(REIP_REG_21__SCAN_IN), .ZN(n5071) );
  OAI21_X1 U5994 ( .B1(n5550), .B2(n6510), .A(n5071), .ZN(n4967) );
  AOI21_X1 U5995 ( .B1(n5517), .B2(n5163), .A(n4967), .ZN(n4968) );
  OAI211_X1 U5996 ( .C1(n5692), .C2(n5196), .A(n4969), .B(n4968), .ZN(U2965)
         );
  XNOR2_X1 U5997 ( .A(n4971), .B(n4970), .ZN(n5094) );
  NOR2_X1 U5998 ( .A1(n5612), .A2(n6307), .ZN(n5088) );
  AOI21_X1 U5999 ( .B1(n5536), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5088), 
        .ZN(n4972) );
  OAI21_X1 U6000 ( .B1(n5176), .B2(n5546), .A(n4972), .ZN(n4973) );
  AOI21_X1 U6001 ( .B1(n5200), .B2(n5702), .A(n4973), .ZN(n4974) );
  OAI21_X1 U6002 ( .B1(n5555), .B2(n5094), .A(n4974), .ZN(U2966) );
  OAI21_X1 U6003 ( .B1(n4975), .B2(n6476), .A(n4935), .ZN(n4976) );
  XNOR2_X1 U6004 ( .A(n4976), .B(n5203), .ZN(n5102) );
  NAND2_X1 U6005 ( .A1(n5630), .A2(REIP_REG_19__SCAN_IN), .ZN(n5097) );
  OAI21_X1 U6006 ( .B1(n5550), .B2(n4977), .A(n5097), .ZN(n4980) );
  NOR2_X1 U6007 ( .A1(n4978), .A2(n5692), .ZN(n4979) );
  AOI211_X1 U6008 ( .C1(n5517), .C2(n4981), .A(n4980), .B(n4979), .ZN(n4982)
         );
  OAI21_X1 U6009 ( .B1(n5555), .B2(n5102), .A(n4982), .ZN(U2967) );
  XNOR2_X1 U6010 ( .A(n5203), .B(n6497), .ZN(n4984) );
  XNOR2_X1 U6011 ( .A(n4983), .B(n4984), .ZN(n5112) );
  NOR2_X1 U6012 ( .A1(n5612), .A2(n6300), .ZN(n5108) );
  AND2_X1 U6013 ( .A1(n5536), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4985)
         );
  AOI211_X1 U6014 ( .C1(n5517), .C2(n4986), .A(n5108), .B(n4985), .ZN(n4988)
         );
  NAND2_X1 U6015 ( .A1(n5407), .A2(n5702), .ZN(n4987) );
  OAI211_X1 U6016 ( .C1(n5112), .C2(n5555), .A(n4988), .B(n4987), .ZN(U2970)
         );
  XNOR2_X1 U6017 ( .A(n5203), .B(n5240), .ZN(n4990) );
  XNOR2_X1 U6018 ( .A(n4989), .B(n4990), .ZN(n5237) );
  NAND2_X1 U6019 ( .A1(n5237), .A2(n5541), .ZN(n4994) );
  OAI22_X1 U6020 ( .A1(n5550), .A2(n3699), .B1(n5612), .B2(n6440), .ZN(n4991)
         );
  AOI21_X1 U6021 ( .B1(n5517), .B2(n4992), .A(n4991), .ZN(n4993) );
  OAI211_X1 U6022 ( .C1(n5692), .C2(n4995), .A(n4994), .B(n4993), .ZN(U2971)
         );
  INV_X1 U6023 ( .A(n4997), .ZN(n5001) );
  NOR2_X1 U6024 ( .A1(n4998), .A2(n5585), .ZN(n4999) );
  AOI211_X1 U6025 ( .C1(n5001), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5000), .B(n4999), .ZN(n5005) );
  INV_X1 U6026 ( .A(n5024), .ZN(n5013) );
  NAND3_X1 U6027 ( .A1(n5013), .A2(n5003), .A3(n5002), .ZN(n5004) );
  OAI211_X1 U6028 ( .C1(n5006), .C2(n5654), .A(n5005), .B(n5004), .ZN(U2989)
         );
  INV_X1 U6029 ( .A(n5037), .ZN(n5043) );
  OAI21_X1 U6030 ( .B1(n5007), .B2(n5572), .A(n5043), .ZN(n5021) );
  NOR2_X1 U6031 ( .A1(n5008), .A2(n5585), .ZN(n5009) );
  AOI211_X1 U6032 ( .C1(n5021), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5010), .B(n5009), .ZN(n5015) );
  NAND3_X1 U6033 ( .A1(n5013), .A2(n5012), .A3(n5011), .ZN(n5014) );
  OAI211_X1 U6034 ( .C1(n5016), .C2(n5654), .A(n5015), .B(n5014), .ZN(U2990)
         );
  NAND2_X1 U6035 ( .A1(n5017), .A2(n5636), .ZN(n5023) );
  NOR2_X1 U6036 ( .A1(n5018), .A2(n5585), .ZN(n5019) );
  AOI211_X1 U6037 ( .C1(n5021), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5020), .B(n5019), .ZN(n5022) );
  OAI211_X1 U6038 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5024), .A(n5023), .B(n5022), .ZN(U2991) );
  NAND2_X1 U6039 ( .A1(n5025), .A2(n3438), .ZN(n5038) );
  AOI21_X1 U6040 ( .B1(n5038), .B2(n5043), .A(n5026), .ZN(n5031) );
  NOR4_X1 U6041 ( .A1(n5090), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5027), 
        .A4(n3438), .ZN(n5030) );
  OAI21_X1 U6042 ( .B1(n5117), .B2(n5585), .A(n5028), .ZN(n5029) );
  NOR3_X1 U6043 ( .A1(n5031), .A2(n5030), .A3(n5029), .ZN(n5032) );
  OAI21_X1 U6044 ( .B1(n5033), .B2(n5654), .A(n5032), .ZN(U2992) );
  INV_X1 U6045 ( .A(n5034), .ZN(n5040) );
  OAI21_X1 U6046 ( .B1(n5126), .B2(n5585), .A(n5035), .ZN(n5036) );
  AOI21_X1 U6047 ( .B1(n5037), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5036), 
        .ZN(n5039) );
  OAI211_X1 U6048 ( .C1(n5040), .C2(n5654), .A(n5039), .B(n5038), .ZN(U2993)
         );
  INV_X1 U6049 ( .A(n5041), .ZN(n5047) );
  NOR2_X1 U6050 ( .A1(n5090), .A2(n5091), .ZN(n5059) );
  INV_X1 U6051 ( .A(n5042), .ZN(n5060) );
  NAND3_X1 U6052 ( .A1(n5059), .A2(n5060), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5045) );
  AOI21_X1 U6053 ( .B1(n5045), .B2(n5044), .A(n5043), .ZN(n5046) );
  AOI211_X1 U6054 ( .C1(n5649), .C2(n5134), .A(n5047), .B(n5046), .ZN(n5048)
         );
  OAI21_X1 U6055 ( .B1(n5049), .B2(n5654), .A(n5048), .ZN(U2994) );
  NOR2_X1 U6056 ( .A1(n5050), .A2(n5053), .ZN(n5051) );
  AOI211_X1 U6057 ( .C1(n5649), .C2(n5141), .A(n5052), .B(n5051), .ZN(n5055)
         );
  NAND3_X1 U6058 ( .A1(n5059), .A2(n5060), .A3(n5053), .ZN(n5054) );
  OAI211_X1 U6059 ( .C1(n5056), .C2(n5654), .A(n5055), .B(n5054), .ZN(U2995)
         );
  INV_X1 U6060 ( .A(n5057), .ZN(n5073) );
  OAI21_X1 U6061 ( .B1(n5585), .B2(n5159), .A(n5058), .ZN(n5063) );
  INV_X1 U6062 ( .A(n5059), .ZN(n5076) );
  NOR3_X1 U6063 ( .A1(n5076), .A2(n5061), .A3(n5060), .ZN(n5062) );
  AOI211_X1 U6064 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5073), .A(n5063), .B(n5062), .ZN(n5064) );
  OAI21_X1 U6065 ( .B1(n5065), .B2(n5654), .A(n5064), .ZN(U2996) );
  NAND2_X1 U6066 ( .A1(n5066), .A2(n5636), .ZN(n5075) );
  INV_X1 U6067 ( .A(n5067), .ZN(n5070) );
  NAND2_X1 U6068 ( .A1(n2974), .A2(n5068), .ZN(n5069) );
  NAND2_X1 U6069 ( .A1(n5070), .A2(n5069), .ZN(n5177) );
  OAI21_X1 U6070 ( .B1(n5585), .B2(n5177), .A(n5071), .ZN(n5072) );
  AOI21_X1 U6071 ( .B1(n5073), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5072), 
        .ZN(n5074) );
  OAI211_X1 U6072 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5076), .A(n5075), .B(n5074), .ZN(U2997) );
  OAI22_X1 U6073 ( .A1(n5079), .A2(n5078), .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5077), .ZN(n5085) );
  INV_X1 U6074 ( .A(n5080), .ZN(n5081) );
  NAND2_X1 U6075 ( .A1(n5569), .A2(n5081), .ZN(n5084) );
  OAI21_X1 U6076 ( .B1(n5228), .B2(n5082), .A(n5571), .ZN(n5083) );
  NAND2_X1 U6077 ( .A1(n5084), .A2(n5083), .ZN(n5231) );
  NOR2_X1 U6078 ( .A1(n5085), .A2(n5231), .ZN(n5098) );
  NOR2_X1 U6079 ( .A1(n5098), .A2(n5086), .ZN(n5087) );
  AOI211_X1 U6080 ( .C1(n5649), .C2(n5089), .A(n5088), .B(n5087), .ZN(n5093)
         );
  INV_X1 U6081 ( .A(n5090), .ZN(n5100) );
  OAI211_X1 U6082 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5100), .B(n5091), .ZN(n5092) );
  OAI211_X1 U6083 ( .C1(n5094), .C2(n5654), .A(n5093), .B(n5092), .ZN(U2998)
         );
  NAND2_X1 U6084 ( .A1(n5649), .A2(n5095), .ZN(n5096) );
  OAI211_X1 U6085 ( .C1(n5098), .C2(n6476), .A(n5097), .B(n5096), .ZN(n5099)
         );
  AOI21_X1 U6086 ( .B1(n5100), .B2(n6476), .A(n5099), .ZN(n5101) );
  OAI21_X1 U6087 ( .B1(n5102), .B2(n5654), .A(n5101), .ZN(U2999) );
  AOI21_X1 U6088 ( .B1(n5103), .B2(n5104), .A(n5558), .ZN(n5241) );
  NOR2_X1 U6089 ( .A1(n5264), .A2(n5104), .ZN(n5235) );
  NAND2_X1 U6090 ( .A1(n5235), .A2(n5105), .ZN(n5106) );
  OAI21_X1 U6091 ( .B1(n5241), .B2(n6497), .A(n5106), .ZN(n5107) );
  OAI21_X1 U6092 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5107), .ZN(n5111) );
  AOI21_X1 U6093 ( .B1(n5649), .B2(n5109), .A(n5108), .ZN(n5110) );
  OAI211_X1 U6094 ( .C1(n5112), .C2(n5654), .A(n5111), .B(n5110), .ZN(U3002)
         );
  AND2_X1 U6095 ( .A1(n5423), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6096 ( .A(n5113), .ZN(n5431) );
  AOI21_X1 U6097 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5114), .A(n5431), .ZN(
        n5116) );
  NAND2_X1 U6098 ( .A1(n5116), .A2(n5115), .ZN(U2788) );
  AOI22_X1 U6099 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5368), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5364), .ZN(n5122) );
  INV_X1 U6100 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6430) );
  NOR2_X1 U6101 ( .A1(n6430), .A2(n5128), .ZN(n5124) );
  AOI21_X1 U6102 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5124), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5119) );
  OAI22_X1 U6103 ( .A1(n5119), .A2(n5118), .B1(n5117), .B2(n5367), .ZN(n5120)
         );
  AOI21_X1 U6104 ( .B1(n5183), .B2(n5351), .A(n5120), .ZN(n5121) );
  OAI211_X1 U6105 ( .C1(n5123), .C2(n5386), .A(n5122), .B(n5121), .ZN(U2801)
         );
  AOI22_X1 U6106 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5368), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5364), .ZN(n5132) );
  INV_X1 U6107 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6314) );
  AOI22_X1 U6108 ( .A1(n5125), .A2(n5340), .B1(n5124), .B2(n6314), .ZN(n5131)
         );
  OAI22_X1 U6109 ( .A1(n5186), .A2(n5164), .B1(n5367), .B2(n5126), .ZN(n5127)
         );
  INV_X1 U6110 ( .A(n5127), .ZN(n5130) );
  NOR2_X1 U6111 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5128), .ZN(n5135) );
  OAI21_X1 U6112 ( .B1(n5135), .B2(n5146), .A(REIP_REG_25__SCAN_IN), .ZN(n5129) );
  NAND4_X1 U6113 ( .A1(n5132), .A2(n5131), .A3(n5130), .A4(n5129), .ZN(U2802)
         );
  AOI22_X1 U6114 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5368), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5364), .ZN(n5139) );
  AOI22_X1 U6115 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5146), .B1(n5133), .B2(
        n5340), .ZN(n5138) );
  AOI22_X1 U6116 ( .A1(n5190), .A2(n5351), .B1(n5377), .B2(n5134), .ZN(n5137)
         );
  INV_X1 U6117 ( .A(n5135), .ZN(n5136) );
  NAND4_X1 U6118 ( .A1(n5139), .A2(n5138), .A3(n5137), .A4(n5136), .ZN(U2803)
         );
  AOI22_X1 U6119 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n5364), .B1(n5140), 
        .B2(n5340), .ZN(n5148) );
  INV_X1 U6120 ( .A(n5141), .ZN(n5142) );
  OAI22_X1 U6121 ( .A1(n5143), .A2(n5164), .B1(n5142), .B2(n5367), .ZN(n5144)
         );
  AOI221_X1 U6122 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5146), .C1(n5145), .C2(
        n5146), .A(n5144), .ZN(n5147) );
  OAI211_X1 U6123 ( .C1(n5149), .C2(n5361), .A(n5148), .B(n5147), .ZN(U2804)
         );
  INV_X1 U6124 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6310) );
  INV_X1 U6125 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5151) );
  OAI22_X1 U6126 ( .A1(n5151), .A2(n5374), .B1(n5386), .B2(n5150), .ZN(n5152)
         );
  AOI21_X1 U6127 ( .B1(n5368), .B2(EBX_REG_22__SCAN_IN), .A(n5152), .ZN(n5153)
         );
  OAI21_X1 U6128 ( .B1(n5171), .B2(n6310), .A(n5153), .ZN(n5154) );
  AOI21_X1 U6129 ( .B1(n5193), .B2(n5351), .A(n5154), .ZN(n5158) );
  INV_X1 U6130 ( .A(n5168), .ZN(n5156) );
  OAI211_X1 U6131 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5156), .B(n5155), .ZN(n5157) );
  OAI211_X1 U6132 ( .C1(n5367), .C2(n5159), .A(n5158), .B(n5157), .ZN(U2805)
         );
  INV_X1 U6133 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5181) );
  AOI22_X1 U6134 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n5364), .B1(
        REIP_REG_21__SCAN_IN), .B2(n5160), .ZN(n5161) );
  OAI21_X1 U6135 ( .B1(n5181), .B2(n5361), .A(n5161), .ZN(n5162) );
  AOI21_X1 U6136 ( .B1(n5163), .B2(n5340), .A(n5162), .ZN(n5167) );
  OAI22_X1 U6137 ( .A1(n5196), .A2(n5164), .B1(n5367), .B2(n5177), .ZN(n5165)
         );
  INV_X1 U6138 ( .A(n5165), .ZN(n5166) );
  OAI211_X1 U6139 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5168), .A(n5167), .B(n5166), .ZN(U2806) );
  AOI22_X1 U6140 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5368), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5364), .ZN(n5175) );
  AOI21_X1 U6141 ( .B1(n5169), .B2(REIP_REG_19__SCAN_IN), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5172) );
  OAI22_X1 U6142 ( .A1(n5172), .A2(n5171), .B1(n5367), .B2(n5170), .ZN(n5173)
         );
  AOI21_X1 U6143 ( .B1(n5200), .B2(n5351), .A(n5173), .ZN(n5174) );
  OAI211_X1 U6144 ( .C1(n5176), .C2(n5386), .A(n5175), .B(n5174), .ZN(U2807)
         );
  OAI22_X1 U6145 ( .A1(n5196), .A2(n4891), .B1(n5178), .B2(n5177), .ZN(n5179)
         );
  INV_X1 U6146 ( .A(n5179), .ZN(n5180) );
  OAI21_X1 U6147 ( .B1(n5398), .B2(n5181), .A(n5180), .ZN(U2838) );
  AOI22_X1 U6148 ( .A1(n5183), .A2(n5406), .B1(n5405), .B2(DATAI_26_), .ZN(
        n5185) );
  AOI22_X1 U6149 ( .A1(n5409), .A2(DATAI_10_), .B1(n5408), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6150 ( .A1(n5185), .A2(n5184), .ZN(U2865) );
  INV_X1 U6151 ( .A(n5186), .ZN(n5187) );
  AOI22_X1 U6152 ( .A1(n5187), .A2(n5406), .B1(n5405), .B2(DATAI_25_), .ZN(
        n5189) );
  AOI22_X1 U6153 ( .A1(n5409), .A2(DATAI_9_), .B1(n5408), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6154 ( .A1(n5189), .A2(n5188), .ZN(U2866) );
  AOI22_X1 U6155 ( .A1(n5190), .A2(n5406), .B1(n5405), .B2(DATAI_24_), .ZN(
        n5192) );
  AOI22_X1 U6156 ( .A1(n5409), .A2(DATAI_8_), .B1(n5408), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6157 ( .A1(n5192), .A2(n5191), .ZN(U2867) );
  AOI22_X1 U6158 ( .A1(n5193), .A2(n5406), .B1(n5405), .B2(DATAI_22_), .ZN(
        n5195) );
  AOI22_X1 U6159 ( .A1(n5409), .A2(DATAI_6_), .B1(n5408), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6160 ( .A1(n5195), .A2(n5194), .ZN(U2869) );
  INV_X1 U6161 ( .A(n5196), .ZN(n5197) );
  AOI22_X1 U6162 ( .A1(n5197), .A2(n5406), .B1(n5405), .B2(DATAI_21_), .ZN(
        n5199) );
  AOI22_X1 U6163 ( .A1(n5409), .A2(DATAI_5_), .B1(n5408), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6164 ( .A1(n5199), .A2(n5198), .ZN(U2870) );
  AOI22_X1 U6165 ( .A1(n5200), .A2(n5406), .B1(n5405), .B2(DATAI_20_), .ZN(
        n5202) );
  AOI22_X1 U6166 ( .A1(n5409), .A2(DATAI_4_), .B1(n5408), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6167 ( .A1(n5202), .A2(n5201), .ZN(U2871) );
  AOI22_X1 U6168 ( .A1(n5630), .A2(REIP_REG_18__SCAN_IN), .B1(n5536), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5209) );
  NAND3_X1 U6169 ( .A1(n4983), .A2(n5204), .A3(n6497), .ZN(n5210) );
  NOR3_X1 U6170 ( .A1(n4983), .A2(n5204), .A3(n6497), .ZN(n5212) );
  NAND2_X1 U6171 ( .A1(n5212), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5205) );
  OAI21_X1 U6172 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5210), .A(n5205), 
        .ZN(n5206) );
  XNOR2_X1 U6173 ( .A(n5206), .B(n5223), .ZN(n5221) );
  AOI22_X1 U6174 ( .A1(n5221), .A2(n5541), .B1(n5702), .B2(n5399), .ZN(n5208)
         );
  OAI211_X1 U6175 ( .C1(n5546), .C2(n5301), .A(n5209), .B(n5208), .ZN(U2968)
         );
  INV_X1 U6176 ( .A(n5210), .ZN(n5211) );
  NOR2_X1 U6177 ( .A1(n5212), .A2(n5211), .ZN(n5213) );
  XNOR2_X1 U6178 ( .A(n5213), .B(n5228), .ZN(n5234) );
  AOI22_X1 U6179 ( .A1(n5630), .A2(REIP_REG_17__SCAN_IN), .B1(n5536), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5216) );
  AOI22_X1 U6180 ( .A1(n5402), .A2(n5702), .B1(n5517), .B2(n5214), .ZN(n5215)
         );
  OAI211_X1 U6181 ( .C1(n5234), .C2(n5555), .A(n5216), .B(n5215), .ZN(U2969)
         );
  AOI22_X1 U6182 ( .A1(n5630), .A2(REIP_REG_13__SCAN_IN), .B1(n5536), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5220) );
  XNOR2_X1 U6183 ( .A(n5217), .B(n5218), .ZN(n5260) );
  AOI22_X1 U6184 ( .A1(n5260), .A2(n5541), .B1(n5702), .B2(n5388), .ZN(n5219)
         );
  OAI211_X1 U6185 ( .C1(n5546), .C2(n5320), .A(n5220), .B(n5219), .ZN(U2973)
         );
  AOI22_X1 U6186 ( .A1(n5221), .A2(n5636), .B1(n5649), .B2(n5298), .ZN(n5227)
         );
  NAND2_X1 U6187 ( .A1(n5630), .A2(REIP_REG_18__SCAN_IN), .ZN(n5226) );
  OAI221_X1 U6188 ( .B1(n5231), .B2(n5222), .C1(n5231), .C2(n5228), .A(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5225) );
  NAND3_X1 U6189 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5229), .A3(n5223), .ZN(n5224) );
  NAND4_X1 U6190 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(U3000)
         );
  AOI22_X1 U6191 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5630), .B1(n5229), .B2(
        n5228), .ZN(n5233) );
  AOI22_X1 U6192 ( .A1(n5231), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n5649), .B2(n5230), .ZN(n5232) );
  OAI211_X1 U6193 ( .C1(n5234), .C2(n5654), .A(n5233), .B(n5232), .ZN(U3001)
         );
  AOI22_X1 U6194 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5630), .B1(n5235), .B2(
        n5240), .ZN(n5239) );
  AOI22_X1 U6195 ( .A1(n5237), .A2(n5636), .B1(n5649), .B2(n5236), .ZN(n5238)
         );
  OAI211_X1 U6196 ( .C1(n5241), .C2(n5240), .A(n5239), .B(n5238), .ZN(U3003)
         );
  INV_X1 U6197 ( .A(n5264), .ZN(n5557) );
  NAND2_X1 U6198 ( .A1(n5247), .A2(n5557), .ZN(n5253) );
  AOI21_X1 U6199 ( .B1(n5243), .B2(n5242), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5250) );
  INV_X1 U6200 ( .A(n5651), .ZN(n5246) );
  AOI21_X1 U6201 ( .B1(n5244), .B2(n5254), .A(n5558), .ZN(n5245) );
  OAI21_X1 U6202 ( .B1(n5247), .B2(n5246), .A(n5245), .ZN(n5259) );
  OAI22_X1 U6203 ( .A1(n5248), .A2(n5654), .B1(n5585), .B2(n5303), .ZN(n5249)
         );
  AOI221_X1 U6204 ( .B1(n5250), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .C1(
        n5259), .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5249), .ZN(n5252) );
  NAND2_X1 U6205 ( .A1(n5630), .A2(REIP_REG_14__SCAN_IN), .ZN(n5251) );
  OAI211_X1 U6206 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n5253), .A(n5252), .B(n5251), .ZN(U3004) );
  OR2_X1 U6207 ( .A1(n5254), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5263)
         );
  AND2_X1 U6208 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  NOR2_X1 U6209 ( .A1(n5258), .A2(n5257), .ZN(n5387) );
  AOI22_X1 U6210 ( .A1(n5649), .A2(n5387), .B1(n5630), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5262) );
  AOI22_X1 U6211 ( .A1(n5260), .A2(n5636), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5259), .ZN(n5261) );
  OAI211_X1 U6212 ( .C1(n5264), .C2(n5263), .A(n5262), .B(n5261), .ZN(U3005)
         );
  INV_X1 U6213 ( .A(n5265), .ZN(n5267) );
  NAND4_X1 U6214 ( .A1(n5267), .A2(n5266), .A3(n6252), .A4(n5354), .ZN(n5268)
         );
  OAI21_X1 U6215 ( .B1(n6340), .B2(n4299), .A(n5268), .ZN(U3455) );
  INV_X1 U6216 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6459) );
  AOI21_X1 U6217 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6459), .A(n6523), .ZN(n5276) );
  INV_X1 U6218 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5269) );
  AOI21_X1 U6219 ( .B1(n5276), .B2(n5269), .A(n6376), .ZN(U2789) );
  NAND2_X1 U6220 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5270), .ZN(n5274) );
  INV_X1 U6221 ( .A(n5271), .ZN(n5272) );
  OAI21_X1 U6222 ( .B1(n5272), .B2(n6236), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5273) );
  OAI21_X1 U6223 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5274), .A(n5273), .ZN(
        U2790) );
  INV_X2 U6224 ( .A(n6376), .ZN(n6543) );
  NOR2_X1 U6225 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5277) );
  OAI21_X1 U6226 ( .B1(n5277), .B2(D_C_N_REG_SCAN_IN), .A(n6543), .ZN(n5275)
         );
  OAI21_X1 U6227 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6543), .A(n5275), .ZN(
        U2791) );
  NOR2_X1 U6228 ( .A1(n6376), .A2(n5276), .ZN(n6328) );
  OAI21_X1 U6229 ( .B1(n5277), .B2(BS16_N), .A(n6328), .ZN(n6326) );
  OAI21_X1 U6230 ( .B1(n6328), .B2(n6363), .A(n6326), .ZN(U2792) );
  OAI21_X1 U6231 ( .B1(n5278), .B2(n6229), .A(n5555), .ZN(U2793) );
  NOR4_X1 U6232 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5282) );
  NOR4_X1 U6233 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5281) );
  NOR4_X1 U6234 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5280) );
  NOR4_X1 U6235 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5279) );
  NAND4_X1 U6236 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n5288)
         );
  NOR4_X1 U6237 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n5286) );
  AOI211_X1 U6238 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_10__SCAN_IN), .B(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n5285) );
  NOR4_X1 U6239 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5284) );
  NOR4_X1 U6240 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5283) );
  NAND4_X1 U6241 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n5287)
         );
  NOR2_X1 U6242 ( .A1(n5288), .A2(n5287), .ZN(n6357) );
  INV_X1 U6243 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5290) );
  NOR3_X1 U6244 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5291) );
  OAI21_X1 U6245 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5291), .A(n6357), .ZN(n5289)
         );
  OAI21_X1 U6246 ( .B1(n6357), .B2(n5290), .A(n5289), .ZN(U2794) );
  INV_X1 U6247 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6327) );
  AOI21_X1 U6248 ( .B1(n6353), .B2(n6327), .A(n5291), .ZN(n5293) );
  INV_X1 U6249 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5292) );
  INV_X1 U6250 ( .A(n6357), .ZN(n6360) );
  AOI22_X1 U6251 ( .A1(n6357), .A2(n5293), .B1(n5292), .B2(n6360), .ZN(U2795)
         );
  AOI21_X1 U6252 ( .B1(n5364), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5344), 
        .ZN(n5294) );
  OAI221_X1 U6253 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5296), .C1(n6303), .C2(
        n5295), .A(n5294), .ZN(n5297) );
  AOI21_X1 U6254 ( .B1(EBX_REG_18__SCAN_IN), .B2(n5368), .A(n5297), .ZN(n5300)
         );
  AOI22_X1 U6255 ( .A1(n5399), .A2(n5351), .B1(n5377), .B2(n5298), .ZN(n5299)
         );
  OAI211_X1 U6256 ( .C1(n5301), .C2(n5386), .A(n5300), .B(n5299), .ZN(U2809)
         );
  AND2_X1 U6257 ( .A1(n5357), .A2(n5302), .ZN(n5313) );
  AOI21_X1 U6258 ( .B1(REIP_REG_13__SCAN_IN), .B2(n5313), .A(
        REIP_REG_14__SCAN_IN), .ZN(n5311) );
  OAI22_X1 U6259 ( .A1(n5304), .A2(n5374), .B1(n5367), .B2(n5303), .ZN(n5305)
         );
  AOI211_X1 U6260 ( .C1(n5368), .C2(EBX_REG_14__SCAN_IN), .A(n5344), .B(n5305), 
        .ZN(n5310) );
  INV_X1 U6261 ( .A(n5306), .ZN(n5308) );
  AOI22_X1 U6262 ( .A1(n5308), .A2(n5351), .B1(n5340), .B2(n5307), .ZN(n5309)
         );
  OAI211_X1 U6263 ( .C1(n5312), .C2(n5311), .A(n5310), .B(n5309), .ZN(U2813)
         );
  INV_X1 U6264 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6296) );
  AOI22_X1 U6265 ( .A1(n5377), .A2(n5387), .B1(n5313), .B2(n6296), .ZN(n5315)
         );
  AOI21_X1 U6266 ( .B1(n5364), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5344), 
        .ZN(n5314) );
  OAI211_X1 U6267 ( .C1(n5390), .C2(n5361), .A(n5315), .B(n5314), .ZN(n5316)
         );
  AOI21_X1 U6268 ( .B1(n5388), .B2(n5351), .A(n5316), .ZN(n5319) );
  OAI21_X1 U6269 ( .B1(n5317), .B2(n5324), .A(REIP_REG_13__SCAN_IN), .ZN(n5318) );
  OAI211_X1 U6270 ( .C1(n5386), .C2(n5320), .A(n5319), .B(n5318), .ZN(U2814)
         );
  NAND3_X1 U6271 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n5330), .ZN(n5329) );
  AOI21_X1 U6272 ( .B1(n5323), .B2(n5322), .A(n5321), .ZN(n5556) );
  AOI22_X1 U6273 ( .A1(n5377), .A2(n5556), .B1(REIP_REG_11__SCAN_IN), .B2(
        n5324), .ZN(n5325) );
  OAI21_X1 U6274 ( .B1(n5392), .B2(n5361), .A(n5325), .ZN(n5326) );
  AOI211_X1 U6275 ( .C1(n5364), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5344), 
        .B(n5326), .ZN(n5328) );
  AOI22_X1 U6276 ( .A1(n5518), .A2(n5351), .B1(n5340), .B2(n5516), .ZN(n5327)
         );
  OAI211_X1 U6277 ( .C1(REIP_REG_11__SCAN_IN), .C2(n5329), .A(n5328), .B(n5327), .ZN(U2816) );
  INV_X1 U6278 ( .A(n5330), .ZN(n5343) );
  INV_X1 U6279 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6290) );
  OR2_X1 U6280 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  AND2_X1 U6281 ( .A1(n5334), .A2(n5333), .ZN(n5578) );
  AOI22_X1 U6282 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5368), .B1(n5377), .B2(n5578), 
        .ZN(n5335) );
  OAI21_X1 U6283 ( .B1(n6290), .B2(n5336), .A(n5335), .ZN(n5337) );
  AOI211_X1 U6284 ( .C1(n5364), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5344), 
        .B(n5337), .ZN(n5342) );
  INV_X1 U6285 ( .A(n5338), .ZN(n5395) );
  AOI22_X1 U6286 ( .A1(n5395), .A2(n5351), .B1(n5340), .B2(n5339), .ZN(n5341)
         );
  OAI211_X1 U6287 ( .C1(REIP_REG_9__SCAN_IN), .C2(n5343), .A(n5342), .B(n5341), 
        .ZN(U2818) );
  AOI21_X1 U6288 ( .B1(n5364), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5344), 
        .ZN(n5347) );
  INV_X1 U6289 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6285) );
  NAND3_X1 U6290 ( .A1(n5357), .A2(n5345), .A3(n6285), .ZN(n5346) );
  OAI211_X1 U6291 ( .C1(n5348), .C2(n5367), .A(n5347), .B(n5346), .ZN(n5349)
         );
  AOI21_X1 U6292 ( .B1(EBX_REG_6__SCAN_IN), .B2(n5368), .A(n5349), .ZN(n5353)
         );
  AOI22_X1 U6293 ( .A1(n5522), .A2(n5351), .B1(REIP_REG_6__SCAN_IN), .B2(n5350), .ZN(n5352) );
  OAI211_X1 U6294 ( .C1(n5526), .C2(n5386), .A(n5353), .B(n5352), .ZN(U2821)
         );
  AOI22_X1 U6295 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5355), .B1(n5354), .B2(n5378), .ZN(n5366) );
  INV_X1 U6296 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6283) );
  NAND3_X1 U6297 ( .A1(n5357), .A2(n6283), .A3(n5356), .ZN(n5358) );
  OAI211_X1 U6298 ( .C1(n5361), .C2(n5360), .A(n5359), .B(n5358), .ZN(n5363)
         );
  OAI22_X1 U6299 ( .A1(n5531), .A2(n5382), .B1(n5535), .B2(n5386), .ZN(n5362)
         );
  AOI211_X1 U6300 ( .C1(PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n5364), .A(n5363), 
        .B(n5362), .ZN(n5365) );
  OAI211_X1 U6301 ( .C1(n5367), .C2(n5611), .A(n5366), .B(n5365), .ZN(U2823)
         );
  NAND2_X1 U6302 ( .A1(n5368), .A2(EBX_REG_1__SCAN_IN), .ZN(n5369) );
  AND2_X1 U6303 ( .A1(n5370), .A2(n5369), .ZN(n5385) );
  INV_X1 U6304 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U6305 ( .A1(n5371), .A2(REIP_REG_1__SCAN_IN), .ZN(n5372) );
  OAI21_X1 U6306 ( .B1(n5374), .B2(n5373), .A(n5372), .ZN(n5375) );
  AOI21_X1 U6307 ( .B1(n5377), .B2(n5376), .A(n5375), .ZN(n5380) );
  NAND2_X1 U6308 ( .A1(n5378), .A2(n5797), .ZN(n5379) );
  OAI211_X1 U6309 ( .C1(n5382), .C2(n5381), .A(n5380), .B(n5379), .ZN(n5383)
         );
  INV_X1 U6310 ( .A(n5383), .ZN(n5384) );
  OAI211_X1 U6311 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n5386), .A(n5385), 
        .B(n5384), .ZN(U2826) );
  AOI22_X1 U6312 ( .A1(n5388), .A2(n5394), .B1(n5393), .B2(n5387), .ZN(n5389)
         );
  OAI21_X1 U6313 ( .B1(n5398), .B2(n5390), .A(n5389), .ZN(U2846) );
  AOI22_X1 U6314 ( .A1(n5518), .A2(n5394), .B1(n5393), .B2(n5556), .ZN(n5391)
         );
  OAI21_X1 U6315 ( .B1(n5398), .B2(n5392), .A(n5391), .ZN(U2848) );
  AOI22_X1 U6316 ( .A1(n5395), .A2(n5394), .B1(n5393), .B2(n5578), .ZN(n5396)
         );
  OAI21_X1 U6317 ( .B1(n5398), .B2(n5397), .A(n5396), .ZN(U2850) );
  AOI22_X1 U6318 ( .A1(n5399), .A2(n5406), .B1(n5405), .B2(DATAI_18_), .ZN(
        n5401) );
  AOI22_X1 U6319 ( .A1(n5409), .A2(DATAI_2_), .B1(n5408), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U6320 ( .A1(n5401), .A2(n5400), .ZN(U2873) );
  AOI22_X1 U6321 ( .A1(n5402), .A2(n5406), .B1(n5405), .B2(DATAI_17_), .ZN(
        n5404) );
  AOI22_X1 U6322 ( .A1(n5409), .A2(DATAI_1_), .B1(n5408), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6323 ( .A1(n5404), .A2(n5403), .ZN(U2874) );
  AOI22_X1 U6324 ( .A1(n5407), .A2(n5406), .B1(n5405), .B2(DATAI_16_), .ZN(
        n5411) );
  AOI22_X1 U6325 ( .A1(n5409), .A2(DATAI_0_), .B1(n5408), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6326 ( .A1(n5411), .A2(n5410), .ZN(U2875) );
  INV_X1 U6327 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6437) );
  AOI22_X1 U6328 ( .A1(n6237), .A2(LWORD_REG_15__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5413) );
  OAI21_X1 U6329 ( .B1(n6437), .B2(n5430), .A(n5413), .ZN(U2908) );
  INV_X1 U6330 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5508) );
  AOI22_X1 U6331 ( .A1(n6237), .A2(LWORD_REG_14__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5414) );
  OAI21_X1 U6332 ( .B1(n5508), .B2(n5430), .A(n5414), .ZN(U2909) );
  INV_X1 U6333 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5504) );
  AOI22_X1 U6334 ( .A1(n6237), .A2(LWORD_REG_13__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5415) );
  OAI21_X1 U6335 ( .B1(n5504), .B2(n5430), .A(n5415), .ZN(U2910) );
  INV_X1 U6336 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5501) );
  AOI22_X1 U6337 ( .A1(n6237), .A2(LWORD_REG_12__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5416) );
  OAI21_X1 U6338 ( .B1(n5501), .B2(n5430), .A(n5416), .ZN(U2911) );
  INV_X1 U6339 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5498) );
  AOI22_X1 U6340 ( .A1(n6237), .A2(LWORD_REG_11__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5417) );
  OAI21_X1 U6341 ( .B1(n5498), .B2(n5430), .A(n5417), .ZN(U2912) );
  INV_X1 U6342 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6443) );
  AOI22_X1 U6343 ( .A1(n6237), .A2(LWORD_REG_10__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5418) );
  OAI21_X1 U6344 ( .B1(n6443), .B2(n5430), .A(n5418), .ZN(U2913) );
  INV_X1 U6345 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5492) );
  AOI22_X1 U6346 ( .A1(n6237), .A2(LWORD_REG_9__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5419) );
  OAI21_X1 U6347 ( .B1(n5492), .B2(n5430), .A(n5419), .ZN(U2914) );
  INV_X1 U6348 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5489) );
  AOI22_X1 U6349 ( .A1(n6237), .A2(LWORD_REG_8__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5420) );
  OAI21_X1 U6350 ( .B1(n5489), .B2(n5430), .A(n5420), .ZN(U2915) );
  AOI22_X1 U6351 ( .A1(n6237), .A2(LWORD_REG_7__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5421) );
  OAI21_X1 U6352 ( .B1(n3510), .B2(n5430), .A(n5421), .ZN(U2916) );
  AOI22_X1 U6353 ( .A1(n6237), .A2(LWORD_REG_6__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5422) );
  OAI21_X1 U6354 ( .B1(n4389), .B2(n5430), .A(n5422), .ZN(U2917) );
  AOI22_X1 U6355 ( .A1(n6237), .A2(LWORD_REG_5__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5424) );
  OAI21_X1 U6356 ( .B1(n5482), .B2(n5430), .A(n5424), .ZN(U2918) );
  AOI22_X1 U6357 ( .A1(n6237), .A2(LWORD_REG_4__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5425) );
  OAI21_X1 U6358 ( .B1(n5479), .B2(n5430), .A(n5425), .ZN(U2919) );
  AOI22_X1 U6359 ( .A1(n6237), .A2(LWORD_REG_3__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5426) );
  OAI21_X1 U6360 ( .B1(n6489), .B2(n5430), .A(n5426), .ZN(U2920) );
  AOI22_X1 U6361 ( .A1(n6237), .A2(LWORD_REG_2__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5427) );
  OAI21_X1 U6362 ( .B1(n5474), .B2(n5430), .A(n5427), .ZN(U2921) );
  AOI22_X1 U6363 ( .A1(n6237), .A2(LWORD_REG_1__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5428) );
  OAI21_X1 U6364 ( .B1(n5471), .B2(n5430), .A(n5428), .ZN(U2922) );
  AOI22_X1 U6365 ( .A1(n6237), .A2(LWORD_REG_0__SCAN_IN), .B1(n5423), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5429) );
  OAI21_X1 U6366 ( .B1(n5468), .B2(n5430), .A(n5429), .ZN(U2923) );
  OAI21_X1 U6367 ( .B1(n6364), .B2(n6271), .A(n5431), .ZN(n5496) );
  INV_X1 U6368 ( .A(n5463), .ZN(n5509) );
  AND2_X1 U6369 ( .A1(n5509), .A2(DATAI_0_), .ZN(n5466) );
  AOI21_X1 U6370 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n5506), .A(n5466), .ZN(n5432) );
  OAI21_X1 U6371 ( .B1(n5433), .B2(n5511), .A(n5432), .ZN(U2924) );
  AND2_X1 U6372 ( .A1(n5509), .A2(DATAI_1_), .ZN(n5469) );
  AOI21_X1 U6373 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n5506), .A(n5469), .ZN(n5434) );
  OAI21_X1 U6374 ( .B1(n5435), .B2(n5511), .A(n5434), .ZN(U2925) );
  AND2_X1 U6375 ( .A1(n5509), .A2(DATAI_2_), .ZN(n5472) );
  AOI21_X1 U6376 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n5506), .A(n5472), .ZN(n5436) );
  OAI21_X1 U6377 ( .B1(n5437), .B2(n5511), .A(n5436), .ZN(U2926) );
  AND2_X1 U6378 ( .A1(n5509), .A2(DATAI_3_), .ZN(n5475) );
  AOI21_X1 U6379 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n5506), .A(n5475), .ZN(n5438) );
  OAI21_X1 U6380 ( .B1(n5439), .B2(n5511), .A(n5438), .ZN(U2927) );
  AND2_X1 U6381 ( .A1(n5509), .A2(DATAI_4_), .ZN(n5477) );
  AOI21_X1 U6382 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n5506), .A(n5477), .ZN(n5440) );
  OAI21_X1 U6383 ( .B1(n3775), .B2(n5511), .A(n5440), .ZN(U2928) );
  AND2_X1 U6384 ( .A1(n5509), .A2(DATAI_5_), .ZN(n5480) );
  AOI21_X1 U6385 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n5506), .A(n5480), .ZN(n5441) );
  OAI21_X1 U6386 ( .B1(n6441), .B2(n5511), .A(n5441), .ZN(U2929) );
  NOR2_X1 U6387 ( .A1(n5463), .A2(n5442), .ZN(n5483) );
  AOI21_X1 U6388 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n5506), .A(n5483), .ZN(n5443) );
  OAI21_X1 U6389 ( .B1(n5444), .B2(n5511), .A(n5443), .ZN(U2930) );
  AND2_X1 U6390 ( .A1(n5509), .A2(DATAI_7_), .ZN(n5485) );
  AOI21_X1 U6391 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n5506), .A(n5485), .ZN(n5445) );
  OAI21_X1 U6392 ( .B1(n5446), .B2(n5511), .A(n5445), .ZN(U2931) );
  INV_X1 U6393 ( .A(DATAI_8_), .ZN(n5447) );
  NOR2_X1 U6394 ( .A1(n5463), .A2(n5447), .ZN(n5487) );
  AOI21_X1 U6395 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n5506), .A(n5487), .ZN(n5448) );
  OAI21_X1 U6396 ( .B1(n6453), .B2(n5511), .A(n5448), .ZN(U2932) );
  INV_X1 U6397 ( .A(DATAI_9_), .ZN(n5449) );
  NOR2_X1 U6398 ( .A1(n5463), .A2(n5449), .ZN(n5490) );
  AOI21_X1 U6399 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n5506), .A(n5490), .ZN(n5450) );
  OAI21_X1 U6400 ( .B1(n3876), .B2(n5511), .A(n5450), .ZN(U2933) );
  INV_X1 U6401 ( .A(DATAI_10_), .ZN(n5451) );
  NOR2_X1 U6402 ( .A1(n5463), .A2(n5451), .ZN(n5493) );
  AOI21_X1 U6403 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n5506), .A(n5493), .ZN(
        n5452) );
  OAI21_X1 U6404 ( .B1(n5453), .B2(n5511), .A(n5452), .ZN(U2934) );
  INV_X1 U6405 ( .A(DATAI_11_), .ZN(n5454) );
  NOR2_X1 U6406 ( .A1(n5463), .A2(n5454), .ZN(n5495) );
  AOI21_X1 U6407 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n5506), .A(n5495), .ZN(
        n5455) );
  OAI21_X1 U6408 ( .B1(n5456), .B2(n5511), .A(n5455), .ZN(U2935) );
  INV_X1 U6409 ( .A(DATAI_12_), .ZN(n5457) );
  NOR2_X1 U6410 ( .A1(n5463), .A2(n5457), .ZN(n5499) );
  AOI21_X1 U6411 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n5496), .A(n5499), .ZN(
        n5458) );
  OAI21_X1 U6412 ( .B1(n6526), .B2(n5511), .A(n5458), .ZN(U2936) );
  INV_X1 U6413 ( .A(DATAI_13_), .ZN(n5459) );
  NOR2_X1 U6414 ( .A1(n5463), .A2(n5459), .ZN(n5502) );
  AOI21_X1 U6415 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n5496), .A(n5502), .ZN(
        n5460) );
  OAI21_X1 U6416 ( .B1(n5461), .B2(n5511), .A(n5460), .ZN(U2937) );
  INV_X1 U6417 ( .A(DATAI_14_), .ZN(n5462) );
  NOR2_X1 U6418 ( .A1(n5463), .A2(n5462), .ZN(n5505) );
  AOI21_X1 U6419 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n5496), .A(n5505), .ZN(
        n5464) );
  OAI21_X1 U6420 ( .B1(n5465), .B2(n5511), .A(n5464), .ZN(U2938) );
  AOI21_X1 U6421 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n5506), .A(n5466), .ZN(n5467) );
  OAI21_X1 U6422 ( .B1(n5468), .B2(n5511), .A(n5467), .ZN(U2939) );
  AOI21_X1 U6423 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n5506), .A(n5469), .ZN(n5470) );
  OAI21_X1 U6424 ( .B1(n5471), .B2(n5511), .A(n5470), .ZN(U2940) );
  AOI21_X1 U6425 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n5506), .A(n5472), .ZN(n5473) );
  OAI21_X1 U6426 ( .B1(n5474), .B2(n5511), .A(n5473), .ZN(U2941) );
  AOI21_X1 U6427 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n5506), .A(n5475), .ZN(n5476) );
  OAI21_X1 U6428 ( .B1(n6489), .B2(n5511), .A(n5476), .ZN(U2942) );
  AOI21_X1 U6429 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n5506), .A(n5477), .ZN(n5478) );
  OAI21_X1 U6430 ( .B1(n5479), .B2(n5511), .A(n5478), .ZN(U2943) );
  AOI21_X1 U6431 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n5506), .A(n5480), .ZN(n5481) );
  OAI21_X1 U6432 ( .B1(n5482), .B2(n5511), .A(n5481), .ZN(U2944) );
  AOI21_X1 U6433 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n5496), .A(n5483), .ZN(n5484) );
  OAI21_X1 U6434 ( .B1(n4389), .B2(n5511), .A(n5484), .ZN(U2945) );
  AOI21_X1 U6435 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n5496), .A(n5485), .ZN(n5486) );
  OAI21_X1 U6436 ( .B1(n3510), .B2(n5511), .A(n5486), .ZN(U2946) );
  AOI21_X1 U6437 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n5496), .A(n5487), .ZN(n5488) );
  OAI21_X1 U6438 ( .B1(n5489), .B2(n5511), .A(n5488), .ZN(U2947) );
  AOI21_X1 U6439 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n5496), .A(n5490), .ZN(n5491) );
  OAI21_X1 U6440 ( .B1(n5492), .B2(n5511), .A(n5491), .ZN(U2948) );
  AOI21_X1 U6441 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n5496), .A(n5493), .ZN(
        n5494) );
  OAI21_X1 U6442 ( .B1(n6443), .B2(n5511), .A(n5494), .ZN(U2949) );
  AOI21_X1 U6443 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n5496), .A(n5495), .ZN(
        n5497) );
  OAI21_X1 U6444 ( .B1(n5498), .B2(n5511), .A(n5497), .ZN(U2950) );
  AOI21_X1 U6445 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n5506), .A(n5499), .ZN(
        n5500) );
  OAI21_X1 U6446 ( .B1(n5501), .B2(n5511), .A(n5500), .ZN(U2951) );
  AOI21_X1 U6447 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n5496), .A(n5502), .ZN(
        n5503) );
  OAI21_X1 U6448 ( .B1(n5504), .B2(n5511), .A(n5503), .ZN(U2952) );
  AOI21_X1 U6449 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n5506), .A(n5505), .ZN(
        n5507) );
  OAI21_X1 U6450 ( .B1(n5508), .B2(n5511), .A(n5507), .ZN(U2953) );
  AOI22_X1 U6451 ( .A1(n5496), .A2(LWORD_REG_15__SCAN_IN), .B1(n5509), .B2(
        DATAI_15_), .ZN(n5510) );
  OAI21_X1 U6452 ( .B1(n6437), .B2(n5511), .A(n5510), .ZN(U2954) );
  NAND2_X1 U6453 ( .A1(n5512), .A2(n5513), .ZN(n5515) );
  XNOR2_X1 U6454 ( .A(n5203), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5514)
         );
  XNOR2_X1 U6455 ( .A(n5515), .B(n5514), .ZN(n5561) );
  AOI22_X1 U6456 ( .A1(n5630), .A2(REIP_REG_11__SCAN_IN), .B1(n5536), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5520) );
  AOI22_X1 U6457 ( .A1(n5518), .A2(n5702), .B1(n5517), .B2(n5516), .ZN(n5519)
         );
  OAI211_X1 U6458 ( .C1(n5561), .C2(n5555), .A(n5520), .B(n5519), .ZN(U2975)
         );
  AOI22_X1 U6459 ( .A1(n5630), .A2(REIP_REG_6__SCAN_IN), .B1(n5536), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5525) );
  INV_X1 U6460 ( .A(n5521), .ZN(n5523) );
  AOI22_X1 U6461 ( .A1(n5523), .A2(n5541), .B1(n5702), .B2(n5522), .ZN(n5524)
         );
  OAI211_X1 U6462 ( .C1(n5546), .C2(n5526), .A(n5525), .B(n5524), .ZN(U2980)
         );
  AOI22_X1 U6463 ( .A1(n5630), .A2(REIP_REG_4__SCAN_IN), .B1(n5536), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5534) );
  OR2_X1 U6464 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  NAND2_X1 U6465 ( .A1(n5527), .A2(n5530), .ZN(n5616) );
  OAI22_X1 U6466 ( .A1(n5616), .A2(n5555), .B1(n5531), .B2(n5692), .ZN(n5532)
         );
  INV_X1 U6467 ( .A(n5532), .ZN(n5533) );
  OAI211_X1 U6468 ( .C1(n5546), .C2(n5535), .A(n5534), .B(n5533), .ZN(U2982)
         );
  AOI22_X1 U6469 ( .A1(n5630), .A2(REIP_REG_2__SCAN_IN), .B1(n5536), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5544) );
  INV_X1 U6470 ( .A(n5537), .ZN(n5542) );
  XOR2_X1 U6471 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .B(n5538), .Z(n5540) );
  XNOR2_X1 U6472 ( .A(n5540), .B(n5539), .ZN(n5637) );
  AOI22_X1 U6473 ( .A1(n5542), .A2(n5702), .B1(n5637), .B2(n5541), .ZN(n5543)
         );
  OAI211_X1 U6474 ( .C1(n5546), .C2(n5545), .A(n5544), .B(n5543), .ZN(U2984)
         );
  OAI21_X1 U6475 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5548), .A(n5547), 
        .ZN(n5655) );
  INV_X1 U6476 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6359) );
  NOR2_X1 U6477 ( .A1(n5612), .A2(n6359), .ZN(n5646) );
  INV_X1 U6478 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5549) );
  AOI21_X1 U6479 ( .B1(n5551), .B2(n5550), .A(n5549), .ZN(n5552) );
  AOI211_X1 U6480 ( .C1(n5553), .C2(n5702), .A(n5646), .B(n5552), .ZN(n5554)
         );
  OAI21_X1 U6481 ( .B1(n5555), .B2(n5655), .A(n5554), .ZN(U2986) );
  AOI22_X1 U6482 ( .A1(n5649), .A2(n5556), .B1(n5630), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5560) );
  AOI22_X1 U6483 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5558), .B1(n5557), .B2(n3422), .ZN(n5559) );
  OAI211_X1 U6484 ( .C1(n5561), .C2(n5654), .A(n5560), .B(n5559), .ZN(U3007)
         );
  INV_X1 U6485 ( .A(n5562), .ZN(n5564) );
  NOR2_X1 U6486 ( .A1(n5564), .A2(n5563), .ZN(n5596) );
  NAND2_X1 U6487 ( .A1(n5588), .A2(n5596), .ZN(n5583) );
  AOI22_X1 U6488 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n3421), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5565), .ZN(n5576) );
  AOI21_X1 U6489 ( .B1(n5567), .B2(n5649), .A(n5566), .ZN(n5575) );
  AOI22_X1 U6490 ( .A1(n5571), .A2(n5570), .B1(n5569), .B2(n5568), .ZN(n5600)
         );
  OAI21_X1 U6491 ( .B1(n5572), .B2(n5588), .A(n5600), .ZN(n5579) );
  AOI22_X1 U6492 ( .A1(n5573), .A2(n5636), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5579), .ZN(n5574) );
  OAI211_X1 U6493 ( .C1(n5583), .C2(n5576), .A(n5575), .B(n5574), .ZN(U3008)
         );
  AOI21_X1 U6494 ( .B1(n5649), .B2(n5578), .A(n5577), .ZN(n5582) );
  AOI22_X1 U6495 ( .A1(n5580), .A2(n5636), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n5579), .ZN(n5581) );
  OAI211_X1 U6496 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n5583), .A(n5582), 
        .B(n5581), .ZN(U3009) );
  OAI222_X1 U6497 ( .A1(n5586), .A2(n5585), .B1(n5612), .B2(n6288), .C1(n5654), 
        .C2(n5584), .ZN(n5587) );
  INV_X1 U6498 ( .A(n5587), .ZN(n5591) );
  INV_X1 U6499 ( .A(n5588), .ZN(n5589) );
  OAI211_X1 U6500 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5596), .B(n5589), .ZN(n5590) );
  OAI211_X1 U6501 ( .C1(n5600), .C2(n5592), .A(n5591), .B(n5590), .ZN(U3010)
         );
  AOI21_X1 U6502 ( .B1(n5649), .B2(n5594), .A(n5593), .ZN(n5599) );
  INV_X1 U6503 ( .A(n5595), .ZN(n5597) );
  AOI22_X1 U6504 ( .A1(n5597), .A2(n5636), .B1(n5596), .B2(n6482), .ZN(n5598)
         );
  OAI211_X1 U6505 ( .C1(n5600), .C2(n6482), .A(n5599), .B(n5598), .ZN(U3011)
         );
  AOI21_X1 U6506 ( .B1(n5610), .B2(n5625), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n5607) );
  INV_X1 U6507 ( .A(n5601), .ZN(n5604) );
  INV_X1 U6508 ( .A(n5602), .ZN(n5603) );
  AOI22_X1 U6509 ( .A1(n5604), .A2(n5636), .B1(n5649), .B2(n5603), .ZN(n5606)
         );
  NAND2_X1 U6510 ( .A1(n5630), .A2(REIP_REG_5__SCAN_IN), .ZN(n5605) );
  OAI211_X1 U6511 ( .C1(n5608), .C2(n5607), .A(n5606), .B(n5605), .ZN(U3013)
         );
  AOI21_X1 U6512 ( .B1(n5632), .B2(n5634), .A(n5635), .ZN(n5629) );
  AOI211_X1 U6513 ( .C1(n5628), .C2(n5620), .A(n5610), .B(n5609), .ZN(n5618)
         );
  INV_X1 U6514 ( .A(n5611), .ZN(n5614) );
  NOR2_X1 U6515 ( .A1(n5612), .A2(n6283), .ZN(n5613) );
  AOI21_X1 U6516 ( .B1(n5649), .B2(n5614), .A(n5613), .ZN(n5615) );
  OAI21_X1 U6517 ( .B1(n5616), .B2(n5654), .A(n5615), .ZN(n5617) );
  NOR2_X1 U6518 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  OAI21_X1 U6519 ( .B1(n5629), .B2(n5620), .A(n5619), .ZN(U3014) );
  AOI21_X1 U6520 ( .B1(n5649), .B2(n5622), .A(n5621), .ZN(n5627) );
  INV_X1 U6521 ( .A(n5623), .ZN(n5624) );
  AOI22_X1 U6522 ( .A1(n5625), .A2(n5628), .B1(n5624), .B2(n5636), .ZN(n5626)
         );
  OAI211_X1 U6523 ( .C1(n5629), .C2(n5628), .A(n5627), .B(n5626), .ZN(U3015)
         );
  AOI22_X1 U6524 ( .A1(n5649), .A2(n5631), .B1(n5630), .B2(REIP_REG_2__SCAN_IN), .ZN(n5643) );
  OAI221_X1 U6525 ( .B1(n5634), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .C1(n5634), .C2(n5633), .A(n5632), .ZN(n5642) );
  AOI22_X1 U6526 ( .A1(n5637), .A2(n5636), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n5635), .ZN(n5641) );
  INV_X1 U6527 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5638) );
  NAND3_X1 U6528 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5639), .A3(n5638), 
        .ZN(n5640) );
  NAND4_X1 U6529 ( .A1(n5643), .A2(n5642), .A3(n5641), .A4(n5640), .ZN(U3016)
         );
  INV_X1 U6530 ( .A(n5644), .ZN(n5648) );
  OR2_X1 U6531 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  AOI21_X1 U6532 ( .B1(n5649), .B2(n5648), .A(n5647), .ZN(n5653) );
  OAI21_X1 U6533 ( .B1(n5651), .B2(n5650), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5652) );
  OAI211_X1 U6534 ( .C1(n5655), .C2(n5654), .A(n5653), .B(n5652), .ZN(U3018)
         );
  NOR2_X1 U6535 ( .A1(n5656), .A2(n6348), .ZN(U3019) );
  INV_X1 U6536 ( .A(DATAI_24_), .ZN(n5657) );
  NOR2_X1 U6537 ( .A1(n5692), .A2(n5657), .ZN(n6158) );
  INV_X1 U6538 ( .A(n6158), .ZN(n6115) );
  AND2_X1 U6539 ( .A1(n4338), .A2(n5917), .ZN(n5658) );
  NAND2_X1 U6540 ( .A1(n5663), .A2(n5658), .ZN(n6150) );
  NOR2_X2 U6541 ( .A1(n5659), .A2(n5703), .ZN(n6149) );
  NAND2_X1 U6542 ( .A1(n2965), .A2(n5855), .ZN(n5949) );
  NOR2_X1 U6543 ( .A1(n4264), .A2(n5949), .ZN(n5711) );
  INV_X1 U6544 ( .A(n5711), .ZN(n5660) );
  AND2_X1 U6545 ( .A1(n5665), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6105) );
  INV_X1 U6546 ( .A(n6105), .ZN(n6049) );
  NOR2_X1 U6547 ( .A1(n5914), .A2(n5913), .ZN(n5666) );
  INV_X1 U6548 ( .A(n5666), .ZN(n5799) );
  OAI22_X1 U6549 ( .A1(n5660), .A2(n6370), .B1(n6049), .B2(n5799), .ZN(n5706)
         );
  NOR2_X2 U6550 ( .A1(n5704), .A2(n5662), .ZN(n6148) );
  NAND3_X1 U6551 ( .A1(n3479), .A2(n6213), .A3(n6218), .ZN(n5715) );
  NOR2_X1 U6552 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5715), .ZN(n5705)
         );
  AOI22_X1 U6553 ( .A1(n6149), .A2(n5706), .B1(n6148), .B2(n5705), .ZN(n5672)
         );
  NAND2_X1 U6554 ( .A1(n5712), .A2(n6071), .ZN(n5732) );
  INV_X1 U6555 ( .A(n6192), .ZN(n6204) );
  NOR3_X1 U6556 ( .A1(n5734), .A2(n6204), .A3(n6370), .ZN(n5664) );
  NOR2_X1 U6557 ( .A1(n5664), .A2(n5919), .ZN(n5669) );
  INV_X1 U6558 ( .A(n5705), .ZN(n5667) );
  NOR2_X1 U6559 ( .A1(n5665), .A2(n3558), .ZN(n5923) );
  OAI21_X1 U6560 ( .B1(n5666), .B2(n3558), .A(n5921), .ZN(n5802) );
  AOI211_X1 U6561 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5667), .A(n5923), .B(
        n5802), .ZN(n5668) );
  INV_X1 U6562 ( .A(DATAI_16_), .ZN(n5670) );
  NOR2_X2 U6563 ( .A1(n5692), .A2(n5670), .ZN(n6112) );
  AOI22_X1 U6564 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n5708), .B1(n6112), 
        .B2(n5734), .ZN(n5671) );
  OAI211_X1 U6565 ( .C1(n6115), .C2(n6192), .A(n5672), .B(n5671), .ZN(U3020)
         );
  INV_X1 U6566 ( .A(DATAI_25_), .ZN(n5673) );
  NOR2_X1 U6567 ( .A1(n5692), .A2(n5673), .ZN(n6164) );
  INV_X1 U6568 ( .A(n6164), .ZN(n6119) );
  NOR2_X2 U6569 ( .A1(n6474), .A2(n5703), .ZN(n6163) );
  NOR2_X2 U6570 ( .A1(n5704), .A2(n3160), .ZN(n6162) );
  AOI22_X1 U6571 ( .A1(n6163), .A2(n5706), .B1(n6162), .B2(n5705), .ZN(n5676)
         );
  INV_X1 U6572 ( .A(DATAI_17_), .ZN(n5674) );
  AOI22_X1 U6573 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n5708), .B1(n6116), 
        .B2(n5734), .ZN(n5675) );
  OAI211_X1 U6574 ( .C1(n6119), .C2(n6192), .A(n5676), .B(n5675), .ZN(U3021)
         );
  INV_X1 U6575 ( .A(DATAI_26_), .ZN(n5677) );
  NOR2_X1 U6576 ( .A1(n5692), .A2(n5677), .ZN(n6170) );
  INV_X1 U6577 ( .A(n6170), .ZN(n6123) );
  NOR2_X2 U6578 ( .A1(n5678), .A2(n5703), .ZN(n6169) );
  NOR2_X2 U6579 ( .A1(n5704), .A2(n3150), .ZN(n6168) );
  AOI22_X1 U6580 ( .A1(n6169), .A2(n5706), .B1(n6168), .B2(n5705), .ZN(n5681)
         );
  INV_X1 U6581 ( .A(DATAI_18_), .ZN(n5679) );
  NOR2_X2 U6582 ( .A1(n5692), .A2(n5679), .ZN(n6120) );
  AOI22_X1 U6583 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n5708), .B1(n6120), 
        .B2(n5734), .ZN(n5680) );
  OAI211_X1 U6584 ( .C1(n6123), .C2(n6192), .A(n5681), .B(n5680), .ZN(U3022)
         );
  INV_X1 U6585 ( .A(DATAI_27_), .ZN(n5682) );
  NOR2_X1 U6586 ( .A1(n5692), .A2(n5682), .ZN(n6176) );
  INV_X1 U6587 ( .A(n6176), .ZN(n6127) );
  NOR2_X2 U6588 ( .A1(n5683), .A2(n5703), .ZN(n6175) );
  NOR2_X2 U6589 ( .A1(n5704), .A2(n5684), .ZN(n6174) );
  AOI22_X1 U6590 ( .A1(n6175), .A2(n5706), .B1(n6174), .B2(n5705), .ZN(n5687)
         );
  INV_X1 U6591 ( .A(DATAI_19_), .ZN(n5685) );
  NOR2_X1 U6592 ( .A1(n5692), .A2(n5685), .ZN(n6124) );
  AOI22_X1 U6593 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n5708), .B1(n6124), 
        .B2(n5734), .ZN(n5686) );
  OAI211_X1 U6594 ( .C1(n6127), .C2(n6192), .A(n5687), .B(n5686), .ZN(U3023)
         );
  INV_X1 U6595 ( .A(DATAI_28_), .ZN(n5688) );
  NOR2_X1 U6596 ( .A1(n5692), .A2(n5688), .ZN(n6182) );
  INV_X1 U6597 ( .A(n6182), .ZN(n6131) );
  NOR2_X2 U6598 ( .A1(n5689), .A2(n5703), .ZN(n6181) );
  NOR2_X2 U6599 ( .A1(n5704), .A2(n5690), .ZN(n6180) );
  AOI22_X1 U6600 ( .A1(n6181), .A2(n5706), .B1(n6180), .B2(n5705), .ZN(n5694)
         );
  INV_X1 U6601 ( .A(DATAI_20_), .ZN(n5691) );
  NOR2_X1 U6602 ( .A1(n5692), .A2(n5691), .ZN(n6128) );
  AOI22_X1 U6603 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5708), .B1(n6128), 
        .B2(n5734), .ZN(n5693) );
  OAI211_X1 U6604 ( .C1(n6131), .C2(n6192), .A(n5694), .B(n5693), .ZN(U3024)
         );
  INV_X1 U6605 ( .A(DATAI_29_), .ZN(n5695) );
  NOR2_X1 U6606 ( .A1(n5692), .A2(n5695), .ZN(n6189) );
  INV_X1 U6607 ( .A(n6189), .ZN(n6135) );
  NOR2_X2 U6608 ( .A1(n5696), .A2(n5703), .ZN(n6187) );
  NOR2_X2 U6609 ( .A1(n5704), .A2(n3146), .ZN(n6186) );
  AOI22_X1 U6610 ( .A1(n6187), .A2(n5706), .B1(n6186), .B2(n5705), .ZN(n5699)
         );
  INV_X1 U6611 ( .A(DATAI_21_), .ZN(n5697) );
  NOR2_X1 U6612 ( .A1(n5692), .A2(n5697), .ZN(n6132) );
  AOI22_X1 U6613 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n5708), .B1(n6132), 
        .B2(n5734), .ZN(n5698) );
  OAI211_X1 U6614 ( .C1(n6135), .C2(n6192), .A(n5699), .B(n5698), .ZN(U3025)
         );
  NAND2_X1 U6615 ( .A1(n5702), .A2(DATAI_30_), .ZN(n6199) );
  NOR2_X2 U6616 ( .A1(n5704), .A2(n3131), .ZN(n6195) );
  AOI22_X1 U6617 ( .A1(n6195), .A2(n5705), .B1(n6194), .B2(n5706), .ZN(n5701)
         );
  AOI22_X1 U6618 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n5708), .B1(n6196), 
        .B2(n5734), .ZN(n5700) );
  OAI211_X1 U6619 ( .C1(n6199), .C2(n6192), .A(n5701), .B(n5700), .ZN(U3026)
         );
  NAND2_X1 U6620 ( .A1(n5702), .A2(DATAI_31_), .ZN(n6210) );
  NOR2_X2 U6621 ( .A1(n6479), .A2(n5703), .ZN(n6203) );
  NOR2_X2 U6622 ( .A1(n5704), .A2(n3132), .ZN(n6200) );
  AOI22_X1 U6623 ( .A1(n6203), .A2(n5706), .B1(n6200), .B2(n5705), .ZN(n5710)
         );
  INV_X1 U6624 ( .A(DATAI_23_), .ZN(n5707) );
  NOR2_X2 U6625 ( .A1(n5692), .A2(n5707), .ZN(n6205) );
  AOI22_X1 U6626 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n5708), .B1(n6205), 
        .B2(n5734), .ZN(n5709) );
  OAI211_X1 U6627 ( .C1(n6210), .C2(n6192), .A(n5710), .B(n5709), .ZN(U3027)
         );
  NOR2_X1 U6628 ( .A1(n6349), .A2(n5715), .ZN(n5733) );
  AOI22_X1 U6629 ( .A1(n5739), .A2(n6112), .B1(n6148), .B2(n5733), .ZN(n5719)
         );
  OAI21_X1 U6630 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6331), .A(n5921), 
        .ZN(n6014) );
  INV_X1 U6631 ( .A(n6014), .ZN(n6156) );
  INV_X1 U6632 ( .A(n5948), .ZN(n6347) );
  AOI21_X1 U6633 ( .B1(n5711), .B2(n6347), .A(n5733), .ZN(n5716) );
  AOI21_X1 U6634 ( .B1(n5712), .B2(STATEBS16_REG_SCAN_IN), .A(n6370), .ZN(
        n5714) );
  AOI22_X1 U6635 ( .A1(n5716), .A2(n5714), .B1(n6370), .B2(n5715), .ZN(n5713)
         );
  NAND2_X1 U6636 ( .A1(n6156), .A2(n5713), .ZN(n5736) );
  INV_X1 U6637 ( .A(n5714), .ZN(n5717) );
  OAI22_X1 U6638 ( .A1(n5717), .A2(n5716), .B1(n3558), .B2(n5715), .ZN(n5735)
         );
  AOI22_X1 U6639 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5736), .B1(n6149), 
        .B2(n5735), .ZN(n5718) );
  OAI211_X1 U6640 ( .C1(n6115), .C2(n5732), .A(n5719), .B(n5718), .ZN(U3028)
         );
  AOI22_X1 U6641 ( .A1(n5739), .A2(n6116), .B1(n6162), .B2(n5733), .ZN(n5721)
         );
  AOI22_X1 U6642 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5736), .B1(n6163), 
        .B2(n5735), .ZN(n5720) );
  OAI211_X1 U6643 ( .C1(n6119), .C2(n5732), .A(n5721), .B(n5720), .ZN(U3029)
         );
  INV_X1 U6644 ( .A(n6120), .ZN(n6173) );
  AOI22_X1 U6645 ( .A1(n5734), .A2(n6170), .B1(n6168), .B2(n5733), .ZN(n5723)
         );
  AOI22_X1 U6646 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5736), .B1(n6169), 
        .B2(n5735), .ZN(n5722) );
  OAI211_X1 U6647 ( .C1(n5761), .C2(n6173), .A(n5723), .B(n5722), .ZN(U3030)
         );
  INV_X1 U6648 ( .A(n6124), .ZN(n6179) );
  AOI22_X1 U6649 ( .A1(n5734), .A2(n6176), .B1(n6174), .B2(n5733), .ZN(n5725)
         );
  AOI22_X1 U6650 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5736), .B1(n6175), 
        .B2(n5735), .ZN(n5724) );
  OAI211_X1 U6651 ( .C1(n5761), .C2(n6179), .A(n5725), .B(n5724), .ZN(U3031)
         );
  INV_X1 U6652 ( .A(n6128), .ZN(n6185) );
  AOI22_X1 U6653 ( .A1(n5734), .A2(n6182), .B1(n6180), .B2(n5733), .ZN(n5727)
         );
  AOI22_X1 U6654 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5736), .B1(n6181), 
        .B2(n5735), .ZN(n5726) );
  OAI211_X1 U6655 ( .C1(n5761), .C2(n6185), .A(n5727), .B(n5726), .ZN(U3032)
         );
  INV_X1 U6656 ( .A(n6132), .ZN(n6193) );
  AOI22_X1 U6657 ( .A1(n5734), .A2(n6189), .B1(n6186), .B2(n5733), .ZN(n5729)
         );
  AOI22_X1 U6658 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5736), .B1(n6187), 
        .B2(n5735), .ZN(n5728) );
  OAI211_X1 U6659 ( .C1(n5761), .C2(n6193), .A(n5729), .B(n5728), .ZN(U3033)
         );
  AOI22_X1 U6660 ( .A1(n5739), .A2(n6196), .B1(n6195), .B2(n5733), .ZN(n5731)
         );
  AOI22_X1 U6661 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5736), .B1(n6194), 
        .B2(n5735), .ZN(n5730) );
  OAI211_X1 U6662 ( .C1(n6199), .C2(n5732), .A(n5731), .B(n5730), .ZN(U3034)
         );
  INV_X1 U6663 ( .A(n6205), .ZN(n5912) );
  INV_X1 U6664 ( .A(n6210), .ZN(n5905) );
  AOI22_X1 U6665 ( .A1(n5734), .A2(n5905), .B1(n6200), .B2(n5733), .ZN(n5738)
         );
  AOI22_X1 U6666 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5736), .B1(n6203), 
        .B2(n5735), .ZN(n5737) );
  OAI211_X1 U6667 ( .C1(n5761), .C2(n5912), .A(n5738), .B(n5737), .ZN(U3035)
         );
  AND2_X1 U6668 ( .A1(n2965), .A2(n5797), .ZN(n5982) );
  NAND2_X1 U6669 ( .A1(n6103), .A2(n5982), .ZN(n5767) );
  NAND2_X1 U6670 ( .A1(n6105), .A2(n5914), .ZN(n5986) );
  OAI22_X1 U6671 ( .A1(n5767), .A2(n6370), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n5986), .ZN(n5757) );
  NAND3_X1 U6672 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n3479), .A3(n6213), .ZN(n5772) );
  NOR2_X1 U6673 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5772), .ZN(n5756)
         );
  AOI22_X1 U6674 ( .A1(n6149), .A2(n5757), .B1(n6148), .B2(n5756), .ZN(n5743)
         );
  NAND2_X1 U6675 ( .A1(n5917), .A2(n6071), .ZN(n5979) );
  OAI21_X1 U6676 ( .B1(n5739), .B2(n5791), .A(n6151), .ZN(n5740) );
  NAND2_X1 U6677 ( .A1(n5740), .A2(n5767), .ZN(n5741) );
  OAI21_X1 U6678 ( .B1(n5914), .B2(n3558), .A(n5921), .ZN(n6106) );
  NOR2_X1 U6679 ( .A1(n5923), .A2(n6106), .ZN(n5984) );
  AOI22_X1 U6680 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n5758), .B1(n6112), 
        .B2(n5791), .ZN(n5742) );
  OAI211_X1 U6681 ( .C1(n6115), .C2(n5761), .A(n5743), .B(n5742), .ZN(U3036)
         );
  AOI22_X1 U6682 ( .A1(n6163), .A2(n5757), .B1(n6162), .B2(n5756), .ZN(n5745)
         );
  AOI22_X1 U6683 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n5758), .B1(n5791), 
        .B2(n6116), .ZN(n5744) );
  OAI211_X1 U6684 ( .C1(n5761), .C2(n6119), .A(n5745), .B(n5744), .ZN(U3037)
         );
  AOI22_X1 U6685 ( .A1(n6169), .A2(n5757), .B1(n6168), .B2(n5756), .ZN(n5747)
         );
  AOI22_X1 U6686 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(n5758), .B1(n5791), 
        .B2(n6120), .ZN(n5746) );
  OAI211_X1 U6687 ( .C1(n5761), .C2(n6123), .A(n5747), .B(n5746), .ZN(U3038)
         );
  AOI22_X1 U6688 ( .A1(n6175), .A2(n5757), .B1(n6174), .B2(n5756), .ZN(n5749)
         );
  AOI22_X1 U6689 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(n5758), .B1(n5791), 
        .B2(n6124), .ZN(n5748) );
  OAI211_X1 U6690 ( .C1(n5761), .C2(n6127), .A(n5749), .B(n5748), .ZN(U3039)
         );
  AOI22_X1 U6691 ( .A1(n6181), .A2(n5757), .B1(n6180), .B2(n5756), .ZN(n5751)
         );
  AOI22_X1 U6692 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n5758), .B1(n5791), 
        .B2(n6128), .ZN(n5750) );
  OAI211_X1 U6693 ( .C1(n5761), .C2(n6131), .A(n5751), .B(n5750), .ZN(U3040)
         );
  AOI22_X1 U6694 ( .A1(n6187), .A2(n5757), .B1(n6186), .B2(n5756), .ZN(n5753)
         );
  AOI22_X1 U6695 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n5758), .B1(n5791), 
        .B2(n6132), .ZN(n5752) );
  OAI211_X1 U6696 ( .C1(n5761), .C2(n6135), .A(n5753), .B(n5752), .ZN(U3041)
         );
  AOI22_X1 U6697 ( .A1(n6195), .A2(n5756), .B1(n6194), .B2(n5757), .ZN(n5755)
         );
  AOI22_X1 U6698 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n5758), .B1(n5791), 
        .B2(n6196), .ZN(n5754) );
  OAI211_X1 U6699 ( .C1(n5761), .C2(n6199), .A(n5755), .B(n5754), .ZN(U3042)
         );
  AOI22_X1 U6700 ( .A1(n6203), .A2(n5757), .B1(n6200), .B2(n5756), .ZN(n5760)
         );
  AOI22_X1 U6701 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n5758), .B1(n5791), 
        .B2(n6205), .ZN(n5759) );
  OAI211_X1 U6702 ( .C1(n5761), .C2(n6210), .A(n5760), .B(n5759), .ZN(U3043)
         );
  NOR2_X1 U6703 ( .A1(n6010), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5792)
         );
  NAND2_X1 U6704 ( .A1(n5917), .A2(n6344), .ZN(n6009) );
  INV_X1 U6705 ( .A(n5824), .ZN(n5787) );
  AOI22_X1 U6706 ( .A1(n6148), .A2(n5792), .B1(n5787), .B2(n6112), .ZN(n5776)
         );
  INV_X1 U6707 ( .A(n6011), .ZN(n5763) );
  NAND2_X1 U6708 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  OAI21_X1 U6709 ( .B1(n5766), .B2(n5765), .A(n6345), .ZN(n5773) );
  OR2_X1 U6710 ( .A1(n5767), .A2(n5948), .ZN(n5769) );
  INV_X1 U6711 ( .A(n5792), .ZN(n5768) );
  AND2_X1 U6712 ( .A1(n5769), .A2(n5768), .ZN(n5774) );
  INV_X1 U6713 ( .A(n5774), .ZN(n5771) );
  AOI21_X1 U6714 ( .B1(n6370), .B2(n5772), .A(n6014), .ZN(n5770) );
  OAI21_X1 U6715 ( .B1(n5773), .B2(n5771), .A(n5770), .ZN(n5794) );
  OAI22_X1 U6716 ( .A1(n5774), .A2(n5773), .B1(n3558), .B2(n5772), .ZN(n5793)
         );
  AOI22_X1 U6717 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5794), .B1(n6149), 
        .B2(n5793), .ZN(n5775) );
  OAI211_X1 U6718 ( .C1(n6115), .C2(n5790), .A(n5776), .B(n5775), .ZN(U3044)
         );
  INV_X1 U6719 ( .A(n6116), .ZN(n6167) );
  AOI22_X1 U6720 ( .A1(n6162), .A2(n5792), .B1(n5791), .B2(n6164), .ZN(n5778)
         );
  AOI22_X1 U6721 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5794), .B1(n6163), 
        .B2(n5793), .ZN(n5777) );
  OAI211_X1 U6722 ( .C1(n6167), .C2(n5824), .A(n5778), .B(n5777), .ZN(U3045)
         );
  AOI22_X1 U6723 ( .A1(n6168), .A2(n5792), .B1(n5787), .B2(n6120), .ZN(n5780)
         );
  AOI22_X1 U6724 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5794), .B1(n6169), 
        .B2(n5793), .ZN(n5779) );
  OAI211_X1 U6725 ( .C1(n5790), .C2(n6123), .A(n5780), .B(n5779), .ZN(U3046)
         );
  AOI22_X1 U6726 ( .A1(n6174), .A2(n5792), .B1(n5791), .B2(n6176), .ZN(n5782)
         );
  AOI22_X1 U6727 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n5794), .B1(n6175), 
        .B2(n5793), .ZN(n5781) );
  OAI211_X1 U6728 ( .C1(n6179), .C2(n5824), .A(n5782), .B(n5781), .ZN(U3047)
         );
  AOI22_X1 U6729 ( .A1(n6180), .A2(n5792), .B1(n5791), .B2(n6182), .ZN(n5784)
         );
  AOI22_X1 U6730 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5794), .B1(n6181), 
        .B2(n5793), .ZN(n5783) );
  OAI211_X1 U6731 ( .C1(n6185), .C2(n5824), .A(n5784), .B(n5783), .ZN(U3048)
         );
  AOI22_X1 U6732 ( .A1(n6186), .A2(n5792), .B1(n5787), .B2(n6132), .ZN(n5786)
         );
  AOI22_X1 U6733 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5794), .B1(n6187), 
        .B2(n5793), .ZN(n5785) );
  OAI211_X1 U6734 ( .C1(n5790), .C2(n6135), .A(n5786), .B(n5785), .ZN(U3049)
         );
  AOI22_X1 U6735 ( .A1(n6195), .A2(n5792), .B1(n5787), .B2(n6196), .ZN(n5789)
         );
  AOI22_X1 U6736 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5794), .B1(n6194), 
        .B2(n5793), .ZN(n5788) );
  OAI211_X1 U6737 ( .C1(n5790), .C2(n6199), .A(n5789), .B(n5788), .ZN(U3050)
         );
  AOI22_X1 U6738 ( .A1(n6200), .A2(n5792), .B1(n5791), .B2(n5905), .ZN(n5796)
         );
  AOI22_X1 U6739 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5794), .B1(n6203), 
        .B2(n5793), .ZN(n5795) );
  OAI211_X1 U6740 ( .C1(n5912), .C2(n5824), .A(n5796), .B(n5795), .ZN(U3051)
         );
  INV_X1 U6741 ( .A(n5923), .ZN(n6041) );
  NOR2_X1 U6742 ( .A1(n2965), .A2(n5797), .ZN(n6073) );
  NAND3_X1 U6743 ( .A1(n6103), .A2(n6345), .A3(n6073), .ZN(n5798) );
  OAI21_X1 U6744 ( .B1(n5799), .B2(n6041), .A(n5798), .ZN(n5820) );
  NAND2_X1 U6745 ( .A1(n6218), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6078) );
  OR2_X1 U6746 ( .A1(n6078), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5831)
         );
  NOR2_X1 U6747 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5831), .ZN(n5819)
         );
  AOI22_X1 U6748 ( .A1(n6149), .A2(n5820), .B1(n6148), .B2(n5819), .ZN(n5806)
         );
  AOI21_X1 U6749 ( .B1(n5854), .B2(n5824), .A(n6363), .ZN(n5800) );
  AOI211_X1 U6750 ( .C1(n5801), .C2(n6073), .A(n6370), .B(n5800), .ZN(n5803)
         );
  NOR3_X1 U6751 ( .A1(n5803), .A2(n6105), .A3(n5802), .ZN(n5804) );
  AOI22_X1 U6752 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n5821), .B1(n6112), 
        .B2(n5844), .ZN(n5805) );
  OAI211_X1 U6753 ( .C1(n6115), .C2(n5824), .A(n5806), .B(n5805), .ZN(U3052)
         );
  AOI22_X1 U6754 ( .A1(n6163), .A2(n5820), .B1(n6162), .B2(n5819), .ZN(n5808)
         );
  AOI22_X1 U6755 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n5821), .B1(n6116), 
        .B2(n5844), .ZN(n5807) );
  OAI211_X1 U6756 ( .C1(n6119), .C2(n5824), .A(n5808), .B(n5807), .ZN(U3053)
         );
  AOI22_X1 U6757 ( .A1(n6169), .A2(n5820), .B1(n6168), .B2(n5819), .ZN(n5810)
         );
  AOI22_X1 U6758 ( .A1(INSTQUEUE_REG_4__2__SCAN_IN), .A2(n5821), .B1(n6120), 
        .B2(n5844), .ZN(n5809) );
  OAI211_X1 U6759 ( .C1(n6123), .C2(n5824), .A(n5810), .B(n5809), .ZN(U3054)
         );
  AOI22_X1 U6760 ( .A1(n6175), .A2(n5820), .B1(n6174), .B2(n5819), .ZN(n5812)
         );
  AOI22_X1 U6761 ( .A1(INSTQUEUE_REG_4__3__SCAN_IN), .A2(n5821), .B1(n6124), 
        .B2(n5844), .ZN(n5811) );
  OAI211_X1 U6762 ( .C1(n6127), .C2(n5824), .A(n5812), .B(n5811), .ZN(U3055)
         );
  AOI22_X1 U6763 ( .A1(n6181), .A2(n5820), .B1(n6180), .B2(n5819), .ZN(n5814)
         );
  AOI22_X1 U6764 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n5821), .B1(n6128), 
        .B2(n5844), .ZN(n5813) );
  OAI211_X1 U6765 ( .C1(n6131), .C2(n5824), .A(n5814), .B(n5813), .ZN(U3056)
         );
  AOI22_X1 U6766 ( .A1(n6187), .A2(n5820), .B1(n6186), .B2(n5819), .ZN(n5816)
         );
  AOI22_X1 U6767 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n5821), .B1(n6132), 
        .B2(n5844), .ZN(n5815) );
  OAI211_X1 U6768 ( .C1(n6135), .C2(n5824), .A(n5816), .B(n5815), .ZN(U3057)
         );
  AOI22_X1 U6769 ( .A1(n6195), .A2(n5819), .B1(n6194), .B2(n5820), .ZN(n5818)
         );
  AOI22_X1 U6770 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(n5821), .B1(n6196), 
        .B2(n5844), .ZN(n5817) );
  OAI211_X1 U6771 ( .C1(n6199), .C2(n5824), .A(n5818), .B(n5817), .ZN(U3058)
         );
  AOI22_X1 U6772 ( .A1(n6203), .A2(n5820), .B1(n6200), .B2(n5819), .ZN(n5823)
         );
  AOI22_X1 U6773 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n5821), .B1(n6205), 
        .B2(n5844), .ZN(n5822) );
  OAI211_X1 U6774 ( .C1(n6210), .C2(n5824), .A(n5823), .B(n5822), .ZN(U3059)
         );
  NOR2_X1 U6775 ( .A1(n6349), .A2(n5831), .ZN(n5849) );
  AOI22_X1 U6776 ( .A1(n5856), .A2(n6112), .B1(n6148), .B2(n5849), .ZN(n5835)
         );
  OAI21_X1 U6777 ( .B1(n5825), .B2(n6363), .A(n6345), .ZN(n5832) );
  NOR2_X1 U6778 ( .A1(n5948), .A2(n5826), .ZN(n5884) );
  NAND2_X1 U6779 ( .A1(n6073), .A2(n5884), .ZN(n5828) );
  INV_X1 U6780 ( .A(n5849), .ZN(n5827) );
  AND2_X1 U6781 ( .A1(n5828), .A2(n5827), .ZN(n5833) );
  INV_X1 U6782 ( .A(n5833), .ZN(n5830) );
  AOI21_X1 U6783 ( .B1(n6370), .B2(n5831), .A(n6014), .ZN(n5829) );
  OAI21_X1 U6784 ( .B1(n5832), .B2(n5830), .A(n5829), .ZN(n5851) );
  OAI22_X1 U6785 ( .A1(n5833), .A2(n5832), .B1(n3558), .B2(n5831), .ZN(n5850)
         );
  AOI22_X1 U6786 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5851), .B1(n6149), 
        .B2(n5850), .ZN(n5834) );
  OAI211_X1 U6787 ( .C1(n6115), .C2(n5854), .A(n5835), .B(n5834), .ZN(U3060)
         );
  AOI22_X1 U6788 ( .A1(n5856), .A2(n6116), .B1(n6162), .B2(n5849), .ZN(n5837)
         );
  AOI22_X1 U6789 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5851), .B1(n6163), 
        .B2(n5850), .ZN(n5836) );
  OAI211_X1 U6790 ( .C1(n6119), .C2(n5854), .A(n5837), .B(n5836), .ZN(U3061)
         );
  AOI22_X1 U6791 ( .A1(n5844), .A2(n6170), .B1(n6168), .B2(n5849), .ZN(n5839)
         );
  AOI22_X1 U6792 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5851), .B1(n6169), 
        .B2(n5850), .ZN(n5838) );
  OAI211_X1 U6793 ( .C1(n6173), .C2(n5880), .A(n5839), .B(n5838), .ZN(U3062)
         );
  AOI22_X1 U6794 ( .A1(n5844), .A2(n6176), .B1(n6174), .B2(n5849), .ZN(n5841)
         );
  AOI22_X1 U6795 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5851), .B1(n6175), 
        .B2(n5850), .ZN(n5840) );
  OAI211_X1 U6796 ( .C1(n6179), .C2(n5880), .A(n5841), .B(n5840), .ZN(U3063)
         );
  AOI22_X1 U6797 ( .A1(n5844), .A2(n6182), .B1(n6180), .B2(n5849), .ZN(n5843)
         );
  AOI22_X1 U6798 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5851), .B1(n6181), 
        .B2(n5850), .ZN(n5842) );
  OAI211_X1 U6799 ( .C1(n6185), .C2(n5880), .A(n5843), .B(n5842), .ZN(U3064)
         );
  AOI22_X1 U6800 ( .A1(n5844), .A2(n6189), .B1(n6186), .B2(n5849), .ZN(n5846)
         );
  AOI22_X1 U6801 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5851), .B1(n6187), 
        .B2(n5850), .ZN(n5845) );
  OAI211_X1 U6802 ( .C1(n6193), .C2(n5880), .A(n5846), .B(n5845), .ZN(U3065)
         );
  AOI22_X1 U6803 ( .A1(n5856), .A2(n6196), .B1(n6195), .B2(n5849), .ZN(n5848)
         );
  AOI22_X1 U6804 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5851), .B1(n6194), 
        .B2(n5850), .ZN(n5847) );
  OAI211_X1 U6805 ( .C1(n6199), .C2(n5854), .A(n5848), .B(n5847), .ZN(U3066)
         );
  AOI22_X1 U6806 ( .A1(n5856), .A2(n6205), .B1(n6200), .B2(n5849), .ZN(n5853)
         );
  AOI22_X1 U6807 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5851), .B1(n6203), 
        .B2(n5850), .ZN(n5852) );
  OAI211_X1 U6808 ( .C1(n6210), .C2(n5854), .A(n5853), .B(n5852), .ZN(U3067)
         );
  OR2_X1 U6809 ( .A1(n2965), .A2(n5855), .ZN(n6109) );
  NAND2_X1 U6810 ( .A1(n6145), .A2(n6345), .ZN(n6104) );
  NAND2_X1 U6811 ( .A1(n5923), .A2(n5914), .ZN(n6102) );
  OAI22_X1 U6812 ( .A1(n6104), .A2(n4264), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6102), .ZN(n5876) );
  NOR2_X1 U6813 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5887), .ZN(n5875)
         );
  AOI22_X1 U6814 ( .A1(n6149), .A2(n5876), .B1(n6148), .B2(n5875), .ZN(n5862)
         );
  OAI21_X1 U6815 ( .B1(n5856), .B2(n5906), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5857) );
  NAND3_X1 U6816 ( .A1(n6109), .A2(n6345), .A3(n5857), .ZN(n5860) );
  INV_X1 U6817 ( .A(n5875), .ZN(n5858) );
  AOI211_X1 U6818 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5858), .A(n6105), .B(
        n6106), .ZN(n5859) );
  NAND3_X1 U6819 ( .A1(n3479), .A2(n5860), .A3(n5859), .ZN(n5877) );
  AOI22_X1 U6820 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n5877), .B1(n6112), 
        .B2(n5906), .ZN(n5861) );
  OAI211_X1 U6821 ( .C1(n6115), .C2(n5880), .A(n5862), .B(n5861), .ZN(U3068)
         );
  AOI22_X1 U6822 ( .A1(n6163), .A2(n5876), .B1(n6162), .B2(n5875), .ZN(n5864)
         );
  AOI22_X1 U6823 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n5877), .B1(n6116), 
        .B2(n5906), .ZN(n5863) );
  OAI211_X1 U6824 ( .C1(n6119), .C2(n5880), .A(n5864), .B(n5863), .ZN(U3069)
         );
  AOI22_X1 U6825 ( .A1(n6169), .A2(n5876), .B1(n6168), .B2(n5875), .ZN(n5866)
         );
  AOI22_X1 U6826 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n5877), .B1(n6120), 
        .B2(n5906), .ZN(n5865) );
  OAI211_X1 U6827 ( .C1(n6123), .C2(n5880), .A(n5866), .B(n5865), .ZN(U3070)
         );
  AOI22_X1 U6828 ( .A1(n6175), .A2(n5876), .B1(n6174), .B2(n5875), .ZN(n5868)
         );
  AOI22_X1 U6829 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n5877), .B1(n6124), 
        .B2(n5906), .ZN(n5867) );
  OAI211_X1 U6830 ( .C1(n6127), .C2(n5880), .A(n5868), .B(n5867), .ZN(U3071)
         );
  AOI22_X1 U6831 ( .A1(n6181), .A2(n5876), .B1(n6180), .B2(n5875), .ZN(n5870)
         );
  AOI22_X1 U6832 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n5877), .B1(n6128), 
        .B2(n5906), .ZN(n5869) );
  OAI211_X1 U6833 ( .C1(n6131), .C2(n5880), .A(n5870), .B(n5869), .ZN(U3072)
         );
  AOI22_X1 U6834 ( .A1(n6187), .A2(n5876), .B1(n6186), .B2(n5875), .ZN(n5872)
         );
  AOI22_X1 U6835 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n5877), .B1(n6132), 
        .B2(n5906), .ZN(n5871) );
  OAI211_X1 U6836 ( .C1(n6135), .C2(n5880), .A(n5872), .B(n5871), .ZN(U3073)
         );
  AOI22_X1 U6837 ( .A1(n6195), .A2(n5875), .B1(n6194), .B2(n5876), .ZN(n5874)
         );
  AOI22_X1 U6838 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n5877), .B1(n6196), 
        .B2(n5906), .ZN(n5873) );
  OAI211_X1 U6839 ( .C1(n6199), .C2(n5880), .A(n5874), .B(n5873), .ZN(U3074)
         );
  AOI22_X1 U6840 ( .A1(n6203), .A2(n5876), .B1(n6200), .B2(n5875), .ZN(n5879)
         );
  AOI22_X1 U6841 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n5877), .B1(n6205), 
        .B2(n5906), .ZN(n5878) );
  OAI211_X1 U6842 ( .C1(n6210), .C2(n5880), .A(n5879), .B(n5878), .ZN(U3075)
         );
  INV_X1 U6843 ( .A(n5881), .ZN(n5907) );
  AOI22_X1 U6844 ( .A1(n6148), .A2(n5907), .B1(n5918), .B2(n6112), .ZN(n5891)
         );
  NOR2_X1 U6845 ( .A1(n5883), .A2(n6370), .ZN(n5886) );
  AOI21_X1 U6846 ( .B1(n6145), .B2(n5884), .A(n5907), .ZN(n5889) );
  AOI22_X1 U6847 ( .A1(n5886), .A2(n5889), .B1(n6370), .B2(n5887), .ZN(n5885)
         );
  NAND2_X1 U6848 ( .A1(n6156), .A2(n5885), .ZN(n5909) );
  INV_X1 U6849 ( .A(n5886), .ZN(n5888) );
  OAI22_X1 U6850 ( .A1(n5889), .A2(n5888), .B1(n3558), .B2(n5887), .ZN(n5908)
         );
  AOI22_X1 U6851 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5909), .B1(n6149), 
        .B2(n5908), .ZN(n5890) );
  OAI211_X1 U6852 ( .C1(n6115), .C2(n5904), .A(n5891), .B(n5890), .ZN(U3076)
         );
  AOI22_X1 U6853 ( .A1(n6162), .A2(n5907), .B1(n5906), .B2(n6164), .ZN(n5893)
         );
  AOI22_X1 U6854 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5909), .B1(n6163), 
        .B2(n5908), .ZN(n5892) );
  OAI211_X1 U6855 ( .C1(n6167), .C2(n5947), .A(n5893), .B(n5892), .ZN(U3077)
         );
  AOI22_X1 U6856 ( .A1(n6168), .A2(n5907), .B1(n5918), .B2(n6120), .ZN(n5895)
         );
  AOI22_X1 U6857 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5909), .B1(n6169), 
        .B2(n5908), .ZN(n5894) );
  OAI211_X1 U6858 ( .C1(n6123), .C2(n5904), .A(n5895), .B(n5894), .ZN(U3078)
         );
  AOI22_X1 U6859 ( .A1(n6174), .A2(n5907), .B1(n5918), .B2(n6124), .ZN(n5897)
         );
  AOI22_X1 U6860 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5909), .B1(n6175), 
        .B2(n5908), .ZN(n5896) );
  OAI211_X1 U6861 ( .C1(n6127), .C2(n5904), .A(n5897), .B(n5896), .ZN(U3079)
         );
  AOI22_X1 U6862 ( .A1(n6180), .A2(n5907), .B1(n5906), .B2(n6182), .ZN(n5899)
         );
  AOI22_X1 U6863 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5909), .B1(n6181), 
        .B2(n5908), .ZN(n5898) );
  OAI211_X1 U6864 ( .C1(n6185), .C2(n5947), .A(n5899), .B(n5898), .ZN(U3080)
         );
  AOI22_X1 U6865 ( .A1(n6186), .A2(n5907), .B1(n5918), .B2(n6132), .ZN(n5901)
         );
  AOI22_X1 U6866 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5909), .B1(n6187), 
        .B2(n5908), .ZN(n5900) );
  OAI211_X1 U6867 ( .C1(n6135), .C2(n5904), .A(n5901), .B(n5900), .ZN(U3081)
         );
  AOI22_X1 U6868 ( .A1(n6195), .A2(n5907), .B1(n5918), .B2(n6196), .ZN(n5903)
         );
  AOI22_X1 U6869 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5909), .B1(n6194), 
        .B2(n5908), .ZN(n5902) );
  OAI211_X1 U6870 ( .C1(n6199), .C2(n5904), .A(n5903), .B(n5902), .ZN(U3082)
         );
  AOI22_X1 U6871 ( .A1(n6200), .A2(n5907), .B1(n5906), .B2(n5905), .ZN(n5911)
         );
  AOI22_X1 U6872 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5909), .B1(n6203), 
        .B2(n5908), .ZN(n5910) );
  OAI211_X1 U6873 ( .C1(n5912), .C2(n5947), .A(n5911), .B(n5910), .ZN(U3083)
         );
  NOR2_X1 U6874 ( .A1(n6103), .A2(n5949), .ZN(n5926) );
  INV_X1 U6875 ( .A(n5926), .ZN(n5916) );
  INV_X1 U6876 ( .A(n5913), .ZN(n5915) );
  NOR2_X1 U6877 ( .A1(n5915), .A2(n5914), .ZN(n5922) );
  INV_X1 U6878 ( .A(n5922), .ZN(n6042) );
  OAI22_X1 U6879 ( .A1(n5916), .A2(n6370), .B1(n6049), .B2(n6042), .ZN(n5943)
         );
  NAND3_X1 U6880 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6213), .A3(n6218), .ZN(n5955) );
  NOR2_X1 U6881 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5955), .ZN(n5942)
         );
  AOI22_X1 U6882 ( .A1(n6149), .A2(n5943), .B1(n6148), .B2(n5942), .ZN(n5929)
         );
  NOR3_X1 U6883 ( .A1(n5968), .A2(n5918), .A3(n6370), .ZN(n5920) );
  NOR2_X1 U6884 ( .A1(n5920), .A2(n5919), .ZN(n5927) );
  INV_X1 U6885 ( .A(n5942), .ZN(n5924) );
  OAI21_X1 U6886 ( .B1(n5922), .B2(n3558), .A(n5921), .ZN(n6047) );
  AOI211_X1 U6887 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5924), .A(n5923), .B(
        n6047), .ZN(n5925) );
  AOI22_X1 U6888 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n5944), .B1(n6112), 
        .B2(n5968), .ZN(n5928) );
  OAI211_X1 U6889 ( .C1(n6115), .C2(n5947), .A(n5929), .B(n5928), .ZN(U3084)
         );
  AOI22_X1 U6890 ( .A1(n6163), .A2(n5943), .B1(n6162), .B2(n5942), .ZN(n5931)
         );
  AOI22_X1 U6891 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n5944), .B1(n6116), 
        .B2(n5968), .ZN(n5930) );
  OAI211_X1 U6892 ( .C1(n6119), .C2(n5947), .A(n5931), .B(n5930), .ZN(U3085)
         );
  AOI22_X1 U6893 ( .A1(n6169), .A2(n5943), .B1(n6168), .B2(n5942), .ZN(n5933)
         );
  AOI22_X1 U6894 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n5944), .B1(n6120), 
        .B2(n5968), .ZN(n5932) );
  OAI211_X1 U6895 ( .C1(n6123), .C2(n5947), .A(n5933), .B(n5932), .ZN(U3086)
         );
  AOI22_X1 U6896 ( .A1(n6175), .A2(n5943), .B1(n6174), .B2(n5942), .ZN(n5935)
         );
  AOI22_X1 U6897 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n5944), .B1(n6124), 
        .B2(n5968), .ZN(n5934) );
  OAI211_X1 U6898 ( .C1(n6127), .C2(n5947), .A(n5935), .B(n5934), .ZN(U3087)
         );
  AOI22_X1 U6899 ( .A1(n6181), .A2(n5943), .B1(n6180), .B2(n5942), .ZN(n5937)
         );
  AOI22_X1 U6900 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n5944), .B1(n6128), 
        .B2(n5968), .ZN(n5936) );
  OAI211_X1 U6901 ( .C1(n6131), .C2(n5947), .A(n5937), .B(n5936), .ZN(U3088)
         );
  AOI22_X1 U6902 ( .A1(n6187), .A2(n5943), .B1(n6186), .B2(n5942), .ZN(n5939)
         );
  AOI22_X1 U6903 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n5944), .B1(n6132), 
        .B2(n5968), .ZN(n5938) );
  OAI211_X1 U6904 ( .C1(n6135), .C2(n5947), .A(n5939), .B(n5938), .ZN(U3089)
         );
  AOI22_X1 U6905 ( .A1(n6195), .A2(n5942), .B1(n6194), .B2(n5943), .ZN(n5941)
         );
  AOI22_X1 U6906 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n5944), .B1(n6196), 
        .B2(n5968), .ZN(n5940) );
  OAI211_X1 U6907 ( .C1(n6199), .C2(n5947), .A(n5941), .B(n5940), .ZN(U3090)
         );
  AOI22_X1 U6908 ( .A1(n6203), .A2(n5943), .B1(n6200), .B2(n5942), .ZN(n5946)
         );
  AOI22_X1 U6909 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n5944), .B1(n6205), 
        .B2(n5968), .ZN(n5945) );
  OAI211_X1 U6910 ( .C1(n6210), .C2(n5947), .A(n5946), .B(n5945), .ZN(U3091)
         );
  NOR2_X1 U6911 ( .A1(n6349), .A2(n5955), .ZN(n5973) );
  AOI22_X1 U6912 ( .A1(n5980), .A2(n6112), .B1(n5973), .B2(n6148), .ZN(n5959)
         );
  NOR2_X1 U6913 ( .A1(n6103), .A2(n5948), .ZN(n6146) );
  INV_X1 U6914 ( .A(n5949), .ZN(n5950) );
  AOI21_X1 U6915 ( .B1(n6146), .B2(n5950), .A(n5973), .ZN(n5957) );
  OR2_X1 U6916 ( .A1(n5951), .A2(n6363), .ZN(n5952) );
  AOI22_X1 U6917 ( .A1(n5957), .A2(n5954), .B1(n6370), .B2(n5955), .ZN(n5953)
         );
  NAND2_X1 U6918 ( .A1(n6156), .A2(n5953), .ZN(n5975) );
  INV_X1 U6919 ( .A(n5954), .ZN(n5956) );
  OAI22_X1 U6920 ( .A1(n5957), .A2(n5956), .B1(n3558), .B2(n5955), .ZN(n5974)
         );
  AOI22_X1 U6921 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5975), .B1(n6149), 
        .B2(n5974), .ZN(n5958) );
  OAI211_X1 U6922 ( .C1(n6115), .C2(n5978), .A(n5959), .B(n5958), .ZN(U3092)
         );
  AOI22_X1 U6923 ( .A1(n5968), .A2(n6164), .B1(n5973), .B2(n6162), .ZN(n5961)
         );
  AOI22_X1 U6924 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5975), .B1(n6163), 
        .B2(n5974), .ZN(n5960) );
  OAI211_X1 U6925 ( .C1(n6167), .C2(n6008), .A(n5961), .B(n5960), .ZN(U3093)
         );
  AOI22_X1 U6926 ( .A1(n5980), .A2(n6120), .B1(n5973), .B2(n6168), .ZN(n5963)
         );
  AOI22_X1 U6927 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5975), .B1(n6169), 
        .B2(n5974), .ZN(n5962) );
  OAI211_X1 U6928 ( .C1(n6123), .C2(n5978), .A(n5963), .B(n5962), .ZN(U3094)
         );
  AOI22_X1 U6929 ( .A1(n5968), .A2(n6176), .B1(n5973), .B2(n6174), .ZN(n5965)
         );
  AOI22_X1 U6930 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5975), .B1(n6175), 
        .B2(n5974), .ZN(n5964) );
  OAI211_X1 U6931 ( .C1(n6179), .C2(n6008), .A(n5965), .B(n5964), .ZN(U3095)
         );
  AOI22_X1 U6932 ( .A1(n5968), .A2(n6182), .B1(n5973), .B2(n6180), .ZN(n5967)
         );
  AOI22_X1 U6933 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5975), .B1(n6181), 
        .B2(n5974), .ZN(n5966) );
  OAI211_X1 U6934 ( .C1(n6185), .C2(n6008), .A(n5967), .B(n5966), .ZN(U3096)
         );
  AOI22_X1 U6935 ( .A1(n5968), .A2(n6189), .B1(n5973), .B2(n6186), .ZN(n5970)
         );
  AOI22_X1 U6936 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5975), .B1(n6187), 
        .B2(n5974), .ZN(n5969) );
  OAI211_X1 U6937 ( .C1(n6193), .C2(n6008), .A(n5970), .B(n5969), .ZN(U3097)
         );
  AOI22_X1 U6938 ( .A1(n5980), .A2(n6196), .B1(n5973), .B2(n6195), .ZN(n5972)
         );
  AOI22_X1 U6939 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5975), .B1(n6194), 
        .B2(n5974), .ZN(n5971) );
  OAI211_X1 U6940 ( .C1(n6199), .C2(n5978), .A(n5972), .B(n5971), .ZN(U3098)
         );
  AOI22_X1 U6941 ( .A1(n5980), .A2(n6205), .B1(n5973), .B2(n6200), .ZN(n5977)
         );
  AOI22_X1 U6942 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5975), .B1(n6203), 
        .B2(n5974), .ZN(n5976) );
  OAI211_X1 U6943 ( .C1(n6210), .C2(n5978), .A(n5977), .B(n5976), .ZN(U3099)
         );
  NAND3_X1 U6944 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6213), .ZN(n6017) );
  NOR2_X1 U6945 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6017), .ZN(n6003)
         );
  AOI22_X1 U6946 ( .A1(n6148), .A2(n6003), .B1(n6030), .B2(n6112), .ZN(n5990)
         );
  OAI21_X1 U6947 ( .B1(n5980), .B2(n6030), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5981) );
  NAND2_X1 U6948 ( .A1(n5981), .A2(n6345), .ZN(n5988) );
  INV_X1 U6949 ( .A(n6003), .ZN(n5983) );
  AOI22_X1 U6950 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n3479), .B1(
        STATE2_REG_3__SCAN_IN), .B2(n5983), .ZN(n5985) );
  OAI211_X1 U6951 ( .C1(n5988), .C2(n6013), .A(n5985), .B(n5984), .ZN(n6005)
         );
  INV_X1 U6952 ( .A(n6013), .ZN(n5987) );
  OAI22_X1 U6953 ( .A1(n5988), .A2(n5987), .B1(n3479), .B2(n5986), .ZN(n6004)
         );
  AOI22_X1 U6954 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6005), .B1(n6149), 
        .B2(n6004), .ZN(n5989) );
  OAI211_X1 U6955 ( .C1(n6115), .C2(n6008), .A(n5990), .B(n5989), .ZN(U3100)
         );
  AOI22_X1 U6956 ( .A1(n6162), .A2(n6003), .B1(n6030), .B2(n6116), .ZN(n5992)
         );
  AOI22_X1 U6957 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6005), .B1(n6163), 
        .B2(n6004), .ZN(n5991) );
  OAI211_X1 U6958 ( .C1(n6119), .C2(n6008), .A(n5992), .B(n5991), .ZN(U3101)
         );
  AOI22_X1 U6959 ( .A1(n6168), .A2(n6003), .B1(n6030), .B2(n6120), .ZN(n5994)
         );
  AOI22_X1 U6960 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6005), .B1(n6169), 
        .B2(n6004), .ZN(n5993) );
  OAI211_X1 U6961 ( .C1(n6123), .C2(n6008), .A(n5994), .B(n5993), .ZN(U3102)
         );
  AOI22_X1 U6962 ( .A1(n6174), .A2(n6003), .B1(n6030), .B2(n6124), .ZN(n5996)
         );
  AOI22_X1 U6963 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6005), .B1(n6175), 
        .B2(n6004), .ZN(n5995) );
  OAI211_X1 U6964 ( .C1(n6127), .C2(n6008), .A(n5996), .B(n5995), .ZN(U3103)
         );
  AOI22_X1 U6965 ( .A1(n6180), .A2(n6003), .B1(n6030), .B2(n6128), .ZN(n5998)
         );
  AOI22_X1 U6966 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6005), .B1(n6181), 
        .B2(n6004), .ZN(n5997) );
  OAI211_X1 U6967 ( .C1(n6131), .C2(n6008), .A(n5998), .B(n5997), .ZN(U3104)
         );
  AOI22_X1 U6968 ( .A1(n6186), .A2(n6003), .B1(n6030), .B2(n6132), .ZN(n6000)
         );
  AOI22_X1 U6969 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6005), .B1(n6187), 
        .B2(n6004), .ZN(n5999) );
  OAI211_X1 U6970 ( .C1(n6135), .C2(n6008), .A(n6000), .B(n5999), .ZN(U3105)
         );
  AOI22_X1 U6971 ( .A1(n6195), .A2(n6003), .B1(n6030), .B2(n6196), .ZN(n6002)
         );
  AOI22_X1 U6972 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6005), .B1(n6194), 
        .B2(n6004), .ZN(n6001) );
  OAI211_X1 U6973 ( .C1(n6199), .C2(n6008), .A(n6002), .B(n6001), .ZN(U3106)
         );
  AOI22_X1 U6974 ( .A1(n6200), .A2(n6003), .B1(n6030), .B2(n6205), .ZN(n6007)
         );
  AOI22_X1 U6975 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6005), .B1(n6203), 
        .B2(n6004), .ZN(n6006) );
  OAI211_X1 U6976 ( .C1(n6210), .C2(n6008), .A(n6007), .B(n6006), .ZN(U3107)
         );
  INV_X1 U6977 ( .A(n6112), .ZN(n6161) );
  NOR2_X1 U6978 ( .A1(n6010), .A2(n3479), .ZN(n6035) );
  AOI22_X1 U6979 ( .A1(n6148), .A2(n6035), .B1(n6030), .B2(n6158), .ZN(n6021)
         );
  OAI21_X1 U6980 ( .B1(n6012), .B2(n6011), .A(n6345), .ZN(n6019) );
  AOI21_X1 U6981 ( .B1(n6013), .B2(n6347), .A(n6035), .ZN(n6018) );
  INV_X1 U6982 ( .A(n6018), .ZN(n6016) );
  AOI21_X1 U6983 ( .B1(n6370), .B2(n6017), .A(n6014), .ZN(n6015) );
  OAI21_X1 U6984 ( .B1(n6019), .B2(n6016), .A(n6015), .ZN(n6037) );
  OAI22_X1 U6985 ( .A1(n6019), .A2(n6018), .B1(n6017), .B2(n3558), .ZN(n6036)
         );
  AOI22_X1 U6986 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6037), .B1(n6149), 
        .B2(n6036), .ZN(n6020) );
  OAI211_X1 U6987 ( .C1(n6161), .C2(n6070), .A(n6021), .B(n6020), .ZN(U3108)
         );
  AOI22_X1 U6988 ( .A1(n6162), .A2(n6035), .B1(n6043), .B2(n6116), .ZN(n6023)
         );
  AOI22_X1 U6989 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6037), .B1(n6163), 
        .B2(n6036), .ZN(n6022) );
  OAI211_X1 U6990 ( .C1(n6119), .C2(n6040), .A(n6023), .B(n6022), .ZN(U3109)
         );
  AOI22_X1 U6991 ( .A1(n6168), .A2(n6035), .B1(n6043), .B2(n6120), .ZN(n6025)
         );
  AOI22_X1 U6992 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6037), .B1(n6169), 
        .B2(n6036), .ZN(n6024) );
  OAI211_X1 U6993 ( .C1(n6123), .C2(n6040), .A(n6025), .B(n6024), .ZN(U3110)
         );
  AOI22_X1 U6994 ( .A1(n6174), .A2(n6035), .B1(n6030), .B2(n6176), .ZN(n6027)
         );
  AOI22_X1 U6995 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6037), .B1(n6175), 
        .B2(n6036), .ZN(n6026) );
  OAI211_X1 U6996 ( .C1(n6179), .C2(n6070), .A(n6027), .B(n6026), .ZN(U3111)
         );
  AOI22_X1 U6997 ( .A1(n6180), .A2(n6035), .B1(n6043), .B2(n6128), .ZN(n6029)
         );
  AOI22_X1 U6998 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6037), .B1(n6181), 
        .B2(n6036), .ZN(n6028) );
  OAI211_X1 U6999 ( .C1(n6131), .C2(n6040), .A(n6029), .B(n6028), .ZN(U3112)
         );
  AOI22_X1 U7000 ( .A1(n6186), .A2(n6035), .B1(n6030), .B2(n6189), .ZN(n6032)
         );
  AOI22_X1 U7001 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6037), .B1(n6187), 
        .B2(n6036), .ZN(n6031) );
  OAI211_X1 U7002 ( .C1(n6193), .C2(n6070), .A(n6032), .B(n6031), .ZN(U3113)
         );
  AOI22_X1 U7003 ( .A1(n6195), .A2(n6035), .B1(n6043), .B2(n6196), .ZN(n6034)
         );
  AOI22_X1 U7004 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6037), .B1(n6194), 
        .B2(n6036), .ZN(n6033) );
  OAI211_X1 U7005 ( .C1(n6199), .C2(n6040), .A(n6034), .B(n6033), .ZN(U3114)
         );
  AOI22_X1 U7006 ( .A1(n6200), .A2(n6035), .B1(n6043), .B2(n6205), .ZN(n6039)
         );
  AOI22_X1 U7007 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6037), .B1(n6203), 
        .B2(n6036), .ZN(n6038) );
  OAI211_X1 U7008 ( .C1(n6210), .C2(n6040), .A(n6039), .B(n6038), .ZN(U3115)
         );
  NAND2_X1 U7009 ( .A1(n6073), .A2(n4264), .ZN(n6044) );
  OAI22_X1 U7010 ( .A1(n6044), .A2(n6370), .B1(n6042), .B2(n6041), .ZN(n6066)
         );
  NOR2_X1 U7011 ( .A1(n3479), .A2(n6078), .ZN(n6075) );
  NAND2_X1 U7012 ( .A1(n6349), .A2(n6075), .ZN(n6048) );
  INV_X1 U7013 ( .A(n6048), .ZN(n6065) );
  AOI22_X1 U7014 ( .A1(n6149), .A2(n6066), .B1(n6148), .B2(n6065), .ZN(n6052)
         );
  OAI21_X1 U7015 ( .B1(n6043), .B2(n6089), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6045) );
  AND3_X1 U7016 ( .A1(n6045), .A2(n6345), .A3(n6044), .ZN(n6046) );
  AOI211_X1 U7017 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6048), .A(n6047), .B(
        n6046), .ZN(n6050) );
  NAND2_X1 U7018 ( .A1(n6050), .A2(n6049), .ZN(n6067) );
  AOI22_X1 U7019 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n6067), .B1(n6112), 
        .B2(n6089), .ZN(n6051) );
  OAI211_X1 U7020 ( .C1(n6115), .C2(n6070), .A(n6052), .B(n6051), .ZN(U3116)
         );
  AOI22_X1 U7021 ( .A1(n6163), .A2(n6066), .B1(n6162), .B2(n6065), .ZN(n6054)
         );
  AOI22_X1 U7022 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n6067), .B1(n6116), 
        .B2(n6089), .ZN(n6053) );
  OAI211_X1 U7023 ( .C1(n6119), .C2(n6070), .A(n6054), .B(n6053), .ZN(U3117)
         );
  AOI22_X1 U7024 ( .A1(n6169), .A2(n6066), .B1(n6168), .B2(n6065), .ZN(n6056)
         );
  AOI22_X1 U7025 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n6067), .B1(n6120), 
        .B2(n6089), .ZN(n6055) );
  OAI211_X1 U7026 ( .C1(n6123), .C2(n6070), .A(n6056), .B(n6055), .ZN(U3118)
         );
  AOI22_X1 U7027 ( .A1(n6175), .A2(n6066), .B1(n6174), .B2(n6065), .ZN(n6058)
         );
  AOI22_X1 U7028 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n6067), .B1(n6124), 
        .B2(n6089), .ZN(n6057) );
  OAI211_X1 U7029 ( .C1(n6127), .C2(n6070), .A(n6058), .B(n6057), .ZN(U3119)
         );
  AOI22_X1 U7030 ( .A1(n6181), .A2(n6066), .B1(n6180), .B2(n6065), .ZN(n6060)
         );
  AOI22_X1 U7031 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n6067), .B1(n6128), 
        .B2(n6089), .ZN(n6059) );
  OAI211_X1 U7032 ( .C1(n6131), .C2(n6070), .A(n6060), .B(n6059), .ZN(U3120)
         );
  AOI22_X1 U7033 ( .A1(n6187), .A2(n6066), .B1(n6186), .B2(n6065), .ZN(n6062)
         );
  AOI22_X1 U7034 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n6067), .B1(n6132), 
        .B2(n6089), .ZN(n6061) );
  OAI211_X1 U7035 ( .C1(n6135), .C2(n6070), .A(n6062), .B(n6061), .ZN(U3121)
         );
  AOI22_X1 U7036 ( .A1(n6195), .A2(n6065), .B1(n6194), .B2(n6066), .ZN(n6064)
         );
  AOI22_X1 U7037 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n6067), .B1(n6196), 
        .B2(n6089), .ZN(n6063) );
  OAI211_X1 U7038 ( .C1(n6199), .C2(n6070), .A(n6064), .B(n6063), .ZN(U3122)
         );
  AOI22_X1 U7039 ( .A1(n6203), .A2(n6066), .B1(n6200), .B2(n6065), .ZN(n6069)
         );
  AOI22_X1 U7040 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n6067), .B1(n6205), 
        .B2(n6089), .ZN(n6068) );
  OAI211_X1 U7041 ( .C1(n6210), .C2(n6070), .A(n6069), .B(n6068), .ZN(U3123)
         );
  AND2_X1 U7042 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6075), .ZN(n6096)
         );
  AOI22_X1 U7043 ( .A1(n6148), .A2(n6096), .B1(n6107), .B2(n6112), .ZN(n6082)
         );
  AOI21_X1 U7044 ( .B1(n6146), .B2(n6073), .A(n6096), .ZN(n6080) );
  NAND3_X1 U7045 ( .A1(n6345), .A2(n6080), .A3(n6076), .ZN(n6074) );
  OAI211_X1 U7046 ( .C1(n6345), .C2(n6075), .A(n6156), .B(n6074), .ZN(n6098)
         );
  NAND2_X1 U7047 ( .A1(n6345), .A2(n6076), .ZN(n6079) );
  NAND2_X1 U7048 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6077) );
  OAI22_X1 U7049 ( .A1(n6080), .A2(n6079), .B1(n6078), .B2(n6077), .ZN(n6097)
         );
  AOI22_X1 U7050 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6098), .B1(n6149), 
        .B2(n6097), .ZN(n6081) );
  OAI211_X1 U7051 ( .C1(n6115), .C2(n6101), .A(n6082), .B(n6081), .ZN(U3124)
         );
  AOI22_X1 U7052 ( .A1(n6162), .A2(n6096), .B1(n6107), .B2(n6116), .ZN(n6084)
         );
  AOI22_X1 U7053 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6098), .B1(n6163), 
        .B2(n6097), .ZN(n6083) );
  OAI211_X1 U7054 ( .C1(n6119), .C2(n6101), .A(n6084), .B(n6083), .ZN(U3125)
         );
  AOI22_X1 U7055 ( .A1(n6168), .A2(n6096), .B1(n6107), .B2(n6120), .ZN(n6086)
         );
  AOI22_X1 U7056 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6098), .B1(n6169), 
        .B2(n6097), .ZN(n6085) );
  OAI211_X1 U7057 ( .C1(n6123), .C2(n6101), .A(n6086), .B(n6085), .ZN(U3126)
         );
  AOI22_X1 U7058 ( .A1(n6174), .A2(n6096), .B1(n6089), .B2(n6176), .ZN(n6088)
         );
  AOI22_X1 U7059 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6098), .B1(n6175), 
        .B2(n6097), .ZN(n6087) );
  OAI211_X1 U7060 ( .C1(n6179), .C2(n6143), .A(n6088), .B(n6087), .ZN(U3127)
         );
  AOI22_X1 U7061 ( .A1(n6180), .A2(n6096), .B1(n6089), .B2(n6182), .ZN(n6091)
         );
  AOI22_X1 U7062 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6098), .B1(n6181), 
        .B2(n6097), .ZN(n6090) );
  OAI211_X1 U7063 ( .C1(n6185), .C2(n6143), .A(n6091), .B(n6090), .ZN(U3128)
         );
  AOI22_X1 U7064 ( .A1(n6186), .A2(n6096), .B1(n6107), .B2(n6132), .ZN(n6093)
         );
  AOI22_X1 U7065 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6098), .B1(n6187), 
        .B2(n6097), .ZN(n6092) );
  OAI211_X1 U7066 ( .C1(n6135), .C2(n6101), .A(n6093), .B(n6092), .ZN(U3129)
         );
  AOI22_X1 U7067 ( .A1(n6195), .A2(n6096), .B1(n6107), .B2(n6196), .ZN(n6095)
         );
  AOI22_X1 U7068 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6098), .B1(n6194), 
        .B2(n6097), .ZN(n6094) );
  OAI211_X1 U7069 ( .C1(n6199), .C2(n6101), .A(n6095), .B(n6094), .ZN(U3130)
         );
  AOI22_X1 U7070 ( .A1(n6200), .A2(n6096), .B1(n6107), .B2(n6205), .ZN(n6100)
         );
  AOI22_X1 U7071 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6098), .B1(n6203), 
        .B2(n6097), .ZN(n6099) );
  OAI211_X1 U7072 ( .C1(n6210), .C2(n6101), .A(n6100), .B(n6099), .ZN(U3131)
         );
  OAI22_X1 U7073 ( .A1(n6104), .A2(n6103), .B1(n3479), .B2(n6102), .ZN(n6139)
         );
  NOR2_X1 U7074 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6147), .ZN(n6138)
         );
  AOI22_X1 U7075 ( .A1(n6149), .A2(n6139), .B1(n6148), .B2(n6138), .ZN(n6114)
         );
  NOR3_X1 U7076 ( .A1(n6106), .A2(n3479), .A3(n6105), .ZN(n6111) );
  OR2_X1 U7077 ( .A1(n6150), .A2(n6344), .ZN(n6209) );
  OAI21_X1 U7078 ( .B1(n6188), .B2(n6107), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6108) );
  NAND3_X1 U7079 ( .A1(n6109), .A2(n6345), .A3(n6108), .ZN(n6110) );
  AOI22_X1 U7080 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6140), .B1(n6112), 
        .B2(n6188), .ZN(n6113) );
  OAI211_X1 U7081 ( .C1(n6115), .C2(n6143), .A(n6114), .B(n6113), .ZN(U3132)
         );
  AOI22_X1 U7082 ( .A1(n6163), .A2(n6139), .B1(n6162), .B2(n6138), .ZN(n6118)
         );
  AOI22_X1 U7083 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6140), .B1(n6116), 
        .B2(n6188), .ZN(n6117) );
  OAI211_X1 U7084 ( .C1(n6119), .C2(n6143), .A(n6118), .B(n6117), .ZN(U3133)
         );
  AOI22_X1 U7085 ( .A1(n6169), .A2(n6139), .B1(n6168), .B2(n6138), .ZN(n6122)
         );
  AOI22_X1 U7086 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6140), .B1(n6120), 
        .B2(n6188), .ZN(n6121) );
  OAI211_X1 U7087 ( .C1(n6123), .C2(n6143), .A(n6122), .B(n6121), .ZN(U3134)
         );
  AOI22_X1 U7088 ( .A1(n6175), .A2(n6139), .B1(n6174), .B2(n6138), .ZN(n6126)
         );
  AOI22_X1 U7089 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6140), .B1(n6124), 
        .B2(n6188), .ZN(n6125) );
  OAI211_X1 U7090 ( .C1(n6127), .C2(n6143), .A(n6126), .B(n6125), .ZN(U3135)
         );
  AOI22_X1 U7091 ( .A1(n6181), .A2(n6139), .B1(n6180), .B2(n6138), .ZN(n6130)
         );
  AOI22_X1 U7092 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6140), .B1(n6128), 
        .B2(n6188), .ZN(n6129) );
  OAI211_X1 U7093 ( .C1(n6131), .C2(n6143), .A(n6130), .B(n6129), .ZN(U3136)
         );
  AOI22_X1 U7094 ( .A1(n6187), .A2(n6139), .B1(n6186), .B2(n6138), .ZN(n6134)
         );
  AOI22_X1 U7095 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6140), .B1(n6132), 
        .B2(n6188), .ZN(n6133) );
  OAI211_X1 U7096 ( .C1(n6135), .C2(n6143), .A(n6134), .B(n6133), .ZN(U3137)
         );
  AOI22_X1 U7097 ( .A1(n6195), .A2(n6138), .B1(n6194), .B2(n6139), .ZN(n6137)
         );
  AOI22_X1 U7098 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6140), .B1(n6196), 
        .B2(n6188), .ZN(n6136) );
  OAI211_X1 U7099 ( .C1(n6199), .C2(n6143), .A(n6137), .B(n6136), .ZN(U3138)
         );
  AOI22_X1 U7100 ( .A1(n6203), .A2(n6139), .B1(n6200), .B2(n6138), .ZN(n6142)
         );
  AOI22_X1 U7101 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6140), .B1(n6205), 
        .B2(n6188), .ZN(n6141) );
  OAI211_X1 U7102 ( .C1(n6210), .C2(n6143), .A(n6142), .B(n6141), .ZN(U3139)
         );
  INV_X1 U7103 ( .A(n6144), .ZN(n6201) );
  AOI21_X1 U7104 ( .B1(n6146), .B2(n6145), .A(n6201), .ZN(n6153) );
  OAI22_X1 U7105 ( .A1(n6153), .A2(n6370), .B1(n6147), .B2(n3558), .ZN(n6202)
         );
  AOI22_X1 U7106 ( .A1(n6149), .A2(n6202), .B1(n6201), .B2(n6148), .ZN(n6160)
         );
  INV_X1 U7107 ( .A(n6150), .ZN(n6152) );
  OAI21_X1 U7108 ( .B1(n6152), .B2(n5692), .A(n6151), .ZN(n6154) );
  NAND2_X1 U7109 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  OAI211_X1 U7110 ( .C1(n6345), .C2(n6157), .A(n6156), .B(n6155), .ZN(n6206)
         );
  AOI22_X1 U7111 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6206), .B1(n6158), 
        .B2(n6188), .ZN(n6159) );
  OAI211_X1 U7112 ( .C1(n6161), .C2(n6192), .A(n6160), .B(n6159), .ZN(U3140)
         );
  AOI22_X1 U7113 ( .A1(n6163), .A2(n6202), .B1(n6201), .B2(n6162), .ZN(n6166)
         );
  AOI22_X1 U7114 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6206), .B1(n6164), 
        .B2(n6188), .ZN(n6165) );
  OAI211_X1 U7115 ( .C1(n6167), .C2(n6192), .A(n6166), .B(n6165), .ZN(U3141)
         );
  AOI22_X1 U7116 ( .A1(n6169), .A2(n6202), .B1(n6201), .B2(n6168), .ZN(n6172)
         );
  AOI22_X1 U7117 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6206), .B1(n6170), 
        .B2(n6188), .ZN(n6171) );
  OAI211_X1 U7118 ( .C1(n6173), .C2(n6192), .A(n6172), .B(n6171), .ZN(U3142)
         );
  AOI22_X1 U7119 ( .A1(n6175), .A2(n6202), .B1(n6201), .B2(n6174), .ZN(n6178)
         );
  AOI22_X1 U7120 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6206), .B1(n6176), 
        .B2(n6188), .ZN(n6177) );
  OAI211_X1 U7121 ( .C1(n6179), .C2(n6192), .A(n6178), .B(n6177), .ZN(U3143)
         );
  AOI22_X1 U7122 ( .A1(n6181), .A2(n6202), .B1(n6201), .B2(n6180), .ZN(n6184)
         );
  AOI22_X1 U7123 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6206), .B1(n6182), 
        .B2(n6188), .ZN(n6183) );
  OAI211_X1 U7124 ( .C1(n6185), .C2(n6192), .A(n6184), .B(n6183), .ZN(U3144)
         );
  AOI22_X1 U7125 ( .A1(n6187), .A2(n6202), .B1(n6201), .B2(n6186), .ZN(n6191)
         );
  AOI22_X1 U7126 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6206), .B1(n6189), 
        .B2(n6188), .ZN(n6190) );
  OAI211_X1 U7127 ( .C1(n6193), .C2(n6192), .A(n6191), .B(n6190), .ZN(U3145)
         );
  AOI22_X1 U7128 ( .A1(n6195), .A2(n6201), .B1(n6194), .B2(n6202), .ZN(n6198)
         );
  AOI22_X1 U7129 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6206), .B1(n6196), 
        .B2(n6204), .ZN(n6197) );
  OAI211_X1 U7130 ( .C1(n6199), .C2(n6209), .A(n6198), .B(n6197), .ZN(U3146)
         );
  AOI22_X1 U7131 ( .A1(n6203), .A2(n6202), .B1(n6201), .B2(n6200), .ZN(n6208)
         );
  AOI22_X1 U7132 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6206), .B1(n6205), 
        .B2(n6204), .ZN(n6207) );
  OAI211_X1 U7133 ( .C1(n6210), .C2(n6209), .A(n6208), .B(n6207), .ZN(U3147)
         );
  NOR2_X1 U7134 ( .A1(n6212), .A2(n6211), .ZN(n6219) );
  OAI22_X1 U7135 ( .A1(n6219), .A2(n6218), .B1(n6220), .B2(n6213), .ZN(n6223)
         );
  AOI22_X1 U7136 ( .A1(n6347), .A2(n6215), .B1(n6214), .B2(n3024), .ZN(n6337)
         );
  NAND2_X1 U7137 ( .A1(n6216), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6343) );
  NAND3_X1 U7138 ( .A1(n6337), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6343), .ZN(n6217) );
  AOI21_X1 U7139 ( .B1(n6219), .B2(n6218), .A(n6217), .ZN(n6222) );
  INV_X1 U7140 ( .A(n6220), .ZN(n6221) );
  OAI22_X1 U7141 ( .A1(n6223), .A2(n6222), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6221), .ZN(n6224) );
  AOI222_X1 U7142 ( .A1(n6225), .A2(n3479), .B1(n6225), .B2(n6224), .C1(n3479), 
        .C2(n6224), .ZN(n6235) );
  INV_X1 U7143 ( .A(n6226), .ZN(n6232) );
  AOI21_X1 U7144 ( .B1(n6229), .B2(n6228), .A(n6227), .ZN(n6231) );
  NOR4_X1 U7145 ( .A1(n6233), .A2(n6232), .A3(n6231), .A4(n6230), .ZN(n6234)
         );
  OAI211_X1 U7146 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n6235), .A(n6244), .B(n6234), .ZN(n6247) );
  OR2_X1 U7147 ( .A1(n6247), .A2(n6236), .ZN(n6242) );
  NAND2_X1 U7148 ( .A1(READY_N), .A2(n6237), .ZN(n6241) );
  NOR2_X1 U7149 ( .A1(n6239), .A2(n6238), .ZN(n6240) );
  AOI21_X1 U7150 ( .B1(n6242), .B2(n6241), .A(n6240), .ZN(n6254) );
  INV_X1 U7151 ( .A(n6254), .ZN(n6330) );
  OAI21_X1 U7152 ( .B1(n6365), .B2(n6333), .A(n6330), .ZN(n6249) );
  NAND3_X1 U7153 ( .A1(n6245), .A2(n6244), .A3(n6243), .ZN(n6350) );
  AOI221_X1 U7154 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6330), .C1(n6271), .C2(
        n6330), .A(n6366), .ZN(n6250) );
  AOI211_X1 U7155 ( .C1(n6251), .C2(n6247), .A(n6246), .B(n6250), .ZN(n6248)
         );
  OAI221_X1 U7156 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6249), .C1(n6366), .C2(
        n6350), .A(n6248), .ZN(U3148) );
  NOR2_X1 U7157 ( .A1(n6250), .A2(n6254), .ZN(n6255) );
  NOR2_X1 U7158 ( .A1(READY_N), .A2(n6366), .ZN(n6258) );
  AOI21_X1 U7159 ( .B1(n6252), .B2(n6258), .A(n6251), .ZN(n6253) );
  OAI22_X1 U7160 ( .A1(n6425), .A2(n6255), .B1(n6254), .B2(n6253), .ZN(n6256)
         );
  OR2_X1 U7161 ( .A1(n6257), .A2(n6256), .ZN(U3149) );
  OAI211_X1 U7162 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6258), .A(n6329), .B(
        n6365), .ZN(n6259) );
  NAND2_X1 U7163 ( .A1(n6260), .A2(n6259), .ZN(U3150) );
  AND2_X1 U7164 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6324), .ZN(U3151) );
  AND2_X1 U7165 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6324), .ZN(U3152) );
  AND2_X1 U7166 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6324), .ZN(U3153) );
  AND2_X1 U7167 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6324), .ZN(U3154) );
  AND2_X1 U7168 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6324), .ZN(U3155) );
  AND2_X1 U7169 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6324), .ZN(U3156) );
  AND2_X1 U7170 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6324), .ZN(U3157) );
  AND2_X1 U7171 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6324), .ZN(U3158) );
  AND2_X1 U7172 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6324), .ZN(U3159) );
  AND2_X1 U7173 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6324), .ZN(U3160) );
  AND2_X1 U7174 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6324), .ZN(U3161) );
  AND2_X1 U7175 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6324), .ZN(U3162) );
  AND2_X1 U7176 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6324), .ZN(U3163) );
  AND2_X1 U7177 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6324), .ZN(U3164) );
  AND2_X1 U7178 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6324), .ZN(U3165) );
  AND2_X1 U7179 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6324), .ZN(U3166) );
  AND2_X1 U7180 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6324), .ZN(U3167) );
  AND2_X1 U7181 ( .A1(n6324), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  AND2_X1 U7182 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6324), .ZN(U3169) );
  AND2_X1 U7183 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6324), .ZN(U3170) );
  AND2_X1 U7184 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6324), .ZN(U3171) );
  AND2_X1 U7185 ( .A1(n6324), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  AND2_X1 U7186 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6324), .ZN(U3173) );
  AND2_X1 U7187 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6324), .ZN(U3174) );
  AND2_X1 U7188 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6324), .ZN(U3175) );
  AND2_X1 U7189 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6324), .ZN(U3176) );
  AND2_X1 U7190 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6324), .ZN(U3177) );
  AND2_X1 U7191 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6324), .ZN(U3178) );
  AND2_X1 U7192 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6324), .ZN(U3179) );
  AND2_X1 U7193 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6324), .ZN(U3180) );
  NOR2_X1 U7194 ( .A1(n6459), .A2(n6267), .ZN(n6268) );
  AOI22_X1 U7195 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6276) );
  AND2_X1 U7196 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6264) );
  INV_X1 U7197 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6262) );
  INV_X1 U7198 ( .A(NA_N), .ZN(n6269) );
  AOI221_X1 U7199 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6269), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6273) );
  AOI221_X1 U7200 ( .B1(n6264), .B2(n6543), .C1(n6262), .C2(n6543), .A(n6273), 
        .ZN(n6261) );
  OAI21_X1 U7201 ( .B1(n6268), .B2(n6276), .A(n6261), .ZN(U3181) );
  NOR2_X1 U7202 ( .A1(n6523), .A2(n6262), .ZN(n6270) );
  NAND2_X1 U7203 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6263) );
  OAI21_X1 U7204 ( .B1(n6270), .B2(n6264), .A(n6263), .ZN(n6265) );
  OAI211_X1 U7205 ( .C1(n6267), .C2(n6271), .A(n6266), .B(n6265), .ZN(U3182)
         );
  AOI21_X1 U7206 ( .B1(n6270), .B2(n6269), .A(n6268), .ZN(n6275) );
  AOI221_X1 U7207 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6271), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6272) );
  AOI221_X1 U7208 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6272), .C2(HOLD), .A(n6523), .ZN(n6274) );
  OAI22_X1 U7209 ( .A1(n6276), .A2(n6275), .B1(n6274), .B2(n6273), .ZN(U3183)
         );
  NOR2_X1 U7210 ( .A1(n6459), .A2(n6543), .ZN(n6542) );
  NOR2_X2 U7211 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6543), .ZN(n6541) );
  AOI22_X1 U7212 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6543), .ZN(n6277) );
  OAI21_X1 U7213 ( .B1(n6353), .B2(n6319), .A(n6277), .ZN(U3184) );
  AOI22_X1 U7214 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6543), .ZN(n6278) );
  OAI21_X1 U7215 ( .B1(n6279), .B2(n6319), .A(n6278), .ZN(U3185) );
  AOI22_X1 U7216 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6543), .ZN(n6280) );
  OAI21_X1 U7217 ( .B1(n6281), .B2(n6319), .A(n6280), .ZN(U3186) );
  AOI22_X1 U7218 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6543), .ZN(n6282) );
  OAI21_X1 U7219 ( .B1(n6283), .B2(n6319), .A(n6282), .ZN(U3187) );
  AOI22_X1 U7220 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6543), .ZN(n6284) );
  OAI21_X1 U7221 ( .B1(n6285), .B2(n6319), .A(n6284), .ZN(U3189) );
  AOI22_X1 U7222 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6543), .ZN(n6286) );
  OAI21_X1 U7223 ( .B1(n4406), .B2(n6319), .A(n6286), .ZN(U3190) );
  AOI22_X1 U7224 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6543), .ZN(n6287) );
  OAI21_X1 U7225 ( .B1(n6288), .B2(n6319), .A(n6287), .ZN(U3191) );
  AOI22_X1 U7226 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6543), .ZN(n6289) );
  OAI21_X1 U7227 ( .B1(n6290), .B2(n6319), .A(n6289), .ZN(U3192) );
  AOI22_X1 U7228 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6543), .ZN(n6291) );
  OAI21_X1 U7229 ( .B1(n6292), .B2(n6319), .A(n6291), .ZN(U3193) );
  INV_X1 U7230 ( .A(n6541), .ZN(n6321) );
  AOI22_X1 U7231 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6543), .ZN(n6293) );
  OAI21_X1 U7232 ( .B1(n4586), .B2(n6321), .A(n6293), .ZN(U3194) );
  AOI22_X1 U7233 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6543), .ZN(n6294) );
  OAI21_X1 U7234 ( .B1(n4586), .B2(n6319), .A(n6294), .ZN(U3195) );
  AOI22_X1 U7235 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6543), .ZN(n6295) );
  OAI21_X1 U7236 ( .B1(n6296), .B2(n6319), .A(n6295), .ZN(U3196) );
  AOI22_X1 U7237 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6543), .ZN(n6297) );
  OAI21_X1 U7238 ( .B1(n6440), .B2(n6321), .A(n6297), .ZN(U3197) );
  AOI22_X1 U7239 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6543), .ZN(n6298) );
  OAI21_X1 U7240 ( .B1(n6300), .B2(n6321), .A(n6298), .ZN(U3198) );
  AOI22_X1 U7241 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6543), .ZN(n6299) );
  OAI21_X1 U7242 ( .B1(n6300), .B2(n6319), .A(n6299), .ZN(U3199) );
  AOI22_X1 U7243 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6543), .ZN(n6301) );
  OAI21_X1 U7244 ( .B1(n6303), .B2(n6321), .A(n6301), .ZN(U3200) );
  AOI22_X1 U7245 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6543), .ZN(n6302) );
  OAI21_X1 U7246 ( .B1(n6303), .B2(n6319), .A(n6302), .ZN(U3201) );
  INV_X1 U7247 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6304) );
  OAI222_X1 U7248 ( .A1(n6319), .A2(n6305), .B1(n6304), .B2(n6376), .C1(n6307), 
        .C2(n6321), .ZN(U3202) );
  AOI22_X1 U7249 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6543), .ZN(n6306) );
  OAI21_X1 U7250 ( .B1(n6307), .B2(n6319), .A(n6306), .ZN(U3203) );
  AOI22_X1 U7251 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6543), .ZN(n6308) );
  OAI21_X1 U7252 ( .B1(n6310), .B2(n6321), .A(n6308), .ZN(U3204) );
  AOI22_X1 U7253 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6543), .ZN(n6309) );
  OAI21_X1 U7254 ( .B1(n6310), .B2(n6319), .A(n6309), .ZN(U3205) );
  AOI22_X1 U7255 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6543), .ZN(n6311) );
  OAI21_X1 U7256 ( .B1(n6430), .B2(n6321), .A(n6311), .ZN(U3206) );
  AOI22_X1 U7257 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6543), .ZN(n6312) );
  OAI21_X1 U7258 ( .B1(n6314), .B2(n6321), .A(n6312), .ZN(U3207) );
  AOI22_X1 U7259 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6543), .ZN(n6313) );
  OAI21_X1 U7260 ( .B1(n6314), .B2(n6319), .A(n6313), .ZN(U3208) );
  AOI22_X1 U7261 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6543), .ZN(n6315) );
  OAI21_X1 U7262 ( .B1(n3930), .B2(n6321), .A(n6315), .ZN(U3209) );
  AOI22_X1 U7263 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6543), .ZN(n6316) );
  OAI21_X1 U7264 ( .B1(n6447), .B2(n6321), .A(n6316), .ZN(U3210) );
  AOI22_X1 U7265 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6543), .ZN(n6317) );
  OAI21_X1 U7266 ( .B1(n6447), .B2(n6319), .A(n6317), .ZN(U3211) );
  AOI22_X1 U7267 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6541), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6543), .ZN(n6318) );
  OAI21_X1 U7268 ( .B1(n6421), .B2(n6319), .A(n6318), .ZN(U3212) );
  AOI22_X1 U7269 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6542), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6543), .ZN(n6320) );
  OAI21_X1 U7270 ( .B1(n6322), .B2(n6321), .A(n6320), .ZN(U3213) );
  MUX2_X1 U7271 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6376), .Z(U3445) );
  MUX2_X1 U7272 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6376), .Z(U3446) );
  MUX2_X1 U7273 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6376), .Z(U3447) );
  MUX2_X1 U7274 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6376), .Z(U3448) );
  INV_X1 U7275 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6325) );
  INV_X1 U7276 ( .A(n6326), .ZN(n6323) );
  AOI21_X1 U7277 ( .B1(n6325), .B2(n6324), .A(n6323), .ZN(U3451) );
  OAI21_X1 U7278 ( .B1(n6328), .B2(n6327), .A(n6326), .ZN(U3452) );
  OAI221_X1 U7279 ( .B1(n6331), .B2(STATE2_REG_0__SCAN_IN), .C1(n6331), .C2(
        n6330), .A(n6329), .ZN(U3453) );
  INV_X1 U7280 ( .A(n6332), .ZN(n6335) );
  OAI22_X1 U7281 ( .A1(n6335), .A2(n6342), .B1(n6334), .B2(n6333), .ZN(n6336)
         );
  MUX2_X1 U7282 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6336), .S(n6340), 
        .Z(U3456) );
  OAI22_X1 U7283 ( .A1(n6337), .A2(n6342), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6425), .ZN(n6339) );
  OAI22_X1 U7284 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6340), .B1(n6339), .B2(n6338), .ZN(n6341) );
  OAI21_X1 U7285 ( .B1(n6343), .B2(n6342), .A(n6341), .ZN(U3461) );
  AOI22_X1 U7286 ( .A1(n6347), .A2(n6346), .B1(n6345), .B2(n6344), .ZN(n6351)
         );
  OAI222_X1 U7287 ( .A1(n6352), .A2(n6351), .B1(n6352), .B2(n6350), .C1(n6349), 
        .C2(n6348), .ZN(U3465) );
  AOI21_X1 U7288 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6354) );
  AOI22_X1 U7289 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6354), .B2(n6353), .ZN(n6356) );
  INV_X1 U7290 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6355) );
  AOI22_X1 U7291 ( .A1(n6357), .A2(n6356), .B1(n6355), .B2(n6360), .ZN(U3468)
         );
  INV_X1 U7292 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6361) );
  NOR2_X1 U7293 ( .A1(n6360), .A2(REIP_REG_1__SCAN_IN), .ZN(n6358) );
  AOI22_X1 U7294 ( .A1(n6361), .A2(n6360), .B1(n6359), .B2(n6358), .ZN(U3469)
         );
  INV_X1 U7295 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6504) );
  MUX2_X1 U7296 ( .A(W_R_N_REG_SCAN_IN), .B(n6504), .S(n6376), .Z(U3470) );
  AOI211_X1 U7297 ( .C1(n6364), .C2(n6363), .A(n3558), .B(n6362), .ZN(n6367)
         );
  OAI21_X1 U7298 ( .B1(n6367), .B2(n6366), .A(n6365), .ZN(n6375) );
  INV_X1 U7299 ( .A(n6368), .ZN(n6373) );
  OAI211_X1 U7300 ( .C1(READY_N), .C2(n6371), .A(n6370), .B(n6369), .ZN(n6372)
         );
  NOR2_X1 U7301 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  MUX2_X1 U7302 ( .A(n6375), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6374), .Z(
        U3472) );
  MUX2_X1 U7303 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6376), .Z(U3473) );
  NAND2_X1 U7304 ( .A1(keyinput29), .A2(keyinput24), .ZN(n6382) );
  NOR2_X1 U7305 ( .A1(keyinput52), .A2(keyinput15), .ZN(n6380) );
  NAND3_X1 U7306 ( .A1(keyinput33), .A2(keyinput59), .A3(keyinput28), .ZN(
        n6378) );
  NAND3_X1 U7307 ( .A1(keyinput23), .A2(keyinput60), .A3(keyinput41), .ZN(
        n6377) );
  NOR4_X1 U7308 ( .A1(keyinput56), .A2(keyinput7), .A3(n6378), .A4(n6377), 
        .ZN(n6379) );
  NAND4_X1 U7309 ( .A1(keyinput14), .A2(keyinput34), .A3(n6380), .A4(n6379), 
        .ZN(n6381) );
  NOR4_X1 U7310 ( .A1(keyinput40), .A2(keyinput9), .A3(n6382), .A4(n6381), 
        .ZN(n6403) );
  NAND4_X1 U7311 ( .A1(keyinput39), .A2(keyinput1), .A3(keyinput45), .A4(
        keyinput26), .ZN(n6384) );
  NAND2_X1 U7312 ( .A1(keyinput22), .A2(keyinput44), .ZN(n6383) );
  NOR4_X1 U7313 ( .A1(keyinput58), .A2(keyinput19), .A3(n6384), .A4(n6383), 
        .ZN(n6402) );
  NAND3_X1 U7314 ( .A1(keyinput18), .A2(keyinput4), .A3(keyinput20), .ZN(n6386) );
  NAND3_X1 U7315 ( .A1(keyinput49), .A2(keyinput57), .A3(keyinput10), .ZN(
        n6385) );
  NOR4_X1 U7316 ( .A1(keyinput11), .A2(keyinput46), .A3(n6386), .A4(n6385), 
        .ZN(n6401) );
  NAND3_X1 U7317 ( .A1(keyinput42), .A2(keyinput51), .A3(keyinput47), .ZN(
        n6399) );
  NAND3_X1 U7318 ( .A1(keyinput63), .A2(keyinput13), .A3(keyinput21), .ZN(
        n6388) );
  NAND3_X1 U7319 ( .A1(keyinput61), .A2(keyinput25), .A3(keyinput27), .ZN(
        n6387) );
  NOR4_X1 U7320 ( .A1(keyinput31), .A2(keyinput62), .A3(n6388), .A4(n6387), 
        .ZN(n6389) );
  NAND4_X1 U7321 ( .A1(keyinput38), .A2(keyinput16), .A3(keyinput32), .A4(
        n6389), .ZN(n6398) );
  NAND2_X1 U7322 ( .A1(keyinput0), .A2(keyinput3), .ZN(n6390) );
  NOR3_X1 U7323 ( .A1(keyinput12), .A2(keyinput6), .A3(n6390), .ZN(n6396) );
  NOR3_X1 U7324 ( .A1(keyinput36), .A2(keyinput54), .A3(keyinput2), .ZN(n6395)
         );
  NAND2_X1 U7325 ( .A1(keyinput35), .A2(keyinput55), .ZN(n6393) );
  INV_X1 U7326 ( .A(keyinput37), .ZN(n6391) );
  NAND4_X1 U7327 ( .A1(keyinput48), .A2(keyinput53), .A3(keyinput30), .A4(
        n6391), .ZN(n6392) );
  NOR4_X1 U7328 ( .A1(keyinput17), .A2(keyinput8), .A3(n6393), .A4(n6392), 
        .ZN(n6394) );
  NAND4_X1 U7329 ( .A1(n6396), .A2(keyinput5), .A3(n6395), .A4(n6394), .ZN(
        n6397) );
  NOR4_X1 U7330 ( .A1(keyinput43), .A2(n6399), .A3(n6398), .A4(n6397), .ZN(
        n6400) );
  NAND4_X1 U7331 ( .A1(n6403), .A2(n6402), .A3(n6401), .A4(n6400), .ZN(n6404)
         );
  NAND2_X1 U7332 ( .A1(keyinput50), .A2(n6404), .ZN(n6540) );
  INV_X1 U7333 ( .A(keyinput38), .ZN(n6407) );
  INV_X1 U7334 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n6405) );
  AOI22_X1 U7335 ( .A1(keyinput50), .A2(n6405), .B1(DATAO_REG_8__SCAN_IN), 
        .B2(n6407), .ZN(n6406) );
  OAI21_X1 U7336 ( .B1(DATAO_REG_8__SCAN_IN), .B2(n6407), .A(n6406), .ZN(n6419) );
  INV_X1 U7337 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6410) );
  INV_X1 U7338 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6409) );
  AOI22_X1 U7339 ( .A1(n6410), .A2(keyinput16), .B1(n6409), .B2(keyinput42), 
        .ZN(n6408) );
  OAI221_X1 U7340 ( .B1(n6410), .B2(keyinput16), .C1(n6409), .C2(keyinput42), 
        .A(n6408), .ZN(n6418) );
  INV_X1 U7341 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6412) );
  AOI22_X1 U7342 ( .A1(n6413), .A2(keyinput51), .B1(n6412), .B2(keyinput47), 
        .ZN(n6411) );
  OAI221_X1 U7343 ( .B1(n6413), .B2(keyinput51), .C1(n6412), .C2(keyinput47), 
        .A(n6411), .ZN(n6417) );
  INV_X1 U7344 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6415) );
  AOI22_X1 U7345 ( .A1(n3510), .A2(keyinput43), .B1(n6415), .B2(keyinput63), 
        .ZN(n6414) );
  OAI221_X1 U7346 ( .B1(n3510), .B2(keyinput43), .C1(n6415), .C2(keyinput63), 
        .A(n6414), .ZN(n6416) );
  NOR4_X1 U7347 ( .A1(n6419), .A2(n6418), .A3(n6417), .A4(n6416), .ZN(n6471)
         );
  INV_X1 U7348 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6422) );
  AOI22_X1 U7349 ( .A1(n6422), .A2(keyinput31), .B1(keyinput13), .B2(n6421), 
        .ZN(n6420) );
  OAI221_X1 U7350 ( .B1(n6422), .B2(keyinput31), .C1(n6421), .C2(keyinput13), 
        .A(n6420), .ZN(n6435) );
  INV_X1 U7351 ( .A(keyinput21), .ZN(n6424) );
  AOI22_X1 U7352 ( .A1(n6425), .A2(keyinput61), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n6424), .ZN(n6423) );
  OAI221_X1 U7353 ( .B1(n6425), .B2(keyinput61), .C1(n6424), .C2(
        DATAO_REG_25__SCAN_IN), .A(n6423), .ZN(n6434) );
  INV_X1 U7354 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6428) );
  INV_X1 U7355 ( .A(keyinput62), .ZN(n6427) );
  AOI22_X1 U7356 ( .A1(n6428), .A2(keyinput25), .B1(ADDRESS_REG_8__SCAN_IN), 
        .B2(n6427), .ZN(n6426) );
  OAI221_X1 U7357 ( .B1(n6428), .B2(keyinput25), .C1(n6427), .C2(
        ADDRESS_REG_8__SCAN_IN), .A(n6426), .ZN(n6433) );
  AOI22_X1 U7358 ( .A1(n6431), .A2(keyinput27), .B1(n6430), .B2(keyinput33), 
        .ZN(n6429) );
  OAI221_X1 U7359 ( .B1(n6431), .B2(keyinput27), .C1(n6430), .C2(keyinput33), 
        .A(n6429), .ZN(n6432) );
  NOR4_X1 U7360 ( .A1(n6435), .A2(n6434), .A3(n6433), .A4(n6432), .ZN(n6470)
         );
  INV_X1 U7361 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6438) );
  AOI22_X1 U7362 ( .A1(n6438), .A2(keyinput59), .B1(keyinput56), .B2(n6437), 
        .ZN(n6436) );
  OAI221_X1 U7363 ( .B1(n6438), .B2(keyinput59), .C1(n6437), .C2(keyinput56), 
        .A(n6436), .ZN(n6451) );
  AOI22_X1 U7364 ( .A1(n6441), .A2(keyinput28), .B1(keyinput29), .B2(n6440), 
        .ZN(n6439) );
  OAI221_X1 U7365 ( .B1(n6441), .B2(keyinput28), .C1(n6440), .C2(keyinput29), 
        .A(n6439), .ZN(n6450) );
  INV_X1 U7366 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6444) );
  AOI22_X1 U7367 ( .A1(n6444), .A2(keyinput24), .B1(keyinput40), .B2(n6443), 
        .ZN(n6442) );
  OAI221_X1 U7368 ( .B1(n6444), .B2(keyinput24), .C1(n6443), .C2(keyinput40), 
        .A(n6442), .ZN(n6449) );
  INV_X1 U7369 ( .A(keyinput9), .ZN(n6446) );
  AOI22_X1 U7370 ( .A1(n6447), .A2(keyinput23), .B1(DATAO_REG_22__SCAN_IN), 
        .B2(n6446), .ZN(n6445) );
  OAI221_X1 U7371 ( .B1(n6447), .B2(keyinput23), .C1(n6446), .C2(
        DATAO_REG_22__SCAN_IN), .A(n6445), .ZN(n6448) );
  NOR4_X1 U7372 ( .A1(n6451), .A2(n6450), .A3(n6449), .A4(n6448), .ZN(n6469)
         );
  AOI22_X1 U7373 ( .A1(n6454), .A2(keyinput60), .B1(keyinput41), .B2(n6453), 
        .ZN(n6452) );
  OAI221_X1 U7374 ( .B1(n6454), .B2(keyinput60), .C1(n6453), .C2(keyinput41), 
        .A(n6452), .ZN(n6467) );
  INV_X1 U7375 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6457) );
  AOI22_X1 U7376 ( .A1(n6457), .A2(keyinput7), .B1(n6456), .B2(keyinput52), 
        .ZN(n6455) );
  OAI221_X1 U7377 ( .B1(n6457), .B2(keyinput7), .C1(n6456), .C2(keyinput52), 
        .A(n6455), .ZN(n6466) );
  INV_X1 U7378 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6460) );
  AOI22_X1 U7379 ( .A1(n6460), .A2(keyinput14), .B1(keyinput15), .B2(n6459), 
        .ZN(n6458) );
  OAI221_X1 U7380 ( .B1(n6460), .B2(keyinput14), .C1(n6459), .C2(keyinput15), 
        .A(n6458), .ZN(n6465) );
  INV_X1 U7381 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6463) );
  INV_X1 U7382 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6462) );
  AOI22_X1 U7383 ( .A1(n6463), .A2(keyinput34), .B1(keyinput11), .B2(n6462), 
        .ZN(n6461) );
  OAI221_X1 U7384 ( .B1(n6463), .B2(keyinput34), .C1(n6462), .C2(keyinput11), 
        .A(n6461), .ZN(n6464) );
  NOR4_X1 U7385 ( .A1(n6467), .A2(n6466), .A3(n6465), .A4(n6464), .ZN(n6468)
         );
  NAND4_X1 U7386 ( .A1(n6471), .A2(n6470), .A3(n6469), .A4(n6468), .ZN(n6539)
         );
  INV_X1 U7387 ( .A(keyinput10), .ZN(n6473) );
  AOI22_X1 U7388 ( .A1(n6474), .A2(keyinput19), .B1(DATAWIDTH_REG_10__SCAN_IN), 
        .B2(n6473), .ZN(n6472) );
  OAI221_X1 U7389 ( .B1(n6474), .B2(keyinput19), .C1(n6473), .C2(
        DATAWIDTH_REG_10__SCAN_IN), .A(n6472), .ZN(n6486) );
  AOI22_X1 U7390 ( .A1(n5462), .A2(keyinput57), .B1(n6476), .B2(keyinput46), 
        .ZN(n6475) );
  OAI221_X1 U7391 ( .B1(n5462), .B2(keyinput57), .C1(n6476), .C2(keyinput46), 
        .A(n6475), .ZN(n6485) );
  INV_X1 U7392 ( .A(keyinput58), .ZN(n6478) );
  AOI22_X1 U7393 ( .A1(n6479), .A2(keyinput12), .B1(ADDRESS_REG_0__SCAN_IN), 
        .B2(n6478), .ZN(n6477) );
  OAI221_X1 U7394 ( .B1(n6479), .B2(keyinput12), .C1(n6478), .C2(
        ADDRESS_REG_0__SCAN_IN), .A(n6477), .ZN(n6484) );
  INV_X1 U7395 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n6481) );
  AOI22_X1 U7396 ( .A1(n6482), .A2(keyinput22), .B1(n6481), .B2(keyinput44), 
        .ZN(n6480) );
  OAI221_X1 U7397 ( .B1(n6482), .B2(keyinput22), .C1(n6481), .C2(keyinput44), 
        .A(n6480), .ZN(n6483) );
  NOR4_X1 U7398 ( .A1(n6486), .A2(n6485), .A3(n6484), .A4(n6483), .ZN(n6537)
         );
  INV_X1 U7399 ( .A(keyinput20), .ZN(n6488) );
  AOI22_X1 U7400 ( .A1(n6489), .A2(keyinput39), .B1(DATAO_REG_19__SCAN_IN), 
        .B2(n6488), .ZN(n6487) );
  OAI221_X1 U7401 ( .B1(n6489), .B2(keyinput39), .C1(n6488), .C2(
        DATAO_REG_19__SCAN_IN), .A(n6487), .ZN(n6502) );
  INV_X1 U7402 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6492) );
  AOI22_X1 U7403 ( .A1(n6492), .A2(keyinput18), .B1(keyinput4), .B2(n6491), 
        .ZN(n6490) );
  OAI221_X1 U7404 ( .B1(n6492), .B2(keyinput18), .C1(n6491), .C2(keyinput4), 
        .A(n6490), .ZN(n6501) );
  INV_X1 U7405 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6495) );
  INV_X1 U7406 ( .A(keyinput26), .ZN(n6494) );
  AOI22_X1 U7407 ( .A1(n6495), .A2(keyinput49), .B1(DATAO_REG_6__SCAN_IN), 
        .B2(n6494), .ZN(n6493) );
  OAI221_X1 U7408 ( .B1(n6495), .B2(keyinput49), .C1(n6494), .C2(
        DATAO_REG_6__SCAN_IN), .A(n6493), .ZN(n6500) );
  INV_X1 U7409 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6498) );
  AOI22_X1 U7410 ( .A1(n6498), .A2(keyinput1), .B1(keyinput45), .B2(n6497), 
        .ZN(n6496) );
  OAI221_X1 U7411 ( .B1(n6498), .B2(keyinput1), .C1(n6497), .C2(keyinput45), 
        .A(n6496), .ZN(n6499) );
  NOR4_X1 U7412 ( .A1(n6502), .A2(n6501), .A3(n6500), .A4(n6499), .ZN(n6536)
         );
  INV_X1 U7413 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6505) );
  AOI22_X1 U7414 ( .A1(n6505), .A2(keyinput8), .B1(keyinput37), .B2(n6504), 
        .ZN(n6503) );
  OAI221_X1 U7415 ( .B1(n6505), .B2(keyinput8), .C1(n6504), .C2(keyinput37), 
        .A(n6503), .ZN(n6517) );
  INV_X1 U7416 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n6508) );
  INV_X1 U7417 ( .A(keyinput35), .ZN(n6507) );
  AOI22_X1 U7418 ( .A1(n6508), .A2(keyinput55), .B1(ADDRESS_REG_18__SCAN_IN), 
        .B2(n6507), .ZN(n6506) );
  OAI221_X1 U7419 ( .B1(n6508), .B2(keyinput55), .C1(n6507), .C2(
        ADDRESS_REG_18__SCAN_IN), .A(n6506), .ZN(n6516) );
  INV_X1 U7420 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6511) );
  AOI22_X1 U7421 ( .A1(n6511), .A2(keyinput32), .B1(keyinput30), .B2(n6510), 
        .ZN(n6509) );
  OAI221_X1 U7422 ( .B1(n6511), .B2(keyinput32), .C1(n6510), .C2(keyinput30), 
        .A(n6509), .ZN(n6515) );
  INV_X1 U7423 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6513) );
  AOI22_X1 U7424 ( .A1(n4844), .A2(keyinput48), .B1(keyinput53), .B2(n6513), 
        .ZN(n6512) );
  OAI221_X1 U7425 ( .B1(n4844), .B2(keyinput48), .C1(n6513), .C2(keyinput53), 
        .A(n6512), .ZN(n6514) );
  NOR4_X1 U7426 ( .A1(n6517), .A2(n6516), .A3(n6515), .A4(n6514), .ZN(n6535)
         );
  INV_X1 U7427 ( .A(keyinput36), .ZN(n6519) );
  AOI22_X1 U7428 ( .A1(n6520), .A2(keyinput54), .B1(DATAWIDTH_REG_14__SCAN_IN), 
        .B2(n6519), .ZN(n6518) );
  OAI221_X1 U7429 ( .B1(n6520), .B2(keyinput54), .C1(n6519), .C2(
        DATAWIDTH_REG_14__SCAN_IN), .A(n6518), .ZN(n6533) );
  INV_X1 U7430 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6522) );
  AOI22_X1 U7431 ( .A1(n6523), .A2(keyinput3), .B1(n6522), .B2(keyinput6), 
        .ZN(n6521) );
  OAI221_X1 U7432 ( .B1(n6523), .B2(keyinput3), .C1(n6522), .C2(keyinput6), 
        .A(n6521), .ZN(n6532) );
  INV_X1 U7433 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6525) );
  AOI22_X1 U7434 ( .A1(n6526), .A2(keyinput0), .B1(n6525), .B2(keyinput5), 
        .ZN(n6524) );
  OAI221_X1 U7435 ( .B1(n6526), .B2(keyinput0), .C1(n6525), .C2(keyinput5), 
        .A(n6524), .ZN(n6531) );
  XOR2_X1 U7436 ( .A(n6527), .B(keyinput17), .Z(n6529) );
  XNOR2_X1 U7437 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput2), .ZN(
        n6528) );
  NAND2_X1 U7438 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  NOR4_X1 U7439 ( .A1(n6533), .A2(n6532), .A3(n6531), .A4(n6530), .ZN(n6534)
         );
  NAND4_X1 U7440 ( .A1(n6537), .A2(n6536), .A3(n6535), .A4(n6534), .ZN(n6538)
         );
  AOI211_X1 U7441 ( .C1(DATAO_REG_9__SCAN_IN), .C2(n6540), .A(n6539), .B(n6538), .ZN(n6545) );
  AOI222_X1 U7442 ( .A1(n6543), .A2(ADDRESS_REG_4__SCAN_IN), .B1(
        REIP_REG_5__SCAN_IN), .B2(n6542), .C1(REIP_REG_6__SCAN_IN), .C2(n6541), 
        .ZN(n6544) );
  XNOR2_X1 U7443 ( .A(n6545), .B(n6544), .ZN(U3188) );
  AND4_X1 U3430 ( .A1(n3087), .A2(n3086), .A3(n3085), .A4(n3084), .ZN(n3088)
         );
  CLKBUF_X2 U3406 ( .A(n3242), .Z(n3230) );
  CLKBUF_X1 U3416 ( .A(n3242), .Z(n4139) );
  CLKBUF_X1 U3436 ( .A(n4845), .Z(n4846) );
  CLKBUF_X1 U3503 ( .A(n3157), .Z(n5690) );
  CLKBUF_X1 U3885 ( .A(n2956), .Z(n3178) );
  CLKBUF_X1 U4130 ( .A(n3159), .Z(n2956) );
endmodule

