

module b22_C_SARLock_k_64_3 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6432, n6433, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331;

  NAND2_X1 U7181 ( .A1(n13263), .A2(n13248), .ZN(n13243) );
  NAND2_X2 U7182 ( .A1(n8983), .A2(n8982), .ZN(n13487) );
  NAND2_X1 U7183 ( .A1(n13718), .A2(n13613), .ZN(n13617) );
  INV_X1 U7184 ( .A(n10692), .ZN(n6937) );
  NAND2_X1 U7185 ( .A1(n11633), .A2(n11630), .ZN(n15070) );
  INV_X1 U7186 ( .A(n9527), .ZN(n11980) );
  INV_X2 U7187 ( .A(n11608), .ZN(n7726) );
  INV_X1 U7188 ( .A(n7677), .ZN(n12862) );
  XNOR2_X2 U7189 ( .A(n7675), .B(P3_IR_REG_29__SCAN_IN), .ZN(n7677) );
  INV_X1 U7190 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8521) );
  OAI21_X1 U7191 ( .B1(n10379), .B2(n7728), .A(n10378), .ZN(n10474) );
  INV_X1 U7192 ( .A(n8493), .ZN(n9795) );
  AND2_X1 U7193 ( .A1(n11457), .A2(n11456), .ZN(n11460) );
  NAND2_X1 U7194 ( .A1(n14339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9191) );
  OR2_X1 U7195 ( .A1(n11970), .A2(n14357), .ZN(n9636) );
  AND2_X1 U7196 ( .A1(n8719), .A2(n8718), .ZN(n7475) );
  OAI21_X1 U7197 ( .B1(n12198), .B2(n6749), .A(n6746), .ZN(n12216) );
  AOI21_X1 U7198 ( .B1(n12294), .B2(n12564), .A(n12163), .ZN(n12264) );
  INV_X1 U7199 ( .A(n11604), .ZN(n9659) );
  INV_X1 U7200 ( .A(n8029), .ZN(n8193) );
  INV_X1 U7201 ( .A(n11754), .ZN(n11748) );
  OAI211_X1 U7202 ( .C1(n10278), .C2(n10176), .A(n7693), .B(n7692), .ZN(n15063) );
  INV_X2 U7203 ( .A(n8537), .ZN(n9073) );
  INV_X1 U7204 ( .A(n9025), .ZN(n8767) );
  NAND2_X1 U7205 ( .A1(n13250), .A2(n13239), .ZN(n13238) );
  NAND2_X1 U7206 ( .A1(n10952), .A2(n14948), .ZN(n11115) );
  INV_X1 U7207 ( .A(n14931), .ZN(n6592) );
  OAI211_X1 U7208 ( .C1(n8493), .C2(n14775), .A(n8545), .B(n8544), .ZN(n10819)
         );
  INV_X1 U7209 ( .A(n8518), .ZN(n9100) );
  INV_X1 U7210 ( .A(n11978), .ZN(n9446) );
  OR2_X1 U7211 ( .A1(n10455), .A2(n10155), .ZN(n14229) );
  OAI21_X2 U7212 ( .B1(n12264), .B2(n12168), .A(n6555), .ZN(n12239) );
  XNOR2_X1 U7213 ( .A(n12162), .B(n12160), .ZN(n12294) );
  AND2_X1 U7214 ( .A1(n6941), .A2(n8231), .ZN(n9891) );
  NAND2_X1 U7215 ( .A1(n12850), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7673) );
  INV_X2 U7216 ( .A(n6439), .ZN(n9833) );
  OR2_X1 U7217 ( .A1(n13243), .A2(n7150), .ZN(n13199) );
  NAND2_X1 U7218 ( .A1(n13573), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8462) );
  INV_X2 U7219 ( .A(n6439), .ZN(n9479) );
  AOI211_X1 U7220 ( .C1(n13492), .C2(n13093), .A(n12949), .B(n12948), .ZN(
        n12953) );
  XNOR2_X1 U7221 ( .A(n9583), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14357) );
  CLKBUF_X3 U7222 ( .A(n10255), .Z(n6433) );
  NAND2_X2 U7223 ( .A1(n7134), .A2(n9243), .ZN(n13870) );
  NOR2_X2 U7225 ( .A1(n13428), .A2(n13434), .ZN(n7144) );
  NAND2_X4 U7226 ( .A1(n7191), .A2(n7190), .ZN(n10597) );
  NOR2_X2 U7227 ( .A1(n10530), .A2(n7324), .ZN(n7323) );
  INV_X4 U7228 ( .A(n13749), .ZN(n13704) );
  NAND2_X4 U7229 ( .A1(n10760), .A2(n13699), .ZN(n13749) );
  NAND2_X1 U7230 ( .A1(n8191), .A2(n8192), .ZN(n6432) );
  NOR4_X2 U7231 ( .A1(n9143), .A2(n9142), .A3(n12118), .A4(n9141), .ZN(n9144)
         );
  INV_X2 U7232 ( .A(n9197), .ZN(n9196) );
  XNOR2_X2 U7233 ( .A(n8437), .B(n8436), .ZN(n9693) );
  OAI211_X2 U7234 ( .C1(n9527), .C2(n9838), .A(n6486), .B(n7178), .ZN(n11832)
         );
  AND2_X2 U7235 ( .A1(n11825), .A2(n11824), .ZN(n10748) );
  XNOR2_X2 U7236 ( .A(n8462), .B(n13574), .ZN(n8467) );
  NOR2_X4 U7237 ( .A1(n7719), .A2(n7574), .ZN(n7770) );
  XNOR2_X2 U7238 ( .A(n9191), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9197) );
  OAI211_X1 U7240 ( .C1(n10317), .C2(n10176), .A(n7725), .B(n7724), .ZN(n15057) );
  XNOR2_X2 U7241 ( .A(n7673), .B(n12851), .ZN(n7678) );
  NAND2_X2 U7242 ( .A1(n11642), .A2(n11632), .ZN(n10546) );
  XNOR2_X2 U7243 ( .A(n8464), .B(n8463), .ZN(n8466) );
  OAI211_X1 U7245 ( .C1(n10179), .C2(n6432), .A(n7701), .B(n7700), .ZN(n10503)
         );
  NAND3_X1 U7247 ( .A1(n8781), .A2(n8564), .A3(n8420), .ZN(n8784) );
  XNOR2_X2 U7248 ( .A(n13487), .B(n12080), .ZN(n13279) );
  XNOR2_X2 U7249 ( .A(n9587), .B(n9586), .ZN(n11981) );
  NAND2_X2 U7250 ( .A1(n9585), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9587) );
  AOI21_X1 U7251 ( .B1(n14342), .B2(n9100), .A(n6575), .ZN(n13458) );
  OAI21_X1 U7252 ( .B1(n13031), .B2(n6640), .A(n6462), .ZN(n12976) );
  NAND2_X1 U7253 ( .A1(n11460), .A2(n11459), .ZN(n12061) );
  OR2_X1 U7254 ( .A1(n14413), .A2(n11897), .ZN(n14225) );
  AND2_X1 U7255 ( .A1(n15010), .A2(n11081), .ZN(n11240) );
  NAND2_X2 U7256 ( .A1(n10438), .A2(n10439), .ZN(n10454) );
  INV_X1 U7257 ( .A(n11993), .ZN(n6438) );
  NAND2_X1 U7258 ( .A1(n9286), .A2(n9285), .ZN(n14724) );
  AOI21_X1 U7259 ( .B1(n8164), .B2(n8165), .A(n6529), .ZN(n7292) );
  INV_X2 U7260 ( .A(n10597), .ZN(n12159) );
  INV_X4 U7261 ( .A(n11903), .ZN(n6435) );
  NAND4_X1 U7262 ( .A1(n8512), .A2(n8511), .A3(n8510), .A4(n8509), .ZN(n13115)
         );
  INV_X1 U7263 ( .A(n13111), .ZN(n10864) );
  NAND4_X1 U7264 ( .A1(n8557), .A2(n8556), .A3(n8555), .A4(n8554), .ZN(n13113)
         );
  NAND2_X1 U7265 ( .A1(n12771), .A2(n10503), .ZN(n12770) );
  INV_X1 U7266 ( .A(n13874), .ZN(n10753) );
  INV_X4 U7267 ( .A(n13752), .ZN(n13608) );
  INV_X2 U7268 ( .A(n12966), .ZN(n12900) );
  INV_X4 U7270 ( .A(n10426), .ZN(n13752) );
  INV_X2 U7271 ( .A(n9122), .ZN(n6436) );
  CLKBUF_X3 U7272 ( .A(n9099), .Z(n6442) );
  NAND2_X1 U7273 ( .A1(n7678), .A2(n12862), .ZN(n11608) );
  NAND2_X1 U7274 ( .A1(n6432), .A2(n9833), .ZN(n7772) );
  NAND2_X1 U7275 ( .A1(n6439), .A2(n9863), .ZN(n9527) );
  INV_X1 U7276 ( .A(n8466), .ZN(n7235) );
  NOR2_X2 U7277 ( .A1(n8143), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8134) );
  INV_X2 U7278 ( .A(n7689), .ZN(n6437) );
  AND3_X1 U7280 ( .A1(n6920), .A2(n7419), .A3(n6545), .ZN(n11797) );
  AND2_X1 U7281 ( .A1(n7277), .A2(n7276), .ZN(n7557) );
  MUX2_X1 U7282 ( .A(n12787), .B(n12786), .S(n15136), .Z(n12788) );
  MUX2_X1 U7283 ( .A(n12707), .B(n12786), .S(n15149), .Z(n12708) );
  NOR2_X1 U7284 ( .A1(n7272), .A2(n7271), .ZN(n7270) );
  NOR2_X1 U7285 ( .A1(n6499), .A2(n6961), .ZN(n6960) );
  NAND2_X1 U7286 ( .A1(n6971), .A2(n6973), .ZN(n9171) );
  AND2_X1 U7287 ( .A1(n14255), .A2(n14254), .ZN(n14256) );
  AOI21_X1 U7288 ( .B1(n14000), .B2(n14403), .A(n13999), .ZN(n14257) );
  NAND2_X1 U7289 ( .A1(n13066), .A2(n6636), .ZN(n12921) );
  AND2_X1 U7290 ( .A1(n14248), .A2(n6556), .ZN(n7082) );
  AOI21_X1 U7291 ( .B1(n6632), .B2(n6447), .A(n6974), .ZN(n6973) );
  NAND2_X1 U7292 ( .A1(n7327), .A2(n6508), .ZN(n13066) );
  OR2_X1 U7293 ( .A1(n14009), .A2(n14008), .ZN(n14251) );
  NAND2_X1 U7294 ( .A1(n7325), .A2(n7328), .ZN(n13067) );
  NOR4_X1 U7295 ( .A1(n12016), .A2(n12013), .A3(n12014), .A4(n12015), .ZN(
        n12017) );
  OR2_X1 U7296 ( .A1(n12905), .A2(n7330), .ZN(n7325) );
  NAND2_X1 U7297 ( .A1(n8128), .A2(n8127), .ZN(n12213) );
  AND2_X1 U7298 ( .A1(n7641), .A2(n11963), .ZN(n6831) );
  AND2_X1 U7299 ( .A1(n7251), .A2(n7250), .ZN(n7244) );
  INV_X1 U7300 ( .A(n7329), .ZN(n7328) );
  OAI21_X1 U7301 ( .B1(n9654), .B2(n9653), .A(n9655), .ZN(n11596) );
  OR2_X1 U7302 ( .A1(n7068), .A2(n7067), .ZN(n7065) );
  AND2_X1 U7303 ( .A1(n12084), .A2(n9127), .ZN(n13207) );
  AOI21_X1 U7304 ( .B1(n14342), .B2(n11980), .A(n11979), .ZN(n14240) );
  NAND2_X1 U7305 ( .A1(n6627), .A2(n9042), .ZN(n13462) );
  NAND2_X1 U7306 ( .A1(n8430), .A2(n8429), .ZN(n13477) );
  NAND3_X1 U7307 ( .A1(n9065), .A2(n9064), .A3(n9063), .ZN(n14342) );
  NAND2_X1 U7308 ( .A1(n12073), .A2(n7459), .ZN(n13331) );
  NAND2_X1 U7309 ( .A1(n12113), .A2(n12112), .ZN(n13254) );
  NAND2_X1 U7310 ( .A1(n7255), .A2(n9128), .ZN(n7254) );
  NAND2_X1 U7311 ( .A1(n9069), .A2(n9068), .ZN(n13465) );
  NAND2_X1 U7312 ( .A1(n9529), .A2(n9528), .ZN(n14264) );
  OAI21_X1 U7313 ( .B1(n8107), .B2(n8106), .A(n8108), .ZN(n8120) );
  AND2_X1 U7314 ( .A1(n7360), .A2(n6806), .ZN(n6805) );
  NAND2_X1 U7315 ( .A1(n13059), .A2(n12887), .ZN(n13031) );
  NAND2_X1 U7316 ( .A1(n13346), .A2(n13347), .ZN(n12073) );
  NAND2_X1 U7317 ( .A1(n7060), .A2(n12071), .ZN(n13346) );
  XNOR2_X1 U7318 ( .A(n9066), .B(n9067), .ZN(n12056) );
  XNOR2_X1 U7319 ( .A(n7507), .B(n6628), .ZN(n11591) );
  NAND2_X1 U7320 ( .A1(n13013), .A2(n6654), .ZN(n13059) );
  NAND2_X1 U7321 ( .A1(n9517), .A2(n9516), .ZN(n14269) );
  AOI21_X1 U7322 ( .B1(n7513), .B2(n7511), .A(n7510), .ZN(n7507) );
  NAND2_X1 U7323 ( .A1(n9504), .A2(n9503), .ZN(n14274) );
  XNOR2_X1 U7324 ( .A(n9035), .B(n9020), .ZN(n11589) );
  AND2_X1 U7325 ( .A1(n8981), .A2(n8980), .ZN(n13587) );
  NAND2_X1 U7326 ( .A1(n8978), .A2(n8979), .ZN(n8980) );
  AOI21_X1 U7327 ( .B1(n13362), .B2(n6711), .A(n6709), .ZN(n6708) );
  XNOR2_X1 U7328 ( .A(n12409), .B(n14391), .ZN(n12390) );
  NAND2_X1 U7329 ( .A1(n7258), .A2(n6710), .ZN(n6709) );
  NAND2_X1 U7330 ( .A1(n8957), .A2(n8956), .ZN(n13492) );
  NAND2_X1 U7331 ( .A1(n12942), .A2(n12870), .ZN(n12872) );
  NAND2_X1 U7332 ( .A1(n8939), .A2(n8938), .ZN(n13498) );
  NOR2_X1 U7333 ( .A1(n13334), .A2(n7460), .ZN(n7459) );
  NAND2_X1 U7334 ( .A1(n12866), .A2(n7334), .ZN(n12942) );
  NAND2_X1 U7335 ( .A1(n6711), .A2(n6472), .ZN(n6710) );
  NAND2_X1 U7336 ( .A1(n7281), .A2(n7280), .ZN(n12627) );
  NAND2_X1 U7337 ( .A1(n13719), .A2(n13720), .ZN(n13718) );
  NAND2_X1 U7338 ( .A1(n9468), .A2(n9467), .ZN(n14288) );
  NAND2_X1 U7339 ( .A1(n8054), .A2(n8053), .ZN(n8065) );
  AOI21_X1 U7340 ( .B1(n7040), .B2(n7042), .A(n6520), .ZN(n7039) );
  NOR2_X1 U7341 ( .A1(n7133), .A2(n7132), .ZN(n7131) );
  NAND2_X1 U7342 ( .A1(n6752), .A2(n6750), .ZN(n12285) );
  OAI21_X1 U7343 ( .B1(n13427), .B2(n12098), .A(n12097), .ZN(n13416) );
  OAI21_X1 U7344 ( .B1(n11587), .B2(n9527), .A(n9459), .ZN(n14293) );
  NAND2_X1 U7345 ( .A1(n7160), .A2(n7159), .ZN(n11472) );
  NAND2_X1 U7346 ( .A1(n8896), .A2(n8895), .ZN(n11587) );
  OAI21_X1 U7347 ( .B1(n13452), .B2(n12095), .A(n12096), .ZN(n13427) );
  OR2_X1 U7348 ( .A1(n14214), .A2(n14508), .ZN(n11901) );
  NOR2_X1 U7349 ( .A1(n14214), .A2(n14222), .ZN(n9400) );
  OR2_X1 U7350 ( .A1(n7514), .A2(n7515), .ZN(n8896) );
  OR2_X1 U7351 ( .A1(n6731), .A2(n6730), .ZN(n13452) );
  NAND2_X1 U7352 ( .A1(n11396), .A2(n9749), .ZN(n11422) );
  NAND2_X1 U7353 ( .A1(n11185), .A2(n11186), .ZN(n11396) );
  NAND2_X1 U7354 ( .A1(n8172), .A2(n14473), .ZN(n7274) );
  NAND2_X1 U7355 ( .A1(n9391), .A2(n9390), .ZN(n14214) );
  XNOR2_X1 U7356 ( .A(n11240), .B(n11241), .ZN(n11082) );
  OR2_X1 U7357 ( .A1(n8401), .A2(n10424), .ZN(n7072) );
  AND2_X1 U7358 ( .A1(n11147), .A2(n9743), .ZN(n11185) );
  OAI22_X1 U7359 ( .A1(n8878), .A2(n8877), .B1(SI_19_), .B2(n8400), .ZN(n8401)
         );
  NAND2_X1 U7360 ( .A1(n9363), .A2(n9362), .ZN(n11897) );
  AOI21_X1 U7361 ( .B1(n8399), .B2(n7026), .A(n7025), .ZN(n8878) );
  NAND2_X1 U7362 ( .A1(n6857), .A2(n6856), .ZN(n15010) );
  XNOR2_X1 U7363 ( .A(n8821), .B(n8820), .ZN(n10337) );
  NAND2_X1 U7364 ( .A1(n8727), .A2(n8726), .ZN(n12092) );
  NAND2_X1 U7365 ( .A1(n8763), .A2(n8819), .ZN(n8821) );
  OR2_X1 U7366 ( .A1(n8762), .A2(n9889), .ZN(n8763) );
  NAND3_X1 U7367 ( .A1(n7291), .A2(n7292), .A3(n8166), .ZN(n11092) );
  NOR2_X1 U7368 ( .A1(n6474), .A2(n11065), .ZN(n11251) );
  AND2_X1 U7369 ( .A1(n7156), .A2(n7155), .ZN(n11075) );
  NOR2_X1 U7370 ( .A1(n12996), .A2(n14885), .ZN(n13046) );
  NAND2_X1 U7371 ( .A1(n8638), .A2(n8637), .ZN(n11109) );
  NAND2_X1 U7372 ( .A1(n6618), .A2(n8375), .ZN(n8719) );
  NAND2_X1 U7373 ( .A1(n10525), .A2(n10524), .ZN(n10523) );
  NAND2_X1 U7374 ( .A1(n9298), .A2(n9297), .ZN(n15310) );
  NAND2_X1 U7375 ( .A1(n8662), .A2(n8661), .ZN(n11232) );
  XNOR2_X1 U7376 ( .A(n8632), .B(n8631), .ZN(n9873) );
  NAND2_X1 U7377 ( .A1(n9272), .A2(n9271), .ZN(n14647) );
  XNOR2_X1 U7378 ( .A(n6933), .B(n10772), .ZN(n10578) );
  NAND2_X1 U7379 ( .A1(n7172), .A2(n7171), .ZN(n6933) );
  INV_X1 U7380 ( .A(n10845), .ZN(n14927) );
  XNOR2_X1 U7381 ( .A(n13113), .B(n10845), .ZN(n10836) );
  AOI21_X1 U7382 ( .B1(n13871), .B2(n13704), .A(n10447), .ZN(n10606) );
  OAI21_X1 U7383 ( .B1(n8591), .B2(n8590), .A(n8592), .ZN(n9859) );
  NAND2_X1 U7384 ( .A1(n7145), .A2(n10658), .ZN(n10673) );
  OR2_X1 U7385 ( .A1(n9248), .A2(n9247), .ZN(n14700) );
  NAND2_X1 U7386 ( .A1(n8592), .A2(n8362), .ZN(n8613) );
  OR2_X1 U7387 ( .A1(n8567), .A2(n8566), .ZN(n10845) );
  OAI211_X1 U7388 ( .C1(n6726), .C2(n6725), .A(n8590), .B(n6723), .ZN(n8592)
         );
  NAND2_X1 U7389 ( .A1(n8214), .A2(n8213), .ZN(n10539) );
  NAND2_X1 U7390 ( .A1(n14906), .A2(n14867), .ZN(n14866) );
  NAND2_X1 U7391 ( .A1(n6530), .A2(n9211), .ZN(n9212) );
  AND4_X1 U7392 ( .A1(n8499), .A2(n8498), .A3(n8497), .A4(n8496), .ZN(n10398)
         );
  AND2_X1 U7393 ( .A1(n6611), .A2(n7090), .ZN(n7089) );
  NAND4_X2 U7394 ( .A1(n7718), .A2(n7717), .A3(n7716), .A4(n7715), .ZN(n15067)
         );
  OR2_X1 U7395 ( .A1(n10376), .A2(n10375), .ZN(n10480) );
  INV_X1 U7396 ( .A(n7498), .ZN(n7092) );
  NAND3_X2 U7397 ( .A1(n7349), .A2(n7348), .A3(n7346), .ZN(n12966) );
  AND3_X1 U7398 ( .A1(n7761), .A2(n7760), .A3(n7759), .ZN(n11007) );
  NAND4_X1 U7399 ( .A1(n7786), .A2(n7785), .A3(n7784), .A4(n7783), .ZN(n12358)
         );
  NAND2_X1 U7401 ( .A1(n6516), .A2(n9222), .ZN(n13872) );
  OR2_X2 U7402 ( .A1(n11823), .A2(n10457), .ZN(n13754) );
  NAND4_X2 U7403 ( .A1(n9232), .A2(n9231), .A3(n9230), .A4(n9229), .ZN(n13871)
         );
  NAND2_X1 U7404 ( .A1(n9694), .A2(n10655), .ZN(n9122) );
  XNOR2_X1 U7405 ( .A(n7993), .B(n7992), .ZN(n12459) );
  NAND2_X1 U7406 ( .A1(n8467), .A2(n8466), .ZN(n8507) );
  OAI21_X1 U7407 ( .B1(n6476), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7993) );
  CLKBUF_X1 U7408 ( .A(n11970), .Z(n6895) );
  NAND2_X2 U7409 ( .A1(n9863), .A2(n9833), .ZN(n11978) );
  OAI21_X1 U7410 ( .B1(n7502), .B2(n7500), .A(n8367), .ZN(n7499) );
  INV_X2 U7411 ( .A(n11603), .ZN(n9662) );
  AND2_X4 U7412 ( .A1(n9196), .A2(n11592), .ZN(n9228) );
  NAND2_X4 U7413 ( .A1(n9197), .A2(n9195), .ZN(n9520) );
  NAND2_X2 U7414 ( .A1(n9641), .A2(n14344), .ZN(n9863) );
  AND2_X1 U7415 ( .A1(n8205), .A2(n8204), .ZN(n8231) );
  NAND2_X1 U7416 ( .A1(n8210), .A2(n6475), .ZN(n11104) );
  AND2_X2 U7417 ( .A1(n7678), .A2(n7677), .ZN(n11603) );
  NAND2_X1 U7418 ( .A1(n8440), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8437) );
  INV_X1 U7419 ( .A(n8449), .ZN(n11137) );
  MUX2_X1 U7420 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8209), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8210) );
  XNOR2_X1 U7421 ( .A(n6610), .B(n7671), .ZN(n8192) );
  AND2_X1 U7422 ( .A1(n9578), .A2(n9579), .ZN(n14350) );
  XNOR2_X1 U7423 ( .A(n9194), .B(n9193), .ZN(n11592) );
  XNOR2_X1 U7424 ( .A(n8439), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8449) );
  NAND2_X1 U7425 ( .A1(n8630), .A2(SI_8_), .ZN(n7501) );
  XNOR2_X1 U7426 ( .A(n9207), .B(n9206), .ZN(n9641) );
  OAI21_X1 U7427 ( .B1(n9479), .B2(n6901), .A(n6900), .ZN(n8354) );
  OR2_X1 U7428 ( .A1(n9205), .A2(n9192), .ZN(n9207) );
  NAND2_X1 U7429 ( .A1(n9152), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U7430 ( .A1(n8444), .A2(n8443), .ZN(n11586) );
  NAND2_X1 U7431 ( .A1(n6930), .A2(n7895), .ZN(n7936) );
  NAND2_X1 U7432 ( .A1(n6911), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U7433 ( .A1(n6919), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U7434 ( .A1(n8204), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6610) );
  MUX2_X1 U7435 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8442), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8444) );
  NOR2_X1 U7436 ( .A1(n9575), .A2(n9189), .ZN(n9577) );
  AND2_X1 U7437 ( .A1(n7579), .A2(n7655), .ZN(n7310) );
  AND2_X1 U7438 ( .A1(n6452), .A2(n8426), .ZN(n7463) );
  XNOR2_X1 U7439 ( .A(n7720), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10317) );
  AND2_X1 U7440 ( .A1(n8424), .A2(n6544), .ZN(n7269) );
  OAI21_X1 U7441 ( .B1(n7721), .B2(n6691), .A(n7738), .ZN(n6690) );
  INV_X2 U7442 ( .A(n6437), .ZN(n6439) );
  AND2_X1 U7443 ( .A1(n7581), .A2(n7580), .ZN(n7579) );
  OAI211_X1 U7444 ( .C1(n7707), .C2(n7176), .A(n7708), .B(n7175), .ZN(n10255)
         );
  NAND2_X1 U7445 ( .A1(n6630), .A2(n6629), .ZN(n7689) );
  AND2_X1 U7446 ( .A1(n6494), .A2(n9181), .ZN(n6767) );
  AND2_X1 U7447 ( .A1(n7582), .A2(n7670), .ZN(n7581) );
  AND2_X1 U7448 ( .A1(n9224), .A2(n9176), .ZN(n7355) );
  AND2_X1 U7449 ( .A1(n9209), .A2(n6768), .ZN(n6765) );
  AND4_X1 U7450 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n9149), .ZN(n8424)
         );
  AND2_X1 U7451 ( .A1(n8233), .A2(n7669), .ZN(n7582) );
  NAND2_X1 U7452 ( .A1(n9188), .A2(n9187), .ZN(n9189) );
  INV_X4 U7453 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7454 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7661) );
  INV_X1 U7455 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7577) );
  INV_X4 U7456 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7457 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n7234) );
  INV_X1 U7458 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7660) );
  NOR2_X1 U7459 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7233) );
  NOR2_X1 U7460 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7232) );
  NOR3_X1 U7461 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .A3(
        P2_IR_REG_16__SCAN_IN), .ZN(n8420) );
  NOR2_X1 U7462 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n7015) );
  NOR2_X1 U7463 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7016) );
  NOR2_X1 U7464 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7017) );
  INV_X1 U7465 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8436) );
  INV_X1 U7466 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6738) );
  OR2_X4 U7467 ( .A1(n9109), .A2(n7348), .ZN(n8728) );
  AND3_X1 U7468 ( .A1(n13216), .A2(n13215), .A3(n13214), .ZN(n13466) );
  NOR2_X2 U7469 ( .A1(n14269), .A2(n14073), .ZN(n14055) );
  NOR2_X2 U7470 ( .A1(n13376), .A2(n13522), .ZN(n6887) );
  CLKBUF_X1 U7471 ( .A(n9641), .Z(n6440) );
  NOR2_X2 U7472 ( .A1(n13304), .A2(n13492), .ZN(n6889) );
  NAND2_X1 U7474 ( .A1(n8493), .A2(n6439), .ZN(n9099) );
  NOR2_X2 U7475 ( .A1(n8562), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8564) );
  XNOR2_X2 U7476 ( .A(n8428), .B(n8427), .ZN(n13579) );
  INV_X1 U7477 ( .A(n7678), .ZN(n7676) );
  OR2_X1 U7478 ( .A1(n12213), .A2(n12478), .ZN(n11751) );
  NAND2_X1 U7479 ( .A1(n13458), .A2(n9108), .ZN(n9121) );
  NAND2_X1 U7480 ( .A1(n13213), .A2(n7153), .ZN(n7152) );
  NOR2_X1 U7481 ( .A1(n13462), .A2(n13472), .ZN(n7153) );
  INV_X1 U7482 ( .A(n7069), .ZN(n7067) );
  OR2_X1 U7483 ( .A1(n14100), .A2(n13862), .ZN(n9628) );
  NAND2_X1 U7484 ( .A1(n9019), .A2(n9018), .ZN(n9035) );
  NAND2_X1 U7485 ( .A1(n8411), .A2(SI_24_), .ZN(n8414) );
  NAND2_X1 U7486 ( .A1(n6842), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7157) );
  INV_X1 U7487 ( .A(n10578), .ZN(n6842) );
  NAND2_X1 U7488 ( .A1(n7348), .A2(n7347), .ZN(n7346) );
  NOR2_X1 U7489 ( .A1(n9693), .A2(n10655), .ZN(n7347) );
  INV_X1 U7490 ( .A(n13301), .ZN(n13040) );
  AOI21_X1 U7491 ( .B1(n7249), .B2(n7251), .A(n7248), .ZN(n7247) );
  NOR2_X1 U7492 ( .A1(n13234), .A2(n13073), .ZN(n7248) );
  NAND2_X1 U7493 ( .A1(n6704), .A2(n12102), .ZN(n13363) );
  NAND2_X1 U7494 ( .A1(n6700), .A2(n6458), .ZN(n6704) );
  NOR2_X1 U7495 ( .A1(n11874), .A2(n11875), .ZN(n7609) );
  NAND2_X1 U7496 ( .A1(n11899), .A2(n14235), .ZN(n7595) );
  MUX2_X1 U7497 ( .A(n14405), .B(n11898), .S(n11903), .Z(n11899) );
  NAND2_X1 U7498 ( .A1(n6810), .A2(n6963), .ZN(n11931) );
  INV_X1 U7499 ( .A(n6964), .ZN(n6963) );
  NAND2_X1 U7500 ( .A1(n6812), .A2(n6811), .ZN(n6810) );
  OAI21_X1 U7501 ( .B1(n11928), .B2(n14147), .A(n11927), .ZN(n6964) );
  NAND2_X1 U7502 ( .A1(n11814), .A2(n11813), .ZN(n11947) );
  NAND2_X1 U7503 ( .A1(n14274), .A2(n6435), .ZN(n11814) );
  INV_X1 U7504 ( .A(n12074), .ZN(n7458) );
  NOR2_X1 U7505 ( .A1(n12070), .A2(n7059), .ZN(n7058) );
  INV_X1 U7506 ( .A(n12069), .ZN(n7059) );
  NOR2_X1 U7507 ( .A1(n14147), .A2(n7604), .ZN(n7603) );
  INV_X1 U7508 ( .A(n11817), .ZN(n7604) );
  NAND2_X1 U7509 ( .A1(n6622), .A2(n6621), .ZN(n8411) );
  NAND2_X1 U7510 ( .A1(n6623), .A2(n7495), .ZN(n6622) );
  AOI21_X1 U7511 ( .B1(n8741), .B2(n7480), .A(n7479), .ZN(n7478) );
  INV_X1 U7512 ( .A(n8379), .ZN(n7480) );
  INV_X1 U7513 ( .A(n8383), .ZN(n7479) );
  INV_X1 U7514 ( .A(n7499), .ZN(n7498) );
  NOR2_X1 U7515 ( .A1(n8249), .A2(n8250), .ZN(n8251) );
  INV_X1 U7516 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U7517 ( .A1(n12525), .A2(n12536), .ZN(n11629) );
  NAND2_X1 U7518 ( .A1(n6521), .A2(n8181), .ZN(n7306) );
  OR2_X1 U7519 ( .A1(n12540), .A2(n12549), .ZN(n8078) );
  OR2_X1 U7520 ( .A1(n12298), .A2(n12564), .ZN(n11731) );
  OR2_X1 U7521 ( .A1(n12837), .A2(n12659), .ZN(n11704) );
  NAND2_X1 U7522 ( .A1(n8171), .A2(n12309), .ZN(n7275) );
  INV_X1 U7523 ( .A(n12909), .ZN(n7330) );
  NAND2_X1 U7524 ( .A1(n7328), .A2(n7330), .ZN(n7326) );
  INV_X1 U7525 ( .A(n9014), .ZN(n7550) );
  INV_X1 U7526 ( .A(n9013), .ZN(n7552) );
  NAND2_X1 U7527 ( .A1(n6978), .A2(n6977), .ZN(n6976) );
  NAND2_X1 U7528 ( .A1(n6482), .A2(n6979), .ZN(n6977) );
  NAND2_X1 U7529 ( .A1(n9086), .A2(n9084), .ZN(n9085) );
  INV_X1 U7530 ( .A(n8467), .ZN(n8465) );
  NOR2_X1 U7531 ( .A1(n12107), .A2(n7259), .ZN(n7258) );
  INV_X1 U7532 ( .A(n12106), .ZN(n7259) );
  INV_X1 U7533 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7230) );
  NOR2_X1 U7534 ( .A1(n11272), .A2(n7375), .ZN(n7374) );
  INV_X1 U7535 ( .A(n11125), .ZN(n7375) );
  XNOR2_X1 U7536 ( .A(n11268), .B(n10692), .ZN(n11275) );
  INV_X1 U7537 ( .A(n11592), .ZN(n9195) );
  NAND2_X1 U7538 ( .A1(n14264), .A2(n13786), .ZN(n7069) );
  NAND2_X1 U7539 ( .A1(n14065), .A2(n7431), .ZN(n7430) );
  INV_X1 U7540 ( .A(n7654), .ZN(n7431) );
  NAND2_X1 U7541 ( .A1(n13650), .A2(n14144), .ZN(n7605) );
  INV_X1 U7542 ( .A(n14293), .ZN(n13650) );
  NAND2_X1 U7543 ( .A1(n14708), .A2(n9263), .ZN(n6781) );
  NAND2_X1 U7544 ( .A1(n10558), .A2(n6783), .ZN(n6782) );
  NOR2_X1 U7545 ( .A1(n9614), .A2(n6784), .ZN(n6783) );
  INV_X1 U7546 ( .A(n9613), .ZN(n6784) );
  OR2_X1 U7547 ( .A1(n13872), .A2(n14692), .ZN(n9610) );
  NAND2_X1 U7548 ( .A1(n9634), .A2(n14071), .ZN(n14073) );
  INV_X1 U7549 ( .A(n14084), .ZN(n7432) );
  NAND2_X1 U7550 ( .A1(n7093), .A2(n9491), .ZN(n14085) );
  NAND2_X1 U7551 ( .A1(n14094), .A2(n9490), .ZN(n7093) );
  NAND2_X1 U7552 ( .A1(n7483), .A2(SI_18_), .ZN(n7026) );
  NOR2_X1 U7553 ( .A1(n7483), .A2(SI_18_), .ZN(n7025) );
  NOR2_X1 U7554 ( .A1(n8696), .A2(n6620), .ZN(n6619) );
  INV_X1 U7555 ( .A(n8369), .ZN(n6620) );
  NOR2_X1 U7556 ( .A1(n12322), .A2(n7205), .ZN(n7204) );
  NOR2_X1 U7557 ( .A1(n12240), .A2(n7207), .ZN(n7205) );
  AND2_X1 U7558 ( .A1(n10538), .A2(n10537), .ZN(n7190) );
  OR2_X1 U7559 ( .A1(n10539), .A2(n11787), .ZN(n7191) );
  OAI21_X1 U7560 ( .B1(n10902), .B2(n6758), .A(n6756), .ZN(n7209) );
  INV_X1 U7561 ( .A(n6757), .ZN(n6756) );
  OAI21_X1 U7562 ( .B1(n6759), .B2(n6758), .A(n11038), .ZN(n6757) );
  INV_X1 U7563 ( .A(n11005), .ZN(n6758) );
  NAND2_X1 U7564 ( .A1(n6694), .A2(n6692), .ZN(n11757) );
  NAND2_X1 U7565 ( .A1(n11756), .A2(n6693), .ZN(n6692) );
  OAI21_X1 U7566 ( .B1(n11752), .B2(n6695), .A(n11784), .ZN(n6694) );
  INV_X1 U7567 ( .A(n11783), .ZN(n6693) );
  NAND2_X1 U7568 ( .A1(n6735), .A2(n7676), .ZN(n6734) );
  OAI21_X1 U7569 ( .B1(n7677), .B2(n7702), .A(n6736), .ZN(n6735) );
  NAND2_X1 U7570 ( .A1(n7677), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n6736) );
  NAND2_X1 U7571 ( .A1(n7157), .A2(n6504), .ZN(n7156) );
  INV_X1 U7572 ( .A(n6933), .ZN(n10778) );
  NOR2_X1 U7573 ( .A1(n11082), .A2(n7844), .ZN(n11242) );
  NOR2_X1 U7574 ( .A1(n6675), .A2(n12402), .ZN(n6669) );
  NOR2_X1 U7575 ( .A1(n12432), .A2(n6932), .ZN(n12434) );
  NOR2_X1 U7576 ( .A1(n12449), .A2(n12637), .ZN(n6932) );
  OR2_X1 U7577 ( .A1(n14431), .A2(n14432), .ZN(n6850) );
  AND2_X1 U7578 ( .A1(n6850), .A2(n6471), .ZN(n14448) );
  OAI21_X1 U7579 ( .B1(n9671), .B2(n9670), .A(n11751), .ZN(n11593) );
  OAI21_X1 U7580 ( .B1(n12525), .B2(n12536), .A(n11629), .ZN(n12521) );
  AND4_X1 U7581 ( .A1(n8017), .A2(n8016), .A3(n8015), .A4(n8014), .ZN(n12563)
         );
  NAND2_X1 U7582 ( .A1(n7985), .A2(n7013), .ZN(n7012) );
  NOR2_X1 U7583 ( .A1(n8006), .A2(n7014), .ZN(n7013) );
  INV_X1 U7584 ( .A(n11711), .ZN(n7014) );
  NAND2_X1 U7585 ( .A1(n12658), .A2(n12657), .ZN(n12656) );
  AOI21_X1 U7586 ( .B1(n7009), .B2(n7568), .A(n11674), .ZN(n7008) );
  INV_X1 U7587 ( .A(n10515), .ZN(n11639) );
  INV_X1 U7588 ( .A(n12459), .ZN(n11785) );
  NAND2_X1 U7589 ( .A1(n9677), .A2(n11628), .ZN(n15072) );
  INV_X1 U7590 ( .A(n6441), .ZN(n7995) );
  INV_X1 U7591 ( .A(n8027), .ZN(n11616) );
  AND2_X1 U7592 ( .A1(n10344), .A2(n9692), .ZN(n10358) );
  AND3_X1 U7593 ( .A1(n8134), .A2(n7310), .A3(n7309), .ZN(n7674) );
  AND2_X1 U7594 ( .A1(n7684), .A2(n7671), .ZN(n7309) );
  NAND2_X1 U7595 ( .A1(n8022), .A2(n7407), .ZN(n8040) );
  INV_X1 U7596 ( .A(n7413), .ZN(n7412) );
  OAI21_X1 U7597 ( .B1(n7972), .B2(n7414), .A(n7989), .ZN(n7413) );
  AND2_X1 U7598 ( .A1(n7931), .A2(n7917), .ZN(n7929) );
  NOR2_X1 U7599 ( .A1(n7417), .A2(n7872), .ZN(n7416) );
  AND2_X1 U7600 ( .A1(n10004), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7872) );
  INV_X1 U7601 ( .A(n7856), .ZN(n7417) );
  AND2_X1 U7602 ( .A1(n7876), .A2(n7217), .ZN(n7216) );
  INV_X1 U7603 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7217) );
  AND2_X1 U7604 ( .A1(n9860), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7790) );
  INV_X1 U7605 ( .A(n7323), .ZN(n7322) );
  NAND2_X1 U7606 ( .A1(n13036), .A2(n6502), .ZN(n12905) );
  OR2_X1 U7607 ( .A1(n12946), .A2(n12950), .ZN(n6940) );
  OR2_X1 U7608 ( .A1(n7468), .A2(n13226), .ZN(n7467) );
  NAND2_X1 U7609 ( .A1(n6531), .A2(n12115), .ZN(n7251) );
  AOI21_X1 U7610 ( .B1(n13296), .B2(n12079), .A(n6444), .ZN(n7438) );
  NAND2_X1 U7611 ( .A1(n13373), .A2(n12067), .ZN(n7461) );
  AOI21_X1 U7612 ( .B1(n6446), .B2(n6703), .A(n6558), .ZN(n6702) );
  INV_X1 U7613 ( .A(n13415), .ZN(n6703) );
  NAND2_X1 U7614 ( .A1(n11382), .A2(n6505), .ZN(n11457) );
  INV_X1 U7615 ( .A(n11451), .ZN(n7045) );
  OR2_X1 U7616 ( .A1(n9834), .A2(n8518), .ZN(n8545) );
  NAND2_X1 U7617 ( .A1(n9158), .A2(n9159), .ZN(n14885) );
  OR2_X1 U7618 ( .A1(n9693), .A2(n13188), .ZN(n10302) );
  NAND2_X1 U7619 ( .A1(n11591), .A2(n9100), .ZN(n6627) );
  AOI21_X1 U7620 ( .B1(n13607), .B2(n13606), .A(n7356), .ZN(n13719) );
  AND2_X1 U7621 ( .A1(n13604), .A2(n13605), .ZN(n7356) );
  NOR2_X1 U7622 ( .A1(n7372), .A2(n15305), .ZN(n7370) );
  INV_X1 U7623 ( .A(n11802), .ZN(n9637) );
  AOI21_X1 U7624 ( .B1(n7102), .B2(n7098), .A(n6445), .ZN(n7097) );
  INV_X1 U7625 ( .A(n7105), .ZN(n7098) );
  NAND2_X1 U7626 ( .A1(n11174), .A2(n9335), .ZN(n11347) );
  AND2_X1 U7627 ( .A1(n11998), .A2(n9619), .ZN(n7614) );
  AND2_X1 U7628 ( .A1(n14613), .A2(n9293), .ZN(n11995) );
  INV_X1 U7629 ( .A(n9863), .ZN(n9445) );
  OR2_X1 U7630 ( .A1(n7181), .A2(n14030), .ZN(n7648) );
  AND2_X1 U7631 ( .A1(n7063), .A2(n7065), .ZN(n6935) );
  AND2_X1 U7632 ( .A1(n9635), .A2(n13985), .ZN(n14245) );
  NAND2_X1 U7633 ( .A1(n7504), .A2(n7508), .ZN(n9094) );
  INV_X1 U7634 ( .A(n7509), .ZN(n7508) );
  OAI21_X1 U7635 ( .B1(n7511), .B2(n7510), .A(n9052), .ZN(n7509) );
  NAND2_X1 U7636 ( .A1(n7487), .A2(n7486), .ZN(n6614) );
  NAND2_X1 U7637 ( .A1(n7487), .A2(n7485), .ZN(n6613) );
  NAND2_X1 U7638 ( .A1(n7515), .A2(n7072), .ZN(n8913) );
  AND2_X1 U7639 ( .A1(n6867), .A2(n6496), .ZN(n8314) );
  AOI21_X1 U7640 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n11074), .A(n8267), .ZN(
        n8281) );
  NOR2_X1 U7641 ( .A1(n8324), .A2(n8323), .ZN(n8267) );
  INV_X1 U7642 ( .A(n14428), .ZN(n7219) );
  OR2_X1 U7643 ( .A1(n12916), .A2(n12917), .ZN(n6636) );
  INV_X1 U7644 ( .A(n6634), .ZN(n6633) );
  OAI22_X1 U7645 ( .A1(n9823), .A2(n9099), .B1(n8518), .B2(n9836), .ZN(n6634)
         );
  NOR2_X1 U7646 ( .A1(n14385), .A2(n14384), .ZN(n14383) );
  NOR2_X1 U7647 ( .A1(n14397), .A2(n14398), .ZN(n14396) );
  INV_X1 U7648 ( .A(n8330), .ZN(n6902) );
  AND2_X1 U7649 ( .A1(n14588), .A2(n7219), .ZN(n6879) );
  INV_X1 U7650 ( .A(n8589), .ZN(n7540) );
  OR2_X1 U7651 ( .A1(n8552), .A2(n8551), .ZN(n8572) );
  AND2_X1 U7652 ( .A1(n8571), .A2(n8570), .ZN(n6995) );
  AOI21_X1 U7653 ( .B1(n7616), .B2(n7618), .A(n7615), .ZN(n11850) );
  NOR2_X1 U7654 ( .A1(n11845), .A2(n11846), .ZN(n7615) );
  AND2_X1 U7655 ( .A1(n7617), .A2(n11843), .ZN(n7616) );
  INV_X1 U7656 ( .A(n8629), .ZN(n6987) );
  AND2_X1 U7657 ( .A1(n8607), .A2(n8629), .ZN(n6986) );
  NAND2_X1 U7658 ( .A1(n6532), .A2(n7607), .ZN(n7606) );
  OR2_X1 U7659 ( .A1(n11879), .A2(n11878), .ZN(n11880) );
  NAND2_X1 U7660 ( .A1(n7538), .A2(n6557), .ZN(n7537) );
  INV_X1 U7661 ( .A(n8694), .ZN(n6990) );
  NAND2_X1 U7662 ( .A1(n7595), .A2(n6481), .ZN(n7586) );
  INV_X1 U7663 ( .A(n11901), .ZN(n7592) );
  NOR2_X1 U7664 ( .A1(n7590), .A2(n11894), .ZN(n7589) );
  AND2_X1 U7665 ( .A1(n11902), .A2(n6435), .ZN(n7593) );
  NOR2_X1 U7666 ( .A1(n8761), .A2(n6968), .ZN(n6967) );
  INV_X1 U7667 ( .A(n7532), .ZN(n6968) );
  AND2_X1 U7668 ( .A1(n8738), .A2(n8739), .ZN(n7535) );
  NAND2_X1 U7669 ( .A1(n7531), .A2(n8761), .ZN(n7530) );
  NAND2_X1 U7670 ( .A1(n7535), .A2(n7532), .ZN(n7531) );
  NAND2_X1 U7671 ( .A1(n7534), .A2(n7533), .ZN(n7532) );
  INV_X1 U7672 ( .A(n8738), .ZN(n7533) );
  INV_X1 U7673 ( .A(n8739), .ZN(n7534) );
  NAND2_X1 U7674 ( .A1(n6836), .A2(n11936), .ZN(n6835) );
  OR2_X1 U7675 ( .A1(n11935), .A2(n7639), .ZN(n7637) );
  NAND2_X1 U7676 ( .A1(n7639), .A2(n11935), .ZN(n7636) );
  NOR2_X1 U7677 ( .A1(n6836), .A2(n11936), .ZN(n6837) );
  AND2_X1 U7678 ( .A1(n8950), .A2(n8951), .ZN(n7529) );
  NAND2_X1 U7679 ( .A1(n7528), .A2(n7527), .ZN(n7526) );
  INV_X1 U7680 ( .A(n8950), .ZN(n7527) );
  INV_X1 U7681 ( .A(n8951), .ZN(n7528) );
  OAI22_X1 U7682 ( .A1(n11946), .A2(n6839), .B1(n11947), .B2(n6838), .ZN(
        n11949) );
  NOR2_X1 U7683 ( .A1(n11945), .A2(n6840), .ZN(n6839) );
  INV_X1 U7684 ( .A(n11945), .ZN(n6838) );
  NOR2_X1 U7685 ( .A1(n11951), .A2(n11948), .ZN(n7628) );
  INV_X1 U7686 ( .A(n7501), .ZN(n7500) );
  AOI21_X1 U7687 ( .B1(n7398), .B2(n7396), .A(n11780), .ZN(n11755) );
  INV_X1 U7688 ( .A(n11746), .ZN(n7397) );
  OR2_X1 U7689 ( .A1(n11050), .A2(n6609), .ZN(n11657) );
  NOR2_X1 U7690 ( .A1(n7458), .A2(n7057), .ZN(n7056) );
  INV_X1 U7691 ( .A(n13347), .ZN(n7057) );
  INV_X1 U7692 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9402) );
  OAI21_X1 U7693 ( .B1(n9479), .B2(n6626), .A(n6625), .ZN(n6624) );
  NAND2_X1 U7694 ( .A1(n9479), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U7695 ( .A1(n7503), .A2(n15221), .ZN(n7502) );
  INV_X1 U7696 ( .A(n8630), .ZN(n7503) );
  NAND2_X1 U7697 ( .A1(n6696), .A2(n11781), .ZN(n6695) );
  NAND2_X1 U7698 ( .A1(n11755), .A2(n11754), .ZN(n6696) );
  NAND2_X1 U7699 ( .A1(n10281), .A2(n10280), .ZN(n10318) );
  NAND2_X1 U7700 ( .A1(n7173), .A2(n10483), .ZN(n7172) );
  OAI21_X1 U7701 ( .B1(n15018), .B2(n11070), .A(n15003), .ZN(n11254) );
  OAI21_X1 U7702 ( .B1(n11480), .B2(n11257), .A(n11479), .ZN(n12375) );
  NOR2_X1 U7703 ( .A1(n12453), .A2(n12435), .ZN(n7170) );
  OR2_X1 U7704 ( .A1(n12496), .A2(n12507), .ZN(n11740) );
  INV_X1 U7705 ( .A(n12560), .ZN(n7308) );
  INV_X1 U7706 ( .A(n7000), .ZN(n6605) );
  INV_X1 U7707 ( .A(n7289), .ZN(n7288) );
  OAI21_X1 U7708 ( .B1(n8168), .B2(n7290), .A(n11674), .ZN(n7289) );
  INV_X1 U7709 ( .A(n8170), .ZN(n7290) );
  OR2_X1 U7710 ( .A1(n12688), .A2(n14473), .ZN(n11684) );
  NAND2_X1 U7711 ( .A1(n11305), .A2(n8164), .ZN(n7291) );
  NAND2_X1 U7712 ( .A1(n11050), .A2(n6609), .ZN(n11661) );
  INV_X1 U7713 ( .A(n11632), .ZN(n7572) );
  NAND2_X1 U7714 ( .A1(n15068), .A2(n12780), .ZN(n11632) );
  INV_X1 U7715 ( .A(n15068), .ZN(n6912) );
  INV_X1 U7716 ( .A(n11793), .ZN(n8151) );
  NAND2_X1 U7717 ( .A1(n8134), .A2(n7310), .ZN(n8204) );
  INV_X1 U7718 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U7719 ( .A1(n6687), .A2(n8066), .ZN(n8067) );
  NAND2_X1 U7720 ( .A1(n8065), .A2(n8064), .ZN(n6687) );
  NAND2_X1 U7721 ( .A1(n6686), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8080) );
  INV_X1 U7722 ( .A(n8067), .ZN(n6686) );
  NAND2_X1 U7723 ( .A1(n6699), .A2(n7410), .ZN(n8020) );
  AOI21_X1 U7724 ( .B1(n7412), .B2(n7414), .A(n7411), .ZN(n7410) );
  NAND2_X1 U7725 ( .A1(n7973), .A2(n7412), .ZN(n6699) );
  INV_X1 U7726 ( .A(n8008), .ZN(n7411) );
  NOR2_X1 U7727 ( .A1(n7936), .A2(n7935), .ZN(n7956) );
  INV_X1 U7728 ( .A(n7890), .ZN(n7418) );
  INV_X1 U7729 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7824) );
  INV_X1 U7730 ( .A(n7405), .ZN(n7404) );
  OAI21_X1 U7731 ( .B1(n7805), .B2(n7406), .A(n7822), .ZN(n7405) );
  INV_X1 U7732 ( .A(n7808), .ZN(n7406) );
  INV_X1 U7733 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U7734 ( .A1(n9111), .A2(n13097), .ZN(n7474) );
  AOI21_X1 U7735 ( .B1(n11204), .B2(P2_REG1_REG_14__SCAN_IN), .A(n11203), .ZN(
        n11205) );
  OR2_X1 U7736 ( .A1(n8940), .A2(n13037), .ZN(n8960) );
  INV_X1 U7737 ( .A(n7457), .ZN(n7456) );
  OAI21_X1 U7738 ( .B1(n7459), .B2(n7458), .A(n12075), .ZN(n7457) );
  NOR2_X1 U7739 ( .A1(n7041), .A2(n13439), .ZN(n7038) );
  INV_X1 U7740 ( .A(n7042), .ZN(n7041) );
  AOI21_X1 U7741 ( .B1(n7455), .B2(n14494), .A(n13442), .ZN(n7454) );
  XNOR2_X1 U7742 ( .A(n11232), .B(n13108), .ZN(n11155) );
  AND2_X1 U7743 ( .A1(n7445), .A2(n14856), .ZN(n7442) );
  NAND2_X1 U7744 ( .A1(n7449), .A2(n7450), .ZN(n7448) );
  AND2_X1 U7745 ( .A1(n12083), .A2(n7022), .ZN(n7021) );
  NAND2_X1 U7746 ( .A1(n13226), .A2(n7023), .ZN(n7022) );
  INV_X1 U7747 ( .A(n12082), .ZN(n7023) );
  OR2_X1 U7748 ( .A1(n13465), .A2(n12926), .ZN(n12084) );
  NOR2_X1 U7749 ( .A1(n6789), .A2(n11128), .ZN(n11271) );
  INV_X1 U7750 ( .A(n13774), .ZN(n7364) );
  AOI22_X1 U7751 ( .A1(n13873), .A2(n10426), .B1(n9212), .B2(n13699), .ZN(
        n10431) );
  OAI21_X1 U7752 ( .B1(n11964), .B2(n6830), .A(n6828), .ZN(n11972) );
  AOI21_X1 U7753 ( .B1(n6831), .B2(n6829), .A(n6449), .ZN(n6828) );
  NOR2_X1 U7754 ( .A1(n6510), .A2(n6831), .ZN(n6830) );
  OR2_X1 U7755 ( .A1(n9520), .A2(n10761), .ZN(n9200) );
  AND2_X1 U7756 ( .A1(n6959), .A2(n14084), .ZN(n6771) );
  AND2_X1 U7757 ( .A1(n12009), .A2(n6495), .ZN(n6772) );
  AND2_X1 U7758 ( .A1(n14117), .A2(n13863), .ZN(n7596) );
  NOR2_X1 U7759 ( .A1(n14126), .A2(n7601), .ZN(n7600) );
  INV_X1 U7760 ( .A(n11926), .ZN(n7601) );
  NOR2_X1 U7761 ( .A1(n9441), .A2(n7103), .ZN(n7102) );
  INV_X1 U7762 ( .A(n9431), .ZN(n7103) );
  NAND2_X1 U7763 ( .A1(n6936), .A2(n10751), .ZN(n11824) );
  AND2_X2 U7764 ( .A1(n11970), .A2(n11981), .ZN(n11823) );
  NAND2_X1 U7765 ( .A1(n14159), .A2(n7603), .ZN(n7602) );
  NAND2_X1 U7766 ( .A1(n6763), .A2(n9622), .ZN(n14401) );
  NOR2_X1 U7767 ( .A1(n9067), .A2(n7512), .ZN(n7511) );
  INV_X1 U7768 ( .A(n9037), .ZN(n7512) );
  INV_X1 U7769 ( .A(n9041), .ZN(n7510) );
  INV_X1 U7770 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9188) );
  INV_X1 U7771 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9187) );
  AOI21_X1 U7772 ( .B1(n8402), .B2(n6617), .A(n6616), .ZN(n6615) );
  INV_X1 U7773 ( .A(n8406), .ZN(n6616) );
  NOR2_X1 U7774 ( .A1(n8405), .A2(n8893), .ZN(n6617) );
  NAND2_X1 U7775 ( .A1(n8404), .A2(SI_21_), .ZN(n8406) );
  XNOR2_X1 U7776 ( .A(n8400), .B(SI_19_), .ZN(n8877) );
  NAND2_X1 U7777 ( .A1(n8398), .A2(n8397), .ZN(n8399) );
  NOR2_X1 U7778 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9178) );
  NOR2_X1 U7779 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n9177) );
  AOI21_X1 U7780 ( .B1(n6524), .B2(n7478), .A(n6464), .ZN(n7476) );
  AOI21_X1 U7781 ( .B1(n7476), .B2(n7477), .A(n7081), .ZN(n7080) );
  INV_X1 U7782 ( .A(n8390), .ZN(n7081) );
  NAND2_X1 U7783 ( .A1(n7478), .A2(n6479), .ZN(n7477) );
  AND2_X1 U7784 ( .A1(n8379), .A2(n8378), .ZN(n8718) );
  INV_X1 U7785 ( .A(n7475), .ZN(n8717) );
  AOI21_X1 U7786 ( .B1(n7089), .B2(n7092), .A(n8675), .ZN(n7088) );
  XNOR2_X1 U7787 ( .A(n6624), .B(SI_9_), .ZN(n8658) );
  OAI21_X1 U7788 ( .B1(n8364), .B2(n7091), .A(n7502), .ZN(n6728) );
  OR2_X1 U7789 ( .A1(n9296), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U7790 ( .A1(n8613), .A2(n8364), .ZN(n8366) );
  OAI21_X1 U7791 ( .B1(n6437), .B2(n8347), .A(n8346), .ZN(n8348) );
  XNOR2_X1 U7792 ( .A(n6962), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n8292) );
  INV_X1 U7793 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n6962) );
  OAI21_X1 U7794 ( .B1(n8292), .B2(n8293), .A(n8245), .ZN(n8246) );
  NAND2_X1 U7795 ( .A1(n8244), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n8245) );
  INV_X1 U7796 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8244) );
  OAI21_X1 U7797 ( .B1(n8288), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6519), .ZN(
        n6859) );
  XNOR2_X1 U7798 ( .A(n6859), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n8287) );
  OAI22_X1 U7799 ( .A1(n8306), .A2(n8257), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n8256), .ZN(n8258) );
  AND2_X1 U7800 ( .A1(n8256), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n8257) );
  INV_X1 U7801 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n8256) );
  AOI21_X1 U7802 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n8262), .A(n8261), .ZN(
        n8285) );
  NOR2_X1 U7803 ( .A1(n8313), .A2(n8312), .ZN(n8261) );
  NAND2_X1 U7804 ( .A1(n11663), .A2(n11664), .ZN(n11658) );
  OR2_X1 U7805 ( .A1(n7979), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8000) );
  AOI21_X1 U7806 ( .B1(n7200), .B2(n7202), .A(n6500), .ZN(n7198) );
  INV_X1 U7807 ( .A(n7203), .ZN(n7202) );
  INV_X1 U7808 ( .A(n12275), .ZN(n6749) );
  NOR2_X1 U7809 ( .A1(n6518), .A2(n6747), .ZN(n6746) );
  NAND2_X1 U7810 ( .A1(n12334), .A2(n12659), .ZN(n6743) );
  AND2_X1 U7811 ( .A1(n10904), .A2(n10901), .ZN(n6759) );
  INV_X1 U7812 ( .A(n6743), .ZN(n6742) );
  OR2_X1 U7813 ( .A1(n12334), .A2(n12659), .ZN(n6744) );
  NAND2_X1 U7814 ( .A1(n7883), .A2(n11483), .ZN(n7906) );
  INV_X1 U7815 ( .A(n11536), .ZN(n6755) );
  INV_X1 U7816 ( .A(n7213), .ZN(n7212) );
  OAI21_X1 U7817 ( .B1(n7215), .B2(n7214), .A(n12133), .ZN(n7213) );
  INV_X1 U7818 ( .A(n12138), .ZN(n6751) );
  AND3_X1 U7819 ( .A1(n7863), .A2(n6566), .A3(n7862), .ZN(n12302) );
  OR2_X1 U7820 ( .A1(n7906), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7923) );
  AOI22_X1 U7821 ( .A1(n12461), .A2(n11624), .B1(n11623), .B2(n12348), .ZN(
        n11783) );
  OAI21_X1 U7822 ( .B1(n6433), .B2(n10188), .A(n7645), .ZN(n10189) );
  NAND2_X1 U7823 ( .A1(n10260), .A2(n10261), .ZN(n10281) );
  XNOR2_X1 U7824 ( .A(n10318), .B(n10317), .ZN(n10282) );
  NAND2_X1 U7825 ( .A1(n10282), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10320) );
  OAI21_X1 U7826 ( .B1(n10572), .B2(n7762), .A(n10571), .ZN(n10771) );
  INV_X1 U7827 ( .A(n10781), .ZN(n7155) );
  NAND2_X1 U7828 ( .A1(n14985), .A2(n14986), .ZN(n15013) );
  NOR2_X1 U7829 ( .A1(n15011), .A2(n15012), .ZN(n6681) );
  NOR2_X1 U7830 ( .A1(n15011), .A2(n6683), .ZN(n6682) );
  INV_X1 U7831 ( .A(n14986), .ZN(n6683) );
  INV_X1 U7832 ( .A(n11245), .ZN(n7159) );
  NAND2_X1 U7833 ( .A1(n6858), .A2(n12370), .ZN(n7158) );
  NAND2_X1 U7834 ( .A1(n7158), .A2(n12398), .ZN(n12409) );
  NAND2_X1 U7835 ( .A1(n6671), .A2(n14391), .ZN(n6670) );
  NAND2_X1 U7836 ( .A1(n12400), .A2(n6672), .ZN(n6668) );
  NOR2_X1 U7837 ( .A1(n6673), .A2(n14391), .ZN(n6672) );
  INV_X1 U7838 ( .A(n12399), .ZN(n6673) );
  OR2_X1 U7839 ( .A1(n12390), .A2(n12391), .ZN(n6855) );
  NAND2_X1 U7840 ( .A1(n6938), .A2(n7561), .ZN(n12506) );
  AOI21_X1 U7841 ( .B1(n11777), .B2(n12534), .A(n7562), .ZN(n7561) );
  INV_X1 U7842 ( .A(n11629), .ZN(n7562) );
  NAND2_X1 U7843 ( .A1(n12506), .A2(n12505), .ZN(n12504) );
  AND2_X1 U7844 ( .A1(n8091), .A2(n8090), .ZN(n12519) );
  NOR2_X1 U7845 ( .A1(n12521), .A2(n12522), .ZN(n11777) );
  NAND2_X1 U7846 ( .A1(n12532), .A2(n7303), .ZN(n12520) );
  AND3_X1 U7847 ( .A1(n8077), .A2(n8076), .A3(n8075), .ZN(n12536) );
  NAND2_X1 U7848 ( .A1(n8050), .A2(n11731), .ZN(n12532) );
  AND2_X1 U7849 ( .A1(n11731), .A2(n11732), .ZN(n12551) );
  NAND2_X1 U7850 ( .A1(n7308), .A2(n7307), .ZN(n12558) );
  NAND2_X1 U7851 ( .A1(n7012), .A2(n7011), .ZN(n12580) );
  NOR2_X1 U7852 ( .A1(n12572), .A2(n8007), .ZN(n7011) );
  OR2_X1 U7853 ( .A1(n8012), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U7854 ( .A1(n7566), .A2(n7564), .ZN(n7985) );
  NOR2_X1 U7855 ( .A1(n7296), .A2(n7565), .ZN(n7564) );
  INV_X1 U7856 ( .A(n11715), .ZN(n7565) );
  NAND2_X1 U7857 ( .A1(n12611), .A2(n12610), .ZN(n7566) );
  OR2_X1 U7858 ( .A1(n12828), .A2(n12628), .ZN(n11715) );
  AND4_X1 U7859 ( .A1(n8005), .A2(n8004), .A3(n8003), .A4(n8002), .ZN(n12604)
         );
  AND4_X1 U7860 ( .A1(n7946), .A2(n7945), .A3(n7944), .A4(n7943), .ZN(n12615)
         );
  NAND2_X1 U7861 ( .A1(n12614), .A2(n12613), .ZN(n12612) );
  AND4_X1 U7862 ( .A1(n7984), .A2(n7983), .A3(n7982), .A4(n7981), .ZN(n12618)
         );
  OR2_X1 U7863 ( .A1(n7941), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7963) );
  AOI21_X1 U7864 ( .B1(n7002), .B2(n7003), .A(n7001), .ZN(n7000) );
  NOR2_X1 U7865 ( .A1(n7578), .A2(n7912), .ZN(n7002) );
  NOR2_X1 U7866 ( .A1(n6999), .A2(n7912), .ZN(n6998) );
  INV_X1 U7867 ( .A(n7003), .ZN(n6999) );
  AND2_X1 U7868 ( .A1(n12644), .A2(n7283), .ZN(n7282) );
  NAND2_X1 U7869 ( .A1(n7284), .A2(n8175), .ZN(n7283) );
  INV_X1 U7870 ( .A(n12657), .ZN(n7284) );
  INV_X1 U7871 ( .A(n8175), .ZN(n7285) );
  NAND2_X1 U7872 ( .A1(n12656), .A2(n8175), .ZN(n12645) );
  AOI21_X1 U7873 ( .B1(n7578), .B2(n7005), .A(n7004), .ZN(n7003) );
  NAND2_X1 U7874 ( .A1(n12670), .A2(n8174), .ZN(n12658) );
  OR2_X1 U7875 ( .A1(n14468), .A2(n14479), .ZN(n11687) );
  NAND2_X1 U7876 ( .A1(n12672), .A2(n12671), .ZN(n12670) );
  OAI21_X1 U7877 ( .B1(n14472), .B2(n14471), .A(n11684), .ZN(n12682) );
  NAND2_X1 U7878 ( .A1(n12682), .A2(n12683), .ZN(n12681) );
  AOI21_X1 U7879 ( .B1(n8166), .B2(n7567), .A(n7010), .ZN(n7009) );
  INV_X1 U7880 ( .A(n11673), .ZN(n7010) );
  AND2_X1 U7881 ( .A1(n11672), .A2(n11673), .ZN(n11760) );
  AND3_X1 U7882 ( .A1(n7813), .A2(n7812), .A3(n7811), .ZN(n11410) );
  NAND2_X1 U7883 ( .A1(n7558), .A2(n11661), .ZN(n6608) );
  NAND2_X1 U7884 ( .A1(n11767), .A2(n7018), .ZN(n7558) );
  NAND2_X1 U7885 ( .A1(n11653), .A2(n8160), .ZN(n7018) );
  INV_X1 U7886 ( .A(n11658), .ZN(n11763) );
  NAND2_X1 U7887 ( .A1(n8199), .A2(n11748), .ZN(n15046) );
  NAND2_X1 U7888 ( .A1(n10503), .A2(n6910), .ZN(n12777) );
  INV_X1 U7889 ( .A(n12771), .ZN(n6910) );
  NAND2_X1 U7890 ( .A1(n11599), .A2(n11598), .ZN(n11613) );
  OR2_X1 U7891 ( .A1(n7674), .A2(n7937), .ZN(n7675) );
  NAND2_X1 U7892 ( .A1(n8124), .A2(n8123), .ZN(n9654) );
  NAND2_X1 U7893 ( .A1(n6908), .A2(n6907), .ZN(n8096) );
  INV_X1 U7894 ( .A(n8093), .ZN(n6907) );
  OAI21_X1 U7895 ( .B1(n8079), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8080), .ZN(
        n8094) );
  OR2_X1 U7896 ( .A1(n8135), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n8138) );
  OR2_X1 U7897 ( .A1(n8020), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U7898 ( .A1(n8019), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8022) );
  XNOR2_X1 U7899 ( .A(n8020), .B(n11588), .ZN(n8019) );
  AND2_X1 U7900 ( .A1(n8008), .A2(n7988), .ZN(n7989) );
  INV_X1 U7901 ( .A(n7986), .ZN(n7414) );
  AND2_X1 U7902 ( .A1(n7986), .A2(n7971), .ZN(n7972) );
  NAND2_X1 U7903 ( .A1(n7970), .A2(n7969), .ZN(n7973) );
  NAND2_X1 U7904 ( .A1(n7973), .A2(n7972), .ZN(n7987) );
  NAND2_X1 U7905 ( .A1(n7953), .A2(n7952), .ZN(n7970) );
  AOI21_X1 U7906 ( .B1(n7929), .B2(n7393), .A(n7392), .ZN(n7391) );
  INV_X1 U7907 ( .A(n7931), .ZN(n7392) );
  INV_X1 U7908 ( .A(n7915), .ZN(n7393) );
  INV_X1 U7909 ( .A(n7929), .ZN(n7394) );
  NAND2_X1 U7910 ( .A1(n6697), .A2(n7900), .ZN(n7914) );
  NAND2_X1 U7911 ( .A1(n6698), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6697) );
  AND2_X1 U7912 ( .A1(n7915), .A2(n7901), .ZN(n7913) );
  INV_X1 U7913 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U7914 ( .A1(n7894), .A2(n10123), .ZN(n7900) );
  NAND2_X1 U7915 ( .A1(n7893), .A2(n7892), .ZN(n7894) );
  INV_X1 U7916 ( .A(n7667), .ZN(n7876) );
  NAND2_X1 U7917 ( .A1(n7855), .A2(n7854), .ZN(n7857) );
  XNOR2_X1 U7918 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7822) );
  INV_X1 U7919 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U7920 ( .A1(n7777), .A2(n7776), .ZN(n7791) );
  NAND2_X1 U7921 ( .A1(n7661), .A2(n7577), .ZN(n7575) );
  NAND2_X1 U7922 ( .A1(n7576), .A2(n7661), .ZN(n7733) );
  INV_X1 U7923 ( .A(n7719), .ZN(n7576) );
  NAND2_X1 U7924 ( .A1(n6738), .A2(n7176), .ZN(n7708) );
  NAND2_X1 U7925 ( .A1(n8491), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7705) );
  XNOR2_X1 U7926 ( .A(n10942), .B(n12966), .ZN(n9736) );
  AND2_X1 U7927 ( .A1(n6926), .A2(n9757), .ZN(n6653) );
  INV_X1 U7928 ( .A(n9780), .ZN(n6926) );
  INV_X1 U7929 ( .A(n13106), .ZN(n11455) );
  NAND2_X1 U7930 ( .A1(n8456), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8940) );
  INV_X1 U7931 ( .A(n8918), .ZN(n8456) );
  INV_X1 U7932 ( .A(n12894), .ZN(n7345) );
  INV_X1 U7933 ( .A(n12890), .ZN(n6639) );
  AND2_X1 U7934 ( .A1(n11151), .A2(n10927), .ZN(n6655) );
  INV_X1 U7935 ( .A(n9727), .ZN(n7324) );
  INV_X1 U7936 ( .A(n10508), .ZN(n7321) );
  NAND2_X1 U7937 ( .A1(n12976), .A2(n12899), .ZN(n12904) );
  AND2_X1 U7938 ( .A1(n6922), .A2(n12881), .ZN(n6654) );
  INV_X1 U7939 ( .A(n13061), .ZN(n6922) );
  AND2_X1 U7940 ( .A1(n13077), .A2(n12915), .ZN(n7331) );
  NAND2_X1 U7941 ( .A1(n7543), .A2(n7542), .ZN(n9051) );
  OAI22_X1 U7942 ( .A1(n6997), .A2(n6996), .B1(n7544), .B2(n7547), .ZN(n7543)
         );
  AND2_X1 U7943 ( .A1(n7548), .A2(n7549), .ZN(n7547) );
  AND2_X1 U7944 ( .A1(n6975), .A2(n6447), .ZN(n6972) );
  INV_X1 U7945 ( .A(n6976), .ZN(n6975) );
  OAI211_X1 U7946 ( .C1(n6976), .C2(n6527), .A(n7469), .B(n7472), .ZN(n6632)
         );
  NAND2_X1 U7947 ( .A1(n9116), .A2(n9092), .ZN(n7472) );
  OR2_X1 U7948 ( .A1(n9025), .A2(n10199), .ZN(n8499) );
  OR2_X1 U7949 ( .A1(n8986), .A2(n8495), .ZN(n8497) );
  INV_X1 U7950 ( .A(n13207), .ZN(n13205) );
  NOR2_X1 U7951 ( .A1(n7253), .A2(n12114), .ZN(n7252) );
  INV_X1 U7952 ( .A(n12115), .ZN(n7253) );
  INV_X1 U7953 ( .A(n12058), .ZN(n13250) );
  AND2_X1 U7954 ( .A1(n12081), .A2(n9129), .ZN(n13257) );
  NAND2_X1 U7955 ( .A1(n6889), .A2(n6888), .ZN(n13273) );
  AND2_X1 U7956 ( .A1(n7029), .A2(n6548), .ZN(n7036) );
  NAND2_X1 U7957 ( .A1(n7438), .A2(n7439), .ZN(n7029) );
  NAND2_X1 U7958 ( .A1(n13497), .A2(n12108), .ZN(n13292) );
  AOI21_X1 U7959 ( .B1(n7258), .B2(n12105), .A(n6463), .ZN(n7257) );
  NAND2_X1 U7960 ( .A1(n7437), .A2(n13310), .ZN(n13299) );
  INV_X1 U7961 ( .A(n7147), .ZN(n13320) );
  NAND2_X1 U7962 ( .A1(n6701), .A2(n6446), .ZN(n6700) );
  INV_X1 U7963 ( .A(n13416), .ZN(n6701) );
  NAND2_X1 U7964 ( .A1(n13416), .A2(n13415), .ZN(n12100) );
  OR2_X1 U7965 ( .A1(n7454), .A2(n7453), .ZN(n7452) );
  NOR2_X1 U7966 ( .A1(n14494), .A2(n7455), .ZN(n7453) );
  NAND2_X1 U7967 ( .A1(n7454), .A2(n13434), .ZN(n7451) );
  INV_X1 U7968 ( .A(n13105), .ZN(n13421) );
  NAND2_X1 U7969 ( .A1(n13440), .A2(n13451), .ZN(n12063) );
  OR2_X1 U7970 ( .A1(n11105), .A2(n11109), .ZN(n11108) );
  OR2_X1 U7971 ( .A1(n10938), .A2(n10946), .ZN(n11111) );
  NAND2_X1 U7972 ( .A1(n10937), .A2(n10936), .ZN(n10938) );
  NAND2_X1 U7973 ( .A1(n7241), .A2(n7239), .ZN(n10959) );
  NOR2_X1 U7974 ( .A1(n7447), .A2(n7240), .ZN(n7239) );
  INV_X1 U7975 ( .A(n10858), .ZN(n7240) );
  INV_X1 U7976 ( .A(n14885), .ZN(n13441) );
  NAND2_X1 U7977 ( .A1(n10398), .A2(n14879), .ZN(n10295) );
  NAND2_X1 U7978 ( .A1(n13465), .A2(n14930), .ZN(n6948) );
  NAND2_X2 U7979 ( .A1(n9022), .A2(n9021), .ZN(n13472) );
  AND2_X1 U7980 ( .A1(n9769), .A2(n9768), .ZN(n14891) );
  AND2_X1 U7981 ( .A1(n9157), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9690) );
  AND2_X1 U7982 ( .A1(n7269), .A2(n7268), .ZN(n7267) );
  INV_X1 U7983 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7268) );
  INV_X1 U7984 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9149) );
  OAI21_X1 U7985 ( .B1(n8440), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9147) );
  INV_X1 U7986 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9146) );
  AND2_X1 U7987 ( .A1(n7353), .A2(n8431), .ZN(n7352) );
  INV_X1 U7988 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8431) );
  XNOR2_X1 U7989 ( .A(n8445), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10655) );
  INV_X1 U7990 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U7991 ( .A1(n13818), .A2(n13671), .ZN(n13728) );
  INV_X1 U7992 ( .A(n14406), .ZN(n11552) );
  AND2_X1 U7993 ( .A1(n6818), .A2(n13712), .ZN(n6443) );
  OR2_X1 U7994 ( .A1(n13838), .A2(n13709), .ZN(n6818) );
  INV_X1 U7995 ( .A(n6937), .ZN(n13750) );
  OR2_X1 U7996 ( .A1(n13618), .A2(n13848), .ZN(n7384) );
  AND2_X1 U7997 ( .A1(n13618), .A2(n13848), .ZN(n7383) );
  INV_X1 U7998 ( .A(n7374), .ZN(n7367) );
  AOI21_X1 U7999 ( .B1(n13704), .B2(n13874), .A(n7386), .ZN(n10147) );
  INV_X1 U8000 ( .A(n10145), .ZN(n7386) );
  AOI21_X1 U8001 ( .B1(n13700), .B2(n10896), .A(n10144), .ZN(n10145) );
  AND2_X1 U8002 ( .A1(n13662), .A2(n13811), .ZN(n6809) );
  INV_X1 U8003 ( .A(n13648), .ZN(n6807) );
  INV_X1 U8004 ( .A(n6809), .ZN(n6808) );
  AND2_X1 U8005 ( .A1(n13820), .A2(n7361), .ZN(n7360) );
  NAND2_X1 U8006 ( .A1(n7363), .A2(n13662), .ZN(n7361) );
  NAND2_X1 U8007 ( .A1(n13837), .A2(n13838), .ZN(n13836) );
  INV_X1 U8008 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n13883) );
  NOR2_X1 U8009 ( .A1(n13991), .A2(n13985), .ZN(n13986) );
  NAND2_X1 U8010 ( .A1(n6774), .A2(n6515), .ZN(n7066) );
  NAND2_X1 U8011 ( .A1(n14032), .A2(n14033), .ZN(n14031) );
  OAI21_X1 U8012 ( .B1(n14085), .B2(n6525), .A(n7427), .ZN(n14052) );
  NAND2_X1 U8013 ( .A1(n7430), .A2(n9515), .ZN(n7427) );
  INV_X1 U8014 ( .A(n7430), .ZN(n7428) );
  AND2_X1 U8015 ( .A1(n9628), .A2(n9489), .ZN(n14103) );
  NAND2_X1 U8016 ( .A1(n14133), .A2(n6487), .ZN(n14118) );
  NOR2_X1 U8017 ( .A1(n6778), .A2(n14111), .ZN(n6777) );
  INV_X1 U8018 ( .A(n7061), .ZN(n6778) );
  OR2_X1 U8019 ( .A1(n7600), .A2(n7597), .ZN(n7061) );
  INV_X1 U8020 ( .A(n7605), .ZN(n7597) );
  NAND2_X1 U8021 ( .A1(n14159), .A2(n7598), .ZN(n6779) );
  INV_X1 U8022 ( .A(n7102), .ZN(n7099) );
  AND3_X1 U8023 ( .A1(n9456), .A2(n9455), .A3(n9454), .ZN(n14164) );
  NAND2_X1 U8024 ( .A1(n14311), .A2(n14195), .ZN(n9627) );
  NOR2_X1 U8025 ( .A1(n9430), .A2(n7106), .ZN(n7105) );
  INV_X1 U8026 ( .A(n9416), .ZN(n7106) );
  NAND2_X1 U8027 ( .A1(n14205), .A2(n6560), .ZN(n14192) );
  INV_X1 U8028 ( .A(n12004), .ZN(n14193) );
  AOI21_X1 U8029 ( .B1(n7421), .B2(n7131), .A(n9400), .ZN(n7129) );
  INV_X1 U8030 ( .A(n7131), .ZN(n7130) );
  NAND2_X1 U8031 ( .A1(n7625), .A2(n7624), .ZN(n6786) );
  AND2_X1 U8032 ( .A1(n11900), .A2(n9625), .ZN(n7624) );
  NAND2_X1 U8033 ( .A1(n6786), .A2(n6785), .ZN(n14205) );
  AND2_X1 U8034 ( .A1(n7133), .A2(n11893), .ZN(n6785) );
  AOI21_X1 U8035 ( .B1(n6453), .B2(n7119), .A(n6511), .ZN(n7115) );
  INV_X1 U8036 ( .A(n12000), .ZN(n14400) );
  NAND2_X1 U8037 ( .A1(n14554), .A2(n11552), .ZN(n7120) );
  AND4_X1 U8038 ( .A1(n9319), .A2(n9318), .A3(n9317), .A4(n9316), .ZN(n14618)
         );
  NAND2_X1 U8039 ( .A1(n6764), .A2(n11997), .ZN(n11025) );
  AND2_X1 U8040 ( .A1(n11995), .A2(n9616), .ZN(n7623) );
  NAND2_X1 U8041 ( .A1(n6782), .A2(n6781), .ZN(n14638) );
  NOR2_X1 U8042 ( .A1(n7114), .A2(n9265), .ZN(n7113) );
  INV_X1 U8043 ( .A(n9249), .ZN(n7114) );
  NAND2_X1 U8044 ( .A1(n10558), .A2(n9613), .ZN(n10639) );
  NAND2_X1 U8045 ( .A1(n9238), .A2(n9237), .ZN(n10733) );
  AND2_X1 U8046 ( .A1(n9610), .A2(n9609), .ZN(n11989) );
  AND2_X1 U8047 ( .A1(n9833), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U8048 ( .A1(n9863), .A2(n7424), .ZN(n7423) );
  NOR2_X1 U8049 ( .A1(n9836), .A2(n9479), .ZN(n7424) );
  OR2_X1 U8050 ( .A1(n11984), .A2(n13877), .ZN(n14617) );
  INV_X1 U8051 ( .A(n14403), .ZN(n14639) );
  INV_X1 U8052 ( .A(n14619), .ZN(n14127) );
  INV_X1 U8053 ( .A(n14617), .ZN(n14404) );
  INV_X1 U8054 ( .A(n13991), .ZN(n14243) );
  NAND2_X1 U8055 ( .A1(n9632), .A2(n9631), .ZN(n14403) );
  INV_X1 U8056 ( .A(n14085), .ZN(n7433) );
  NAND2_X1 U8057 ( .A1(n10151), .A2(n10150), .ZN(n14723) );
  INV_X1 U8058 ( .A(n9094), .ZN(n9058) );
  AND2_X1 U8059 ( .A1(n9206), .A2(n9203), .ZN(n7622) );
  XNOR2_X1 U8060 ( .A(n9098), .B(n9097), .ZN(n11806) );
  AND4_X1 U8061 ( .A1(n9185), .A2(n9184), .A3(n9443), .A4(n9586), .ZN(n9186)
         );
  INV_X1 U8062 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9206) );
  NAND2_X1 U8063 ( .A1(n7494), .A2(n7493), .ZN(n7492) );
  INV_X1 U8064 ( .A(n8415), .ZN(n7494) );
  INV_X1 U8065 ( .A(n8998), .ZN(n7490) );
  NAND2_X1 U8066 ( .A1(n8408), .A2(SI_22_), .ZN(n8410) );
  INV_X1 U8067 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9572) );
  INV_X1 U8068 ( .A(n6894), .ZN(n9584) );
  NAND2_X1 U8069 ( .A1(n8402), .A2(n8403), .ZN(n7515) );
  INV_X1 U8070 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9442) );
  INV_X1 U8071 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9443) );
  INV_X1 U8072 ( .A(n8855), .ZN(n7483) );
  OR2_X1 U8073 ( .A1(n8399), .A2(n10142), .ZN(n7482) );
  NAND2_X1 U8074 ( .A1(n8399), .A2(n10142), .ZN(n7484) );
  INV_X1 U8075 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9176) );
  NOR2_X2 U8076 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9209) );
  XNOR2_X1 U8077 ( .A(n8292), .B(n6950), .ZN(n8294) );
  INV_X1 U8078 ( .A(n8293), .ZN(n6950) );
  XNOR2_X1 U8079 ( .A(n8287), .B(n13935), .ZN(n8301) );
  NAND2_X1 U8080 ( .A1(n15314), .A2(n8300), .ZN(n8302) );
  INV_X1 U8081 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n13962) );
  NAND2_X1 U8082 ( .A1(n14392), .A2(n8316), .ZN(n8318) );
  OAI21_X1 U8083 ( .B1(n8266), .B2(n15023), .A(n8265), .ZN(n8324) );
  OAI21_X1 U8084 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n8269), .A(n8268), .ZN(
        n8327) );
  AND2_X1 U8085 ( .A1(n6880), .A2(n14577), .ZN(n8329) );
  OAI21_X1 U8086 ( .B1(n14578), .B2(n14579), .A(n15245), .ZN(n6880) );
  NAND2_X1 U8087 ( .A1(n8056), .A2(n8055), .ZN(n12540) );
  INV_X1 U8088 ( .A(n10598), .ZN(n7210) );
  AND2_X1 U8089 ( .A1(n6886), .A2(n10585), .ZN(n10548) );
  INV_X1 U8090 ( .A(n12353), .ZN(n12564) );
  NAND2_X1 U8091 ( .A1(n8028), .A2(n6578), .ZN(n12565) );
  NAND2_X1 U8092 ( .A1(n10902), .A2(n6759), .ZN(n11006) );
  NAND2_X1 U8093 ( .A1(n8043), .A2(n8042), .ZN(n12298) );
  INV_X1 U8094 ( .A(n12339), .ZN(n12324) );
  NAND2_X1 U8095 ( .A1(n10359), .A2(n10358), .ZN(n12332) );
  OAI21_X1 U8096 ( .B1(n11757), .B2(n10538), .A(n11790), .ZN(n6939) );
  INV_X1 U8097 ( .A(n15069), .ZN(n15048) );
  INV_X1 U8098 ( .A(n12615), .ZN(n12646) );
  XNOR2_X1 U8099 ( .A(n10256), .B(n6433), .ZN(n10258) );
  OR2_X1 U8100 ( .A1(n10373), .A2(n10372), .ZN(n6661) );
  AND2_X1 U8101 ( .A1(n6667), .A2(n6666), .ZN(n10569) );
  NAND2_X1 U8102 ( .A1(n6664), .A2(n6662), .ZN(n6667) );
  AND2_X1 U8103 ( .A1(n6847), .A2(n15019), .ZN(n6846) );
  OR2_X1 U8104 ( .A1(n6471), .A2(n6931), .ZN(n6847) );
  AND2_X1 U8105 ( .A1(n6471), .A2(n6931), .ZN(n6845) );
  XNOR2_X1 U8106 ( .A(n12446), .B(n12445), .ZN(n6657) );
  AND2_X1 U8107 ( .A1(P3_U3897), .A2(n8191), .ZN(n15015) );
  OAI211_X1 U8108 ( .C1(n14448), .C2(n7164), .A(n7161), .B(n6660), .ZN(n6659)
         );
  NAND2_X1 U8109 ( .A1(n7165), .A2(n7169), .ZN(n7164) );
  INV_X1 U8110 ( .A(n12460), .ZN(n6660) );
  AOI21_X1 U8111 ( .B1(n7299), .B2(n12476), .A(n6522), .ZN(n7297) );
  XNOR2_X1 U8112 ( .A(n11593), .B(n9673), .ZN(n12050) );
  NAND2_X1 U8113 ( .A1(n15058), .A2(n14477), .ZN(n12691) );
  AND2_X1 U8114 ( .A1(n15091), .A2(n12045), .ZN(n15059) );
  NAND2_X1 U8115 ( .A1(n7557), .A2(n15136), .ZN(n7279) );
  NAND2_X1 U8116 ( .A1(n8011), .A2(n8010), .ZN(n12815) );
  NAND2_X1 U8117 ( .A1(n7940), .A2(n7939), .ZN(n12831) );
  NAND2_X1 U8118 ( .A1(n7920), .A2(n7919), .ZN(n12837) );
  OR2_X1 U8119 ( .A1(n15137), .A2(n15111), .ZN(n12846) );
  NAND2_X1 U8120 ( .A1(n13050), .A2(n13051), .ZN(n13049) );
  NOR2_X1 U8121 ( .A1(n7338), .A2(n13082), .ZN(n7337) );
  OAI21_X1 U8122 ( .B1(n7342), .B2(n7341), .A(n7339), .ZN(n7338) );
  NAND2_X1 U8123 ( .A1(n7340), .A2(n12964), .ZN(n7339) );
  OR2_X1 U8124 ( .A1(n12920), .A2(n12968), .ZN(n7343) );
  NAND2_X1 U8125 ( .A1(n8804), .A2(n8803), .ZN(n13533) );
  NAND2_X1 U8126 ( .A1(n8787), .A2(n8786), .ZN(n13527) );
  NAND2_X1 U8127 ( .A1(n9715), .A2(n6651), .ZN(n6648) );
  INV_X1 U8128 ( .A(n13445), .ZN(n12059) );
  NAND2_X1 U8129 ( .A1(n8701), .A2(n8700), .ZN(n13549) );
  OR2_X1 U8130 ( .A1(n14349), .A2(n8518), .ZN(n8430) );
  XNOR2_X1 U8131 ( .A(n12872), .B(n12873), .ZN(n13086) );
  INV_X1 U8132 ( .A(n13082), .ZN(n13085) );
  NAND2_X1 U8133 ( .A1(n9783), .A2(n14881), .ZN(n13093) );
  NAND2_X1 U8134 ( .A1(n9029), .A2(n9028), .ZN(n13241) );
  NAND2_X1 U8135 ( .A1(n8473), .A2(n8472), .ZN(n13259) );
  NAND2_X1 U8136 ( .A1(n8992), .A2(n8991), .ZN(n13258) );
  NAND2_X1 U8137 ( .A1(n8966), .A2(n8965), .ZN(n13301) );
  INV_X1 U8138 ( .A(n12120), .ZN(n7273) );
  NAND2_X1 U8139 ( .A1(n7260), .A2(n12106), .ZN(n13319) );
  OR2_X1 U8140 ( .A1(n13330), .A2(n12105), .ZN(n7260) );
  NAND2_X1 U8141 ( .A1(n13331), .A2(n12074), .ZN(n13314) );
  NAND2_X1 U8142 ( .A1(n12073), .A2(n12072), .ZN(n13333) );
  NAND2_X1 U8143 ( .A1(n8861), .A2(n8860), .ZN(n13522) );
  INV_X1 U8144 ( .A(n14865), .ZN(n14881) );
  INV_X1 U8145 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13574) );
  AND2_X1 U8146 ( .A1(n6488), .A2(n7555), .ZN(n7554) );
  AND2_X1 U8147 ( .A1(n8461), .A2(n7556), .ZN(n7555) );
  NAND2_X1 U8148 ( .A1(n9480), .A2(n8936), .ZN(n7027) );
  INV_X1 U8149 ( .A(n10655), .ZN(n13188) );
  INV_X1 U8150 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U8151 ( .A1(n11356), .A2(n6792), .ZN(n11551) );
  NAND2_X1 U8152 ( .A1(n11355), .A2(n11354), .ZN(n6792) );
  NAND2_X1 U8153 ( .A1(n9326), .A2(n9325), .ZN(n14741) );
  NAND2_X1 U8154 ( .A1(n7371), .A2(n7369), .ZN(n15304) );
  AND2_X1 U8155 ( .A1(n11565), .A2(n11564), .ZN(n7359) );
  NAND2_X1 U8156 ( .A1(n9408), .A2(n9407), .ZN(n14518) );
  NAND2_X1 U8157 ( .A1(n6795), .A2(n10454), .ZN(n6794) );
  NAND2_X1 U8158 ( .A1(n6802), .A2(n10689), .ZN(n6799) );
  NAND2_X1 U8159 ( .A1(n11279), .A2(n11278), .ZN(n11356) );
  NAND2_X1 U8160 ( .A1(n9228), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U8161 ( .A1(n9228), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U8162 ( .A1(n9228), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U8163 ( .A1(n9228), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9501) );
  AOI21_X1 U8164 ( .B1(n9228), .B2(P1_REG0_REG_4__SCAN_IN), .A(n7135), .ZN(
        n7134) );
  OAI21_X1 U8165 ( .B1(n10615), .B2(n9520), .A(n6892), .ZN(n7135) );
  AOI21_X1 U8166 ( .B1(n14245), .B2(n14633), .A(n9650), .ZN(n9651) );
  NAND2_X1 U8167 ( .A1(n14009), .A2(n14008), .ZN(n14250) );
  OR2_X1 U8168 ( .A1(n14349), .A2(n9527), .ZN(n9529) );
  NAND2_X1 U8169 ( .A1(n9493), .A2(n9492), .ZN(n14089) );
  NAND2_X1 U8170 ( .A1(n14542), .A2(n7131), .ZN(n14207) );
  NAND2_X1 U8171 ( .A1(n9646), .A2(n14229), .ZN(n14231) );
  OAI211_X1 U8172 ( .C1(n14250), .C2(n7128), .A(n7126), .B(n7123), .ZN(n14244)
         );
  NAND2_X1 U8173 ( .A1(n12015), .A2(n7127), .ZN(n7126) );
  INV_X1 U8174 ( .A(n12015), .ZN(n7128) );
  NAND2_X1 U8175 ( .A1(n14250), .A2(n7125), .ZN(n7123) );
  NAND2_X1 U8176 ( .A1(n14751), .A2(n14748), .ZN(n7124) );
  INV_X1 U8177 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10554) );
  NAND2_X1 U8178 ( .A1(n6865), .A2(n6864), .ZN(n6863) );
  NOR2_X1 U8179 ( .A1(n8308), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U8180 ( .A1(n14383), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6860) );
  NOR2_X1 U8181 ( .A1(n14396), .A2(n8322), .ZN(n14568) );
  OR2_X1 U8182 ( .A1(n14568), .A2(n14567), .ZN(n7220) );
  AND2_X1 U8183 ( .A1(n7220), .A2(n6913), .ZN(n14570) );
  INV_X1 U8184 ( .A(n14571), .ZN(n6890) );
  NAND2_X1 U8185 ( .A1(n8329), .A2(n8328), .ZN(n14584) );
  NAND2_X1 U8186 ( .A1(n14584), .A2(n14585), .ZN(n14581) );
  NAND2_X1 U8187 ( .A1(n6915), .A2(n6914), .ZN(n14583) );
  INV_X1 U8188 ( .A(n8328), .ZN(n6914) );
  INV_X1 U8189 ( .A(n8329), .ZN(n6915) );
  NAND2_X1 U8190 ( .A1(n6874), .A2(n6873), .ZN(n6875) );
  INV_X1 U8191 ( .A(n6878), .ZN(n6873) );
  AOI21_X1 U8192 ( .B1(n6877), .B2(n6878), .A(P2_ADDR_REG_18__SCAN_IN), .ZN(
        n6868) );
  XNOR2_X1 U8193 ( .A(n8342), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n8343) );
  AOI21_X1 U8194 ( .B1(n8728), .B2(n13116), .A(n8490), .ZN(n8527) );
  AND2_X1 U8195 ( .A1(n10297), .A2(n6436), .ZN(n8490) );
  NAND2_X1 U8196 ( .A1(n7540), .A2(n6480), .ZN(n7539) );
  OR2_X1 U8197 ( .A1(n8571), .A2(n8570), .ZN(n6994) );
  NAND2_X1 U8198 ( .A1(n11874), .A2(n11875), .ZN(n7610) );
  INV_X1 U8199 ( .A(n11855), .ZN(n6825) );
  NAND2_X1 U8200 ( .A1(n11857), .A2(n14615), .ZN(n7608) );
  INV_X1 U8201 ( .A(n7609), .ZN(n7607) );
  INV_X1 U8202 ( .A(n8628), .ZN(n6988) );
  NAND2_X1 U8203 ( .A1(n11883), .A2(n7613), .ZN(n7612) );
  NAND2_X1 U8204 ( .A1(n11901), .A2(n11903), .ZN(n7590) );
  NOR2_X1 U8205 ( .A1(n8693), .A2(n6990), .ZN(n6989) );
  INV_X1 U8206 ( .A(n11896), .ZN(n7591) );
  OAI21_X1 U8207 ( .B1(n6970), .B2(n6969), .A(n6966), .ZN(n8843) );
  INV_X1 U8208 ( .A(n8760), .ZN(n6969) );
  NOR2_X1 U8209 ( .A1(n11924), .A2(n14147), .ZN(n6811) );
  OAI21_X1 U8210 ( .B1(n11931), .B2(n11930), .A(n11929), .ZN(n11933) );
  AND2_X1 U8211 ( .A1(n8909), .A2(n8910), .ZN(n7522) );
  NAND2_X1 U8212 ( .A1(n6992), .A2(n6561), .ZN(n8911) );
  NAND2_X1 U8213 ( .A1(n7521), .A2(n7520), .ZN(n7519) );
  INV_X1 U8214 ( .A(n8909), .ZN(n7520) );
  INV_X1 U8215 ( .A(n8910), .ZN(n7521) );
  AND2_X1 U8216 ( .A1(n6833), .A2(n11941), .ZN(n6832) );
  NAND2_X1 U8217 ( .A1(n6837), .A2(n6835), .ZN(n6833) );
  INV_X1 U8218 ( .A(n11941), .ZN(n6927) );
  INV_X1 U8219 ( .A(n11947), .ZN(n6840) );
  INV_X1 U8220 ( .A(n15070), .ZN(n11762) );
  NAND2_X1 U8221 ( .A1(n7400), .A2(n6492), .ZN(n7399) );
  AOI21_X1 U8222 ( .B1(n8952), .B2(n7526), .A(n7524), .ZN(n7523) );
  NAND2_X1 U8223 ( .A1(n8973), .A2(n7525), .ZN(n7524) );
  NAND2_X1 U8224 ( .A1(n7529), .A2(n7526), .ZN(n7525) );
  INV_X1 U8225 ( .A(n7628), .ZN(n7627) );
  OAI21_X1 U8226 ( .B1(n11949), .B2(n7628), .A(n7629), .ZN(n11954) );
  NAND2_X1 U8227 ( .A1(n11967), .A2(n7642), .ZN(n7641) );
  NAND2_X1 U8228 ( .A1(n7496), .A2(n10856), .ZN(n7495) );
  INV_X1 U8229 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7228) );
  INV_X1 U8230 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7229) );
  NAND2_X1 U8231 ( .A1(n11962), .A2(n11960), .ZN(n7635) );
  INV_X1 U8232 ( .A(n11967), .ZN(n7640) );
  NAND2_X1 U8233 ( .A1(n11810), .A2(n11811), .ZN(n11968) );
  AND2_X1 U8234 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9250) );
  AOI21_X1 U8235 ( .B1(n7078), .B2(n7080), .A(n7077), .ZN(n7076) );
  INV_X1 U8236 ( .A(n7651), .ZN(n7077) );
  INV_X1 U8237 ( .A(n7476), .ZN(n7078) );
  INV_X1 U8238 ( .A(n7080), .ZN(n7079) );
  INV_X1 U8239 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6768) );
  INV_X1 U8240 ( .A(n12219), .ZN(n7208) );
  AND2_X1 U8241 ( .A1(n12275), .A2(n6748), .ZN(n6747) );
  INV_X1 U8242 ( .A(n12153), .ZN(n6748) );
  AND2_X1 U8243 ( .A1(n11750), .A2(n11751), .ZN(n7395) );
  OR3_X1 U8244 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n10501), .ZN(n7645) );
  OAI21_X1 U8245 ( .B1(n10278), .B2(n10263), .A(n10277), .ZN(n10323) );
  NAND2_X1 U8246 ( .A1(n10479), .A2(n7174), .ZN(n7173) );
  INV_X1 U8247 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11483) );
  OAI21_X1 U8248 ( .B1(n12449), .B2(n12448), .A(n12447), .ZN(n12451) );
  INV_X1 U8249 ( .A(n7170), .ZN(n7168) );
  INV_X1 U8250 ( .A(n11739), .ZN(n6599) );
  OR2_X1 U8251 ( .A1(n8099), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8114) );
  NOR2_X1 U8252 ( .A1(n7563), .A2(n7560), .ZN(n7559) );
  INV_X1 U8253 ( .A(n11731), .ZN(n7560) );
  INV_X1 U8254 ( .A(n11777), .ZN(n7563) );
  NAND2_X1 U8255 ( .A1(n8072), .A2(n8071), .ZN(n8084) );
  OR2_X1 U8256 ( .A1(n8057), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8073) );
  OR2_X1 U8257 ( .A1(n12565), .A2(n12574), .ZN(n11727) );
  INV_X1 U8258 ( .A(n11760), .ZN(n8168) );
  INV_X1 U8259 ( .A(n8051), .ZN(n7409) );
  OR2_X1 U8260 ( .A1(n7809), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7820) );
  NOR2_X1 U8261 ( .A1(n8769), .A2(n15198), .ZN(n8768) );
  OAI21_X1 U8262 ( .B1(n6456), .B2(n7330), .A(n12985), .ZN(n7329) );
  OAI21_X1 U8263 ( .B1(n7545), .B2(n7549), .A(n9016), .ZN(n7541) );
  NAND2_X1 U8264 ( .A1(n7546), .A2(n9017), .ZN(n7545) );
  NAND2_X1 U8265 ( .A1(n7551), .A2(n7549), .ZN(n7546) );
  AND2_X1 U8266 ( .A1(n9013), .A2(n9014), .ZN(n7551) );
  INV_X1 U8267 ( .A(n9089), .ZN(n7470) );
  NOR2_X1 U8268 ( .A1(n9087), .A2(n9088), .ZN(n7471) );
  NOR2_X1 U8269 ( .A1(n7252), .A2(n13226), .ZN(n7249) );
  NAND2_X1 U8270 ( .A1(n7056), .A2(n7054), .ZN(n7053) );
  INV_X1 U8271 ( .A(n12071), .ZN(n7054) );
  NOR2_X1 U8272 ( .A1(n7055), .A2(n7052), .ZN(n7051) );
  INV_X1 U8273 ( .A(n7058), .ZN(n7052) );
  INV_X1 U8274 ( .A(n7056), .ZN(n7055) );
  INV_X1 U8275 ( .A(n12072), .ZN(n7460) );
  INV_X1 U8276 ( .A(n6712), .ZN(n6711) );
  OAI21_X1 U8277 ( .B1(n12103), .B2(n6472), .A(n12104), .ZN(n6712) );
  NAND2_X1 U8278 ( .A1(n8455), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8899) );
  AND2_X1 U8279 ( .A1(n8805), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8788) );
  AND2_X1 U8280 ( .A1(n8768), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8805) );
  NOR2_X1 U8281 ( .A1(n12065), .A2(n7043), .ZN(n7042) );
  INV_X1 U8282 ( .A(n7451), .ZN(n7043) );
  INV_X1 U8283 ( .A(n7452), .ZN(n7040) );
  NAND2_X1 U8284 ( .A1(n6591), .A2(n6590), .ZN(n13428) );
  INV_X1 U8285 ( .A(n13447), .ZN(n6591) );
  NAND2_X1 U8286 ( .A1(n7461), .A2(n7058), .ZN(n7060) );
  INV_X1 U8287 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6631) );
  INV_X1 U8288 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7353) );
  INV_X1 U8289 ( .A(n14514), .ZN(n7382) );
  AOI21_X1 U8290 ( .B1(n7380), .B2(n7383), .A(n13795), .ZN(n7379) );
  INV_X1 U8291 ( .A(n10610), .ZN(n6803) );
  AND2_X1 U8292 ( .A1(n9494), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9505) );
  NOR2_X1 U8293 ( .A1(n14095), .A2(n14089), .ZN(n14071) );
  NAND2_X1 U8294 ( .A1(n7096), .A2(n14147), .ZN(n7095) );
  NAND2_X1 U8295 ( .A1(n7097), .A2(n7099), .ZN(n7096) );
  NOR2_X1 U8296 ( .A1(n14214), .A2(n14518), .ZN(n7183) );
  NAND2_X1 U8297 ( .A1(n7122), .A2(n7120), .ZN(n7118) );
  INV_X1 U8298 ( .A(n7120), .ZN(n7119) );
  NOR2_X1 U8299 ( .A1(n11882), .A2(n7187), .ZN(n7186) );
  INV_X1 U8300 ( .A(n7188), .ZN(n7187) );
  NAND2_X1 U8301 ( .A1(n7108), .A2(n7110), .ZN(n7107) );
  NAND2_X1 U8302 ( .A1(n7113), .A2(n6438), .ZN(n7108) );
  NAND2_X1 U8303 ( .A1(n7112), .A2(n6438), .ZN(n7110) );
  AND2_X1 U8304 ( .A1(n7064), .A2(n12011), .ZN(n7063) );
  NOR2_X1 U8305 ( .A1(n7506), .A2(n7510), .ZN(n7505) );
  INV_X1 U8306 ( .A(n9034), .ZN(n7506) );
  INV_X1 U8307 ( .A(n8417), .ZN(n7491) );
  INV_X1 U8308 ( .A(n8411), .ZN(n8412) );
  NAND2_X1 U8309 ( .A1(n6894), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7365) );
  INV_X1 U8310 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9183) );
  INV_X1 U8311 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U8312 ( .A1(n7024), .A2(n7073), .ZN(n8780) );
  AOI21_X1 U8313 ( .B1(n7076), .B2(n7079), .A(n7074), .ZN(n7073) );
  NAND2_X1 U8314 ( .A1(n7475), .A2(n7076), .ZN(n7024) );
  INV_X1 U8315 ( .A(n8394), .ZN(n7074) );
  NAND2_X1 U8316 ( .A1(n6448), .A2(n9181), .ZN(n9387) );
  INV_X1 U8317 ( .A(n8388), .ZN(n8820) );
  INV_X1 U8318 ( .A(n6612), .ZN(n6611) );
  NAND2_X1 U8319 ( .A1(n7498), .A2(n7091), .ZN(n7090) );
  OAI21_X1 U8320 ( .B1(n7499), .B2(n7501), .A(n6526), .ZN(n6612) );
  NAND2_X1 U8321 ( .A1(n7689), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6716) );
  AOI21_X1 U8322 ( .B1(n8246), .B2(n7225), .A(n7224), .ZN(n8248) );
  AND2_X1 U8323 ( .A1(n13883), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7224) );
  INV_X1 U8324 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n8247) );
  NOR2_X1 U8325 ( .A1(n8260), .A2(n8259), .ZN(n8313) );
  NOR2_X1 U8326 ( .A1(n8311), .A2(n13962), .ZN(n8259) );
  OAI21_X1 U8327 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n8264), .A(n8263), .ZN(
        n8283) );
  OAI21_X1 U8328 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n12396), .A(n8273), .ZN(
        n8275) );
  AOI21_X1 U8329 ( .B1(n7204), .B2(n7207), .A(n6528), .ZN(n7203) );
  AND2_X1 U8330 ( .A1(n12127), .A2(n12190), .ZN(n7215) );
  AOI21_X1 U8331 ( .B1(n7203), .B2(n7201), .A(n6484), .ZN(n7200) );
  INV_X1 U8332 ( .A(n7204), .ZN(n7201) );
  OR2_X1 U8333 ( .A1(n12780), .A2(n10597), .ZN(n10541) );
  NAND2_X1 U8334 ( .A1(n6753), .A2(n6755), .ZN(n12128) );
  INV_X1 U8335 ( .A(n11535), .ZN(n6753) );
  NAND2_X1 U8336 ( .A1(n12216), .A2(n12158), .ZN(n12162) );
  NAND2_X1 U8337 ( .A1(n12189), .A2(n12132), .ZN(n12227) );
  AND2_X1 U8338 ( .A1(n11611), .A2(n11610), .ZN(n11624) );
  OR2_X1 U8339 ( .A1(n10189), .A2(n7702), .ZN(n10259) );
  AND2_X1 U8340 ( .A1(n6685), .A2(n6684), .ZN(n10256) );
  NAND2_X1 U8341 ( .A1(n11248), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n6684) );
  OR2_X1 U8342 ( .A1(n11248), .A2(n7702), .ZN(n6685) );
  XNOR2_X1 U8343 ( .A(n10278), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10261) );
  NAND2_X1 U8344 ( .A1(n10259), .A2(n7645), .ZN(n10260) );
  XNOR2_X1 U8345 ( .A(n10323), .B(n10317), .ZN(n10325) );
  OR2_X1 U8346 ( .A1(n10327), .A2(n10326), .ZN(n10378) );
  AND2_X1 U8347 ( .A1(n10320), .A2(n10319), .ZN(n10322) );
  NOR2_X1 U8348 ( .A1(n10322), .A2(n10321), .ZN(n10376) );
  NOR2_X1 U8349 ( .A1(n10476), .A2(n10477), .ZN(n10570) );
  NAND2_X1 U8350 ( .A1(n10373), .A2(n6473), .ZN(n6664) );
  AOI21_X1 U8351 ( .B1(n10372), .B2(n6473), .A(n6663), .ZN(n6662) );
  INV_X1 U8352 ( .A(n10472), .ZN(n6663) );
  XNOR2_X1 U8353 ( .A(n11068), .B(n11078), .ZN(n14997) );
  NOR2_X1 U8354 ( .A1(n11075), .A2(n7154), .ZN(n11077) );
  NOR2_X1 U8355 ( .A1(n11067), .A2(n11099), .ZN(n7154) );
  OAI21_X1 U8356 ( .B1(n11067), .B2(n7796), .A(n11066), .ZN(n11068) );
  NAND2_X1 U8357 ( .A1(n14997), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n14996) );
  XNOR2_X1 U8358 ( .A(n11254), .B(n11241), .ZN(n11071) );
  NAND2_X1 U8359 ( .A1(n11071), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n11255) );
  OR2_X1 U8360 ( .A1(n11242), .A2(n11243), .ZN(n7160) );
  XNOR2_X1 U8361 ( .A(n12375), .B(n12365), .ZN(n11481) );
  NAND2_X1 U8362 ( .A1(n11481), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12376) );
  OR2_X1 U8363 ( .A1(n12361), .A2(n12362), .ZN(n6858) );
  AND2_X1 U8364 ( .A1(n6677), .A2(n6676), .ZN(n12441) );
  NAND2_X1 U8365 ( .A1(n6483), .A2(n12414), .ZN(n6676) );
  NOR2_X1 U8366 ( .A1(n7163), .A2(n6470), .ZN(n7162) );
  INV_X1 U8367 ( .A(n7165), .ZN(n7163) );
  NOR2_X1 U8368 ( .A1(n15001), .A2(n7166), .ZN(n7165) );
  INV_X1 U8369 ( .A(n7167), .ZN(n7166) );
  AOI22_X1 U8370 ( .A1(n6470), .A2(n14447), .B1(n12444), .B2(n7170), .ZN(n7167) );
  NAND2_X1 U8371 ( .A1(n6931), .A2(n12444), .ZN(n7169) );
  NOR2_X1 U8372 ( .A1(n12206), .A2(n7300), .ZN(n7299) );
  INV_X1 U8373 ( .A(n8190), .ZN(n7300) );
  INV_X1 U8374 ( .A(n7299), .ZN(n7298) );
  AND2_X1 U8375 ( .A1(n11781), .A2(n11620), .ZN(n9672) );
  NAND2_X1 U8376 ( .A1(n12475), .A2(n11747), .ZN(n9671) );
  NAND2_X1 U8377 ( .A1(n7301), .A2(n7299), .ZN(n9652) );
  OAI21_X1 U8378 ( .B1(n12504), .B2(n6601), .A(n6598), .ZN(n12477) );
  INV_X1 U8379 ( .A(n11740), .ZN(n6601) );
  AOI21_X1 U8380 ( .B1(n11740), .B2(n6600), .A(n6599), .ZN(n6598) );
  INV_X1 U8381 ( .A(n8092), .ZN(n6600) );
  XNOR2_X1 U8382 ( .A(n12511), .B(n12519), .ZN(n12503) );
  OAI21_X1 U8383 ( .B1(n12560), .B2(n7305), .A(n7302), .ZN(n8183) );
  AOI21_X1 U8384 ( .B1(n7304), .B2(n7306), .A(n7303), .ZN(n7302) );
  OAI21_X1 U8385 ( .B1(n7308), .B2(n7306), .A(n7304), .ZN(n12531) );
  NAND2_X1 U8386 ( .A1(n7999), .A2(n7998), .ZN(n8012) );
  INV_X1 U8387 ( .A(n8000), .ZN(n7999) );
  AOI21_X1 U8388 ( .B1(n7294), .B2(n12610), .A(n6513), .ZN(n7293) );
  AOI21_X1 U8389 ( .B1(n7282), .B2(n7285), .A(n6512), .ZN(n7280) );
  NAND2_X1 U8390 ( .A1(n12658), .A2(n7282), .ZN(n7281) );
  NAND2_X1 U8391 ( .A1(n7922), .A2(n7921), .ZN(n7941) );
  INV_X1 U8392 ( .A(n7923), .ZN(n7922) );
  OAI21_X1 U8393 ( .B1(n12682), .B2(n6605), .A(n6603), .ZN(n6606) );
  INV_X1 U8394 ( .A(n6604), .ZN(n6603) );
  OAI21_X1 U8395 ( .B1(n6998), .B2(n6605), .A(n12641), .ZN(n6604) );
  NAND2_X1 U8396 ( .A1(n7275), .A2(n7274), .ZN(n12684) );
  OR2_X1 U8397 ( .A1(n7827), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7846) );
  OR2_X1 U8398 ( .A1(n7846), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7866) );
  AOI21_X1 U8399 ( .B1(n7288), .B2(n7290), .A(n6491), .ZN(n7286) );
  NAND2_X1 U8400 ( .A1(n11223), .A2(n8170), .ZN(n11367) );
  NAND2_X1 U8401 ( .A1(n8169), .A2(n8168), .ZN(n11223) );
  NOR2_X1 U8402 ( .A1(n7780), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7798) );
  AND2_X1 U8403 ( .A1(n7798), .A2(n7797), .ZN(n7814) );
  NAND2_X1 U8404 ( .A1(n7291), .A2(n7292), .ZN(n11090) );
  INV_X1 U8405 ( .A(n11332), .ZN(n11767) );
  OR2_X1 U8406 ( .A1(n7763), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U8407 ( .A1(n15025), .A2(n11653), .ZN(n11333) );
  NAND2_X1 U8408 ( .A1(n7744), .A2(n11650), .ZN(n15026) );
  NAND2_X1 U8409 ( .A1(n15026), .A2(n15028), .ZN(n15025) );
  INV_X1 U8410 ( .A(n8160), .ZN(n15028) );
  NAND2_X1 U8411 ( .A1(n11642), .A2(n7572), .ZN(n7571) );
  AND2_X1 U8412 ( .A1(n15084), .A2(n8151), .ZN(n15132) );
  AND2_X1 U8413 ( .A1(n10177), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9692) );
  INV_X1 U8414 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7672) );
  INV_X1 U8415 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7580) );
  INV_X1 U8416 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7684) );
  INV_X1 U8417 ( .A(n8192), .ZN(n11058) );
  NAND2_X1 U8418 ( .A1(n8068), .A2(n8080), .ZN(n8079) );
  NOR2_X1 U8419 ( .A1(n6909), .A2(n7667), .ZN(n7668) );
  AND2_X1 U8420 ( .A1(n7969), .A2(n7951), .ZN(n7952) );
  INV_X1 U8421 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7933) );
  INV_X1 U8422 ( .A(n7902), .ZN(n6930) );
  AOI21_X1 U8423 ( .B1(n7404), .B2(n7406), .A(n6564), .ZN(n7402) );
  NAND2_X1 U8424 ( .A1(n7806), .A2(n7404), .ZN(n7401) );
  INV_X1 U8425 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7787) );
  XNOR2_X1 U8426 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7773) );
  XNOR2_X1 U8427 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7754) );
  NAND2_X1 U8428 ( .A1(n8453), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8684) );
  INV_X1 U8429 ( .A(n12968), .ZN(n7340) );
  XNOR2_X1 U8430 ( .A(n12966), .B(n10297), .ZN(n9701) );
  OR2_X1 U8431 ( .A1(n9003), .A2(n9002), .ZN(n9005) );
  INV_X1 U8432 ( .A(n8960), .ZN(n8457) );
  OR2_X1 U8433 ( .A1(n8984), .A2(n13019), .ZN(n9003) );
  INV_X1 U8434 ( .A(n9710), .ZN(n6651) );
  OR2_X1 U8435 ( .A1(n8751), .A2(n8750), .ZN(n8769) );
  NAND2_X1 U8436 ( .A1(n8788), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8862) );
  OR2_X1 U8437 ( .A1(n8862), .A2(n13170), .ZN(n8883) );
  NAND2_X1 U8438 ( .A1(n10507), .A2(n10508), .ZN(n10506) );
  AND2_X1 U8439 ( .A1(n8474), .A2(n9693), .ZN(n9694) );
  AOI222_X1 U8440 ( .A1(n8767), .A2(P2_REG2_REG_31__SCAN_IN), .B1(n9073), .B2(
        P2_REG1_REG_31__SCAN_IN), .C1(n9074), .C2(P2_REG0_REG_31__SCAN_IN), 
        .ZN(n9108) );
  NAND2_X1 U8441 ( .A1(n9074), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8481) );
  AOI21_X1 U8442 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n10134), .A(n10133), .ZN(
        n10136) );
  AOI21_X1 U8443 ( .B1(n10631), .B2(P2_REG1_REG_13__SCAN_IN), .A(n10630), .ZN(
        n10632) );
  NOR2_X1 U8444 ( .A1(n11207), .A2(n13147), .ZN(n11209) );
  AOI21_X1 U8445 ( .B1(n13166), .B2(P2_REG1_REG_17__SCAN_IN), .A(n13165), .ZN(
        n13167) );
  NAND2_X1 U8446 ( .A1(n7151), .A2(n9125), .ZN(n7150) );
  INV_X1 U8447 ( .A(n7152), .ZN(n7151) );
  INV_X1 U8448 ( .A(n13498), .ZN(n7146) );
  NAND2_X1 U8449 ( .A1(n7149), .A2(n7148), .ZN(n13338) );
  OAI21_X1 U8450 ( .B1(n13362), .B2(n6472), .A(n6711), .ZN(n13330) );
  INV_X1 U8451 ( .A(n7144), .ZN(n13429) );
  NOR2_X1 U8452 ( .A1(n12092), .A2(n13445), .ZN(n6730) );
  NOR2_X1 U8453 ( .A1(n12094), .A2(n12093), .ZN(n6731) );
  NAND2_X1 U8454 ( .A1(n11465), .A2(n14500), .ZN(n13447) );
  OR2_X1 U8455 ( .A1(n8730), .A2(n8729), .ZN(n8751) );
  OR2_X1 U8456 ( .A1(n8684), .A2(n8683), .ZN(n8704) );
  NAND2_X1 U8457 ( .A1(n8454), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8730) );
  INV_X1 U8458 ( .A(n8704), .ZN(n8454) );
  AOI21_X1 U8459 ( .B1(n7264), .B2(n7262), .A(n6493), .ZN(n6707) );
  INV_X1 U8460 ( .A(n11110), .ZN(n7262) );
  INV_X1 U8461 ( .A(n7142), .ZN(n11163) );
  OR2_X1 U8462 ( .A1(n8641), .A2(n8640), .ZN(n8665) );
  OAI211_X1 U8463 ( .C1(n7443), .C2(n10863), .A(n10941), .B(n7441), .ZN(n10945) );
  NAND2_X1 U8464 ( .A1(n7448), .A2(n7446), .ZN(n10970) );
  NAND2_X1 U8465 ( .A1(n7448), .A2(n10861), .ZN(n10968) );
  NAND2_X1 U8466 ( .A1(n6593), .A2(n6592), .ZN(n10960) );
  NAND2_X1 U8467 ( .A1(n10660), .A2(n10659), .ZN(n10811) );
  OAI22_X1 U8468 ( .A1(n10296), .A2(n14869), .B1(n13116), .B2(n10297), .ZN(
        n10657) );
  NAND2_X1 U8469 ( .A1(n7021), .A2(n7250), .ZN(n7019) );
  OAI21_X1 U8470 ( .B1(n9694), .B2(n7350), .A(n13188), .ZN(n14922) );
  NOR2_X1 U8471 ( .A1(n8474), .A2(n9693), .ZN(n7350) );
  INV_X1 U8472 ( .A(n8936), .ZN(n7497) );
  NAND2_X1 U8473 ( .A1(n8433), .A2(n8432), .ZN(n8443) );
  OR2_X1 U8474 ( .A1(n8799), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8801) );
  OR2_X1 U8475 ( .A1(n8746), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8825) );
  OR2_X1 U8476 ( .A1(n8633), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8635) );
  OR2_X1 U8477 ( .A1(n8635), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8676) );
  AND2_X1 U8478 ( .A1(n10452), .A2(n10453), .ZN(n7354) );
  NAND2_X1 U8479 ( .A1(n11127), .A2(n7374), .ZN(n7371) );
  INV_X1 U8480 ( .A(n7372), .ZN(n7369) );
  NAND2_X1 U8481 ( .A1(n6798), .A2(n6800), .ZN(n6795) );
  NAND2_X1 U8482 ( .A1(n7354), .A2(n10689), .ZN(n6800) );
  NOR2_X1 U8483 ( .A1(n9410), .A2(n9409), .ZN(n9424) );
  OAI21_X1 U8484 ( .B1(n7378), .B2(n13617), .A(n7376), .ZN(n13793) );
  AOI21_X1 U8485 ( .B1(n7379), .B2(n7381), .A(n7377), .ZN(n7376) );
  INV_X1 U8486 ( .A(n7379), .ZN(n7378) );
  INV_X1 U8487 ( .A(n13794), .ZN(n7377) );
  NAND2_X1 U8488 ( .A1(n7354), .A2(n6803), .ZN(n6798) );
  NAND2_X1 U8489 ( .A1(n6797), .A2(n6803), .ZN(n6796) );
  INV_X1 U8490 ( .A(n10609), .ZN(n6797) );
  NOR2_X1 U8491 ( .A1(n9461), .A2(n9460), .ZN(n9469) );
  AND2_X1 U8492 ( .A1(n9353), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U8493 ( .A1(n13655), .A2(n7362), .ZN(n13772) );
  OR2_X1 U8494 ( .A1(n9328), .A2(n9327), .ZN(n9337) );
  NOR2_X1 U8495 ( .A1(n9337), .A2(n9336), .ZN(n9353) );
  OR2_X1 U8496 ( .A1(n9393), .A2(n9392), .ZN(n9410) );
  OR2_X1 U8497 ( .A1(n9380), .A2(n9379), .ZN(n9393) );
  NAND2_X1 U8498 ( .A1(n11972), .A2(n11973), .ZN(n11976) );
  NAND2_X1 U8499 ( .A1(n9228), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n11803) );
  AND4_X1 U8500 ( .A1(n9385), .A2(n9384), .A3(n9383), .A4(n9382), .ZN(n13850)
         );
  AND4_X1 U8501 ( .A1(n9305), .A2(n9304), .A3(n9303), .A4(n9302), .ZN(n11266)
         );
  OR2_X1 U8502 ( .A1(n9254), .A2(n9928), .ZN(n6892) );
  NAND2_X1 U8503 ( .A1(n9228), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9199) );
  OR2_X1 U8504 ( .A1(n9254), .A2(n9929), .ZN(n9201) );
  OR2_X1 U8505 ( .A1(n11802), .A2(n9955), .ZN(n9198) );
  NAND2_X1 U8506 ( .A1(n7137), .A2(n7136), .ZN(n14009) );
  NAND2_X1 U8507 ( .A1(n7140), .A2(n9549), .ZN(n7136) );
  AND2_X1 U8508 ( .A1(n14032), .A2(n9549), .ZN(n7138) );
  OR2_X1 U8509 ( .A1(n14252), .A2(n7182), .ZN(n14001) );
  NAND2_X1 U8510 ( .A1(n14055), .A2(n13847), .ZN(n14038) );
  NAND2_X1 U8511 ( .A1(n14032), .A2(n7069), .ZN(n7064) );
  NAND2_X1 U8512 ( .A1(n14051), .A2(n7070), .ZN(n7068) );
  NAND2_X1 U8513 ( .A1(n14044), .A2(n7070), .ZN(n14028) );
  NAND2_X1 U8514 ( .A1(n14030), .A2(n14404), .ZN(n6953) );
  NAND2_X1 U8515 ( .A1(n6769), .A2(n6770), .ZN(n14046) );
  OR2_X1 U8516 ( .A1(n6958), .A2(n6772), .ZN(n6770) );
  AND2_X1 U8517 ( .A1(n9505), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9519) );
  OAI21_X1 U8518 ( .B1(n14159), .B2(n6776), .A(n6775), .ZN(n6780) );
  INV_X1 U8519 ( .A(n6777), .ZN(n6776) );
  AOI21_X1 U8520 ( .B1(n6777), .B2(n7599), .A(n7596), .ZN(n6775) );
  NAND2_X1 U8521 ( .A1(n7177), .A2(n14100), .ZN(n14095) );
  NAND2_X1 U8522 ( .A1(n9424), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9452) );
  NAND2_X1 U8523 ( .A1(n14209), .A2(n6455), .ZN(n14174) );
  NAND2_X1 U8524 ( .A1(n14209), .A2(n9633), .ZN(n14210) );
  INV_X1 U8525 ( .A(n9386), .ZN(n7132) );
  NAND2_X1 U8526 ( .A1(n7625), .A2(n9625), .ZN(n14220) );
  NAND2_X1 U8527 ( .A1(n6762), .A2(n9623), .ZN(n11495) );
  NAND3_X1 U8528 ( .A1(n14629), .A2(n7186), .A3(n7185), .ZN(n14413) );
  NAND2_X1 U8529 ( .A1(n14629), .A2(n7186), .ZN(n14412) );
  NAND2_X1 U8530 ( .A1(n14629), .A2(n11873), .ZN(n11177) );
  NAND2_X1 U8531 ( .A1(n14624), .A2(n11868), .ZN(n11027) );
  AND2_X1 U8532 ( .A1(n14631), .A2(n14737), .ZN(n14629) );
  NOR2_X1 U8533 ( .A1(n14648), .A2(n14724), .ZN(n14631) );
  NAND2_X1 U8534 ( .A1(n10736), .A2(n9611), .ZN(n10556) );
  NAND2_X1 U8535 ( .A1(n10736), .A2(n6893), .ZN(n10558) );
  AND2_X1 U8536 ( .A1(n9612), .A2(n9611), .ZN(n6893) );
  XNOR2_X1 U8537 ( .A(n13870), .B(n10616), .ZN(n11990) );
  INV_X1 U8538 ( .A(n14700), .ZN(n10616) );
  NOR2_X1 U8539 ( .A1(n10744), .A2(n14700), .ZN(n10645) );
  OR2_X1 U8540 ( .A1(n10885), .A2(n11839), .ZN(n10744) );
  NAND2_X1 U8541 ( .A1(n10737), .A2(n11987), .ZN(n10736) );
  NAND2_X1 U8542 ( .A1(n10878), .A2(n9610), .ZN(n10737) );
  XNOR2_X1 U8543 ( .A(n13871), .B(n11839), .ZN(n11987) );
  NAND2_X1 U8544 ( .A1(n7179), .A2(n14692), .ZN(n10885) );
  INV_X1 U8545 ( .A(n10883), .ZN(n7179) );
  AND2_X1 U8546 ( .A1(n11822), .A2(n11824), .ZN(n10879) );
  NAND2_X1 U8547 ( .A1(n11989), .A2(n10879), .ZN(n10878) );
  NOR2_X1 U8548 ( .A1(n12015), .A2(n7127), .ZN(n7125) );
  INV_X1 U8549 ( .A(n9562), .ZN(n7127) );
  NAND2_X1 U8550 ( .A1(n7602), .A2(n11926), .ZN(n14125) );
  NAND2_X1 U8551 ( .A1(n9448), .A2(n9447), .ZN(n14299) );
  INV_X1 U8553 ( .A(n14723), .ZN(n14743) );
  INV_X1 U8554 ( .A(n9636), .ZN(n10167) );
  AND2_X1 U8555 ( .A1(n7622), .A2(n9190), .ZN(n7619) );
  INV_X1 U8556 ( .A(n9052), .ZN(n6628) );
  AND2_X1 U8557 ( .A1(n9186), .A2(n7435), .ZN(n7434) );
  XNOR2_X1 U8558 ( .A(n9580), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9593) );
  XNOR2_X1 U8559 ( .A(n9581), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9594) );
  XNOR2_X1 U8560 ( .A(n9574), .B(n9573), .ZN(n9865) );
  INV_X1 U8561 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9573) );
  NOR2_X1 U8562 ( .A1(n9571), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n6788) );
  OR2_X1 U8563 ( .A1(n9405), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U8564 ( .A1(n7075), .A2(n7080), .ZN(n8798) );
  NAND2_X1 U8565 ( .A1(n7475), .A2(n7476), .ZN(n7075) );
  XNOR2_X1 U8566 ( .A(n9376), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10716) );
  NAND2_X1 U8567 ( .A1(n8742), .A2(n8741), .ZN(n8744) );
  NAND2_X1 U8568 ( .A1(n8717), .A2(n8379), .ZN(n8742) );
  OR2_X1 U8569 ( .A1(n9346), .A2(n9345), .ZN(n9350) );
  NAND2_X1 U8570 ( .A1(n8370), .A2(n8369), .ZN(n8697) );
  OAI21_X1 U8571 ( .B1(n8613), .B2(n7091), .A(n6727), .ZN(n6729) );
  INV_X1 U8572 ( .A(n6728), .ZN(n6727) );
  NAND2_X1 U8573 ( .A1(n8366), .A2(n8365), .ZN(n8632) );
  XNOR2_X1 U8574 ( .A(n8613), .B(n8612), .ZN(n9868) );
  OR2_X1 U8575 ( .A1(n9388), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U8576 ( .A1(n7689), .A2(n8344), .ZN(n6715) );
  INV_X1 U8577 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n15209) );
  NOR2_X1 U8578 ( .A1(n8295), .A2(n15329), .ZN(n8296) );
  INV_X1 U8579 ( .A(n8246), .ZN(n8291) );
  INV_X1 U8580 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U8581 ( .A1(n15317), .A2(n8303), .ZN(n8305) );
  NOR2_X1 U8582 ( .A1(n8255), .A2(n8254), .ZN(n8306) );
  INV_X1 U8583 ( .A(n6859), .ZN(n8253) );
  NOR2_X1 U8584 ( .A1(n14394), .A2(n8319), .ZN(n8320) );
  INV_X1 U8585 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6884) );
  OAI21_X1 U8586 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n8271), .A(n8270), .ZN(
        n8280) );
  NAND2_X1 U8587 ( .A1(n14588), .A2(n6461), .ZN(n6874) );
  AND2_X1 U8588 ( .A1(n14586), .A2(n6877), .ZN(n6871) );
  AND2_X1 U8589 ( .A1(n14588), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6876) );
  NOR2_X1 U8590 ( .A1(n14428), .A2(n11444), .ZN(n6878) );
  XNOR2_X1 U8591 ( .A(n12264), .B(n12263), .ZN(n6761) );
  NAND2_X1 U8592 ( .A1(n12128), .A2(n7215), .ZN(n12189) );
  NAND2_X1 U8593 ( .A1(n7211), .A2(n10596), .ZN(n10599) );
  OAI21_X1 U8594 ( .B1(n7198), .B2(n7206), .A(n7194), .ZN(n7193) );
  NAND2_X1 U8595 ( .A1(n7198), .A2(n7195), .ZN(n7194) );
  NAND2_X1 U8596 ( .A1(n7196), .A2(n12207), .ZN(n7195) );
  INV_X1 U8597 ( .A(n7200), .ZN(n7196) );
  NAND2_X1 U8598 ( .A1(n7198), .A2(n12207), .ZN(n7197) );
  OR2_X1 U8599 ( .A1(n6441), .A2(n12122), .ZN(n8127) );
  NAND2_X1 U8600 ( .A1(n12274), .A2(n12156), .ZN(n12218) );
  NAND2_X1 U8601 ( .A1(n6739), .A2(n6743), .ZN(n12248) );
  NAND2_X1 U8602 ( .A1(n12336), .A2(n6744), .ZN(n6739) );
  OAI21_X1 U8603 ( .B1(n12336), .B2(n6742), .A(n6740), .ZN(n6745) );
  INV_X1 U8604 ( .A(n6741), .ZN(n6740) );
  OAI21_X1 U8605 ( .B1(n6744), .B2(n6742), .A(n12246), .ZN(n6741) );
  AOI21_X1 U8606 ( .B1(n12264), .B2(n6760), .A(n6562), .ZN(n12268) );
  NAND2_X1 U8607 ( .A1(n12164), .A2(n12549), .ZN(n6760) );
  AND2_X1 U8608 ( .A1(n10902), .A2(n10901), .ZN(n10903) );
  NAND2_X1 U8609 ( .A1(n12276), .A2(n12275), .ZN(n12274) );
  NAND2_X1 U8610 ( .A1(n12198), .A2(n12153), .ZN(n12276) );
  AOI21_X1 U8611 ( .B1(n7212), .B2(n6754), .A(n6751), .ZN(n6750) );
  NAND2_X1 U8612 ( .A1(n11535), .A2(n7212), .ZN(n6752) );
  NAND2_X1 U8613 ( .A1(n6755), .A2(n12132), .ZN(n6754) );
  AND4_X1 U8614 ( .A1(n7852), .A2(n7851), .A3(n7850), .A4(n7849), .ZN(n12309)
         );
  NAND2_X1 U8615 ( .A1(n7209), .A2(n11042), .ZN(n11043) );
  AOI21_X1 U8616 ( .B1(n12483), .B2(n8193), .A(n8119), .ZN(n12328) );
  NAND2_X1 U8617 ( .A1(n10550), .A2(n15066), .ZN(n12327) );
  INV_X1 U8618 ( .A(n7207), .ZN(n6956) );
  NAND2_X1 U8619 ( .A1(n8098), .A2(n6580), .ZN(n12496) );
  NAND2_X1 U8620 ( .A1(n15083), .A2(n10353), .ZN(n12330) );
  INV_X1 U8621 ( .A(n12332), .ZN(n12337) );
  INV_X1 U8622 ( .A(n11624), .ZN(n12463) );
  AND2_X1 U8623 ( .A1(n11611), .A2(n8198), .ZN(n12210) );
  INV_X1 U8624 ( .A(n12328), .ZN(n12490) );
  OR2_X1 U8625 ( .A1(n10344), .A2(n12848), .ZN(n12352) );
  INV_X1 U8626 ( .A(n12563), .ZN(n12590) );
  INV_X1 U8627 ( .A(n12604), .ZN(n12355) );
  INV_X1 U8628 ( .A(n12309), .ZN(n12688) );
  OR2_X1 U8629 ( .A1(n8029), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U8630 ( .A1(n7678), .A2(n6733), .ZN(n6737) );
  NOR2_X1 U8631 ( .A1(n7677), .A2(n7703), .ZN(n6733) );
  CLKBUF_X1 U8632 ( .A(n12771), .Z(n6905) );
  INV_X1 U8633 ( .A(n7157), .ZN(n10780) );
  NAND2_X1 U8634 ( .A1(n10773), .A2(n10774), .ZN(n10775) );
  AOI21_X1 U8635 ( .B1(n10770), .B2(n10769), .A(n6665), .ZN(n11055) );
  INV_X1 U8636 ( .A(n7156), .ZN(n10782) );
  XNOR2_X1 U8637 ( .A(n11077), .B(n11078), .ZN(n14983) );
  NOR2_X1 U8638 ( .A1(n14983), .A2(n14984), .ZN(n14982) );
  INV_X1 U8639 ( .A(n6681), .ZN(n6678) );
  INV_X1 U8640 ( .A(n7160), .ZN(n11246) );
  XNOR2_X1 U8641 ( .A(n12360), .B(n12365), .ZN(n11473) );
  NOR2_X1 U8642 ( .A1(n11473), .A2(n7882), .ZN(n12361) );
  INV_X1 U8643 ( .A(n7158), .ZN(n12389) );
  INV_X1 U8644 ( .A(n6858), .ZN(n12363) );
  OAI21_X1 U8645 ( .B1(n12390), .B2(n6853), .A(n6851), .ZN(n12432) );
  OR2_X1 U8646 ( .A1(n12412), .A2(n12391), .ZN(n6853) );
  NAND2_X1 U8647 ( .A1(n12411), .A2(n6852), .ZN(n6851) );
  INV_X1 U8648 ( .A(n12412), .ZN(n6852) );
  INV_X1 U8649 ( .A(n12411), .ZN(n6854) );
  NAND2_X1 U8650 ( .A1(n11602), .A2(n11601), .ZN(n14478) );
  NAND2_X1 U8651 ( .A1(n12504), .A2(n8092), .ZN(n12492) );
  NAND2_X1 U8652 ( .A1(n12520), .A2(n11777), .ZN(n12523) );
  NAND2_X1 U8653 ( .A1(n12558), .A2(n8181), .ZN(n12547) );
  AND2_X1 U8654 ( .A1(n12577), .A2(n12576), .ZN(n12735) );
  AND2_X1 U8655 ( .A1(n7012), .A2(n11719), .ZN(n12582) );
  NAND2_X1 U8656 ( .A1(n7985), .A2(n11711), .ZN(n12586) );
  NAND2_X1 U8657 ( .A1(n7566), .A2(n11715), .ZN(n12599) );
  NAND2_X1 U8658 ( .A1(n12612), .A2(n8177), .ZN(n12600) );
  NAND2_X1 U8659 ( .A1(n6602), .A2(n7000), .ZN(n12642) );
  NAND2_X1 U8660 ( .A1(n12682), .A2(n6998), .ZN(n6602) );
  OAI21_X1 U8661 ( .B1(n12658), .B2(n7285), .A(n7282), .ZN(n12643) );
  OAI21_X1 U8662 ( .B1(n12682), .B2(n7006), .A(n7003), .ZN(n12655) );
  NAND2_X1 U8663 ( .A1(n12681), .A2(n11687), .ZN(n12669) );
  OAI21_X1 U8664 ( .B1(n11089), .B2(n7568), .A(n7009), .ZN(n11366) );
  NAND2_X1 U8665 ( .A1(n11089), .A2(n11761), .ZN(n7569) );
  AND2_X1 U8666 ( .A1(n6608), .A2(n6607), .ZN(n11304) );
  INV_X1 U8667 ( .A(n11050), .ZN(n15112) );
  AND2_X1 U8668 ( .A1(n15091), .A2(n15090), .ZN(n12544) );
  AND2_X1 U8669 ( .A1(n15084), .A2(n11639), .ZN(n15090) );
  INV_X1 U8670 ( .A(n15053), .ZN(n15083) );
  OR2_X1 U8671 ( .A1(n8027), .A2(n9832), .ZN(n7700) );
  NAND2_X1 U8672 ( .A1(n15149), .A2(n14477), .ZN(n12769) );
  NAND2_X1 U8673 ( .A1(n7960), .A2(n7959), .ZN(n12828) );
  NAND2_X1 U8674 ( .A1(n7905), .A2(n7904), .ZN(n12841) );
  OAI22_X1 U8675 ( .A1(n11613), .A2(n11612), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n11807), .ZN(n11615) );
  INV_X1 U8676 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12851) );
  NAND2_X1 U8677 ( .A1(n8040), .A2(n8039), .ZN(n8052) );
  NOR2_X1 U8678 ( .A1(n8142), .A2(n8141), .ZN(n11793) );
  NAND2_X1 U8679 ( .A1(n8137), .A2(n8138), .ZN(n10515) );
  NAND2_X1 U8680 ( .A1(n8022), .A2(n8021), .ZN(n8025) );
  INV_X1 U8681 ( .A(SI_20_), .ZN(n10424) );
  INV_X1 U8682 ( .A(n8019), .ZN(n8018) );
  OAI21_X1 U8683 ( .B1(n7973), .B2(n7414), .A(n7412), .ZN(n8009) );
  NAND2_X1 U8684 ( .A1(n7987), .A2(n7986), .ZN(n7990) );
  INV_X1 U8685 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7992) );
  INV_X1 U8686 ( .A(SI_17_), .ZN(n10078) );
  NAND2_X1 U8687 ( .A1(n7389), .A2(n7391), .ZN(n7948) );
  OR2_X1 U8688 ( .A1(n7916), .A2(n7394), .ZN(n7389) );
  NAND2_X1 U8689 ( .A1(n7916), .A2(n7915), .ZN(n7930) );
  INV_X1 U8690 ( .A(SI_14_), .ZN(n9889) );
  INV_X1 U8691 ( .A(SI_13_), .ZN(n14377) );
  NAND2_X1 U8692 ( .A1(n7900), .A2(n6698), .ZN(n7899) );
  NAND2_X1 U8693 ( .A1(n7415), .A2(n7874), .ZN(n7891) );
  INV_X1 U8694 ( .A(SI_12_), .ZN(n9862) );
  NAND2_X1 U8695 ( .A1(n7770), .A2(n7876), .ZN(n7218) );
  NAND2_X1 U8696 ( .A1(n7857), .A2(n7856), .ZN(n7873) );
  XNOR2_X1 U8697 ( .A(n7836), .B(P3_IR_REG_10__SCAN_IN), .ZN(n15018) );
  NAND2_X1 U8698 ( .A1(n7403), .A2(n7808), .ZN(n7823) );
  NAND2_X1 U8699 ( .A1(n7806), .A2(n7805), .ZN(n7403) );
  INV_X1 U8700 ( .A(n10772), .ZN(n10779) );
  AND2_X1 U8701 ( .A1(n7737), .A2(n7736), .ZN(n10379) );
  NAND2_X1 U8702 ( .A1(n7176), .A2(n7937), .ZN(n7175) );
  NAND2_X1 U8703 ( .A1(n7317), .A2(n7319), .ZN(n10680) );
  AOI21_X1 U8704 ( .B1(n7321), .B2(n7323), .A(n7320), .ZN(n7319) );
  OR2_X1 U8705 ( .A1(n10507), .A2(n7322), .ZN(n7317) );
  NAND2_X1 U8706 ( .A1(n6635), .A2(n7341), .ZN(n12930) );
  INV_X1 U8707 ( .A(n12921), .ZN(n6635) );
  NAND2_X1 U8708 ( .A1(n13472), .A2(n13093), .ZN(n12929) );
  AND2_X1 U8709 ( .A1(n12937), .A2(n12865), .ZN(n7334) );
  OR2_X1 U8710 ( .A1(n10366), .A2(n9700), .ZN(n10400) );
  NAND2_X1 U8711 ( .A1(n13028), .A2(n6639), .ZN(n6638) );
  NOR2_X1 U8712 ( .A1(n12974), .A2(n7345), .ZN(n7344) );
  NAND2_X1 U8713 ( .A1(n13034), .A2(n12894), .ZN(n12975) );
  NAND2_X1 U8714 ( .A1(n7315), .A2(n13005), .ZN(n13013) );
  NAND2_X1 U8715 ( .A1(n6647), .A2(n7314), .ZN(n13010) );
  AND2_X1 U8716 ( .A1(n12875), .A2(n7316), .ZN(n7314) );
  INV_X1 U8717 ( .A(n12995), .ZN(n7316) );
  NAND2_X1 U8718 ( .A1(n12905), .A2(n7332), .ZN(n13014) );
  OR2_X1 U8719 ( .A1(n9789), .A2(n9788), .ZN(n12996) );
  INV_X1 U8720 ( .A(n6643), .ZN(n6642) );
  NAND2_X1 U8721 ( .A1(n9738), .A2(n10927), .ZN(n11141) );
  NAND2_X1 U8722 ( .A1(n6637), .A2(n13028), .ZN(n13034) );
  NAND2_X1 U8723 ( .A1(n13031), .A2(n12890), .ZN(n6637) );
  NAND2_X1 U8724 ( .A1(n11430), .A2(n9757), .ZN(n9779) );
  XNOR2_X1 U8725 ( .A(n12904), .B(n12902), .ZN(n13035) );
  INV_X1 U8726 ( .A(n10658), .ZN(n13048) );
  NAND2_X1 U8727 ( .A1(n13013), .A2(n12881), .ZN(n13062) );
  NAND2_X1 U8728 ( .A1(n10506), .A2(n9727), .ZN(n10531) );
  OAI21_X2 U8729 ( .B1(n9859), .B2(n8518), .A(n8596), .ZN(n10965) );
  AND2_X1 U8730 ( .A1(n9145), .A2(n11137), .ZN(n9164) );
  INV_X1 U8731 ( .A(n9086), .ZN(n9143) );
  INV_X1 U8732 ( .A(n9123), .ZN(n6974) );
  OR2_X2 U8733 ( .A1(n9799), .A2(n9691), .ZN(n13117) );
  OR2_X1 U8734 ( .A1(n14830), .A2(n14829), .ZN(n14832) );
  OAI21_X1 U8735 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n14839), .A(n14832), .ZN(
        n10092) );
  INV_X1 U8736 ( .A(n7465), .ZN(n7464) );
  NAND2_X1 U8737 ( .A1(n13225), .A2(n7467), .ZN(n7466) );
  NAND2_X1 U8738 ( .A1(n7246), .A2(n7251), .ZN(n13224) );
  NAND2_X1 U8739 ( .A1(n7245), .A2(n7252), .ZN(n7246) );
  INV_X1 U8740 ( .A(n13254), .ZN(n7245) );
  NAND2_X1 U8741 ( .A1(n7035), .A2(n7036), .ZN(n13270) );
  NAND2_X1 U8742 ( .A1(n13299), .A2(n12079), .ZN(n13283) );
  NAND2_X1 U8743 ( .A1(n7256), .A2(n6501), .ZN(n13497) );
  NAND2_X1 U8744 ( .A1(n7256), .A2(n7257), .ZN(n13311) );
  AND2_X1 U8745 ( .A1(n13303), .A2(n13302), .ZN(n13503) );
  NAND2_X1 U8746 ( .A1(n13362), .A2(n12103), .ZN(n13345) );
  NAND2_X1 U8747 ( .A1(n7461), .A2(n12069), .ZN(n13359) );
  NAND2_X1 U8748 ( .A1(n6700), .A2(n6702), .ZN(n13384) );
  NAND2_X1 U8749 ( .A1(n12100), .A2(n6446), .ZN(n13391) );
  NAND2_X1 U8750 ( .A1(n12100), .A2(n12099), .ZN(n13389) );
  NAND2_X1 U8751 ( .A1(n7044), .A2(n7451), .ZN(n13407) );
  NAND2_X1 U8752 ( .A1(n12063), .A2(n7452), .ZN(n7044) );
  NAND2_X1 U8753 ( .A1(n12063), .A2(n12062), .ZN(n13420) );
  NAND2_X1 U8754 ( .A1(n11382), .A2(n11381), .ZN(n11384) );
  NAND2_X1 U8755 ( .A1(n11111), .A2(n11110), .ZN(n11154) );
  NAND2_X1 U8756 ( .A1(n7241), .A2(n10858), .ZN(n10957) );
  INV_X1 U8757 ( .A(n9124), .ZN(n14880) );
  NOR2_X1 U8758 ( .A1(n6594), .A2(n7049), .ZN(n7048) );
  INV_X1 U8759 ( .A(n13463), .ZN(n6594) );
  INV_X1 U8760 ( .A(n6947), .ZN(n6946) );
  NAND2_X1 U8761 ( .A1(n6722), .A2(n6721), .ZN(n13558) );
  OR2_X1 U8762 ( .A1(n13480), .A2(n14934), .ZN(n6722) );
  AND2_X1 U8763 ( .A1(n13478), .A2(n13479), .ZN(n6721) );
  OR2_X1 U8764 ( .A1(n13508), .A2(n13507), .ZN(n13563) );
  INV_X1 U8765 ( .A(n14892), .ZN(n14893) );
  AND2_X1 U8766 ( .A1(n9799), .A2(n9690), .ZN(n14895) );
  INV_X1 U8767 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8463) );
  AOI21_X1 U8768 ( .B1(n8425), .B2(n7269), .A(n8438), .ZN(n6652) );
  XNOR2_X1 U8769 ( .A(n9150), .B(n9149), .ZN(n13591) );
  INV_X1 U8770 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10396) );
  INV_X1 U8771 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10335) );
  INV_X1 U8772 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10405) );
  INV_X1 U8773 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10339) );
  INV_X1 U8774 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10076) );
  INV_X1 U8775 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n15222) );
  INV_X1 U8776 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9860) );
  INV_X1 U8777 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9828) );
  INV_X1 U8778 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9825) );
  XNOR2_X1 U8779 ( .A(n8489), .B(n8488), .ZN(n10079) );
  OAI21_X1 U8780 ( .B1(n11127), .B2(n11126), .A(n11125), .ZN(n11273) );
  NAND2_X1 U8781 ( .A1(n13836), .A2(n13710), .ZN(n13711) );
  NAND2_X1 U8782 ( .A1(n6817), .A2(n6443), .ZN(n13748) );
  NAND2_X1 U8783 ( .A1(n10454), .A2(n7354), .ZN(n10611) );
  NAND2_X1 U8784 ( .A1(n6816), .A2(n6815), .ZN(n13758) );
  AOI21_X1 U8785 ( .B1(n6443), .B2(n13709), .A(n13747), .ZN(n6815) );
  XNOR2_X1 U8786 ( .A(n13756), .B(n13755), .ZN(n13757) );
  NAND2_X1 U8787 ( .A1(n13655), .A2(n13654), .ZN(n13775) );
  AOI21_X1 U8788 ( .B1(n13617), .B2(n7384), .A(n7383), .ZN(n14513) );
  OAI21_X1 U8789 ( .B1(n6798), .B2(n6793), .A(n6796), .ZN(n10688) );
  INV_X1 U8790 ( .A(n10454), .ZN(n6793) );
  NOR2_X1 U8791 ( .A1(n6943), .A2(n6942), .ZN(n11279) );
  AOI21_X1 U8792 ( .B1(n7370), .B2(n7367), .A(n6523), .ZN(n7366) );
  NAND2_X1 U8793 ( .A1(n13740), .A2(n13648), .ZN(n13812) );
  NAND2_X1 U8794 ( .A1(n11573), .A2(n7358), .ZN(n7357) );
  INV_X1 U8795 ( .A(n11575), .ZN(n7358) );
  NAND2_X1 U8796 ( .A1(n6809), .A2(n6807), .ZN(n6806) );
  NAND2_X1 U8797 ( .A1(n13772), .A2(n13662), .ZN(n13819) );
  AOI21_X1 U8798 ( .B1(n11551), .B2(n11550), .A(n6921), .ZN(n14523) );
  AND2_X1 U8799 ( .A1(n11548), .A2(n11549), .ZN(n6921) );
  NAND2_X1 U8800 ( .A1(n14523), .A2(n14524), .ZN(n14522) );
  NAND2_X1 U8801 ( .A1(n10157), .A2(n10153), .ZN(n15306) );
  XNOR2_X1 U8802 ( .A(n13617), .B(n13618), .ZN(n13849) );
  AND2_X1 U8803 ( .A1(n10919), .A2(n14723), .ZN(n15311) );
  NOR2_X1 U8804 ( .A1(n10155), .A2(n10458), .ZN(n12040) );
  INV_X1 U8805 ( .A(n12043), .ZN(n6904) );
  NAND2_X1 U8806 ( .A1(n9228), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9513) );
  NAND2_X1 U8807 ( .A1(n9228), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9487) );
  INV_X1 U8808 ( .A(n11266), .ZN(n13867) );
  NAND4_X1 U8809 ( .A1(n9291), .A2(n9290), .A3(n9289), .A4(n9288), .ZN(n14620)
         );
  NAND2_X1 U8810 ( .A1(n9228), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9222) );
  OR2_X1 U8811 ( .A1(n9254), .A2(n9934), .ZN(n9220) );
  OR2_X1 U8812 ( .A1(n9882), .A2(n10146), .ZN(n13878) );
  OR2_X1 U8813 ( .A1(n11802), .A2(n10893), .ZN(n9214) );
  OR2_X1 U8814 ( .A1(n9520), .A2(n10892), .ZN(n9216) );
  AND2_X1 U8815 ( .A1(n9215), .A2(n9217), .ZN(n6906) );
  NAND2_X1 U8816 ( .A1(n11809), .A2(n11808), .ZN(n13991) );
  NAND2_X1 U8817 ( .A1(n13998), .A2(n13997), .ZN(n13999) );
  NAND2_X1 U8818 ( .A1(n14031), .A2(n7139), .ZN(n14015) );
  AND2_X1 U8819 ( .A1(n14031), .A2(n9537), .ZN(n14016) );
  AOI21_X1 U8820 ( .B1(n6954), .B2(n14403), .A(n6951), .ZN(n14266) );
  NAND2_X1 U8821 ( .A1(n6953), .A2(n6952), .ZN(n6951) );
  XNOR2_X1 U8822 ( .A(n14028), .B(n14027), .ZN(n6954) );
  NAND2_X1 U8823 ( .A1(n14029), .A2(n14619), .ZN(n6952) );
  NAND2_X1 U8824 ( .A1(n13587), .A2(n11980), .ZN(n9504) );
  NAND2_X1 U8825 ( .A1(n7429), .A2(n7428), .ZN(n14064) );
  AND2_X1 U8826 ( .A1(n6773), .A2(n6495), .ZN(n14061) );
  NAND2_X1 U8827 ( .A1(n14078), .A2(n14084), .ZN(n6773) );
  NAND2_X1 U8828 ( .A1(n14133), .A2(n9466), .ZN(n14120) );
  NAND2_X1 U8829 ( .A1(n6779), .A2(n7061), .ZN(n14110) );
  AND2_X1 U8830 ( .A1(n6779), .A2(n6777), .ZN(n14109) );
  OAI21_X1 U8831 ( .B1(n9417), .B2(n7099), .A(n7097), .ZN(n14146) );
  NAND2_X1 U8832 ( .A1(n14159), .A2(n11817), .ZN(n14143) );
  NAND2_X1 U8833 ( .A1(n7104), .A2(n9431), .ZN(n14158) );
  NAND2_X1 U8834 ( .A1(n9417), .A2(n7105), .ZN(n7104) );
  AND2_X1 U8835 ( .A1(n14192), .A2(n9626), .ZN(n14181) );
  NAND2_X1 U8836 ( .A1(n9417), .A2(n9416), .ZN(n14173) );
  AND2_X1 U8837 ( .A1(n14205), .A2(n11901), .ZN(n14194) );
  NAND2_X1 U8838 ( .A1(n9372), .A2(n7420), .ZN(n14542) );
  NAND2_X1 U8839 ( .A1(n7117), .A2(n7120), .ZN(n14399) );
  NAND2_X1 U8840 ( .A1(n11347), .A2(n7121), .ZN(n7117) );
  AND2_X1 U8841 ( .A1(n11025), .A2(n9619), .ZN(n11171) );
  NAND2_X1 U8842 ( .A1(n9617), .A2(n9616), .ZN(n10800) );
  NAND2_X1 U8843 ( .A1(n7111), .A2(n9264), .ZN(n14637) );
  NAND2_X1 U8844 ( .A1(n10555), .A2(n7113), .ZN(n7111) );
  NAND2_X1 U8845 ( .A1(n10555), .A2(n9249), .ZN(n10638) );
  INV_X1 U8846 ( .A(n14216), .ZN(n14633) );
  NAND2_X1 U8847 ( .A1(n9863), .A2(n7426), .ZN(n7425) );
  INV_X1 U8848 ( .A(n10750), .ZN(n10896) );
  INV_X1 U8849 ( .A(n14190), .ZN(n14646) );
  NAND2_X1 U8850 ( .A1(n7085), .A2(n14748), .ZN(n7084) );
  INV_X1 U8851 ( .A(n14244), .ZN(n7085) );
  INV_X2 U8852 ( .A(n14749), .ZN(n14751) );
  NAND2_X1 U8853 ( .A1(n9865), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9882) );
  NAND2_X1 U8854 ( .A1(n9058), .A2(n7657), .ZN(n9064) );
  AND2_X1 U8855 ( .A1(n7622), .A2(n7621), .ZN(n7620) );
  NOR2_X1 U8856 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n7621) );
  XNOR2_X1 U8857 ( .A(n9204), .B(n9203), .ZN(n14344) );
  NAND2_X1 U8858 ( .A1(n8980), .A2(n7487), .ZN(n7489) );
  NAND2_X1 U8859 ( .A1(n8937), .A2(n8410), .ZN(n8955) );
  NAND2_X1 U8860 ( .A1(n9582), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U8861 ( .A1(n8913), .A2(n8912), .ZN(n8915) );
  XNOR2_X1 U8862 ( .A(n9444), .B(n9443), .ZN(n11525) );
  NAND2_X1 U8863 ( .A1(n7482), .A2(n7484), .ZN(n8856) );
  INV_X1 U8864 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10388) );
  INV_X1 U8865 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10312) );
  INV_X1 U8866 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10390) );
  INV_X1 U8867 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10338) );
  INV_X1 U8868 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10074) );
  INV_X1 U8869 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10004) );
  INV_X1 U8870 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9926) );
  INV_X1 U8871 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9857) );
  NAND2_X1 U8872 ( .A1(n7355), .A2(n9209), .ZN(n9244) );
  INV_X1 U8873 ( .A(n8513), .ZN(n8515) );
  XNOR2_X1 U8874 ( .A(n8294), .B(n9802), .ZN(n15330) );
  OAI21_X1 U8875 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14366), .A(n14367), .ZN(
        n15325) );
  XNOR2_X1 U8876 ( .A(n7221), .B(n8302), .ZN(n15319) );
  XNOR2_X1 U8877 ( .A(n8305), .B(n8304), .ZN(n14385) );
  NOR2_X1 U8878 ( .A1(n15322), .A2(n6862), .ZN(n6861) );
  INV_X1 U8879 ( .A(n6866), .ZN(n6862) );
  XNOR2_X1 U8880 ( .A(n8314), .B(n7226), .ZN(n14393) );
  INV_X1 U8881 ( .A(n8315), .ZN(n7226) );
  NAND2_X1 U8882 ( .A1(n14393), .A2(n14828), .ZN(n14392) );
  XNOR2_X1 U8883 ( .A(n8318), .B(n8317), .ZN(n14395) );
  NOR2_X1 U8884 ( .A1(n14395), .A2(n14849), .ZN(n14394) );
  OR2_X1 U8885 ( .A1(n14571), .A2(n6884), .ZN(n6883) );
  NAND2_X1 U8886 ( .A1(n14575), .A2(n14574), .ZN(n14573) );
  NAND2_X1 U8887 ( .A1(n14578), .A2(n14579), .ZN(n14577) );
  NAND2_X1 U8888 ( .A1(n11006), .A2(n11005), .ZN(n11039) );
  NAND2_X1 U8889 ( .A1(n6661), .A2(n6473), .ZN(n10473) );
  AND2_X1 U8890 ( .A1(n14460), .A2(n14461), .ZN(n6848) );
  OR2_X1 U8891 ( .A1(n14431), .A2(n6589), .ZN(n6844) );
  INV_X1 U8892 ( .A(n6659), .ZN(n6658) );
  NAND2_X1 U8893 ( .A1(n6460), .A2(n15007), .ZN(n6918) );
  NAND2_X1 U8894 ( .A1(n6657), .A2(n15015), .ZN(n6656) );
  AND2_X1 U8895 ( .A1(n7277), .A2(n9667), .ZN(n12044) );
  NAND2_X1 U8896 ( .A1(n7279), .A2(n7278), .ZN(n9689) );
  NAND2_X1 U8897 ( .A1(n15137), .A2(n9688), .ZN(n7278) );
  OAI222_X1 U8898 ( .A1(P3_U3151), .A2(n10577), .B1(n14378), .B2(n9830), .C1(
        n9829), .C2(n14376), .ZN(P3_U3289) );
  NAND2_X1 U8899 ( .A1(n13049), .A2(n9710), .ZN(n10519) );
  NAND2_X1 U8900 ( .A1(n7337), .A2(n7343), .ZN(n7336) );
  INV_X1 U8901 ( .A(n6647), .ZN(n13095) );
  MUX2_X1 U8902 ( .A(n13190), .B(n13189), .S(n13188), .Z(n13192) );
  OAI21_X1 U8903 ( .B1(n7656), .B2(n14871), .A(n7270), .ZN(P2_U3236) );
  AND2_X1 U8904 ( .A1(n13461), .A2(n14850), .ZN(n7271) );
  OAI21_X1 U8905 ( .B1(n13464), .B2(n13456), .A(n7273), .ZN(n7272) );
  NAND2_X1 U8906 ( .A1(n6898), .A2(n6897), .ZN(P2_U3528) );
  NAND2_X1 U8907 ( .A1(n14971), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U8908 ( .A1(n6899), .A2(n14974), .ZN(n6898) );
  NAND2_X1 U8909 ( .A1(n7048), .A2(n13464), .ZN(n6899) );
  AOI21_X1 U8910 ( .B1(n7049), .B2(n14959), .A(n6469), .ZN(n6595) );
  NAND2_X1 U8911 ( .A1(n6720), .A2(n6719), .ZN(P2_U3493) );
  NAND2_X1 U8912 ( .A1(n14958), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U8913 ( .A1(n13558), .A2(n14959), .ZN(n6720) );
  NAND2_X1 U8914 ( .A1(n8937), .A2(n7027), .ZN(n11493) );
  OAI21_X1 U8915 ( .B1(n14249), .B2(n14656), .A(n6960), .ZN(P1_U3356) );
  AND2_X1 U8916 ( .A1(n7083), .A2(n6556), .ZN(n14249) );
  INV_X1 U8917 ( .A(n9651), .ZN(n6961) );
  OAI21_X1 U8918 ( .B1(n7422), .B2(n14749), .A(n6923), .ZN(P1_U3525) );
  INV_X1 U8919 ( .A(n6924), .ZN(n6923) );
  OAI21_X1 U8920 ( .B1(n14244), .B2(n7124), .A(n6577), .ZN(n6924) );
  OAI21_X1 U8921 ( .B1(n12125), .B2(n11585), .A(n7630), .ZN(P1_U3325) );
  INV_X1 U8922 ( .A(n7631), .ZN(n7630) );
  INV_X1 U8923 ( .A(n7220), .ZN(n14566) );
  INV_X1 U8924 ( .A(n14570), .ZN(n6882) );
  INV_X1 U8925 ( .A(n14583), .ZN(n14582) );
  AND2_X1 U8926 ( .A1(n6879), .A2(n14586), .ZN(n14426) );
  XNOR2_X1 U8927 ( .A(n8343), .B(n8337), .ZN(n7222) );
  AND2_X1 U8928 ( .A1(n13492), .A2(n13040), .ZN(n6444) );
  AND2_X1 U8929 ( .A1(n7101), .A2(n7100), .ZN(n6445) );
  INV_X1 U8930 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8438) );
  AND2_X1 U8931 ( .A1(n12099), .A2(n13395), .ZN(n6446) );
  INV_X1 U8932 ( .A(n14214), .ZN(n9633) );
  OR2_X1 U8933 ( .A1(n7473), .A2(n9119), .ZN(n6447) );
  AOI21_X1 U8934 ( .B1(n11806), .B2(n9100), .A(n6583), .ZN(n9125) );
  INV_X1 U8935 ( .A(n14362), .ZN(n6877) );
  INV_X1 U8936 ( .A(n7568), .ZN(n7567) );
  NAND2_X1 U8937 ( .A1(n11668), .A2(n11672), .ZN(n7568) );
  AND3_X1 U8938 ( .A1(n9180), .A2(n9344), .A3(n9179), .ZN(n6448) );
  AND2_X1 U8939 ( .A1(n11966), .A2(n7640), .ZN(n6449) );
  AND2_X1 U8940 ( .A1(n8891), .A2(n8890), .ZN(n6450) );
  AND2_X1 U8941 ( .A1(n6794), .A2(n6506), .ZN(n6451) );
  AND2_X1 U8942 ( .A1(n8424), .A2(n7556), .ZN(n6452) );
  AND2_X1 U8943 ( .A1(n14400), .A2(n7118), .ZN(n6453) );
  AND2_X1 U8944 ( .A1(n13847), .A2(n7181), .ZN(n6454) );
  INV_X1 U8945 ( .A(n12534), .ZN(n7303) );
  AND2_X1 U8946 ( .A1(n7183), .A2(n14311), .ZN(n6455) );
  NOR2_X1 U8947 ( .A1(n13015), .A2(n7333), .ZN(n6456) );
  INV_X1 U8948 ( .A(n11745), .ZN(n12476) );
  NAND2_X1 U8949 ( .A1(n9010), .A2(n9009), .ZN(n13240) );
  AND2_X1 U8950 ( .A1(n10965), .A2(n10864), .ZN(n6457) );
  NAND4_X1 U8951 ( .A1(n9201), .A2(n9200), .A3(n9199), .A4(n9198), .ZN(n13873)
         );
  AND2_X1 U8952 ( .A1(n6702), .A2(n12101), .ZN(n6458) );
  AND2_X1 U8953 ( .A1(n9239), .A2(n11990), .ZN(n6459) );
  NAND2_X1 U8954 ( .A1(n9634), .A2(n13860), .ZN(n6959) );
  XOR2_X1 U8955 ( .A(n12456), .B(n12455), .Z(n6460) );
  OR2_X1 U8956 ( .A1(n7219), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6461) );
  AND2_X1 U8957 ( .A1(n7344), .A2(n6638), .ZN(n6462) );
  AND2_X1 U8958 ( .A1(n7261), .A2(n13336), .ZN(n6463) );
  INV_X1 U8959 ( .A(n7264), .ZN(n7263) );
  NOR2_X1 U8960 ( .A1(n11155), .A2(n7265), .ZN(n7264) );
  OR2_X1 U8961 ( .A1(n8822), .A2(n8389), .ZN(n6464) );
  INV_X1 U8962 ( .A(n8673), .ZN(n7538) );
  AND2_X1 U8963 ( .A1(n11653), .A2(n11650), .ZN(n6465) );
  AND3_X1 U8964 ( .A1(n9190), .A2(n7436), .A3(n9206), .ZN(n6466) );
  NAND2_X1 U8965 ( .A1(n8105), .A2(n8104), .ZN(n12350) );
  INV_X1 U8966 ( .A(n12350), .ZN(n12507) );
  AND2_X1 U8967 ( .A1(n6454), .A2(n7180), .ZN(n6467) );
  AND2_X1 U8968 ( .A1(n11687), .A2(n11688), .ZN(n12683) );
  INV_X1 U8969 ( .A(n12683), .ZN(n7005) );
  NAND2_X1 U8970 ( .A1(n12963), .A2(n12968), .ZN(n7342) );
  NAND2_X1 U8971 ( .A1(n8081), .A2(n6579), .ZN(n12511) );
  INV_X1 U8972 ( .A(n12511), .ZN(n7400) );
  INV_X1 U8973 ( .A(n14183), .ZN(n7100) );
  NAND2_X1 U8974 ( .A1(n8425), .A2(n6452), .ZN(n6468) );
  AND2_X1 U8975 ( .A1(n9167), .A2(n8449), .ZN(n9158) );
  NAND2_X1 U8976 ( .A1(n8681), .A2(n8680), .ZN(n11380) );
  INV_X1 U8977 ( .A(n11380), .ZN(n7141) );
  AND2_X1 U8978 ( .A1(n14958), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6469) );
  AND2_X1 U8979 ( .A1(n12438), .A2(n7168), .ZN(n6470) );
  NAND2_X1 U8980 ( .A1(n8111), .A2(n8110), .ZN(n12482) );
  OR2_X1 U8981 ( .A1(n14435), .A2(n12434), .ZN(n6471) );
  NAND2_X1 U8982 ( .A1(n9378), .A2(n9377), .ZN(n14233) );
  AND2_X1 U8983 ( .A1(n13516), .A2(n13100), .ZN(n6472) );
  AND2_X1 U8984 ( .A1(n8134), .A2(n7655), .ZN(n8141) );
  OR2_X1 U8985 ( .A1(n10371), .A2(n10370), .ZN(n6473) );
  NAND2_X2 U8986 ( .A1(n11811), .A2(n9606), .ZN(n10692) );
  AND2_X1 U8987 ( .A1(n6680), .A2(n6679), .ZN(n6474) );
  NAND2_X1 U8988 ( .A1(n7914), .A2(n7913), .ZN(n7916) );
  NAND2_X1 U8989 ( .A1(n8141), .A2(n7582), .ZN(n6475) );
  OR2_X1 U8990 ( .A1(n7975), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6476) );
  INV_X1 U8991 ( .A(n12920), .ZN(n7341) );
  NAND2_X1 U8992 ( .A1(n8070), .A2(n8069), .ZN(n12525) );
  XNOR2_X1 U8993 ( .A(n13472), .B(n13241), .ZN(n13226) );
  INV_X1 U8994 ( .A(n13226), .ZN(n7250) );
  NAND2_X1 U8995 ( .A1(n8141), .A2(n7581), .ZN(n8202) );
  AND2_X1 U8996 ( .A1(n12905), .A2(n6456), .ZN(n6477) );
  NOR2_X1 U8997 ( .A1(n12014), .A2(n12020), .ZN(n6478) );
  AND2_X1 U8998 ( .A1(n8414), .A2(n7490), .ZN(n7487) );
  NAND2_X1 U8999 ( .A1(n9551), .A2(n9550), .ZN(n14252) );
  INV_X1 U9000 ( .A(n12207), .ZN(n7206) );
  OR2_X1 U9001 ( .A1(n8820), .A2(SI_14_), .ZN(n6479) );
  AND2_X1 U9002 ( .A1(n8588), .A2(n8587), .ZN(n6480) );
  OR2_X1 U9003 ( .A1(n11895), .A2(n7592), .ZN(n6481) );
  INV_X1 U9004 ( .A(n7429), .ZN(n14083) );
  NAND2_X1 U9005 ( .A1(n7433), .A2(n7432), .ZN(n7429) );
  NAND2_X1 U9006 ( .A1(n13812), .A2(n13811), .ZN(n13655) );
  AND2_X1 U9007 ( .A1(n9031), .A2(n9030), .ZN(n6482) );
  NOR2_X1 U9008 ( .A1(n7719), .A2(n7575), .ZN(n7735) );
  OAI21_X1 U9009 ( .B1(n7791), .B2(n7790), .A(n7792), .ZN(n7806) );
  AND2_X1 U9010 ( .A1(n12400), .A2(n12399), .ZN(n6483) );
  XOR2_X1 U9011 ( .A(n12205), .B(n12490), .Z(n6484) );
  AND2_X1 U9012 ( .A1(n7355), .A2(n6765), .ZN(n6485) );
  OR2_X1 U9013 ( .A1(n9863), .A2(n13890), .ZN(n6486) );
  INV_X1 U9014 ( .A(n7446), .ZN(n7445) );
  AND2_X1 U9015 ( .A1(n7447), .A2(n10861), .ZN(n7446) );
  AND2_X1 U9016 ( .A1(n14111), .A2(n9466), .ZN(n6487) );
  INV_X1 U9017 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7312) );
  AND2_X1 U9018 ( .A1(n8426), .A2(n8427), .ZN(n6488) );
  OR3_X1 U9019 ( .A1(n11911), .A2(n11910), .A3(n11919), .ZN(n6489) );
  OR2_X1 U9020 ( .A1(n8493), .A2(n14766), .ZN(n6490) );
  INV_X1 U9021 ( .A(n13859), .ZN(n13786) );
  INV_X1 U9022 ( .A(n8358), .ZN(n6726) );
  XNOR2_X1 U9023 ( .A(n14264), .B(n13859), .ZN(n14027) );
  INV_X1 U9024 ( .A(n8365), .ZN(n7091) );
  INV_X1 U9025 ( .A(n14208), .ZN(n7133) );
  NAND2_X1 U9026 ( .A1(n8617), .A2(n8616), .ZN(n10942) );
  INV_X1 U9027 ( .A(n10503), .ZN(n12055) );
  AND2_X1 U9028 ( .A1(n14467), .A2(n12193), .ZN(n6491) );
  INV_X1 U9029 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7671) );
  AND2_X1 U9030 ( .A1(n9312), .A2(n9311), .ZN(n11873) );
  INV_X1 U9031 ( .A(n11873), .ZN(n7189) );
  NAND2_X1 U9032 ( .A1(n9539), .A2(n9538), .ZN(n14022) );
  INV_X1 U9033 ( .A(n14022), .ZN(n7181) );
  INV_X1 U9034 ( .A(n12062), .ZN(n7455) );
  AND2_X1 U9035 ( .A1(n9423), .A2(n9422), .ZN(n14311) );
  INV_X1 U9036 ( .A(n14311), .ZN(n7184) );
  AND2_X1 U9037 ( .A1(n12489), .A2(n11748), .ZN(n6492) );
  NAND2_X1 U9038 ( .A1(n8766), .A2(n8765), .ZN(n13434) );
  INV_X1 U9039 ( .A(n11965), .ZN(n6829) );
  AND2_X1 U9040 ( .A1(n11232), .A2(n13108), .ZN(n6493) );
  AND3_X1 U9041 ( .A1(n9402), .A2(n9183), .A3(n9182), .ZN(n6494) );
  INV_X1 U9042 ( .A(n7071), .ZN(n7070) );
  NOR2_X1 U9043 ( .A1(n9629), .A2(n14029), .ZN(n7071) );
  NAND2_X1 U9044 ( .A1(n6713), .A2(SI_1_), .ZN(n8345) );
  NAND2_X1 U9045 ( .A1(n14089), .A2(n13821), .ZN(n6495) );
  INV_X1 U9046 ( .A(n7473), .ZN(n9117) );
  OR2_X1 U9047 ( .A1(n8309), .A2(n8310), .ZN(n6496) );
  AND4_X1 U9048 ( .A1(n7355), .A2(n6765), .A3(n6494), .A4(n9181), .ZN(n6497)
         );
  NAND4_X1 U9049 ( .A1(n8521), .A2(n8489), .A3(n7313), .A4(n7312), .ZN(n8562)
         );
  OR2_X1 U9050 ( .A1(n13477), .A2(n13259), .ZN(n6498) );
  XNOR2_X1 U9051 ( .A(n12119), .B(n12118), .ZN(n7656) );
  INV_X1 U9052 ( .A(n11882), .ZN(n14554) );
  NAND2_X1 U9053 ( .A1(n9349), .A2(n9348), .ZN(n11882) );
  AND2_X1 U9054 ( .A1(n14358), .A2(n9863), .ZN(n14283) );
  NAND2_X1 U9055 ( .A1(n9209), .A2(n9224), .ZN(n9233) );
  NAND2_X1 U9056 ( .A1(n8519), .A2(n8521), .ZN(n8538) );
  NOR2_X1 U9057 ( .A1(n14244), .A2(n14202), .ZN(n6499) );
  INV_X1 U9058 ( .A(n7381), .ZN(n7380) );
  OAI21_X1 U9059 ( .B1(n7383), .B2(n7384), .A(n7382), .ZN(n7381) );
  INV_X1 U9060 ( .A(n6889), .ZN(n13287) );
  AND2_X1 U9061 ( .A1(n12205), .A2(n12328), .ZN(n6500) );
  AND2_X1 U9062 ( .A1(n13296), .A2(n7257), .ZN(n6501) );
  NAND2_X1 U9063 ( .A1(n7605), .A2(n7603), .ZN(n7599) );
  NAND2_X1 U9064 ( .A1(n14055), .A2(n6454), .ZN(n7182) );
  AND2_X1 U9065 ( .A1(n12945), .A2(n6940), .ZN(n6502) );
  AND2_X1 U9066 ( .A1(n7602), .A2(n7600), .ZN(n6503) );
  INV_X1 U9067 ( .A(n11938), .ZN(n6836) );
  OR2_X1 U9068 ( .A1(n10779), .A2(n10778), .ZN(n6504) );
  AND2_X1 U9069 ( .A1(n7045), .A2(n11381), .ZN(n6505) );
  AND2_X1 U9070 ( .A1(n6799), .A2(n6796), .ZN(n6506) );
  INV_X1 U9071 ( .A(n7305), .ZN(n7304) );
  OAI22_X1 U9072 ( .A1(n7307), .A2(n7306), .B1(n12808), .B2(n12564), .ZN(n7305) );
  AND2_X1 U9073 ( .A1(n7301), .A2(n8190), .ZN(n6507) );
  AND2_X1 U9074 ( .A1(n7326), .A2(n7331), .ZN(n6508) );
  OR2_X1 U9075 ( .A1(n9686), .A2(n12210), .ZN(n11781) );
  INV_X1 U9076 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7556) );
  INV_X1 U9077 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8427) );
  OR2_X1 U9078 ( .A1(n13112), .A2(n14931), .ZN(n6509) );
  AND2_X1 U9079 ( .A1(n7641), .A2(n6829), .ZN(n6510) );
  AND2_X1 U9080 ( .A1(n11668), .A2(n11669), .ZN(n11761) );
  INV_X1 U9081 ( .A(n11761), .ZN(n8166) );
  NOR2_X1 U9082 ( .A1(n14410), .A2(n14527), .ZN(n6511) );
  NOR2_X1 U9083 ( .A1(n12837), .A2(n12250), .ZN(n6512) );
  NOR2_X1 U9084 ( .A1(n12313), .A2(n12589), .ZN(n6513) );
  INV_X1 U9085 ( .A(n7578), .ZN(n7006) );
  AND2_X1 U9086 ( .A1(n11693), .A2(n11687), .ZN(n7578) );
  OR2_X1 U9087 ( .A1(n7593), .A2(n7589), .ZN(n6514) );
  INV_X1 U9088 ( .A(n12079), .ZN(n7439) );
  NOR2_X1 U9089 ( .A1(n7071), .A2(n7067), .ZN(n6515) );
  AND3_X1 U9090 ( .A1(n9221), .A2(n9219), .A3(n9220), .ZN(n6516) );
  OR2_X1 U9091 ( .A1(n6781), .A2(n6438), .ZN(n6517) );
  NAND2_X1 U9092 ( .A1(n7208), .A2(n12156), .ZN(n6518) );
  OR2_X1 U9093 ( .A1(n8251), .A2(n8252), .ZN(n6519) );
  NOR2_X1 U9094 ( .A1(n13538), .A2(n13423), .ZN(n6520) );
  OR2_X1 U9095 ( .A1(n12298), .A2(n12353), .ZN(n6521) );
  AND2_X1 U9096 ( .A1(n11751), .A2(n11749), .ZN(n12206) );
  AND2_X1 U9097 ( .A1(n12213), .A2(n12349), .ZN(n6522) );
  NOR2_X1 U9098 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n8519) );
  INV_X1 U9099 ( .A(n7486), .ZN(n8978) );
  NAND2_X1 U9100 ( .A1(n8414), .A2(n8413), .ZN(n7486) );
  NAND2_X1 U9101 ( .A1(n7550), .A2(n7552), .ZN(n7549) );
  AND2_X1 U9102 ( .A1(n11276), .A2(n11275), .ZN(n6523) );
  AND2_X1 U9103 ( .A1(n11711), .A2(n11714), .ZN(n12601) );
  INV_X1 U9104 ( .A(n12601), .ZN(n7296) );
  AND2_X1 U9105 ( .A1(n11756), .A2(n11622), .ZN(n11784) );
  AND2_X1 U9106 ( .A1(n7481), .A2(n6479), .ZN(n6524) );
  NAND2_X1 U9107 ( .A1(n9515), .A2(n7432), .ZN(n6525) );
  NAND2_X1 U9108 ( .A1(n6624), .A2(SI_9_), .ZN(n6526) );
  INV_X1 U9109 ( .A(n7421), .ZN(n7420) );
  NAND2_X1 U9110 ( .A1(n14219), .A2(n9371), .ZN(n7421) );
  OR2_X1 U9111 ( .A1(n6482), .A2(n6979), .ZN(n6527) );
  AND2_X1 U9112 ( .A1(n8449), .A2(n11586), .ZN(n8474) );
  INV_X1 U9113 ( .A(n8474), .ZN(n7348) );
  AND2_X1 U9114 ( .A1(n12170), .A2(n12507), .ZN(n6528) );
  INV_X1 U9115 ( .A(n7122), .ZN(n7121) );
  NOR2_X1 U9116 ( .A1(n14554), .A2(n11552), .ZN(n7122) );
  INV_X1 U9117 ( .A(n11966), .ZN(n7642) );
  AND2_X1 U9118 ( .A1(n12358), .A2(n11293), .ZN(n6529) );
  AND2_X1 U9119 ( .A1(n7425), .A2(n7423), .ZN(n6530) );
  NAND2_X1 U9120 ( .A1(n6498), .A2(n7254), .ZN(n6531) );
  INV_X1 U9121 ( .A(n6802), .ZN(n6801) );
  NAND2_X1 U9122 ( .A1(n10609), .A2(n10610), .ZN(n6802) );
  INV_X1 U9123 ( .A(n7363), .ZN(n7362) );
  NAND2_X1 U9124 ( .A1(n7364), .A2(n13654), .ZN(n7363) );
  INV_X1 U9125 ( .A(n7140), .ZN(n7139) );
  NAND2_X1 U9126 ( .A1(n9548), .A2(n9537), .ZN(n7140) );
  OR2_X1 U9127 ( .A1(n12461), .A2(n11624), .ZN(n11756) );
  NAND2_X1 U9128 ( .A1(n11872), .A2(n7610), .ZN(n6532) );
  OR2_X1 U9129 ( .A1(n8493), .A2(n10079), .ZN(n6533) );
  XNOR2_X1 U9130 ( .A(n7365), .B(P1_IR_REG_21__SCAN_IN), .ZN(n11970) );
  AND2_X1 U9131 ( .A1(n7200), .A2(n7206), .ZN(n6534) );
  NAND3_X1 U9132 ( .A1(n6906), .A2(n9214), .A3(n9216), .ZN(n13874) );
  AND3_X1 U9133 ( .A1(n7711), .A2(n7710), .A3(n7709), .ZN(n12780) );
  AND2_X1 U9134 ( .A1(n8629), .A2(n8610), .ZN(n6535) );
  OAI21_X1 U9135 ( .B1(n8366), .B2(n7092), .A(n7089), .ZN(n8674) );
  INV_X1 U9136 ( .A(n8741), .ZN(n7481) );
  AND2_X1 U9137 ( .A1(n7337), .A2(n7342), .ZN(n6536) );
  OR2_X1 U9138 ( .A1(n6441), .A2(SI_10_), .ZN(n6537) );
  OR2_X1 U9139 ( .A1(n6441), .A2(n9829), .ZN(n6538) );
  INV_X1 U9140 ( .A(n7333), .ZN(n7332) );
  AND2_X1 U9141 ( .A1(n13048), .A2(n6436), .ZN(n6539) );
  NOR2_X1 U9142 ( .A1(n7609), .A2(n7608), .ZN(n6540) );
  AND2_X1 U9143 ( .A1(n11375), .A2(n10936), .ZN(n6541) );
  INV_X1 U9144 ( .A(n9264), .ZN(n7112) );
  AND2_X1 U9145 ( .A1(n9186), .A2(n6466), .ZN(n6542) );
  AND2_X1 U9146 ( .A1(n11045), .A2(n11042), .ZN(n6543) );
  AND2_X1 U9147 ( .A1(n6488), .A2(n7556), .ZN(n6544) );
  NAND2_X1 U9148 ( .A1(n11757), .A2(n15084), .ZN(n6545) );
  AND2_X1 U9149 ( .A1(n6855), .A2(n6854), .ZN(n6546) );
  AND2_X1 U9150 ( .A1(n7456), .A2(n7053), .ZN(n6547) );
  OR2_X1 U9151 ( .A1(n13492), .A2(n13040), .ZN(n6548) );
  INV_X1 U9152 ( .A(n14252), .ZN(n14006) );
  AND2_X1 U9153 ( .A1(n6455), .A2(n7101), .ZN(n6549) );
  INV_X1 U9154 ( .A(n6959), .ZN(n6958) );
  INV_X1 U9155 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9203) );
  INV_X1 U9156 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U9157 ( .A1(n13487), .A2(n12080), .ZN(n6550) );
  OR2_X1 U9158 ( .A1(n6890), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6551) );
  OR2_X1 U9159 ( .A1(n7540), .A2(n6480), .ZN(n6552) );
  OR2_X1 U9160 ( .A1(n7538), .A2(n6557), .ZN(n6553) );
  INV_X1 U9161 ( .A(n7295), .ZN(n7294) );
  NAND2_X1 U9162 ( .A1(n7296), .A2(n8177), .ZN(n7295) );
  INV_X1 U9163 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9190) );
  INV_X1 U9164 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9586) );
  INV_X1 U9165 ( .A(n14525), .ZN(n6791) );
  INV_X1 U9166 ( .A(n9693), .ZN(n9167) );
  NAND2_X1 U9167 ( .A1(n13086), .A2(n12871), .ZN(n6647) );
  INV_X1 U9168 ( .A(n13028), .ZN(n6640) );
  AND2_X1 U9169 ( .A1(n11727), .A2(n11728), .ZN(n12561) );
  INV_X1 U9170 ( .A(n12561), .ZN(n7307) );
  NAND2_X1 U9171 ( .A1(n8917), .A2(n8916), .ZN(n13325) );
  INV_X1 U9172 ( .A(n13325), .ZN(n7261) );
  INV_X1 U9173 ( .A(n13487), .ZN(n6888) );
  NAND2_X1 U9174 ( .A1(n9001), .A2(n9000), .ZN(n13482) );
  INV_X1 U9175 ( .A(n13482), .ZN(n7255) );
  AND2_X1 U9176 ( .A1(n14209), .A2(n7183), .ZN(n6554) );
  OR2_X1 U9177 ( .A1(n14135), .A2(n14134), .ZN(n14133) );
  INV_X1 U9178 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6901) );
  AND2_X1 U9179 ( .A1(n12166), .A2(n12167), .ZN(n6555) );
  OAI21_X1 U9180 ( .B1(n9372), .B2(n7130), .A(n7129), .ZN(n14187) );
  NAND2_X1 U9181 ( .A1(n7287), .A2(n7286), .ZN(n14465) );
  NAND2_X1 U9182 ( .A1(n7116), .A2(n7115), .ZN(n11498) );
  INV_X1 U9183 ( .A(n11692), .ZN(n7004) );
  AND3_X1 U9184 ( .A1(n8063), .A2(n8062), .A3(n8061), .ZN(n12549) );
  INV_X1 U9185 ( .A(n11703), .ZN(n7001) );
  NAND2_X1 U9186 ( .A1(n6786), .A2(n11893), .ZN(n14203) );
  OAI21_X1 U9187 ( .B1(n12926), .B2(n13422), .A(n12087), .ZN(n12088) );
  NAND2_X1 U9188 ( .A1(n13858), .A2(n14619), .ZN(n6556) );
  NAND2_X1 U9189 ( .A1(n9570), .A2(n9569), .ZN(n14247) );
  INV_X1 U9190 ( .A(n14247), .ZN(n7180) );
  NAND2_X1 U9191 ( .A1(n9372), .A2(n9371), .ZN(n14234) );
  AND2_X1 U9192 ( .A1(n8672), .A2(n8671), .ZN(n6557) );
  AND2_X1 U9193 ( .A1(n13533), .A2(n13103), .ZN(n6558) );
  INV_X1 U9194 ( .A(n6766), .ZN(n9420) );
  AND2_X1 U9195 ( .A1(n7370), .A2(n7371), .ZN(n6559) );
  INV_X1 U9196 ( .A(n12132), .ZN(n7214) );
  INV_X1 U9197 ( .A(n6887), .ZN(n13365) );
  AND2_X1 U9198 ( .A1(n14193), .A2(n11901), .ZN(n6560) );
  INV_X1 U9199 ( .A(n7177), .ZN(n14114) );
  NOR2_X1 U9200 ( .A1(n14136), .A2(n14288), .ZN(n7177) );
  OR2_X1 U9201 ( .A1(n8892), .A2(n6450), .ZN(n6561) );
  AND2_X1 U9202 ( .A1(n12263), .A2(n12265), .ZN(n6562) );
  INV_X1 U9203 ( .A(n7149), .ZN(n13354) );
  AND2_X1 U9204 ( .A1(n6887), .A2(n6597), .ZN(n7149) );
  AND2_X1 U9205 ( .A1(n12612), .A2(n7294), .ZN(n6563) );
  INV_X1 U9206 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10125) );
  INV_X1 U9207 ( .A(n8893), .ZN(n8403) );
  AND2_X1 U9208 ( .A1(n7824), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6564) );
  INV_X1 U9209 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7313) );
  AND2_X1 U9210 ( .A1(n7892), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6565) );
  OR2_X1 U9211 ( .A1(n6441), .A2(SI_11_), .ZN(n6566) );
  AND2_X1 U9212 ( .A1(n14542), .A2(n9386), .ZN(n6567) );
  INV_X1 U9213 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6626) );
  AND2_X1 U9214 ( .A1(n14180), .A2(n9626), .ZN(n6568) );
  AND2_X1 U9215 ( .A1(n7418), .A2(n7874), .ZN(n6569) );
  OR2_X1 U9216 ( .A1(n7613), .A2(n11883), .ZN(n6570) );
  AND2_X1 U9217 ( .A1(n12929), .A2(n12928), .ZN(n6571) );
  NAND2_X1 U9218 ( .A1(n8892), .A2(n6450), .ZN(n6572) );
  AND2_X1 U9219 ( .A1(n6882), .A2(n6890), .ZN(n6573) );
  INV_X1 U9220 ( .A(n14375), .ZN(n11241) );
  NAND2_X1 U9221 ( .A1(n6459), .A2(n10733), .ZN(n10555) );
  AND2_X1 U9222 ( .A1(n8238), .A2(n8237), .ZN(n15137) );
  NAND2_X1 U9223 ( .A1(n9352), .A2(n9351), .ZN(n14410) );
  INV_X1 U9224 ( .A(n14410), .ZN(n7185) );
  NAND2_X1 U9225 ( .A1(n8749), .A2(n8748), .ZN(n13543) );
  INV_X1 U9226 ( .A(n13543), .ZN(n6590) );
  NAND2_X1 U9227 ( .A1(n9434), .A2(n9433), .ZN(n14306) );
  INV_X1 U9228 ( .A(n14306), .ZN(n7101) );
  OAI211_X1 U9229 ( .C1(n6438), .C2(n6782), .A(n6517), .B(n7623), .ZN(n10801)
         );
  AND2_X1 U9230 ( .A1(n14629), .A2(n7188), .ZN(n6574) );
  NOR2_X1 U9231 ( .A1(n6442), .A2(n15195), .ZN(n6575) );
  NAND2_X1 U9232 ( .A1(n8881), .A2(n8880), .ZN(n13516) );
  INV_X1 U9233 ( .A(n13516), .ZN(n6597) );
  NAND2_X1 U9234 ( .A1(n7569), .A2(n11668), .ZN(n11220) );
  NAND2_X1 U9235 ( .A1(n8828), .A2(n8827), .ZN(n13538) );
  INV_X1 U9236 ( .A(n13538), .ZN(n7143) );
  NAND2_X1 U9237 ( .A1(n12459), .A2(n10536), .ZN(n10538) );
  NAND2_X1 U9238 ( .A1(n8898), .A2(n8897), .ZN(n13511) );
  INV_X1 U9239 ( .A(n13511), .ZN(n7148) );
  INV_X1 U9240 ( .A(n8979), .ZN(n7485) );
  OR2_X1 U9241 ( .A1(n14761), .A2(n9564), .ZN(n6576) );
  INV_X1 U9242 ( .A(n8953), .ZN(n7496) );
  OR2_X1 U9243 ( .A1(n14751), .A2(n9563), .ZN(n6577) );
  OR2_X1 U9244 ( .A1(n6441), .A2(n10516), .ZN(n6578) );
  OR2_X1 U9245 ( .A1(n6441), .A2(n7493), .ZN(n6579) );
  OR2_X1 U9246 ( .A1(n6441), .A2(n11449), .ZN(n6580) );
  AND2_X1 U9247 ( .A1(n10611), .A2(n6801), .ZN(n6581) );
  OR2_X1 U9248 ( .A1(n14982), .A2(n11079), .ZN(n6857) );
  INV_X1 U9249 ( .A(n6675), .ZN(n6674) );
  NOR2_X1 U9250 ( .A1(n12399), .A2(n12414), .ZN(n6675) );
  AND2_X1 U9251 ( .A1(n6680), .A2(n6678), .ZN(n6582) );
  NOR2_X1 U9252 ( .A1(n6442), .A2(n12124), .ZN(n6583) );
  INV_X1 U9253 ( .A(SI_18_), .ZN(n10142) );
  AND2_X1 U9254 ( .A1(n7409), .A2(n8039), .ZN(n6584) );
  AND2_X1 U9255 ( .A1(n12128), .A2(n12127), .ZN(n6585) );
  OR2_X1 U9256 ( .A1(n7496), .A2(n10856), .ZN(n6586) );
  AND2_X1 U9257 ( .A1(n7495), .A2(n7497), .ZN(n6587) );
  AND2_X1 U9258 ( .A1(n7491), .A2(n7492), .ZN(n7488) );
  AND2_X1 U9259 ( .A1(n14878), .A2(n9788), .ZN(n14930) );
  INV_X1 U9260 ( .A(n14930), .ZN(n14953) );
  INV_X1 U9261 ( .A(n15029), .ZN(n6609) );
  AND2_X2 U9262 ( .A1(n10874), .A2(n10309), .ZN(n14974) );
  XNOR2_X1 U9263 ( .A(n13114), .B(n10819), .ZN(n10817) );
  AND2_X2 U9264 ( .A1(n10874), .A2(n14894), .ZN(n14959) );
  INV_X1 U9265 ( .A(n10843), .ZN(n6593) );
  INV_X1 U9266 ( .A(n15009), .ZN(n6856) );
  INV_X1 U9267 ( .A(n14447), .ZN(n6931) );
  INV_X1 U9268 ( .A(n9732), .ZN(n7320) );
  AND2_X1 U9269 ( .A1(n10733), .A2(n9239), .ZN(n6588) );
  OR2_X1 U9270 ( .A1(n6931), .A2(n14432), .ZN(n6589) );
  INV_X1 U9271 ( .A(SI_25_), .ZN(n7493) );
  INV_X1 U9272 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6965) );
  AOI22_X1 U9273 ( .A1(n13227), .A2(n13441), .B1(n13444), .B2(n13259), .ZN(
        n7465) );
  OAI22_X1 U9274 ( .A1(n10569), .A2(n10568), .B1(n10567), .B2(n10577), .ZN(
        n10770) );
  NAND2_X1 U9275 ( .A1(n10577), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7171) );
  INV_X2 U9276 ( .A(n14759), .ZN(n14761) );
  NOR2_X2 U9277 ( .A1(n11386), .A2(n13549), .ZN(n11465) );
  AND2_X2 U9278 ( .A1(n10869), .A2(n14856), .ZN(n10952) );
  NOR2_X1 U9279 ( .A1(n10960), .A2(n10965), .ZN(n10869) );
  OAI21_X1 U9280 ( .B1(n13463), .B2(n14958), .A(n6595), .ZN(n6596) );
  INV_X1 U9281 ( .A(n6596), .ZN(n7046) );
  NOR2_X2 U9282 ( .A1(n13338), .A2(n13325), .ZN(n7147) );
  NOR2_X2 U9283 ( .A1(n13273), .A2(n13482), .ZN(n13263) );
  INV_X2 U9284 ( .A(n14906), .ZN(n10297) );
  INV_X1 U9285 ( .A(n14866), .ZN(n7145) );
  AND2_X2 U9286 ( .A1(n6633), .A2(n6533), .ZN(n14906) );
  NAND2_X1 U9287 ( .A1(n6606), .A2(n11704), .ZN(n12632) );
  NAND3_X1 U9288 ( .A1(n6608), .A2(n11763), .A3(n6607), .ZN(n7795) );
  NAND3_X1 U9289 ( .A1(n7744), .A2(n11661), .A3(n6465), .ZN(n6607) );
  AOI21_X1 U9290 ( .B1(n12050), .B2(n15102), .A(n9668), .ZN(n7276) );
  NAND2_X1 U9291 ( .A1(n11657), .A2(n11661), .ZN(n11332) );
  NAND3_X1 U9292 ( .A1(n6614), .A2(n6613), .A3(n7488), .ZN(n9019) );
  OAI21_X1 U9293 ( .B1(n7072), .B2(n8405), .A(n6615), .ZN(n8408) );
  NAND2_X1 U9294 ( .A1(n8370), .A2(n6619), .ZN(n6618) );
  NAND3_X1 U9295 ( .A1(n7028), .A2(n8410), .A3(n7497), .ZN(n8937) );
  NAND3_X1 U9296 ( .A1(n7028), .A2(n8410), .A3(n6587), .ZN(n6621) );
  NAND2_X1 U9297 ( .A1(n8410), .A2(n6586), .ZN(n6623) );
  NAND4_X1 U9298 ( .A1(n6631), .A2(n7688), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n6629) );
  NAND4_X1 U9299 ( .A1(n13193), .A2(n7687), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n7686), .ZN(n6630) );
  NAND2_X2 U9300 ( .A1(n8493), .A2(n9833), .ZN(n8518) );
  NAND3_X1 U9301 ( .A1(n6644), .A2(n6642), .A3(n6641), .ZN(n10930) );
  NAND3_X1 U9302 ( .A1(n10679), .A2(n7321), .A3(n7323), .ZN(n6641) );
  OAI21_X1 U9303 ( .B1(n7318), .B2(n9732), .A(n9737), .ZN(n6643) );
  NAND3_X1 U9304 ( .A1(n10523), .A2(n6645), .A3(n10679), .ZN(n6644) );
  NOR2_X1 U9305 ( .A1(n7322), .A2(n6646), .ZN(n6645) );
  NAND2_X1 U9306 ( .A1(n10523), .A2(n9721), .ZN(n10507) );
  INV_X1 U9307 ( .A(n9721), .ZN(n6646) );
  NAND2_X1 U9308 ( .A1(n6647), .A2(n12875), .ZN(n12994) );
  NAND3_X1 U9309 ( .A1(n6650), .A2(n6649), .A3(n6648), .ZN(n10525) );
  NAND3_X1 U9310 ( .A1(n13050), .A2(n9715), .A3(n13051), .ZN(n6649) );
  NAND2_X1 U9311 ( .A1(n10518), .A2(n9715), .ZN(n6650) );
  XNOR2_X2 U9312 ( .A(n6652), .B(P2_IR_REG_28__SCAN_IN), .ZN(n9159) );
  INV_X2 U9313 ( .A(n8784), .ZN(n8425) );
  NAND2_X1 U9314 ( .A1(n11430), .A2(n6653), .ZN(n12866) );
  NAND3_X1 U9315 ( .A1(n9738), .A2(n9739), .A3(n6655), .ZN(n11147) );
  NAND3_X1 U9316 ( .A1(n6918), .A2(n6658), .A3(n6656), .ZN(P3_U3201) );
  AND2_X1 U9317 ( .A1(n10768), .A2(n10779), .ZN(n6665) );
  NAND2_X1 U9318 ( .A1(n10470), .A2(n10471), .ZN(n6666) );
  INV_X1 U9319 ( .A(n12400), .ZN(n6671) );
  NAND3_X1 U9320 ( .A1(n6670), .A2(n6674), .A3(n6668), .ZN(n12401) );
  NAND3_X1 U9321 ( .A1(n6670), .A2(n6669), .A3(n6668), .ZN(n6677) );
  INV_X1 U9322 ( .A(n6677), .ZN(n12413) );
  NOR2_X1 U9323 ( .A1(n6681), .A2(n11064), .ZN(n6679) );
  NAND2_X1 U9324 ( .A1(n14985), .A2(n6682), .ZN(n6680) );
  NAND2_X1 U9325 ( .A1(n6688), .A2(n7723), .ZN(n7739) );
  NAND2_X1 U9326 ( .A1(n7722), .A2(n7721), .ZN(n6688) );
  OAI21_X1 U9327 ( .B1(n7722), .B2(n6691), .A(n6689), .ZN(n7741) );
  INV_X1 U9328 ( .A(n6690), .ZN(n6689) );
  INV_X1 U9329 ( .A(n7723), .ZN(n6691) );
  NAND2_X1 U9330 ( .A1(n7387), .A2(n7691), .ZN(n7722) );
  NAND2_X1 U9331 ( .A1(n7893), .A2(n6565), .ZN(n6698) );
  OAI211_X1 U9332 ( .C1(n6707), .C2(n11378), .A(n6705), .B(n11377), .ZN(n11452) );
  NAND3_X1 U9333 ( .A1(n7264), .A2(n10937), .A3(n6541), .ZN(n6705) );
  NAND2_X1 U9334 ( .A1(n6706), .A2(n6707), .ZN(n11376) );
  OR2_X1 U9335 ( .A1(n7263), .A2(n10938), .ZN(n6706) );
  INV_X1 U9336 ( .A(n6708), .ZN(n7256) );
  NAND2_X1 U9337 ( .A1(n6716), .A2(n6945), .ZN(n6713) );
  NAND3_X1 U9338 ( .A1(n8345), .A2(n6717), .A3(n8483), .ZN(n8487) );
  AND2_X1 U9339 ( .A1(n6715), .A2(n6714), .ZN(n8483) );
  AOI21_X1 U9340 ( .B1(n6437), .B2(n8491), .A(n9831), .ZN(n6714) );
  NAND2_X1 U9341 ( .A1(n8345), .A2(n6717), .ZN(n8485) );
  NAND3_X1 U9342 ( .A1(n6716), .A2(n6945), .A3(n6718), .ZN(n6717) );
  INV_X1 U9343 ( .A(SI_1_), .ZN(n6718) );
  NAND2_X1 U9344 ( .A1(n8561), .A2(n8356), .ZN(n8580) );
  NAND2_X1 U9345 ( .A1(n8561), .A2(n6724), .ZN(n6723) );
  AND2_X1 U9346 ( .A1(n8359), .A2(n8356), .ZN(n6724) );
  INV_X1 U9347 ( .A(n8359), .ZN(n6725) );
  NAND2_X1 U9348 ( .A1(n8582), .A2(n8359), .ZN(n8591) );
  NAND2_X1 U9349 ( .A1(n8580), .A2(n6726), .ZN(n8582) );
  NAND2_X1 U9350 ( .A1(n6729), .A2(n7501), .ZN(n8659) );
  NAND2_X1 U9351 ( .A1(n11454), .A2(n11453), .ZN(n12094) );
  OAI21_X1 U9352 ( .B1(n13254), .B2(n12114), .A(n7254), .ZN(n13249) );
  NAND2_X2 U9353 ( .A1(n6732), .A2(n6737), .ZN(n15068) );
  NAND2_X2 U9354 ( .A1(n7676), .A2(n7677), .ZN(n8029) );
  NAND2_X2 U9355 ( .A1(n7676), .A2(n12862), .ZN(n11604) );
  AND2_X1 U9356 ( .A1(n7704), .A2(n6734), .ZN(n6732) );
  NAND3_X2 U9357 ( .A1(n6738), .A2(n7176), .A3(n7660), .ZN(n7719) );
  NAND2_X1 U9358 ( .A1(n6745), .A2(n12247), .ZN(n12258) );
  NAND2_X1 U9359 ( .A1(n12285), .A2(n12283), .ZN(n12141) );
  XNOR2_X1 U9360 ( .A(n6761), .B(n12549), .ZN(n12188) );
  NAND2_X1 U9361 ( .A1(n14401), .A2(n12000), .ZN(n6762) );
  NAND2_X1 U9362 ( .A1(n11345), .A2(n9621), .ZN(n6763) );
  INV_X1 U9363 ( .A(n11027), .ZN(n6764) );
  NAND2_X1 U9364 ( .A1(n9618), .A2(n14615), .ZN(n14624) );
  NAND3_X1 U9365 ( .A1(n6485), .A2(n6448), .A3(n6767), .ZN(n6766) );
  NAND3_X1 U9366 ( .A1(n6497), .A2(n9186), .A3(n6448), .ZN(n9575) );
  NAND2_X1 U9367 ( .A1(n14078), .A2(n6771), .ZN(n6769) );
  INV_X1 U9368 ( .A(n14046), .ZN(n6774) );
  INV_X1 U9369 ( .A(n6780), .ZN(n14102) );
  NAND2_X1 U9370 ( .A1(n14638), .A2(n11993), .ZN(n9617) );
  NAND2_X1 U9371 ( .A1(n7086), .A2(n14403), .ZN(n7083) );
  AND2_X1 U9372 ( .A1(n7083), .A2(n7082), .ZN(n7422) );
  NAND2_X1 U9373 ( .A1(n6787), .A2(n14761), .ZN(n6934) );
  NAND3_X1 U9374 ( .A1(n7083), .A2(n7082), .A3(n7084), .ZN(n6787) );
  INV_X1 U9375 ( .A(n6788), .ZN(n9585) );
  NAND2_X1 U9376 ( .A1(n6788), .A2(n9586), .ZN(n6894) );
  AND2_X1 U9377 ( .A1(n14724), .A2(n13608), .ZN(n6789) );
  AOI21_X1 U9378 ( .B1(n14741), .B2(n13699), .A(n6790), .ZN(n11358) );
  NOR2_X1 U9379 ( .A1(n6791), .A2(n13752), .ZN(n6790) );
  AOI21_X1 U9380 ( .B1(n14741), .B2(n10426), .A(n11357), .ZN(n11546) );
  AOI21_X1 U9381 ( .B1(n14410), .B2(n10426), .A(n11563), .ZN(n11575) );
  AOI21_X1 U9382 ( .B1(n11897), .B2(n10426), .A(n11576), .ZN(n13602) );
  AOI21_X1 U9383 ( .B1(n14518), .B2(n10426), .A(n13622), .ZN(n13623) );
  AOI21_X1 U9384 ( .B1(n14299), .B2(n10426), .A(n13641), .ZN(n13646) );
  AOI21_X1 U9385 ( .B1(n14288), .B2(n10426), .A(n13659), .ZN(n13660) );
  OR2_X1 U9386 ( .A1(n13740), .A2(n6808), .ZN(n6804) );
  NAND2_X1 U9387 ( .A1(n6804), .A2(n6805), .ZN(n13818) );
  NAND2_X1 U9388 ( .A1(n6813), .A2(n6489), .ZN(n6812) );
  NAND2_X1 U9389 ( .A1(n6814), .A2(n11912), .ZN(n6813) );
  NAND2_X1 U9390 ( .A1(n7587), .A2(n7588), .ZN(n6814) );
  NAND2_X1 U9391 ( .A1(n13837), .A2(n6443), .ZN(n6816) );
  OR2_X1 U9392 ( .A1(n13837), .A2(n13709), .ZN(n6817) );
  NAND2_X1 U9393 ( .A1(n6819), .A2(n12042), .ZN(P1_U3242) );
  NAND2_X1 U9394 ( .A1(n6820), .A2(n6904), .ZN(n6819) );
  NAND4_X1 U9395 ( .A1(n7583), .A2(n6823), .A3(n12038), .A4(n6821), .ZN(n6820)
         );
  NAND2_X1 U9396 ( .A1(n6822), .A2(n6478), .ZN(n6821) );
  INV_X1 U9397 ( .A(n7584), .ZN(n6822) );
  NAND2_X1 U9398 ( .A1(n6824), .A2(n6478), .ZN(n6823) );
  INV_X1 U9399 ( .A(n7585), .ZN(n6824) );
  NAND2_X1 U9400 ( .A1(n11852), .A2(n11851), .ZN(n11856) );
  NAND3_X1 U9401 ( .A1(n11852), .A2(n11851), .A3(n6825), .ZN(n6827) );
  NAND2_X1 U9402 ( .A1(n6826), .A2(n7606), .ZN(n11879) );
  NAND3_X1 U9403 ( .A1(n11858), .A2(n6540), .A3(n6827), .ZN(n6826) );
  MUX2_X1 U9404 ( .A(n11827), .B(n11826), .S(n11903), .Z(n11828) );
  INV_X4 U9405 ( .A(n11815), .ZN(n11903) );
  MUX2_X1 U9406 ( .A(n11981), .B(n6895), .S(n11968), .Z(n11815) );
  OAI21_X1 U9407 ( .B1(n11937), .B2(n6837), .A(n6835), .ZN(n11942) );
  NAND2_X1 U9408 ( .A1(n6834), .A2(n6832), .ZN(n11940) );
  NAND2_X1 U9409 ( .A1(n11937), .A2(n6835), .ZN(n6834) );
  XNOR2_X2 U9410 ( .A(n6841), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U9411 ( .A1(n7708), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U9412 ( .A1(n6845), .A2(n6850), .ZN(n6843) );
  NAND3_X1 U9413 ( .A1(n6846), .A2(n6844), .A3(n6843), .ZN(n6849) );
  INV_X1 U9414 ( .A(n6850), .ZN(n14430) );
  NAND2_X1 U9415 ( .A1(n6849), .A2(n6848), .ZN(P3_U3200) );
  INV_X1 U9416 ( .A(n6855), .ZN(n12410) );
  INV_X1 U9417 ( .A(n14383), .ZN(n6865) );
  NAND3_X1 U9418 ( .A1(n6863), .A2(n6866), .A3(n6860), .ZN(n15323) );
  NAND3_X1 U9419 ( .A1(n6863), .A2(n6861), .A3(n6860), .ZN(n6867) );
  NOR2_X1 U9420 ( .A1(n14383), .A2(n8308), .ZN(n8309) );
  NAND2_X1 U9421 ( .A1(n8308), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6866) );
  INV_X1 U9422 ( .A(n6867), .ZN(n15321) );
  OR2_X1 U9423 ( .A1(n14586), .A2(n6878), .ZN(n6872) );
  NAND3_X1 U9424 ( .A1(n6870), .A2(n6869), .A3(n6868), .ZN(n7223) );
  NAND2_X1 U9425 ( .A1(n6879), .A2(n6871), .ZN(n6869) );
  NAND2_X1 U9426 ( .A1(n6876), .A2(n6871), .ZN(n6870) );
  NAND2_X1 U9427 ( .A1(n6875), .A2(n6872), .ZN(n14363) );
  NAND2_X1 U9428 ( .A1(n14586), .A2(n14588), .ZN(n14427) );
  NAND2_X1 U9429 ( .A1(n6881), .A2(n6551), .ZN(n14575) );
  NAND3_X1 U9430 ( .A1(n7220), .A2(n6913), .A3(n6883), .ZN(n6881) );
  NAND2_X1 U9431 ( .A1(n14589), .A2(n14590), .ZN(n14586) );
  OAI21_X1 U9432 ( .B1(n14575), .B2(n14574), .A(n6965), .ZN(n6885) );
  NAND2_X1 U9433 ( .A1(n14573), .A2(n6885), .ZN(n14578) );
  NAND2_X1 U9434 ( .A1(n10592), .A2(n10593), .ZN(n7211) );
  NAND2_X1 U9435 ( .A1(n12141), .A2(n12284), .ZN(n12178) );
  NAND2_X1 U9436 ( .A1(n11289), .A2(n11288), .ZN(n11290) );
  NAND2_X1 U9437 ( .A1(n12256), .A2(n12147), .ZN(n12316) );
  NAND2_X1 U9438 ( .A1(n11533), .A2(n11532), .ZN(n11535) );
  NAND2_X1 U9439 ( .A1(n10542), .A2(n15068), .ZN(n6886) );
  NAND2_X1 U9440 ( .A1(n11412), .A2(n11411), .ZN(n11533) );
  NAND2_X1 U9442 ( .A1(n7638), .A2(n7637), .ZN(n11937) );
  NAND2_X1 U9443 ( .A1(n7633), .A2(n7635), .ZN(n11964) );
  NAND2_X1 U9444 ( .A1(n13468), .A2(n6946), .ZN(n13556) );
  OAI211_X1 U9445 ( .C1(n14934), .C2(n13470), .A(n13469), .B(n6948), .ZN(n6947) );
  NAND2_X1 U9446 ( .A1(n14363), .A2(n14362), .ZN(n14361) );
  NAND2_X1 U9447 ( .A1(n14581), .A2(n14583), .ZN(n8331) );
  XNOR2_X1 U9448 ( .A(n6891), .B(n7222), .ZN(SUB_1596_U4) );
  NAND2_X1 U9449 ( .A1(n7223), .A2(n14361), .ZN(n6891) );
  NAND2_X1 U9450 ( .A1(n6896), .A2(n6877), .ZN(n6917) );
  NAND2_X1 U9451 ( .A1(n9420), .A2(n9442), .ZN(n9571) );
  NAND2_X1 U9452 ( .A1(n13827), .A2(n13645), .ZN(n13740) );
  NAND2_X1 U9453 ( .A1(n13727), .A2(n13680), .ZN(n13804) );
  NAND2_X1 U9454 ( .A1(n13783), .A2(n13698), .ZN(n13837) );
  INV_X1 U9455 ( .A(n14363), .ZN(n6896) );
  OAI21_X1 U9456 ( .B1(n13464), .B2(n14958), .A(n7046), .ZN(P2_U3496) );
  NAND2_X1 U9457 ( .A1(n14179), .A2(n9627), .ZN(n14161) );
  AOI22_X1 U9458 ( .A1(n13995), .A2(n13994), .B1(n14252), .B2(n13753), .ZN(
        n9630) );
  NOR2_X1 U9459 ( .A1(n10916), .A2(n10915), .ZN(n11126) );
  NAND2_X1 U9460 ( .A1(n11574), .A2(n7357), .ZN(n13607) );
  OAI22_X1 U9461 ( .A1(n11272), .A2(n7373), .B1(n11270), .B2(n11271), .ZN(
        n7372) );
  AOI21_X1 U9462 ( .B1(n12921), .B2(n12920), .A(n13082), .ZN(n12931) );
  NAND2_X1 U9463 ( .A1(n6903), .A2(n6902), .ZN(n14589) );
  NAND2_X1 U9464 ( .A1(n15319), .A2(n15318), .ZN(n15317) );
  XNOR2_X1 U9465 ( .A(n8320), .B(n8321), .ZN(n14397) );
  NAND2_X1 U9466 ( .A1(n11126), .A2(n11125), .ZN(n7373) );
  NAND2_X1 U9467 ( .A1(n14522), .A2(n7359), .ZN(n11574) );
  INV_X1 U9468 ( .A(n7370), .ZN(n7368) );
  NAND2_X1 U9469 ( .A1(n7489), .A2(n7492), .ZN(n8418) );
  NAND2_X1 U9470 ( .A1(n8407), .A2(n8041), .ZN(n7028) );
  OAI21_X1 U9471 ( .B1(n7033), .B2(n7438), .A(n6550), .ZN(n7032) );
  INV_X1 U9472 ( .A(n7032), .ZN(n7031) );
  NAND2_X1 U9473 ( .A1(n10400), .A2(n7311), .ZN(n10399) );
  NAND3_X1 U9474 ( .A1(n7015), .A2(n7016), .A3(n7017), .ZN(n7667) );
  NAND2_X1 U9475 ( .A1(n7668), .A2(n7770), .ZN(n8143) );
  NAND2_X1 U9476 ( .A1(n7199), .A2(n7203), .ZN(n6944) );
  INV_X1 U9477 ( .A(n6939), .ZN(n6920) );
  NAND2_X1 U9478 ( .A1(n7401), .A2(n7402), .ZN(n7839) );
  OAI21_X1 U9479 ( .B1(n10597), .B2(n15068), .A(n11642), .ZN(n10540) );
  INV_X1 U9480 ( .A(n8094), .ZN(n6908) );
  NAND2_X1 U9481 ( .A1(n11789), .A2(n11788), .ZN(n11790) );
  NAND2_X1 U9482 ( .A1(n12930), .A2(n12931), .ZN(n6925) );
  NAND2_X1 U9483 ( .A1(n6437), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6900) );
  INV_X1 U9484 ( .A(n10398), .ZN(n13118) );
  NAND2_X1 U9485 ( .A1(n7242), .A2(n6509), .ZN(n7241) );
  NAND2_X1 U9486 ( .A1(n10959), .A2(n10859), .ZN(n10860) );
  INV_X1 U9487 ( .A(n7366), .ZN(n6942) );
  INV_X1 U9488 ( .A(n8331), .ZN(n6903) );
  OAI21_X1 U9489 ( .B1(n8821), .B2(n8820), .A(n8819), .ZN(n8824) );
  NAND2_X1 U9490 ( .A1(n7626), .A2(n7627), .ZN(n11957) );
  AOI21_X1 U9491 ( .B1(n10544), .B2(n10597), .A(n10543), .ZN(n10545) );
  NAND2_X1 U9492 ( .A1(n7475), .A2(n8741), .ZN(n6929) );
  NAND2_X1 U9493 ( .A1(n11290), .A2(n11406), .ZN(n11409) );
  NAND2_X1 U9494 ( .A1(n12200), .A2(n12199), .ZN(n12198) );
  INV_X1 U9495 ( .A(n12777), .ZN(n7573) );
  AOI21_X1 U9496 ( .B1(n7594), .B2(n7591), .A(n6514), .ZN(n7588) );
  INV_X1 U9497 ( .A(n7599), .ZN(n7598) );
  NAND2_X1 U9498 ( .A1(n14192), .A2(n6568), .ZN(n14179) );
  NAND2_X1 U9499 ( .A1(n6929), .A2(n7478), .ZN(n8762) );
  NAND2_X1 U9500 ( .A1(n8513), .A2(n8349), .ZN(n8516) );
  INV_X1 U9501 ( .A(n7595), .ZN(n7594) );
  NAND2_X1 U9502 ( .A1(n6928), .A2(n6927), .ZN(n11943) );
  NAND2_X1 U9503 ( .A1(n7650), .A2(n11791), .ZN(n7419) );
  NAND4_X1 U9504 ( .A1(n7663), .A2(n7664), .A3(n7666), .A4(n7665), .ZN(n6909)
         );
  NAND3_X1 U9505 ( .A1(n8134), .A2(n7310), .A3(n7671), .ZN(n6911) );
  NAND3_X1 U9506 ( .A1(n7211), .A2(n10596), .A3(n7210), .ZN(n10902) );
  NAND2_X1 U9507 ( .A1(n12316), .A2(n12315), .ZN(n12314) );
  NAND2_X1 U9508 ( .A1(n12258), .A2(n12257), .ZN(n12256) );
  NAND2_X2 U9509 ( .A1(n8152), .A2(n6912), .ZN(n11642) );
  NAND2_X1 U9510 ( .A1(n8325), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U9511 ( .A1(n6917), .A2(n14361), .ZN(n6916) );
  XNOR2_X1 U9512 ( .A(n8248), .B(n8247), .ZN(n8289) );
  INV_X1 U9513 ( .A(n8301), .ZN(n7221) );
  XNOR2_X1 U9514 ( .A(n6916), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9515 ( .A1(n10753), .A2(n10896), .ZN(n11819) );
  NAND2_X1 U9516 ( .A1(n13204), .A2(n13205), .ZN(n12117) );
  NAND2_X1 U9517 ( .A1(n7243), .A2(n7247), .ZN(n13204) );
  NAND2_X1 U9518 ( .A1(n8516), .A2(n8350), .ZN(n8541) );
  INV_X1 U9519 ( .A(n11942), .ZN(n6928) );
  INV_X4 U9520 ( .A(n13754), .ZN(n13699) );
  AOI21_X2 U9521 ( .B1(n6451), .B2(n10913), .A(n10912), .ZN(n11127) );
  NAND2_X1 U9522 ( .A1(n9577), .A2(n7619), .ZN(n6919) );
  AOI21_X1 U9523 ( .B1(n7391), .B2(n7394), .A(n7947), .ZN(n7390) );
  XNOR2_X1 U9524 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7706) );
  NAND2_X1 U9525 ( .A1(n8096), .A2(n8095), .ZN(n8107) );
  NAND2_X1 U9526 ( .A1(n12176), .A2(n12143), .ZN(n12336) );
  NAND2_X1 U9527 ( .A1(n12239), .A2(n7204), .ZN(n7199) );
  NAND2_X1 U9528 ( .A1(n8040), .A2(n6584), .ZN(n8054) );
  XNOR2_X1 U9529 ( .A(n8120), .B(n8109), .ZN(n11490) );
  XNOR2_X1 U9530 ( .A(n6944), .B(n6484), .ZN(n12175) );
  NOR2_X1 U9531 ( .A1(n11127), .A2(n7368), .ZN(n6943) );
  INV_X1 U9532 ( .A(n8441), .ZN(n8433) );
  NAND2_X1 U9533 ( .A1(n8435), .A2(n8434), .ZN(n8440) );
  NAND2_X1 U9534 ( .A1(n6925), .A2(n6571), .ZN(P2_U3186) );
  XNOR2_X1 U9535 ( .A(n8251), .B(n8252), .ZN(n8288) );
  NAND2_X1 U9536 ( .A1(n12905), .A2(n7328), .ZN(n7327) );
  NAND2_X1 U9537 ( .A1(n13035), .A2(n12901), .ZN(n13036) );
  NAND2_X1 U9538 ( .A1(n6934), .A2(n6576), .ZN(P1_U3557) );
  NAND2_X1 U9539 ( .A1(n11975), .A2(n11974), .ZN(n7584) );
  AOI211_X2 U9540 ( .C1(n13462), .C2(n13216), .A(n9733), .B(n13200), .ZN(
        n13461) );
  NAND2_X1 U9541 ( .A1(n7144), .A2(n7143), .ZN(n13410) );
  NAND2_X1 U9542 ( .A1(n7142), .A2(n7141), .ZN(n11386) );
  NAND2_X1 U9543 ( .A1(n7147), .A2(n7146), .ZN(n13304) );
  NAND2_X1 U9544 ( .A1(n13398), .A2(n13382), .ZN(n13376) );
  AND3_X2 U9545 ( .A1(n7462), .A2(n6490), .A3(n8523), .ZN(n10658) );
  NAND2_X1 U9546 ( .A1(n12178), .A2(n12177), .ZN(n12176) );
  NAND2_X1 U9547 ( .A1(n11409), .A2(n11408), .ZN(n11412) );
  NAND2_X1 U9548 ( .A1(n8141), .A2(n8233), .ZN(n8208) );
  NAND2_X1 U9549 ( .A1(n7066), .A2(n6935), .ZN(n7062) );
  NAND2_X1 U9550 ( .A1(n14161), .A2(n14160), .ZN(n14159) );
  NAND2_X1 U9551 ( .A1(n11025), .A2(n7614), .ZN(n11170) );
  NAND2_X1 U9552 ( .A1(n13764), .A2(n10437), .ZN(n10438) );
  CLKBUF_X2 U9553 ( .A(n13873), .Z(n6936) );
  XNOR2_X1 U9554 ( .A(n10431), .B(n6937), .ZN(n10433) );
  NAND2_X1 U9555 ( .A1(n7559), .A2(n8050), .ZN(n6938) );
  NAND2_X1 U9556 ( .A1(n7415), .A2(n6569), .ZN(n7893) );
  INV_X1 U9557 ( .A(n8021), .ZN(n7408) );
  INV_X1 U9558 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7687) );
  INV_X1 U9559 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9560 ( .A1(n13010), .A2(n12877), .ZN(n7315) );
  NAND2_X1 U9561 ( .A1(n8211), .A2(n11219), .ZN(n6941) );
  NAND2_X1 U9562 ( .A1(n7468), .A2(n13226), .ZN(n13225) );
  NAND2_X1 U9563 ( .A1(n6437), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6945) );
  NAND2_X1 U9564 ( .A1(n7036), .A2(n7034), .ZN(n7033) );
  NAND2_X1 U9565 ( .A1(n13766), .A2(n13765), .ZN(n13764) );
  XNOR2_X1 U9566 ( .A(n8299), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15315) );
  XNOR2_X1 U9567 ( .A(n8288), .B(n6949), .ZN(n8299) );
  INV_X1 U9568 ( .A(n8290), .ZN(n7225) );
  NAND2_X1 U9569 ( .A1(n15315), .A2(n15316), .ZN(n15314) );
  NOR2_X1 U9570 ( .A1(n7656), .A2(n14934), .ZN(n7049) );
  NAND2_X1 U9571 ( .A1(n11819), .A2(n11825), .ZN(n11822) );
  NAND2_X1 U9572 ( .A1(n14102), .A2(n14103), .ZN(n14101) );
  NOR2_X1 U9573 ( .A1(n8289), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n8249) );
  XNOR2_X1 U9574 ( .A(n6955), .B(n12322), .ZN(n12333) );
  NAND2_X1 U9575 ( .A1(n6957), .A2(n6956), .ZN(n6955) );
  NAND2_X1 U9576 ( .A1(n12239), .A2(n12240), .ZN(n6957) );
  NAND2_X2 U9577 ( .A1(n9197), .A2(n11592), .ZN(n11802) );
  NAND2_X1 U9578 ( .A1(n11495), .A2(n9624), .ZN(n7625) );
  NAND2_X1 U9579 ( .A1(n14101), .A2(n9628), .ZN(n14078) );
  NAND2_X1 U9580 ( .A1(n7062), .A2(n7648), .ZN(n13995) );
  INV_X1 U9581 ( .A(n10679), .ZN(n7318) );
  NAND2_X1 U9582 ( .A1(n11976), .A2(n11977), .ZN(n7585) );
  NAND2_X1 U9583 ( .A1(n6436), .A2(n13116), .ZN(n8505) );
  NAND3_X1 U9584 ( .A1(n6436), .A2(n14867), .A3(n13118), .ZN(n8502) );
  OAI21_X1 U9585 ( .B1(n8740), .B2(n7535), .A(n6967), .ZN(n6966) );
  AOI21_X1 U9586 ( .B1(n8740), .B2(n7532), .A(n7530), .ZN(n6970) );
  NAND2_X1 U9587 ( .A1(n9051), .A2(n6972), .ZN(n6971) );
  NOR2_X1 U9588 ( .A1(n9085), .A2(n9089), .ZN(n6978) );
  INV_X1 U9589 ( .A(n9032), .ZN(n6979) );
  NAND2_X1 U9590 ( .A1(n6983), .A2(n6980), .ZN(n8652) );
  NAND3_X1 U9591 ( .A1(n6982), .A2(n6981), .A3(n6987), .ZN(n6980) );
  NAND2_X1 U9592 ( .A1(n8611), .A2(n8610), .ZN(n6981) );
  NAND2_X1 U9593 ( .A1(n8608), .A2(n8607), .ZN(n6982) );
  NAND3_X1 U9594 ( .A1(n6985), .A2(n6984), .A3(n6988), .ZN(n6983) );
  NAND2_X1 U9595 ( .A1(n8611), .A2(n6535), .ZN(n6984) );
  NAND2_X1 U9596 ( .A1(n8608), .A2(n6986), .ZN(n6985) );
  OAI22_X1 U9597 ( .A1(n8695), .A2(n6989), .B1(n8694), .B2(n6991), .ZN(n8714)
         );
  NOR2_X1 U9598 ( .A1(n8714), .A2(n8713), .ZN(n8715) );
  INV_X1 U9599 ( .A(n8693), .ZN(n6991) );
  NAND3_X1 U9600 ( .A1(n8876), .A2(n8875), .A3(n6572), .ZN(n6992) );
  OAI211_X1 U9601 ( .C1(n8572), .C2(n6995), .A(n6552), .B(n6994), .ZN(n6993)
         );
  NAND2_X1 U9602 ( .A1(n6993), .A2(n7539), .ZN(n8609) );
  NOR2_X1 U9603 ( .A1(n8997), .A2(n8996), .ZN(n6996) );
  AOI21_X1 U9604 ( .B1(n8997), .B2(n8996), .A(n8995), .ZN(n6997) );
  NAND2_X1 U9605 ( .A1(n7007), .A2(n7008), .ZN(n7843) );
  NAND2_X1 U9606 ( .A1(n11089), .A2(n7009), .ZN(n7007) );
  NAND2_X1 U9607 ( .A1(n13238), .A2(n12082), .ZN(n7468) );
  OAI21_X1 U9608 ( .B1(n13238), .B2(n7250), .A(n7021), .ZN(n13206) );
  NAND3_X1 U9609 ( .A1(n7020), .A2(n12084), .A3(n7019), .ZN(n12085) );
  NAND2_X1 U9610 ( .A1(n13238), .A2(n7021), .ZN(n7020) );
  NAND3_X1 U9611 ( .A1(n7482), .A2(n7483), .A3(n7484), .ZN(n8858) );
  NAND3_X1 U9612 ( .A1(n8937), .A2(n7027), .A3(n9100), .ZN(n8939) );
  NAND2_X1 U9613 ( .A1(n7028), .A2(n8410), .ZN(n9480) );
  OR2_X1 U9614 ( .A1(n7437), .A2(n7033), .ZN(n7030) );
  NAND2_X1 U9615 ( .A1(n7030), .A2(n7031), .ZN(n13256) );
  INV_X1 U9616 ( .A(n13279), .ZN(n7034) );
  NAND2_X1 U9617 ( .A1(n7437), .A2(n7438), .ZN(n7035) );
  NAND2_X1 U9618 ( .A1(n13440), .A2(n7038), .ZN(n7037) );
  NAND2_X1 U9619 ( .A1(n7037), .A2(n7039), .ZN(n13394) );
  XNOR2_X1 U9620 ( .A(n12085), .B(n12118), .ZN(n7047) );
  AOI21_X2 U9621 ( .B1(n7047), .B2(n14882), .A(n12088), .ZN(n13464) );
  NAND2_X1 U9622 ( .A1(n7461), .A2(n7051), .ZN(n7050) );
  NAND2_X1 U9623 ( .A1(n7050), .A2(n6547), .ZN(n12077) );
  NAND3_X1 U9624 ( .A1(n7066), .A2(n7065), .A3(n7064), .ZN(n14012) );
  NAND2_X1 U9625 ( .A1(n14046), .A2(n14045), .ZN(n14044) );
  INV_X1 U9626 ( .A(n14027), .ZN(n14032) );
  INV_X1 U9627 ( .A(n7072), .ZN(n7514) );
  NAND2_X1 U9628 ( .A1(n7072), .A2(n8402), .ZN(n8894) );
  XNOR2_X1 U9629 ( .A(n9630), .B(n12015), .ZN(n7086) );
  NAND2_X1 U9630 ( .A1(n7087), .A2(n7088), .ZN(n8370) );
  NAND2_X1 U9631 ( .A1(n8366), .A2(n7089), .ZN(n7087) );
  NAND2_X1 U9632 ( .A1(n14052), .A2(n14051), .ZN(n14050) );
  NAND2_X1 U9633 ( .A1(n9228), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9567) );
  AOI21_X1 U9634 ( .B1(n9417), .B2(n7097), .A(n7095), .ZN(n7094) );
  INV_X1 U9635 ( .A(n7094), .ZN(n9458) );
  NAND2_X1 U9636 ( .A1(n7109), .A2(n7107), .ZN(n9283) );
  NAND3_X1 U9637 ( .A1(n6459), .A2(n9264), .A3(n10733), .ZN(n7109) );
  NAND2_X1 U9638 ( .A1(n11347), .A2(n6453), .ZN(n7116) );
  NAND2_X1 U9639 ( .A1(n14033), .A2(n7138), .ZN(n7137) );
  NOR2_X2 U9640 ( .A1(n11115), .A2(n11232), .ZN(n7142) );
  NOR2_X2 U9641 ( .A1(n13410), .A2(n13533), .ZN(n13398) );
  NOR2_X1 U9642 ( .A1(n13243), .A2(n7152), .ZN(n13200) );
  NOR2_X1 U9643 ( .A1(n13243), .A2(n13472), .ZN(n13230) );
  OR3_X1 U9644 ( .A1(n13243), .A2(n13465), .A3(n13472), .ZN(n13216) );
  NAND2_X1 U9645 ( .A1(n14448), .A2(n7162), .ZN(n7161) );
  INV_X1 U9646 ( .A(n7173), .ZN(n10485) );
  INV_X1 U9647 ( .A(n7172), .ZN(n10576) );
  NAND2_X1 U9648 ( .A1(n10480), .A2(n10481), .ZN(n7174) );
  INV_X2 U9649 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7176) );
  OR2_X1 U9650 ( .A1(n11978), .A2(n8347), .ZN(n7178) );
  NAND3_X1 U9651 ( .A1(n6467), .A2(n14006), .A3(n14055), .ZN(n13985) );
  INV_X1 U9652 ( .A(n7182), .ZN(n14018) );
  NAND2_X1 U9653 ( .A1(n6549), .A2(n14209), .ZN(n14165) );
  NOR2_X1 U9654 ( .A1(n14741), .A2(n7189), .ZN(n7188) );
  NAND2_X1 U9655 ( .A1(n12239), .A2(n6534), .ZN(n7192) );
  OAI211_X1 U9656 ( .C1(n12239), .C2(n7197), .A(n7192), .B(n7193), .ZN(n12215)
         );
  AND2_X1 U9657 ( .A1(n12169), .A2(n12519), .ZN(n7207) );
  NAND2_X1 U9658 ( .A1(n7209), .A2(n6543), .ZN(n11289) );
  NAND2_X1 U9659 ( .A1(n7770), .A2(n7216), .ZN(n7902) );
  NAND2_X1 U9660 ( .A1(n7218), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7877) );
  NOR2_X2 U9661 ( .A1(n8721), .A2(n7227), .ZN(n8781) );
  NAND4_X1 U9662 ( .A1(n7231), .A2(n7230), .A3(n7229), .A4(n7228), .ZN(n7227)
         );
  INV_X1 U9663 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7231) );
  NAND3_X1 U9664 ( .A1(n7234), .A2(n7233), .A3(n7232), .ZN(n8721) );
  NAND2_X4 U9665 ( .A1(n7235), .A2(n8465), .ZN(n8986) );
  NAND2_X1 U9666 ( .A1(n7235), .A2(n8467), .ZN(n8537) );
  NAND2_X1 U9667 ( .A1(n10817), .A2(n10812), .ZN(n7236) );
  NAND3_X1 U9668 ( .A1(n7237), .A2(n10813), .A3(n7236), .ZN(n10815) );
  NAND3_X1 U9669 ( .A1(n10660), .A2(n10812), .A3(n10659), .ZN(n7237) );
  NAND2_X1 U9670 ( .A1(n7238), .A2(n10812), .ZN(n10835) );
  NAND2_X1 U9671 ( .A1(n10811), .A2(n10810), .ZN(n7238) );
  INV_X1 U9672 ( .A(n10857), .ZN(n7242) );
  NAND2_X1 U9673 ( .A1(n13254), .A2(n7244), .ZN(n7243) );
  AND2_X1 U9674 ( .A1(n10946), .A2(n11110), .ZN(n7265) );
  NAND2_X1 U9675 ( .A1(n8425), .A2(n7267), .ZN(n7266) );
  NAND2_X1 U9676 ( .A1(n8425), .A2(n8424), .ZN(n9154) );
  NAND3_X1 U9677 ( .A1(n7275), .A2(n7274), .A3(n7005), .ZN(n12686) );
  NAND2_X1 U9678 ( .A1(n9669), .A2(n15072), .ZN(n7277) );
  NAND2_X1 U9679 ( .A1(n8169), .A2(n7288), .ZN(n7287) );
  OAI21_X1 U9680 ( .B1(n12614), .B2(n7295), .A(n7293), .ZN(n8178) );
  OAI21_X1 U9681 ( .B1(n12474), .B2(n7298), .A(n7297), .ZN(n9658) );
  NAND2_X1 U9682 ( .A1(n12474), .A2(n11745), .ZN(n7301) );
  NAND2_X1 U9683 ( .A1(n10860), .A2(n10865), .ZN(n10937) );
  NAND2_X1 U9684 ( .A1(n12111), .A2(n12110), .ZN(n13278) );
  NAND2_X1 U9685 ( .A1(n12686), .A2(n8173), .ZN(n12672) );
  NAND2_X1 U9686 ( .A1(n12587), .A2(n8179), .ZN(n12573) );
  OAI21_X2 U9687 ( .B1(n12488), .B2(n8189), .A(n8188), .ZN(n12474) );
  NAND2_X1 U9688 ( .A1(n11644), .A2(n11645), .ZN(n15041) );
  NAND2_X1 U9689 ( .A1(n12573), .A2(n12572), .ZN(n12571) );
  NAND2_X1 U9690 ( .A1(n12588), .A2(n7644), .ZN(n12587) );
  NAND4_X2 U9691 ( .A1(n7769), .A2(n7768), .A3(n7767), .A4(n7766), .ZN(n15029)
         );
  NOR2_X2 U9692 ( .A1(n10673), .A2(n10819), .ZN(n10842) );
  NAND2_X1 U9693 ( .A1(n11092), .A2(n8167), .ZN(n11221) );
  NAND2_X1 U9694 ( .A1(n8193), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7683) );
  INV_X1 U9695 ( .A(n11221), .ZN(n8169) );
  NAND2_X1 U9696 ( .A1(n8187), .A2(n8186), .ZN(n12488) );
  OR2_X1 U9697 ( .A1(n9025), .A2(n8477), .ZN(n8482) );
  XNOR2_X2 U9698 ( .A(n13116), .B(n10297), .ZN(n10296) );
  OAI21_X1 U9699 ( .B1(n10400), .B2(n7311), .A(n10399), .ZN(n10401) );
  XNOR2_X1 U9700 ( .A(n9701), .B(n9702), .ZN(n7311) );
  NOR2_X1 U9701 ( .A1(n12906), .A2(n12907), .ZN(n7333) );
  NAND2_X1 U9702 ( .A1(n12921), .A2(n6536), .ZN(n7335) );
  OAI211_X1 U9703 ( .C1(n12921), .C2(n7336), .A(n7335), .B(n12973), .ZN(
        P2_U3192) );
  NAND3_X1 U9704 ( .A1(n9693), .A2(n8474), .A3(n13188), .ZN(n7349) );
  NAND4_X1 U9705 ( .A1(n8781), .A2(n8564), .A3(n7352), .A4(n8420), .ZN(n8441)
         );
  NAND4_X1 U9706 ( .A1(n8781), .A2(n8564), .A3(n8420), .A4(n7353), .ZN(n7351)
         );
  OAI21_X1 U9707 ( .B1(n13617), .B2(n7383), .A(n7380), .ZN(n7385) );
  INV_X1 U9708 ( .A(n7385), .ZN(n14512) );
  NAND2_X1 U9709 ( .A1(n7690), .A2(n7706), .ZN(n7387) );
  NAND2_X1 U9710 ( .A1(n7388), .A2(n7390), .ZN(n7950) );
  NAND2_X1 U9711 ( .A1(n7916), .A2(n7391), .ZN(n7388) );
  NOR2_X1 U9712 ( .A1(n11755), .A2(n7395), .ZN(n11752) );
  NAND2_X1 U9713 ( .A1(n12476), .A2(n7397), .ZN(n7396) );
  NAND3_X1 U9714 ( .A1(n11744), .A2(n11743), .A3(n7399), .ZN(n7398) );
  NOR2_X1 U9715 ( .A1(n7408), .A2(n8024), .ZN(n7407) );
  NAND2_X1 U9716 ( .A1(n7857), .A2(n7416), .ZN(n7415) );
  INV_X1 U9717 ( .A(n9212), .ZN(n10751) );
  NOR2_X1 U9718 ( .A1(n14083), .A2(n7654), .ZN(n14066) );
  AND2_X1 U9719 ( .A1(n9420), .A2(n7434), .ZN(n9205) );
  NOR2_X1 U9720 ( .A1(n9189), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U9721 ( .A1(n9420), .A2(n6542), .ZN(n9202) );
  INV_X1 U9722 ( .A(n9189), .ZN(n7436) );
  INV_X1 U9723 ( .A(n13297), .ZN(n7437) );
  INV_X1 U9724 ( .A(n10967), .ZN(n7447) );
  INV_X1 U9725 ( .A(n10863), .ZN(n7449) );
  NAND2_X1 U9726 ( .A1(n7440), .A2(n7444), .ZN(n10943) );
  NAND2_X1 U9727 ( .A1(n10863), .A2(n7446), .ZN(n7440) );
  NAND2_X1 U9728 ( .A1(n7442), .A2(n7444), .ZN(n7441) );
  NAND2_X1 U9729 ( .A1(n7444), .A2(n14856), .ZN(n7443) );
  AOI21_X2 U9730 ( .B1(n10862), .B2(n7446), .A(n6457), .ZN(n7444) );
  INV_X1 U9731 ( .A(n10862), .ZN(n7450) );
  XNOR2_X2 U9732 ( .A(n10658), .B(n13115), .ZN(n10661) );
  OR2_X1 U9733 ( .A1(n6442), .A2(n9824), .ZN(n7462) );
  NAND2_X1 U9734 ( .A1(n8425), .A2(n7463), .ZN(n9152) );
  AOI21_X2 U9735 ( .B1(n7466), .B2(n14882), .A(n7464), .ZN(n13474) );
  NAND3_X1 U9736 ( .A1(n9086), .A2(n7471), .A3(n7470), .ZN(n7469) );
  OAI21_X1 U9737 ( .B1(n9125), .B2(n9122), .A(n7474), .ZN(n7473) );
  NAND2_X1 U9738 ( .A1(n8980), .A2(n8414), .ZN(n8999) );
  NAND2_X1 U9739 ( .A1(n9035), .A2(n9034), .ZN(n7513) );
  NAND2_X1 U9740 ( .A1(n9035), .A2(n7505), .ZN(n7504) );
  NAND2_X1 U9741 ( .A1(n7513), .A2(n9037), .ZN(n9066) );
  OAI21_X1 U9742 ( .B1(n8911), .B2(n7522), .A(n7519), .ZN(n8930) );
  INV_X1 U9743 ( .A(n7516), .ZN(n8929) );
  AOI21_X1 U9744 ( .B1(n8911), .B2(n7519), .A(n7517), .ZN(n7516) );
  NAND2_X1 U9745 ( .A1(n7518), .A2(n8931), .ZN(n7517) );
  NAND2_X1 U9746 ( .A1(n7522), .A2(n7519), .ZN(n7518) );
  OAI21_X1 U9747 ( .B1(n8952), .B2(n7529), .A(n7526), .ZN(n8972) );
  INV_X1 U9748 ( .A(n7523), .ZN(n8971) );
  NAND3_X1 U9749 ( .A1(n8657), .A2(n6553), .A3(n8656), .ZN(n7536) );
  NAND2_X1 U9750 ( .A1(n7536), .A2(n7537), .ZN(n8695) );
  INV_X1 U9751 ( .A(n8609), .ZN(n8611) );
  INV_X1 U9752 ( .A(n7541), .ZN(n7544) );
  AOI22_X1 U9753 ( .A1(n7545), .A2(n9016), .B1(n7547), .B2(n7551), .ZN(n7542)
         );
  INV_X1 U9754 ( .A(n9017), .ZN(n7548) );
  INV_X1 U9755 ( .A(n9154), .ZN(n7553) );
  NAND2_X1 U9756 ( .A1(n7553), .A2(n7554), .ZN(n13573) );
  MUX2_X1 U9757 ( .A(n9685), .B(n7557), .S(n15149), .Z(n9687) );
  NAND2_X1 U9758 ( .A1(n12777), .A2(n11642), .ZN(n7570) );
  OR2_X2 U9759 ( .A1(n12772), .A2(n15063), .ZN(n11630) );
  NAND4_X1 U9760 ( .A1(n7570), .A2(n7571), .A3(n11630), .A4(n11633), .ZN(n7712) );
  NAND2_X1 U9761 ( .A1(n10544), .A2(n11642), .ZN(n15062) );
  NAND2_X1 U9762 ( .A1(n7573), .A2(n11632), .ZN(n10544) );
  NAND3_X1 U9763 ( .A1(n7661), .A2(n7577), .A3(n7662), .ZN(n7574) );
  NAND3_X1 U9764 ( .A1(n7585), .A2(n7584), .A3(n12037), .ZN(n7583) );
  NAND3_X1 U9765 ( .A1(n11892), .A2(n11891), .A3(n7586), .ZN(n7587) );
  NAND3_X1 U9766 ( .A1(n11881), .A2(n11880), .A3(n6570), .ZN(n7611) );
  NAND2_X1 U9767 ( .A1(n7611), .A2(n7612), .ZN(n11887) );
  INV_X1 U9768 ( .A(n11884), .ZN(n7613) );
  NAND2_X1 U9769 ( .A1(n11845), .A2(n11846), .ZN(n7617) );
  NAND3_X1 U9770 ( .A1(n11838), .A2(n11837), .A3(n11987), .ZN(n7618) );
  NAND2_X1 U9771 ( .A1(n9577), .A2(n7620), .ZN(n14339) );
  NAND2_X1 U9772 ( .A1(n10801), .A2(n14613), .ZN(n9618) );
  NAND2_X1 U9773 ( .A1(n11951), .A2(n11948), .ZN(n7629) );
  NAND2_X1 U9774 ( .A1(n11949), .A2(n7629), .ZN(n7626) );
  NAND2_X4 U9775 ( .A1(n9196), .A2(n9195), .ZN(n9254) );
  OAI22_X1 U9776 ( .A1(n9196), .A2(P1_U3086), .B1(n11807), .B2(n14353), .ZN(
        n7631) );
  NAND2_X1 U9777 ( .A1(n11961), .A2(n7632), .ZN(n7634) );
  INV_X1 U9778 ( .A(n11960), .ZN(n7632) );
  NAND3_X1 U9779 ( .A1(n11959), .A2(n7634), .A3(n11958), .ZN(n7633) );
  NAND3_X1 U9780 ( .A1(n11933), .A2(n11932), .A3(n7636), .ZN(n7638) );
  INV_X1 U9781 ( .A(n11934), .ZN(n7639) );
  INV_X1 U9782 ( .A(n14465), .ZN(n8172) );
  NAND2_X1 U9783 ( .A1(n14257), .A2(n14256), .ZN(n14323) );
  NAND2_X1 U9784 ( .A1(n9213), .A2(n9212), .ZN(n11825) );
  NAND4_X4 U9785 ( .A1(n8482), .A2(n8481), .A3(n8480), .A4(n8479), .ZN(n13116)
         );
  INV_X1 U9786 ( .A(n11819), .ZN(n11820) );
  NOR2_X1 U9787 ( .A1(n11593), .A2(n11753), .ZN(n11626) );
  OAI21_X1 U9788 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(n9174) );
  OR2_X1 U9789 ( .A1(n9171), .A2(n9124), .ZN(n9165) );
  OR2_X1 U9790 ( .A1(n11850), .A2(n11849), .ZN(n11851) );
  NAND2_X1 U9791 ( .A1(n15054), .A2(n11644), .ZN(n11015) );
  INV_X1 U9792 ( .A(n11995), .ZN(n10799) );
  OR2_X1 U9793 ( .A1(n12210), .A2(n15046), .ZN(n7643) );
  NAND2_X1 U9794 ( .A1(n11718), .A2(n11719), .ZN(n7644) );
  OR3_X1 U9795 ( .A1(n12053), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n7646) );
  AND2_X1 U9796 ( .A1(n8200), .A2(n7643), .ZN(n7647) );
  OR2_X1 U9797 ( .A1(n12048), .A2(n12769), .ZN(n7649) );
  XOR2_X1 U9798 ( .A(n11627), .B(n12459), .Z(n7650) );
  INV_X1 U9799 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U9800 ( .A1(n9079), .A2(n9078), .ZN(n13227) );
  INV_X1 U9801 ( .A(n13227), .ZN(n12926) );
  INV_X1 U9802 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n8347) );
  INV_X1 U9803 ( .A(SI_24_), .ZN(n15242) );
  AND2_X1 U9804 ( .A1(n8394), .A2(n8393), .ZN(n7651) );
  OR2_X1 U9805 ( .A1(n15310), .A2(n13867), .ZN(n7652) );
  OR2_X1 U9806 ( .A1(n12048), .A2(n12846), .ZN(n7653) );
  AND2_X1 U9807 ( .A1(n14089), .A2(n13861), .ZN(n7654) );
  INV_X1 U9808 ( .A(n13444), .ZN(n13422) );
  NAND2_X2 U9809 ( .A1(n10502), .A2(n15083), .ZN(n15091) );
  NOR2_X1 U9810 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n7655) );
  INV_X1 U9811 ( .A(n10426), .ZN(n10430) );
  INV_X1 U9812 ( .A(n12011), .ZN(n9548) );
  AND2_X1 U9813 ( .A1(n9059), .A2(n9096), .ZN(n7657) );
  AND2_X1 U9814 ( .A1(n8851), .A2(n8841), .ZN(n7658) );
  INV_X1 U9815 ( .A(n12302), .ZN(n14473) );
  OR2_X1 U9816 ( .A1(n9168), .A2(n13188), .ZN(n7659) );
  NAND2_X2 U9817 ( .A1(n10654), .A2(n14881), .ZN(n13402) );
  AOI21_X1 U9818 ( .B1(n13115), .B2(n8728), .A(n6539), .ZN(n8532) );
  INV_X1 U9819 ( .A(n8868), .ZN(n8869) );
  INV_X1 U9820 ( .A(n8931), .ZN(n8932) );
  OR4_X1 U9821 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n8223) );
  INV_X1 U9822 ( .A(n8073), .ZN(n8072) );
  INV_X1 U9823 ( .A(n11990), .ZN(n9612) );
  INV_X1 U9824 ( .A(n13873), .ZN(n9213) );
  NOR2_X1 U9825 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9344) );
  INV_X1 U9826 ( .A(n8031), .ZN(n8030) );
  INV_X1 U9827 ( .A(n7963), .ZN(n7962) );
  NAND2_X1 U9828 ( .A1(n8083), .A2(n8082), .ZN(n8099) );
  INV_X1 U9829 ( .A(n11719), .ZN(n8007) );
  INV_X1 U9830 ( .A(n7866), .ZN(n7865) );
  OR2_X1 U9831 ( .A1(n12359), .A2(n15035), .ZN(n11653) );
  INV_X1 U9832 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7669) );
  INV_X1 U9833 ( .A(n9005), .ZN(n8458) );
  INV_X1 U9834 ( .A(n8665), .ZN(n8453) );
  AND2_X1 U9835 ( .A1(n13207), .A2(n13208), .ZN(n12083) );
  INV_X1 U9836 ( .A(n8883), .ZN(n8455) );
  INV_X1 U9837 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8683) );
  INV_X1 U9838 ( .A(n8721), .ZN(n8722) );
  INV_X1 U9839 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15248) );
  INV_X1 U9840 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n15198) );
  AND2_X1 U9841 ( .A1(n10457), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10144) );
  AND2_X1 U9842 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n9483), .ZN(n9494) );
  INV_X1 U9843 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9299) );
  AND2_X1 U9844 ( .A1(n9250), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9273) );
  INV_X1 U9845 ( .A(n14274), .ZN(n9634) );
  INV_X1 U9846 ( .A(SI_11_), .ZN(n8371) );
  NAND2_X1 U9847 ( .A1(n6437), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8346) );
  INV_X1 U9848 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U9849 ( .A1(n8030), .A2(n15248), .ZN(n8044) );
  INV_X1 U9850 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U9851 ( .A1(n7962), .A2(n7961), .ZN(n7979) );
  NAND2_X1 U9852 ( .A1(n7865), .A2(n7864), .ZN(n7884) );
  OR2_X1 U9853 ( .A1(n12357), .A2(n11410), .ZN(n11668) );
  INV_X1 U9854 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7955) );
  OR3_X1 U9855 ( .A1(n9070), .A2(n12922), .A3(n12969), .ZN(n9071) );
  NAND2_X1 U9856 ( .A1(n8458), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U9857 ( .A1(n8457), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8984) );
  OR2_X1 U9858 ( .A1(n8899), .A2(n13024), .ZN(n8918) );
  OR2_X1 U9859 ( .A1(n14923), .A2(n8449), .ZN(n10307) );
  INV_X1 U9860 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9327) );
  INV_X1 U9861 ( .A(n9482), .ZN(n9483) );
  AND2_X1 U9862 ( .A1(n9273), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9287) );
  NOR2_X1 U9863 ( .A1(n14299), .A2(n14165), .ZN(n14149) );
  INV_X1 U9864 ( .A(n14209), .ZN(n14226) );
  INV_X1 U9865 ( .A(n11981), .ZN(n12018) );
  AND2_X1 U9866 ( .A1(n8383), .A2(n8382), .ZN(n8741) );
  NAND2_X1 U9867 ( .A1(n7814), .A2(n11537), .ZN(n7827) );
  OR2_X1 U9868 ( .A1(n8044), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U9869 ( .A1(n10545), .A2(n10548), .ZN(n10586) );
  NAND2_X1 U9870 ( .A1(n10550), .A2(n15069), .ZN(n12340) );
  INV_X1 U9871 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11537) );
  INV_X1 U9872 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11074) );
  OR2_X1 U9873 ( .A1(n8129), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12046) );
  INV_X1 U9874 ( .A(n9667), .ZN(n9668) );
  AND2_X1 U9875 ( .A1(n11740), .A2(n11739), .ZN(n12491) );
  AND2_X1 U9876 ( .A1(n10498), .A2(n10497), .ZN(n10499) );
  OR2_X1 U9877 ( .A1(n6441), .A2(n11491), .ZN(n8110) );
  OR2_X1 U9878 ( .A1(n6441), .A2(n8041), .ZN(n8042) );
  INV_X1 U9879 ( .A(SI_15_), .ZN(n8384) );
  AND3_X1 U9880 ( .A1(n7881), .A2(n7880), .A3(n7879), .ZN(n14479) );
  INV_X1 U9881 ( .A(n11007), .ZN(n15035) );
  INV_X1 U9882 ( .A(n11018), .ZN(n11759) );
  INV_X1 U9883 ( .A(n15072), .ZN(n15043) );
  INV_X1 U9884 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U9885 ( .A1(n7841), .A2(n7840), .ZN(n7855) );
  INV_X1 U9886 ( .A(n12927), .ZN(n12928) );
  AND2_X1 U9887 ( .A1(n9005), .A2(n9004), .ZN(n13264) );
  INV_X1 U9888 ( .A(n8986), .ZN(n9043) );
  AND2_X1 U9889 ( .A1(n10413), .A2(n10412), .ZN(n10417) );
  AND2_X1 U9890 ( .A1(n9804), .A2(n9803), .ZN(n9812) );
  INV_X1 U9891 ( .A(n13159), .ZN(n13166) );
  NAND2_X1 U9892 ( .A1(n13097), .A2(n13195), .ZN(n12087) );
  INV_X1 U9893 ( .A(n11155), .ZN(n11153) );
  NAND2_X1 U9894 ( .A1(n13402), .A2(n10671), .ZN(n14874) );
  INV_X1 U9895 ( .A(n14882), .ZN(n13424) );
  NAND2_X1 U9896 ( .A1(n9693), .A2(n14880), .ZN(n14923) );
  INV_X1 U9897 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8432) );
  OR2_X1 U9898 ( .A1(n8724), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8746) );
  OR2_X1 U9899 ( .A1(n9452), .A2(n9451), .ZN(n9461) );
  INV_X1 U9900 ( .A(n14195), .ZN(n14511) );
  INV_X1 U9901 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15228) );
  OR2_X1 U9902 ( .A1(n10233), .A2(n10232), .ZN(n10250) );
  INV_X1 U9903 ( .A(n11320), .ZN(n11322) );
  NOR2_X1 U9904 ( .A1(n9636), .A2(n12018), .ZN(n10143) );
  NAND2_X1 U9905 ( .A1(n14030), .A2(n14619), .ZN(n13997) );
  INV_X1 U9906 ( .A(n12009), .ZN(n14065) );
  INV_X1 U9907 ( .A(n14283), .ZN(n14100) );
  AOI21_X1 U9908 ( .B1(n9307), .B2(n7652), .A(n9306), .ZN(n11031) );
  AND2_X1 U9909 ( .A1(n11868), .A2(n11864), .ZN(n14615) );
  INV_X1 U9910 ( .A(n14708), .ZN(n10704) );
  OR2_X1 U9911 ( .A1(n14656), .A2(n10151), .ZN(n14190) );
  NAND2_X1 U9912 ( .A1(n9591), .A2(n9593), .ZN(n9877) );
  NOR2_X1 U9913 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n8287), .ZN(n8254) );
  INV_X1 U9914 ( .A(n12340), .ZN(n12323) );
  INV_X1 U9915 ( .A(n12327), .ZN(n12344) );
  AOI21_X1 U9916 ( .B1(n12468), .B2(n8193), .A(n8133), .ZN(n12478) );
  AND4_X1 U9917 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), .ZN(n12574)
         );
  INV_X1 U9918 ( .A(n14989), .ZN(n15017) );
  INV_X1 U9919 ( .A(n14976), .ZN(n15007) );
  AND3_X1 U9920 ( .A1(n6432), .A2(n10190), .A3(n11748), .ZN(n15069) );
  NAND2_X1 U9921 ( .A1(n8150), .A2(n8149), .ZN(n15031) );
  NOR2_X1 U9922 ( .A1(n10502), .A2(n15084), .ZN(n15058) );
  AND2_X1 U9923 ( .A1(n10351), .A2(n15084), .ZN(n15053) );
  INV_X1 U9924 ( .A(n15111), .ZN(n14477) );
  NAND2_X1 U9925 ( .A1(n8151), .A2(n10515), .ZN(n15111) );
  OR2_X1 U9926 ( .A1(n15031), .A2(n15132), .ZN(n15102) );
  INV_X1 U9927 ( .A(n15046), .ZN(n15066) );
  NAND2_X1 U9928 ( .A1(n8217), .A2(n8216), .ZN(n10496) );
  INV_X1 U9929 ( .A(n13091), .ZN(n13070) );
  INV_X1 U9930 ( .A(n12996), .ZN(n13089) );
  NAND2_X1 U9931 ( .A1(n10365), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13091) );
  INV_X1 U9932 ( .A(n13039), .ZN(n13078) );
  NAND2_X1 U9933 ( .A1(n9171), .A2(n7659), .ZN(n9169) );
  OR2_X1 U9934 ( .A1(n13069), .A2(n8986), .ZN(n8473) );
  INV_X1 U9935 ( .A(n14794), .ZN(n14840) );
  INV_X1 U9936 ( .A(n14844), .ZN(n14816) );
  AND2_X1 U9937 ( .A1(n9158), .A2(n9790), .ZN(n13444) );
  INV_X1 U9938 ( .A(n14868), .ZN(n14850) );
  AND2_X1 U9939 ( .A1(n14895), .A2(n9782), .ZN(n14865) );
  AND3_X1 U9940 ( .A1(n13501), .A2(n13500), .A3(n13499), .ZN(n13502) );
  AND2_X1 U9941 ( .A1(n14922), .A2(n14923), .ZN(n14934) );
  AND2_X1 U9942 ( .A1(n10653), .A2(n10308), .ZN(n10874) );
  OR3_X1 U9943 ( .A1(n13591), .A2(n13583), .A3(n13585), .ZN(n9799) );
  AND2_X1 U9944 ( .A1(n9833), .A2(P2_U3088), .ZN(n13577) );
  NOR2_X1 U9945 ( .A1(n11281), .A2(n14127), .ZN(n14526) );
  INV_X1 U9946 ( .A(n11281), .ZN(n15299) );
  INV_X1 U9947 ( .A(n15306), .ZN(n14532) );
  AND4_X1 U9948 ( .A1(n9399), .A2(n9398), .A3(n9397), .A4(n9396), .ZN(n14508)
         );
  INV_X1 U9949 ( .A(n14604), .ZN(n13976) );
  INV_X1 U9950 ( .A(n13926), .ZN(n14607) );
  INV_X1 U9951 ( .A(n11525), .ZN(n14230) );
  AND2_X1 U9952 ( .A1(n10149), .A2(n13877), .ZN(n14619) );
  INV_X1 U9953 ( .A(n14202), .ZN(n14634) );
  NAND2_X1 U9954 ( .A1(n9595), .A2(n9879), .ZN(n10171) );
  AND2_X1 U9955 ( .A1(n10756), .A2(n14729), .ZN(n14703) );
  INV_X1 U9956 ( .A(n14703), .ZN(n14748) );
  OR2_X1 U9957 ( .A1(n9882), .A2(n10457), .ZN(n10155) );
  INV_X1 U9958 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9193) );
  AND2_X1 U9959 ( .A1(n9406), .A2(n9418), .ZN(n10982) );
  INV_X1 U9960 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9224) );
  AND2_X1 U9961 ( .A1(n6439), .A2(P1_U3086), .ZN(n14341) );
  AND2_X1 U9962 ( .A1(n10186), .A2(n10185), .ZN(n14995) );
  AND2_X1 U9963 ( .A1(n10350), .A2(n10349), .ZN(n12339) );
  INV_X1 U9964 ( .A(n12519), .ZN(n12489) );
  INV_X1 U9965 ( .A(n12618), .ZN(n12589) );
  INV_X1 U9966 ( .A(n14995), .ZN(n15024) );
  OR2_X1 U9967 ( .A1(n10191), .A2(n10190), .ZN(n15001) );
  INV_X1 U9968 ( .A(n15059), .ZN(n12697) );
  INV_X1 U9969 ( .A(n12213), .ZN(n12704) );
  INV_X2 U9970 ( .A(n15147), .ZN(n15149) );
  OR2_X1 U9971 ( .A1(n10493), .A2(n9684), .ZN(n15147) );
  INV_X1 U9972 ( .A(n12298), .ZN(n12808) );
  INV_X2 U9973 ( .A(n15137), .ZN(n15136) );
  INV_X1 U9974 ( .A(n9692), .ZN(n12848) );
  INV_X1 U9975 ( .A(n8231), .ZN(n11450) );
  INV_X1 U9976 ( .A(SI_16_), .ZN(n10070) );
  INV_X1 U9977 ( .A(n11067), .ZN(n11076) );
  NAND2_X1 U9978 ( .A1(n9479), .A2(P3_U3151), .ZN(n14376) );
  INV_X1 U9979 ( .A(n13093), .ZN(n13023) );
  OR2_X1 U9980 ( .A1(n9789), .A2(n9778), .ZN(n13082) );
  INV_X1 U9981 ( .A(n9107), .ZN(n13097) );
  NAND2_X1 U9982 ( .A1(n8947), .A2(n8946), .ZN(n13098) );
  AND2_X1 U9983 ( .A1(n11202), .A2(n11201), .ZN(n11440) );
  NAND2_X1 U9984 ( .A1(n13402), .A2(n13188), .ZN(n14868) );
  INV_X1 U9985 ( .A(n13402), .ZN(n13456) );
  NAND2_X1 U9986 ( .A1(n13402), .A2(n10656), .ZN(n14871) );
  INV_X1 U9987 ( .A(n13402), .ZN(n14890) );
  INV_X1 U9988 ( .A(n14974), .ZN(n14971) );
  INV_X1 U9989 ( .A(n14959), .ZN(n14958) );
  NOR2_X1 U9990 ( .A1(n14897), .A2(n14891), .ZN(n14892) );
  AND2_X1 U9991 ( .A1(n14895), .A2(n10651), .ZN(n14896) );
  INV_X1 U9992 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13581) );
  AND2_X1 U9993 ( .A1(n10462), .A2(n12043), .ZN(n15303) );
  INV_X1 U9994 ( .A(n15311), .ZN(n14530) );
  NAND4_X1 U9995 ( .A1(n9547), .A2(n9546), .A3(n9545), .A4(n9544), .ZN(n14030)
         );
  OR2_X1 U9996 ( .A1(n9429), .A2(n9428), .ZN(n14195) );
  INV_X1 U9997 ( .A(n14618), .ZN(n13866) );
  OR2_X1 U9998 ( .A1(n14596), .A2(n13877), .ZN(n14602) );
  INV_X1 U9999 ( .A(n14594), .ZN(n14611) );
  INV_X1 U10000 ( .A(n14231), .ZN(n14625) );
  OR2_X1 U10001 ( .A1(n14656), .A2(n9608), .ZN(n14202) );
  INV_X2 U10002 ( .A(n14231), .ZN(n14656) );
  OR2_X1 U10003 ( .A1(n10172), .A2(n10171), .ZN(n14759) );
  OR2_X1 U10004 ( .A1(n10172), .A2(n10164), .ZN(n14749) );
  INV_X1 U10005 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10851) );
  INV_X1 U10006 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10123) );
  INV_X2 U10007 ( .A(n12352), .ZN(P3_U3897) );
  INV_X1 U10008 ( .A(n13117), .ZN(P2_U3947) );
  INV_X1 U10009 ( .A(n13878), .ZN(P1_U4016) );
  NOR2_X1 U10010 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), 
        .ZN(n7666) );
  NOR2_X1 U10011 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n7665) );
  NOR2_X1 U10012 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), 
        .ZN(n7664) );
  NOR2_X1 U10013 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), 
        .ZN(n7663) );
  NAND2_X1 U10014 ( .A1(n7674), .A2(n7672), .ZN(n12850) );
  INV_X1 U10015 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15080) );
  OR2_X1 U10016 ( .A1(n11604), .A2(n15080), .ZN(n7682) );
  INV_X1 U10017 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10263) );
  OR2_X1 U10018 ( .A1(n9662), .A2(n10263), .ZN(n7681) );
  INV_X1 U10019 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n7679) );
  OR2_X1 U10020 ( .A1(n11608), .A2(n7679), .ZN(n7680) );
  NAND4_X2 U10021 ( .A1(n7683), .A2(n7682), .A3(n7681), .A4(n7680), .ZN(n12772) );
  XNOR2_X2 U10022 ( .A(n7685), .B(n7684), .ZN(n8191) );
  INV_X1 U10023 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7686) );
  NAND2_X4 U10024 ( .A1(n10176), .A2(n6439), .ZN(n8027) );
  INV_X1 U10025 ( .A(n7705), .ZN(n7690) );
  INV_X1 U10026 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9823) );
  NAND2_X1 U10027 ( .A1(n9823), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7691) );
  XNOR2_X1 U10028 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7721) );
  XNOR2_X1 U10029 ( .A(n7722), .B(n7721), .ZN(n9849) );
  OR2_X1 U10030 ( .A1(n8027), .A2(n9849), .ZN(n7693) );
  OR2_X1 U10031 ( .A1(n6441), .A2(SI_2_), .ZN(n7692) );
  NAND2_X1 U10032 ( .A1(n12772), .A2(n15063), .ZN(n11633) );
  NAND2_X1 U10033 ( .A1(n7726), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7698) );
  INV_X1 U10034 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10501) );
  OR2_X1 U10035 ( .A1(n11604), .A2(n10501), .ZN(n7697) );
  INV_X1 U10036 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n12053) );
  OR2_X1 U10037 ( .A1(n9662), .A2(n12053), .ZN(n7696) );
  INV_X1 U10038 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n7694) );
  OR2_X1 U10039 ( .A1(n8029), .A2(n7694), .ZN(n7695) );
  NAND4_X1 U10040 ( .A1(n7698), .A2(n7697), .A3(n7696), .A4(n7695), .ZN(n12771) );
  INV_X1 U10041 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10179) );
  INV_X1 U10042 ( .A(SI_0_), .ZN(n9831) );
  OR2_X1 U10043 ( .A1(n6441), .A2(n9831), .ZN(n7701) );
  INV_X1 U10044 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8344) );
  NAND2_X1 U10045 ( .A1(n8344), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7699) );
  AND2_X1 U10046 ( .A1(n7705), .A2(n7699), .ZN(n9832) );
  INV_X1 U10047 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n7702) );
  INV_X1 U10048 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15082) );
  NAND2_X1 U10049 ( .A1(n11603), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7704) );
  INV_X1 U10050 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7703) );
  OR2_X1 U10051 ( .A1(n7772), .A2(n6718), .ZN(n7711) );
  XNOR2_X1 U10052 ( .A(n7705), .B(n7706), .ZN(n9826) );
  OR2_X1 U10053 ( .A1(n8027), .A2(n9826), .ZN(n7710) );
  NAND2_X1 U10054 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n7707) );
  OR2_X1 U10055 ( .A1(n10176), .A2(n6433), .ZN(n7709) );
  NAND2_X1 U10056 ( .A1(n7712), .A2(n11630), .ZN(n15056) );
  NAND2_X1 U10057 ( .A1(n11603), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7718) );
  INV_X1 U10058 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n7713) );
  OR2_X1 U10059 ( .A1(n11604), .A2(n7713), .ZN(n7716) );
  INV_X1 U10060 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n7714) );
  OR2_X1 U10061 ( .A1(n11608), .A2(n7714), .ZN(n7715) );
  NAND2_X1 U10062 ( .A1(n7719), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7720) );
  INV_X1 U10063 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9824) );
  NAND2_X1 U10064 ( .A1(n9824), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7723) );
  XNOR2_X1 U10065 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7738) );
  XNOR2_X1 U10066 ( .A(n7739), .B(n7738), .ZN(n9853) );
  OR2_X1 U10067 ( .A1(n8027), .A2(n9853), .ZN(n7725) );
  OR2_X1 U10068 ( .A1(n6441), .A2(SI_3_), .ZN(n7724) );
  NAND2_X1 U10069 ( .A1(n15067), .A2(n15057), .ZN(n11645) );
  INV_X1 U10070 ( .A(n15041), .ZN(n15055) );
  NAND2_X1 U10071 ( .A1(n15056), .A2(n15055), .ZN(n15054) );
  NAND2_X1 U10072 ( .A1(n7726), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7732) );
  INV_X1 U10073 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10374) );
  OR2_X1 U10074 ( .A1(n11604), .A2(n10374), .ZN(n7731) );
  NOR2_X1 U10075 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7747) );
  AND2_X1 U10076 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7727) );
  NOR2_X1 U10077 ( .A1(n7747), .A2(n7727), .ZN(n11016) );
  OR2_X1 U10078 ( .A1(n8029), .A2(n11016), .ZN(n7730) );
  INV_X1 U10079 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n7728) );
  OR2_X1 U10080 ( .A1(n9662), .A2(n7728), .ZN(n7729) );
  NAND4_X1 U10081 ( .A1(n7732), .A2(n7731), .A3(n7730), .A4(n7729), .ZN(n15030) );
  NAND2_X1 U10082 ( .A1(n7733), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7734) );
  MUX2_X1 U10083 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7734), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7737) );
  INV_X1 U10084 ( .A(n7735), .ZN(n7736) );
  NAND2_X1 U10085 ( .A1(n9825), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U10086 ( .A1(n7741), .A2(n7740), .ZN(n7755) );
  XNOR2_X1 U10087 ( .A(n7755), .B(n7754), .ZN(n9847) );
  OR2_X1 U10088 ( .A1(n8027), .A2(n9847), .ZN(n7743) );
  OR2_X1 U10089 ( .A1(n6441), .A2(SI_4_), .ZN(n7742) );
  OAI211_X1 U10090 ( .C1(n10379), .C2(n6432), .A(n7743), .B(n7742), .ZN(n15103) );
  OR2_X1 U10091 ( .A1(n15030), .A2(n15103), .ZN(n11650) );
  NAND2_X1 U10092 ( .A1(n15030), .A2(n15103), .ZN(n11649) );
  NAND2_X1 U10093 ( .A1(n11650), .A2(n11649), .ZN(n11018) );
  NAND2_X1 U10094 ( .A1(n11015), .A2(n11759), .ZN(n7744) );
  NAND2_X1 U10095 ( .A1(n11603), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7753) );
  INV_X1 U10096 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n7745) );
  OR2_X1 U10097 ( .A1(n11604), .A2(n7745), .ZN(n7752) );
  NAND2_X1 U10098 ( .A1(n7747), .A2(n7746), .ZN(n7763) );
  OR2_X1 U10099 ( .A1(n7747), .A2(n7746), .ZN(n7748) );
  AND2_X1 U10100 ( .A1(n7763), .A2(n7748), .ZN(n11008) );
  OR2_X1 U10101 ( .A1(n8029), .A2(n11008), .ZN(n7751) );
  INV_X1 U10102 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n7749) );
  OR2_X1 U10103 ( .A1(n11608), .A2(n7749), .ZN(n7750) );
  NAND4_X1 U10104 ( .A1(n7753), .A2(n7752), .A3(n7751), .A4(n7750), .ZN(n12359) );
  OR2_X1 U10105 ( .A1(n6441), .A2(SI_5_), .ZN(n7761) );
  NAND2_X1 U10106 ( .A1(n7755), .A2(n7754), .ZN(n7757) );
  NAND2_X1 U10107 ( .A1(n9828), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U10108 ( .A1(n7757), .A2(n7756), .ZN(n7774) );
  XNOR2_X1 U10109 ( .A(n7774), .B(n7773), .ZN(n9855) );
  OR2_X1 U10110 ( .A1(n8027), .A2(n9855), .ZN(n7760) );
  OR2_X1 U10111 ( .A1(n7735), .A2(n7937), .ZN(n7758) );
  XNOR2_X1 U10112 ( .A(n7758), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10471) );
  OR2_X1 U10113 ( .A1(n10176), .A2(n10471), .ZN(n7759) );
  NAND2_X1 U10114 ( .A1(n12359), .A2(n15035), .ZN(n11654) );
  NAND2_X1 U10115 ( .A1(n11653), .A2(n11654), .ZN(n8160) );
  NAND2_X1 U10116 ( .A1(n9659), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7769) );
  INV_X1 U10117 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n7762) );
  OR2_X1 U10118 ( .A1(n9662), .A2(n7762), .ZN(n7768) );
  NAND2_X1 U10119 ( .A1(n7763), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7764) );
  AND2_X1 U10120 ( .A1(n7780), .A2(n7764), .ZN(n11334) );
  OR2_X1 U10121 ( .A1(n8029), .A2(n11334), .ZN(n7767) );
  INV_X1 U10122 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n7765) );
  OR2_X1 U10123 ( .A1(n11608), .A2(n7765), .ZN(n7766) );
  OR2_X1 U10124 ( .A1(n7770), .A2(n7937), .ZN(n7771) );
  XNOR2_X1 U10125 ( .A(n7771), .B(n7787), .ZN(n10577) );
  INV_X1 U10126 ( .A(SI_6_), .ZN(n9829) );
  NAND2_X1 U10127 ( .A1(n7774), .A2(n7773), .ZN(n7777) );
  INV_X1 U10128 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U10129 ( .A1(n7775), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7776) );
  XNOR2_X1 U10130 ( .A(n9860), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7778) );
  XNOR2_X1 U10131 ( .A(n7791), .B(n7778), .ZN(n9830) );
  OR2_X1 U10132 ( .A1(n8027), .A2(n9830), .ZN(n7779) );
  OAI211_X1 U10133 ( .C1(n10176), .C2(n10577), .A(n6538), .B(n7779), .ZN(
        n11050) );
  NAND2_X1 U10134 ( .A1(n7726), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7786) );
  INV_X1 U10135 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11311) );
  OR2_X1 U10136 ( .A1(n11604), .A2(n11311), .ZN(n7785) );
  AND2_X1 U10137 ( .A1(n7780), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7781) );
  NOR2_X1 U10138 ( .A1(n7798), .A2(n7781), .ZN(n11313) );
  OR2_X1 U10139 ( .A1(n8029), .A2(n11313), .ZN(n7784) );
  INV_X1 U10140 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n7782) );
  OR2_X1 U10141 ( .A1(n9662), .A2(n7782), .ZN(n7783) );
  NAND2_X1 U10142 ( .A1(n7770), .A2(n7787), .ZN(n7809) );
  NAND2_X1 U10143 ( .A1(n7809), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7789) );
  INV_X1 U10144 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7788) );
  XNOR2_X1 U10145 ( .A(n7789), .B(n7788), .ZN(n10772) );
  NAND2_X1 U10146 ( .A1(n9857), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7792) );
  XNOR2_X1 U10147 ( .A(n7807), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n7804) );
  XNOR2_X1 U10148 ( .A(n7806), .B(n7804), .ZN(n9851) );
  OR2_X1 U10149 ( .A1(n8027), .A2(n9851), .ZN(n7794) );
  OR2_X1 U10150 ( .A1(n6441), .A2(SI_7_), .ZN(n7793) );
  OAI211_X1 U10151 ( .C1(n10779), .C2(n10176), .A(n7794), .B(n7793), .ZN(
        n11312) );
  OR2_X1 U10152 ( .A1(n12358), .A2(n11312), .ZN(n11663) );
  NAND2_X1 U10153 ( .A1(n12358), .A2(n11312), .ZN(n11664) );
  NAND2_X1 U10154 ( .A1(n7795), .A2(n11663), .ZN(n11089) );
  NAND2_X1 U10155 ( .A1(n7726), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7803) );
  INV_X1 U10156 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11099) );
  OR2_X1 U10157 ( .A1(n11604), .A2(n11099), .ZN(n7802) );
  INV_X1 U10158 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n7796) );
  OR2_X1 U10159 ( .A1(n9662), .A2(n7796), .ZN(n7801) );
  NOR2_X1 U10160 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  OR2_X1 U10161 ( .A1(n7814), .A2(n7799), .ZN(n11097) );
  INV_X1 U10162 ( .A(n11097), .ZN(n11419) );
  OR2_X1 U10163 ( .A1(n8029), .A2(n11419), .ZN(n7800) );
  NAND4_X1 U10164 ( .A1(n7803), .A2(n7802), .A3(n7801), .A4(n7800), .ZN(n12357) );
  INV_X1 U10165 ( .A(SI_8_), .ZN(n15221) );
  OR2_X1 U10166 ( .A1(n6441), .A2(n15221), .ZN(n7813) );
  INV_X1 U10167 ( .A(n7804), .ZN(n7805) );
  NAND2_X1 U10168 ( .A1(n7807), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7808) );
  XNOR2_X1 U10169 ( .A(n7823), .B(n7822), .ZN(n9827) );
  OR2_X1 U10170 ( .A1(n8027), .A2(n9827), .ZN(n7812) );
  NAND2_X1 U10171 ( .A1(n7820), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7810) );
  XNOR2_X1 U10172 ( .A(n7810), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11067) );
  OR2_X1 U10173 ( .A1(n10176), .A2(n11076), .ZN(n7811) );
  NAND2_X1 U10174 ( .A1(n12357), .A2(n11410), .ZN(n11669) );
  NAND2_X1 U10175 ( .A1(n7726), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7819) );
  INV_X1 U10176 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14984) );
  OR2_X1 U10177 ( .A1(n11604), .A2(n14984), .ZN(n7818) );
  OR2_X1 U10178 ( .A1(n7814), .A2(n11537), .ZN(n7815) );
  AND2_X1 U10179 ( .A1(n7827), .A2(n7815), .ZN(n11227) );
  OR2_X1 U10180 ( .A1(n8029), .A2(n11227), .ZN(n7817) );
  INV_X1 U10181 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15145) );
  OR2_X1 U10182 ( .A1(n9662), .A2(n15145), .ZN(n7816) );
  NAND4_X1 U10183 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .ZN(n12356) );
  NOR2_X1 U10184 ( .A1(n7820), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7835) );
  OR2_X1 U10185 ( .A1(n7835), .A2(n7937), .ZN(n7821) );
  INV_X1 U10186 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7834) );
  XNOR2_X1 U10187 ( .A(n7821), .B(n7834), .ZN(n14990) );
  INV_X1 U10188 ( .A(n14990), .ZN(n11078) );
  XNOR2_X1 U10189 ( .A(n6626), .B(P1_DATAO_REG_9__SCAN_IN), .ZN(n7837) );
  XNOR2_X1 U10190 ( .A(n7839), .B(n7837), .ZN(n14371) );
  OR2_X1 U10191 ( .A1(n8027), .A2(n14371), .ZN(n7826) );
  OR2_X1 U10192 ( .A1(n6441), .A2(SI_9_), .ZN(n7825) );
  OAI211_X1 U10193 ( .C1(n11078), .C2(n10176), .A(n7826), .B(n7825), .ZN(
        n11529) );
  OR2_X1 U10194 ( .A1(n12356), .A2(n11529), .ZN(n11672) );
  NAND2_X1 U10195 ( .A1(n12356), .A2(n11529), .ZN(n11673) );
  NAND2_X1 U10196 ( .A1(n9659), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7833) );
  INV_X1 U10197 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11070) );
  OR2_X1 U10198 ( .A1(n9662), .A2(n11070), .ZN(n7832) );
  NAND2_X1 U10199 ( .A1(n7827), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7828) );
  AND2_X1 U10200 ( .A1(n7846), .A2(n7828), .ZN(n12196) );
  OR2_X1 U10201 ( .A1(n8029), .A2(n12196), .ZN(n7831) );
  INV_X1 U10202 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n7829) );
  OR2_X1 U10203 ( .A1(n11608), .A2(n7829), .ZN(n7830) );
  NAND4_X1 U10204 ( .A1(n7833), .A2(n7832), .A3(n7831), .A4(n7830), .ZN(n14467) );
  NAND2_X1 U10205 ( .A1(n7835), .A2(n7834), .ZN(n7859) );
  NAND2_X1 U10206 ( .A1(n7859), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7836) );
  INV_X1 U10207 ( .A(n7837), .ZN(n7838) );
  NAND2_X1 U10208 ( .A1(n7839), .A2(n7838), .ZN(n7841) );
  NAND2_X1 U10209 ( .A1(n6626), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7840) );
  XNOR2_X1 U10210 ( .A(n9926), .B(P1_DATAO_REG_10__SCAN_IN), .ZN(n7853) );
  XNOR2_X1 U10211 ( .A(n7855), .B(n7853), .ZN(n9845) );
  OR2_X1 U10212 ( .A1(n8027), .A2(n9845), .ZN(n7842) );
  OAI211_X1 U10213 ( .C1(n15018), .C2(n6432), .A(n7842), .B(n6537), .ZN(n12129) );
  OR2_X1 U10214 ( .A1(n14467), .A2(n12129), .ZN(n11677) );
  NAND2_X1 U10215 ( .A1(n14467), .A2(n12129), .ZN(n11678) );
  NAND2_X1 U10216 ( .A1(n11677), .A2(n11678), .ZN(n11674) );
  INV_X1 U10217 ( .A(n11674), .ZN(n11764) );
  NAND2_X1 U10218 ( .A1(n7843), .A2(n11678), .ZN(n14472) );
  NAND2_X1 U10219 ( .A1(n7726), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7852) );
  INV_X1 U10220 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n7844) );
  OR2_X1 U10221 ( .A1(n11604), .A2(n7844), .ZN(n7851) );
  INV_X1 U10222 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n7845) );
  OR2_X1 U10223 ( .A1(n9662), .A2(n7845), .ZN(n7850) );
  NAND2_X1 U10224 ( .A1(n7846), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7847) );
  NAND2_X1 U10225 ( .A1(n7866), .A2(n7847), .ZN(n14470) );
  INV_X1 U10226 ( .A(n14470), .ZN(n7848) );
  OR2_X1 U10227 ( .A1(n8029), .A2(n7848), .ZN(n7849) );
  INV_X1 U10228 ( .A(n7853), .ZN(n7854) );
  NAND2_X1 U10229 ( .A1(n9926), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7856) );
  XNOR2_X1 U10230 ( .A(n15222), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n7858) );
  XNOR2_X1 U10231 ( .A(n7873), .B(n7858), .ZN(n14373) );
  OR2_X1 U10232 ( .A1(n8027), .A2(n14373), .ZN(n7863) );
  OAI21_X1 U10233 ( .B1(n7859), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7861) );
  INV_X1 U10234 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7860) );
  XNOR2_X1 U10235 ( .A(n7861), .B(n7860), .ZN(n14375) );
  OR2_X1 U10236 ( .A1(n6432), .A2(n11241), .ZN(n7862) );
  NAND2_X1 U10237 ( .A1(n12688), .A2(n14473), .ZN(n11683) );
  NAND2_X1 U10238 ( .A1(n11684), .A2(n11683), .ZN(n14471) );
  NAND2_X1 U10239 ( .A1(n7726), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7871) );
  INV_X1 U10240 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12693) );
  OR2_X1 U10241 ( .A1(n11604), .A2(n12693), .ZN(n7870) );
  INV_X1 U10242 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U10243 ( .A1(n7866), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7867) );
  AND2_X1 U10244 ( .A1(n7884), .A2(n7867), .ZN(n12692) );
  OR2_X1 U10245 ( .A1(n8029), .A2(n12692), .ZN(n7869) );
  INV_X1 U10246 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11257) );
  OR2_X1 U10247 ( .A1(n9662), .A2(n11257), .ZN(n7868) );
  NAND4_X1 U10248 ( .A1(n7871), .A2(n7870), .A3(n7869), .A4(n7868), .ZN(n14468) );
  NAND2_X1 U10249 ( .A1(n15222), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U10250 ( .A1(n10074), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U10251 ( .A1(n10076), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U10252 ( .A1(n7892), .A2(n7875), .ZN(n7890) );
  XNOR2_X1 U10253 ( .A(n7891), .B(n7890), .ZN(n9861) );
  OR2_X1 U10254 ( .A1(n8027), .A2(n9861), .ZN(n7881) );
  OR2_X1 U10255 ( .A1(n6441), .A2(n9862), .ZN(n7880) );
  MUX2_X1 U10256 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7877), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7878) );
  NAND2_X1 U10257 ( .A1(n7878), .A2(n7902), .ZN(n11478) );
  OR2_X1 U10258 ( .A1(n10176), .A2(n11478), .ZN(n7879) );
  NAND2_X1 U10259 ( .A1(n14468), .A2(n14479), .ZN(n11688) );
  NAND2_X1 U10260 ( .A1(n7726), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7889) );
  INV_X1 U10261 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n7882) );
  OR2_X1 U10262 ( .A1(n11604), .A2(n7882), .ZN(n7888) );
  INV_X1 U10263 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12767) );
  OR2_X1 U10264 ( .A1(n9662), .A2(n12767), .ZN(n7887) );
  INV_X1 U10265 ( .A(n7884), .ZN(n7883) );
  NAND2_X1 U10266 ( .A1(n7884), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7885) );
  AND2_X1 U10267 ( .A1(n7906), .A2(n7885), .ZN(n12676) );
  OR2_X1 U10268 ( .A1(n8029), .A2(n12676), .ZN(n7886) );
  NAND4_X1 U10269 ( .A1(n7889), .A2(n7888), .A3(n7887), .A4(n7886), .ZN(n12687) );
  XNOR2_X1 U10270 ( .A(n7899), .B(n10125), .ZN(n14379) );
  NAND2_X1 U10271 ( .A1(n14379), .A2(n11616), .ZN(n7898) );
  INV_X1 U10272 ( .A(n10176), .ZN(n7994) );
  NAND2_X1 U10273 ( .A1(n7902), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7896) );
  INV_X1 U10274 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7895) );
  XNOR2_X1 U10275 ( .A(n7896), .B(n7895), .ZN(n14382) );
  AOI22_X1 U10276 ( .A1(n7995), .A2(n14377), .B1(n7994), .B2(n14382), .ZN(
        n7897) );
  NAND2_X1 U10277 ( .A1(n7898), .A2(n7897), .ZN(n12845) );
  OR2_X1 U10278 ( .A1(n12687), .A2(n12845), .ZN(n11693) );
  NAND2_X1 U10279 ( .A1(n12687), .A2(n12845), .ZN(n11692) );
  NAND2_X1 U10280 ( .A1(n10338), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U10281 ( .A1(n10339), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7901) );
  XNOR2_X1 U10282 ( .A(n7914), .B(n7913), .ZN(n9890) );
  NAND2_X1 U10283 ( .A1(n9890), .A2(n11616), .ZN(n7905) );
  NAND2_X1 U10284 ( .A1(n7936), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7903) );
  XNOR2_X1 U10285 ( .A(n7903), .B(n7934), .ZN(n12368) );
  AOI22_X1 U10286 ( .A1(n7995), .A2(n9889), .B1(n7994), .B2(n12368), .ZN(n7904) );
  NAND2_X1 U10287 ( .A1(n9659), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7911) );
  INV_X1 U10288 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12839) );
  OR2_X1 U10289 ( .A1(n11608), .A2(n12839), .ZN(n7910) );
  NAND2_X1 U10290 ( .A1(n7906), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7907) );
  AND2_X1 U10291 ( .A1(n7923), .A2(n7907), .ZN(n12662) );
  OR2_X1 U10292 ( .A1(n8029), .A2(n12662), .ZN(n7909) );
  INV_X1 U10293 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12763) );
  OR2_X1 U10294 ( .A1(n9662), .A2(n12763), .ZN(n7908) );
  NAND4_X1 U10295 ( .A1(n7911), .A2(n7910), .A3(n7909), .A4(n7908), .ZN(n12673) );
  NAND2_X1 U10296 ( .A1(n12841), .A2(n12673), .ZN(n11698) );
  INV_X1 U10297 ( .A(n11698), .ZN(n7912) );
  OR2_X1 U10298 ( .A1(n12841), .A2(n12673), .ZN(n11703) );
  NAND2_X1 U10299 ( .A1(n10390), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U10300 ( .A1(n10405), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n7917) );
  XNOR2_X1 U10301 ( .A(n7930), .B(n7929), .ZN(n14386) );
  NAND2_X1 U10302 ( .A1(n14386), .A2(n11616), .ZN(n7920) );
  OAI21_X1 U10303 ( .B1(n7936), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7918) );
  XNOR2_X1 U10304 ( .A(n7918), .B(n7933), .ZN(n14391) );
  AOI22_X1 U10305 ( .A1(n7995), .A2(n8384), .B1(n7994), .B2(n14391), .ZN(n7919) );
  NAND2_X1 U10306 ( .A1(n7726), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7928) );
  INV_X1 U10307 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12391) );
  OR2_X1 U10308 ( .A1(n11604), .A2(n12391), .ZN(n7927) );
  INV_X1 U10309 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10310 ( .A1(n7923), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7924) );
  AND2_X1 U10311 ( .A1(n7941), .A2(n7924), .ZN(n12649) );
  OR2_X1 U10312 ( .A1(n8029), .A2(n12649), .ZN(n7926) );
  INV_X1 U10313 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12759) );
  OR2_X1 U10314 ( .A1(n9662), .A2(n12759), .ZN(n7925) );
  NAND4_X1 U10315 ( .A1(n7928), .A2(n7927), .A3(n7926), .A4(n7925), .ZN(n12659) );
  NAND2_X1 U10316 ( .A1(n12837), .A2(n12659), .ZN(n11697) );
  NAND2_X1 U10317 ( .A1(n11704), .A2(n11697), .ZN(n12644) );
  INV_X1 U10318 ( .A(n12644), .ZN(n12641) );
  NAND2_X1 U10319 ( .A1(n10312), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10320 ( .A1(n10335), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n7932) );
  NAND2_X1 U10321 ( .A1(n7949), .A2(n7932), .ZN(n7947) );
  XNOR2_X1 U10322 ( .A(n7948), .B(n7947), .ZN(n10069) );
  NAND2_X1 U10323 ( .A1(n10069), .A2(n11616), .ZN(n7940) );
  NAND2_X1 U10324 ( .A1(n7934), .A2(n7933), .ZN(n7935) );
  OR2_X1 U10325 ( .A1(n7956), .A2(n7937), .ZN(n7938) );
  XNOR2_X1 U10326 ( .A(n7938), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U10327 ( .A1(n7995), .A2(SI_16_), .B1(n7994), .B2(n12449), .ZN(
        n7939) );
  NAND2_X1 U10328 ( .A1(n7726), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7946) );
  INV_X1 U10329 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12637) );
  OR2_X1 U10330 ( .A1(n11604), .A2(n12637), .ZN(n7945) );
  NAND2_X1 U10331 ( .A1(n7941), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7942) );
  AND2_X1 U10332 ( .A1(n7963), .A2(n7942), .ZN(n12636) );
  OR2_X1 U10333 ( .A1(n8029), .A2(n12636), .ZN(n7944) );
  INV_X1 U10334 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12448) );
  OR2_X1 U10335 ( .A1(n9662), .A2(n12448), .ZN(n7943) );
  OR2_X1 U10336 ( .A1(n12831), .A2(n12615), .ZN(n11696) );
  NAND2_X1 U10337 ( .A1(n12831), .A2(n12615), .ZN(n11702) );
  NAND2_X1 U10338 ( .A1(n11696), .A2(n11702), .ZN(n12626) );
  INV_X1 U10339 ( .A(n12626), .ZN(n12631) );
  NAND2_X1 U10340 ( .A1(n12632), .A2(n12631), .ZN(n12634) );
  NAND2_X1 U10341 ( .A1(n12634), .A2(n11702), .ZN(n12611) );
  NAND2_X1 U10342 ( .A1(n7950), .A2(n7949), .ZN(n7953) );
  NAND2_X1 U10343 ( .A1(n10388), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U10344 ( .A1(n10396), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7951) );
  OR2_X1 U10345 ( .A1(n7953), .A2(n7952), .ZN(n7954) );
  NAND2_X1 U10346 ( .A1(n7970), .A2(n7954), .ZN(n10077) );
  NAND2_X1 U10347 ( .A1(n10077), .A2(n11616), .ZN(n7960) );
  NAND2_X1 U10348 ( .A1(n7956), .A2(n7955), .ZN(n7975) );
  NAND2_X1 U10349 ( .A1(n7975), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7958) );
  INV_X1 U10350 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7957) );
  XNOR2_X1 U10351 ( .A(n7958), .B(n7957), .ZN(n12450) );
  AOI22_X1 U10352 ( .A1(n7995), .A2(n10078), .B1(n7994), .B2(n12450), .ZN(
        n7959) );
  NAND2_X1 U10353 ( .A1(n7726), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7968) );
  INV_X1 U10354 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14432) );
  OR2_X1 U10355 ( .A1(n11604), .A2(n14432), .ZN(n7967) );
  INV_X1 U10356 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U10357 ( .A1(n7963), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7964) );
  AND2_X1 U10358 ( .A1(n7979), .A2(n7964), .ZN(n12619) );
  OR2_X1 U10359 ( .A1(n8029), .A2(n12619), .ZN(n7966) );
  INV_X1 U10360 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12749) );
  OR2_X1 U10361 ( .A1(n9662), .A2(n12749), .ZN(n7965) );
  NAND4_X1 U10362 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n12628) );
  NAND2_X1 U10363 ( .A1(n12828), .A2(n12628), .ZN(n11712) );
  NAND2_X1 U10364 ( .A1(n11715), .A2(n11712), .ZN(n12613) );
  INV_X1 U10365 ( .A(n12613), .ZN(n12610) );
  NAND2_X1 U10366 ( .A1(n10554), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10367 ( .A1(n10565), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7971) );
  OR2_X1 U10368 ( .A1(n7973), .A2(n7972), .ZN(n7974) );
  NAND2_X1 U10369 ( .A1(n7987), .A2(n7974), .ZN(n10141) );
  OR2_X1 U10370 ( .A1(n10141), .A2(n8027), .ZN(n7978) );
  NAND2_X1 U10371 ( .A1(n6476), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7976) );
  XNOR2_X1 U10372 ( .A(n7976), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U10373 ( .A1(n7995), .A2(SI_18_), .B1(n7994), .B2(n12453), .ZN(
        n7977) );
  NAND2_X1 U10374 ( .A1(n7978), .A2(n7977), .ZN(n12313) );
  NAND2_X1 U10375 ( .A1(n9659), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7984) );
  INV_X1 U10376 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12745) );
  OR2_X1 U10377 ( .A1(n9662), .A2(n12745), .ZN(n7983) );
  NAND2_X1 U10378 ( .A1(n7979), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7980) );
  AND2_X1 U10379 ( .A1(n8000), .A2(n7980), .ZN(n12317) );
  OR2_X1 U10380 ( .A1(n8029), .A2(n12317), .ZN(n7982) );
  INV_X1 U10381 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12822) );
  OR2_X1 U10382 ( .A1(n11608), .A2(n12822), .ZN(n7981) );
  OR2_X1 U10383 ( .A1(n12313), .A2(n12618), .ZN(n11711) );
  NAND2_X1 U10384 ( .A1(n12313), .A2(n12618), .ZN(n11714) );
  NAND2_X1 U10385 ( .A1(n10851), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8008) );
  INV_X1 U10386 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10853) );
  NAND2_X1 U10387 ( .A1(n10853), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n7988) );
  OR2_X1 U10388 ( .A1(n7990), .A2(n7989), .ZN(n7991) );
  NAND2_X1 U10389 ( .A1(n8009), .A2(n7991), .ZN(n10224) );
  OR2_X1 U10390 ( .A1(n10224), .A2(n8027), .ZN(n7997) );
  AOI22_X1 U10391 ( .A1(n7995), .A2(SI_19_), .B1(n11785), .B2(n7994), .ZN(
        n7996) );
  NAND2_X1 U10392 ( .A1(n7997), .A2(n7996), .ZN(n12197) );
  NAND2_X1 U10393 ( .A1(n7726), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8005) );
  INV_X1 U10394 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12594) );
  OR2_X1 U10395 ( .A1(n11604), .A2(n12594), .ZN(n8004) );
  INV_X1 U10396 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U10397 ( .A1(n8000), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8001) );
  AND2_X1 U10398 ( .A1(n8012), .A2(n8001), .ZN(n12593) );
  OR2_X1 U10399 ( .A1(n8029), .A2(n12593), .ZN(n8003) );
  INV_X1 U10400 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12741) );
  OR2_X1 U10401 ( .A1(n9662), .A2(n12741), .ZN(n8002) );
  OR2_X1 U10402 ( .A1(n12197), .A2(n12604), .ZN(n11718) );
  INV_X1 U10403 ( .A(n11718), .ZN(n8006) );
  NAND2_X1 U10404 ( .A1(n12197), .A2(n12604), .ZN(n11719) );
  INV_X1 U10405 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11014) );
  XNOR2_X1 U10406 ( .A(n8018), .B(n11014), .ZN(n10423) );
  NAND2_X1 U10407 ( .A1(n10423), .A2(n11616), .ZN(n8011) );
  OR2_X1 U10408 ( .A1(n6441), .A2(n10424), .ZN(n8010) );
  NAND2_X1 U10409 ( .A1(n11603), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8017) );
  INV_X1 U10410 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12579) );
  OR2_X1 U10411 ( .A1(n11604), .A2(n12579), .ZN(n8016) );
  NAND2_X1 U10412 ( .A1(n8012), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8013) );
  AND2_X1 U10413 ( .A1(n8031), .A2(n8013), .ZN(n12578) );
  OR2_X1 U10414 ( .A1(n12578), .A2(n8029), .ZN(n8015) );
  INV_X1 U10415 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n15180) );
  OR2_X1 U10416 ( .A1(n11608), .A2(n15180), .ZN(n8014) );
  XNOR2_X1 U10417 ( .A(n12815), .B(n12563), .ZN(n12572) );
  INV_X1 U10418 ( .A(n12572), .ZN(n12581) );
  OR2_X1 U10419 ( .A1(n12815), .A2(n12563), .ZN(n11723) );
  NAND2_X1 U10420 ( .A1(n12580), .A2(n11723), .ZN(n12557) );
  INV_X1 U10421 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U10422 ( .A1(n11136), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8039) );
  INV_X1 U10423 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U10424 ( .A1(n11139), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8023) );
  NAND2_X1 U10425 ( .A1(n8039), .A2(n8023), .ZN(n8024) );
  NAND2_X1 U10426 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  NAND2_X1 U10427 ( .A1(n8040), .A2(n8026), .ZN(n10517) );
  OR2_X1 U10428 ( .A1(n10517), .A2(n8027), .ZN(n8028) );
  INV_X1 U10429 ( .A(SI_21_), .ZN(n10516) );
  NAND2_X1 U10430 ( .A1(n8031), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10431 ( .A1(n8044), .A2(n8032), .ZN(n12566) );
  NAND2_X1 U10432 ( .A1(n8193), .A2(n12566), .ZN(n8037) );
  INV_X1 U10433 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12810) );
  OR2_X1 U10434 ( .A1(n11608), .A2(n12810), .ZN(n8036) );
  INV_X1 U10435 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n8033) );
  OR2_X1 U10436 ( .A1(n11604), .A2(n8033), .ZN(n8035) );
  INV_X1 U10437 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12731) );
  OR2_X1 U10438 ( .A1(n9662), .A2(n12731), .ZN(n8034) );
  NAND2_X1 U10439 ( .A1(n12565), .A2(n12574), .ZN(n11728) );
  NAND2_X1 U10440 ( .A1(n12557), .A2(n11728), .ZN(n8038) );
  NAND2_X1 U10441 ( .A1(n8038), .A2(n11727), .ZN(n12550) );
  INV_X1 U10442 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11494) );
  XNOR2_X1 U10443 ( .A(n11494), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8051) );
  XNOR2_X1 U10444 ( .A(n8052), .B(n8051), .ZN(n10621) );
  NAND2_X1 U10445 ( .A1(n10621), .A2(n11616), .ZN(n8043) );
  INV_X1 U10446 ( .A(SI_22_), .ZN(n8041) );
  NAND2_X1 U10447 ( .A1(n8044), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U10448 ( .A1(n8057), .A2(n8045), .ZN(n12552) );
  NAND2_X1 U10449 ( .A1(n12552), .A2(n8193), .ZN(n8049) );
  NAND2_X1 U10450 ( .A1(n9659), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10451 ( .A1(n11603), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10452 ( .A1(n7726), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8046) );
  NAND4_X1 U10453 ( .A1(n8049), .A2(n8048), .A3(n8047), .A4(n8046), .ZN(n12353) );
  NAND2_X1 U10454 ( .A1(n12298), .A2(n12564), .ZN(n11732) );
  NAND2_X1 U10455 ( .A1(n12550), .A2(n11732), .ZN(n8050) );
  NAND2_X1 U10456 ( .A1(n11494), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8053) );
  XNOR2_X1 U10457 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8064) );
  XNOR2_X1 U10458 ( .A(n8065), .B(n8064), .ZN(n10854) );
  NAND2_X1 U10459 ( .A1(n10854), .A2(n11616), .ZN(n8056) );
  INV_X1 U10460 ( .A(SI_23_), .ZN(n10856) );
  OR2_X1 U10461 ( .A1(n6441), .A2(n10856), .ZN(n8055) );
  NAND2_X1 U10462 ( .A1(n8057), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U10463 ( .A1(n8073), .A2(n8058), .ZN(n12541) );
  NAND2_X1 U10464 ( .A1(n12541), .A2(n8193), .ZN(n8063) );
  NAND2_X1 U10465 ( .A1(n7726), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10466 ( .A1(n9659), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8059) );
  AND2_X1 U10467 ( .A1(n8060), .A2(n8059), .ZN(n8062) );
  NAND2_X1 U10468 ( .A1(n11603), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U10469 ( .A1(n12540), .A2(n12549), .ZN(n11775) );
  NAND2_X1 U10470 ( .A1(n8078), .A2(n11775), .ZN(n12534) );
  INV_X1 U10471 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U10472 ( .A1(n11510), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8066) );
  INV_X1 U10473 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13589) );
  NAND2_X1 U10474 ( .A1(n8067), .A2(n13589), .ZN(n8068) );
  INV_X1 U10475 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14354) );
  XNOR2_X1 U10476 ( .A(n8079), .B(n14354), .ZN(n11102) );
  NAND2_X1 U10477 ( .A1(n11102), .A2(n11616), .ZN(n8070) );
  OR2_X1 U10478 ( .A1(n6441), .A2(n15242), .ZN(n8069) );
  INV_X1 U10479 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10480 ( .A1(n8073), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10481 ( .A1(n8084), .A2(n8074), .ZN(n12526) );
  NAND2_X1 U10482 ( .A1(n12526), .A2(n8193), .ZN(n8077) );
  AOI22_X1 U10483 ( .A1(n7726), .A2(P3_REG0_REG_24__SCAN_IN), .B1(n9659), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U10484 ( .A1(n11603), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8075) );
  INV_X1 U10485 ( .A(n8078), .ZN(n12522) );
  INV_X1 U10486 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13586) );
  XNOR2_X1 U10487 ( .A(n13586), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8093) );
  XNOR2_X1 U10488 ( .A(n8094), .B(n8093), .ZN(n11217) );
  NAND2_X1 U10489 ( .A1(n11217), .A2(n11616), .ZN(n8081) );
  INV_X1 U10490 ( .A(n8084), .ZN(n8083) );
  INV_X1 U10491 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8082) );
  NAND2_X1 U10492 ( .A1(n8084), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8085) );
  NAND2_X1 U10493 ( .A1(n8099), .A2(n8085), .ZN(n12512) );
  NAND2_X1 U10494 ( .A1(n12512), .A2(n8193), .ZN(n8091) );
  INV_X1 U10495 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U10496 ( .A1(n11603), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10497 ( .A1(n7726), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8086) );
  OAI211_X1 U10498 ( .C1(n11604), .C2(n8088), .A(n8087), .B(n8086), .ZN(n8089)
         );
  INV_X1 U10499 ( .A(n8089), .ZN(n8090) );
  INV_X1 U10500 ( .A(n12503), .ZN(n12505) );
  NAND2_X1 U10501 ( .A1(n12511), .A2(n12519), .ZN(n8092) );
  NAND2_X1 U10502 ( .A1(n13586), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8095) );
  INV_X1 U10503 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13582) );
  INV_X1 U10504 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14347) );
  AOI22_X1 U10505 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13582), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14347), .ZN(n8097) );
  XNOR2_X1 U10506 ( .A(n8107), .B(n8097), .ZN(n11447) );
  NAND2_X1 U10507 ( .A1(n11447), .A2(n11616), .ZN(n8098) );
  INV_X1 U10508 ( .A(SI_26_), .ZN(n11449) );
  NAND2_X1 U10509 ( .A1(n8099), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8100) );
  NAND2_X1 U10510 ( .A1(n8114), .A2(n8100), .ZN(n12497) );
  NAND2_X1 U10511 ( .A1(n12497), .A2(n8193), .ZN(n8105) );
  INV_X1 U10512 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12711) );
  NAND2_X1 U10513 ( .A1(n9659), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U10514 ( .A1(n7726), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8101) );
  OAI211_X1 U10515 ( .C1(n12711), .C2(n9662), .A(n8102), .B(n8101), .ZN(n8103)
         );
  INV_X1 U10516 ( .A(n8103), .ZN(n8104) );
  NAND2_X1 U10517 ( .A1(n12496), .A2(n12507), .ZN(n11739) );
  NOR2_X1 U10518 ( .A1(n14347), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10519 ( .A1(n14347), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8108) );
  XNOR2_X1 U10520 ( .A(n13581), .B(P2_DATAO_REG_27__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U10521 ( .A1(n11490), .A2(n11616), .ZN(n8111) );
  INV_X1 U10522 ( .A(SI_27_), .ZN(n11491) );
  INV_X1 U10523 ( .A(n8114), .ZN(n8113) );
  INV_X1 U10524 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U10525 ( .A1(n8113), .A2(n8112), .ZN(n8129) );
  NAND2_X1 U10526 ( .A1(n8114), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U10527 ( .A1(n8129), .A2(n8115), .ZN(n12483) );
  INV_X1 U10528 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8118) );
  NAND2_X1 U10529 ( .A1(n11603), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U10530 ( .A1(n7726), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8116) );
  OAI211_X1 U10531 ( .C1(n11604), .C2(n8118), .A(n8117), .B(n8116), .ZN(n8119)
         );
  OR2_X1 U10532 ( .A1(n12482), .A2(n12328), .ZN(n11742) );
  NAND2_X1 U10533 ( .A1(n12482), .A2(n12328), .ZN(n11747) );
  NAND2_X1 U10534 ( .A1(n11742), .A2(n11747), .ZN(n11745) );
  NAND2_X1 U10535 ( .A1(n12477), .A2(n12476), .ZN(n12475) );
  INV_X1 U10536 ( .A(n8120), .ZN(n8122) );
  INV_X1 U10537 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11590) );
  NAND2_X1 U10538 ( .A1(n11590), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U10539 ( .A1(n8122), .A2(n8121), .ZN(n8124) );
  NAND2_X1 U10540 ( .A1(n13581), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8123) );
  INV_X1 U10541 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n12057) );
  INV_X1 U10542 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14346) );
  AOI22_X1 U10543 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n12057), .B2(n14346), .ZN(n8125) );
  INV_X1 U10544 ( .A(n8125), .ZN(n8126) );
  XNOR2_X1 U10545 ( .A(n9654), .B(n8126), .ZN(n12121) );
  NAND2_X1 U10546 ( .A1(n12121), .A2(n11616), .ZN(n8128) );
  INV_X1 U10547 ( .A(SI_28_), .ZN(n12122) );
  NAND2_X1 U10548 ( .A1(n8129), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8130) );
  NAND2_X1 U10549 ( .A1(n12046), .A2(n8130), .ZN(n12468) );
  INV_X1 U10550 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12702) );
  NAND2_X1 U10551 ( .A1(n7726), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8132) );
  NAND2_X1 U10552 ( .A1(n9659), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8131) );
  OAI211_X1 U10553 ( .C1(n12702), .C2(n9662), .A(n8132), .B(n8131), .ZN(n8133)
         );
  NAND2_X1 U10554 ( .A1(n12213), .A2(n12478), .ZN(n11749) );
  XNOR2_X1 U10555 ( .A(n9671), .B(n12206), .ZN(n12467) );
  INV_X1 U10556 ( .A(n8134), .ZN(n8135) );
  NAND2_X1 U10557 ( .A1(n8135), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8136) );
  MUX2_X1 U10558 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8136), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n8137) );
  NAND2_X1 U10559 ( .A1(n12459), .A2(n10515), .ZN(n8147) );
  NAND2_X1 U10560 ( .A1(n8138), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8139) );
  MUX2_X1 U10561 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8139), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8140) );
  INV_X1 U10562 ( .A(n8140), .ZN(n8142) );
  NAND2_X1 U10563 ( .A1(n8143), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8144) );
  MUX2_X1 U10564 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8144), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8145) );
  NAND2_X1 U10565 ( .A1(n8145), .A2(n8135), .ZN(n10536) );
  AND2_X1 U10566 ( .A1(n10515), .A2(n10536), .ZN(n9678) );
  XNOR2_X1 U10567 ( .A(n8151), .B(n9678), .ZN(n8146) );
  NAND2_X1 U10568 ( .A1(n8147), .A2(n8146), .ZN(n10354) );
  INV_X1 U10569 ( .A(n10538), .ZN(n11758) );
  NAND3_X1 U10570 ( .A1(n10354), .A2(n11758), .A3(n15111), .ZN(n8150) );
  NOR2_X1 U10571 ( .A1(n8151), .A2(n10536), .ZN(n8148) );
  AND2_X1 U10572 ( .A1(n12459), .A2(n8148), .ZN(n10494) );
  INV_X1 U10573 ( .A(n10494), .ZN(n8149) );
  AND2_X1 U10574 ( .A1(n11785), .A2(n10536), .ZN(n15084) );
  NAND2_X1 U10575 ( .A1(n10546), .A2(n12770), .ZN(n8154) );
  INV_X1 U10576 ( .A(n12780), .ZN(n8152) );
  OR2_X1 U10577 ( .A1(n15068), .A2(n8152), .ZN(n8153) );
  NAND2_X1 U10578 ( .A1(n8154), .A2(n8153), .ZN(n15071) );
  NAND2_X1 U10579 ( .A1(n15071), .A2(n15070), .ZN(n15040) );
  INV_X1 U10580 ( .A(n15063), .ZN(n8155) );
  OR2_X1 U10581 ( .A1(n12772), .A2(n8155), .ZN(n15042) );
  AND2_X1 U10582 ( .A1(n15041), .A2(n15042), .ZN(n8156) );
  NAND2_X1 U10583 ( .A1(n15040), .A2(n8156), .ZN(n15039) );
  INV_X1 U10584 ( .A(n15057), .ZN(n10603) );
  NAND2_X1 U10585 ( .A1(n15067), .A2(n10603), .ZN(n8157) );
  NAND2_X1 U10586 ( .A1(n15039), .A2(n8157), .ZN(n11017) );
  NAND2_X1 U10587 ( .A1(n11017), .A2(n11018), .ZN(n8159) );
  INV_X1 U10588 ( .A(n15103), .ZN(n10909) );
  NAND2_X1 U10589 ( .A1(n15030), .A2(n10909), .ZN(n8158) );
  NAND2_X1 U10590 ( .A1(n8159), .A2(n8158), .ZN(n11305) );
  NAND2_X1 U10591 ( .A1(n15029), .A2(n11050), .ZN(n8161) );
  NAND2_X1 U10592 ( .A1(n8160), .A2(n8161), .ZN(n8165) );
  INV_X1 U10593 ( .A(n8161), .ZN(n11306) );
  NOR2_X1 U10594 ( .A1(n12359), .A2(n11007), .ZN(n11336) );
  NAND2_X1 U10595 ( .A1(n11336), .A2(n8161), .ZN(n8162) );
  OAI211_X1 U10596 ( .C1(n11332), .C2(n11306), .A(n11658), .B(n8162), .ZN(
        n8163) );
  INV_X1 U10597 ( .A(n8163), .ZN(n8164) );
  INV_X1 U10598 ( .A(n11312), .ZN(n11293) );
  INV_X1 U10599 ( .A(n11410), .ZN(n11416) );
  OR2_X1 U10600 ( .A1(n12357), .A2(n11416), .ZN(n8167) );
  INV_X1 U10601 ( .A(n11529), .ZN(n11541) );
  NAND2_X1 U10602 ( .A1(n12356), .A2(n11541), .ZN(n8170) );
  INV_X1 U10603 ( .A(n12129), .ZN(n12193) );
  NAND2_X1 U10604 ( .A1(n14465), .A2(n12302), .ZN(n8171) );
  INV_X1 U10605 ( .A(n14479), .ZN(n12236) );
  NAND2_X1 U10606 ( .A1(n14468), .A2(n12236), .ZN(n8173) );
  NAND2_X1 U10607 ( .A1(n11693), .A2(n11692), .ZN(n12671) );
  INV_X1 U10608 ( .A(n12845), .ZN(n12291) );
  NAND2_X1 U10609 ( .A1(n12687), .A2(n12291), .ZN(n8174) );
  NAND2_X1 U10610 ( .A1(n11703), .A2(n11698), .ZN(n12657) );
  INV_X1 U10611 ( .A(n12673), .ZN(n12341) );
  OR2_X1 U10612 ( .A1(n12841), .A2(n12341), .ZN(n8175) );
  INV_X1 U10613 ( .A(n12659), .ZN(n12250) );
  NAND2_X1 U10614 ( .A1(n12627), .A2(n12626), .ZN(n12625) );
  NAND2_X1 U10615 ( .A1(n12831), .A2(n12646), .ZN(n8176) );
  NAND2_X1 U10616 ( .A1(n12625), .A2(n8176), .ZN(n12614) );
  INV_X1 U10617 ( .A(n12628), .ZN(n12603) );
  OR2_X1 U10618 ( .A1(n12828), .A2(n12603), .ZN(n8177) );
  INV_X1 U10619 ( .A(n8178), .ZN(n12588) );
  NAND2_X1 U10620 ( .A1(n12197), .A2(n12355), .ZN(n8179) );
  NAND2_X1 U10621 ( .A1(n12815), .A2(n12590), .ZN(n8180) );
  NAND2_X1 U10622 ( .A1(n12571), .A2(n8180), .ZN(n12560) );
  INV_X1 U10623 ( .A(n12574), .ZN(n12354) );
  OR2_X1 U10624 ( .A1(n12565), .A2(n12354), .ZN(n8181) );
  INV_X1 U10625 ( .A(n12549), .ZN(n12265) );
  NAND2_X1 U10626 ( .A1(n12540), .A2(n12265), .ZN(n8182) );
  NAND2_X1 U10627 ( .A1(n8183), .A2(n8182), .ZN(n12517) );
  NAND2_X1 U10628 ( .A1(n12517), .A2(n12521), .ZN(n8185) );
  INV_X1 U10629 ( .A(n12536), .ZN(n12351) );
  NAND2_X1 U10630 ( .A1(n12525), .A2(n12351), .ZN(n8184) );
  NAND2_X1 U10631 ( .A1(n8185), .A2(n8184), .ZN(n12502) );
  NAND2_X1 U10632 ( .A1(n12502), .A2(n12503), .ZN(n8187) );
  NAND2_X1 U10633 ( .A1(n12511), .A2(n12489), .ZN(n8186) );
  AND2_X1 U10634 ( .A1(n12496), .A2(n12350), .ZN(n8189) );
  OR2_X1 U10635 ( .A1(n12496), .A2(n12350), .ZN(n8188) );
  OR2_X1 U10636 ( .A1(n12482), .A2(n12490), .ZN(n8190) );
  INV_X1 U10637 ( .A(n12206), .ZN(n11780) );
  NAND2_X1 U10638 ( .A1(n11785), .A2(n11793), .ZN(n9677) );
  INV_X1 U10639 ( .A(n10536), .ZN(n8228) );
  NAND2_X1 U10640 ( .A1(n11639), .A2(n8228), .ZN(n11628) );
  OAI211_X1 U10641 ( .C1(n6507), .C2(n11780), .A(n15072), .B(n9652), .ZN(n8201) );
  INV_X1 U10642 ( .A(n8191), .ZN(n9665) );
  NAND2_X1 U10643 ( .A1(n9665), .A2(n11058), .ZN(n10190) );
  NAND2_X2 U10644 ( .A1(n11793), .A2(n11639), .ZN(n11754) );
  NAND2_X1 U10645 ( .A1(n12490), .A2(n15069), .ZN(n8200) );
  INV_X1 U10646 ( .A(n12046), .ZN(n8194) );
  NAND2_X1 U10647 ( .A1(n8194), .A2(n8193), .ZN(n11611) );
  INV_X1 U10648 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U10649 ( .A1(n7726), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8196) );
  NAND2_X1 U10650 ( .A1(n9659), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8195) );
  OAI211_X1 U10651 ( .C1(n9662), .C2(n9685), .A(n8196), .B(n8195), .ZN(n8197)
         );
  INV_X1 U10652 ( .A(n8197), .ZN(n8198) );
  NAND2_X1 U10653 ( .A1(n10176), .A2(n10190), .ZN(n8199) );
  NAND2_X1 U10654 ( .A1(n8201), .A2(n7647), .ZN(n12471) );
  AOI21_X1 U10655 ( .B1(n12467), .B2(n15102), .A(n12471), .ZN(n12701) );
  NAND2_X1 U10656 ( .A1(n8202), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8203) );
  MUX2_X1 U10657 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8203), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8205) );
  NAND2_X1 U10658 ( .A1(n6475), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8206) );
  MUX2_X1 U10659 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8206), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8207) );
  NAND2_X1 U10660 ( .A1(n8207), .A2(n8202), .ZN(n11219) );
  NAND2_X1 U10661 ( .A1(n8208), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8209) );
  XNOR2_X1 U10662 ( .A(n11104), .B(P3_B_REG_SCAN_IN), .ZN(n8211) );
  INV_X1 U10663 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8212) );
  NAND2_X1 U10664 ( .A1(n9891), .A2(n8212), .ZN(n8214) );
  NAND2_X1 U10665 ( .A1(n11450), .A2(n11104), .ZN(n8213) );
  INV_X1 U10666 ( .A(n10539), .ZN(n12849) );
  INV_X1 U10667 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U10668 ( .A1(n9891), .A2(n8215), .ZN(n8217) );
  NAND2_X1 U10669 ( .A1(n11450), .A2(n11219), .ZN(n8216) );
  INV_X1 U10670 ( .A(n10496), .ZN(n12847) );
  NOR4_X1 U10671 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8226) );
  NOR4_X1 U10672 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8221) );
  NOR4_X1 U10673 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8220) );
  NOR4_X1 U10674 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8219) );
  NOR4_X1 U10675 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8218) );
  NAND4_X1 U10676 ( .A1(n8221), .A2(n8220), .A3(n8219), .A4(n8218), .ZN(n8222)
         );
  NOR4_X1 U10677 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n8223), .A4(n8222), .ZN(n8225) );
  NOR4_X1 U10678 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n8224) );
  NAND3_X1 U10679 ( .A1(n8226), .A2(n8225), .A3(n8224), .ZN(n8227) );
  NAND2_X1 U10680 ( .A1(n9891), .A2(n8227), .ZN(n9674) );
  NAND3_X1 U10681 ( .A1(n12849), .A2(n12847), .A3(n9674), .ZN(n10357) );
  NAND2_X1 U10682 ( .A1(n10515), .A2(n8228), .ZN(n11787) );
  OR2_X1 U10683 ( .A1(n9677), .A2(n11787), .ZN(n10355) );
  INV_X1 U10684 ( .A(n10354), .ZN(n8229) );
  NAND3_X1 U10685 ( .A1(n10496), .A2(n10539), .A3(n9674), .ZN(n10356) );
  OAI22_X1 U10686 ( .A1(n10357), .A2(n10355), .B1(n8229), .B2(n10356), .ZN(
        n8235) );
  NOR2_X1 U10687 ( .A1(n11219), .A2(n11104), .ZN(n8230) );
  NAND2_X1 U10688 ( .A1(n8231), .A2(n8230), .ZN(n10344) );
  INV_X1 U10689 ( .A(n8141), .ZN(n8232) );
  NAND2_X1 U10690 ( .A1(n8232), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8234) );
  XNOR2_X1 U10691 ( .A(n8234), .B(n8233), .ZN(n10177) );
  NAND2_X1 U10692 ( .A1(n8235), .A2(n10358), .ZN(n8238) );
  INV_X1 U10693 ( .A(n10357), .ZN(n8236) );
  NAND2_X1 U10694 ( .A1(n10358), .A2(n11758), .ZN(n11792) );
  NOR2_X1 U10695 ( .A1(n11792), .A2(n11754), .ZN(n10348) );
  NAND2_X1 U10696 ( .A1(n8236), .A2(n10348), .ZN(n8237) );
  OR2_X1 U10697 ( .A1(n12701), .A2(n15137), .ZN(n8242) );
  INV_X1 U10698 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8239) );
  OAI22_X1 U10699 ( .A1(n12704), .A2(n12846), .B1(n15136), .B2(n8239), .ZN(
        n8240) );
  INV_X1 U10700 ( .A(n8240), .ZN(n8241) );
  NAND2_X1 U10701 ( .A1(n8242), .A2(n8241), .ZN(P3_U3455) );
  INV_X1 U10702 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n12425) );
  NAND2_X1 U10703 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n12425), .ZN(n8243) );
  OAI21_X1 U10704 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n12425), .A(n8243), .ZN(
        n8276) );
  INV_X1 U10705 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12396) );
  XNOR2_X1 U10706 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n8278) );
  INV_X1 U10707 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12383) );
  INV_X1 U10708 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8271) );
  XNOR2_X1 U10709 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8326) );
  INV_X1 U10710 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n8269) );
  XNOR2_X1 U10711 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8282) );
  INV_X1 U10712 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n8264) );
  XNOR2_X1 U10713 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8286) );
  INV_X1 U10714 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U10715 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n15209), .ZN(n8293) );
  XNOR2_X1 U10716 ( .A(n13883), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n8290) );
  NOR2_X1 U10717 ( .A1(n8248), .A2(n8247), .ZN(n8250) );
  INV_X1 U10718 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n10381) );
  NOR2_X1 U10719 ( .A1(n8253), .A2(n10381), .ZN(n8255) );
  NOR2_X1 U10720 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n8258), .ZN(n8260) );
  XNOR2_X1 U10721 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n8258), .ZN(n8311) );
  XOR2_X1 U10722 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n8312) );
  NAND2_X1 U10723 ( .A1(n8286), .A2(n8285), .ZN(n8263) );
  NOR2_X1 U10724 ( .A1(n15228), .A2(n8283), .ZN(n8266) );
  INV_X1 U10725 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15023) );
  NAND2_X1 U10726 ( .A1(n15228), .A2(n8283), .ZN(n8265) );
  INV_X1 U10727 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10039) );
  XOR2_X1 U10728 ( .A(n11074), .B(n10039), .Z(n8323) );
  NAND2_X1 U10729 ( .A1(n8282), .A2(n8281), .ZN(n8268) );
  NAND2_X1 U10730 ( .A1(n8326), .A2(n8327), .ZN(n8270) );
  XNOR2_X1 U10731 ( .A(n12383), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n8279) );
  NOR2_X1 U10732 ( .A1(n8280), .A2(n8279), .ZN(n8272) );
  AOI21_X1 U10733 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n12383), .A(n8272), .ZN(
        n8277) );
  NAND2_X1 U10734 ( .A1(n8278), .A2(n8277), .ZN(n8273) );
  NOR2_X1 U10735 ( .A1(n8276), .A2(n8275), .ZN(n8274) );
  AOI21_X1 U10736 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n12425), .A(n8274), .ZN(
        n8332) );
  XOR2_X1 U10737 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n8332), .Z(n8334) );
  XNOR2_X1 U10738 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n8334), .ZN(n14428) );
  XNOR2_X1 U10739 ( .A(n8276), .B(n8275), .ZN(n8330) );
  XNOR2_X1 U10740 ( .A(n8278), .B(n8277), .ZN(n8328) );
  XNOR2_X1 U10741 ( .A(n8280), .B(n8279), .ZN(n14579) );
  XOR2_X1 U10742 ( .A(n8282), .B(n8281), .Z(n14571) );
  XNOR2_X1 U10743 ( .A(n15228), .B(n8283), .ZN(n8284) );
  XNOR2_X1 U10744 ( .A(n8284), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n8321) );
  XOR2_X1 U10745 ( .A(n8286), .B(n8285), .Z(n8317) );
  INV_X1 U10746 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n13935) );
  INV_X1 U10747 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14801) );
  NAND2_X1 U10748 ( .A1(n8299), .A2(n14801), .ZN(n8300) );
  XOR2_X1 U10749 ( .A(n8289), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15326) );
  XOR2_X1 U10750 ( .A(n8291), .B(n8290), .Z(n8297) );
  INV_X1 U10751 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9802) );
  NOR2_X1 U10752 ( .A1(n8294), .A2(n9802), .ZN(n8295) );
  OAI21_X1 U10753 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n15209), .A(n8293), .ZN(
        n15320) );
  NAND2_X1 U10754 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15320), .ZN(n15331) );
  NOR2_X1 U10755 ( .A1(n15331), .A2(n15330), .ZN(n15329) );
  NOR2_X1 U10756 ( .A1(n8297), .A2(n8296), .ZN(n14366) );
  NAND2_X1 U10757 ( .A1(n8297), .A2(n8296), .ZN(n14367) );
  NAND2_X1 U10758 ( .A1(n15326), .A2(n15325), .ZN(n8298) );
  NOR2_X1 U10759 ( .A1(n15326), .A2(n15325), .ZN(n15324) );
  AOI21_X1 U10760 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n8298), .A(n15324), .ZN(
        n15316) );
  NAND2_X1 U10761 ( .A1(n8301), .A2(n8302), .ZN(n8303) );
  INV_X1 U10762 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15318) );
  INV_X1 U10763 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8304) );
  NOR2_X1 U10764 ( .A1(n8305), .A2(n8304), .ZN(n8308) );
  XNOR2_X1 U10765 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n8307) );
  XNOR2_X1 U10766 ( .A(n8307), .B(n8306), .ZN(n14384) );
  INV_X1 U10767 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n8310) );
  XNOR2_X1 U10768 ( .A(n8311), .B(n13962), .ZN(n15322) );
  XNOR2_X1 U10769 ( .A(n8313), .B(n8312), .ZN(n8315) );
  NAND2_X1 U10770 ( .A1(n8314), .A2(n8315), .ZN(n8316) );
  INV_X1 U10771 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14828) );
  NOR2_X1 U10772 ( .A1(n8317), .A2(n8318), .ZN(n8319) );
  INV_X1 U10773 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14849) );
  NOR2_X1 U10774 ( .A1(n8321), .A2(n8320), .ZN(n8322) );
  INV_X1 U10775 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14398) );
  XNOR2_X1 U10776 ( .A(n8324), .B(n8323), .ZN(n14567) );
  NAND2_X1 U10777 ( .A1(n14568), .A2(n14567), .ZN(n8325) );
  XOR2_X1 U10778 ( .A(n8327), .B(n8326), .Z(n14574) );
  INV_X1 U10779 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14585) );
  NAND2_X1 U10780 ( .A1(n8330), .A2(n8331), .ZN(n14588) );
  INV_X1 U10781 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14590) );
  INV_X1 U10782 ( .A(n8332), .ZN(n8333) );
  NOR2_X1 U10783 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n8333), .ZN(n8336) );
  INV_X1 U10784 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14438) );
  NOR2_X1 U10785 ( .A1(n14438), .A2(n8334), .ZN(n8335) );
  NOR2_X1 U10786 ( .A1(n8336), .A2(n8335), .ZN(n8339) );
  INV_X1 U10787 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n8341) );
  XNOR2_X1 U10788 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n8341), .ZN(n8338) );
  XOR2_X1 U10789 ( .A(n8339), .B(n8338), .Z(n14362) );
  XNOR2_X1 U10790 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n8337) );
  NOR2_X1 U10791 ( .A1(n8339), .A2(n8338), .ZN(n8340) );
  AOI21_X1 U10792 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n8341), .A(n8340), .ZN(
        n8342) );
  NAND2_X1 U10793 ( .A1(n8487), .A2(n8345), .ZN(n8513) );
  NAND2_X1 U10794 ( .A1(n8348), .A2(SI_2_), .ZN(n8350) );
  OAI21_X1 U10795 ( .B1(n8348), .B2(SI_2_), .A(n8350), .ZN(n8514) );
  INV_X1 U10796 ( .A(n8514), .ZN(n8349) );
  MUX2_X1 U10797 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n6437), .Z(n8351) );
  NAND2_X1 U10798 ( .A1(n8351), .A2(SI_3_), .ZN(n8353) );
  OAI21_X1 U10799 ( .B1(n8351), .B2(SI_3_), .A(n8353), .ZN(n8352) );
  INV_X1 U10800 ( .A(n8352), .ZN(n8540) );
  NAND2_X1 U10801 ( .A1(n8541), .A2(n8540), .ZN(n8543) );
  NAND2_X1 U10802 ( .A1(n8543), .A2(n8353), .ZN(n8559) );
  NAND2_X1 U10803 ( .A1(n8354), .A2(SI_4_), .ZN(n8356) );
  OAI21_X1 U10804 ( .B1(n8354), .B2(SI_4_), .A(n8356), .ZN(n8355) );
  INV_X1 U10805 ( .A(n8355), .ZN(n8558) );
  NAND2_X1 U10806 ( .A1(n8559), .A2(n8558), .ZN(n8561) );
  MUX2_X1 U10807 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6437), .Z(n8357) );
  NAND2_X1 U10808 ( .A1(n8357), .A2(SI_5_), .ZN(n8359) );
  OAI21_X1 U10809 ( .B1(n8357), .B2(SI_5_), .A(n8359), .ZN(n8358) );
  MUX2_X1 U10810 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9479), .Z(n8360) );
  NAND2_X1 U10811 ( .A1(n8360), .A2(SI_6_), .ZN(n8362) );
  OAI21_X1 U10812 ( .B1(SI_6_), .B2(n8360), .A(n8362), .ZN(n8361) );
  INV_X1 U10813 ( .A(n8361), .ZN(n8590) );
  MUX2_X1 U10814 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9479), .Z(n8363) );
  NAND2_X1 U10815 ( .A1(n8363), .A2(SI_7_), .ZN(n8365) );
  OAI21_X1 U10816 ( .B1(n8363), .B2(SI_7_), .A(n8365), .ZN(n8612) );
  INV_X1 U10817 ( .A(n8612), .ZN(n8364) );
  MUX2_X1 U10818 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9479), .Z(n8630) );
  INV_X1 U10819 ( .A(n8658), .ZN(n8367) );
  MUX2_X1 U10820 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9479), .Z(n8368) );
  XNOR2_X1 U10821 ( .A(n8368), .B(SI_10_), .ZN(n8675) );
  NAND2_X1 U10822 ( .A1(n8368), .A2(SI_10_), .ZN(n8369) );
  MUX2_X1 U10823 ( .A(n10004), .B(n15222), .S(n9833), .Z(n8372) );
  NAND2_X1 U10824 ( .A1(n8372), .A2(n8371), .ZN(n8375) );
  INV_X1 U10825 ( .A(n8372), .ZN(n8373) );
  NAND2_X1 U10826 ( .A1(n8373), .A2(SI_11_), .ZN(n8374) );
  NAND2_X1 U10827 ( .A1(n8375), .A2(n8374), .ZN(n8696) );
  MUX2_X1 U10828 ( .A(n10074), .B(n10076), .S(n9479), .Z(n8376) );
  NAND2_X1 U10829 ( .A1(n8376), .A2(n9862), .ZN(n8379) );
  INV_X1 U10830 ( .A(n8376), .ZN(n8377) );
  NAND2_X1 U10831 ( .A1(n8377), .A2(SI_12_), .ZN(n8378) );
  MUX2_X1 U10832 ( .A(n10123), .B(n10125), .S(n9833), .Z(n8380) );
  NAND2_X1 U10833 ( .A1(n8380), .A2(n14377), .ZN(n8383) );
  INV_X1 U10834 ( .A(n8380), .ZN(n8381) );
  NAND2_X1 U10835 ( .A1(n8381), .A2(SI_13_), .ZN(n8382) );
  MUX2_X1 U10836 ( .A(n10338), .B(n10339), .S(n9833), .Z(n8388) );
  MUX2_X1 U10837 ( .A(n10390), .B(n10405), .S(n9479), .Z(n8385) );
  NAND2_X1 U10838 ( .A1(n8385), .A2(n8384), .ZN(n8390) );
  INV_X1 U10839 ( .A(n8385), .ZN(n8386) );
  NAND2_X1 U10840 ( .A1(n8386), .A2(SI_15_), .ZN(n8387) );
  NAND2_X1 U10841 ( .A1(n8390), .A2(n8387), .ZN(n8822) );
  NOR2_X1 U10842 ( .A1(n8388), .A2(n9889), .ZN(n8389) );
  MUX2_X1 U10843 ( .A(n10312), .B(n10335), .S(n9833), .Z(n8391) );
  NAND2_X1 U10844 ( .A1(n8391), .A2(n10070), .ZN(n8394) );
  INV_X1 U10845 ( .A(n8391), .ZN(n8392) );
  NAND2_X1 U10846 ( .A1(n8392), .A2(SI_16_), .ZN(n8393) );
  MUX2_X1 U10847 ( .A(n10388), .B(n10396), .S(n9479), .Z(n8778) );
  INV_X1 U10848 ( .A(n8778), .ZN(n8395) );
  NAND2_X1 U10849 ( .A1(n8395), .A2(SI_17_), .ZN(n8396) );
  NAND2_X1 U10850 ( .A1(n8780), .A2(n8396), .ZN(n8398) );
  NAND2_X1 U10851 ( .A1(n8778), .A2(n10078), .ZN(n8397) );
  MUX2_X1 U10852 ( .A(n10554), .B(n10565), .S(n9833), .Z(n8855) );
  MUX2_X1 U10853 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9479), .Z(n8400) );
  NAND2_X1 U10854 ( .A1(n8401), .A2(n10424), .ZN(n8402) );
  INV_X1 U10855 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11588) );
  MUX2_X1 U10856 ( .A(n11014), .B(n11588), .S(n9479), .Z(n8893) );
  MUX2_X1 U10857 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9833), .Z(n8404) );
  OAI21_X1 U10858 ( .B1(SI_21_), .B2(n8404), .A(n8406), .ZN(n8405) );
  INV_X1 U10859 ( .A(n8405), .ZN(n8912) );
  INV_X1 U10860 ( .A(n8408), .ZN(n8407) );
  INV_X1 U10861 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8409) );
  MUX2_X1 U10862 ( .A(n8409), .B(n11494), .S(n9479), .Z(n8936) );
  MUX2_X1 U10863 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9833), .Z(n8953) );
  NAND2_X1 U10864 ( .A1(n8412), .A2(n15242), .ZN(n8413) );
  MUX2_X1 U10865 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9833), .Z(n8979) );
  MUX2_X1 U10866 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9833), .Z(n8415) );
  XNOR2_X1 U10867 ( .A(n8415), .B(SI_25_), .ZN(n8998) );
  MUX2_X1 U10868 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n9479), .Z(n8416) );
  NAND2_X1 U10869 ( .A1(n8416), .A2(SI_26_), .ZN(n9018) );
  OAI21_X1 U10870 ( .B1(SI_26_), .B2(n8416), .A(n9018), .ZN(n8417) );
  NAND2_X1 U10871 ( .A1(n8418), .A2(n8417), .ZN(n8419) );
  NAND2_X1 U10872 ( .A1(n9019), .A2(n8419), .ZN(n14349) );
  NOR2_X1 U10873 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n8423) );
  NOR2_X1 U10874 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8422) );
  NOR2_X1 U10875 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8421) );
  NAND2_X2 U10876 ( .A1(n9159), .A2(n13579), .ZN(n8493) );
  OR2_X1 U10877 ( .A1(n6442), .A2(n13582), .ZN(n8429) );
  INV_X1 U10878 ( .A(n8443), .ZN(n8435) );
  INV_X1 U10879 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U10880 ( .A1(n8443), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8439) );
  XNOR2_X1 U10881 ( .A(n9147), .B(n9146), .ZN(n9157) );
  NAND2_X1 U10882 ( .A1(n9158), .A2(n9157), .ZN(n9797) );
  NAND2_X1 U10883 ( .A1(n8441), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10884 ( .A1(n7351), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10885 ( .A1(n11586), .A2(n13188), .ZN(n9788) );
  NAND2_X1 U10886 ( .A1(n8449), .A2(n9788), .ZN(n8446) );
  NAND2_X1 U10887 ( .A1(n9797), .A2(n8446), .ZN(n8448) );
  NAND2_X1 U10888 ( .A1(n11586), .A2(n10655), .ZN(n9124) );
  NAND2_X1 U10889 ( .A1(n9167), .A2(n14880), .ZN(n8447) );
  NAND2_X1 U10890 ( .A1(n8448), .A2(n8447), .ZN(n9109) );
  INV_X1 U10891 ( .A(n8728), .ZN(n8887) );
  NAND2_X1 U10892 ( .A1(n13477), .A2(n8728), .ZN(n8476) );
  NAND2_X1 U10893 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8574) );
  INV_X1 U10894 ( .A(n8574), .ZN(n8450) );
  NAND2_X1 U10895 ( .A1(n8450), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8598) );
  INV_X1 U10896 ( .A(n8598), .ZN(n8451) );
  NAND2_X1 U10897 ( .A1(n8451), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8620) );
  INV_X1 U10898 ( .A(n8620), .ZN(n8452) );
  NAND2_X1 U10899 ( .A1(n8452), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8641) );
  INV_X1 U10900 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8640) );
  INV_X1 U10901 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8729) );
  INV_X1 U10902 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n13170) );
  INV_X1 U10903 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13024) );
  INV_X1 U10904 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13037) );
  INV_X1 U10905 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13019) );
  INV_X1 U10906 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9002) );
  INV_X1 U10907 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8459) );
  NAND2_X1 U10908 ( .A1(n9005), .A2(n8459), .ZN(n8460) );
  NAND2_X1 U10909 ( .A1(n9070), .A2(n8460), .ZN(n13069) );
  NOR2_X1 U10910 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .ZN(n8461) );
  INV_X1 U10911 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8470) );
  NAND2_X4 U10912 ( .A1(n8465), .A2(n8466), .ZN(n9025) );
  NAND2_X1 U10913 ( .A1(n9073), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8469) );
  INV_X4 U10914 ( .A(n8507), .ZN(n9074) );
  NAND2_X1 U10915 ( .A1(n9074), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8468) );
  OAI211_X1 U10916 ( .C1(n8470), .C2(n9025), .A(n8469), .B(n8468), .ZN(n8471)
         );
  INV_X1 U10917 ( .A(n8471), .ZN(n8472) );
  INV_X1 U10918 ( .A(n9122), .ZN(n8958) );
  NAND2_X1 U10919 ( .A1(n13259), .A2(n8958), .ZN(n8475) );
  NAND2_X1 U10920 ( .A1(n8476), .A2(n8475), .ZN(n9017) );
  INV_X1 U10921 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8477) );
  INV_X1 U10922 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9818) );
  OR2_X1 U10923 ( .A1(n8986), .A2(n9818), .ZN(n8480) );
  INV_X1 U10924 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8478) );
  OR2_X1 U10925 ( .A1(n8537), .A2(n8478), .ZN(n8479) );
  INV_X1 U10926 ( .A(n8483), .ZN(n8484) );
  NAND2_X1 U10927 ( .A1(n8485), .A2(n8484), .ZN(n8486) );
  NAND2_X1 U10928 ( .A1(n8487), .A2(n8486), .ZN(n9836) );
  INV_X1 U10929 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10930 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8488) );
  NAND2_X1 U10931 ( .A1(n9833), .A2(SI_0_), .ZN(n8492) );
  XNOR2_X1 U10932 ( .A(n8491), .B(n8492), .ZN(n13593) );
  MUX2_X1 U10933 ( .A(n7313), .B(n13593), .S(n8493), .Z(n14867) );
  INV_X1 U10934 ( .A(n14867), .ZN(n14879) );
  NAND2_X1 U10935 ( .A1(n9693), .A2(n10655), .ZN(n8494) );
  AND2_X1 U10936 ( .A1(n8494), .A2(n8474), .ZN(n8500) );
  AOI21_X1 U10937 ( .B1(n14879), .B2(n9122), .A(n8500), .ZN(n8503) );
  INV_X1 U10938 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U10939 ( .A1(n9074), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8498) );
  INV_X1 U10940 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8495) );
  OR2_X1 U10941 ( .A1(n8537), .A2(n14960), .ZN(n8496) );
  NAND2_X1 U10942 ( .A1(n14879), .A2(n8500), .ZN(n8501) );
  OAI211_X1 U10943 ( .C1(n8503), .C2(n13118), .A(n8502), .B(n8501), .ZN(n8526)
         );
  NAND2_X1 U10944 ( .A1(n8728), .A2(n10297), .ZN(n8504) );
  NAND2_X1 U10945 ( .A1(n8505), .A2(n8504), .ZN(n8506) );
  OAI21_X1 U10946 ( .B1(n8527), .B2(n8526), .A(n8506), .ZN(n8530) );
  NAND2_X1 U10947 ( .A1(n8767), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8512) );
  INV_X1 U10948 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10995) );
  OR2_X1 U10949 ( .A1(n8986), .A2(n10995), .ZN(n8511) );
  INV_X1 U10950 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8508) );
  OR2_X1 U10951 ( .A1(n8507), .A2(n8508), .ZN(n8510) );
  INV_X1 U10952 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10082) );
  OR2_X1 U10953 ( .A1(n8537), .A2(n10082), .ZN(n8509) );
  NAND2_X1 U10954 ( .A1(n13115), .A2(n6436), .ZN(n8525) );
  NAND2_X1 U10955 ( .A1(n8515), .A2(n8514), .ZN(n8517) );
  NAND2_X1 U10956 ( .A1(n8517), .A2(n8516), .ZN(n9838) );
  OR2_X1 U10957 ( .A1(n8518), .A2(n9838), .ZN(n8523) );
  INV_X1 U10958 ( .A(n8519), .ZN(n8520) );
  NAND2_X1 U10959 ( .A1(n8520), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8522) );
  XNOR2_X1 U10960 ( .A(n8522), .B(n8521), .ZN(n14766) );
  NAND2_X1 U10961 ( .A1(n8728), .A2(n13048), .ZN(n8524) );
  NAND2_X1 U10962 ( .A1(n8525), .A2(n8524), .ZN(n8531) );
  NAND2_X1 U10963 ( .A1(n8531), .A2(n8532), .ZN(n8529) );
  NAND2_X1 U10964 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  NAND3_X1 U10965 ( .A1(n8530), .A2(n8529), .A3(n8528), .ZN(n8536) );
  INV_X1 U10966 ( .A(n8531), .ZN(n8534) );
  INV_X1 U10967 ( .A(n8532), .ZN(n8533) );
  NAND2_X1 U10968 ( .A1(n8534), .A2(n8533), .ZN(n8535) );
  NAND2_X1 U10969 ( .A1(n8536), .A2(n8535), .ZN(n8550) );
  NAND2_X1 U10970 ( .A1(n9074), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n10294) );
  OR2_X1 U10971 ( .A1(n8986), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10293) );
  INV_X1 U10972 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10669) );
  OR2_X1 U10973 ( .A1(n9025), .A2(n10669), .ZN(n10292) );
  INV_X1 U10974 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10084) );
  OR2_X1 U10975 ( .A1(n8537), .A2(n10084), .ZN(n10291) );
  NAND4_X1 U10976 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n13114) );
  NAND2_X1 U10977 ( .A1(n13114), .A2(n8728), .ZN(n8547) );
  NAND2_X1 U10978 ( .A1(n8538), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8539) );
  XNOR2_X1 U10979 ( .A(n8539), .B(n7312), .ZN(n14775) );
  OR2_X1 U10980 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U10981 ( .A1(n8543), .A2(n8542), .ZN(n9834) );
  OR2_X1 U10982 ( .A1(n6442), .A2(n9825), .ZN(n8544) );
  NAND2_X1 U10983 ( .A1(n10819), .A2(n6436), .ZN(n8546) );
  NAND2_X1 U10984 ( .A1(n8547), .A2(n8546), .ZN(n8549) );
  AOI22_X1 U10985 ( .A1(n13114), .A2(n6436), .B1(n10819), .B2(n8728), .ZN(
        n8548) );
  AOI21_X1 U10986 ( .B1(n8550), .B2(n8549), .A(n8548), .ZN(n8552) );
  NOR2_X1 U10987 ( .A1(n8550), .A2(n8549), .ZN(n8551) );
  NAND2_X1 U10988 ( .A1(n9073), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8557) );
  INV_X1 U10989 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8553) );
  OR2_X1 U10990 ( .A1(n8507), .A2(n8553), .ZN(n8556) );
  OAI21_X1 U10991 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8574), .ZN(n10846) );
  OR2_X1 U10992 ( .A1(n8986), .A2(n10846), .ZN(n8555) );
  INV_X1 U10993 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10841) );
  OR2_X1 U10994 ( .A1(n9025), .A2(n10841), .ZN(n8554) );
  NAND2_X1 U10995 ( .A1(n13113), .A2(n8958), .ZN(n8569) );
  OR2_X1 U10996 ( .A1(n8559), .A2(n8558), .ZN(n8560) );
  NAND2_X1 U10997 ( .A1(n8561), .A2(n8560), .ZN(n9844) );
  NOR2_X1 U10998 ( .A1(n9844), .A2(n8518), .ZN(n8567) );
  NAND2_X1 U10999 ( .A1(n8562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8563) );
  MUX2_X1 U11000 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8563), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8565) );
  INV_X1 U11001 ( .A(n8564), .ZN(n8583) );
  NAND2_X1 U11002 ( .A1(n8565), .A2(n8583), .ZN(n14793) );
  OAI22_X1 U11003 ( .A1(n6442), .A2(n9828), .B1(n8493), .B2(n14793), .ZN(n8566) );
  NAND2_X1 U11004 ( .A1(n8728), .A2(n10845), .ZN(n8568) );
  NAND2_X1 U11005 ( .A1(n8569), .A2(n8568), .ZN(n8571) );
  AOI22_X1 U11006 ( .A1(n13113), .A2(n8728), .B1(n6436), .B2(n10845), .ZN(
        n8570) );
  NAND2_X1 U11007 ( .A1(n9074), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8579) );
  INV_X1 U11008 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10087) );
  OR2_X1 U11009 ( .A1(n8537), .A2(n10087), .ZN(n8578) );
  INV_X1 U11010 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11011 ( .A1(n8574), .A2(n8573), .ZN(n8575) );
  NAND2_X1 U11012 ( .A1(n8598), .A2(n8575), .ZN(n10831) );
  OR2_X1 U11013 ( .A1(n8986), .A2(n10831), .ZN(n8577) );
  INV_X1 U11014 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10829) );
  OR2_X1 U11015 ( .A1(n9025), .A2(n10829), .ZN(n8576) );
  NAND4_X1 U11016 ( .A1(n8579), .A2(n8578), .A3(n8577), .A4(n8576), .ZN(n13112) );
  NAND2_X1 U11017 ( .A1(n13112), .A2(n8728), .ZN(n8588) );
  OR2_X1 U11018 ( .A1(n8580), .A2(n6726), .ZN(n8581) );
  NAND2_X1 U11019 ( .A1(n8582), .A2(n8581), .ZN(n9841) );
  OR2_X1 U11020 ( .A1(n9841), .A2(n8518), .ZN(n8586) );
  INV_X2 U11021 ( .A(n6442), .ZN(n8879) );
  NAND2_X1 U11022 ( .A1(n8583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8584) );
  XNOR2_X1 U11023 ( .A(n8584), .B(P2_IR_REG_5__SCAN_IN), .ZN(n14808) );
  AOI22_X1 U11024 ( .A1(n8879), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9795), .B2(
        n14808), .ZN(n8585) );
  NAND2_X1 U11025 ( .A1(n8586), .A2(n8585), .ZN(n14931) );
  INV_X1 U11026 ( .A(n9122), .ZN(n9081) );
  NAND2_X1 U11027 ( .A1(n14931), .A2(n9081), .ZN(n8587) );
  AOI22_X1 U11028 ( .A1(n8958), .A2(n13112), .B1(n14931), .B2(n8728), .ZN(
        n8589) );
  INV_X1 U11029 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8593) );
  AND2_X1 U11030 ( .A1(n8564), .A2(n8593), .ZN(n8782) );
  INV_X1 U11031 ( .A(n8782), .ZN(n8594) );
  NAND2_X1 U11032 ( .A1(n8594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8595) );
  XNOR2_X1 U11033 ( .A(n8595), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U11034 ( .A1(n8879), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9795), .B2(
        n13124), .ZN(n8596) );
  NAND2_X1 U11035 ( .A1(n9073), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U11036 ( .A1(n9074), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8602) );
  INV_X1 U11037 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11038 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U11039 ( .A1(n8620), .A2(n8599), .ZN(n10963) );
  OR2_X1 U11040 ( .A1(n8986), .A2(n10963), .ZN(n8601) );
  INV_X1 U11041 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10102) );
  OR2_X1 U11042 ( .A1(n9025), .A2(n10102), .ZN(n8600) );
  NAND4_X1 U11043 ( .A1(n8603), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n13111) );
  AOI22_X1 U11044 ( .A1(n10965), .A2(n8728), .B1(n6436), .B2(n13111), .ZN(
        n8610) );
  INV_X1 U11045 ( .A(n8610), .ZN(n8604) );
  NAND2_X1 U11046 ( .A1(n8609), .A2(n8604), .ZN(n8608) );
  NAND2_X1 U11047 ( .A1(n10965), .A2(n8958), .ZN(n8606) );
  NAND2_X1 U11048 ( .A1(n13111), .A2(n8728), .ZN(n8605) );
  NAND2_X1 U11049 ( .A1(n8606), .A2(n8605), .ZN(n8607) );
  NAND2_X1 U11050 ( .A1(n9868), .A2(n9100), .ZN(n8617) );
  INV_X1 U11051 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U11052 ( .A1(n8782), .A2(n8614), .ZN(n8633) );
  NAND2_X1 U11053 ( .A1(n8633), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8615) );
  XNOR2_X1 U11054 ( .A(n8615), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U11055 ( .A1(n8879), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9795), .B2(
        n13136), .ZN(n8616) );
  NAND2_X1 U11056 ( .A1(n10942), .A2(n8958), .ZN(n8627) );
  NAND2_X1 U11057 ( .A1(n9073), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8625) );
  INV_X1 U11058 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8618) );
  OR2_X1 U11059 ( .A1(n8507), .A2(n8618), .ZN(n8624) );
  INV_X1 U11060 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U11061 ( .A1(n8620), .A2(n8619), .ZN(n8621) );
  NAND2_X1 U11062 ( .A1(n8641), .A2(n8621), .ZN(n14852) );
  OR2_X1 U11063 ( .A1(n8986), .A2(n14852), .ZN(n8623) );
  INV_X1 U11064 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10105) );
  OR2_X1 U11065 ( .A1(n9025), .A2(n10105), .ZN(n8622) );
  NAND4_X1 U11066 ( .A1(n8625), .A2(n8624), .A3(n8623), .A4(n8622), .ZN(n13110) );
  NAND2_X1 U11067 ( .A1(n13110), .A2(n8728), .ZN(n8626) );
  NAND2_X1 U11068 ( .A1(n8627), .A2(n8626), .ZN(n8629) );
  AOI22_X1 U11069 ( .A1(n10942), .A2(n8728), .B1(n6436), .B2(n13110), .ZN(
        n8628) );
  XNOR2_X1 U11070 ( .A(n8630), .B(SI_8_), .ZN(n8631) );
  NAND2_X1 U11071 ( .A1(n9873), .A2(n9100), .ZN(n8638) );
  NAND2_X1 U11072 ( .A1(n8635), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8634) );
  MUX2_X1 U11073 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8634), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8636) );
  NAND2_X1 U11074 ( .A1(n8636), .A2(n8676), .ZN(n10109) );
  INV_X1 U11075 ( .A(n10109), .ZN(n14822) );
  AOI22_X1 U11076 ( .A1(n8879), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9795), .B2(
        n14822), .ZN(n8637) );
  NAND2_X1 U11077 ( .A1(n11109), .A2(n8728), .ZN(n8648) );
  NAND2_X1 U11078 ( .A1(n9073), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8646) );
  INV_X1 U11079 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8639) );
  OR2_X1 U11080 ( .A1(n8507), .A2(n8639), .ZN(n8645) );
  NAND2_X1 U11081 ( .A1(n8641), .A2(n8640), .ZN(n8642) );
  NAND2_X1 U11082 ( .A1(n8665), .A2(n8642), .ZN(n10950) );
  OR2_X1 U11083 ( .A1(n8986), .A2(n10950), .ZN(n8644) );
  INV_X1 U11084 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10951) );
  OR2_X1 U11085 ( .A1(n9025), .A2(n10951), .ZN(n8643) );
  NAND4_X1 U11086 ( .A1(n8646), .A2(n8645), .A3(n8644), .A4(n8643), .ZN(n13109) );
  NAND2_X1 U11087 ( .A1(n13109), .A2(n9081), .ZN(n8647) );
  NAND2_X1 U11088 ( .A1(n8648), .A2(n8647), .ZN(n8653) );
  NAND2_X1 U11089 ( .A1(n8652), .A2(n8653), .ZN(n8651) );
  INV_X1 U11090 ( .A(n13109), .ZN(n11146) );
  NAND2_X1 U11091 ( .A1(n11109), .A2(n9081), .ZN(n8649) );
  OAI21_X1 U11092 ( .B1(n11146), .B2(n8887), .A(n8649), .ZN(n8650) );
  NAND2_X1 U11093 ( .A1(n8651), .A2(n8650), .ZN(n8657) );
  INV_X1 U11094 ( .A(n8652), .ZN(n8655) );
  INV_X1 U11095 ( .A(n8653), .ZN(n8654) );
  NAND2_X1 U11096 ( .A1(n8655), .A2(n8654), .ZN(n8656) );
  XNOR2_X1 U11097 ( .A(n8659), .B(n8658), .ZN(n9884) );
  NAND2_X1 U11098 ( .A1(n9884), .A2(n9100), .ZN(n8662) );
  NAND2_X1 U11099 ( .A1(n8676), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8660) );
  XNOR2_X1 U11100 ( .A(n8660), .B(P2_IR_REG_9__SCAN_IN), .ZN(n14839) );
  AOI22_X1 U11101 ( .A1(n8879), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9795), .B2(
        n14839), .ZN(n8661) );
  NAND2_X1 U11102 ( .A1(n11232), .A2(n9081), .ZN(n8672) );
  NAND2_X1 U11103 ( .A1(n9074), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8670) );
  INV_X1 U11104 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8663) );
  OR2_X1 U11105 ( .A1(n8537), .A2(n8663), .ZN(n8669) );
  INV_X1 U11106 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U11107 ( .A1(n8665), .A2(n8664), .ZN(n8666) );
  NAND2_X1 U11108 ( .A1(n8684), .A2(n8666), .ZN(n11142) );
  OR2_X1 U11109 ( .A1(n8986), .A2(n11142), .ZN(n8668) );
  INV_X1 U11110 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10111) );
  OR2_X1 U11111 ( .A1(n9025), .A2(n10111), .ZN(n8667) );
  NAND4_X1 U11112 ( .A1(n8670), .A2(n8669), .A3(n8668), .A4(n8667), .ZN(n13108) );
  NAND2_X1 U11113 ( .A1(n13108), .A2(n8728), .ZN(n8671) );
  AOI22_X1 U11114 ( .A1(n11232), .A2(n8728), .B1(n8958), .B2(n13108), .ZN(
        n8673) );
  XNOR2_X1 U11115 ( .A(n8674), .B(n8675), .ZN(n9922) );
  NAND2_X1 U11116 ( .A1(n9922), .A2(n9100), .ZN(n8681) );
  INV_X1 U11117 ( .A(n8676), .ZN(n8678) );
  INV_X1 U11118 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U11119 ( .A1(n8678), .A2(n8677), .ZN(n8698) );
  NAND2_X1 U11120 ( .A1(n8698), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8679) );
  XNOR2_X1 U11121 ( .A(n8679), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U11122 ( .A1(n8879), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9795), 
        .B2(n10134), .ZN(n8680) );
  NAND2_X1 U11123 ( .A1(n11380), .A2(n8728), .ZN(n8691) );
  NAND2_X1 U11124 ( .A1(n9073), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8689) );
  INV_X1 U11125 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8682) );
  OR2_X1 U11126 ( .A1(n8507), .A2(n8682), .ZN(n8688) );
  NAND2_X1 U11127 ( .A1(n8684), .A2(n8683), .ZN(n8685) );
  NAND2_X1 U11128 ( .A1(n8704), .A2(n8685), .ZN(n11187) );
  OR2_X1 U11129 ( .A1(n8986), .A2(n11187), .ZN(n8687) );
  INV_X1 U11130 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11162) );
  OR2_X1 U11131 ( .A1(n9025), .A2(n11162), .ZN(n8686) );
  NAND4_X1 U11132 ( .A1(n8689), .A2(n8688), .A3(n8687), .A4(n8686), .ZN(n13107) );
  NAND2_X1 U11133 ( .A1(n13107), .A2(n6436), .ZN(n8690) );
  NAND2_X1 U11134 ( .A1(n8691), .A2(n8690), .ZN(n8694) );
  INV_X1 U11135 ( .A(n13107), .ZN(n11397) );
  NAND2_X1 U11136 ( .A1(n11380), .A2(n8958), .ZN(n8692) );
  OAI21_X1 U11137 ( .B1(n11397), .B2(n8887), .A(n8692), .ZN(n8693) );
  XNOR2_X1 U11138 ( .A(n8697), .B(n8696), .ZN(n10002) );
  NAND2_X1 U11139 ( .A1(n10002), .A2(n9100), .ZN(n8701) );
  OAI21_X1 U11140 ( .B1(n8698), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8699) );
  XNOR2_X1 U11141 ( .A(n8699), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U11142 ( .A1(n8879), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9795), 
        .B2(n10211), .ZN(n8700) );
  NAND2_X1 U11143 ( .A1(n13549), .A2(n8958), .ZN(n8711) );
  NAND2_X1 U11144 ( .A1(n9073), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8709) );
  INV_X1 U11145 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8702) );
  OR2_X1 U11146 ( .A1(n8507), .A2(n8702), .ZN(n8708) );
  INV_X1 U11147 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U11148 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  NAND2_X1 U11149 ( .A1(n8730), .A2(n8705), .ZN(n11395) );
  OR2_X1 U11150 ( .A1(n8986), .A2(n11395), .ZN(n8707) );
  INV_X1 U11151 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11388) );
  OR2_X1 U11152 ( .A1(n9025), .A2(n11388), .ZN(n8706) );
  NAND4_X1 U11153 ( .A1(n8709), .A2(n8708), .A3(n8707), .A4(n8706), .ZN(n13106) );
  NAND2_X1 U11154 ( .A1(n13106), .A2(n8728), .ZN(n8710) );
  NAND2_X1 U11155 ( .A1(n8711), .A2(n8710), .ZN(n8713) );
  AOI22_X1 U11156 ( .A1(n13549), .A2(n8728), .B1(n6436), .B2(n13106), .ZN(
        n8712) );
  AOI21_X1 U11157 ( .B1(n8714), .B2(n8713), .A(n8712), .ZN(n8716) );
  OR2_X1 U11158 ( .A1(n8716), .A2(n8715), .ZN(n8740) );
  OR2_X1 U11159 ( .A1(n8719), .A2(n8718), .ZN(n8720) );
  NAND2_X1 U11160 ( .A1(n8717), .A2(n8720), .ZN(n10072) );
  NAND2_X1 U11161 ( .A1(n10072), .A2(n9100), .ZN(n8727) );
  NAND2_X1 U11162 ( .A1(n8782), .A2(n8722), .ZN(n8724) );
  NAND2_X1 U11163 ( .A1(n8724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8723) );
  MUX2_X1 U11164 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8723), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8725) );
  AND2_X1 U11165 ( .A1(n8725), .A2(n8746), .ZN(n10408) );
  AOI22_X1 U11166 ( .A1(n8879), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9795), 
        .B2(n10408), .ZN(n8726) );
  NAND2_X1 U11167 ( .A1(n12092), .A2(n8728), .ZN(n8737) );
  NAND2_X1 U11168 ( .A1(n9074), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8735) );
  INV_X1 U11169 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11464) );
  OR2_X1 U11170 ( .A1(n9025), .A2(n11464), .ZN(n8734) );
  NAND2_X1 U11171 ( .A1(n8730), .A2(n8729), .ZN(n8731) );
  NAND2_X1 U11172 ( .A1(n8751), .A2(n8731), .ZN(n11463) );
  OR2_X1 U11173 ( .A1(n8986), .A2(n11463), .ZN(n8733) );
  INV_X1 U11174 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10206) );
  OR2_X1 U11175 ( .A1(n8537), .A2(n10206), .ZN(n8732) );
  NAND4_X1 U11176 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n13445) );
  NAND2_X1 U11177 ( .A1(n13445), .A2(n8958), .ZN(n8736) );
  NAND2_X1 U11178 ( .A1(n8737), .A2(n8736), .ZN(n8739) );
  AOI22_X1 U11179 ( .A1(n12092), .A2(n8958), .B1(n13445), .B2(n8728), .ZN(
        n8738) );
  OR2_X1 U11180 ( .A1(n8742), .A2(n8741), .ZN(n8743) );
  NAND2_X1 U11181 ( .A1(n8744), .A2(n8743), .ZN(n10122) );
  NAND2_X1 U11182 ( .A1(n10122), .A2(n9100), .ZN(n8749) );
  NAND2_X1 U11183 ( .A1(n8746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8745) );
  MUX2_X1 U11184 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8745), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8747) );
  NAND2_X1 U11185 ( .A1(n8747), .A2(n8825), .ZN(n10414) );
  INV_X1 U11186 ( .A(n10414), .ZN(n10631) );
  AOI22_X1 U11187 ( .A1(n8879), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9795), 
        .B2(n10631), .ZN(n8748) );
  NAND2_X1 U11188 ( .A1(n13543), .A2(n8958), .ZN(n8758) );
  NAND2_X1 U11189 ( .A1(n9074), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11190 ( .A1(n8751), .A2(n8750), .ZN(n8752) );
  NAND2_X1 U11191 ( .A1(n8769), .A2(n8752), .ZN(n13448) );
  OR2_X1 U11192 ( .A1(n8986), .A2(n13448), .ZN(n8755) );
  INV_X1 U11193 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10415) );
  OR2_X1 U11194 ( .A1(n9025), .A2(n10415), .ZN(n8754) );
  INV_X1 U11195 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10406) );
  OR2_X1 U11196 ( .A1(n8537), .A2(n10406), .ZN(n8753) );
  NAND4_X1 U11197 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), .ZN(n13105) );
  NAND2_X1 U11198 ( .A1(n13105), .A2(n8728), .ZN(n8757) );
  NAND2_X1 U11199 ( .A1(n8758), .A2(n8757), .ZN(n8761) );
  NAND2_X1 U11200 ( .A1(n13543), .A2(n8728), .ZN(n8759) );
  OAI21_X1 U11201 ( .B1(n13421), .B2(n9122), .A(n8759), .ZN(n8760) );
  NAND2_X1 U11202 ( .A1(n8762), .A2(n9889), .ZN(n8819) );
  NAND2_X1 U11203 ( .A1(n10337), .A2(n9100), .ZN(n8766) );
  NAND2_X1 U11204 ( .A1(n8825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8764) );
  XNOR2_X1 U11205 ( .A(n8764), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U11206 ( .A1(n8879), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9795), 
        .B2(n11204), .ZN(n8765) );
  NAND2_X1 U11207 ( .A1(n13434), .A2(n8728), .ZN(n8776) );
  NAND2_X1 U11208 ( .A1(n9074), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8774) );
  INV_X1 U11209 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n13431) );
  OR2_X1 U11210 ( .A1(n9025), .A2(n13431), .ZN(n8773) );
  INV_X1 U11211 ( .A(n8768), .ZN(n8830) );
  NAND2_X1 U11212 ( .A1(n8769), .A2(n15198), .ZN(n8770) );
  NAND2_X1 U11213 ( .A1(n8830), .A2(n8770), .ZN(n13430) );
  OR2_X1 U11214 ( .A1(n8986), .A2(n13430), .ZN(n8772) );
  INV_X1 U11215 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10628) );
  OR2_X1 U11216 ( .A1(n8537), .A2(n10628), .ZN(n8771) );
  NAND4_X1 U11217 ( .A1(n8774), .A2(n8773), .A3(n8772), .A4(n8771), .ZN(n13442) );
  NAND2_X1 U11218 ( .A1(n13442), .A2(n6436), .ZN(n8775) );
  NAND2_X1 U11219 ( .A1(n8776), .A2(n8775), .ZN(n8842) );
  AOI22_X1 U11220 ( .A1(n13434), .A2(n8958), .B1(n13442), .B2(n8728), .ZN(
        n8777) );
  AOI21_X1 U11221 ( .B1(n8843), .B2(n8842), .A(n8777), .ZN(n8854) );
  XNOR2_X1 U11222 ( .A(n8778), .B(SI_17_), .ZN(n8779) );
  XNOR2_X1 U11223 ( .A(n8780), .B(n8779), .ZN(n10387) );
  NAND2_X1 U11224 ( .A1(n10387), .A2(n9100), .ZN(n8787) );
  NAND2_X1 U11225 ( .A1(n8782), .A2(n8781), .ZN(n8799) );
  NAND2_X1 U11226 ( .A1(n8801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8783) );
  MUX2_X1 U11227 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8783), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8785) );
  NAND2_X1 U11228 ( .A1(n8785), .A2(n8784), .ZN(n13159) );
  AOI22_X1 U11229 ( .A1(n8879), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9795), 
        .B2(n13166), .ZN(n8786) );
  INV_X1 U11230 ( .A(n8788), .ZN(n8807) );
  INV_X1 U11231 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U11232 ( .A1(n8807), .A2(n8789), .ZN(n8790) );
  NAND2_X1 U11233 ( .A1(n8862), .A2(n8790), .ZN(n13379) );
  OR2_X1 U11234 ( .A1(n13379), .A2(n8986), .ZN(n8794) );
  NAND2_X1 U11235 ( .A1(n9073), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U11236 ( .A1(n9074), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U11237 ( .A1(n8767), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8791) );
  NAND4_X1 U11238 ( .A1(n8794), .A2(n8793), .A3(n8792), .A4(n8791), .ZN(n13102) );
  AOI22_X1 U11239 ( .A1(n13527), .A2(n8728), .B1(n8958), .B2(n13102), .ZN(
        n8797) );
  NAND2_X1 U11240 ( .A1(n13527), .A2(n9081), .ZN(n8796) );
  NAND2_X1 U11241 ( .A1(n13102), .A2(n8728), .ZN(n8795) );
  NAND2_X1 U11242 ( .A1(n8796), .A2(n8795), .ZN(n8848) );
  NAND2_X1 U11243 ( .A1(n8797), .A2(n8848), .ZN(n8818) );
  XNOR2_X1 U11244 ( .A(n8798), .B(n7651), .ZN(n10311) );
  NAND2_X1 U11245 ( .A1(n10311), .A2(n9100), .ZN(n8804) );
  NAND2_X1 U11246 ( .A1(n8799), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8800) );
  MUX2_X1 U11247 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8800), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8802) );
  AND2_X1 U11248 ( .A1(n8802), .A2(n8801), .ZN(n11434) );
  AOI22_X1 U11249 ( .A1(n8879), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9795), 
        .B2(n11434), .ZN(n8803) );
  INV_X1 U11250 ( .A(n8805), .ZN(n8832) );
  INV_X1 U11251 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U11252 ( .A1(n8832), .A2(n15197), .ZN(n8806) );
  NAND2_X1 U11253 ( .A1(n8807), .A2(n8806), .ZN(n13400) );
  OR2_X1 U11254 ( .A1(n13400), .A2(n8986), .ZN(n8813) );
  INV_X1 U11255 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8808) );
  OR2_X1 U11256 ( .A1(n8537), .A2(n8808), .ZN(n8812) );
  INV_X1 U11257 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8809) );
  OR2_X1 U11258 ( .A1(n8507), .A2(n8809), .ZN(n8811) );
  INV_X1 U11259 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13401) );
  OR2_X1 U11260 ( .A1(n9025), .A2(n13401), .ZN(n8810) );
  NAND4_X1 U11261 ( .A1(n8813), .A2(n8812), .A3(n8811), .A4(n8810), .ZN(n13103) );
  AND2_X1 U11262 ( .A1(n13103), .A2(n6436), .ZN(n8814) );
  AOI21_X1 U11263 ( .B1(n13533), .B2(n8728), .A(n8814), .ZN(n8845) );
  NAND2_X1 U11264 ( .A1(n13533), .A2(n9081), .ZN(n8816) );
  NAND2_X1 U11265 ( .A1(n13103), .A2(n8728), .ZN(n8815) );
  NAND2_X1 U11266 ( .A1(n8816), .A2(n8815), .ZN(n8844) );
  NAND2_X1 U11267 ( .A1(n8845), .A2(n8844), .ZN(n8817) );
  AND2_X1 U11268 ( .A1(n8818), .A2(n8817), .ZN(n8851) );
  INV_X1 U11269 ( .A(n8822), .ZN(n8823) );
  XNOR2_X1 U11270 ( .A(n8824), .B(n8823), .ZN(n10389) );
  NAND2_X1 U11271 ( .A1(n10389), .A2(n9100), .ZN(n8828) );
  OAI21_X1 U11272 ( .B1(n8825), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8826) );
  XNOR2_X1 U11273 ( .A(n8826), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U11274 ( .A1(n8879), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9795), 
        .B2(n11198), .ZN(n8827) );
  NAND2_X1 U11275 ( .A1(n9074), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8837) );
  INV_X1 U11276 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11206) );
  OR2_X1 U11277 ( .A1(n8537), .A2(n11206), .ZN(n8836) );
  INV_X1 U11278 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8829) );
  NAND2_X1 U11279 ( .A1(n8830), .A2(n8829), .ZN(n8831) );
  NAND2_X1 U11280 ( .A1(n8832), .A2(n8831), .ZN(n13412) );
  OR2_X1 U11281 ( .A1(n8986), .A2(n13412), .ZN(n8835) );
  INV_X1 U11282 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8833) );
  OR2_X1 U11283 ( .A1(n9025), .A2(n8833), .ZN(n8834) );
  NAND4_X1 U11284 ( .A1(n8837), .A2(n8836), .A3(n8835), .A4(n8834), .ZN(n13104) );
  AND2_X1 U11285 ( .A1(n13104), .A2(n6436), .ZN(n8838) );
  AOI21_X1 U11286 ( .B1(n13538), .B2(n8728), .A(n8838), .ZN(n8847) );
  NAND2_X1 U11287 ( .A1(n13538), .A2(n9081), .ZN(n8840) );
  NAND2_X1 U11288 ( .A1(n13104), .A2(n8728), .ZN(n8839) );
  NAND2_X1 U11289 ( .A1(n8840), .A2(n8839), .ZN(n8846) );
  NAND2_X1 U11290 ( .A1(n8847), .A2(n8846), .ZN(n8841) );
  OAI21_X1 U11291 ( .B1(n8843), .B2(n8842), .A(n7658), .ZN(n8853) );
  OAI22_X1 U11292 ( .A1(n8847), .A2(n8846), .B1(n8845), .B2(n8844), .ZN(n8850)
         );
  INV_X1 U11293 ( .A(n8848), .ZN(n8849) );
  OR2_X1 U11294 ( .A1(n13527), .A2(n13102), .ZN(n12102) );
  AOI22_X1 U11295 ( .A1(n8851), .A2(n8850), .B1(n8849), .B2(n12102), .ZN(n8852) );
  OAI21_X1 U11296 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(n8871) );
  NAND2_X1 U11297 ( .A1(n8856), .A2(n8855), .ZN(n8857) );
  NAND2_X1 U11298 ( .A1(n8858), .A2(n8857), .ZN(n10566) );
  OR2_X1 U11299 ( .A1(n10566), .A2(n8518), .ZN(n8861) );
  NAND2_X1 U11300 ( .A1(n8784), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8859) );
  XNOR2_X1 U11301 ( .A(n8859), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13162) );
  AOI22_X1 U11302 ( .A1(n8879), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9795), 
        .B2(n13162), .ZN(n8860) );
  NAND2_X1 U11303 ( .A1(n13522), .A2(n8728), .ZN(n8867) );
  NAND2_X1 U11304 ( .A1(n8862), .A2(n13170), .ZN(n8863) );
  NAND2_X1 U11305 ( .A1(n8883), .A2(n8863), .ZN(n13366) );
  AOI22_X1 U11306 ( .A1(n9073), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9074), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U11307 ( .A1(n8767), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8864) );
  OAI211_X1 U11308 ( .C1(n13366), .C2(n8986), .A(n8865), .B(n8864), .ZN(n13101) );
  NAND2_X1 U11309 ( .A1(n13101), .A2(n8958), .ZN(n8866) );
  NAND2_X1 U11310 ( .A1(n8867), .A2(n8866), .ZN(n8872) );
  NAND2_X1 U11311 ( .A1(n8871), .A2(n8872), .ZN(n8870) );
  AOI22_X1 U11312 ( .A1(n13522), .A2(n8958), .B1(n13101), .B2(n8728), .ZN(
        n8868) );
  NAND2_X1 U11313 ( .A1(n8870), .A2(n8869), .ZN(n8876) );
  INV_X1 U11314 ( .A(n8871), .ZN(n8874) );
  INV_X1 U11315 ( .A(n8872), .ZN(n8873) );
  NAND2_X1 U11316 ( .A1(n8874), .A2(n8873), .ZN(n8875) );
  XNOR2_X1 U11317 ( .A(n8878), .B(n8877), .ZN(n10850) );
  NAND2_X1 U11318 ( .A1(n10850), .A2(n9100), .ZN(n8881) );
  AOI22_X1 U11319 ( .A1(n8879), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10655), 
        .B2(n9795), .ZN(n8880) );
  NAND2_X1 U11320 ( .A1(n13516), .A2(n9081), .ZN(n8889) );
  INV_X1 U11321 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13355) );
  INV_X1 U11322 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U11323 ( .A1(n8883), .A2(n8882), .ZN(n8884) );
  NAND2_X1 U11324 ( .A1(n8899), .A2(n8884), .ZN(n13352) );
  OR2_X1 U11325 ( .A1(n13352), .A2(n8986), .ZN(n8886) );
  AOI22_X1 U11326 ( .A1(n9073), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9074), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n8885) );
  OAI211_X1 U11327 ( .C1(n9025), .C2(n13355), .A(n8886), .B(n8885), .ZN(n13100) );
  NAND2_X1 U11328 ( .A1(n13100), .A2(n8728), .ZN(n8888) );
  NAND2_X1 U11329 ( .A1(n8889), .A2(n8888), .ZN(n8892) );
  NAND2_X1 U11330 ( .A1(n13516), .A2(n8728), .ZN(n8891) );
  NAND2_X1 U11331 ( .A1(n13100), .A2(n9081), .ZN(n8890) );
  NAND2_X1 U11332 ( .A1(n8894), .A2(n8893), .ZN(n8895) );
  OR2_X1 U11333 ( .A1(n11587), .A2(n8518), .ZN(n8898) );
  OR2_X1 U11334 ( .A1(n6442), .A2(n11588), .ZN(n8897) );
  NAND2_X1 U11335 ( .A1(n13511), .A2(n8728), .ZN(n8908) );
  NAND2_X1 U11336 ( .A1(n8899), .A2(n13024), .ZN(n8900) );
  AND2_X1 U11337 ( .A1(n8918), .A2(n8900), .ZN(n13340) );
  NAND2_X1 U11338 ( .A1(n13340), .A2(n9043), .ZN(n8906) );
  INV_X1 U11339 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U11340 ( .A1(n9073), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U11341 ( .A1(n9074), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8901) );
  OAI211_X1 U11342 ( .C1(n8903), .C2(n9025), .A(n8902), .B(n8901), .ZN(n8904)
         );
  INV_X1 U11343 ( .A(n8904), .ZN(n8905) );
  NAND2_X1 U11344 ( .A1(n8906), .A2(n8905), .ZN(n13099) );
  NAND2_X1 U11345 ( .A1(n13099), .A2(n8958), .ZN(n8907) );
  NAND2_X1 U11346 ( .A1(n8908), .A2(n8907), .ZN(n8910) );
  AOI22_X1 U11347 ( .A1(n13511), .A2(n9081), .B1(n13099), .B2(n8728), .ZN(
        n8909) );
  OR2_X1 U11348 ( .A1(n8913), .A2(n8912), .ZN(n8914) );
  NAND2_X1 U11349 ( .A1(n8915), .A2(n8914), .ZN(n11138) );
  OR2_X1 U11350 ( .A1(n11138), .A2(n8518), .ZN(n8917) );
  OR2_X1 U11351 ( .A1(n6442), .A2(n11139), .ZN(n8916) );
  NAND2_X1 U11352 ( .A1(n13325), .A2(n6436), .ZN(n8926) );
  INV_X1 U11353 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12979) );
  NAND2_X1 U11354 ( .A1(n8918), .A2(n12979), .ZN(n8919) );
  NAND2_X1 U11355 ( .A1(n8940), .A2(n8919), .ZN(n13322) );
  OR2_X1 U11356 ( .A1(n13322), .A2(n8986), .ZN(n8924) );
  INV_X1 U11357 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13323) );
  NAND2_X1 U11358 ( .A1(n9074), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U11359 ( .A1(n9073), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8920) );
  OAI211_X1 U11360 ( .C1(n13323), .C2(n9025), .A(n8921), .B(n8920), .ZN(n8922)
         );
  INV_X1 U11361 ( .A(n8922), .ZN(n8923) );
  NAND2_X1 U11362 ( .A1(n8924), .A2(n8923), .ZN(n13300) );
  NAND2_X1 U11363 ( .A1(n13300), .A2(n8728), .ZN(n8925) );
  NAND2_X1 U11364 ( .A1(n8926), .A2(n8925), .ZN(n8931) );
  INV_X1 U11365 ( .A(n13300), .ZN(n13336) );
  NAND2_X1 U11366 ( .A1(n13325), .A2(n8728), .ZN(n8927) );
  OAI21_X1 U11367 ( .B1(n13336), .B2(n9122), .A(n8927), .ZN(n8928) );
  NAND2_X1 U11368 ( .A1(n8929), .A2(n8928), .ZN(n8935) );
  INV_X1 U11369 ( .A(n8930), .ZN(n8933) );
  NAND2_X1 U11370 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  NAND2_X1 U11371 ( .A1(n8935), .A2(n8934), .ZN(n8952) );
  OR2_X1 U11372 ( .A1(n6442), .A2(n11494), .ZN(n8938) );
  NAND2_X1 U11373 ( .A1(n13498), .A2(n8728), .ZN(n8949) );
  NAND2_X1 U11374 ( .A1(n8940), .A2(n13037), .ZN(n8941) );
  AND2_X1 U11375 ( .A1(n8960), .A2(n8941), .ZN(n13306) );
  NAND2_X1 U11376 ( .A1(n13306), .A2(n9043), .ZN(n8947) );
  INV_X1 U11377 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U11378 ( .A1(n9073), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8943) );
  NAND2_X1 U11379 ( .A1(n9074), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8942) );
  OAI211_X1 U11380 ( .C1(n8944), .C2(n9025), .A(n8943), .B(n8942), .ZN(n8945)
         );
  INV_X1 U11381 ( .A(n8945), .ZN(n8946) );
  NAND2_X1 U11382 ( .A1(n13098), .A2(n6436), .ZN(n8948) );
  NAND2_X1 U11383 ( .A1(n8949), .A2(n8948), .ZN(n8951) );
  AOI22_X1 U11384 ( .A1(n13498), .A2(n8958), .B1(n13098), .B2(n8728), .ZN(
        n8950) );
  XNOR2_X1 U11385 ( .A(n8953), .B(SI_23_), .ZN(n8954) );
  XNOR2_X1 U11386 ( .A(n8955), .B(n8954), .ZN(n11507) );
  NAND2_X1 U11387 ( .A1(n11507), .A2(n9100), .ZN(n8957) );
  OR2_X1 U11388 ( .A1(n6442), .A2(n11510), .ZN(n8956) );
  NAND2_X1 U11389 ( .A1(n13492), .A2(n8958), .ZN(n8968) );
  INV_X1 U11390 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U11391 ( .A1(n8960), .A2(n8959), .ZN(n8961) );
  NAND2_X1 U11392 ( .A1(n8984), .A2(n8961), .ZN(n12943) );
  OR2_X1 U11393 ( .A1(n12943), .A2(n8986), .ZN(n8966) );
  INV_X1 U11394 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n15283) );
  NAND2_X1 U11395 ( .A1(n9073), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U11396 ( .A1(n8767), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8962) );
  OAI211_X1 U11397 ( .C1(n8507), .C2(n15283), .A(n8963), .B(n8962), .ZN(n8964)
         );
  INV_X1 U11398 ( .A(n8964), .ZN(n8965) );
  NAND2_X1 U11399 ( .A1(n13301), .A2(n8728), .ZN(n8967) );
  NAND2_X1 U11400 ( .A1(n8968), .A2(n8967), .ZN(n8973) );
  NAND2_X1 U11401 ( .A1(n13492), .A2(n8728), .ZN(n8969) );
  OAI21_X1 U11402 ( .B1(n13040), .B2(n9122), .A(n8969), .ZN(n8970) );
  NAND2_X1 U11403 ( .A1(n8971), .A2(n8970), .ZN(n8977) );
  INV_X1 U11404 ( .A(n8972), .ZN(n8975) );
  INV_X1 U11405 ( .A(n8973), .ZN(n8974) );
  NAND2_X1 U11406 ( .A1(n8975), .A2(n8974), .ZN(n8976) );
  NAND2_X1 U11407 ( .A1(n8977), .A2(n8976), .ZN(n8997) );
  NAND2_X1 U11408 ( .A1(n7486), .A2(n7485), .ZN(n8981) );
  NAND2_X1 U11409 ( .A1(n13587), .A2(n9100), .ZN(n8983) );
  OR2_X1 U11410 ( .A1(n6442), .A2(n13589), .ZN(n8982) );
  NAND2_X1 U11411 ( .A1(n13487), .A2(n8728), .ZN(n8994) );
  NAND2_X1 U11412 ( .A1(n8984), .A2(n13019), .ZN(n8985) );
  NAND2_X1 U11413 ( .A1(n9003), .A2(n8985), .ZN(n13275) );
  OR2_X1 U11414 ( .A1(n13275), .A2(n8986), .ZN(n8992) );
  INV_X1 U11415 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8989) );
  NAND2_X1 U11416 ( .A1(n9073), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U11417 ( .A1(n9074), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8987) );
  OAI211_X1 U11418 ( .C1(n8989), .C2(n9025), .A(n8988), .B(n8987), .ZN(n8990)
         );
  INV_X1 U11419 ( .A(n8990), .ZN(n8991) );
  NAND2_X1 U11420 ( .A1(n13258), .A2(n9081), .ZN(n8993) );
  NAND2_X1 U11421 ( .A1(n8994), .A2(n8993), .ZN(n8996) );
  AOI22_X1 U11422 ( .A1(n13487), .A2(n9081), .B1(n13258), .B2(n8728), .ZN(
        n8995) );
  XNOR2_X1 U11423 ( .A(n8999), .B(n8998), .ZN(n13584) );
  NAND2_X1 U11424 ( .A1(n13584), .A2(n9100), .ZN(n9001) );
  OR2_X1 U11425 ( .A1(n6442), .A2(n13586), .ZN(n9000) );
  NAND2_X1 U11426 ( .A1(n13482), .A2(n9081), .ZN(n9012) );
  NAND2_X1 U11427 ( .A1(n9003), .A2(n9002), .ZN(n9004) );
  NAND2_X1 U11428 ( .A1(n13264), .A2(n9043), .ZN(n9010) );
  INV_X1 U11429 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n15257) );
  NAND2_X1 U11430 ( .A1(n9074), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U11431 ( .A1(n8767), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9006) );
  OAI211_X1 U11432 ( .C1(n8537), .C2(n15257), .A(n9007), .B(n9006), .ZN(n9008)
         );
  INV_X1 U11433 ( .A(n9008), .ZN(n9009) );
  NAND2_X1 U11434 ( .A1(n13240), .A2(n8728), .ZN(n9011) );
  NAND2_X1 U11435 ( .A1(n9012), .A2(n9011), .ZN(n9014) );
  AOI22_X1 U11436 ( .A1(n13482), .A2(n8728), .B1(n6436), .B2(n13240), .ZN(
        n9013) );
  INV_X1 U11437 ( .A(n13259), .ZN(n12923) );
  NAND2_X1 U11438 ( .A1(n13477), .A2(n9081), .ZN(n9015) );
  OAI21_X1 U11439 ( .B1(n12923), .B2(n8887), .A(n9015), .ZN(n9016) );
  MUX2_X1 U11440 ( .A(n11590), .B(n13581), .S(n9479), .Z(n9033) );
  INV_X1 U11441 ( .A(n9033), .ZN(n9036) );
  XNOR2_X1 U11442 ( .A(n9036), .B(SI_27_), .ZN(n9020) );
  NAND2_X1 U11443 ( .A1(n11589), .A2(n9100), .ZN(n9022) );
  OR2_X1 U11444 ( .A1(n6442), .A2(n13581), .ZN(n9021) );
  NAND2_X1 U11445 ( .A1(n13472), .A2(n6436), .ZN(n9031) );
  XNOR2_X1 U11446 ( .A(n9070), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13231) );
  NAND2_X1 U11447 ( .A1(n13231), .A2(n9043), .ZN(n9029) );
  INV_X1 U11448 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9026) );
  NAND2_X1 U11449 ( .A1(n9074), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U11450 ( .A1(n9073), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9023) );
  OAI211_X1 U11451 ( .C1(n9026), .C2(n9025), .A(n9024), .B(n9023), .ZN(n9027)
         );
  INV_X1 U11452 ( .A(n9027), .ZN(n9028) );
  NAND2_X1 U11453 ( .A1(n13241), .A2(n8728), .ZN(n9030) );
  AOI22_X1 U11454 ( .A1(n13472), .A2(n8728), .B1(n9081), .B2(n13241), .ZN(
        n9032) );
  NAND2_X1 U11455 ( .A1(n9033), .A2(n11491), .ZN(n9034) );
  NAND2_X1 U11456 ( .A1(n9036), .A2(SI_27_), .ZN(n9037) );
  MUX2_X1 U11457 ( .A(n14346), .B(n12057), .S(n9479), .Z(n9038) );
  NAND2_X1 U11458 ( .A1(n9038), .A2(n12122), .ZN(n9041) );
  INV_X1 U11459 ( .A(n9038), .ZN(n9039) );
  NAND2_X1 U11460 ( .A1(n9039), .A2(SI_28_), .ZN(n9040) );
  NAND2_X1 U11461 ( .A1(n9041), .A2(n9040), .ZN(n9067) );
  INV_X1 U11462 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11597) );
  INV_X1 U11463 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11798) );
  MUX2_X1 U11464 ( .A(n11597), .B(n11798), .S(n9833), .Z(n9053) );
  XNOR2_X1 U11465 ( .A(n9053), .B(SI_29_), .ZN(n9052) );
  OR2_X1 U11466 ( .A1(n6442), .A2(n11798), .ZN(n9042) );
  INV_X1 U11467 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12922) );
  INV_X1 U11468 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n12969) );
  INV_X1 U11469 ( .A(n9071), .ZN(n12089) );
  NAND2_X1 U11470 ( .A1(n12089), .A2(n9043), .ZN(n9049) );
  INV_X1 U11471 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U11472 ( .A1(n8767), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U11473 ( .A1(n9074), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9044) );
  OAI211_X1 U11474 ( .C1(n9046), .C2(n8537), .A(n9045), .B(n9044), .ZN(n9047)
         );
  INV_X1 U11475 ( .A(n9047), .ZN(n9048) );
  NAND2_X1 U11476 ( .A1(n9049), .A2(n9048), .ZN(n13209) );
  AOI22_X1 U11477 ( .A1(n13462), .A2(n8728), .B1(n6436), .B2(n13209), .ZN(
        n9113) );
  INV_X1 U11478 ( .A(n13209), .ZN(n9126) );
  NAND2_X1 U11479 ( .A1(n13462), .A2(n8958), .ZN(n9050) );
  INV_X1 U11480 ( .A(n9157), .ZN(n9796) );
  OAI211_X1 U11481 ( .C1(n9126), .C2(n8887), .A(n9050), .B(n9796), .ZN(n9112)
         );
  NOR2_X1 U11482 ( .A1(n9113), .A2(n9112), .ZN(n9089) );
  INV_X1 U11483 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11807) );
  INV_X1 U11484 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12124) );
  MUX2_X1 U11485 ( .A(n11807), .B(n12124), .S(n9833), .Z(n9056) );
  INV_X1 U11486 ( .A(SI_30_), .ZN(n12859) );
  NAND2_X1 U11487 ( .A1(n9056), .A2(n12859), .ZN(n9095) );
  INV_X1 U11488 ( .A(SI_29_), .ZN(n12863) );
  NAND2_X1 U11489 ( .A1(n9053), .A2(n12863), .ZN(n9093) );
  NAND2_X1 U11490 ( .A1(n9095), .A2(n9093), .ZN(n9061) );
  MUX2_X1 U11491 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9479), .Z(n9054) );
  INV_X1 U11492 ( .A(SI_31_), .ZN(n12852) );
  XNOR2_X1 U11493 ( .A(n9054), .B(n12852), .ZN(n9059) );
  NOR2_X1 U11494 ( .A1(n9061), .A2(n9059), .ZN(n9055) );
  NAND2_X1 U11495 ( .A1(n9094), .A2(n9055), .ZN(n9065) );
  INV_X1 U11496 ( .A(n9056), .ZN(n9057) );
  NAND2_X1 U11497 ( .A1(n9057), .A2(SI_30_), .ZN(n9096) );
  INV_X1 U11498 ( .A(n9059), .ZN(n9062) );
  XNOR2_X1 U11499 ( .A(n9059), .B(n9096), .ZN(n9060) );
  OAI21_X1 U11500 ( .B1(n9062), .B2(n9061), .A(n9060), .ZN(n9063) );
  INV_X1 U11501 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n15195) );
  OAI21_X1 U11502 ( .B1(n13458), .B2(n9108), .A(n9121), .ZN(n9086) );
  NAND2_X1 U11503 ( .A1(n12056), .A2(n9100), .ZN(n9069) );
  OR2_X1 U11504 ( .A1(n6442), .A2(n12057), .ZN(n9068) );
  OAI21_X1 U11505 ( .B1(n9070), .B2(n12922), .A(n12969), .ZN(n9072) );
  NAND2_X1 U11506 ( .A1(n9072), .A2(n9071), .ZN(n13218) );
  OR2_X1 U11507 ( .A1(n13218), .A2(n8986), .ZN(n9079) );
  INV_X1 U11508 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13217) );
  NAND2_X1 U11509 ( .A1(n9073), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U11510 ( .A1(n9074), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9075) );
  OAI211_X1 U11511 ( .C1(n13217), .C2(n9025), .A(n9076), .B(n9075), .ZN(n9077)
         );
  INV_X1 U11512 ( .A(n9077), .ZN(n9078) );
  AND2_X1 U11513 ( .A1(n13227), .A2(n8728), .ZN(n9080) );
  AOI21_X1 U11514 ( .B1(n13465), .B2(n6436), .A(n9080), .ZN(n9088) );
  NAND2_X1 U11515 ( .A1(n13465), .A2(n8728), .ZN(n9083) );
  NAND2_X1 U11516 ( .A1(n13227), .A2(n9081), .ZN(n9082) );
  NAND2_X1 U11517 ( .A1(n9083), .A2(n9082), .ZN(n9087) );
  NAND2_X1 U11518 ( .A1(n9088), .A2(n9087), .ZN(n9084) );
  INV_X1 U11519 ( .A(n13458), .ZN(n9090) );
  NAND2_X1 U11520 ( .A1(n9090), .A2(n8728), .ZN(n9091) );
  OAI211_X1 U11521 ( .C1(n9108), .C2(n9122), .A(n9121), .B(n9091), .ZN(n9092)
         );
  NAND2_X1 U11522 ( .A1(n9094), .A2(n9093), .ZN(n9098) );
  AND2_X1 U11523 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  INV_X1 U11524 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9101) );
  OR2_X1 U11525 ( .A1(n8537), .A2(n9101), .ZN(n9106) );
  INV_X1 U11526 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9102) );
  OR2_X1 U11527 ( .A1(n9025), .A2(n9102), .ZN(n9105) );
  INV_X1 U11528 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9103) );
  OR2_X1 U11529 ( .A1(n8507), .A2(n9103), .ZN(n9104) );
  AND3_X1 U11530 ( .A1(n9106), .A2(n9105), .A3(n9104), .ZN(n9107) );
  OAI22_X1 U11531 ( .A1(n9125), .A2(n8887), .B1(n9107), .B2(n9122), .ZN(n9118)
         );
  INV_X1 U11532 ( .A(n9108), .ZN(n13196) );
  NAND2_X1 U11533 ( .A1(n13196), .A2(n8728), .ZN(n9120) );
  INV_X1 U11534 ( .A(n9109), .ZN(n9110) );
  NAND2_X1 U11535 ( .A1(n9120), .A2(n9110), .ZN(n9111) );
  INV_X1 U11536 ( .A(n9112), .ZN(n9115) );
  INV_X1 U11537 ( .A(n9113), .ZN(n9114) );
  OAI22_X1 U11538 ( .A1(n9118), .A2(n9117), .B1(n9115), .B2(n9114), .ZN(n9116)
         );
  INV_X1 U11539 ( .A(n9118), .ZN(n9119) );
  OAI211_X1 U11540 ( .C1(n13458), .C2(n9122), .A(n9121), .B(n9120), .ZN(n9123)
         );
  XNOR2_X1 U11541 ( .A(n9125), .B(n13097), .ZN(n9142) );
  XNOR2_X1 U11542 ( .A(n13462), .B(n9126), .ZN(n12118) );
  NAND2_X1 U11543 ( .A1(n13465), .A2(n12926), .ZN(n9127) );
  INV_X1 U11544 ( .A(n13240), .ZN(n9128) );
  NAND2_X1 U11545 ( .A1(n13482), .A2(n9128), .ZN(n12081) );
  OR2_X1 U11546 ( .A1(n13482), .A2(n9128), .ZN(n9129) );
  INV_X1 U11547 ( .A(n13477), .ZN(n13248) );
  NAND2_X1 U11548 ( .A1(n13248), .A2(n13259), .ZN(n9130) );
  NAND2_X1 U11549 ( .A1(n13477), .A2(n12923), .ZN(n12082) );
  NAND2_X1 U11550 ( .A1(n9130), .A2(n12082), .ZN(n12058) );
  XNOR2_X1 U11551 ( .A(n13492), .B(n13040), .ZN(n13291) );
  INV_X1 U11552 ( .A(n13258), .ZN(n12080) );
  XNOR2_X1 U11553 ( .A(n13498), .B(n13098), .ZN(n13310) );
  INV_X1 U11554 ( .A(n13099), .ZN(n13350) );
  NAND2_X1 U11555 ( .A1(n13511), .A2(n13350), .ZN(n12074) );
  OR2_X1 U11556 ( .A1(n13511), .A2(n13350), .ZN(n9131) );
  NAND2_X1 U11557 ( .A1(n12074), .A2(n9131), .ZN(n13334) );
  INV_X1 U11558 ( .A(n13104), .ZN(n13423) );
  XNOR2_X1 U11559 ( .A(n13538), .B(n13423), .ZN(n13415) );
  INV_X1 U11560 ( .A(n13101), .ZN(n13349) );
  XNOR2_X1 U11561 ( .A(n13522), .B(n13349), .ZN(n13364) );
  NAND2_X1 U11562 ( .A1(n13527), .A2(n13102), .ZN(n12101) );
  NAND2_X1 U11563 ( .A1(n12102), .A2(n12101), .ZN(n13383) );
  XNOR2_X1 U11564 ( .A(n13543), .B(n13421), .ZN(n13439) );
  XNOR2_X1 U11565 ( .A(n12092), .B(n12059), .ZN(n11458) );
  XNOR2_X1 U11566 ( .A(n13549), .B(n11455), .ZN(n11451) );
  XNOR2_X1 U11567 ( .A(n10965), .B(n10864), .ZN(n10967) );
  INV_X1 U11568 ( .A(n13110), .ZN(n10941) );
  XNOR2_X1 U11569 ( .A(n10942), .B(n10941), .ZN(n10865) );
  NAND2_X1 U11570 ( .A1(n13118), .A2(n14867), .ZN(n10369) );
  NAND2_X1 U11571 ( .A1(n10369), .A2(n10295), .ZN(n14902) );
  NOR3_X1 U11572 ( .A1(n10661), .A2(n11586), .A3(n14902), .ZN(n9132) );
  NAND4_X1 U11573 ( .A1(n9132), .A2(n10836), .A3(n10817), .A4(n10296), .ZN(
        n9133) );
  XNOR2_X1 U11574 ( .A(n6592), .B(n13112), .ZN(n10816) );
  NOR4_X1 U11575 ( .A1(n10967), .A2(n10865), .A3(n9133), .A4(n10816), .ZN(
        n9134) );
  XNOR2_X1 U11576 ( .A(n11380), .B(n13107), .ZN(n11378) );
  XNOR2_X1 U11577 ( .A(n11109), .B(n13109), .ZN(n10946) );
  NAND4_X1 U11578 ( .A1(n9134), .A2(n11378), .A3(n11155), .A4(n10946), .ZN(
        n9135) );
  NOR4_X1 U11579 ( .A1(n13439), .A2(n11458), .A3(n11451), .A4(n9135), .ZN(
        n9136) );
  XNOR2_X1 U11580 ( .A(n13533), .B(n13103), .ZN(n13388) );
  XNOR2_X1 U11581 ( .A(n13434), .B(n13442), .ZN(n13426) );
  NAND4_X1 U11582 ( .A1(n13383), .A2(n9136), .A3(n13388), .A4(n13426), .ZN(
        n9137) );
  NOR4_X1 U11583 ( .A1(n13334), .A2(n13415), .A3(n13364), .A4(n9137), .ZN(
        n9138) );
  XNOR2_X1 U11584 ( .A(n13516), .B(n13100), .ZN(n13347) );
  XNOR2_X1 U11585 ( .A(n13325), .B(n13300), .ZN(n13318) );
  NAND4_X1 U11586 ( .A1(n13310), .A2(n9138), .A3(n13347), .A4(n13318), .ZN(
        n9139) );
  NOR4_X1 U11587 ( .A1(n12058), .A2(n13291), .A3(n13279), .A4(n9139), .ZN(
        n9140) );
  NAND4_X1 U11588 ( .A1(n13207), .A2(n13257), .A3(n9140), .A4(n13226), .ZN(
        n9141) );
  XOR2_X1 U11589 ( .A(n10655), .B(n9144), .Z(n9145) );
  NAND2_X1 U11590 ( .A1(n9796), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11508) );
  NAND2_X1 U11591 ( .A1(n9147), .A2(n9146), .ZN(n9148) );
  NAND2_X1 U11592 ( .A1(n9148), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U11593 ( .A1(n6468), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9151) );
  MUX2_X1 U11594 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9151), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9153) );
  NAND2_X1 U11595 ( .A1(n9153), .A2(n9152), .ZN(n13583) );
  NAND2_X1 U11596 ( .A1(n9154), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9155) );
  MUX2_X1 U11597 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9155), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9156) );
  NAND2_X1 U11598 ( .A1(n9156), .A2(n6468), .ZN(n13585) );
  INV_X1 U11599 ( .A(n13579), .ZN(n12086) );
  INV_X1 U11600 ( .A(n9159), .ZN(n9790) );
  INV_X1 U11601 ( .A(n9788), .ZN(n9160) );
  NAND4_X1 U11602 ( .A1(n14895), .A2(n12086), .A3(n13444), .A4(n9160), .ZN(
        n9161) );
  OAI211_X1 U11603 ( .C1(n9167), .C2(n11508), .A(n9161), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9162) );
  INV_X1 U11604 ( .A(n9162), .ZN(n9163) );
  AOI21_X1 U11605 ( .B1(n9165), .B2(n9164), .A(n9163), .ZN(n9175) );
  INV_X1 U11606 ( .A(n9694), .ZN(n9166) );
  OAI211_X1 U11607 ( .C1(n10655), .C2(n11137), .A(n9166), .B(n9788), .ZN(n9170) );
  MUX2_X1 U11608 ( .A(n11137), .B(n9693), .S(n11586), .Z(n9168) );
  INV_X1 U11609 ( .A(n11508), .ZN(n9172) );
  NOR2_X1 U11610 ( .A1(n9172), .A2(P2_B_REG_SCAN_IN), .ZN(n9173) );
  AOI21_X1 U11611 ( .B1(n9175), .B2(n9174), .A(n9173), .ZN(P2_U3328) );
  AND2_X1 U11612 ( .A1(n9178), .A2(n9177), .ZN(n9181) );
  NOR2_X1 U11613 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9180) );
  NOR2_X1 U11614 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .ZN(n9179) );
  NOR2_X1 U11615 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9185) );
  NOR2_X1 U11616 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9184) );
  INV_X1 U11617 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9192) );
  INV_X1 U11618 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9929) );
  INV_X1 U11619 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10761) );
  INV_X1 U11620 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9955) );
  NAND2_X1 U11621 ( .A1(n9202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9204) );
  INV_X1 U11622 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9837) );
  NAND2_X1 U11623 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9208) );
  MUX2_X1 U11624 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9208), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9210) );
  INV_X1 U11625 ( .A(n9209), .ZN(n9223) );
  NAND2_X1 U11626 ( .A1(n9210), .A2(n9223), .ZN(n10033) );
  OR2_X1 U11627 ( .A1(n9863), .A2(n10033), .ZN(n9211) );
  NAND2_X1 U11628 ( .A1(n9228), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9217) );
  INV_X1 U11629 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10892) );
  INV_X1 U11630 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14592) );
  OR2_X1 U11631 ( .A1(n9254), .A2(n14592), .ZN(n9215) );
  INV_X1 U11632 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10893) );
  INV_X1 U11633 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13879) );
  NOR2_X1 U11634 ( .A1(n9833), .A2(n9831), .ZN(n9218) );
  XNOR2_X1 U11635 ( .A(n9218), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14359) );
  MUX2_X1 U11636 ( .A(n13879), .B(n14359), .S(n9863), .Z(n10750) );
  NAND2_X1 U11637 ( .A1(n13874), .A2(n10896), .ZN(n10166) );
  INV_X1 U11638 ( .A(n10166), .ZN(n10749) );
  OAI22_X1 U11639 ( .A1(n10748), .A2(n10749), .B1(n6936), .B2(n9212), .ZN(
        n10877) );
  INV_X1 U11640 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13882) );
  OR2_X1 U11641 ( .A1(n9520), .A2(n13882), .ZN(n9221) );
  INV_X1 U11642 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9934) );
  INV_X1 U11643 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9960) );
  OR2_X1 U11644 ( .A1(n11802), .A2(n9960), .ZN(n9219) );
  NAND2_X1 U11645 ( .A1(n9223), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9225) );
  XNOR2_X1 U11646 ( .A(n9225), .B(n9224), .ZN(n13890) );
  NOR2_X1 U11647 ( .A1(n13872), .A2(n11832), .ZN(n9227) );
  NAND2_X1 U11648 ( .A1(n13872), .A2(n11832), .ZN(n9226) );
  OAI21_X1 U11649 ( .B1(n10877), .B2(n9227), .A(n9226), .ZN(n10735) );
  INV_X1 U11650 ( .A(n10735), .ZN(n9238) );
  NAND2_X1 U11651 ( .A1(n9228), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9232) );
  INV_X1 U11652 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10742) );
  OR2_X1 U11653 ( .A1(n11802), .A2(n10742), .ZN(n9231) );
  OR2_X1 U11654 ( .A1(n9254), .A2(n13907), .ZN(n9230) );
  OR2_X1 U11655 ( .A1(n9520), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U11656 ( .A1(n9233), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9234) );
  XNOR2_X1 U11657 ( .A(n9234), .B(n9176), .ZN(n13906) );
  OR2_X1 U11658 ( .A1(n9834), .A2(n9527), .ZN(n9236) );
  INV_X1 U11659 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9835) );
  OR2_X1 U11660 ( .A1(n11978), .A2(n9835), .ZN(n9235) );
  OAI211_X1 U11661 ( .C1(n9863), .C2(n13906), .A(n9236), .B(n9235), .ZN(n11839) );
  INV_X1 U11662 ( .A(n11987), .ZN(n9237) );
  OR2_X1 U11663 ( .A1(n13871), .A2(n11839), .ZN(n9239) );
  INV_X1 U11664 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9954) );
  OR2_X1 U11665 ( .A1(n11802), .A2(n9954), .ZN(n9243) );
  INV_X1 U11666 ( .A(n9250), .ZN(n9252) );
  INV_X1 U11667 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9241) );
  INV_X1 U11668 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9240) );
  NAND2_X1 U11669 ( .A1(n9241), .A2(n9240), .ZN(n9242) );
  NAND2_X1 U11670 ( .A1(n9252), .A2(n9242), .ZN(n10615) );
  INV_X1 U11671 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U11672 ( .A1(n9844), .A2(n9527), .ZN(n9248) );
  NAND2_X1 U11673 ( .A1(n9244), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9245) );
  MUX2_X1 U11674 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9245), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9246) );
  INV_X1 U11675 ( .A(n6485), .ZN(n9388) );
  NAND2_X1 U11676 ( .A1(n9246), .A2(n9388), .ZN(n13928) );
  OAI22_X1 U11677 ( .A1(n11978), .A2(n6901), .B1(n9863), .B2(n13928), .ZN(
        n9247) );
  NAND2_X1 U11678 ( .A1(n13870), .A2(n14700), .ZN(n9249) );
  NAND2_X1 U11679 ( .A1(n9228), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9259) );
  INV_X1 U11680 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10643) );
  OR2_X1 U11681 ( .A1(n11802), .A2(n10643), .ZN(n9258) );
  INV_X1 U11682 ( .A(n9273), .ZN(n9275) );
  INV_X1 U11683 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U11684 ( .A1(n9252), .A2(n9251), .ZN(n9253) );
  NAND2_X1 U11685 ( .A1(n9275), .A2(n9253), .ZN(n10703) );
  OR2_X1 U11686 ( .A1(n9520), .A2(n10703), .ZN(n9257) );
  INV_X1 U11687 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9255) );
  OR2_X1 U11688 ( .A1(n9254), .A2(n9255), .ZN(n9256) );
  NAND4_X1 U11689 ( .A1(n9259), .A2(n9258), .A3(n9257), .A4(n9256), .ZN(n13869) );
  OR2_X1 U11690 ( .A1(n9841), .A2(n9527), .ZN(n9262) );
  NAND2_X1 U11691 ( .A1(n9388), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9260) );
  XNOR2_X1 U11692 ( .A(n9260), .B(P1_IR_REG_5__SCAN_IN), .ZN(n13941) );
  AOI22_X1 U11693 ( .A1(n9446), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9445), .B2(
        n13941), .ZN(n9261) );
  NAND2_X1 U11694 ( .A1(n9262), .A2(n9261), .ZN(n14708) );
  AND2_X1 U11695 ( .A1(n13869), .A2(n14708), .ZN(n9265) );
  INV_X1 U11696 ( .A(n13869), .ZN(n9263) );
  NAND2_X1 U11697 ( .A1(n9263), .A2(n10704), .ZN(n9264) );
  OR2_X1 U11698 ( .A1(n9859), .A2(n9527), .ZN(n9272) );
  NAND2_X1 U11699 ( .A1(n9267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9266) );
  MUX2_X1 U11700 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9266), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n9270) );
  INV_X1 U11701 ( .A(n9267), .ZN(n9269) );
  INV_X1 U11702 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U11703 ( .A1(n9269), .A2(n9268), .ZN(n9296) );
  NAND2_X1 U11704 ( .A1(n9270), .A2(n9296), .ZN(n13951) );
  INV_X1 U11705 ( .A(n13951), .ZN(n9971) );
  AOI22_X1 U11706 ( .A1(n9446), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9445), .B2(
        n9971), .ZN(n9271) );
  NAND2_X1 U11707 ( .A1(n9228), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9281) );
  INV_X1 U11708 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9968) );
  OR2_X1 U11709 ( .A1(n11802), .A2(n9968), .ZN(n9280) );
  INV_X1 U11710 ( .A(n9287), .ZN(n9277) );
  INV_X1 U11711 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9274) );
  NAND2_X1 U11712 ( .A1(n9275), .A2(n9274), .ZN(n9276) );
  NAND2_X1 U11713 ( .A1(n9277), .A2(n9276), .ZN(n14643) );
  OR2_X1 U11714 ( .A1(n9520), .A2(n14643), .ZN(n9279) );
  INV_X1 U11715 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9941) );
  OR2_X1 U11716 ( .A1(n9254), .A2(n9941), .ZN(n9278) );
  NAND4_X1 U11717 ( .A1(n9281), .A2(n9280), .A3(n9279), .A4(n9278), .ZN(n13868) );
  XNOR2_X1 U11718 ( .A(n14647), .B(n13868), .ZN(n11993) );
  OR2_X1 U11719 ( .A1(n14647), .A2(n13868), .ZN(n9282) );
  NAND2_X1 U11720 ( .A1(n9283), .A2(n9282), .ZN(n10798) );
  NAND2_X1 U11721 ( .A1(n9868), .A2(n11980), .ZN(n9286) );
  NAND2_X1 U11722 ( .A1(n9296), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9284) );
  XNOR2_X1 U11723 ( .A(n9284), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13970) );
  AOI22_X1 U11724 ( .A1(n9446), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9445), .B2(
        n13970), .ZN(n9285) );
  NAND2_X1 U11725 ( .A1(n9228), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9291) );
  INV_X1 U11726 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9942) );
  OR2_X1 U11727 ( .A1(n9254), .A2(n9942), .ZN(n9290) );
  NAND2_X1 U11728 ( .A1(n9287), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9300) );
  OAI21_X1 U11729 ( .B1(n9287), .B2(P1_REG3_REG_7__SCAN_IN), .A(n9300), .ZN(
        n11124) );
  OR2_X1 U11730 ( .A1(n9520), .A2(n11124), .ZN(n9289) );
  INV_X1 U11731 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10805) );
  OR2_X1 U11732 ( .A1(n11802), .A2(n10805), .ZN(n9288) );
  INV_X1 U11733 ( .A(n14620), .ZN(n9292) );
  OR2_X1 U11734 ( .A1(n14724), .A2(n9292), .ZN(n14613) );
  NAND2_X1 U11735 ( .A1(n14724), .A2(n9292), .ZN(n9293) );
  NAND2_X1 U11736 ( .A1(n10798), .A2(n10799), .ZN(n9295) );
  OR2_X1 U11737 ( .A1(n14724), .A2(n14620), .ZN(n9294) );
  NAND2_X1 U11738 ( .A1(n9295), .A2(n9294), .ZN(n14627) );
  INV_X1 U11739 ( .A(n14627), .ZN(n9307) );
  NAND2_X1 U11740 ( .A1(n9873), .A2(n11980), .ZN(n9298) );
  NAND2_X1 U11741 ( .A1(n9346), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9309) );
  XNOR2_X1 U11742 ( .A(n9309), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U11743 ( .A1(n9446), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9445), .B2(
        n9991), .ZN(n9297) );
  NAND2_X1 U11744 ( .A1(n9228), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9305) );
  INV_X1 U11745 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9974) );
  OR2_X1 U11746 ( .A1(n11802), .A2(n9974), .ZN(n9304) );
  AND2_X1 U11747 ( .A1(n9300), .A2(n9299), .ZN(n9301) );
  NOR2_X1 U11748 ( .A1(n9300), .A2(n9299), .ZN(n9313) );
  OR2_X1 U11749 ( .A1(n9301), .A2(n9313), .ZN(n15302) );
  OR2_X1 U11750 ( .A1(n9520), .A2(n15302), .ZN(n9303) );
  INV_X1 U11751 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9927) );
  OR2_X1 U11752 ( .A1(n9254), .A2(n9927), .ZN(n9302) );
  NAND2_X1 U11753 ( .A1(n15310), .A2(n13867), .ZN(n11859) );
  INV_X1 U11754 ( .A(n11859), .ZN(n9306) );
  NAND2_X1 U11755 ( .A1(n9884), .A2(n11980), .ZN(n9312) );
  INV_X1 U11756 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U11757 ( .A1(n9309), .A2(n9308), .ZN(n9310) );
  NAND2_X1 U11758 ( .A1(n9310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9322) );
  XNOR2_X1 U11759 ( .A(n9322), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10014) );
  AOI22_X1 U11760 ( .A1(n9446), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9445), .B2(
        n10014), .ZN(n9311) );
  NAND2_X1 U11761 ( .A1(n9228), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9319) );
  INV_X1 U11762 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9992) );
  OR2_X1 U11763 ( .A1(n11802), .A2(n9992), .ZN(n9318) );
  NAND2_X1 U11764 ( .A1(n9313), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9328) );
  OR2_X1 U11765 ( .A1(n9313), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9314) );
  NAND2_X1 U11766 ( .A1(n9328), .A2(n9314), .ZN(n11032) );
  OR2_X1 U11767 ( .A1(n9520), .A2(n11032), .ZN(n9317) );
  INV_X1 U11768 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9315) );
  OR2_X1 U11769 ( .A1(n9254), .A2(n9315), .ZN(n9316) );
  XNOR2_X1 U11770 ( .A(n7189), .B(n13866), .ZN(n11997) );
  INV_X1 U11771 ( .A(n11997), .ZN(n11030) );
  NAND2_X1 U11772 ( .A1(n11031), .A2(n11030), .ZN(n11029) );
  NAND2_X1 U11773 ( .A1(n11873), .A2(n14618), .ZN(n9320) );
  NAND2_X1 U11774 ( .A1(n11029), .A2(n9320), .ZN(n11176) );
  NAND2_X1 U11775 ( .A1(n9922), .A2(n11980), .ZN(n9326) );
  INV_X1 U11776 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9321) );
  NAND2_X1 U11777 ( .A1(n9322), .A2(n9321), .ZN(n9323) );
  NAND2_X1 U11778 ( .A1(n9323), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9324) );
  XNOR2_X1 U11779 ( .A(n9324), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10041) );
  AOI22_X1 U11780 ( .A1(n9446), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9445), 
        .B2(n10041), .ZN(n9325) );
  NAND2_X1 U11781 ( .A1(n9228), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U11782 ( .A1(n9328), .A2(n9327), .ZN(n9329) );
  NAND2_X1 U11783 ( .A1(n9337), .A2(n9329), .ZN(n11362) );
  OR2_X1 U11784 ( .A1(n9520), .A2(n11362), .ZN(n9333) );
  INV_X1 U11785 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9330) );
  OR2_X1 U11786 ( .A1(n9254), .A2(n9330), .ZN(n9332) );
  INV_X1 U11787 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11179) );
  OR2_X1 U11788 ( .A1(n11802), .A2(n11179), .ZN(n9331) );
  NAND4_X1 U11789 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n14525) );
  XNOR2_X1 U11790 ( .A(n14741), .B(n14525), .ZN(n11998) );
  INV_X1 U11791 ( .A(n11998), .ZN(n11175) );
  NAND2_X1 U11792 ( .A1(n11176), .A2(n11175), .ZN(n11174) );
  OR2_X1 U11793 ( .A1(n14741), .A2(n14525), .ZN(n9335) );
  NAND2_X1 U11794 ( .A1(n9228), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9342) );
  INV_X1 U11795 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9336) );
  AND2_X1 U11796 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  OR2_X1 U11797 ( .A1(n9338), .A2(n9353), .ZN(n14536) );
  OR2_X1 U11798 ( .A1(n9520), .A2(n14536), .ZN(n9341) );
  INV_X1 U11799 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10034) );
  OR2_X1 U11800 ( .A1(n9254), .A2(n10034), .ZN(n9340) );
  INV_X1 U11801 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10042) );
  OR2_X1 U11802 ( .A1(n11802), .A2(n10042), .ZN(n9339) );
  NAND4_X1 U11803 ( .A1(n9342), .A2(n9341), .A3(n9340), .A4(n9339), .ZN(n14406) );
  NAND2_X1 U11804 ( .A1(n10002), .A2(n11980), .ZN(n9349) );
  INV_X1 U11805 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U11806 ( .A1(n9344), .A2(n9343), .ZN(n9345) );
  NAND2_X1 U11807 ( .A1(n9350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9347) );
  XNOR2_X1 U11808 ( .A(n9347), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10058) );
  AOI22_X1 U11809 ( .A1(n9446), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9445), 
        .B2(n10058), .ZN(n9348) );
  NAND2_X1 U11810 ( .A1(n10072), .A2(n11980), .ZN(n9352) );
  OAI21_X1 U11811 ( .B1(n9350), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9360) );
  XNOR2_X1 U11812 ( .A(n9360), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U11813 ( .A1(n9446), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9445), 
        .B2(n10229), .ZN(n9351) );
  NAND2_X1 U11814 ( .A1(n9228), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9358) );
  INV_X1 U11815 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10052) );
  OR2_X1 U11816 ( .A1(n11802), .A2(n10052), .ZN(n9357) );
  NOR2_X1 U11817 ( .A1(n9353), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9354) );
  OR2_X1 U11818 ( .A1(n9364), .A2(n9354), .ZN(n14408) );
  OR2_X1 U11819 ( .A1(n9520), .A2(n14408), .ZN(n9356) );
  OR2_X1 U11820 ( .A1(n9254), .A2(n14424), .ZN(n9355) );
  NAND4_X1 U11821 ( .A1(n9358), .A2(n9357), .A3(n9356), .A4(n9355), .ZN(n14527) );
  XNOR2_X1 U11822 ( .A(n14410), .B(n14527), .ZN(n12000) );
  NAND2_X1 U11823 ( .A1(n10122), .A2(n11980), .ZN(n9363) );
  INV_X1 U11824 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U11825 ( .A1(n9360), .A2(n9359), .ZN(n9361) );
  NAND2_X1 U11826 ( .A1(n9361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9374) );
  XNOR2_X1 U11827 ( .A(n9374), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U11828 ( .A1(n9446), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9445), 
        .B2(n10244), .ZN(n9362) );
  NAND2_X1 U11829 ( .A1(n9228), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9370) );
  INV_X1 U11830 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11500) );
  OR2_X1 U11831 ( .A1(n11802), .A2(n11500), .ZN(n9369) );
  NAND2_X1 U11832 ( .A1(n9364), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9380) );
  OR2_X1 U11833 ( .A1(n9364), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9365) );
  NAND2_X1 U11834 ( .A1(n9380), .A2(n9365), .ZN(n11581) );
  OR2_X1 U11835 ( .A1(n9520), .A2(n11581), .ZN(n9368) );
  INV_X1 U11836 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9366) );
  OR2_X1 U11837 ( .A1(n9254), .A2(n9366), .ZN(n9367) );
  NAND4_X1 U11838 ( .A1(n9370), .A2(n9369), .A3(n9368), .A4(n9367), .ZN(n14405) );
  INV_X1 U11839 ( .A(n14405), .ZN(n11568) );
  XNOR2_X1 U11840 ( .A(n11897), .B(n11568), .ZN(n12002) );
  NAND2_X1 U11841 ( .A1(n11498), .A2(n12002), .ZN(n9372) );
  OR2_X1 U11842 ( .A1(n11897), .A2(n14405), .ZN(n9371) );
  NAND2_X1 U11843 ( .A1(n10337), .A2(n11980), .ZN(n9378) );
  INV_X1 U11844 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U11845 ( .A1(n9374), .A2(n9373), .ZN(n9375) );
  NAND2_X1 U11846 ( .A1(n9375), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9376) );
  AOI22_X1 U11847 ( .A1(n9445), .A2(n10716), .B1(n9446), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9377) );
  NAND2_X1 U11848 ( .A1(n9228), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9385) );
  INV_X1 U11849 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10710) );
  OR2_X1 U11850 ( .A1(n9254), .A2(n10710), .ZN(n9384) );
  INV_X1 U11851 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9379) );
  NAND2_X1 U11852 ( .A1(n9380), .A2(n9379), .ZN(n9381) );
  NAND2_X1 U11853 ( .A1(n9393), .A2(n9381), .ZN(n14228) );
  OR2_X1 U11854 ( .A1(n9520), .A2(n14228), .ZN(n9383) );
  INV_X1 U11855 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10245) );
  OR2_X1 U11856 ( .A1(n11802), .A2(n10245), .ZN(n9382) );
  OR2_X1 U11857 ( .A1(n14233), .A2(n13850), .ZN(n11900) );
  NAND2_X1 U11858 ( .A1(n14233), .A2(n13850), .ZN(n11893) );
  NAND2_X1 U11859 ( .A1(n11900), .A2(n11893), .ZN(n14219) );
  INV_X1 U11860 ( .A(n14219), .ZN(n14235) );
  INV_X1 U11861 ( .A(n13850), .ZN(n13865) );
  NAND2_X1 U11862 ( .A1(n14233), .A2(n13865), .ZN(n9386) );
  NAND2_X1 U11863 ( .A1(n10389), .A2(n11980), .ZN(n9391) );
  OR2_X1 U11864 ( .A1(n9388), .A2(n9387), .ZN(n9401) );
  NAND2_X1 U11865 ( .A1(n9401), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9389) );
  XNOR2_X1 U11866 ( .A(n9389), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U11867 ( .A1(n9446), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9445), 
        .B2(n10719), .ZN(n9390) );
  NAND2_X1 U11868 ( .A1(n9228), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9399) );
  INV_X1 U11869 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n14212) );
  OR2_X1 U11870 ( .A1(n11802), .A2(n14212), .ZN(n9398) );
  INV_X1 U11871 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U11872 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U11873 ( .A1(n9410), .A2(n9394), .ZN(n14211) );
  OR2_X1 U11874 ( .A1(n9520), .A2(n14211), .ZN(n9397) );
  INV_X1 U11875 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9395) );
  OR2_X1 U11876 ( .A1(n9254), .A2(n9395), .ZN(n9396) );
  NAND2_X1 U11877 ( .A1(n14214), .A2(n14508), .ZN(n11904) );
  NAND2_X1 U11878 ( .A1(n11901), .A2(n11904), .ZN(n14208) );
  INV_X1 U11879 ( .A(n14508), .ZN(n14222) );
  NAND2_X1 U11880 ( .A1(n10311), .A2(n11980), .ZN(n9408) );
  INV_X1 U11881 ( .A(n9401), .ZN(n9403) );
  NAND2_X1 U11882 ( .A1(n9403), .A2(n9402), .ZN(n9405) );
  NAND2_X1 U11883 ( .A1(n9405), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9404) );
  MUX2_X1 U11884 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9404), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9406) );
  AOI22_X1 U11885 ( .A1(n9446), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9445), 
        .B2(n10982), .ZN(n9407) );
  INV_X1 U11886 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9409) );
  AND2_X1 U11887 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  OR2_X1 U11888 ( .A1(n9411), .A2(n9424), .ZN(n14521) );
  INV_X1 U11889 ( .A(n14521), .ZN(n14197) );
  INV_X1 U11890 ( .A(n9520), .ZN(n9471) );
  NAND2_X1 U11891 ( .A1(n14197), .A2(n9471), .ZN(n9415) );
  NAND2_X1 U11892 ( .A1(n9228), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9414) );
  INV_X1 U11893 ( .A(n9254), .ZN(n9463) );
  NAND2_X1 U11894 ( .A1(n9463), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11895 ( .A1(n9637), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9412) );
  NAND4_X1 U11896 ( .A1(n9415), .A2(n9414), .A3(n9413), .A4(n9412), .ZN(n14182) );
  INV_X1 U11897 ( .A(n14182), .ZN(n13851) );
  XNOR2_X1 U11898 ( .A(n14518), .B(n13851), .ZN(n12004) );
  NAND2_X1 U11899 ( .A1(n14187), .A2(n12004), .ZN(n9417) );
  OR2_X1 U11900 ( .A1(n14518), .A2(n14182), .ZN(n9416) );
  NAND2_X1 U11901 ( .A1(n10387), .A2(n11980), .ZN(n9423) );
  NAND2_X1 U11902 ( .A1(n9418), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9419) );
  MUX2_X1 U11903 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9419), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9421) );
  NAND2_X1 U11904 ( .A1(n9421), .A2(n6766), .ZN(n11320) );
  AOI22_X1 U11905 ( .A1(n9446), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9445), 
        .B2(n11322), .ZN(n9422) );
  OR2_X1 U11906 ( .A1(n9424), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U11907 ( .A1(n9452), .A2(n9425), .ZN(n14175) );
  INV_X1 U11908 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9426) );
  OAI22_X1 U11909 ( .A1(n14175), .A2(n9520), .B1(n9254), .B2(n9426), .ZN(n9429) );
  INV_X1 U11910 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14176) );
  NAND2_X1 U11911 ( .A1(n9228), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9427) );
  OAI21_X1 U11912 ( .B1(n14176), .B2(n11802), .A(n9427), .ZN(n9428) );
  AND2_X1 U11913 ( .A1(n14311), .A2(n14511), .ZN(n9430) );
  OR2_X1 U11914 ( .A1(n14311), .A2(n14511), .ZN(n9431) );
  OR2_X1 U11915 ( .A1(n10566), .A2(n9527), .ZN(n9434) );
  NAND2_X1 U11916 ( .A1(n6766), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9432) );
  XNOR2_X1 U11917 ( .A(n9432), .B(P1_IR_REG_18__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U11918 ( .A1(n9446), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9445), 
        .B2(n11515), .ZN(n9433) );
  XNOR2_X1 U11919 ( .A(n9452), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14167) );
  NAND2_X1 U11920 ( .A1(n14167), .A2(n9471), .ZN(n9440) );
  INV_X1 U11921 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U11922 ( .A1(n9637), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U11923 ( .A1(n9228), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9435) );
  OAI211_X1 U11924 ( .C1(n9437), .C2(n9254), .A(n9436), .B(n9435), .ZN(n9438)
         );
  INV_X1 U11925 ( .A(n9438), .ZN(n9439) );
  NAND2_X1 U11926 ( .A1(n9440), .A2(n9439), .ZN(n14183) );
  AND2_X1 U11927 ( .A1(n14306), .A2(n14183), .ZN(n9441) );
  NAND2_X1 U11928 ( .A1(n10850), .A2(n11980), .ZN(n9448) );
  NAND2_X1 U11929 ( .A1(n9571), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9444) );
  AOI22_X1 U11930 ( .A1(n9446), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14230), 
        .B2(n9445), .ZN(n9447) );
  INV_X1 U11931 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9450) );
  INV_X1 U11932 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9449) );
  OAI21_X1 U11933 ( .B1(n9452), .B2(n9450), .A(n9449), .ZN(n9453) );
  NAND2_X1 U11934 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n9451) );
  AND2_X1 U11935 ( .A1(n9453), .A2(n9461), .ZN(n14150) );
  NAND2_X1 U11936 ( .A1(n14150), .A2(n9471), .ZN(n9456) );
  AOI22_X1 U11937 ( .A1(n9637), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9228), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U11938 ( .A1(n9463), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9454) );
  OR2_X1 U11939 ( .A1(n14299), .A2(n14164), .ZN(n11925) );
  NAND2_X1 U11940 ( .A1(n14299), .A2(n14164), .ZN(n11926) );
  NAND2_X1 U11941 ( .A1(n11925), .A2(n11926), .ZN(n14147) );
  INV_X1 U11942 ( .A(n14164), .ZN(n13864) );
  OR2_X1 U11943 ( .A1(n14299), .A2(n13864), .ZN(n9457) );
  NAND2_X1 U11944 ( .A1(n9458), .A2(n9457), .ZN(n14135) );
  OR2_X1 U11945 ( .A1(n11978), .A2(n11014), .ZN(n9459) );
  INV_X1 U11946 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9460) );
  AND2_X1 U11947 ( .A1(n9461), .A2(n9460), .ZN(n9462) );
  OR2_X1 U11948 ( .A1(n9462), .A2(n9469), .ZN(n14131) );
  AOI22_X1 U11949 ( .A1(n9637), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9228), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U11950 ( .A1(n9463), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9464) );
  OAI211_X1 U11951 ( .C1(n14131), .C2(n9520), .A(n9465), .B(n9464), .ZN(n14144) );
  INV_X1 U11952 ( .A(n14144), .ZN(n13649) );
  XNOR2_X1 U11953 ( .A(n14293), .B(n13649), .ZN(n14126) );
  INV_X1 U11954 ( .A(n14126), .ZN(n14134) );
  OR2_X1 U11955 ( .A1(n13650), .A2(n13649), .ZN(n9466) );
  OR2_X1 U11956 ( .A1(n11138), .A2(n9527), .ZN(n9468) );
  OR2_X1 U11957 ( .A1(n11978), .A2(n11136), .ZN(n9467) );
  OR2_X1 U11958 ( .A1(n9469), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U11959 ( .A1(n9469), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9482) );
  AND2_X1 U11960 ( .A1(n9470), .A2(n9482), .ZN(n14115) );
  NAND2_X1 U11961 ( .A1(n14115), .A2(n9471), .ZN(n9477) );
  INV_X1 U11962 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U11963 ( .A1(n9228), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U11964 ( .A1(n9637), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9472) );
  OAI211_X1 U11965 ( .C1(n9254), .C2(n9474), .A(n9473), .B(n9472), .ZN(n9475)
         );
  INV_X1 U11966 ( .A(n9475), .ZN(n9476) );
  NAND2_X1 U11967 ( .A1(n9477), .A2(n9476), .ZN(n13863) );
  INV_X1 U11968 ( .A(n13863), .ZN(n14128) );
  XNOR2_X1 U11969 ( .A(n14288), .B(n14128), .ZN(n14111) );
  INV_X1 U11970 ( .A(n14111), .ZN(n14121) );
  OR2_X1 U11971 ( .A1(n14288), .A2(n13863), .ZN(n9478) );
  NAND2_X1 U11972 ( .A1(n14118), .A2(n9478), .ZN(n14094) );
  OR2_X1 U11973 ( .A1(n9480), .A2(n9833), .ZN(n9481) );
  XNOR2_X1 U11974 ( .A(n9481), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14358) );
  NAND2_X1 U11975 ( .A1(n9637), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9488) );
  INV_X1 U11976 ( .A(n9494), .ZN(n9496) );
  OAI21_X1 U11977 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n9483), .A(n9496), .ZN(
        n14097) );
  OR2_X1 U11978 ( .A1(n9520), .A2(n14097), .ZN(n9486) );
  INV_X1 U11979 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9484) );
  OR2_X1 U11980 ( .A1(n9254), .A2(n9484), .ZN(n9485) );
  NAND4_X1 U11981 ( .A1(n9488), .A2(n9487), .A3(n9486), .A4(n9485), .ZN(n13862) );
  NAND2_X1 U11982 ( .A1(n14100), .A2(n13862), .ZN(n9489) );
  INV_X1 U11983 ( .A(n14103), .ZN(n9490) );
  OR2_X1 U11984 ( .A1(n14283), .A2(n13862), .ZN(n9491) );
  NAND2_X1 U11985 ( .A1(n11507), .A2(n11980), .ZN(n9493) );
  INV_X1 U11986 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11506) );
  OR2_X1 U11987 ( .A1(n11978), .A2(n11506), .ZN(n9492) );
  NAND2_X1 U11988 ( .A1(n9637), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9502) );
  INV_X1 U11989 ( .A(n9505), .ZN(n9507) );
  INV_X1 U11990 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U11991 ( .A1(n9496), .A2(n9495), .ZN(n9497) );
  NAND2_X1 U11992 ( .A1(n9507), .A2(n9497), .ZN(n14087) );
  OR2_X1 U11993 ( .A1(n9520), .A2(n14087), .ZN(n9500) );
  INV_X1 U11994 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9498) );
  OR2_X1 U11995 ( .A1(n9254), .A2(n9498), .ZN(n9499) );
  NAND4_X1 U11996 ( .A1(n9502), .A2(n9501), .A3(n9500), .A4(n9499), .ZN(n13861) );
  XNOR2_X1 U11997 ( .A(n14089), .B(n13861), .ZN(n14084) );
  OR2_X1 U11998 ( .A1(n11978), .A2(n14354), .ZN(n9503) );
  NAND2_X1 U11999 ( .A1(n9637), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9514) );
  INV_X1 U12000 ( .A(n9519), .ZN(n9509) );
  INV_X1 U12001 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9506) );
  NAND2_X1 U12002 ( .A1(n9507), .A2(n9506), .ZN(n9508) );
  NAND2_X1 U12003 ( .A1(n9509), .A2(n9508), .ZN(n14069) );
  OR2_X1 U12004 ( .A1(n9520), .A2(n14069), .ZN(n9512) );
  INV_X1 U12005 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9510) );
  OR2_X1 U12006 ( .A1(n9254), .A2(n9510), .ZN(n9511) );
  NAND4_X1 U12007 ( .A1(n9514), .A2(n9513), .A3(n9512), .A4(n9511), .ZN(n13860) );
  XNOR2_X1 U12008 ( .A(n14274), .B(n13860), .ZN(n12009) );
  OR2_X1 U12009 ( .A1(n14274), .A2(n13860), .ZN(n9515) );
  NAND2_X1 U12010 ( .A1(n13584), .A2(n11980), .ZN(n9517) );
  INV_X1 U12011 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15215) );
  OR2_X1 U12012 ( .A1(n11978), .A2(n15215), .ZN(n9516) );
  NAND2_X1 U12013 ( .A1(n9228), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9525) );
  INV_X1 U12014 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9518) );
  OR2_X1 U12015 ( .A1(n9254), .A2(n9518), .ZN(n9524) );
  NAND2_X1 U12016 ( .A1(n9519), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9530) );
  OAI21_X1 U12017 ( .B1(n9519), .B2(P1_REG3_REG_25__SCAN_IN), .A(n9530), .ZN(
        n14049) );
  OR2_X1 U12018 ( .A1(n9520), .A2(n14049), .ZN(n9523) );
  INV_X1 U12019 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9521) );
  OR2_X1 U12020 ( .A1(n11802), .A2(n9521), .ZN(n9522) );
  NAND4_X1 U12021 ( .A1(n9525), .A2(n9524), .A3(n9523), .A4(n9522), .ZN(n14029) );
  XNOR2_X1 U12022 ( .A(n14269), .B(n14029), .ZN(n14045) );
  INV_X1 U12023 ( .A(n14045), .ZN(n14051) );
  NAND2_X1 U12024 ( .A1(n14269), .A2(n14029), .ZN(n9526) );
  NAND2_X1 U12025 ( .A1(n14050), .A2(n9526), .ZN(n14033) );
  OR2_X1 U12026 ( .A1(n11978), .A2(n14347), .ZN(n9528) );
  NAND2_X1 U12027 ( .A1(n9637), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9536) );
  INV_X1 U12028 ( .A(n9530), .ZN(n9531) );
  NAND2_X1 U12029 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n9531), .ZN(n9542) );
  OAI21_X1 U12030 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n9531), .A(n9542), .ZN(
        n14035) );
  OR2_X1 U12031 ( .A1(n9520), .A2(n14035), .ZN(n9534) );
  INV_X1 U12032 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9532) );
  OR2_X1 U12033 ( .A1(n9254), .A2(n9532), .ZN(n9533) );
  NAND4_X1 U12034 ( .A1(n9536), .A2(n9535), .A3(n9534), .A4(n9533), .ZN(n13859) );
  NAND2_X1 U12035 ( .A1(n14264), .A2(n13859), .ZN(n9537) );
  NAND2_X1 U12036 ( .A1(n11589), .A2(n11980), .ZN(n9539) );
  OR2_X1 U12037 ( .A1(n11978), .A2(n11590), .ZN(n9538) );
  NAND2_X1 U12038 ( .A1(n9637), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9547) );
  INV_X1 U12039 ( .A(n9542), .ZN(n9540) );
  NAND2_X1 U12040 ( .A1(n9540), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9554) );
  INV_X1 U12041 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U12042 ( .A1(n9542), .A2(n9541), .ZN(n9543) );
  NAND2_X1 U12043 ( .A1(n9554), .A2(n9543), .ZN(n14020) );
  OR2_X1 U12044 ( .A1(n9520), .A2(n14020), .ZN(n9545) );
  INV_X1 U12045 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n15207) );
  OR2_X1 U12046 ( .A1(n9254), .A2(n15207), .ZN(n9544) );
  XNOR2_X1 U12047 ( .A(n14022), .B(n14030), .ZN(n12011) );
  OR2_X1 U12048 ( .A1(n14022), .A2(n14030), .ZN(n9549) );
  NAND2_X1 U12049 ( .A1(n12056), .A2(n11980), .ZN(n9551) );
  OR2_X1 U12050 ( .A1(n11978), .A2(n14346), .ZN(n9550) );
  NAND2_X1 U12051 ( .A1(n9637), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9560) );
  INV_X1 U12052 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15278) );
  INV_X1 U12053 ( .A(n9554), .ZN(n9552) );
  NAND2_X1 U12054 ( .A1(n9552), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9645) );
  INV_X1 U12055 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9553) );
  NAND2_X1 U12056 ( .A1(n9554), .A2(n9553), .ZN(n9555) );
  NAND2_X1 U12057 ( .A1(n9645), .A2(n9555), .ZN(n14003) );
  OR2_X1 U12058 ( .A1(n9520), .A2(n14003), .ZN(n9558) );
  INV_X1 U12059 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9556) );
  OR2_X1 U12060 ( .A1(n9254), .A2(n9556), .ZN(n9557) );
  NAND4_X1 U12061 ( .A1(n9560), .A2(n9559), .A3(n9558), .A4(n9557), .ZN(n13858) );
  NAND2_X1 U12062 ( .A1(n14252), .A2(n13858), .ZN(n9562) );
  OR2_X1 U12063 ( .A1(n14252), .A2(n13858), .ZN(n9561) );
  NAND2_X1 U12064 ( .A1(n9562), .A2(n9561), .ZN(n13994) );
  INV_X1 U12065 ( .A(n13994), .ZN(n14008) );
  NAND2_X1 U12066 ( .A1(n9637), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9568) );
  INV_X1 U12067 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9563) );
  OR2_X1 U12068 ( .A1(n9520), .A2(n9645), .ZN(n9566) );
  INV_X1 U12069 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9564) );
  OR2_X1 U12070 ( .A1(n9254), .A2(n9564), .ZN(n9565) );
  NAND4_X1 U12071 ( .A1(n9568), .A2(n9567), .A3(n9566), .A4(n9565), .ZN(n13996) );
  NAND2_X1 U12072 ( .A1(n11591), .A2(n11980), .ZN(n9570) );
  OR2_X1 U12073 ( .A1(n11978), .A2(n11597), .ZN(n9569) );
  XOR2_X1 U12074 ( .A(n13996), .B(n14247), .Z(n12015) );
  NAND2_X1 U12075 ( .A1(n9584), .A2(n9572), .ZN(n9582) );
  OAI21_X1 U12076 ( .B1(n9582), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9574) );
  OAI21_X1 U12077 ( .B1(n9575), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9576) );
  MUX2_X1 U12078 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9576), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9578) );
  INV_X1 U12079 ( .A(n9577), .ZN(n9579) );
  NAND2_X1 U12080 ( .A1(n9579), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9580) );
  NAND2_X1 U12081 ( .A1(n9575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9581) );
  AND3_X2 U12082 ( .A1(n14350), .A2(n9593), .A3(n9594), .ZN(n10457) );
  NAND2_X1 U12083 ( .A1(n14357), .A2(n6895), .ZN(n11984) );
  INV_X1 U12084 ( .A(n11984), .ZN(n10149) );
  NAND2_X1 U12085 ( .A1(n11981), .A2(n11525), .ZN(n9588) );
  AND2_X1 U12086 ( .A1(n10149), .A2(n9588), .ZN(n10458) );
  INV_X1 U12087 ( .A(P1_B_REG_SCAN_IN), .ZN(n9642) );
  NOR2_X1 U12088 ( .A1(n14350), .A2(n9642), .ZN(n9589) );
  MUX2_X1 U12089 ( .A(n9589), .B(n9642), .S(n9594), .Z(n9590) );
  INV_X1 U12090 ( .A(n9590), .ZN(n9591) );
  OR2_X1 U12091 ( .A1(n9877), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9592) );
  OR2_X1 U12092 ( .A1(n9593), .A2(n14350), .ZN(n9881) );
  NAND2_X1 U12093 ( .A1(n9592), .A2(n9881), .ZN(n10162) );
  INV_X1 U12094 ( .A(n10162), .ZN(n10148) );
  OR2_X1 U12095 ( .A1(n9877), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9595) );
  INV_X1 U12096 ( .A(n9593), .ZN(n14348) );
  INV_X1 U12097 ( .A(n9594), .ZN(n14355) );
  NAND2_X1 U12098 ( .A1(n14348), .A2(n14355), .ZN(n9879) );
  NOR4_X1 U12099 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9604) );
  NOR4_X1 U12100 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9603) );
  INV_X1 U12101 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15193) );
  INV_X1 U12102 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15214) );
  INV_X1 U12103 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15243) );
  INV_X1 U12104 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14683) );
  NAND4_X1 U12105 ( .A1(n15193), .A2(n15214), .A3(n15243), .A4(n14683), .ZN(
        n9601) );
  NOR4_X1 U12106 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n9599) );
  NOR4_X1 U12107 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9598) );
  NOR4_X1 U12108 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n9597) );
  NOR4_X1 U12109 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9596) );
  NAND4_X1 U12110 ( .A1(n9599), .A2(n9598), .A3(n9597), .A4(n9596), .ZN(n9600)
         );
  NOR4_X1 U12111 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n9601), .A4(n9600), .ZN(n9602) );
  AND3_X1 U12112 ( .A1(n9604), .A2(n9603), .A3(n9602), .ZN(n9605) );
  OR2_X1 U12113 ( .A1(n9877), .A2(n9605), .ZN(n10163) );
  NAND4_X1 U12114 ( .A1(n12040), .A2(n10148), .A3(n10171), .A4(n10163), .ZN(
        n9646) );
  NAND2_X1 U12115 ( .A1(n14725), .A2(n14230), .ZN(n10455) );
  AND2_X1 U12116 ( .A1(n11984), .A2(n11525), .ZN(n9607) );
  NAND2_X1 U12117 ( .A1(n14357), .A2(n11525), .ZN(n11811) );
  INV_X1 U12118 ( .A(n11823), .ZN(n9606) );
  NAND2_X1 U12119 ( .A1(n9607), .A2(n13750), .ZN(n10756) );
  NAND2_X1 U12120 ( .A1(n11823), .A2(n14230), .ZN(n11985) );
  AND2_X1 U12121 ( .A1(n10756), .A2(n11985), .ZN(n9608) );
  INV_X1 U12122 ( .A(n14269), .ZN(n9629) );
  INV_X1 U12123 ( .A(n14288), .ZN(n14117) );
  INV_X2 U12124 ( .A(n11832), .ZN(n14692) );
  NAND2_X1 U12125 ( .A1(n13872), .A2(n14692), .ZN(n9609) );
  INV_X1 U12126 ( .A(n11839), .ZN(n11840) );
  OR2_X1 U12127 ( .A1(n13871), .A2(n11840), .ZN(n9611) );
  NAND2_X1 U12128 ( .A1(n13870), .A2(n10616), .ZN(n9613) );
  AND2_X1 U12129 ( .A1(n10704), .A2(n13869), .ZN(n9614) );
  INV_X1 U12130 ( .A(n13868), .ZN(n9615) );
  NAND2_X1 U12131 ( .A1(n14647), .A2(n9615), .ZN(n9616) );
  OR2_X1 U12132 ( .A1(n15310), .A2(n11266), .ZN(n11868) );
  NAND2_X1 U12133 ( .A1(n15310), .A2(n11266), .ZN(n11864) );
  OR2_X1 U12134 ( .A1(n11873), .A2(n13866), .ZN(n9619) );
  OR2_X1 U12135 ( .A1(n14741), .A2(n6791), .ZN(n9620) );
  NAND2_X1 U12136 ( .A1(n11170), .A2(n9620), .ZN(n11345) );
  NAND2_X1 U12137 ( .A1(n11882), .A2(n11552), .ZN(n9621) );
  OR2_X1 U12138 ( .A1(n11882), .A2(n11552), .ZN(n9622) );
  INV_X1 U12139 ( .A(n14527), .ZN(n11496) );
  OR2_X1 U12140 ( .A1(n14410), .A2(n11496), .ZN(n9623) );
  INV_X1 U12141 ( .A(n12002), .ZN(n9624) );
  OR2_X1 U12142 ( .A1(n11897), .A2(n11568), .ZN(n9625) );
  NAND2_X1 U12143 ( .A1(n14518), .A2(n13851), .ZN(n9626) );
  XNOR2_X1 U12144 ( .A(n7184), .B(n14511), .ZN(n14172) );
  INV_X1 U12145 ( .A(n14172), .ZN(n14180) );
  XNOR2_X1 U12146 ( .A(n14306), .B(n14183), .ZN(n14160) );
  OR2_X1 U12147 ( .A1(n14306), .A2(n7100), .ZN(n11817) );
  INV_X1 U12148 ( .A(n13861), .ZN(n13821) );
  INV_X1 U12149 ( .A(n13858), .ZN(n13753) );
  NAND2_X1 U12150 ( .A1(n14357), .A2(n14230), .ZN(n9632) );
  NAND2_X1 U12151 ( .A1(n6895), .A2(n12018), .ZN(n9631) );
  INV_X1 U12152 ( .A(n14344), .ZN(n13877) );
  INV_X1 U12153 ( .A(n14264), .ZN(n13847) );
  NAND2_X1 U12154 ( .A1(n10751), .A2(n10750), .ZN(n10883) );
  NAND2_X1 U12155 ( .A1(n10645), .A2(n10704), .ZN(n10646) );
  OR2_X1 U12156 ( .A1(n10646), .A2(n14647), .ZN(n14648) );
  INV_X1 U12157 ( .A(n15310), .ZN(n14737) );
  NOR2_X2 U12158 ( .A1(n14225), .A2(n14233), .ZN(n14209) );
  NAND2_X1 U12159 ( .A1(n13650), .A2(n14149), .ZN(n14136) );
  INV_X1 U12160 ( .A(n14725), .ZN(n14715) );
  AOI21_X1 U12161 ( .B1(n14001), .B2(n14247), .A(n14715), .ZN(n9635) );
  OR2_X1 U12162 ( .A1(n9646), .A2(n14230), .ZN(n14216) );
  NAND2_X1 U12163 ( .A1(n10167), .A2(n12018), .ZN(n10151) );
  INV_X1 U12164 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12165 ( .A1(n9637), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U12166 ( .A1(n9228), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9638) );
  OAI211_X1 U12167 ( .C1(n9254), .C2(n9640), .A(n9639), .B(n9638), .ZN(n13857)
         );
  INV_X1 U12168 ( .A(n13857), .ZN(n9644) );
  NOR2_X1 U12169 ( .A1(n6440), .A2(n9642), .ZN(n9643) );
  OR2_X1 U12170 ( .A1(n14617), .A2(n9643), .ZN(n13981) );
  NOR2_X1 U12171 ( .A1(n9644), .A2(n13981), .ZN(n14246) );
  INV_X1 U12172 ( .A(n14246), .ZN(n9647) );
  OAI22_X1 U12173 ( .A1(n9647), .A2(n9646), .B1(n9645), .B2(n14229), .ZN(n9648) );
  AOI21_X1 U12174 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14625), .A(n9648), .ZN(
        n9649) );
  OAI21_X1 U12175 ( .B1(n7180), .B2(n14190), .A(n9649), .ZN(n9650) );
  INV_X1 U12176 ( .A(n12478), .ZN(n12349) );
  AND2_X1 U12177 ( .A1(n12057), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U12178 ( .A1(n14346), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9655) );
  XNOR2_X1 U12179 ( .A(n11798), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n11594) );
  XNOR2_X1 U12180 ( .A(n11596), .B(n11594), .ZN(n12860) );
  NAND2_X1 U12181 ( .A1(n12860), .A2(n11616), .ZN(n9657) );
  OR2_X1 U12182 ( .A1(n6441), .A2(n12863), .ZN(n9656) );
  NAND2_X1 U12183 ( .A1(n9657), .A2(n9656), .ZN(n9686) );
  NAND2_X1 U12184 ( .A1(n9686), .A2(n12210), .ZN(n11620) );
  XNOR2_X1 U12185 ( .A(n9658), .B(n9672), .ZN(n9669) );
  INV_X1 U12186 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n15240) );
  NAND2_X1 U12187 ( .A1(n7726), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U12188 ( .A1(n9659), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9660) );
  OAI211_X1 U12189 ( .C1(n15240), .C2(n9662), .A(n9661), .B(n9660), .ZN(n9663)
         );
  INV_X1 U12190 ( .A(n9663), .ZN(n9664) );
  NAND2_X1 U12191 ( .A1(n11611), .A2(n9664), .ZN(n12348) );
  AND2_X1 U12192 ( .A1(n9665), .A2(P3_B_REG_SCAN_IN), .ZN(n9666) );
  NOR2_X1 U12193 ( .A1(n15046), .A2(n9666), .ZN(n12462) );
  AOI22_X1 U12194 ( .A1(n15069), .A2(n12349), .B1(n12348), .B2(n12462), .ZN(
        n9667) );
  INV_X1 U12195 ( .A(n11749), .ZN(n9670) );
  INV_X1 U12196 ( .A(n9672), .ZN(n9673) );
  XNOR2_X1 U12197 ( .A(n10539), .B(n12847), .ZN(n9676) );
  AND2_X1 U12198 ( .A1(n10358), .A2(n9674), .ZN(n9675) );
  NAND2_X1 U12199 ( .A1(n9676), .A2(n9675), .ZN(n10493) );
  NAND2_X1 U12200 ( .A1(n12847), .A2(n11758), .ZN(n9683) );
  OAI211_X1 U12201 ( .C1(n11793), .C2(n9678), .A(n10538), .B(n9677), .ZN(n9679) );
  INV_X1 U12202 ( .A(n9679), .ZN(n9680) );
  NAND2_X1 U12203 ( .A1(n10496), .A2(n9680), .ZN(n9681) );
  OAI21_X1 U12204 ( .B1(n10496), .B2(n10494), .A(n9681), .ZN(n9682) );
  MUX2_X1 U12205 ( .A(n9683), .B(n9682), .S(n11754), .Z(n9684) );
  INV_X1 U12206 ( .A(n9686), .ZN(n12048) );
  NAND2_X1 U12207 ( .A1(n9687), .A2(n7649), .ZN(P3_U3488) );
  INV_X1 U12208 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U12209 ( .A1(n9689), .A2(n7653), .ZN(P3_U3456) );
  INV_X1 U12210 ( .A(n10457), .ZN(n10146) );
  INV_X1 U12211 ( .A(n9690), .ZN(n9691) );
  INV_X2 U12212 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  XNOR2_X1 U12213 ( .A(n13543), .B(n12966), .ZN(n9695) );
  NAND2_X1 U12214 ( .A1(n9693), .A2(n11137), .ZN(n9781) );
  INV_X1 U12215 ( .A(n11586), .ZN(n10300) );
  OR2_X2 U12216 ( .A1(n9781), .A2(n10300), .ZN(n9733) );
  AND2_X1 U12217 ( .A1(n13105), .A2(n9733), .ZN(n9696) );
  NAND2_X1 U12218 ( .A1(n9695), .A2(n9696), .ZN(n12865) );
  INV_X1 U12219 ( .A(n9695), .ZN(n12934) );
  INV_X1 U12220 ( .A(n9696), .ZN(n9697) );
  NAND2_X1 U12221 ( .A1(n12934), .A2(n9697), .ZN(n9698) );
  NAND2_X1 U12222 ( .A1(n12865), .A2(n9698), .ZN(n9780) );
  OR2_X1 U12223 ( .A1(n14867), .A2(n9733), .ZN(n9699) );
  NAND2_X1 U12224 ( .A1(n10295), .A2(n9699), .ZN(n10366) );
  AND2_X1 U12225 ( .A1(n12966), .A2(n14867), .ZN(n9700) );
  NAND2_X1 U12226 ( .A1(n13116), .A2(n9733), .ZN(n9702) );
  INV_X1 U12227 ( .A(n9701), .ZN(n9703) );
  NAND2_X1 U12228 ( .A1(n9703), .A2(n9702), .ZN(n9704) );
  NAND2_X1 U12229 ( .A1(n10399), .A2(n9704), .ZN(n13050) );
  XNOR2_X1 U12230 ( .A(n12966), .B(n10658), .ZN(n9706) );
  NAND2_X1 U12231 ( .A1(n13115), .A2(n12864), .ZN(n9705) );
  NAND2_X1 U12232 ( .A1(n9706), .A2(n9705), .ZN(n9710) );
  INV_X1 U12233 ( .A(n9705), .ZN(n9708) );
  INV_X1 U12234 ( .A(n9706), .ZN(n9707) );
  NAND2_X1 U12235 ( .A1(n9708), .A2(n9707), .ZN(n9709) );
  AND2_X1 U12236 ( .A1(n9710), .A2(n9709), .ZN(n13051) );
  INV_X1 U12237 ( .A(n10819), .ZN(n14914) );
  XNOR2_X1 U12238 ( .A(n12966), .B(n14914), .ZN(n9712) );
  NAND2_X1 U12239 ( .A1(n13114), .A2(n12864), .ZN(n9711) );
  XNOR2_X1 U12240 ( .A(n9712), .B(n9711), .ZN(n10518) );
  INV_X1 U12241 ( .A(n9711), .ZN(n9714) );
  INV_X1 U12242 ( .A(n9712), .ZN(n9713) );
  NAND2_X1 U12243 ( .A1(n9714), .A2(n9713), .ZN(n9715) );
  XNOR2_X1 U12244 ( .A(n12900), .B(n10845), .ZN(n9717) );
  NAND2_X1 U12245 ( .A1(n13113), .A2(n12864), .ZN(n9716) );
  NAND2_X1 U12246 ( .A1(n9717), .A2(n9716), .ZN(n9721) );
  INV_X1 U12247 ( .A(n9716), .ZN(n9719) );
  INV_X1 U12248 ( .A(n9717), .ZN(n9718) );
  NAND2_X1 U12249 ( .A1(n9719), .A2(n9718), .ZN(n9720) );
  AND2_X1 U12250 ( .A1(n9721), .A2(n9720), .ZN(n10524) );
  XNOR2_X1 U12251 ( .A(n14931), .B(n12900), .ZN(n9722) );
  NAND2_X1 U12252 ( .A1(n13112), .A2(n12864), .ZN(n9723) );
  NAND2_X1 U12253 ( .A1(n9722), .A2(n9723), .ZN(n9727) );
  INV_X1 U12254 ( .A(n9722), .ZN(n9725) );
  INV_X1 U12255 ( .A(n9723), .ZN(n9724) );
  NAND2_X1 U12256 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  AND2_X1 U12257 ( .A1(n9727), .A2(n9726), .ZN(n10508) );
  XNOR2_X1 U12258 ( .A(n10965), .B(n12900), .ZN(n9728) );
  NAND2_X1 U12259 ( .A1(n13111), .A2(n12864), .ZN(n9729) );
  XNOR2_X1 U12260 ( .A(n9728), .B(n9729), .ZN(n10530) );
  INV_X1 U12261 ( .A(n9728), .ZN(n9731) );
  INV_X1 U12262 ( .A(n9729), .ZN(n9730) );
  NAND2_X1 U12263 ( .A1(n9731), .A2(n9730), .ZN(n9732) );
  NAND2_X1 U12264 ( .A1(n13110), .A2(n9733), .ZN(n9734) );
  XNOR2_X1 U12265 ( .A(n9736), .B(n9734), .ZN(n10679) );
  INV_X1 U12266 ( .A(n9734), .ZN(n9735) );
  NAND2_X1 U12267 ( .A1(n9736), .A2(n9735), .ZN(n9737) );
  XNOR2_X1 U12268 ( .A(n11109), .B(n12966), .ZN(n10928) );
  NAND2_X1 U12269 ( .A1(n10930), .A2(n10928), .ZN(n9738) );
  AND2_X1 U12270 ( .A1(n13109), .A2(n9733), .ZN(n10929) );
  NAND2_X1 U12271 ( .A1(n10928), .A2(n10929), .ZN(n10927) );
  NAND2_X1 U12272 ( .A1(n10930), .A2(n10929), .ZN(n9739) );
  XNOR2_X1 U12273 ( .A(n11232), .B(n12966), .ZN(n9740) );
  NAND2_X1 U12274 ( .A1(n13108), .A2(n9733), .ZN(n9741) );
  XNOR2_X1 U12275 ( .A(n9740), .B(n9741), .ZN(n11151) );
  INV_X1 U12276 ( .A(n9740), .ZN(n9742) );
  NAND2_X1 U12277 ( .A1(n9742), .A2(n9741), .ZN(n9743) );
  XNOR2_X1 U12278 ( .A(n11380), .B(n12966), .ZN(n9744) );
  AND2_X1 U12279 ( .A1(n13107), .A2(n9733), .ZN(n9745) );
  NAND2_X1 U12280 ( .A1(n9744), .A2(n9745), .ZN(n9748) );
  INV_X1 U12281 ( .A(n9744), .ZN(n11398) );
  INV_X1 U12282 ( .A(n9745), .ZN(n9746) );
  NAND2_X1 U12283 ( .A1(n11398), .A2(n9746), .ZN(n9747) );
  AND2_X1 U12284 ( .A1(n9748), .A2(n9747), .ZN(n11186) );
  XNOR2_X1 U12285 ( .A(n13549), .B(n12966), .ZN(n11423) );
  NAND2_X1 U12286 ( .A1(n13106), .A2(n9733), .ZN(n9750) );
  XNOR2_X1 U12287 ( .A(n11423), .B(n9750), .ZN(n11401) );
  AND2_X1 U12288 ( .A1(n11401), .A2(n9748), .ZN(n9749) );
  INV_X1 U12289 ( .A(n11423), .ZN(n9751) );
  NAND2_X1 U12290 ( .A1(n9751), .A2(n9750), .ZN(n9752) );
  NAND2_X1 U12291 ( .A1(n11422), .A2(n9752), .ZN(n9753) );
  XNOR2_X1 U12292 ( .A(n12092), .B(n12966), .ZN(n9754) );
  NAND2_X1 U12293 ( .A1(n13445), .A2(n12864), .ZN(n9755) );
  XNOR2_X1 U12294 ( .A(n9754), .B(n9755), .ZN(n11424) );
  NAND2_X1 U12295 ( .A1(n9753), .A2(n11424), .ZN(n11430) );
  INV_X1 U12296 ( .A(n9754), .ZN(n9756) );
  NAND2_X1 U12297 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  NOR4_X1 U12298 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n9766) );
  INV_X1 U12299 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15183) );
  INV_X1 U12300 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15210) );
  INV_X1 U12301 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15246) );
  INV_X1 U12302 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15268) );
  NAND4_X1 U12303 ( .A1(n15183), .A2(n15210), .A3(n15246), .A4(n15268), .ZN(
        n9763) );
  NOR4_X1 U12304 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n9761) );
  NOR4_X1 U12305 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9760) );
  NOR4_X1 U12306 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9759) );
  NOR4_X1 U12307 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9758) );
  NAND4_X1 U12308 ( .A1(n9761), .A2(n9760), .A3(n9759), .A4(n9758), .ZN(n9762)
         );
  NOR4_X1 U12309 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n9763), .A4(n9762), .ZN(n9765) );
  NOR4_X1 U12310 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9764) );
  NAND3_X1 U12311 ( .A1(n9766), .A2(n9765), .A3(n9764), .ZN(n9770) );
  INV_X1 U12312 ( .A(n13583), .ZN(n9769) );
  XNOR2_X1 U12313 ( .A(n13591), .B(P2_B_REG_SCAN_IN), .ZN(n9767) );
  NAND2_X1 U12314 ( .A1(n13585), .A2(n9767), .ZN(n9768) );
  AND2_X1 U12315 ( .A1(n9770), .A2(n14891), .ZN(n10306) );
  INV_X1 U12316 ( .A(n10306), .ZN(n9776) );
  NAND2_X1 U12317 ( .A1(n13591), .A2(n13583), .ZN(n9772) );
  INV_X1 U12318 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15212) );
  NAND2_X1 U12319 ( .A1(n14891), .A2(n15212), .ZN(n9771) );
  NAND2_X1 U12320 ( .A1(n9772), .A2(n9771), .ZN(n14894) );
  INV_X1 U12321 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14898) );
  NAND2_X1 U12322 ( .A1(n14891), .A2(n14898), .ZN(n9774) );
  NAND2_X1 U12323 ( .A1(n13583), .A2(n13585), .ZN(n9773) );
  NAND2_X1 U12324 ( .A1(n9774), .A2(n9773), .ZN(n10651) );
  NOR2_X1 U12325 ( .A1(n14894), .A2(n10651), .ZN(n9775) );
  NAND2_X1 U12326 ( .A1(n9776), .A2(n9775), .ZN(n9784) );
  INV_X1 U12327 ( .A(n9784), .ZN(n9777) );
  NAND2_X1 U12328 ( .A1(n9777), .A2(n14895), .ZN(n9789) );
  INV_X1 U12329 ( .A(n9781), .ZN(n14878) );
  OR2_X1 U12330 ( .A1(n14930), .A2(n9158), .ZN(n9778) );
  INV_X1 U12331 ( .A(n12866), .ZN(n12936) );
  AOI211_X1 U12332 ( .C1(n9780), .C2(n9779), .A(n13082), .B(n12936), .ZN(n9794) );
  OR2_X1 U12333 ( .A1(n9781), .A2(n11586), .ZN(n10670) );
  OR2_X1 U12334 ( .A1(n9789), .A2(n10670), .ZN(n9783) );
  INV_X1 U12335 ( .A(n10307), .ZN(n9782) );
  NOR2_X1 U12336 ( .A1(n6590), .A2(n13023), .ZN(n9793) );
  NAND2_X1 U12337 ( .A1(n9784), .A2(n10307), .ZN(n9787) );
  AND2_X1 U12338 ( .A1(n9158), .A2(n9788), .ZN(n10305) );
  NOR2_X1 U12339 ( .A1(n10305), .A2(n9796), .ZN(n9785) );
  AND2_X1 U12340 ( .A1(n9799), .A2(n9785), .ZN(n9786) );
  NAND2_X1 U12341 ( .A1(n9787), .A2(n9786), .ZN(n10365) );
  OAI22_X1 U12342 ( .A1(n13091), .A2(n13448), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8750), .ZN(n9792) );
  INV_X1 U12343 ( .A(n13046), .ZN(n13072) );
  INV_X1 U12344 ( .A(n13442), .ZN(n12064) );
  NAND2_X1 U12345 ( .A1(n13089), .A2(n13444), .ZN(n13039) );
  OAI22_X1 U12346 ( .A1(n13072), .A2(n12064), .B1(n12059), .B2(n13039), .ZN(
        n9791) );
  OR4_X1 U12347 ( .A1(n9794), .A2(n9793), .A3(n9792), .A4(n9791), .ZN(P2_U3206) );
  OAI21_X1 U12348 ( .B1(n9799), .B2(n9796), .A(n9795), .ZN(n9801) );
  INV_X1 U12349 ( .A(n9797), .ZN(n9798) );
  NAND2_X1 U12350 ( .A1(n9799), .A2(n9798), .ZN(n9800) );
  NAND2_X1 U12351 ( .A1(n9801), .A2(n9800), .ZN(n9817) );
  AND2_X1 U12352 ( .A1(n9817), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14762) );
  INV_X1 U12353 ( .A(n14762), .ZN(n14848) );
  NOR2_X1 U12354 ( .A1(n9802), .A2(n14848), .ZN(n9822) );
  INV_X1 U12355 ( .A(n9817), .ZN(n9804) );
  NOR2_X1 U12356 ( .A1(n9159), .A2(P2_U3088), .ZN(n9803) );
  INV_X1 U12357 ( .A(n9812), .ZN(n9805) );
  NOR2_X2 U12358 ( .A1(n9805), .A2(n13579), .ZN(n14838) );
  INV_X1 U12359 ( .A(n14838), .ZN(n13176) );
  XNOR2_X1 U12360 ( .A(n10079), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n9807) );
  AND2_X1 U12361 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9806) );
  NAND2_X1 U12362 ( .A1(n9807), .A2(n9806), .ZN(n10096) );
  INV_X1 U12363 ( .A(n10096), .ZN(n9809) );
  AOI21_X1 U12364 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(P2_REG2_REG_0__SCAN_IN), 
        .A(n9807), .ZN(n9808) );
  NOR3_X1 U12365 ( .A1(n13176), .A2(n9809), .A3(n9808), .ZN(n9821) );
  NAND2_X1 U12366 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9815) );
  XNOR2_X1 U12367 ( .A(n10079), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9811) );
  INV_X1 U12368 ( .A(n9811), .ZN(n9814) );
  INV_X1 U12369 ( .A(n9815), .ZN(n9810) );
  NAND2_X1 U12370 ( .A1(n9811), .A2(n9810), .ZN(n10081) );
  INV_X1 U12371 ( .A(n10081), .ZN(n9813) );
  NAND2_X1 U12372 ( .A1(n9812), .A2(n13579), .ZN(n14844) );
  AOI211_X1 U12373 ( .C1(n9815), .C2(n9814), .A(n9813), .B(n14844), .ZN(n9820)
         );
  NAND2_X1 U12374 ( .A1(n9159), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9816) );
  OR2_X1 U12375 ( .A1(n9817), .A2(n9816), .ZN(n14794) );
  OAI22_X1 U12376 ( .A1(n14794), .A2(n10079), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9818), .ZN(n9819) );
  OR4_X1 U12377 ( .A1(n9822), .A2(n9821), .A3(n9820), .A4(n9819), .ZN(P2_U3215) );
  NAND2_X2 U12378 ( .A1(n6439), .A2(P2_U3088), .ZN(n13588) );
  INV_X2 U12379 ( .A(n13577), .ZN(n13590) );
  OAI222_X1 U12380 ( .A1(n13588), .A2(n9823), .B1(n13590), .B2(n9836), .C1(
        n10079), .C2(P2_U3088), .ZN(P2_U3326) );
  OAI222_X1 U12381 ( .A1(P2_U3088), .A2(n14766), .B1(n13590), .B2(n9838), .C1(
        n9824), .C2(n13588), .ZN(P2_U3325) );
  INV_X1 U12382 ( .A(n13588), .ZN(n9839) );
  OAI222_X1 U12383 ( .A1(n13588), .A2(n9825), .B1(n13590), .B2(n9834), .C1(
        n14775), .C2(P2_U3088), .ZN(P2_U3324) );
  NOR2_X2 U12384 ( .A1(n9833), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14388) );
  INV_X1 U12385 ( .A(n14388), .ZN(n14378) );
  OAI222_X1 U12386 ( .A1(n14378), .A2(n9826), .B1(n14376), .B2(n6718), .C1(
        P3_U3151), .C2(n6433), .ZN(P3_U3294) );
  OAI222_X1 U12387 ( .A1(n14378), .A2(n9827), .B1(n14376), .B2(n15221), .C1(
        P3_U3151), .C2(n11076), .ZN(P3_U3287) );
  OAI222_X1 U12388 ( .A1(n13588), .A2(n9828), .B1(n13590), .B2(n9844), .C1(
        n14793), .C2(P2_U3088), .ZN(P2_U3323) );
  OAI222_X1 U12389 ( .A1(P3_U3151), .A2(n10179), .B1(n14378), .B2(n9832), .C1(
        n9831), .C2(n14376), .ZN(P3_U3295) );
  NAND2_X2 U12390 ( .A1(n9479), .A2(P1_U3086), .ZN(n14353) );
  OAI222_X1 U12391 ( .A1(n14353), .A2(n9835), .B1(n13906), .B2(P1_U3086), .C1(
        n11585), .C2(n9834), .ZN(P1_U3352) );
  OAI222_X1 U12392 ( .A1(n14353), .A2(n9837), .B1(n10033), .B2(P1_U3086), .C1(
        n11585), .C2(n9836), .ZN(P1_U3354) );
  OAI222_X1 U12393 ( .A1(n14353), .A2(n8347), .B1(n13890), .B2(P1_U3086), .C1(
        n11585), .C2(n9838), .ZN(P1_U3353) );
  AOI22_X1 U12394 ( .A1(n14808), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n9839), .ZN(n9840) );
  OAI21_X1 U12395 ( .B1(n9841), .B2(n13590), .A(n9840), .ZN(P2_U3322) );
  INV_X1 U12396 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9843) );
  INV_X1 U12397 ( .A(n13941), .ZN(n9842) );
  OAI222_X1 U12398 ( .A1(n14353), .A2(n9843), .B1(n9842), .B2(P1_U3086), .C1(
        n11585), .C2(n9841), .ZN(P1_U3350) );
  INV_X2 U12399 ( .A(n14341), .ZN(n11585) );
  OAI222_X1 U12400 ( .A1(n11585), .A2(n9844), .B1(n13928), .B2(P1_U3086), .C1(
        n6901), .C2(n14353), .ZN(P1_U3351) );
  INV_X1 U12401 ( .A(n14376), .ZN(n14387) );
  AOI222_X1 U12402 ( .A1(n9845), .A2(n14388), .B1(SI_10_), .B2(n14387), .C1(
        n15018), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9846) );
  INV_X1 U12403 ( .A(n9846), .ZN(P3_U3285) );
  AOI222_X1 U12404 ( .A1(n9847), .A2(n14388), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10379), .C1(SI_4_), .C2(n14387), .ZN(n9848) );
  INV_X1 U12405 ( .A(n9848), .ZN(P3_U3291) );
  AOI222_X1 U12406 ( .A1(n9849), .A2(n14388), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10278), .C1(SI_2_), .C2(n14387), .ZN(n9850) );
  INV_X1 U12407 ( .A(n9850), .ZN(P3_U3293) );
  AOI222_X1 U12408 ( .A1(n9851), .A2(n14388), .B1(n10779), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_7_), .C2(n14387), .ZN(n9852) );
  INV_X1 U12409 ( .A(n9852), .ZN(P3_U3288) );
  AOI222_X1 U12410 ( .A1(n9853), .A2(n14388), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10317), .C1(SI_3_), .C2(n14387), .ZN(n9854) );
  INV_X1 U12411 ( .A(n9854), .ZN(P3_U3292) );
  AOI222_X1 U12412 ( .A1(n9855), .A2(n14388), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10471), .C1(SI_5_), .C2(n14387), .ZN(n9856) );
  INV_X1 U12413 ( .A(n9856), .ZN(P3_U3290) );
  OAI222_X1 U12414 ( .A1(n11585), .A2(n9859), .B1(n13951), .B2(P1_U3086), .C1(
        n9857), .C2(n14353), .ZN(P1_U3349) );
  INV_X1 U12415 ( .A(n13124), .ZN(n9858) );
  OAI222_X1 U12416 ( .A1(n13588), .A2(n9860), .B1(n13590), .B2(n9859), .C1(
        n9858), .C2(P2_U3088), .ZN(P2_U3321) );
  OAI222_X1 U12417 ( .A1(P3_U3151), .A2(n11478), .B1(n14376), .B2(n9862), .C1(
        n14378), .C2(n9861), .ZN(P3_U3283) );
  NAND2_X1 U12418 ( .A1(n10149), .A2(n9865), .ZN(n9864) );
  AND2_X1 U12419 ( .A1(n9864), .A2(n9863), .ZN(n9950) );
  INV_X1 U12420 ( .A(n9950), .ZN(n9867) );
  INV_X1 U12421 ( .A(n9865), .ZN(n9866) );
  NAND2_X1 U12422 ( .A1(n9866), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12043) );
  NAND2_X1 U12423 ( .A1(n10155), .A2(n12043), .ZN(n9949) );
  AND2_X1 U12424 ( .A1(n9867), .A2(n9949), .ZN(n14594) );
  NOR2_X1 U12425 ( .A1(n14594), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12426 ( .A(n9868), .ZN(n9871) );
  INV_X1 U12427 ( .A(n14353), .ZN(n9885) );
  AOI22_X1 U12428 ( .A1(n13970), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9885), .ZN(n9869) );
  OAI21_X1 U12429 ( .B1(n9871), .B2(n11585), .A(n9869), .ZN(P1_U3348) );
  INV_X1 U12430 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9872) );
  INV_X1 U12431 ( .A(n13136), .ZN(n9870) );
  OAI222_X1 U12432 ( .A1(n13588), .A2(n9872), .B1(n13590), .B2(n9871), .C1(
        P2_U3088), .C2(n9870), .ZN(P2_U3320) );
  INV_X1 U12433 ( .A(n9873), .ZN(n9875) );
  AOI22_X1 U12434 ( .A1(n9991), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9885), .ZN(n9874) );
  OAI21_X1 U12435 ( .B1(n9875), .B2(n11585), .A(n9874), .ZN(P1_U3347) );
  INV_X1 U12436 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9876) );
  OAI222_X1 U12437 ( .A1(n13588), .A2(n9876), .B1(n13590), .B2(n9875), .C1(
        P2_U3088), .C2(n10109), .ZN(P2_U3319) );
  INV_X1 U12438 ( .A(n9877), .ZN(n9878) );
  NOR2_X4 U12439 ( .A1(n10155), .A2(n9878), .ZN(n14684) );
  OAI22_X1 U12440 ( .A1(n14684), .A2(P1_D_REG_0__SCAN_IN), .B1(n9882), .B2(
        n9879), .ZN(n9880) );
  INV_X1 U12441 ( .A(n9880), .ZN(P1_U3445) );
  OAI22_X1 U12442 ( .A1(n14684), .A2(P1_D_REG_1__SCAN_IN), .B1(n9882), .B2(
        n9881), .ZN(n9883) );
  INV_X1 U12443 ( .A(n9883), .ZN(P1_U3446) );
  INV_X1 U12444 ( .A(n9884), .ZN(n9887) );
  AOI22_X1 U12445 ( .A1(n10014), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9885), .ZN(n9886) );
  OAI21_X1 U12446 ( .B1(n9887), .B2(n11585), .A(n9886), .ZN(P1_U3346) );
  INV_X1 U12447 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9888) );
  INV_X1 U12448 ( .A(n14839), .ZN(n10112) );
  OAI222_X1 U12449 ( .A1(n13588), .A2(n9888), .B1(n13590), .B2(n9887), .C1(
        P2_U3088), .C2(n10112), .ZN(P2_U3318) );
  OAI222_X1 U12450 ( .A1(n12368), .A2(P3_U3151), .B1(n14378), .B2(n9890), .C1(
        n9889), .C2(n14376), .ZN(P3_U3281) );
  NOR2_X1 U12451 ( .A1(n9891), .A2(n12848), .ZN(n9893) );
  INV_X1 U12452 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9892) );
  NOR2_X1 U12453 ( .A1(n9921), .A2(n9892), .ZN(P3_U3239) );
  CLKBUF_X1 U12454 ( .A(n9893), .Z(n9921) );
  INV_X1 U12455 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9894) );
  NOR2_X1 U12456 ( .A1(n9921), .A2(n9894), .ZN(P3_U3247) );
  INV_X1 U12457 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9895) );
  NOR2_X1 U12458 ( .A1(n9893), .A2(n9895), .ZN(P3_U3242) );
  INV_X1 U12459 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9896) );
  NOR2_X1 U12460 ( .A1(n9921), .A2(n9896), .ZN(P3_U3253) );
  INV_X1 U12461 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9897) );
  NOR2_X1 U12462 ( .A1(n9893), .A2(n9897), .ZN(P3_U3243) );
  INV_X1 U12463 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9898) );
  NOR2_X1 U12464 ( .A1(n9893), .A2(n9898), .ZN(P3_U3245) );
  INV_X1 U12465 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9899) );
  NOR2_X1 U12466 ( .A1(n9921), .A2(n9899), .ZN(P3_U3246) );
  INV_X1 U12467 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9900) );
  NOR2_X1 U12468 ( .A1(n9921), .A2(n9900), .ZN(P3_U3249) );
  INV_X1 U12469 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9901) );
  NOR2_X1 U12470 ( .A1(n9921), .A2(n9901), .ZN(P3_U3248) );
  INV_X1 U12471 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9902) );
  NOR2_X1 U12472 ( .A1(n9921), .A2(n9902), .ZN(P3_U3254) );
  INV_X1 U12473 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9903) );
  NOR2_X1 U12474 ( .A1(n9893), .A2(n9903), .ZN(P3_U3235) );
  INV_X1 U12475 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9904) );
  NOR2_X1 U12476 ( .A1(n9893), .A2(n9904), .ZN(P3_U3240) );
  INV_X1 U12477 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9905) );
  NOR2_X1 U12478 ( .A1(n9893), .A2(n9905), .ZN(P3_U3241) );
  INV_X1 U12479 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9906) );
  NOR2_X1 U12480 ( .A1(n9921), .A2(n9906), .ZN(P3_U3261) );
  INV_X1 U12481 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n15254) );
  NOR2_X1 U12482 ( .A1(n9893), .A2(n15254), .ZN(P3_U3260) );
  INV_X1 U12483 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U12484 ( .A1(n9893), .A2(n9907), .ZN(P3_U3244) );
  INV_X1 U12485 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U12486 ( .A1(n9893), .A2(n9908), .ZN(P3_U3258) );
  INV_X1 U12487 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9909) );
  NOR2_X1 U12488 ( .A1(n9893), .A2(n9909), .ZN(P3_U3234) );
  INV_X1 U12489 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9910) );
  NOR2_X1 U12490 ( .A1(n9921), .A2(n9910), .ZN(P3_U3256) );
  INV_X1 U12491 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9911) );
  NOR2_X1 U12492 ( .A1(n9921), .A2(n9911), .ZN(P3_U3255) );
  INV_X1 U12493 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n15256) );
  NOR2_X1 U12494 ( .A1(n9921), .A2(n15256), .ZN(P3_U3251) );
  INV_X1 U12495 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U12496 ( .A1(n9921), .A2(n9912), .ZN(P3_U3250) );
  INV_X1 U12497 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9913) );
  NOR2_X1 U12498 ( .A1(n9921), .A2(n9913), .ZN(P3_U3252) );
  INV_X1 U12499 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9914) );
  NOR2_X1 U12500 ( .A1(n9893), .A2(n9914), .ZN(P3_U3236) );
  INV_X1 U12501 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9915) );
  NOR2_X1 U12502 ( .A1(n9921), .A2(n9915), .ZN(P3_U3237) );
  INV_X1 U12503 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9916) );
  NOR2_X1 U12504 ( .A1(n9921), .A2(n9916), .ZN(P3_U3257) );
  INV_X1 U12505 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U12506 ( .A1(n9921), .A2(n9917), .ZN(P3_U3238) );
  INV_X1 U12507 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U12508 ( .A1(n9921), .A2(n9918), .ZN(P3_U3263) );
  INV_X1 U12509 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9919) );
  NOR2_X1 U12510 ( .A1(n9921), .A2(n9919), .ZN(P3_U3262) );
  INV_X1 U12511 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U12512 ( .A1(n9921), .A2(n9920), .ZN(P3_U3259) );
  INV_X1 U12513 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9924) );
  INV_X1 U12514 ( .A(n9922), .ZN(n9925) );
  INV_X1 U12515 ( .A(n10134), .ZN(n9923) );
  OAI222_X1 U12516 ( .A1(n13588), .A2(n9924), .B1(n13590), .B2(n9925), .C1(
        P2_U3088), .C2(n9923), .ZN(P2_U3317) );
  INV_X1 U12517 ( .A(n10041), .ZN(n10023) );
  OAI222_X1 U12518 ( .A1(n14353), .A2(n9926), .B1(n11585), .B2(n9925), .C1(
        P1_U3086), .C2(n10023), .ZN(P1_U3345) );
  MUX2_X1 U12519 ( .A(n9927), .B(P1_REG1_REG_8__SCAN_IN), .S(n9991), .Z(n9948)
         );
  MUX2_X1 U12520 ( .A(n9928), .B(P1_REG1_REG_4__SCAN_IN), .S(n13928), .Z(n9938) );
  MUX2_X1 U12521 ( .A(n9929), .B(P1_REG1_REG_1__SCAN_IN), .S(n10033), .Z(n9931) );
  AND2_X1 U12522 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9930) );
  NAND2_X1 U12523 ( .A1(n9931), .A2(n9930), .ZN(n13888) );
  INV_X1 U12524 ( .A(n10033), .ZN(n9957) );
  NAND2_X1 U12525 ( .A1(n9957), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n13887) );
  NAND2_X1 U12526 ( .A1(n13888), .A2(n13887), .ZN(n9933) );
  MUX2_X1 U12527 ( .A(n9934), .B(P1_REG1_REG_2__SCAN_IN), .S(n13890), .Z(n9932) );
  NAND2_X1 U12528 ( .A1(n9933), .A2(n9932), .ZN(n13910) );
  OR2_X1 U12529 ( .A1(n13890), .A2(n9934), .ZN(n13909) );
  NAND2_X1 U12530 ( .A1(n13910), .A2(n13909), .ZN(n9936) );
  MUX2_X1 U12531 ( .A(n13907), .B(P1_REG1_REG_3__SCAN_IN), .S(n13906), .Z(
        n9935) );
  NAND2_X1 U12532 ( .A1(n9936), .A2(n9935), .ZN(n13916) );
  OR2_X1 U12533 ( .A1(n13906), .A2(n13907), .ZN(n13915) );
  NAND2_X1 U12534 ( .A1(n13916), .A2(n13915), .ZN(n9937) );
  NAND2_X1 U12535 ( .A1(n9938), .A2(n9937), .ZN(n13919) );
  INV_X1 U12536 ( .A(n13928), .ZN(n9965) );
  NAND2_X1 U12537 ( .A1(n9965), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9939) );
  AND2_X1 U12538 ( .A1(n13919), .A2(n9939), .ZN(n13938) );
  MUX2_X1 U12539 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9255), .S(n13941), .Z(
        n13939) );
  NAND2_X1 U12540 ( .A1(n13938), .A2(n13939), .ZN(n13937) );
  OR2_X1 U12541 ( .A1(n13941), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9940) );
  AND2_X1 U12542 ( .A1(n13937), .A2(n9940), .ZN(n13957) );
  MUX2_X1 U12543 ( .A(n9941), .B(P1_REG1_REG_6__SCAN_IN), .S(n13951), .Z(
        n13956) );
  NAND2_X1 U12544 ( .A1(n13957), .A2(n13956), .ZN(n13967) );
  NAND2_X1 U12545 ( .A1(n9971), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U12546 ( .A1(n13967), .A2(n13966), .ZN(n9944) );
  MUX2_X1 U12547 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9942), .S(n13970), .Z(n9943) );
  NAND2_X1 U12548 ( .A1(n9944), .A2(n9943), .ZN(n13969) );
  NAND2_X1 U12549 ( .A1(n13970), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9945) );
  NAND2_X1 U12550 ( .A1(n13969), .A2(n9945), .ZN(n9947) );
  OR2_X1 U12551 ( .A1(n9947), .A2(n9948), .ZN(n9987) );
  INV_X1 U12552 ( .A(n9987), .ZN(n9946) );
  AOI21_X1 U12553 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(n9982) );
  NAND2_X1 U12554 ( .A1(n9950), .A2(n9949), .ZN(n14596) );
  INV_X1 U12555 ( .A(n6440), .ZN(n12039) );
  OR2_X1 U12556 ( .A1(n14596), .A2(n12039), .ZN(n13926) );
  NOR2_X1 U12557 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9299), .ZN(n9953) );
  INV_X1 U12558 ( .A(n9991), .ZN(n9951) );
  NOR2_X1 U12559 ( .A1(n14602), .A2(n9951), .ZN(n9952) );
  AOI211_X1 U12560 ( .C1(n14594), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9953), .B(
        n9952), .ZN(n9981) );
  OR3_X1 U12561 ( .A1(n14596), .A2(n6440), .A3(n14344), .ZN(n14604) );
  MUX2_X1 U12562 ( .A(n9954), .B(P1_REG2_REG_4__SCAN_IN), .S(n13928), .Z(n9964) );
  MUX2_X1 U12563 ( .A(n9955), .B(P1_REG2_REG_1__SCAN_IN), .S(n10033), .Z(n9956) );
  AND2_X1 U12564 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10024) );
  NAND2_X1 U12565 ( .A1(n9956), .A2(n10024), .ZN(n13893) );
  NAND2_X1 U12566 ( .A1(n9957), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n13892) );
  NAND2_X1 U12567 ( .A1(n13893), .A2(n13892), .ZN(n9959) );
  MUX2_X1 U12568 ( .A(n9960), .B(P1_REG2_REG_2__SCAN_IN), .S(n13890), .Z(n9958) );
  NAND2_X1 U12569 ( .A1(n9959), .A2(n9958), .ZN(n13904) );
  OR2_X1 U12570 ( .A1(n13890), .A2(n9960), .ZN(n13903) );
  NAND2_X1 U12571 ( .A1(n13904), .A2(n13903), .ZN(n9962) );
  MUX2_X1 U12572 ( .A(n10742), .B(P1_REG2_REG_3__SCAN_IN), .S(n13906), .Z(
        n9961) );
  NAND2_X1 U12573 ( .A1(n9962), .A2(n9961), .ZN(n13921) );
  OR2_X1 U12574 ( .A1(n13906), .A2(n10742), .ZN(n13920) );
  NAND2_X1 U12575 ( .A1(n13921), .A2(n13920), .ZN(n9963) );
  NAND2_X1 U12576 ( .A1(n9964), .A2(n9963), .ZN(n13944) );
  NAND2_X1 U12577 ( .A1(n9965), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13943) );
  NAND2_X1 U12578 ( .A1(n13944), .A2(n13943), .ZN(n9967) );
  MUX2_X1 U12579 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10643), .S(n13941), .Z(
        n9966) );
  NAND2_X1 U12580 ( .A1(n9967), .A2(n9966), .ZN(n13953) );
  NAND2_X1 U12581 ( .A1(n13941), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n13952) );
  NAND2_X1 U12582 ( .A1(n13953), .A2(n13952), .ZN(n9970) );
  MUX2_X1 U12583 ( .A(n9968), .B(P1_REG2_REG_6__SCAN_IN), .S(n13951), .Z(n9969) );
  NAND2_X1 U12584 ( .A1(n9970), .A2(n9969), .ZN(n13973) );
  NAND2_X1 U12585 ( .A1(n9971), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n13972) );
  NAND2_X1 U12586 ( .A1(n13973), .A2(n13972), .ZN(n9973) );
  MUX2_X1 U12587 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10805), .S(n13970), .Z(
        n9972) );
  NAND2_X1 U12588 ( .A1(n9973), .A2(n9972), .ZN(n13975) );
  NAND2_X1 U12589 ( .A1(n13970), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9978) );
  NAND2_X1 U12590 ( .A1(n13975), .A2(n9978), .ZN(n9976) );
  MUX2_X1 U12591 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9974), .S(n9991), .Z(n9975)
         );
  NAND2_X1 U12592 ( .A1(n9976), .A2(n9975), .ZN(n9997) );
  MUX2_X1 U12593 ( .A(n9974), .B(P1_REG2_REG_8__SCAN_IN), .S(n9991), .Z(n9977)
         );
  NAND3_X1 U12594 ( .A1(n13975), .A2(n9978), .A3(n9977), .ZN(n9979) );
  NAND3_X1 U12595 ( .A1(n13976), .A2(n9997), .A3(n9979), .ZN(n9980) );
  OAI211_X1 U12596 ( .C1(n9982), .C2(n13926), .A(n9981), .B(n9980), .ZN(
        P1_U3251) );
  OR2_X1 U12597 ( .A1(n9991), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U12598 ( .A1(n9987), .A2(n9985), .ZN(n9983) );
  MUX2_X1 U12599 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9315), .S(n10014), .Z(n9984) );
  NAND2_X1 U12600 ( .A1(n9983), .A2(n9984), .ZN(n10008) );
  INV_X1 U12601 ( .A(n9984), .ZN(n9986) );
  NAND3_X1 U12602 ( .A1(n9987), .A2(n9986), .A3(n9985), .ZN(n9988) );
  AND2_X1 U12603 ( .A1(n10008), .A2(n9988), .ZN(n10001) );
  INV_X1 U12604 ( .A(n14602), .ZN(n13964) );
  INV_X1 U12605 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U12606 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11280) );
  OAI21_X1 U12607 ( .B1(n14611), .B2(n9989), .A(n11280), .ZN(n9990) );
  AOI21_X1 U12608 ( .B1(n10014), .B2(n13964), .A(n9990), .ZN(n10000) );
  NAND2_X1 U12609 ( .A1(n9991), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U12610 ( .A1(n9997), .A2(n9996), .ZN(n9994) );
  MUX2_X1 U12611 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9992), .S(n10014), .Z(n9993) );
  NAND2_X1 U12612 ( .A1(n9994), .A2(n9993), .ZN(n10019) );
  MUX2_X1 U12613 ( .A(n9992), .B(P1_REG2_REG_9__SCAN_IN), .S(n10014), .Z(n9995) );
  NAND3_X1 U12614 ( .A1(n9997), .A2(n9996), .A3(n9995), .ZN(n9998) );
  NAND3_X1 U12615 ( .A1(n13976), .A2(n10019), .A3(n9998), .ZN(n9999) );
  OAI211_X1 U12616 ( .C1(n10001), .C2(n13926), .A(n10000), .B(n9999), .ZN(
        P1_U3252) );
  INV_X1 U12617 ( .A(n10002), .ZN(n10006) );
  INV_X1 U12618 ( .A(n10058), .ZN(n10003) );
  OAI222_X1 U12619 ( .A1(n14353), .A2(n10004), .B1(n11585), .B2(n10006), .C1(
        P1_U3086), .C2(n10003), .ZN(P1_U3344) );
  INV_X1 U12620 ( .A(n10211), .ZN(n10005) );
  OAI222_X1 U12621 ( .A1(n13588), .A2(n15222), .B1(n13590), .B2(n10006), .C1(
        P2_U3088), .C2(n10005), .ZN(P2_U3316) );
  AND2_X1 U12622 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11360) );
  OR2_X1 U12623 ( .A1(n10014), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U12624 ( .A1(n10008), .A2(n10007), .ZN(n10010) );
  MUX2_X1 U12625 ( .A(n9330), .B(P1_REG1_REG_10__SCAN_IN), .S(n10041), .Z(
        n10009) );
  AOI21_X1 U12626 ( .B1(n10010), .B2(n10009), .A(n13926), .ZN(n10011) );
  OR2_X1 U12627 ( .A1(n10010), .A2(n10009), .ZN(n10036) );
  NAND2_X1 U12628 ( .A1(n10011), .A2(n10036), .ZN(n10012) );
  OAI21_X1 U12629 ( .B1(n15228), .B2(n14611), .A(n10012), .ZN(n10013) );
  NOR2_X1 U12630 ( .A1(n11360), .A2(n10013), .ZN(n10022) );
  NAND2_X1 U12631 ( .A1(n10014), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10018) );
  NAND2_X1 U12632 ( .A1(n10019), .A2(n10018), .ZN(n10016) );
  MUX2_X1 U12633 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11179), .S(n10041), .Z(
        n10015) );
  NAND2_X1 U12634 ( .A1(n10016), .A2(n10015), .ZN(n10047) );
  MUX2_X1 U12635 ( .A(n11179), .B(P1_REG2_REG_10__SCAN_IN), .S(n10041), .Z(
        n10017) );
  NAND3_X1 U12636 ( .A1(n10019), .A2(n10018), .A3(n10017), .ZN(n10020) );
  NAND3_X1 U12637 ( .A1(n13976), .A2(n10047), .A3(n10020), .ZN(n10021) );
  OAI211_X1 U12638 ( .C1(n14602), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        P1_U3253) );
  INV_X1 U12639 ( .A(n10024), .ZN(n13876) );
  MUX2_X1 U12640 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9955), .S(n10033), .Z(
        n10026) );
  INV_X1 U12641 ( .A(n13893), .ZN(n10025) );
  AOI211_X1 U12642 ( .C1(n13876), .C2(n10026), .A(n10025), .B(n14604), .ZN(
        n10030) );
  MUX2_X1 U12643 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9929), .S(n10033), .Z(
        n10027) );
  OAI21_X1 U12644 ( .B1(n14592), .B2(n13879), .A(n10027), .ZN(n10028) );
  AND3_X1 U12645 ( .A1(n14607), .A2(n13888), .A3(n10028), .ZN(n10029) );
  NOR2_X1 U12646 ( .A1(n10030), .A2(n10029), .ZN(n10032) );
  AOI22_X1 U12647 ( .A1(n14594), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10031) );
  OAI211_X1 U12648 ( .C1(n10033), .C2(n14602), .A(n10032), .B(n10031), .ZN(
        P1_U3244) );
  MUX2_X1 U12649 ( .A(n10034), .B(P1_REG1_REG_11__SCAN_IN), .S(n10058), .Z(
        n10038) );
  NAND2_X1 U12650 ( .A1(n10041), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10035) );
  NAND2_X1 U12651 ( .A1(n10036), .A2(n10035), .ZN(n10037) );
  NOR2_X1 U12652 ( .A1(n10037), .A2(n10038), .ZN(n10061) );
  AOI21_X1 U12653 ( .B1(n10038), .B2(n10037), .A(n10061), .ZN(n10051) );
  NAND2_X1 U12654 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14534)
         );
  OAI21_X1 U12655 ( .B1(n14611), .B2(n10039), .A(n14534), .ZN(n10040) );
  AOI21_X1 U12656 ( .B1(n10058), .B2(n13964), .A(n10040), .ZN(n10050) );
  NAND2_X1 U12657 ( .A1(n10041), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10046) );
  NAND2_X1 U12658 ( .A1(n10047), .A2(n10046), .ZN(n10044) );
  MUX2_X1 U12659 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10042), .S(n10058), .Z(
        n10043) );
  NAND2_X1 U12660 ( .A1(n10044), .A2(n10043), .ZN(n10054) );
  MUX2_X1 U12661 ( .A(n10042), .B(P1_REG2_REG_11__SCAN_IN), .S(n10058), .Z(
        n10045) );
  NAND3_X1 U12662 ( .A1(n10047), .A2(n10046), .A3(n10045), .ZN(n10048) );
  NAND3_X1 U12663 ( .A1(n10054), .A2(n13976), .A3(n10048), .ZN(n10049) );
  OAI211_X1 U12664 ( .C1(n10051), .C2(n13926), .A(n10050), .B(n10049), .ZN(
        P1_U3254) );
  MUX2_X1 U12665 ( .A(n10052), .B(P1_REG2_REG_12__SCAN_IN), .S(n10229), .Z(
        n10057) );
  NAND2_X1 U12666 ( .A1(n10058), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U12667 ( .A1(n10054), .A2(n10053), .ZN(n10056) );
  OR2_X1 U12668 ( .A1(n10056), .A2(n10057), .ZN(n10231) );
  INV_X1 U12669 ( .A(n10231), .ZN(n10055) );
  AOI21_X1 U12670 ( .B1(n10057), .B2(n10056), .A(n10055), .ZN(n10068) );
  NOR2_X1 U12671 ( .A1(n10058), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10059) );
  INV_X1 U12672 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14424) );
  MUX2_X1 U12673 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n14424), .S(n10229), .Z(
        n10060) );
  OAI21_X1 U12674 ( .B1(n10061), .B2(n10059), .A(n10060), .ZN(n10225) );
  INV_X1 U12675 ( .A(n10225), .ZN(n10063) );
  NOR3_X1 U12676 ( .A1(n10061), .A2(n10060), .A3(n10059), .ZN(n10062) );
  OAI21_X1 U12677 ( .B1(n10063), .B2(n10062), .A(n14607), .ZN(n10067) );
  INV_X1 U12678 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11567) );
  NOR2_X1 U12679 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11567), .ZN(n10065) );
  INV_X1 U12680 ( .A(n10229), .ZN(n10073) );
  NOR2_X1 U12681 ( .A1(n14602), .A2(n10073), .ZN(n10064) );
  AOI211_X1 U12682 ( .C1(n14594), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n10065), 
        .B(n10064), .ZN(n10066) );
  OAI211_X1 U12683 ( .C1(n10068), .C2(n14604), .A(n10067), .B(n10066), .ZN(
        P1_U3255) );
  INV_X1 U12684 ( .A(n12449), .ZN(n12433) );
  INV_X1 U12685 ( .A(n10069), .ZN(n10071) );
  OAI222_X1 U12686 ( .A1(n12433), .A2(P3_U3151), .B1(n14378), .B2(n10071), 
        .C1(n10070), .C2(n14376), .ZN(P3_U3279) );
  INV_X1 U12687 ( .A(n10072), .ZN(n10075) );
  OAI222_X1 U12688 ( .A1(n14353), .A2(n10074), .B1(n11585), .B2(n10075), .C1(
        P1_U3086), .C2(n10073), .ZN(P1_U3343) );
  INV_X1 U12689 ( .A(n10408), .ZN(n10411) );
  OAI222_X1 U12690 ( .A1(n13588), .A2(n10076), .B1(n13590), .B2(n10075), .C1(
        P2_U3088), .C2(n10411), .ZN(P2_U3315) );
  OAI222_X1 U12691 ( .A1(P3_U3151), .A2(n12450), .B1(n14376), .B2(n10078), 
        .C1(n14378), .C2(n10077), .ZN(P3_U3278) );
  MUX2_X1 U12692 ( .A(n14972), .B(P2_REG1_REG_10__SCAN_IN), .S(n10134), .Z(
        n10093) );
  INV_X1 U12693 ( .A(n10079), .ZN(n10094) );
  NAND2_X1 U12694 ( .A1(n10094), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10080) );
  NAND2_X1 U12695 ( .A1(n10081), .A2(n10080), .ZN(n14764) );
  XNOR2_X1 U12696 ( .A(n14766), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n14765) );
  NAND2_X1 U12697 ( .A1(n14764), .A2(n14765), .ZN(n14763) );
  OR2_X1 U12698 ( .A1(n14766), .A2(n10082), .ZN(n10083) );
  NAND2_X1 U12699 ( .A1(n14763), .A2(n10083), .ZN(n14777) );
  XNOR2_X1 U12700 ( .A(n14775), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n14778) );
  NAND2_X1 U12701 ( .A1(n14777), .A2(n14778), .ZN(n14776) );
  OR2_X1 U12702 ( .A1(n14775), .A2(n10084), .ZN(n10085) );
  NAND2_X1 U12703 ( .A1(n14776), .A2(n10085), .ZN(n14789) );
  XNOR2_X1 U12704 ( .A(n14793), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n14790) );
  NAND2_X1 U12705 ( .A1(n14789), .A2(n14790), .ZN(n14788) );
  INV_X1 U12706 ( .A(n14793), .ZN(n10100) );
  NAND2_X1 U12707 ( .A1(n10100), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10086) );
  NAND2_X1 U12708 ( .A1(n14788), .A2(n10086), .ZN(n14803) );
  XNOR2_X1 U12709 ( .A(n14808), .B(n10087), .ZN(n14804) );
  NAND2_X1 U12710 ( .A1(n14803), .A2(n14804), .ZN(n14802) );
  NAND2_X1 U12711 ( .A1(n14808), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10088) );
  NAND2_X1 U12712 ( .A1(n14802), .A2(n10088), .ZN(n13120) );
  INV_X1 U12713 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14967) );
  MUX2_X1 U12714 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n14967), .S(n13124), .Z(
        n13121) );
  NAND2_X1 U12715 ( .A1(n13120), .A2(n13121), .ZN(n13119) );
  NAND2_X1 U12716 ( .A1(n13124), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U12717 ( .A1(n13119), .A2(n10089), .ZN(n13133) );
  INV_X1 U12718 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10873) );
  MUX2_X1 U12719 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10873), .S(n13136), .Z(
        n13134) );
  NAND2_X1 U12720 ( .A1(n13133), .A2(n13134), .ZN(n13132) );
  NAND2_X1 U12721 ( .A1(n13136), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U12722 ( .A1(n13132), .A2(n10090), .ZN(n14817) );
  INV_X1 U12723 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14969) );
  MUX2_X1 U12724 ( .A(n14969), .B(P2_REG1_REG_8__SCAN_IN), .S(n10109), .Z(
        n14818) );
  NAND2_X1 U12725 ( .A1(n14817), .A2(n14818), .ZN(n14815) );
  NAND2_X1 U12726 ( .A1(n14822), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U12727 ( .A1(n14815), .A2(n10091), .ZN(n14830) );
  MUX2_X1 U12728 ( .A(n8663), .B(P2_REG1_REG_9__SCAN_IN), .S(n14839), .Z(
        n14829) );
  NOR2_X1 U12729 ( .A1(n10092), .A2(n10093), .ZN(n10133) );
  AOI211_X1 U12730 ( .C1(n10093), .C2(n10092), .A(n14844), .B(n10133), .ZN(
        n10121) );
  INV_X1 U12731 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10097) );
  MUX2_X1 U12732 ( .A(n10097), .B(P2_REG2_REG_2__SCAN_IN), .S(n14766), .Z(
        n14770) );
  NAND2_X1 U12733 ( .A1(n10094), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U12734 ( .A1(n10096), .A2(n10095), .ZN(n14771) );
  NAND2_X1 U12735 ( .A1(n14770), .A2(n14771), .ZN(n14769) );
  OR2_X1 U12736 ( .A1(n14766), .A2(n10097), .ZN(n10098) );
  NAND2_X1 U12737 ( .A1(n14769), .A2(n10098), .ZN(n14785) );
  MUX2_X1 U12738 ( .A(n10669), .B(P2_REG2_REG_3__SCAN_IN), .S(n14775), .Z(
        n14784) );
  NAND2_X1 U12739 ( .A1(n14785), .A2(n14784), .ZN(n14783) );
  OR2_X1 U12740 ( .A1(n14775), .A2(n10669), .ZN(n10099) );
  NAND2_X1 U12741 ( .A1(n14783), .A2(n10099), .ZN(n14798) );
  MUX2_X1 U12742 ( .A(n10841), .B(P2_REG2_REG_4__SCAN_IN), .S(n14793), .Z(
        n14797) );
  NAND2_X1 U12743 ( .A1(n14798), .A2(n14797), .ZN(n14796) );
  NAND2_X1 U12744 ( .A1(n10100), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10101) );
  NAND2_X1 U12745 ( .A1(n14796), .A2(n10101), .ZN(n14811) );
  MUX2_X1 U12746 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10829), .S(n14808), .Z(
        n14810) );
  NAND2_X1 U12747 ( .A1(n14811), .A2(n14810), .ZN(n14809) );
  NAND2_X1 U12748 ( .A1(n14808), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13126) );
  NAND2_X1 U12749 ( .A1(n14809), .A2(n13126), .ZN(n10104) );
  MUX2_X1 U12750 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10102), .S(n13124), .Z(
        n10103) );
  NAND2_X1 U12751 ( .A1(n10104), .A2(n10103), .ZN(n13139) );
  NAND2_X1 U12752 ( .A1(n13124), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13138) );
  NAND2_X1 U12753 ( .A1(n13139), .A2(n13138), .ZN(n10107) );
  MUX2_X1 U12754 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10105), .S(n13136), .Z(
        n10106) );
  NAND2_X1 U12755 ( .A1(n10107), .A2(n10106), .ZN(n13141) );
  NAND2_X1 U12756 ( .A1(n13136), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10108) );
  NAND2_X1 U12757 ( .A1(n13141), .A2(n10108), .ZN(n14825) );
  MUX2_X1 U12758 ( .A(n10951), .B(P2_REG2_REG_8__SCAN_IN), .S(n10109), .Z(
        n14824) );
  NAND2_X1 U12759 ( .A1(n14825), .A2(n14824), .ZN(n14823) );
  NAND2_X1 U12760 ( .A1(n14822), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10110) );
  NAND2_X1 U12761 ( .A1(n14823), .A2(n10110), .ZN(n14834) );
  MUX2_X1 U12762 ( .A(n10111), .B(P2_REG2_REG_9__SCAN_IN), .S(n14839), .Z(
        n14833) );
  OR2_X1 U12763 ( .A1(n14834), .A2(n14833), .ZN(n14836) );
  NAND2_X1 U12764 ( .A1(n10112), .A2(n10111), .ZN(n10113) );
  NAND2_X1 U12765 ( .A1(n14836), .A2(n10113), .ZN(n10115) );
  INV_X1 U12766 ( .A(n10115), .ZN(n10117) );
  MUX2_X1 U12767 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n11162), .S(n10134), .Z(
        n10116) );
  MUX2_X1 U12768 ( .A(n11162), .B(P2_REG2_REG_10__SCAN_IN), .S(n10134), .Z(
        n10114) );
  OR2_X1 U12769 ( .A1(n10115), .A2(n10114), .ZN(n10127) );
  OAI211_X1 U12770 ( .C1(n10117), .C2(n10116), .A(n14838), .B(n10127), .ZN(
        n10119) );
  AND2_X1 U12771 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11190) );
  AOI21_X1 U12772 ( .B1(n14840), .B2(n10134), .A(n11190), .ZN(n10118) );
  OAI211_X1 U12773 ( .C1(n14848), .C2(n14398), .A(n10119), .B(n10118), .ZN(
        n10120) );
  OR2_X1 U12774 ( .A1(n10121), .A2(n10120), .ZN(P2_U3224) );
  INV_X1 U12775 ( .A(n10122), .ZN(n10124) );
  INV_X1 U12776 ( .A(n10244), .ZN(n10239) );
  OAI222_X1 U12777 ( .A1(n14353), .A2(n10123), .B1(n11585), .B2(n10124), .C1(
        P1_U3086), .C2(n10239), .ZN(P1_U3342) );
  OAI222_X1 U12778 ( .A1(n13588), .A2(n10125), .B1(n13590), .B2(n10124), .C1(
        P2_U3088), .C2(n10414), .ZN(P2_U3314) );
  NAND2_X1 U12779 ( .A1(n10134), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10126) );
  AND2_X1 U12780 ( .A1(n10127), .A2(n10126), .ZN(n10129) );
  MUX2_X1 U12781 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11388), .S(n10211), .Z(
        n10128) );
  NAND2_X1 U12782 ( .A1(n10129), .A2(n10128), .ZN(n10217) );
  OAI21_X1 U12783 ( .B1(n10129), .B2(n10128), .A(n10217), .ZN(n10139) );
  INV_X1 U12784 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U12785 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11393)
         );
  INV_X1 U12786 ( .A(n11393), .ZN(n10130) );
  AOI21_X1 U12787 ( .B1(n14840), .B2(n10211), .A(n10130), .ZN(n10131) );
  OAI21_X1 U12788 ( .B1(n14848), .B2(n10132), .A(n10131), .ZN(n10138) );
  MUX2_X1 U12789 ( .A(n13553), .B(P2_REG1_REG_11__SCAN_IN), .S(n10211), .Z(
        n10135) );
  NOR2_X1 U12790 ( .A1(n10136), .A2(n10135), .ZN(n10208) );
  AOI211_X1 U12791 ( .C1(n10136), .C2(n10135), .A(n14844), .B(n10208), .ZN(
        n10137) );
  AOI211_X1 U12792 ( .C1(n14838), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10140) );
  INV_X1 U12793 ( .A(n10140), .ZN(P2_U3225) );
  INV_X1 U12794 ( .A(n12453), .ZN(n14449) );
  OAI222_X1 U12795 ( .A1(P3_U3151), .A2(n14449), .B1(n14376), .B2(n10142), 
        .C1(n14378), .C2(n10141), .ZN(P3_U3277) );
  NAND2_X1 U12796 ( .A1(n10143), .A2(n11525), .ZN(n10760) );
  AND2_X2 U12797 ( .A1(n10146), .A2(n11823), .ZN(n10426) );
  OAI222_X1 U12798 ( .A1(n13754), .A2(n10750), .B1(n13752), .B2(n10753), .C1(
        n10146), .C2(n14592), .ZN(n10435) );
  NAND2_X1 U12799 ( .A1(n10147), .A2(n10435), .ZN(n10434) );
  OAI21_X1 U12800 ( .B1(n10147), .B2(n10435), .A(n10434), .ZN(n13875) );
  INV_X1 U12801 ( .A(n10171), .ZN(n10164) );
  NAND3_X1 U12802 ( .A1(n10164), .A2(n10148), .A3(n10163), .ZN(n10456) );
  INV_X1 U12803 ( .A(n10456), .ZN(n10157) );
  OR2_X1 U12804 ( .A1(n10155), .A2(n10149), .ZN(n10152) );
  NAND2_X1 U12805 ( .A1(n10167), .A2(n14230), .ZN(n10150) );
  NOR2_X1 U12806 ( .A1(n10152), .A2(n14723), .ZN(n10153) );
  INV_X1 U12807 ( .A(n12040), .ZN(n10154) );
  OR2_X1 U12808 ( .A1(n10456), .A2(n10154), .ZN(n11281) );
  NOR2_X1 U12809 ( .A1(n11281), .A2(n14617), .ZN(n14528) );
  AOI22_X1 U12810 ( .A1(n13875), .A2(n14532), .B1(n14528), .B2(n6936), .ZN(
        n10161) );
  INV_X1 U12811 ( .A(n10155), .ZN(n10156) );
  NAND2_X1 U12812 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  NAND2_X1 U12813 ( .A1(n10158), .A2(n14229), .ZN(n10919) );
  INV_X1 U12814 ( .A(n10458), .ZN(n10159) );
  NAND2_X1 U12815 ( .A1(n10919), .A2(n10159), .ZN(n13768) );
  AOI22_X1 U12816 ( .A1(n15311), .A2(n10896), .B1(n13768), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U12817 ( .A1(n10161), .A2(n10160), .ZN(P1_U3232) );
  NAND4_X1 U12818 ( .A1(n12040), .A2(n10163), .A3(n10162), .A4(n10455), .ZN(
        n10172) );
  INV_X1 U12819 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10170) );
  OR3_X1 U12820 ( .A1(n14357), .A2(n12018), .A3(n11525), .ZN(n14729) );
  OR2_X1 U12821 ( .A1(n13874), .A2(n10896), .ZN(n10165) );
  NAND2_X1 U12822 ( .A1(n10166), .A2(n10165), .ZN(n11988) );
  INV_X1 U12823 ( .A(n11988), .ZN(n10895) );
  AOI22_X1 U12824 ( .A1(n10895), .A2(n14403), .B1(n14404), .B2(n6936), .ZN(
        n10899) );
  NAND2_X1 U12825 ( .A1(n10896), .A2(n10167), .ZN(n10168) );
  OAI211_X1 U12826 ( .C1(n14703), .C2(n11988), .A(n10899), .B(n10168), .ZN(
        n10173) );
  NAND2_X1 U12827 ( .A1(n10173), .A2(n14751), .ZN(n10169) );
  OAI21_X1 U12828 ( .B1(n14751), .B2(n10170), .A(n10169), .ZN(P1_U3459) );
  NAND2_X1 U12829 ( .A1(n10173), .A2(n14761), .ZN(n10174) );
  OAI21_X1 U12830 ( .B1(n14761), .B2(n14592), .A(n10174), .ZN(P1_U3528) );
  NAND2_X1 U12831 ( .A1(n11748), .A2(n10177), .ZN(n10175) );
  AND2_X1 U12832 ( .A1(n10176), .A2(n10175), .ZN(n10184) );
  INV_X1 U12833 ( .A(n10358), .ZN(n10178) );
  OR2_X1 U12834 ( .A1(n10177), .A2(P3_U3151), .ZN(n11796) );
  NAND2_X1 U12835 ( .A1(n10178), .A2(n11796), .ZN(n10185) );
  NAND2_X1 U12836 ( .A1(n10184), .A2(n10185), .ZN(n10191) );
  MUX2_X1 U12837 ( .A(n12352), .B(n10191), .S(n8191), .Z(n14989) );
  OR2_X1 U12838 ( .A1(n10191), .A2(n11058), .ZN(n14976) );
  AND2_X1 U12839 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10179), .ZN(n10180) );
  OAI21_X1 U12840 ( .B1(n6433), .B2(n10180), .A(n7646), .ZN(n10182) );
  INV_X1 U12841 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10181) );
  OR2_X1 U12842 ( .A1(n10182), .A2(n10181), .ZN(n10264) );
  NAND2_X1 U12843 ( .A1(n10182), .A2(n10181), .ZN(n10183) );
  NAND2_X1 U12844 ( .A1(n10264), .A2(n10183), .ZN(n10195) );
  INV_X1 U12845 ( .A(n10184), .ZN(n10186) );
  NAND2_X1 U12846 ( .A1(n14995), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10187) );
  OAI21_X1 U12847 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n15082), .A(n10187), .ZN(
        n10194) );
  NOR2_X1 U12848 ( .A1(n10501), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10188) );
  NAND2_X1 U12849 ( .A1(n10189), .A2(n7702), .ZN(n10192) );
  AOI21_X1 U12850 ( .B1(n10259), .B2(n10192), .A(n15001), .ZN(n10193) );
  AOI211_X1 U12851 ( .C1(n15007), .C2(n10195), .A(n10194), .B(n10193), .ZN(
        n10198) );
  INV_X2 U12852 ( .A(n11058), .ZN(n11248) );
  MUX2_X1 U12853 ( .A(n10501), .B(n12053), .S(n11248), .Z(n14975) );
  AND2_X1 U12854 ( .A1(n14975), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14979) );
  XNOR2_X1 U12855 ( .A(n10258), .B(n14979), .ZN(n10196) );
  NAND2_X1 U12856 ( .A1(n10196), .A2(n15015), .ZN(n10197) );
  OAI211_X1 U12857 ( .C1(n14989), .C2(n6433), .A(n10198), .B(n10197), .ZN(
        P3_U3183) );
  INV_X1 U12858 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14960) );
  AOI22_X1 U12859 ( .A1(n14816), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n14838), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10203) );
  NAND2_X1 U12860 ( .A1(n14838), .A2(n10199), .ZN(n10200) );
  OAI211_X1 U12861 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14844), .A(n10200), .B(
        n14794), .ZN(n10201) );
  INV_X1 U12862 ( .A(n10201), .ZN(n10202) );
  MUX2_X1 U12863 ( .A(n10203), .B(n10202), .S(P2_IR_REG_0__SCAN_IN), .Z(n10205) );
  NAND2_X1 U12864 ( .A1(n14762), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n10204) );
  OAI211_X1 U12865 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n8495), .A(n10205), .B(
        n10204), .ZN(P2_U3214) );
  NOR2_X1 U12866 ( .A1(n10411), .A2(n10206), .ZN(n10207) );
  AOI21_X1 U12867 ( .B1(n10206), .B2(n10411), .A(n10207), .ZN(n10210) );
  AOI21_X1 U12868 ( .B1(n10211), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10208), 
        .ZN(n10209) );
  NAND2_X1 U12869 ( .A1(n10209), .A2(n10210), .ZN(n10407) );
  OAI21_X1 U12870 ( .B1(n10210), .B2(n10209), .A(n10407), .ZN(n10222) );
  OR2_X1 U12871 ( .A1(n10211), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10215) );
  NAND2_X1 U12872 ( .A1(n10217), .A2(n10215), .ZN(n10213) );
  NAND2_X1 U12873 ( .A1(n10408), .A2(n11464), .ZN(n10212) );
  OAI21_X1 U12874 ( .B1(n10408), .B2(n11464), .A(n10212), .ZN(n10214) );
  NAND2_X1 U12875 ( .A1(n10213), .A2(n10214), .ZN(n10413) );
  INV_X1 U12876 ( .A(n10214), .ZN(n10216) );
  NAND3_X1 U12877 ( .A1(n10217), .A2(n10216), .A3(n10215), .ZN(n10218) );
  AOI21_X1 U12878 ( .B1(n10413), .B2(n10218), .A(n13176), .ZN(n10221) );
  NAND2_X1 U12879 ( .A1(n14762), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n10219) );
  NAND2_X1 U12880 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11420)
         );
  OAI211_X1 U12881 ( .C1(n14794), .C2(n10411), .A(n10219), .B(n11420), .ZN(
        n10220) );
  AOI211_X1 U12882 ( .C1(n10222), .C2(n14816), .A(n10221), .B(n10220), .ZN(
        n10223) );
  INV_X1 U12883 ( .A(n10223), .ZN(P2_U3226) );
  INV_X1 U12884 ( .A(SI_19_), .ZN(n15270) );
  OAI222_X1 U12885 ( .A1(n14376), .A2(n15270), .B1(P3_U3151), .B2(n12459), 
        .C1(n14378), .C2(n10224), .ZN(P3_U3276) );
  OAI21_X1 U12886 ( .B1(n10229), .B2(P1_REG1_REG_12__SCAN_IN), .A(n10225), 
        .ZN(n10227) );
  MUX2_X1 U12887 ( .A(n9366), .B(P1_REG1_REG_13__SCAN_IN), .S(n10244), .Z(
        n10226) );
  NOR2_X1 U12888 ( .A1(n10227), .A2(n10226), .ZN(n10240) );
  AOI211_X1 U12889 ( .C1(n10227), .C2(n10226), .A(n13926), .B(n10240), .ZN(
        n10228) );
  INV_X1 U12890 ( .A(n10228), .ZN(n10238) );
  NAND2_X1 U12891 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11579)
         );
  MUX2_X1 U12892 ( .A(n11500), .B(P1_REG2_REG_13__SCAN_IN), .S(n10244), .Z(
        n10232) );
  OR2_X1 U12893 ( .A1(n10229), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U12894 ( .A1(n10231), .A2(n10230), .ZN(n10233) );
  AOI21_X1 U12895 ( .B1(n10232), .B2(n10233), .A(n14604), .ZN(n10234) );
  NAND2_X1 U12896 ( .A1(n10234), .A2(n10250), .ZN(n10235) );
  NAND2_X1 U12897 ( .A1(n11579), .A2(n10235), .ZN(n10236) );
  AOI21_X1 U12898 ( .B1(n14594), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10236), 
        .ZN(n10237) );
  OAI211_X1 U12899 ( .C1(n14602), .C2(n10239), .A(n10238), .B(n10237), .ZN(
        P1_U3256) );
  AOI21_X1 U12900 ( .B1(n10244), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10240), 
        .ZN(n10712) );
  XNOR2_X1 U12901 ( .A(n10716), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10241) );
  XNOR2_X1 U12902 ( .A(n10712), .B(n10241), .ZN(n10254) );
  NAND2_X1 U12903 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13722)
         );
  INV_X1 U12904 ( .A(n13722), .ZN(n10243) );
  INV_X1 U12905 ( .A(n10716), .ZN(n10709) );
  NOR2_X1 U12906 ( .A1(n14602), .A2(n10709), .ZN(n10242) );
  AOI211_X1 U12907 ( .C1(n14594), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n10243), 
        .B(n10242), .ZN(n10253) );
  NAND2_X1 U12908 ( .A1(n10244), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10249) );
  NAND2_X1 U12909 ( .A1(n10250), .A2(n10249), .ZN(n10247) );
  MUX2_X1 U12910 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n10245), .S(n10716), .Z(
        n10246) );
  NAND2_X1 U12911 ( .A1(n10247), .A2(n10246), .ZN(n10718) );
  MUX2_X1 U12912 ( .A(n10245), .B(P1_REG2_REG_14__SCAN_IN), .S(n10716), .Z(
        n10248) );
  NAND3_X1 U12913 ( .A1(n10250), .A2(n10249), .A3(n10248), .ZN(n10251) );
  NAND3_X1 U12914 ( .A1(n10718), .A2(n13976), .A3(n10251), .ZN(n10252) );
  OAI211_X1 U12915 ( .C1(n10254), .C2(n13926), .A(n10253), .B(n10252), .ZN(
        P1_U3257) );
  MUX2_X1 U12916 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n11248), .Z(n10274) );
  XOR2_X1 U12917 ( .A(n10278), .B(n10274), .Z(n10275) );
  INV_X1 U12918 ( .A(n6433), .ZN(n10257) );
  AOI22_X1 U12919 ( .A1(n10258), .A2(n14979), .B1(n10257), .B2(n10256), .ZN(
        n10276) );
  XOR2_X1 U12920 ( .A(n10275), .B(n10276), .Z(n10273) );
  INV_X1 U12921 ( .A(n15015), .ZN(n14991) );
  AOI22_X1 U12922 ( .A1(n14995), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10270) );
  INV_X1 U12923 ( .A(n15001), .ZN(n15019) );
  OAI21_X1 U12924 ( .B1(n10261), .B2(n10260), .A(n10281), .ZN(n10262) );
  NAND2_X1 U12925 ( .A1(n15019), .A2(n10262), .ZN(n10269) );
  MUX2_X1 U12926 ( .A(n10263), .B(P3_REG1_REG_2__SCAN_IN), .S(n10278), .Z(
        n10266) );
  NAND2_X1 U12927 ( .A1(n10264), .A2(n7646), .ZN(n10265) );
  NAND2_X1 U12928 ( .A1(n10266), .A2(n10265), .ZN(n10277) );
  OAI21_X1 U12929 ( .B1(n10266), .B2(n10265), .A(n10277), .ZN(n10267) );
  NAND2_X1 U12930 ( .A1(n15007), .A2(n10267), .ZN(n10268) );
  NAND3_X1 U12931 ( .A1(n10270), .A2(n10269), .A3(n10268), .ZN(n10271) );
  AOI21_X1 U12932 ( .B1(n10278), .B2(n15017), .A(n10271), .ZN(n10272) );
  OAI21_X1 U12933 ( .B1(n10273), .B2(n14991), .A(n10272), .ZN(P3_U3184) );
  MUX2_X1 U12934 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n11248), .Z(n10313) );
  XNOR2_X1 U12935 ( .A(n10313), .B(n10317), .ZN(n10315) );
  INV_X1 U12936 ( .A(n10278), .ZN(n10279) );
  OAI22_X1 U12937 ( .A1(n10276), .A2(n10275), .B1(n10274), .B2(n10279), .ZN(
        n10316) );
  XOR2_X1 U12938 ( .A(n10315), .B(n10316), .Z(n10289) );
  XOR2_X1 U12939 ( .A(P3_REG1_REG_3__SCAN_IN), .B(n10325), .Z(n10286) );
  NAND2_X1 U12940 ( .A1(n10279), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10280) );
  OAI21_X1 U12941 ( .B1(n10282), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10320), .ZN(
        n10283) );
  NAND2_X1 U12942 ( .A1(n15019), .A2(n10283), .ZN(n10285) );
  INV_X1 U12943 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15052) );
  NOR2_X1 U12944 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15052), .ZN(n10602) );
  AOI21_X1 U12945 ( .B1(n14995), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10602), .ZN(
        n10284) );
  OAI211_X1 U12946 ( .C1(n10286), .C2(n14976), .A(n10285), .B(n10284), .ZN(
        n10287) );
  AOI21_X1 U12947 ( .B1(n10317), .B2(n15017), .A(n10287), .ZN(n10288) );
  OAI21_X1 U12948 ( .B1(n10289), .B2(n14991), .A(n10288), .ZN(P3_U3185) );
  AND2_X1 U12949 ( .A1(n13118), .A2(n14879), .ZN(n14869) );
  XNOR2_X1 U12950 ( .A(n10657), .B(n10661), .ZN(n10994) );
  INV_X1 U12951 ( .A(n14934), .ZN(n14918) );
  AOI21_X1 U12952 ( .B1(n14866), .B2(n13048), .A(n9733), .ZN(n10290) );
  NAND2_X1 U12953 ( .A1(n10290), .A2(n10673), .ZN(n10999) );
  OAI21_X1 U12954 ( .B1(n10658), .B2(n14953), .A(n10999), .ZN(n10304) );
  AND4_X1 U12955 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n10820) );
  INV_X1 U12956 ( .A(n13116), .ZN(n14886) );
  INV_X1 U12957 ( .A(n10295), .ZN(n14862) );
  NAND2_X1 U12958 ( .A1(n14862), .A2(n10296), .ZN(n10299) );
  NAND2_X1 U12959 ( .A1(n14886), .A2(n10297), .ZN(n10298) );
  NAND2_X1 U12960 ( .A1(n10299), .A2(n10298), .ZN(n10663) );
  XNOR2_X1 U12961 ( .A(n10663), .B(n10661), .ZN(n10303) );
  NAND2_X1 U12962 ( .A1(n8449), .A2(n10300), .ZN(n10301) );
  NAND2_X2 U12963 ( .A1(n10302), .A2(n10301), .ZN(n14882) );
  OAI222_X1 U12964 ( .A1(n14885), .A2(n10820), .B1(n13422), .B2(n14886), .C1(
        n10303), .C2(n13424), .ZN(n11001) );
  AOI211_X1 U12965 ( .C1(n10994), .C2(n14918), .A(n10304), .B(n11001), .ZN(
        n14911) );
  NOR2_X1 U12966 ( .A1(n10306), .A2(n10305), .ZN(n10653) );
  AND2_X1 U12967 ( .A1(n14896), .A2(n10307), .ZN(n10308) );
  INV_X1 U12968 ( .A(n14894), .ZN(n10309) );
  NAND2_X1 U12969 ( .A1(n14971), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10310) );
  OAI21_X1 U12970 ( .B1(n14911), .B2(n14971), .A(n10310), .ZN(P2_U3501) );
  INV_X1 U12971 ( .A(n10311), .ZN(n10336) );
  INV_X1 U12972 ( .A(n10982), .ZN(n10729) );
  OAI222_X1 U12973 ( .A1(n11585), .A2(n10336), .B1(n10729), .B2(P1_U3086), 
        .C1(n10312), .C2(n14353), .ZN(P1_U3339) );
  MUX2_X1 U12974 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n11248), .Z(n10371) );
  XOR2_X1 U12975 ( .A(n10379), .B(n10371), .Z(n10372) );
  INV_X1 U12976 ( .A(n10313), .ZN(n10314) );
  AOI22_X1 U12977 ( .A1(n10316), .A2(n10315), .B1(n10317), .B2(n10314), .ZN(
        n10373) );
  XOR2_X1 U12978 ( .A(n10372), .B(n10373), .Z(n10334) );
  INV_X1 U12979 ( .A(n10317), .ZN(n10324) );
  NAND2_X1 U12980 ( .A1(n10318), .A2(n10324), .ZN(n10319) );
  MUX2_X1 U12981 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10374), .S(n10379), .Z(
        n10321) );
  AOI21_X1 U12982 ( .B1(n10322), .B2(n10321), .A(n10376), .ZN(n10331) );
  AND2_X1 U12983 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U12984 ( .A1(n10325), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n10324), 
        .B2(n10323), .ZN(n10327) );
  MUX2_X1 U12985 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n7728), .S(n10379), .Z(
        n10326) );
  NAND2_X1 U12986 ( .A1(n10327), .A2(n10326), .ZN(n10328) );
  AOI21_X1 U12987 ( .B1(n10378), .B2(n10328), .A(n14976), .ZN(n10329) );
  AOI211_X1 U12988 ( .C1(n14995), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n10908), .B(
        n10329), .ZN(n10330) );
  OAI21_X1 U12989 ( .B1(n10331), .B2(n15001), .A(n10330), .ZN(n10332) );
  AOI21_X1 U12990 ( .B1(n10379), .B2(n15017), .A(n10332), .ZN(n10333) );
  OAI21_X1 U12991 ( .B1(n10334), .B2(n14991), .A(n10333), .ZN(P3_U3186) );
  INV_X1 U12992 ( .A(n11434), .ZN(n11211) );
  OAI222_X1 U12993 ( .A1(P2_U3088), .A2(n11211), .B1(n13590), .B2(n10336), 
        .C1(n10335), .C2(n13588), .ZN(P2_U3311) );
  INV_X1 U12994 ( .A(n10337), .ZN(n10340) );
  OAI222_X1 U12995 ( .A1(n11585), .A2(n10340), .B1(n10709), .B2(P1_U3086), 
        .C1(n10338), .C2(n14353), .ZN(P1_U3341) );
  INV_X1 U12996 ( .A(n11204), .ZN(n10341) );
  OAI222_X1 U12997 ( .A1(P2_U3088), .A2(n10341), .B1(n13590), .B2(n10340), 
        .C1(n10339), .C2(n13588), .ZN(P2_U3313) );
  NAND2_X1 U12998 ( .A1(n10357), .A2(n10354), .ZN(n10345) );
  INV_X1 U12999 ( .A(n10355), .ZN(n10342) );
  NAND2_X1 U13000 ( .A1(n10356), .A2(n10342), .ZN(n10343) );
  NAND2_X1 U13001 ( .A1(n10538), .A2(n11748), .ZN(n10497) );
  NAND4_X1 U13002 ( .A1(n10345), .A2(n10344), .A3(n10343), .A4(n10497), .ZN(
        n10346) );
  NAND2_X1 U13003 ( .A1(n10346), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10350) );
  INV_X1 U13004 ( .A(n11796), .ZN(n10347) );
  AOI21_X1 U13005 ( .B1(n10348), .B2(n10356), .A(n10347), .ZN(n10349) );
  NOR2_X1 U13006 ( .A1(n12324), .A2(P3_U3151), .ZN(n10587) );
  NOR2_X1 U13007 ( .A1(n10356), .A2(n11792), .ZN(n10550) );
  AND2_X1 U13008 ( .A1(n10358), .A2(n14477), .ZN(n10351) );
  INV_X1 U13009 ( .A(n10351), .ZN(n10352) );
  OR2_X1 U13010 ( .A1(n10357), .A2(n10352), .ZN(n10353) );
  AOI22_X1 U13011 ( .A1(n12344), .A2(n15068), .B1(n10503), .B2(n12330), .ZN(
        n10362) );
  NAND2_X1 U13012 ( .A1(n6905), .A2(n12055), .ZN(n11637) );
  AND2_X1 U13013 ( .A1(n12777), .A2(n11637), .ZN(n11769) );
  INV_X1 U13014 ( .A(n11769), .ZN(n10360) );
  NAND2_X1 U13015 ( .A1(n10354), .A2(n15111), .ZN(n10391) );
  OAI22_X1 U13016 ( .A1(n10357), .A2(n10391), .B1(n10356), .B2(n10355), .ZN(
        n10359) );
  NAND2_X1 U13017 ( .A1(n10360), .A2(n12337), .ZN(n10361) );
  OAI211_X1 U13018 ( .C1(n10587), .C2(n7694), .A(n10362), .B(n10361), .ZN(
        P3_U3172) );
  INV_X1 U13019 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n10364) );
  NAND2_X1 U13020 ( .A1(n12265), .A2(P3_U3897), .ZN(n10363) );
  OAI21_X1 U13021 ( .B1(P3_U3897), .B2(n10364), .A(n10363), .ZN(P3_U3514) );
  NAND2_X1 U13022 ( .A1(n13085), .A2(n9733), .ZN(n13075) );
  AOI22_X1 U13023 ( .A1(n13046), .A2(n13116), .B1(n14879), .B2(n13093), .ZN(
        n10368) );
  OR2_X1 U13024 ( .A1(n10365), .A2(P2_U3088), .ZN(n13047) );
  AOI22_X1 U13025 ( .A1(n13085), .A2(n10366), .B1(n13047), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10367) );
  OAI211_X1 U13026 ( .C1(n10369), .C2(n13075), .A(n10368), .B(n10367), .ZN(
        P2_U3204) );
  MUX2_X1 U13027 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n11248), .Z(n10469) );
  XNOR2_X1 U13028 ( .A(n10469), .B(n10471), .ZN(n10472) );
  INV_X1 U13029 ( .A(n10379), .ZN(n10370) );
  XOR2_X1 U13030 ( .A(n10472), .B(n10473), .Z(n10386) );
  NOR2_X1 U13031 ( .A1(n10379), .A2(n10374), .ZN(n10375) );
  XNOR2_X1 U13032 ( .A(n10480), .B(n10471), .ZN(n10377) );
  NAND2_X1 U13033 ( .A1(n10377), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n10479) );
  OAI21_X1 U13034 ( .B1(n10377), .B2(P3_REG2_REG_5__SCAN_IN), .A(n10479), .ZN(
        n10384) );
  INV_X1 U13035 ( .A(n10471), .ZN(n10481) );
  XNOR2_X1 U13036 ( .A(n10474), .B(n10471), .ZN(n10475) );
  XOR2_X1 U13037 ( .A(n10475), .B(P3_REG1_REG_5__SCAN_IN), .Z(n10380) );
  OAI22_X1 U13038 ( .A1(n14989), .A2(n10481), .B1(n10380), .B2(n14976), .ZN(
        n10383) );
  NAND2_X1 U13039 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n11009) );
  OAI21_X1 U13040 ( .B1(n15024), .B2(n10381), .A(n11009), .ZN(n10382) );
  AOI211_X1 U13041 ( .C1(n15019), .C2(n10384), .A(n10383), .B(n10382), .ZN(
        n10385) );
  OAI21_X1 U13042 ( .B1(n10386), .B2(n14991), .A(n10385), .ZN(P3_U3187) );
  INV_X1 U13043 ( .A(n10387), .ZN(n10397) );
  OAI222_X1 U13044 ( .A1(n11585), .A2(n10397), .B1(n11320), .B2(P1_U3086), 
        .C1(n10388), .C2(n14353), .ZN(P1_U3338) );
  INV_X1 U13045 ( .A(n10389), .ZN(n10404) );
  INV_X1 U13046 ( .A(n10719), .ZN(n14603) );
  OAI222_X1 U13047 ( .A1(n11585), .A2(n10404), .B1(n14603), .B2(P1_U3086), 
        .C1(n10390), .C2(n14353), .ZN(P1_U3340) );
  AOI21_X1 U13048 ( .B1(n15043), .B2(n10391), .A(n11769), .ZN(n10392) );
  AOI21_X1 U13049 ( .B1(n15066), .B2(n15068), .A(n10392), .ZN(n12052) );
  INV_X1 U13050 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10393) );
  OAI22_X1 U13051 ( .A1(n12055), .A2(n12846), .B1(n15136), .B2(n10393), .ZN(
        n10394) );
  INV_X1 U13052 ( .A(n10394), .ZN(n10395) );
  OAI21_X1 U13053 ( .B1(n12052), .B2(n15137), .A(n10395), .ZN(P3_U3390) );
  OAI222_X1 U13054 ( .A1(P2_U3088), .A2(n13159), .B1(n13590), .B2(n10397), 
        .C1(n10396), .C2(n13588), .ZN(P2_U3310) );
  INV_X1 U13055 ( .A(n13115), .ZN(n10664) );
  OAI22_X1 U13056 ( .A1(n10398), .A2(n13422), .B1(n10664), .B2(n14885), .ZN(
        n14863) );
  AOI22_X1 U13057 ( .A1(n13089), .A2(n14863), .B1(n13047), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U13058 ( .A1(n13085), .A2(n10401), .ZN(n10402) );
  OAI211_X1 U13059 ( .C1(n14906), .C2(n13023), .A(n10403), .B(n10402), .ZN(
        P2_U3194) );
  INV_X1 U13060 ( .A(n11198), .ZN(n13150) );
  OAI222_X1 U13061 ( .A1(n13588), .A2(n10405), .B1(n13590), .B2(n10404), .C1(
        n13150), .C2(P2_U3088), .ZN(P2_U3312) );
  MUX2_X1 U13062 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n10406), .S(n10414), .Z(
        n10410) );
  OAI21_X1 U13063 ( .B1(n10408), .B2(P2_REG1_REG_12__SCAN_IN), .A(n10407), 
        .ZN(n10409) );
  NOR2_X1 U13064 ( .A1(n10409), .A2(n10410), .ZN(n10630) );
  AOI211_X1 U13065 ( .C1(n10410), .C2(n10409), .A(n14844), .B(n10630), .ZN(
        n10422) );
  NAND2_X1 U13066 ( .A1(n10411), .A2(n11464), .ZN(n10412) );
  MUX2_X1 U13067 ( .A(n10415), .B(P2_REG2_REG_13__SCAN_IN), .S(n10414), .Z(
        n10416) );
  NAND2_X1 U13068 ( .A1(n10417), .A2(n10416), .ZN(n10625) );
  OAI211_X1 U13069 ( .C1(n10417), .C2(n10416), .A(n10625), .B(n14838), .ZN(
        n10420) );
  NOR2_X1 U13070 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8750), .ZN(n10418) );
  AOI21_X1 U13071 ( .B1(n14840), .B2(n10631), .A(n10418), .ZN(n10419) );
  OAI211_X1 U13072 ( .C1(n14848), .C2(n6965), .A(n10420), .B(n10419), .ZN(
        n10421) );
  OR2_X1 U13073 ( .A1(n10422), .A2(n10421), .ZN(P2_U3227) );
  INV_X1 U13074 ( .A(n10423), .ZN(n10425) );
  OAI222_X1 U13075 ( .A1(n14378), .A2(n10425), .B1(n14376), .B2(n10424), .C1(
        P3_U3151), .C2(n10536), .ZN(P3_U3275) );
  INV_X1 U13076 ( .A(n13872), .ZN(n11833) );
  OAI22_X1 U13077 ( .A1(n11833), .A2(n13749), .B1(n14692), .B2(n13752), .ZN(
        n10449) );
  INV_X2 U13078 ( .A(n10430), .ZN(n13700) );
  NAND2_X1 U13079 ( .A1(n13872), .A2(n13700), .ZN(n10428) );
  NAND2_X1 U13080 ( .A1(n11832), .A2(n13699), .ZN(n10427) );
  NAND2_X1 U13081 ( .A1(n10428), .A2(n10427), .ZN(n10429) );
  XNOR2_X1 U13082 ( .A(n10429), .B(n10692), .ZN(n10448) );
  XOR2_X1 U13083 ( .A(n10449), .B(n10448), .Z(n10439) );
  OAI22_X1 U13084 ( .A1(n9213), .A2(n13749), .B1(n10751), .B2(n13752), .ZN(
        n10432) );
  NOR2_X1 U13085 ( .A1(n10433), .A2(n10432), .ZN(n10436) );
  AOI21_X1 U13086 ( .B1(n10433), .B2(n10432), .A(n10436), .ZN(n13766) );
  OAI21_X1 U13087 ( .B1(n10435), .B2(n6937), .A(n10434), .ZN(n13765) );
  INV_X1 U13088 ( .A(n10436), .ZN(n10437) );
  OAI21_X1 U13089 ( .B1(n10439), .B2(n10438), .A(n10454), .ZN(n10440) );
  NAND2_X1 U13090 ( .A1(n10440), .A2(n14532), .ZN(n10443) );
  INV_X1 U13091 ( .A(n13871), .ZN(n10441) );
  OAI22_X1 U13092 ( .A1(n9213), .A2(n14127), .B1(n10441), .B2(n14617), .ZN(
        n10880) );
  AOI22_X1 U13093 ( .A1(n10880), .A2(n15299), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n13768), .ZN(n10442) );
  OAI211_X1 U13094 ( .C1(n14692), .C2(n14530), .A(n10443), .B(n10442), .ZN(
        P1_U3237) );
  NAND2_X1 U13095 ( .A1(n13871), .A2(n13700), .ZN(n10445) );
  NAND2_X1 U13096 ( .A1(n11839), .A2(n13699), .ZN(n10444) );
  NAND2_X1 U13097 ( .A1(n10445), .A2(n10444), .ZN(n10446) );
  XNOR2_X1 U13098 ( .A(n10446), .B(n10692), .ZN(n10608) );
  AND2_X1 U13099 ( .A1(n11839), .A2(n13608), .ZN(n10447) );
  XNOR2_X1 U13100 ( .A(n10608), .B(n10606), .ZN(n10452) );
  INV_X1 U13101 ( .A(n10448), .ZN(n10451) );
  INV_X1 U13102 ( .A(n10449), .ZN(n10450) );
  NAND2_X1 U13103 ( .A1(n10451), .A2(n10450), .ZN(n10453) );
  NAND2_X1 U13104 ( .A1(n10611), .A2(n14532), .ZN(n10468) );
  AOI21_X1 U13105 ( .B1(n10454), .B2(n10453), .A(n10452), .ZN(n10467) );
  NAND2_X1 U13106 ( .A1(n10456), .A2(n10455), .ZN(n10460) );
  NOR2_X1 U13107 ( .A1(n10458), .A2(n10457), .ZN(n10459) );
  NAND2_X1 U13108 ( .A1(n10460), .A2(n10459), .ZN(n10461) );
  NAND2_X1 U13109 ( .A1(n10461), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10462) );
  INV_X1 U13110 ( .A(n15303), .ZN(n13843) );
  NAND2_X1 U13111 ( .A1(n14528), .A2(n13870), .ZN(n10463) );
  NAND2_X1 U13112 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13898) );
  NAND2_X1 U13113 ( .A1(n10463), .A2(n13898), .ZN(n10465) );
  INV_X1 U13114 ( .A(n14526), .ZN(n14509) );
  OAI22_X1 U13115 ( .A1(n14530), .A2(n11840), .B1(n14509), .B2(n11833), .ZN(
        n10464) );
  AOI211_X1 U13116 ( .C1(n9241), .C2(n13843), .A(n10465), .B(n10464), .ZN(
        n10466) );
  OAI21_X1 U13117 ( .B1(n10468), .B2(n10467), .A(n10466), .ZN(P1_U3218) );
  MUX2_X1 U13118 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n11248), .Z(n10567) );
  XNOR2_X1 U13119 ( .A(n10567), .B(n10577), .ZN(n10568) );
  INV_X1 U13120 ( .A(n10469), .ZN(n10470) );
  XOR2_X1 U13121 ( .A(n10568), .B(n10569), .Z(n10492) );
  INV_X1 U13122 ( .A(n10577), .ZN(n10572) );
  MUX2_X1 U13123 ( .A(n7762), .B(P3_REG1_REG_6__SCAN_IN), .S(n10577), .Z(
        n10477) );
  AOI22_X1 U13124 ( .A1(n10475), .A2(P3_REG1_REG_5__SCAN_IN), .B1(n10481), 
        .B2(n10474), .ZN(n10476) );
  AOI21_X1 U13125 ( .B1(n10477), .B2(n10476), .A(n10570), .ZN(n10478) );
  NOR2_X1 U13126 ( .A1(n14976), .A2(n10478), .ZN(n10490) );
  INV_X1 U13127 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10482) );
  MUX2_X1 U13128 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n10482), .S(n10577), .Z(
        n10483) );
  INV_X1 U13129 ( .A(n10483), .ZN(n10484) );
  AOI21_X1 U13130 ( .B1(n10485), .B2(n10484), .A(n10576), .ZN(n10488) );
  NAND2_X1 U13131 ( .A1(n14995), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10487) );
  AND2_X1 U13132 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11049) );
  INV_X1 U13133 ( .A(n11049), .ZN(n10486) );
  OAI211_X1 U13134 ( .C1(n15001), .C2(n10488), .A(n10487), .B(n10486), .ZN(
        n10489) );
  AOI211_X1 U13135 ( .C1(n15017), .C2(n10572), .A(n10490), .B(n10489), .ZN(
        n10491) );
  OAI21_X1 U13136 ( .B1(n10492), .B2(n14991), .A(n10491), .ZN(P3_U3188) );
  INV_X1 U13137 ( .A(n10493), .ZN(n10500) );
  OR2_X1 U13138 ( .A1(n10494), .A2(n11748), .ZN(n10495) );
  XNOR2_X1 U13139 ( .A(n10496), .B(n10495), .ZN(n10498) );
  NAND2_X1 U13140 ( .A1(n10500), .A2(n10499), .ZN(n10502) );
  MUX2_X1 U13141 ( .A(n10501), .B(n12052), .S(n15091), .Z(n10505) );
  INV_X1 U13142 ( .A(n12691), .ZN(n14462) );
  AOI22_X1 U13143 ( .A1(n14462), .A2(n10503), .B1(n15053), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10504) );
  NAND2_X1 U13144 ( .A1(n10505), .A2(n10504), .ZN(P3_U3233) );
  OAI21_X1 U13145 ( .B1(n10508), .B2(n10507), .A(n10506), .ZN(n10509) );
  NAND2_X1 U13146 ( .A1(n10509), .A2(n13085), .ZN(n10514) );
  NAND2_X1 U13147 ( .A1(n13111), .A2(n13441), .ZN(n10511) );
  NAND2_X1 U13148 ( .A1(n13113), .A2(n13444), .ZN(n10510) );
  NAND2_X1 U13149 ( .A1(n10511), .A2(n10510), .ZN(n10827) );
  AND2_X1 U13150 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n14807) );
  OAI22_X1 U13151 ( .A1(n13023), .A2(n6592), .B1(n10831), .B2(n13091), .ZN(
        n10512) );
  AOI211_X1 U13152 ( .C1(n13089), .C2(n10827), .A(n14807), .B(n10512), .ZN(
        n10513) );
  NAND2_X1 U13153 ( .A1(n10514), .A2(n10513), .ZN(P2_U3199) );
  OAI222_X1 U13154 ( .A1(n14378), .A2(n10517), .B1(n14376), .B2(n10516), .C1(
        P3_U3151), .C2(n10515), .ZN(P3_U3274) );
  XNOR2_X1 U13155 ( .A(n10519), .B(n10518), .ZN(n10522) );
  INV_X1 U13156 ( .A(n13113), .ZN(n10823) );
  OAI22_X1 U13157 ( .A1(n10664), .A2(n13422), .B1(n10823), .B2(n14885), .ZN(
        n10667) );
  AND2_X1 U13158 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n14781) );
  OAI22_X1 U13159 ( .A1(n13023), .A2(n14914), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13091), .ZN(n10520) );
  AOI211_X1 U13160 ( .C1(n13089), .C2(n10667), .A(n14781), .B(n10520), .ZN(
        n10521) );
  OAI21_X1 U13161 ( .B1(n10522), .B2(n13082), .A(n10521), .ZN(P2_U3190) );
  OAI21_X1 U13162 ( .B1(n10525), .B2(n10524), .A(n10523), .ZN(n10528) );
  AOI22_X1 U13163 ( .A1(n13444), .A2(n13114), .B1(n13112), .B2(n13441), .ZN(
        n10838) );
  NAND2_X1 U13164 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n14791) );
  OAI21_X1 U13165 ( .B1(n12996), .B2(n10838), .A(n14791), .ZN(n10527) );
  OAI22_X1 U13166 ( .A1(n13023), .A2(n14927), .B1(n13091), .B2(n10846), .ZN(
        n10526) );
  AOI211_X1 U13167 ( .C1(n10528), .C2(n13085), .A(n10527), .B(n10526), .ZN(
        n10529) );
  INV_X1 U13168 ( .A(n10529), .ZN(P2_U3202) );
  XNOR2_X1 U13169 ( .A(n10530), .B(n10531), .ZN(n10535) );
  AOI22_X1 U13170 ( .A1(n13046), .A2(n13110), .B1(n10965), .B2(n13093), .ZN(
        n10534) );
  NAND2_X1 U13171 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13122) );
  OAI21_X1 U13172 ( .B1(n13091), .B2(n10963), .A(n13122), .ZN(n10532) );
  AOI21_X1 U13173 ( .B1(n13078), .B2(n13112), .A(n10532), .ZN(n10533) );
  OAI211_X1 U13174 ( .C1(n10535), .C2(n13082), .A(n10534), .B(n10533), .ZN(
        P2_U3211) );
  NAND2_X1 U13175 ( .A1(n11639), .A2(n10536), .ZN(n10537) );
  NAND2_X1 U13176 ( .A1(n10540), .A2(n10541), .ZN(n10585) );
  INV_X1 U13177 ( .A(n10541), .ZN(n10542) );
  INV_X1 U13178 ( .A(n12770), .ZN(n10543) );
  NAND3_X1 U13179 ( .A1(n10546), .A2(n12777), .A3(n10597), .ZN(n10547) );
  OAI211_X1 U13180 ( .C1(n10548), .C2(n12770), .A(n10586), .B(n10547), .ZN(
        n10549) );
  NAND2_X1 U13181 ( .A1(n10549), .A2(n12337), .ZN(n10553) );
  INV_X1 U13182 ( .A(n12772), .ZN(n15049) );
  INV_X1 U13183 ( .A(n12330), .ZN(n12347) );
  OAI22_X1 U13184 ( .A1(n15049), .A2(n12327), .B1(n12347), .B2(n12780), .ZN(
        n10551) );
  AOI21_X1 U13185 ( .B1(n12323), .B2(n6905), .A(n10551), .ZN(n10552) );
  OAI211_X1 U13186 ( .C1(n10587), .C2(n15082), .A(n10553), .B(n10552), .ZN(
        P3_U3162) );
  INV_X1 U13187 ( .A(n11515), .ZN(n11327) );
  OAI222_X1 U13188 ( .A1(n11585), .A2(n10566), .B1(n11327), .B2(P1_U3086), 
        .C1(n10554), .C2(n14353), .ZN(P1_U3337) );
  OAI21_X1 U13189 ( .B1(n6588), .B2(n11990), .A(n10555), .ZN(n14702) );
  NAND2_X1 U13190 ( .A1(n10556), .A2(n11990), .ZN(n10557) );
  NAND3_X1 U13191 ( .A1(n10558), .A2(n14403), .A3(n10557), .ZN(n10560) );
  AOI22_X1 U13192 ( .A1(n14619), .A2(n13871), .B1(n13869), .B2(n14404), .ZN(
        n10559) );
  NAND2_X1 U13193 ( .A1(n10560), .A2(n10559), .ZN(n14698) );
  MUX2_X1 U13194 ( .A(n14698), .B(P1_REG2_REG_4__SCAN_IN), .S(n14656), .Z(
        n10561) );
  INV_X1 U13195 ( .A(n10561), .ZN(n10564) );
  AOI211_X1 U13196 ( .C1(n14700), .C2(n10744), .A(n14715), .B(n10645), .ZN(
        n14699) );
  OAI22_X1 U13197 ( .A1(n14190), .A2(n10616), .B1(n14229), .B2(n10615), .ZN(
        n10562) );
  AOI21_X1 U13198 ( .B1(n14699), .B2(n14633), .A(n10562), .ZN(n10563) );
  OAI211_X1 U13199 ( .C1(n14202), .C2(n14702), .A(n10564), .B(n10563), .ZN(
        P1_U3289) );
  INV_X1 U13200 ( .A(n13162), .ZN(n13171) );
  OAI222_X1 U13201 ( .A1(P2_U3088), .A2(n13171), .B1(n13590), .B2(n10566), 
        .C1(n10565), .C2(n13588), .ZN(P2_U3309) );
  MUX2_X1 U13202 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n11248), .Z(n10767) );
  XNOR2_X1 U13203 ( .A(n10767), .B(n10779), .ZN(n10769) );
  XOR2_X1 U13204 ( .A(n10769), .B(n10770), .Z(n10584) );
  INV_X1 U13205 ( .A(n10570), .ZN(n10571) );
  XNOR2_X1 U13206 ( .A(n10771), .B(n10779), .ZN(n10573) );
  NAND2_X1 U13207 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10573), .ZN(n10773) );
  OAI21_X1 U13208 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10573), .A(n10773), .ZN(
        n10582) );
  INV_X1 U13209 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10574) );
  NOR2_X1 U13210 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10574), .ZN(n11292) );
  AOI21_X1 U13211 ( .B1(n14995), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11292), .ZN(
        n10575) );
  OAI21_X1 U13212 ( .B1(n14989), .B2(n10772), .A(n10575), .ZN(n10581) );
  AOI21_X1 U13213 ( .B1(n10578), .B2(n11311), .A(n10780), .ZN(n10579) );
  NOR2_X1 U13214 ( .A1(n10579), .A2(n15001), .ZN(n10580) );
  AOI211_X1 U13215 ( .C1(n15007), .C2(n10582), .A(n10581), .B(n10580), .ZN(
        n10583) );
  OAI21_X1 U13216 ( .B1(n10584), .B2(n14991), .A(n10583), .ZN(P3_U3189) );
  XNOR2_X1 U13217 ( .A(n15063), .B(n12159), .ZN(n10594) );
  XNOR2_X1 U13218 ( .A(n10594), .B(n12772), .ZN(n10592) );
  NAND2_X1 U13219 ( .A1(n10586), .A2(n10585), .ZN(n10593) );
  XOR2_X1 U13220 ( .A(n10593), .B(n10592), .Z(n10591) );
  INV_X1 U13221 ( .A(n15067), .ZN(n10906) );
  OAI22_X1 U13222 ( .A1(n10906), .A2(n12327), .B1(n12347), .B2(n15063), .ZN(
        n10589) );
  INV_X1 U13223 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15064) );
  NOR2_X1 U13224 ( .A1(n10587), .A2(n15064), .ZN(n10588) );
  AOI211_X1 U13225 ( .C1(n12323), .C2(n15068), .A(n10589), .B(n10588), .ZN(
        n10590) );
  OAI21_X1 U13226 ( .B1(n10591), .B2(n12332), .A(n10590), .ZN(P3_U3177) );
  INV_X1 U13227 ( .A(n10594), .ZN(n10595) );
  OR2_X1 U13228 ( .A1(n12772), .A2(n10595), .ZN(n10596) );
  XNOR2_X1 U13229 ( .A(n15057), .B(n10597), .ZN(n10900) );
  XNOR2_X1 U13230 ( .A(n10900), .B(n15067), .ZN(n10598) );
  AOI21_X1 U13231 ( .B1(n10599), .B2(n10598), .A(n12332), .ZN(n10600) );
  NAND2_X1 U13232 ( .A1(n10600), .A2(n10902), .ZN(n10605) );
  INV_X1 U13233 ( .A(n15030), .ZN(n15047) );
  OAI22_X1 U13234 ( .A1(n15049), .A2(n12340), .B1(n15047), .B2(n12327), .ZN(
        n10601) );
  AOI211_X1 U13235 ( .C1(n10603), .C2(n12330), .A(n10602), .B(n10601), .ZN(
        n10604) );
  OAI211_X1 U13236 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12339), .A(n10605), .B(
        n10604), .ZN(P3_U3158) );
  INV_X1 U13237 ( .A(n10606), .ZN(n10607) );
  NAND2_X1 U13238 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  AOI22_X1 U13239 ( .A1(n13870), .A2(n13704), .B1(n13608), .B2(n14700), .ZN(
        n10610) );
  NOR2_X1 U13240 ( .A1(n10688), .A2(n6581), .ZN(n10613) );
  AOI22_X1 U13241 ( .A1(n13870), .A2(n13608), .B1(n13699), .B2(n14700), .ZN(
        n10612) );
  XOR2_X1 U13242 ( .A(n10692), .B(n10612), .Z(n10689) );
  XNOR2_X1 U13243 ( .A(n10613), .B(n10689), .ZN(n10620) );
  NAND2_X1 U13244 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13927) );
  NAND2_X1 U13245 ( .A1(n14528), .A2(n13869), .ZN(n10614) );
  OAI211_X1 U13246 ( .C1(n15303), .C2(n10615), .A(n13927), .B(n10614), .ZN(
        n10618) );
  NOR2_X1 U13247 ( .A1(n14530), .A2(n10616), .ZN(n10617) );
  AOI211_X1 U13248 ( .C1(n14526), .C2(n13871), .A(n10618), .B(n10617), .ZN(
        n10619) );
  OAI21_X1 U13249 ( .B1(n10620), .B2(n15306), .A(n10619), .ZN(P1_U3230) );
  INV_X1 U13250 ( .A(n10621), .ZN(n10623) );
  OAI22_X1 U13251 ( .A1(n11793), .A2(P3_U3151), .B1(SI_22_), .B2(n14376), .ZN(
        n10622) );
  AOI21_X1 U13252 ( .B1(n10623), .B2(n14388), .A(n10622), .ZN(P3_U3273) );
  NAND2_X1 U13253 ( .A1(n10631), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10624) );
  NAND2_X1 U13254 ( .A1(n10625), .A2(n10624), .ZN(n11194) );
  XNOR2_X1 U13255 ( .A(n11194), .B(n11204), .ZN(n11195) );
  XNOR2_X1 U13256 ( .A(n11195), .B(n13431), .ZN(n10637) );
  NAND2_X1 U13257 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n12932)
         );
  INV_X1 U13258 ( .A(n12932), .ZN(n10626) );
  AOI21_X1 U13259 ( .B1(n14840), .B2(n11204), .A(n10626), .ZN(n10627) );
  INV_X1 U13260 ( .A(n10627), .ZN(n10635) );
  NOR2_X1 U13261 ( .A1(n11204), .A2(n10628), .ZN(n10629) );
  AOI21_X1 U13262 ( .B1(n11204), .B2(n10628), .A(n10629), .ZN(n10633) );
  NOR2_X1 U13263 ( .A1(n10632), .A2(n10633), .ZN(n11203) );
  AOI211_X1 U13264 ( .C1(n10633), .C2(n10632), .A(n14844), .B(n11203), .ZN(
        n10634) );
  AOI211_X1 U13265 ( .C1(n14762), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n10635), 
        .B(n10634), .ZN(n10636) );
  OAI21_X1 U13266 ( .B1(n10637), .B2(n13176), .A(n10636), .ZN(P2_U3228) );
  XNOR2_X1 U13267 ( .A(n10704), .B(n13869), .ZN(n11991) );
  XNOR2_X1 U13268 ( .A(n10638), .B(n11991), .ZN(n14710) );
  XNOR2_X1 U13269 ( .A(n10639), .B(n11991), .ZN(n10640) );
  NAND2_X1 U13270 ( .A1(n10640), .A2(n14403), .ZN(n10642) );
  AOI22_X1 U13271 ( .A1(n14619), .A2(n13870), .B1(n13868), .B2(n14404), .ZN(
        n10641) );
  NAND2_X1 U13272 ( .A1(n10642), .A2(n10641), .ZN(n14706) );
  INV_X1 U13273 ( .A(n14706), .ZN(n10644) );
  MUX2_X1 U13274 ( .A(n10644), .B(n10643), .S(n14656), .Z(n10650) );
  INV_X1 U13275 ( .A(n10645), .ZN(n10647) );
  INV_X1 U13276 ( .A(n10646), .ZN(n14650) );
  AOI211_X1 U13277 ( .C1(n14708), .C2(n10647), .A(n14715), .B(n14650), .ZN(
        n14707) );
  OAI22_X1 U13278 ( .A1(n14190), .A2(n10704), .B1(n10703), .B2(n14229), .ZN(
        n10648) );
  AOI21_X1 U13279 ( .B1(n14707), .B2(n14633), .A(n10648), .ZN(n10649) );
  OAI211_X1 U13280 ( .C1(n14710), .C2(n14202), .A(n10650), .B(n10649), .ZN(
        P1_U3288) );
  INV_X1 U13281 ( .A(n10651), .ZN(n10652) );
  NAND4_X1 U13282 ( .A1(n10653), .A2(n14895), .A3(n10652), .A4(n14894), .ZN(
        n10654) );
  NAND2_X1 U13283 ( .A1(n8474), .A2(n10655), .ZN(n10940) );
  NAND2_X1 U13284 ( .A1(n14922), .A2(n10940), .ZN(n10656) );
  NAND2_X1 U13285 ( .A1(n10657), .A2(n10661), .ZN(n10660) );
  NAND2_X1 U13286 ( .A1(n10664), .A2(n10658), .ZN(n10659) );
  XNOR2_X1 U13287 ( .A(n10811), .B(n10817), .ZN(n14912) );
  INV_X1 U13288 ( .A(n10661), .ZN(n10662) );
  NAND2_X1 U13289 ( .A1(n10663), .A2(n10662), .ZN(n10666) );
  NAND2_X1 U13290 ( .A1(n10664), .A2(n13048), .ZN(n10665) );
  NAND2_X1 U13291 ( .A1(n10666), .A2(n10665), .ZN(n10818) );
  XNOR2_X1 U13292 ( .A(n10818), .B(n10817), .ZN(n10668) );
  AOI21_X1 U13293 ( .B1(n10668), .B2(n14882), .A(n10667), .ZN(n14915) );
  MUX2_X1 U13294 ( .A(n10669), .B(n14915), .S(n13402), .Z(n10678) );
  INV_X1 U13295 ( .A(n10670), .ZN(n10671) );
  OAI22_X1 U13296 ( .A1(n14874), .A2(n14914), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14881), .ZN(n10676) );
  NAND2_X1 U13297 ( .A1(n10673), .A2(n10819), .ZN(n10672) );
  NAND2_X1 U13298 ( .A1(n10672), .A2(n13215), .ZN(n10674) );
  OR2_X1 U13299 ( .A1(n10674), .A2(n10842), .ZN(n14913) );
  NOR2_X1 U13300 ( .A1(n14868), .A2(n14913), .ZN(n10675) );
  NOR2_X1 U13301 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  OAI211_X1 U13302 ( .C1(n14871), .C2(n14912), .A(n10678), .B(n10677), .ZN(
        P2_U3262) );
  XNOR2_X1 U13303 ( .A(n10680), .B(n10679), .ZN(n10687) );
  NAND2_X1 U13304 ( .A1(n13111), .A2(n13444), .ZN(n10682) );
  NAND2_X1 U13305 ( .A1(n13109), .A2(n13441), .ZN(n10681) );
  AND2_X1 U13306 ( .A1(n10682), .A2(n10681), .ZN(n10866) );
  AND2_X1 U13307 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13135) );
  INV_X1 U13308 ( .A(n13135), .ZN(n10683) );
  OAI21_X1 U13309 ( .B1(n12996), .B2(n10866), .A(n10683), .ZN(n10685) );
  NOR2_X1 U13310 ( .A1(n13091), .A2(n14852), .ZN(n10684) );
  AOI211_X1 U13311 ( .C1(n10942), .C2(n13093), .A(n10685), .B(n10684), .ZN(
        n10686) );
  OAI21_X1 U13312 ( .B1(n10687), .B2(n13082), .A(n10686), .ZN(P2_U3185) );
  NAND2_X1 U13313 ( .A1(n13869), .A2(n13700), .ZN(n10691) );
  NAND2_X1 U13314 ( .A1(n14708), .A2(n13699), .ZN(n10690) );
  NAND2_X1 U13315 ( .A1(n10691), .A2(n10690), .ZN(n10693) );
  XNOR2_X1 U13316 ( .A(n10693), .B(n6937), .ZN(n10696) );
  NAND2_X1 U13317 ( .A1(n13869), .A2(n13704), .ZN(n10695) );
  NAND2_X1 U13318 ( .A1(n14708), .A2(n13700), .ZN(n10694) );
  AND2_X1 U13319 ( .A1(n10695), .A2(n10694), .ZN(n10697) );
  AND2_X1 U13320 ( .A1(n10696), .A2(n10697), .ZN(n10912) );
  INV_X1 U13321 ( .A(n10912), .ZN(n10700) );
  INV_X1 U13322 ( .A(n10696), .ZN(n10699) );
  INV_X1 U13323 ( .A(n10697), .ZN(n10698) );
  NAND2_X1 U13324 ( .A1(n10699), .A2(n10698), .ZN(n10913) );
  NAND2_X1 U13325 ( .A1(n10700), .A2(n10913), .ZN(n10701) );
  XNOR2_X1 U13326 ( .A(n6451), .B(n10701), .ZN(n10708) );
  NAND2_X1 U13327 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13934) );
  NAND2_X1 U13328 ( .A1(n14528), .A2(n13868), .ZN(n10702) );
  OAI211_X1 U13329 ( .C1(n15303), .C2(n10703), .A(n13934), .B(n10702), .ZN(
        n10706) );
  NOR2_X1 U13330 ( .A1(n14530), .A2(n10704), .ZN(n10705) );
  AOI211_X1 U13331 ( .C1(n14526), .C2(n13870), .A(n10706), .B(n10705), .ZN(
        n10707) );
  OAI21_X1 U13332 ( .B1(n10708), .B2(n15306), .A(n10707), .ZN(P1_U3227) );
  XNOR2_X1 U13333 ( .A(n10982), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10715) );
  NAND2_X1 U13334 ( .A1(n10716), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13335 ( .A1(n10712), .A2(n10711), .B1(n10710), .B2(n10709), .ZN(
        n10713) );
  XNOR2_X1 U13336 ( .A(n10713), .B(n14603), .ZN(n14599) );
  NAND2_X1 U13337 ( .A1(n14599), .A2(n9395), .ZN(n14598) );
  OAI21_X1 U13338 ( .B1(n10713), .B2(n10719), .A(n14598), .ZN(n10714) );
  NOR2_X1 U13339 ( .A1(n10714), .A2(n10715), .ZN(n10979) );
  AOI211_X1 U13340 ( .C1(n10715), .C2(n10714), .A(n13926), .B(n10979), .ZN(
        n10732) );
  NAND2_X1 U13341 ( .A1(n10716), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10717) );
  NAND2_X1 U13342 ( .A1(n10718), .A2(n10717), .ZN(n10720) );
  OR2_X1 U13343 ( .A1(n10720), .A2(n10719), .ZN(n10724) );
  INV_X1 U13344 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14189) );
  XNOR2_X1 U13345 ( .A(n10982), .B(n14189), .ZN(n10722) );
  XNOR2_X1 U13346 ( .A(n10720), .B(n10719), .ZN(n14601) );
  NOR2_X1 U13347 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14601), .ZN(n14600) );
  INV_X1 U13348 ( .A(n14600), .ZN(n10723) );
  AND2_X1 U13349 ( .A1(n10722), .A2(n10723), .ZN(n10721) );
  NAND2_X1 U13350 ( .A1(n10724), .A2(n10721), .ZN(n10988) );
  INV_X1 U13351 ( .A(n10988), .ZN(n10726) );
  AOI21_X1 U13352 ( .B1(n10724), .B2(n10723), .A(n10722), .ZN(n10725) );
  NOR3_X1 U13353 ( .A1(n10726), .A2(n10725), .A3(n14604), .ZN(n10731) );
  NAND2_X1 U13354 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14519)
         );
  INV_X1 U13355 ( .A(n14519), .ZN(n10727) );
  AOI21_X1 U13356 ( .B1(n14594), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10727), 
        .ZN(n10728) );
  OAI21_X1 U13357 ( .B1(n10729), .B2(n14602), .A(n10728), .ZN(n10730) );
  OR3_X1 U13358 ( .A1(n10732), .A2(n10731), .A3(n10730), .ZN(P1_U3259) );
  INV_X1 U13359 ( .A(n10733), .ZN(n10734) );
  AOI21_X1 U13360 ( .B1(n11987), .B2(n10735), .A(n10734), .ZN(n10793) );
  OR2_X1 U13361 ( .A1(n14656), .A2(n11985), .ZN(n14411) );
  OAI21_X1 U13362 ( .B1(n10737), .B2(n11987), .A(n10736), .ZN(n10741) );
  INV_X1 U13363 ( .A(n13870), .ZN(n10738) );
  OAI22_X1 U13364 ( .A1(n10738), .A2(n14617), .B1(n11833), .B2(n14127), .ZN(
        n10740) );
  NOR2_X1 U13365 ( .A1(n10793), .A2(n10756), .ZN(n10739) );
  AOI211_X1 U13366 ( .C1(n14403), .C2(n10741), .A(n10740), .B(n10739), .ZN(
        n10792) );
  MUX2_X1 U13367 ( .A(n10742), .B(n10792), .S(n14231), .Z(n10747) );
  AOI21_X1 U13368 ( .B1(n10885), .B2(n11839), .A(n14715), .ZN(n10743) );
  AND2_X1 U13369 ( .A1(n10744), .A2(n10743), .ZN(n10790) );
  OAI22_X1 U13370 ( .A1(n14190), .A2(n11840), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14229), .ZN(n10745) );
  AOI21_X1 U13371 ( .B1(n14633), .B2(n10790), .A(n10745), .ZN(n10746) );
  OAI211_X1 U13372 ( .C1(n10793), .C2(n14411), .A(n10747), .B(n10746), .ZN(
        P1_U3290) );
  XNOR2_X1 U13373 ( .A(n10748), .B(n10749), .ZN(n14690) );
  INV_X1 U13374 ( .A(n14690), .ZN(n10766) );
  OAI21_X1 U13375 ( .B1(n10753), .B2(n14127), .A(n14639), .ZN(n10758) );
  NAND2_X1 U13376 ( .A1(n10748), .A2(n14127), .ZN(n10755) );
  OR2_X1 U13377 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  NAND2_X1 U13378 ( .A1(n10883), .A2(n10752), .ZN(n14687) );
  XNOR2_X1 U13379 ( .A(n14687), .B(n6936), .ZN(n10754) );
  MUX2_X1 U13380 ( .A(n10755), .B(n10754), .S(n10753), .Z(n10757) );
  INV_X1 U13381 ( .A(n10756), .ZN(n14733) );
  AOI22_X1 U13382 ( .A1(n10758), .A2(n10757), .B1(n14690), .B2(n14733), .ZN(
        n10759) );
  INV_X1 U13383 ( .A(n10759), .ZN(n14688) );
  NOR2_X1 U13384 ( .A1(n11833), .A2(n14617), .ZN(n14685) );
  OAI21_X1 U13385 ( .B1(n14688), .B2(n14685), .A(n14231), .ZN(n10765) );
  OR2_X1 U13386 ( .A1(n14656), .A2(n10760), .ZN(n14024) );
  NOR2_X1 U13387 ( .A1(n14024), .A2(n14687), .ZN(n10763) );
  OAI22_X1 U13388 ( .A1(n14231), .A2(n9955), .B1(n10761), .B2(n14229), .ZN(
        n10762) );
  AOI211_X1 U13389 ( .C1(n14646), .C2(n9212), .A(n10763), .B(n10762), .ZN(
        n10764) );
  OAI211_X1 U13390 ( .C1(n10766), .C2(n14411), .A(n10765), .B(n10764), .ZN(
        P1_U3292) );
  MUX2_X1 U13391 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n11248), .Z(n11053) );
  XNOR2_X1 U13392 ( .A(n11053), .B(n11076), .ZN(n11054) );
  INV_X1 U13393 ( .A(n10767), .ZN(n10768) );
  XOR2_X1 U13394 ( .A(n11054), .B(n11055), .Z(n10788) );
  AOI22_X1 U13395 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11076), .B1(n11067), 
        .B2(n7796), .ZN(n10776) );
  NAND2_X1 U13396 ( .A1(n10772), .A2(n10771), .ZN(n10774) );
  NAND2_X1 U13397 ( .A1(n10776), .A2(n10775), .ZN(n11066) );
  OAI21_X1 U13398 ( .B1(n10776), .B2(n10775), .A(n11066), .ZN(n10786) );
  AND2_X1 U13399 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11415) );
  AOI21_X1 U13400 ( .B1(n14995), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11415), .ZN(
        n10777) );
  OAI21_X1 U13401 ( .B1(n14989), .B2(n11076), .A(n10777), .ZN(n10785) );
  AOI22_X1 U13402 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11067), .B1(n11076), 
        .B2(n11099), .ZN(n10781) );
  AOI21_X1 U13403 ( .B1(n10782), .B2(n10781), .A(n11075), .ZN(n10783) );
  NOR2_X1 U13404 ( .A1(n10783), .A2(n15001), .ZN(n10784) );
  AOI211_X1 U13405 ( .C1(n15007), .C2(n10786), .A(n10785), .B(n10784), .ZN(
        n10787) );
  OAI21_X1 U13406 ( .B1(n10788), .B2(n14991), .A(n10787), .ZN(P3_U3190) );
  NAND2_X1 U13407 ( .A1(n12352), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10789) );
  OAI21_X1 U13408 ( .B1(n12210), .B2(n12352), .A(n10789), .ZN(P3_U3520) );
  INV_X1 U13409 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n13907) );
  AOI21_X1 U13410 ( .B1(n11839), .B2(n14723), .A(n10790), .ZN(n10791) );
  OAI211_X1 U13411 ( .C1(n10793), .C2(n14729), .A(n10792), .B(n10791), .ZN(
        n10795) );
  NAND2_X1 U13412 ( .A1(n10795), .A2(n14761), .ZN(n10794) );
  OAI21_X1 U13413 ( .B1(n14761), .B2(n13907), .A(n10794), .ZN(P1_U3531) );
  INV_X1 U13414 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10797) );
  NAND2_X1 U13415 ( .A1(n10795), .A2(n14751), .ZN(n10796) );
  OAI21_X1 U13416 ( .B1(n14751), .B2(n10797), .A(n10796), .ZN(P1_U3468) );
  XNOR2_X1 U13417 ( .A(n10798), .B(n11995), .ZN(n14730) );
  AOI21_X1 U13418 ( .B1(n10800), .B2(n10799), .A(n14639), .ZN(n10804) );
  OR2_X1 U13419 ( .A1(n11266), .A2(n14617), .ZN(n10803) );
  NAND2_X1 U13420 ( .A1(n13868), .A2(n14619), .ZN(n10802) );
  NAND2_X1 U13421 ( .A1(n10803), .A2(n10802), .ZN(n11122) );
  AOI21_X1 U13422 ( .B1(n10804), .B2(n10801), .A(n11122), .ZN(n14728) );
  MUX2_X1 U13423 ( .A(n14728), .B(n10805), .S(n14656), .Z(n10809) );
  AOI21_X1 U13424 ( .B1(n14724), .B2(n14648), .A(n14631), .ZN(n14726) );
  INV_X1 U13425 ( .A(n14024), .ZN(n14652) );
  INV_X1 U13426 ( .A(n14724), .ZN(n10806) );
  OAI22_X1 U13427 ( .A1(n10806), .A2(n14190), .B1(n11124), .B2(n14229), .ZN(
        n10807) );
  AOI21_X1 U13428 ( .B1(n14726), .B2(n14652), .A(n10807), .ZN(n10808) );
  OAI211_X1 U13429 ( .C1(n14202), .C2(n14730), .A(n10809), .B(n10808), .ZN(
        P1_U3286) );
  INV_X1 U13430 ( .A(n10817), .ZN(n10810) );
  NAND2_X1 U13431 ( .A1(n10820), .A2(n14914), .ZN(n10812) );
  INV_X1 U13432 ( .A(n10836), .ZN(n10813) );
  NAND2_X1 U13433 ( .A1(n10823), .A2(n14927), .ZN(n10814) );
  NAND2_X1 U13434 ( .A1(n10815), .A2(n10814), .ZN(n10857) );
  INV_X1 U13435 ( .A(n10816), .ZN(n10826) );
  XNOR2_X1 U13436 ( .A(n10857), .B(n10826), .ZN(n14935) );
  NAND2_X1 U13437 ( .A1(n10818), .A2(n10817), .ZN(n10822) );
  NAND2_X1 U13438 ( .A1(n10820), .A2(n10819), .ZN(n10821) );
  NAND2_X1 U13439 ( .A1(n10822), .A2(n10821), .ZN(n10837) );
  NAND2_X1 U13440 ( .A1(n10837), .A2(n10836), .ZN(n10825) );
  NAND2_X1 U13441 ( .A1(n10823), .A2(n10845), .ZN(n10824) );
  NAND2_X1 U13442 ( .A1(n10825), .A2(n10824), .ZN(n10863) );
  XNOR2_X1 U13443 ( .A(n10863), .B(n10826), .ZN(n10828) );
  AOI21_X1 U13444 ( .B1(n10828), .B2(n14882), .A(n10827), .ZN(n14938) );
  MUX2_X1 U13445 ( .A(n10829), .B(n14938), .S(n13402), .Z(n10834) );
  NAND2_X1 U13446 ( .A1(n10842), .A2(n14927), .ZN(n10843) );
  AOI21_X1 U13447 ( .B1(n10843), .B2(n14931), .A(n9733), .ZN(n10830) );
  AND2_X1 U13448 ( .A1(n10830), .A2(n10960), .ZN(n14933) );
  OAI22_X1 U13449 ( .A1(n14874), .A2(n6592), .B1(n10831), .B2(n14881), .ZN(
        n10832) );
  AOI21_X1 U13450 ( .B1(n14850), .B2(n14933), .A(n10832), .ZN(n10833) );
  OAI211_X1 U13451 ( .C1(n14871), .C2(n14935), .A(n10834), .B(n10833), .ZN(
        P2_U3260) );
  XNOR2_X1 U13452 ( .A(n10835), .B(n10836), .ZN(n14921) );
  XNOR2_X1 U13453 ( .A(n10837), .B(n10836), .ZN(n10840) );
  INV_X1 U13454 ( .A(n10838), .ZN(n10839) );
  AOI21_X1 U13455 ( .B1(n10840), .B2(n14882), .A(n10839), .ZN(n14926) );
  MUX2_X1 U13456 ( .A(n10841), .B(n14926), .S(n13402), .Z(n10849) );
  INV_X1 U13457 ( .A(n10842), .ZN(n10844) );
  AOI211_X1 U13458 ( .C1(n10845), .C2(n10844), .A(n9733), .B(n6593), .ZN(
        n14924) );
  OAI22_X1 U13459 ( .A1(n14874), .A2(n14927), .B1(n14881), .B2(n10846), .ZN(
        n10847) );
  AOI21_X1 U13460 ( .B1(n14924), .B2(n14850), .A(n10847), .ZN(n10848) );
  OAI211_X1 U13461 ( .C1(n14871), .C2(n14921), .A(n10849), .B(n10848), .ZN(
        P2_U3261) );
  INV_X1 U13462 ( .A(n10850), .ZN(n10852) );
  OAI222_X1 U13463 ( .A1(n14353), .A2(n10851), .B1(n11585), .B2(n10852), .C1(
        n11525), .C2(P1_U3086), .ZN(P1_U3336) );
  OAI222_X1 U13464 ( .A1(n13588), .A2(n10853), .B1(n13590), .B2(n10852), .C1(
        P2_U3088), .C2(n13188), .ZN(P2_U3308) );
  NAND2_X1 U13465 ( .A1(n10854), .A2(n14388), .ZN(n10855) );
  OAI211_X1 U13466 ( .C1(n10856), .C2(n14376), .A(n10855), .B(n11796), .ZN(
        P3_U3272) );
  NAND2_X1 U13467 ( .A1(n13112), .A2(n14931), .ZN(n10858) );
  OR2_X1 U13468 ( .A1(n10965), .A2(n13111), .ZN(n10859) );
  OAI21_X1 U13469 ( .B1(n10860), .B2(n10865), .A(n10937), .ZN(n14858) );
  INV_X1 U13470 ( .A(n14858), .ZN(n10871) );
  NOR2_X1 U13471 ( .A1(n6592), .A2(n13112), .ZN(n10862) );
  NAND2_X1 U13472 ( .A1(n6592), .A2(n13112), .ZN(n10861) );
  XOR2_X1 U13473 ( .A(n10865), .B(n10943), .Z(n10868) );
  INV_X1 U13474 ( .A(n10866), .ZN(n10867) );
  AOI21_X1 U13475 ( .B1(n10868), .B2(n14882), .A(n10867), .ZN(n14861) );
  INV_X1 U13476 ( .A(n10869), .ZN(n10961) );
  INV_X1 U13477 ( .A(n10942), .ZN(n14856) );
  AOI211_X1 U13478 ( .C1(n10942), .C2(n10961), .A(n9733), .B(n10952), .ZN(
        n14851) );
  AOI21_X1 U13479 ( .B1(n14930), .B2(n10942), .A(n14851), .ZN(n10870) );
  OAI211_X1 U13480 ( .C1(n14934), .C2(n10871), .A(n14861), .B(n10870), .ZN(
        n10875) );
  NAND2_X1 U13481 ( .A1(n10875), .A2(n14974), .ZN(n10872) );
  OAI21_X1 U13482 ( .B1(n14974), .B2(n10873), .A(n10872), .ZN(P2_U3506) );
  NAND2_X1 U13483 ( .A1(n10875), .A2(n14959), .ZN(n10876) );
  OAI21_X1 U13484 ( .B1(n14959), .B2(n8618), .A(n10876), .ZN(P2_U3451) );
  XOR2_X1 U13485 ( .A(n11989), .B(n10877), .Z(n14696) );
  INV_X1 U13486 ( .A(n14696), .ZN(n10891) );
  OAI21_X1 U13487 ( .B1(n11989), .B2(n10879), .A(n10878), .ZN(n10881) );
  AOI21_X1 U13488 ( .B1(n10881), .B2(n14403), .A(n10880), .ZN(n10882) );
  INV_X1 U13489 ( .A(n10882), .ZN(n14694) );
  NAND2_X1 U13490 ( .A1(n10883), .A2(n11832), .ZN(n10884) );
  NAND2_X1 U13491 ( .A1(n10885), .A2(n10884), .ZN(n14693) );
  NAND2_X1 U13492 ( .A1(n14646), .A2(n11832), .ZN(n10888) );
  NOR2_X1 U13493 ( .A1(n14229), .A2(n13882), .ZN(n10886) );
  AOI21_X1 U13494 ( .B1(n14625), .B2(P1_REG2_REG_2__SCAN_IN), .A(n10886), .ZN(
        n10887) );
  OAI211_X1 U13495 ( .C1(n14693), .C2(n14024), .A(n10888), .B(n10887), .ZN(
        n10889) );
  AOI21_X1 U13496 ( .B1(n14694), .B2(n14231), .A(n10889), .ZN(n10890) );
  OAI21_X1 U13497 ( .B1(n10891), .B2(n14202), .A(n10890), .ZN(P1_U3291) );
  OAI22_X1 U13498 ( .A1(n14231), .A2(n10893), .B1(n10892), .B2(n14229), .ZN(
        n10894) );
  AOI21_X1 U13499 ( .B1(n10895), .B2(n14634), .A(n10894), .ZN(n10898) );
  OAI21_X1 U13500 ( .B1(n14646), .B2(n14652), .A(n10896), .ZN(n10897) );
  OAI211_X1 U13501 ( .C1(n14656), .C2(n10899), .A(n10898), .B(n10897), .ZN(
        P1_U3293) );
  XNOR2_X1 U13502 ( .A(n15103), .B(n12159), .ZN(n11003) );
  XNOR2_X1 U13503 ( .A(n11003), .B(n15030), .ZN(n10904) );
  NAND2_X1 U13504 ( .A1(n10900), .A2(n15067), .ZN(n10901) );
  OAI21_X1 U13505 ( .B1(n10904), .B2(n10903), .A(n11006), .ZN(n10905) );
  NAND2_X1 U13506 ( .A1(n10905), .A2(n12337), .ZN(n10911) );
  INV_X1 U13507 ( .A(n12359), .ZN(n11047) );
  OAI22_X1 U13508 ( .A1(n10906), .A2(n12340), .B1(n11047), .B2(n12327), .ZN(
        n10907) );
  AOI211_X1 U13509 ( .C1(n10909), .C2(n12330), .A(n10908), .B(n10907), .ZN(
        n10910) );
  OAI211_X1 U13510 ( .C1(n11016), .C2(n12339), .A(n10911), .B(n10910), .ZN(
        P3_U3170) );
  AOI22_X1 U13511 ( .A1(n14647), .A2(n13699), .B1(n13608), .B2(n13868), .ZN(
        n10914) );
  XNOR2_X1 U13512 ( .A(n10914), .B(n10692), .ZN(n10916) );
  AOI22_X1 U13513 ( .A1(n14647), .A2(n13608), .B1(n13704), .B2(n13868), .ZN(
        n10915) );
  INV_X1 U13514 ( .A(n11126), .ZN(n10917) );
  NAND2_X1 U13515 ( .A1(n10916), .A2(n10915), .ZN(n11125) );
  NAND2_X1 U13516 ( .A1(n10917), .A2(n11125), .ZN(n10918) );
  XNOR2_X1 U13517 ( .A(n11127), .B(n10918), .ZN(n10925) );
  INV_X1 U13518 ( .A(n10919), .ZN(n13730) );
  NAND2_X1 U13519 ( .A1(n14647), .A2(n14723), .ZN(n14714) );
  NOR2_X1 U13520 ( .A1(n13730), .A2(n14714), .ZN(n10924) );
  NAND2_X1 U13521 ( .A1(n13869), .A2(n14619), .ZN(n10921) );
  NAND2_X1 U13522 ( .A1(n14620), .A2(n14404), .ZN(n10920) );
  NAND2_X1 U13523 ( .A1(n10921), .A2(n10920), .ZN(n14642) );
  AND2_X1 U13524 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n13950) );
  AOI21_X1 U13525 ( .B1(n15299), .B2(n14642), .A(n13950), .ZN(n10922) );
  OAI21_X1 U13526 ( .B1(n15303), .B2(n14643), .A(n10922), .ZN(n10923) );
  AOI211_X1 U13527 ( .C1(n10925), .C2(n14532), .A(n10924), .B(n10923), .ZN(
        n10926) );
  INV_X1 U13528 ( .A(n10926), .ZN(P1_U3239) );
  OAI21_X1 U13529 ( .B1(n10929), .B2(n10928), .A(n10927), .ZN(n10931) );
  XOR2_X1 U13530 ( .A(n10931), .B(n10930), .Z(n10935) );
  AOI22_X1 U13531 ( .A1(n13078), .A2(n13110), .B1(n13046), .B2(n13108), .ZN(
        n10932) );
  NAND2_X1 U13532 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14814) );
  OAI211_X1 U13533 ( .C1(n10950), .C2(n13091), .A(n10932), .B(n14814), .ZN(
        n10933) );
  AOI21_X1 U13534 ( .B1(n11109), .B2(n13093), .A(n10933), .ZN(n10934) );
  OAI21_X1 U13535 ( .B1(n10935), .B2(n13082), .A(n10934), .ZN(P2_U3193) );
  OR2_X1 U13536 ( .A1(n10942), .A2(n13110), .ZN(n10936) );
  NAND2_X1 U13537 ( .A1(n10938), .A2(n10946), .ZN(n10939) );
  NAND2_X1 U13538 ( .A1(n11111), .A2(n10939), .ZN(n14946) );
  INV_X1 U13539 ( .A(n10940), .ZN(n14888) );
  NAND2_X1 U13540 ( .A1(n13402), .A2(n14888), .ZN(n11470) );
  AOI22_X1 U13541 ( .A1(n13444), .A2(n13110), .B1(n13108), .B2(n13441), .ZN(
        n10949) );
  NAND2_X1 U13542 ( .A1(n10943), .A2(n10942), .ZN(n10944) );
  NAND2_X1 U13543 ( .A1(n10945), .A2(n10944), .ZN(n11105) );
  XNOR2_X1 U13544 ( .A(n11105), .B(n10946), .ZN(n10947) );
  NAND2_X1 U13545 ( .A1(n10947), .A2(n14882), .ZN(n10948) );
  OAI211_X1 U13546 ( .C1(n14946), .C2(n14922), .A(n10949), .B(n10948), .ZN(
        n14949) );
  NAND2_X1 U13547 ( .A1(n14949), .A2(n13402), .ZN(n10956) );
  INV_X1 U13548 ( .A(n14874), .ZN(n13433) );
  OAI22_X1 U13549 ( .A1(n13402), .A2(n10951), .B1(n10950), .B2(n14881), .ZN(
        n10954) );
  INV_X1 U13550 ( .A(n11109), .ZN(n14948) );
  OAI211_X1 U13551 ( .C1(n10952), .C2(n14948), .A(n13215), .B(n11115), .ZN(
        n14947) );
  NOR2_X1 U13552 ( .A1(n14947), .A2(n14868), .ZN(n10953) );
  AOI211_X1 U13553 ( .C1(n13433), .C2(n11109), .A(n10954), .B(n10953), .ZN(
        n10955) );
  OAI211_X1 U13554 ( .C1(n14946), .C2(n11470), .A(n10956), .B(n10955), .ZN(
        P2_U3257) );
  INV_X1 U13555 ( .A(n11470), .ZN(n10977) );
  NAND2_X1 U13556 ( .A1(n10957), .A2(n7447), .ZN(n10958) );
  NAND2_X1 U13557 ( .A1(n10959), .A2(n10958), .ZN(n14944) );
  INV_X1 U13558 ( .A(n10965), .ZN(n14941) );
  INV_X1 U13559 ( .A(n10960), .ZN(n10962) );
  OAI211_X1 U13560 ( .C1(n14941), .C2(n10962), .A(n10961), .B(n13215), .ZN(
        n14940) );
  INV_X1 U13561 ( .A(n10963), .ZN(n10964) );
  AOI22_X1 U13562 ( .A1(n13433), .A2(n10965), .B1(n14865), .B2(n10964), .ZN(
        n10966) );
  OAI21_X1 U13563 ( .B1(n14940), .B2(n14868), .A(n10966), .ZN(n10976) );
  INV_X1 U13564 ( .A(n14922), .ZN(n14883) );
  NAND2_X1 U13565 ( .A1(n14944), .A2(n14883), .ZN(n10974) );
  AOI22_X1 U13566 ( .A1(n13444), .A2(n13112), .B1(n13110), .B2(n13441), .ZN(
        n10973) );
  NAND2_X1 U13567 ( .A1(n10968), .A2(n10967), .ZN(n10969) );
  NAND2_X1 U13568 ( .A1(n10970), .A2(n10969), .ZN(n10971) );
  NAND2_X1 U13569 ( .A1(n10971), .A2(n14882), .ZN(n10972) );
  NAND3_X1 U13570 ( .A1(n10974), .A2(n10973), .A3(n10972), .ZN(n14942) );
  MUX2_X1 U13571 ( .A(n14942), .B(P2_REG2_REG_6__SCAN_IN), .S(n14890), .Z(
        n10975) );
  AOI211_X1 U13572 ( .C1(n10977), .C2(n14944), .A(n10976), .B(n10975), .ZN(
        n10978) );
  INV_X1 U13573 ( .A(n10978), .ZN(P2_U3259) );
  AOI21_X1 U13574 ( .B1(n10982), .B2(P1_REG1_REG_16__SCAN_IN), .A(n10979), 
        .ZN(n10981) );
  XNOR2_X1 U13575 ( .A(n11322), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10980) );
  NOR2_X1 U13576 ( .A1(n10981), .A2(n10980), .ZN(n11321) );
  AOI211_X1 U13577 ( .C1(n10981), .C2(n10980), .A(n13926), .B(n11321), .ZN(
        n10993) );
  NAND2_X1 U13578 ( .A1(n10982), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n10984) );
  OAI21_X1 U13579 ( .B1(n11322), .B2(n14176), .A(n10984), .ZN(n10983) );
  AOI21_X1 U13580 ( .B1(n11322), .B2(n14176), .A(n10983), .ZN(n10989) );
  NAND2_X1 U13581 ( .A1(n10988), .A2(n10984), .ZN(n10986) );
  NAND2_X1 U13582 ( .A1(n11320), .A2(n14176), .ZN(n10985) );
  OAI211_X1 U13583 ( .C1(n14176), .C2(n11320), .A(n10986), .B(n10985), .ZN(
        n11319) );
  INV_X1 U13584 ( .A(n11319), .ZN(n10987) );
  AOI211_X1 U13585 ( .C1(n10989), .C2(n10988), .A(n14604), .B(n10987), .ZN(
        n10992) );
  NAND2_X1 U13586 ( .A1(n14594), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n10990) );
  NAND2_X1 U13587 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13798)
         );
  OAI211_X1 U13588 ( .C1(n14602), .C2(n11320), .A(n10990), .B(n13798), .ZN(
        n10991) );
  OR3_X1 U13589 ( .A1(n10993), .A2(n10992), .A3(n10991), .ZN(P1_U3260) );
  INV_X1 U13590 ( .A(n14871), .ZN(n14859) );
  NAND2_X1 U13591 ( .A1(n14859), .A2(n10994), .ZN(n10998) );
  OAI22_X1 U13592 ( .A1(n13402), .A2(n10097), .B1(n10995), .B2(n14881), .ZN(
        n10996) );
  AOI21_X1 U13593 ( .B1(n13433), .B2(n13048), .A(n10996), .ZN(n10997) );
  OAI211_X1 U13594 ( .C1(n10999), .C2(n14868), .A(n10998), .B(n10997), .ZN(
        n11000) );
  AOI21_X1 U13595 ( .B1(n13402), .B2(n11001), .A(n11000), .ZN(n11002) );
  INV_X1 U13596 ( .A(n11002), .ZN(P2_U3263) );
  INV_X1 U13597 ( .A(n11003), .ZN(n11004) );
  OR2_X1 U13598 ( .A1(n15030), .A2(n11004), .ZN(n11005) );
  XNOR2_X1 U13599 ( .A(n11007), .B(n10597), .ZN(n11040) );
  XNOR2_X1 U13600 ( .A(n11040), .B(n12359), .ZN(n11038) );
  XOR2_X1 U13601 ( .A(n11039), .B(n11038), .Z(n11013) );
  INV_X1 U13602 ( .A(n11008), .ZN(n15036) );
  AOI22_X1 U13603 ( .A1(n12323), .A2(n15030), .B1(n12344), .B2(n15029), .ZN(
        n11010) );
  OAI211_X1 U13604 ( .C1(n12347), .C2(n15035), .A(n11010), .B(n11009), .ZN(
        n11011) );
  AOI21_X1 U13605 ( .B1(n15036), .B2(n12324), .A(n11011), .ZN(n11012) );
  OAI21_X1 U13606 ( .B1(n11013), .B2(n12332), .A(n11012), .ZN(P3_U3167) );
  OAI222_X1 U13607 ( .A1(n11585), .A2(n11587), .B1(P1_U3086), .B2(n11981), 
        .C1(n11014), .C2(n14353), .ZN(P1_U3335) );
  XNOR2_X1 U13608 ( .A(n11015), .B(n11759), .ZN(n15106) );
  OAI22_X1 U13609 ( .A1(n12691), .A2(n15103), .B1(n11016), .B2(n15083), .ZN(
        n11023) );
  XNOR2_X1 U13610 ( .A(n11017), .B(n11018), .ZN(n11021) );
  NAND2_X1 U13611 ( .A1(n15106), .A2(n15031), .ZN(n11020) );
  AOI22_X1 U13612 ( .A1(n15069), .A2(n15067), .B1(n12359), .B2(n15066), .ZN(
        n11019) );
  OAI211_X1 U13613 ( .C1(n15043), .C2(n11021), .A(n11020), .B(n11019), .ZN(
        n15104) );
  MUX2_X1 U13614 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n15104), .S(n15091), .Z(
        n11022) );
  AOI211_X1 U13615 ( .C1(n15106), .C2(n12544), .A(n11023), .B(n11022), .ZN(
        n11024) );
  INV_X1 U13616 ( .A(n11024), .ZN(P3_U3229) );
  INV_X1 U13617 ( .A(n11025), .ZN(n11026) );
  AOI21_X1 U13618 ( .B1(n11030), .B2(n11027), .A(n11026), .ZN(n11028) );
  AOI22_X1 U13619 ( .A1(n13867), .A2(n14619), .B1(n14404), .B2(n14525), .ZN(
        n11282) );
  OAI21_X1 U13620 ( .B1(n11028), .B2(n14639), .A(n11282), .ZN(n11297) );
  INV_X1 U13621 ( .A(n11297), .ZN(n11037) );
  OAI21_X1 U13622 ( .B1(n11031), .B2(n11030), .A(n11029), .ZN(n11299) );
  OAI211_X1 U13623 ( .C1(n14629), .C2(n11873), .A(n14725), .B(n11177), .ZN(
        n11296) );
  NOR2_X1 U13624 ( .A1(n11296), .A2(n14216), .ZN(n11035) );
  INV_X1 U13625 ( .A(n11032), .ZN(n11284) );
  INV_X1 U13626 ( .A(n14229), .ZN(n14645) );
  AOI22_X1 U13627 ( .A1(n14625), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11284), 
        .B2(n14645), .ZN(n11033) );
  OAI21_X1 U13628 ( .B1(n11873), .B2(n14190), .A(n11033), .ZN(n11034) );
  AOI211_X1 U13629 ( .C1(n11299), .C2(n14634), .A(n11035), .B(n11034), .ZN(
        n11036) );
  OAI21_X1 U13630 ( .B1(n11037), .B2(n14656), .A(n11036), .ZN(P1_U3284) );
  INV_X1 U13631 ( .A(n11040), .ZN(n11041) );
  OR2_X1 U13632 ( .A1(n11041), .A2(n12359), .ZN(n11042) );
  XNOR2_X1 U13633 ( .A(n11050), .B(n12159), .ZN(n11287) );
  XNOR2_X1 U13634 ( .A(n11287), .B(n15029), .ZN(n11044) );
  AOI21_X1 U13635 ( .B1(n11043), .B2(n11044), .A(n12332), .ZN(n11046) );
  INV_X1 U13636 ( .A(n11044), .ZN(n11045) );
  NAND2_X1 U13637 ( .A1(n11046), .A2(n11289), .ZN(n11052) );
  INV_X1 U13638 ( .A(n12358), .ZN(n11413) );
  OAI22_X1 U13639 ( .A1(n11047), .A2(n12340), .B1(n11413), .B2(n12327), .ZN(
        n11048) );
  AOI211_X1 U13640 ( .C1(n11050), .C2(n12330), .A(n11049), .B(n11048), .ZN(
        n11051) );
  OAI211_X1 U13641 ( .C1(n11334), .C2(n12339), .A(n11052), .B(n11051), .ZN(
        P3_U3179) );
  OAI22_X1 U13642 ( .A1(n11055), .A2(n11054), .B1(n11053), .B2(n11076), .ZN(
        n14985) );
  MUX2_X1 U13643 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n11248), .Z(n11056) );
  NAND2_X1 U13644 ( .A1(n11056), .A2(n14990), .ZN(n14986) );
  INV_X1 U13645 ( .A(n11056), .ZN(n11057) );
  NAND2_X1 U13646 ( .A1(n11057), .A2(n11078), .ZN(n15012) );
  INV_X1 U13647 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11080) );
  MUX2_X1 U13648 ( .A(n11080), .B(n11070), .S(n11248), .Z(n11059) );
  NAND2_X1 U13649 ( .A1(n11059), .A2(n15018), .ZN(n11063) );
  INV_X1 U13650 ( .A(n11059), .ZN(n11061) );
  INV_X1 U13651 ( .A(n15018), .ZN(n11060) );
  NAND2_X1 U13652 ( .A1(n11061), .A2(n11060), .ZN(n11062) );
  NAND2_X1 U13653 ( .A1(n11063), .A2(n11062), .ZN(n15011) );
  INV_X1 U13654 ( .A(n11063), .ZN(n11064) );
  MUX2_X1 U13655 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n11248), .Z(n11247) );
  XNOR2_X1 U13656 ( .A(n11247), .B(n14375), .ZN(n11065) );
  AOI21_X1 U13657 ( .B1(n6474), .B2(n11065), .A(n11251), .ZN(n11088) );
  NAND2_X1 U13658 ( .A1(n14990), .A2(n11068), .ZN(n11069) );
  NAND2_X1 U13659 ( .A1(n11069), .A2(n14996), .ZN(n15005) );
  MUX2_X1 U13660 ( .A(n11070), .B(P3_REG1_REG_10__SCAN_IN), .S(n15018), .Z(
        n15004) );
  NAND2_X1 U13661 ( .A1(n15005), .A2(n15004), .ZN(n15003) );
  OAI21_X1 U13662 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11071), .A(n11255), 
        .ZN(n11086) );
  NAND2_X1 U13663 ( .A1(n15017), .A2(n11241), .ZN(n11073) );
  INV_X1 U13664 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11072) );
  OR2_X1 U13665 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11072), .ZN(n12303) );
  OAI211_X1 U13666 ( .C1(n11074), .C2(n15024), .A(n11073), .B(n12303), .ZN(
        n11085) );
  NOR2_X1 U13667 ( .A1(n11078), .A2(n11077), .ZN(n11079) );
  MUX2_X1 U13668 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n11080), .S(n15018), .Z(
        n15009) );
  OR2_X1 U13669 ( .A1(n15018), .A2(n11080), .ZN(n11081) );
  AOI21_X1 U13670 ( .B1(n7844), .B2(n11082), .A(n11242), .ZN(n11083) );
  NOR2_X1 U13671 ( .A1(n11083), .A2(n15001), .ZN(n11084) );
  AOI211_X1 U13672 ( .C1(n15007), .C2(n11086), .A(n11085), .B(n11084), .ZN(
        n11087) );
  OAI21_X1 U13673 ( .B1(n11088), .B2(n14991), .A(n11087), .ZN(P3_U3193) );
  XNOR2_X1 U13674 ( .A(n11089), .B(n11761), .ZN(n15122) );
  NAND2_X1 U13675 ( .A1(n11090), .A2(n11761), .ZN(n11091) );
  NAND2_X1 U13676 ( .A1(n11092), .A2(n11091), .ZN(n11093) );
  NAND2_X1 U13677 ( .A1(n11093), .A2(n15072), .ZN(n11095) );
  AOI22_X1 U13678 ( .A1(n15069), .A2(n12358), .B1(n12356), .B2(n15066), .ZN(
        n11094) );
  NAND2_X1 U13679 ( .A1(n11095), .A2(n11094), .ZN(n11096) );
  AOI21_X1 U13680 ( .B1(n15122), .B2(n15031), .A(n11096), .ZN(n15124) );
  INV_X2 U13681 ( .A(n15091), .ZN(n15093) );
  NOR2_X1 U13682 ( .A1(n11410), .A2(n15111), .ZN(n15121) );
  AOI22_X1 U13683 ( .A1(n15058), .A2(n15121), .B1(n15053), .B2(n11097), .ZN(
        n11098) );
  OAI21_X1 U13684 ( .B1(n11099), .B2(n15091), .A(n11098), .ZN(n11100) );
  AOI21_X1 U13685 ( .B1(n15122), .B2(n12544), .A(n11100), .ZN(n11101) );
  OAI21_X1 U13686 ( .B1(n15124), .B2(n15093), .A(n11101), .ZN(P3_U3225) );
  INV_X1 U13687 ( .A(n11102), .ZN(n11103) );
  OAI222_X1 U13688 ( .A1(n11104), .A2(P3_U3151), .B1(n14378), .B2(n11103), 
        .C1(n15242), .C2(n14376), .ZN(P3_U3271) );
  NAND2_X1 U13689 ( .A1(n11105), .A2(n11109), .ZN(n11106) );
  NAND2_X1 U13690 ( .A1(n11106), .A2(n13109), .ZN(n11107) );
  NAND2_X1 U13691 ( .A1(n11108), .A2(n11107), .ZN(n11156) );
  XNOR2_X1 U13692 ( .A(n11156), .B(n11153), .ZN(n11114) );
  NAND2_X1 U13693 ( .A1(n11109), .A2(n13109), .ZN(n11110) );
  XNOR2_X1 U13694 ( .A(n11154), .B(n11153), .ZN(n11235) );
  AOI22_X1 U13695 ( .A1(n13444), .A2(n13109), .B1(n13107), .B2(n13441), .ZN(
        n11112) );
  OAI21_X1 U13696 ( .B1(n11235), .B2(n14922), .A(n11112), .ZN(n11113) );
  AOI21_X1 U13697 ( .B1(n11114), .B2(n14882), .A(n11113), .ZN(n11234) );
  INV_X1 U13698 ( .A(n11163), .ZN(n11164) );
  AOI211_X1 U13699 ( .C1(n11232), .C2(n11115), .A(n9733), .B(n11164), .ZN(
        n11231) );
  INV_X1 U13700 ( .A(n11232), .ZN(n11118) );
  INV_X1 U13701 ( .A(n11142), .ZN(n11116) );
  AOI22_X1 U13702 ( .A1(n14890), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11116), 
        .B2(n14865), .ZN(n11117) );
  OAI21_X1 U13703 ( .B1(n11118), .B2(n14874), .A(n11117), .ZN(n11120) );
  NOR2_X1 U13704 ( .A1(n11235), .A2(n11470), .ZN(n11119) );
  AOI211_X1 U13705 ( .C1(n11231), .C2(n14850), .A(n11120), .B(n11119), .ZN(
        n11121) );
  OAI21_X1 U13706 ( .B1(n13456), .B2(n11234), .A(n11121), .ZN(P2_U3256) );
  NAND2_X1 U13707 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13961) );
  NAND2_X1 U13708 ( .A1(n11122), .A2(n15299), .ZN(n11123) );
  OAI211_X1 U13709 ( .C1(n15303), .C2(n11124), .A(n13961), .B(n11123), .ZN(
        n11134) );
  AND2_X1 U13710 ( .A1(n14620), .A2(n13704), .ZN(n11128) );
  NAND2_X1 U13711 ( .A1(n14724), .A2(n13699), .ZN(n11130) );
  NAND2_X1 U13712 ( .A1(n14620), .A2(n13700), .ZN(n11129) );
  NAND2_X1 U13713 ( .A1(n11130), .A2(n11129), .ZN(n11131) );
  XNOR2_X1 U13714 ( .A(n11131), .B(n10692), .ZN(n11269) );
  XOR2_X1 U13715 ( .A(n11269), .B(n11271), .Z(n11272) );
  XNOR2_X1 U13716 ( .A(n11273), .B(n11272), .ZN(n11132) );
  NOR2_X1 U13717 ( .A1(n11132), .A2(n15306), .ZN(n11133) );
  AOI211_X1 U13718 ( .C1(n15311), .C2(n14724), .A(n11134), .B(n11133), .ZN(
        n11135) );
  INV_X1 U13719 ( .A(n11135), .ZN(P1_U3213) );
  INV_X1 U13720 ( .A(n6895), .ZN(n12019) );
  OAI222_X1 U13721 ( .A1(n11585), .A2(n11138), .B1(P1_U3086), .B2(n12019), 
        .C1(n11136), .C2(n14353), .ZN(P1_U3334) );
  OAI222_X1 U13722 ( .A1(n13588), .A2(n11139), .B1(n13590), .B2(n11138), .C1(
        n11137), .C2(P2_U3088), .ZN(P2_U3306) );
  NOR2_X1 U13723 ( .A1(n13075), .A2(n11146), .ZN(n11140) );
  AOI22_X1 U13724 ( .A1(n11141), .A2(n13085), .B1(n11140), .B2(n10930), .ZN(
        n11152) );
  NAND2_X1 U13725 ( .A1(n13046), .A2(n13107), .ZN(n11145) );
  NAND2_X1 U13726 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14846) );
  OAI21_X1 U13727 ( .B1(n13091), .B2(n11142), .A(n14846), .ZN(n11143) );
  INV_X1 U13728 ( .A(n11143), .ZN(n11144) );
  OAI211_X1 U13729 ( .C1(n11146), .C2(n13039), .A(n11145), .B(n11144), .ZN(
        n11149) );
  NOR2_X1 U13730 ( .A1(n11147), .A2(n13082), .ZN(n11148) );
  AOI211_X1 U13731 ( .C1(n11232), .C2(n13093), .A(n11149), .B(n11148), .ZN(
        n11150) );
  OAI21_X1 U13732 ( .B1(n11152), .B2(n11151), .A(n11150), .ZN(P2_U3203) );
  XNOR2_X1 U13733 ( .A(n11376), .B(n11378), .ZN(n14956) );
  INV_X1 U13734 ( .A(n14956), .ZN(n11169) );
  NAND2_X1 U13735 ( .A1(n11156), .A2(n11155), .ZN(n11158) );
  INV_X1 U13736 ( .A(n13108), .ZN(n11188) );
  OR2_X1 U13737 ( .A1(n11232), .A2(n11188), .ZN(n11157) );
  NAND2_X1 U13738 ( .A1(n11158), .A2(n11157), .ZN(n11379) );
  XNOR2_X1 U13739 ( .A(n11379), .B(n11378), .ZN(n11161) );
  AOI22_X1 U13740 ( .A1(n13444), .A2(n13108), .B1(n13106), .B2(n13441), .ZN(
        n11160) );
  NAND2_X1 U13741 ( .A1(n14956), .A2(n14883), .ZN(n11159) );
  OAI211_X1 U13742 ( .C1(n11161), .C2(n13424), .A(n11160), .B(n11159), .ZN(
        n14954) );
  NAND2_X1 U13743 ( .A1(n14954), .A2(n13402), .ZN(n11168) );
  OAI22_X1 U13744 ( .A1(n13402), .A2(n11162), .B1(n11187), .B2(n14881), .ZN(
        n11166) );
  OAI211_X1 U13745 ( .C1(n11164), .C2(n7141), .A(n13215), .B(n11386), .ZN(
        n14952) );
  NOR2_X1 U13746 ( .A1(n14952), .A2(n14868), .ZN(n11165) );
  AOI211_X1 U13747 ( .C1(n13433), .C2(n11380), .A(n11166), .B(n11165), .ZN(
        n11167) );
  OAI211_X1 U13748 ( .C1(n11169), .C2(n11470), .A(n11168), .B(n11167), .ZN(
        P2_U3255) );
  OAI211_X1 U13749 ( .C1(n11171), .C2(n11998), .A(n11170), .B(n14403), .ZN(
        n11173) );
  OR2_X1 U13750 ( .A1(n14618), .A2(n14127), .ZN(n11172) );
  NAND2_X1 U13751 ( .A1(n11173), .A2(n11172), .ZN(n14745) );
  INV_X1 U13752 ( .A(n14745), .ZN(n11184) );
  OAI21_X1 U13753 ( .B1(n11176), .B2(n11175), .A(n11174), .ZN(n14747) );
  AOI211_X1 U13754 ( .C1(n14741), .C2(n11177), .A(n14715), .B(n6574), .ZN(
        n11178) );
  AOI21_X1 U13755 ( .B1(n14404), .B2(n14406), .A(n11178), .ZN(n14742) );
  OAI22_X1 U13756 ( .A1(n14231), .A2(n11179), .B1(n11362), .B2(n14229), .ZN(
        n11180) );
  AOI21_X1 U13757 ( .B1(n14741), .B2(n14646), .A(n11180), .ZN(n11181) );
  OAI21_X1 U13758 ( .B1(n14742), .B2(n14216), .A(n11181), .ZN(n11182) );
  AOI21_X1 U13759 ( .B1(n14747), .B2(n14634), .A(n11182), .ZN(n11183) );
  OAI21_X1 U13760 ( .B1(n14625), .B2(n11184), .A(n11183), .ZN(P1_U3283) );
  OAI211_X1 U13761 ( .C1(n11186), .C2(n11185), .A(n11396), .B(n13085), .ZN(
        n11193) );
  INV_X1 U13762 ( .A(n11187), .ZN(n11191) );
  OAI22_X1 U13763 ( .A1(n13072), .A2(n11455), .B1(n11188), .B2(n13039), .ZN(
        n11189) );
  AOI211_X1 U13764 ( .C1(n11191), .C2(n13070), .A(n11190), .B(n11189), .ZN(
        n11192) );
  OAI211_X1 U13765 ( .C1(n7141), .C2(n13023), .A(n11193), .B(n11192), .ZN(
        P2_U3189) );
  NAND2_X1 U13766 ( .A1(n11204), .A2(n11194), .ZN(n11197) );
  OR2_X1 U13767 ( .A1(n11195), .A2(n13431), .ZN(n11196) );
  NAND2_X1 U13768 ( .A1(n11197), .A2(n11196), .ZN(n11199) );
  NAND2_X1 U13769 ( .A1(n11198), .A2(n11199), .ZN(n11200) );
  XNOR2_X1 U13770 ( .A(n13150), .B(n11199), .ZN(n13154) );
  NAND2_X1 U13771 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n13154), .ZN(n13153) );
  NAND2_X1 U13772 ( .A1(n11200), .A2(n13153), .ZN(n11202) );
  MUX2_X1 U13773 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n13401), .S(n11434), .Z(
        n11201) );
  OAI21_X1 U13774 ( .B1(n11202), .B2(n11201), .A(n14838), .ZN(n11216) );
  NOR2_X1 U13775 ( .A1(n11205), .A2(n13150), .ZN(n11207) );
  XNOR2_X1 U13776 ( .A(n11205), .B(n13150), .ZN(n13146) );
  NOR2_X1 U13777 ( .A1(n11206), .A2(n13146), .ZN(n13147) );
  XNOR2_X1 U13778 ( .A(n11434), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n11208) );
  NOR2_X1 U13779 ( .A1(n11209), .A2(n11208), .ZN(n11431) );
  AOI211_X1 U13780 ( .C1(n11209), .C2(n11208), .A(n14844), .B(n11431), .ZN(
        n11210) );
  INV_X1 U13781 ( .A(n11210), .ZN(n11215) );
  NOR2_X1 U13782 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15197), .ZN(n11213) );
  NOR2_X1 U13783 ( .A1(n14794), .A2(n11211), .ZN(n11212) );
  AOI211_X1 U13784 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n14762), .A(n11213), 
        .B(n11212), .ZN(n11214) );
  OAI211_X1 U13785 ( .C1(n11440), .C2(n11216), .A(n11215), .B(n11214), .ZN(
        P2_U3230) );
  INV_X1 U13786 ( .A(n11217), .ZN(n11218) );
  OAI222_X1 U13787 ( .A1(P3_U3151), .A2(n11219), .B1(n14378), .B2(n11218), 
        .C1(n7493), .C2(n14376), .ZN(P3_U3270) );
  XNOR2_X1 U13788 ( .A(n11220), .B(n11760), .ZN(n15127) );
  NAND2_X1 U13789 ( .A1(n11221), .A2(n11760), .ZN(n11222) );
  NAND3_X1 U13790 ( .A1(n11223), .A2(n15072), .A3(n11222), .ZN(n11225) );
  AOI22_X1 U13791 ( .A1(n15069), .A2(n12357), .B1(n14467), .B2(n15066), .ZN(
        n11224) );
  NAND2_X1 U13792 ( .A1(n11225), .A2(n11224), .ZN(n11226) );
  AOI21_X1 U13793 ( .B1(n15127), .B2(n15031), .A(n11226), .ZN(n15129) );
  NOR2_X1 U13794 ( .A1(n11529), .A2(n15111), .ZN(n15126) );
  INV_X1 U13795 ( .A(n11227), .ZN(n11542) );
  AOI22_X1 U13796 ( .A1(n15058), .A2(n15126), .B1(n15053), .B2(n11542), .ZN(
        n11228) );
  OAI21_X1 U13797 ( .B1(n14984), .B2(n15091), .A(n11228), .ZN(n11229) );
  AOI21_X1 U13798 ( .B1(n15127), .B2(n12544), .A(n11229), .ZN(n11230) );
  OAI21_X1 U13799 ( .B1(n15129), .B2(n15093), .A(n11230), .ZN(P3_U3224) );
  AOI21_X1 U13800 ( .B1(n14930), .B2(n11232), .A(n11231), .ZN(n11233) );
  OAI211_X1 U13801 ( .C1(n11235), .C2(n14923), .A(n11234), .B(n11233), .ZN(
        n11237) );
  NAND2_X1 U13802 ( .A1(n11237), .A2(n14974), .ZN(n11236) );
  OAI21_X1 U13803 ( .B1(n14974), .B2(n8663), .A(n11236), .ZN(P2_U3508) );
  INV_X1 U13804 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11239) );
  NAND2_X1 U13805 ( .A1(n11237), .A2(n14959), .ZN(n11238) );
  OAI21_X1 U13806 ( .B1(n14959), .B2(n11239), .A(n11238), .ZN(P2_U3457) );
  NOR2_X1 U13807 ( .A1(n11241), .A2(n11240), .ZN(n11243) );
  MUX2_X1 U13808 ( .A(n12693), .B(P3_REG2_REG_12__SCAN_IN), .S(n11478), .Z(
        n11245) );
  INV_X1 U13809 ( .A(n11472), .ZN(n11244) );
  AOI21_X1 U13810 ( .B1(n11246), .B2(n11245), .A(n11244), .ZN(n11265) );
  NOR2_X1 U13811 ( .A1(n11247), .A2(n14375), .ZN(n11250) );
  MUX2_X1 U13812 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n11248), .Z(n11475) );
  XNOR2_X1 U13813 ( .A(n11475), .B(n11478), .ZN(n11249) );
  NOR3_X1 U13814 ( .A1(n11251), .A2(n11250), .A3(n11249), .ZN(n11474) );
  INV_X1 U13815 ( .A(n11474), .ZN(n11253) );
  OAI21_X1 U13816 ( .B1(n11251), .B2(n11250), .A(n11249), .ZN(n11252) );
  NAND3_X1 U13817 ( .A1(n11253), .A2(n15015), .A3(n11252), .ZN(n11264) );
  NAND2_X1 U13818 ( .A1(n14375), .A2(n11254), .ZN(n11256) );
  NAND2_X1 U13819 ( .A1(n11256), .A2(n11255), .ZN(n11259) );
  MUX2_X1 U13820 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n11257), .S(n11478), .Z(
        n11258) );
  NAND2_X1 U13821 ( .A1(n11259), .A2(n11258), .ZN(n11479) );
  OAI21_X1 U13822 ( .B1(n11259), .B2(n11258), .A(n11479), .ZN(n11262) );
  AND2_X1 U13823 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12232) );
  AOI21_X1 U13824 ( .B1(n14995), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12232), 
        .ZN(n11260) );
  OAI21_X1 U13825 ( .B1(n14989), .B2(n11478), .A(n11260), .ZN(n11261) );
  AOI21_X1 U13826 ( .B1(n11262), .B2(n15007), .A(n11261), .ZN(n11263) );
  OAI211_X1 U13827 ( .C1(n11265), .C2(n15001), .A(n11264), .B(n11263), .ZN(
        P3_U3194) );
  OAI22_X1 U13828 ( .A1(n14737), .A2(n13752), .B1(n11266), .B2(n13749), .ZN(
        n11274) );
  INV_X1 U13829 ( .A(n11274), .ZN(n11276) );
  NOR2_X1 U13830 ( .A1(n11266), .A2(n13752), .ZN(n11267) );
  AOI21_X1 U13831 ( .B1(n15310), .B2(n13699), .A(n11267), .ZN(n11268) );
  INV_X1 U13832 ( .A(n11269), .ZN(n11270) );
  XOR2_X1 U13833 ( .A(n11274), .B(n11275), .Z(n15305) );
  OAI22_X1 U13834 ( .A1(n11873), .A2(n13752), .B1(n14618), .B2(n13749), .ZN(
        n11354) );
  OAI22_X1 U13835 ( .A1(n11873), .A2(n13754), .B1(n14618), .B2(n13752), .ZN(
        n11277) );
  XNOR2_X1 U13836 ( .A(n11277), .B(n10692), .ZN(n11355) );
  XOR2_X1 U13837 ( .A(n11354), .B(n11355), .Z(n11278) );
  OAI211_X1 U13838 ( .C1(n11279), .C2(n11278), .A(n11356), .B(n14532), .ZN(
        n11286) );
  OAI21_X1 U13839 ( .B1(n11282), .B2(n11281), .A(n11280), .ZN(n11283) );
  AOI21_X1 U13840 ( .B1(n11284), .B2(n13843), .A(n11283), .ZN(n11285) );
  OAI211_X1 U13841 ( .C1(n11873), .C2(n14530), .A(n11286), .B(n11285), .ZN(
        P1_U3231) );
  NAND2_X1 U13842 ( .A1(n11287), .A2(n15029), .ZN(n11288) );
  XNOR2_X1 U13843 ( .A(n11658), .B(n12159), .ZN(n11406) );
  OAI211_X1 U13844 ( .C1(n11290), .C2(n11406), .A(n11409), .B(n12337), .ZN(
        n11295) );
  INV_X1 U13845 ( .A(n12357), .ZN(n11539) );
  OAI22_X1 U13846 ( .A1(n6609), .A2(n12340), .B1(n11539), .B2(n12327), .ZN(
        n11291) );
  AOI211_X1 U13847 ( .C1(n11293), .C2(n12330), .A(n11292), .B(n11291), .ZN(
        n11294) );
  OAI211_X1 U13848 ( .C1(n11313), .C2(n12339), .A(n11295), .B(n11294), .ZN(
        P3_U3153) );
  INV_X1 U13849 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11301) );
  OAI21_X1 U13850 ( .B1(n11873), .B2(n14743), .A(n11296), .ZN(n11298) );
  AOI211_X1 U13851 ( .C1(n14748), .C2(n11299), .A(n11298), .B(n11297), .ZN(
        n11302) );
  OR2_X1 U13852 ( .A1(n11302), .A2(n14749), .ZN(n11300) );
  OAI21_X1 U13853 ( .B1(n14751), .B2(n11301), .A(n11300), .ZN(P1_U3486) );
  OR2_X1 U13854 ( .A1(n11302), .A2(n14759), .ZN(n11303) );
  OAI21_X1 U13855 ( .B1(n14761), .B2(n9315), .A(n11303), .ZN(P1_U3537) );
  XNOR2_X1 U13856 ( .A(n11304), .B(n11763), .ZN(n15119) );
  INV_X1 U13857 ( .A(n15119), .ZN(n11318) );
  INV_X1 U13858 ( .A(n12544), .ZN(n11317) );
  NOR2_X1 U13859 ( .A1(n11305), .A2(n15028), .ZN(n15027) );
  NOR3_X1 U13860 ( .A1(n15027), .A2(n11767), .A3(n11336), .ZN(n11335) );
  NOR2_X1 U13861 ( .A1(n11335), .A2(n11306), .ZN(n11307) );
  XNOR2_X1 U13862 ( .A(n11307), .B(n11763), .ZN(n11309) );
  AOI22_X1 U13863 ( .A1(n15069), .A2(n15029), .B1(n12357), .B2(n15066), .ZN(
        n11308) );
  OAI21_X1 U13864 ( .B1(n11309), .B2(n15043), .A(n11308), .ZN(n11310) );
  AOI21_X1 U13865 ( .B1(n15119), .B2(n15031), .A(n11310), .ZN(n15116) );
  MUX2_X1 U13866 ( .A(n11311), .B(n15116), .S(n15091), .Z(n11316) );
  NOR2_X1 U13867 ( .A1(n11312), .A2(n15111), .ZN(n15118) );
  INV_X1 U13868 ( .A(n11313), .ZN(n11314) );
  AOI22_X1 U13869 ( .A1(n15058), .A2(n15118), .B1(n15053), .B2(n11314), .ZN(
        n11315) );
  OAI211_X1 U13870 ( .C1(n11318), .C2(n11317), .A(n11316), .B(n11315), .ZN(
        P3_U3226) );
  OAI21_X1 U13871 ( .B1(n14176), .B2(n11320), .A(n11319), .ZN(n11516) );
  XNOR2_X1 U13872 ( .A(n11516), .B(n11327), .ZN(n11514) );
  XNOR2_X1 U13873 ( .A(n11514), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n11331) );
  AOI21_X1 U13874 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n11322), .A(n11321), 
        .ZN(n11323) );
  NOR2_X1 U13875 ( .A1(n11323), .A2(n11327), .ZN(n11512) );
  AOI21_X1 U13876 ( .B1(n11323), .B2(n11327), .A(n11512), .ZN(n11325) );
  AND2_X1 U13877 ( .A1(n11325), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n11511) );
  INV_X1 U13878 ( .A(n11511), .ZN(n11324) );
  OAI211_X1 U13879 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11325), .A(n11324), 
        .B(n14607), .ZN(n11330) );
  NAND2_X1 U13880 ( .A1(n14594), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n11326) );
  NAND2_X1 U13881 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13831)
         );
  OAI211_X1 U13882 ( .C1(n14602), .C2(n11327), .A(n11326), .B(n13831), .ZN(
        n11328) );
  INV_X1 U13883 ( .A(n11328), .ZN(n11329) );
  OAI211_X1 U13884 ( .C1(n11331), .C2(n14604), .A(n11330), .B(n11329), .ZN(
        P1_U3261) );
  XNOR2_X1 U13885 ( .A(n11333), .B(n11332), .ZN(n11341) );
  INV_X1 U13886 ( .A(n11341), .ZN(n15115) );
  OAI22_X1 U13887 ( .A1(n12691), .A2(n15112), .B1(n11334), .B2(n15083), .ZN(
        n11343) );
  INV_X1 U13888 ( .A(n15031), .ZN(n15076) );
  INV_X1 U13889 ( .A(n11335), .ZN(n11338) );
  OAI21_X1 U13890 ( .B1(n15027), .B2(n11336), .A(n11767), .ZN(n11337) );
  NAND3_X1 U13891 ( .A1(n11338), .A2(n15072), .A3(n11337), .ZN(n11340) );
  AOI22_X1 U13892 ( .A1(n15069), .A2(n12359), .B1(n12358), .B2(n15066), .ZN(
        n11339) );
  OAI211_X1 U13893 ( .C1(n15076), .C2(n11341), .A(n11340), .B(n11339), .ZN(
        n15113) );
  MUX2_X1 U13894 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n15113), .S(n15091), .Z(
        n11342) );
  AOI211_X1 U13895 ( .C1(n15115), .C2(n12544), .A(n11343), .B(n11342), .ZN(
        n11344) );
  INV_X1 U13896 ( .A(n11344), .ZN(P3_U3227) );
  XNOR2_X1 U13897 ( .A(n11882), .B(n11552), .ZN(n12003) );
  XOR2_X1 U13898 ( .A(n11345), .B(n12003), .Z(n11346) );
  OAI222_X1 U13899 ( .A1(n14617), .A2(n11496), .B1(n11346), .B2(n14639), .C1(
        n14127), .C2(n6791), .ZN(n14555) );
  INV_X1 U13900 ( .A(n14555), .ZN(n11353) );
  XNOR2_X1 U13901 ( .A(n11347), .B(n12003), .ZN(n14557) );
  OAI211_X1 U13902 ( .C1(n6574), .C2(n14554), .A(n14725), .B(n14412), .ZN(
        n14553) );
  NAND2_X1 U13903 ( .A1(n14625), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11348) );
  OAI21_X1 U13904 ( .B1(n14229), .B2(n14536), .A(n11348), .ZN(n11349) );
  AOI21_X1 U13905 ( .B1(n11882), .B2(n14646), .A(n11349), .ZN(n11350) );
  OAI21_X1 U13906 ( .B1(n14553), .B2(n14216), .A(n11350), .ZN(n11351) );
  AOI21_X1 U13907 ( .B1(n14557), .B2(n14634), .A(n11351), .ZN(n11352) );
  OAI21_X1 U13908 ( .B1(n11353), .B2(n14656), .A(n11352), .ZN(P1_U3282) );
  AND2_X1 U13909 ( .A1(n14525), .A2(n13704), .ZN(n11357) );
  XNOR2_X1 U13910 ( .A(n11358), .B(n13750), .ZN(n11547) );
  XOR2_X1 U13911 ( .A(n11546), .B(n11547), .Z(n11550) );
  XNOR2_X1 U13912 ( .A(n11551), .B(n11550), .ZN(n11365) );
  INV_X1 U13913 ( .A(n14528), .ZN(n14510) );
  NOR2_X1 U13914 ( .A1(n14510), .A2(n11552), .ZN(n11359) );
  AOI211_X1 U13915 ( .C1(n14526), .C2(n13866), .A(n11360), .B(n11359), .ZN(
        n11361) );
  OAI21_X1 U13916 ( .B1(n15303), .B2(n11362), .A(n11361), .ZN(n11363) );
  AOI21_X1 U13917 ( .B1(n15311), .B2(n14741), .A(n11363), .ZN(n11364) );
  OAI21_X1 U13918 ( .B1(n11365), .B2(n15306), .A(n11364), .ZN(P1_U3217) );
  XNOR2_X1 U13919 ( .A(n11366), .B(n11674), .ZN(n15133) );
  XNOR2_X1 U13920 ( .A(n11367), .B(n11674), .ZN(n11369) );
  AOI22_X1 U13921 ( .A1(n12688), .A2(n15066), .B1(n15069), .B2(n12356), .ZN(
        n11368) );
  OAI21_X1 U13922 ( .B1(n11369), .B2(n15043), .A(n11368), .ZN(n11370) );
  AOI21_X1 U13923 ( .B1(n15133), .B2(n15031), .A(n11370), .ZN(n15135) );
  NOR2_X1 U13924 ( .A1(n12129), .A2(n15111), .ZN(n15131) );
  INV_X1 U13925 ( .A(n12196), .ZN(n11371) );
  AOI22_X1 U13926 ( .A1(n15058), .A2(n15131), .B1(n15053), .B2(n11371), .ZN(
        n11372) );
  OAI21_X1 U13927 ( .B1(n11080), .B2(n15091), .A(n11372), .ZN(n11373) );
  AOI21_X1 U13928 ( .B1(n15133), .B2(n12544), .A(n11373), .ZN(n11374) );
  OAI21_X1 U13929 ( .B1(n15135), .B2(n15093), .A(n11374), .ZN(P3_U3223) );
  INV_X1 U13930 ( .A(n11378), .ZN(n11375) );
  NAND2_X1 U13931 ( .A1(n11380), .A2(n13107), .ZN(n11377) );
  XNOR2_X1 U13932 ( .A(n11452), .B(n11451), .ZN(n13551) );
  NAND2_X1 U13933 ( .A1(n11379), .A2(n11378), .ZN(n11382) );
  OR2_X1 U13934 ( .A1(n11380), .A2(n11397), .ZN(n11381) );
  INV_X1 U13935 ( .A(n11457), .ZN(n11383) );
  AOI21_X1 U13936 ( .B1(n11451), .B2(n11384), .A(n11383), .ZN(n11385) );
  OAI222_X1 U13937 ( .A1(n14885), .A2(n12059), .B1(n13422), .B2(n11397), .C1(
        n11385), .C2(n13424), .ZN(n13547) );
  NAND2_X1 U13938 ( .A1(n13547), .A2(n13402), .ZN(n11392) );
  AOI211_X1 U13939 ( .C1(n13549), .C2(n11386), .A(n9733), .B(n11465), .ZN(
        n13548) );
  INV_X1 U13940 ( .A(n13549), .ZN(n11387) );
  NOR2_X1 U13941 ( .A1(n11387), .A2(n14874), .ZN(n11390) );
  OAI22_X1 U13942 ( .A1(n13402), .A2(n11388), .B1(n11395), .B2(n14881), .ZN(
        n11389) );
  AOI211_X1 U13943 ( .C1(n13548), .C2(n14850), .A(n11390), .B(n11389), .ZN(
        n11391) );
  OAI211_X1 U13944 ( .C1(n13551), .C2(n14871), .A(n11392), .B(n11391), .ZN(
        P2_U3254) );
  AOI22_X1 U13945 ( .A1(n13078), .A2(n13107), .B1(n13046), .B2(n13445), .ZN(
        n11394) );
  OAI211_X1 U13946 ( .C1(n11395), .C2(n13091), .A(n11394), .B(n11393), .ZN(
        n11404) );
  INV_X1 U13947 ( .A(n11396), .ZN(n11400) );
  NOR3_X1 U13948 ( .A1(n11398), .A2(n11397), .A3(n13075), .ZN(n11399) );
  AOI21_X1 U13949 ( .B1(n11400), .B2(n13085), .A(n11399), .ZN(n11402) );
  NOR2_X1 U13950 ( .A1(n11402), .A2(n11401), .ZN(n11403) );
  AOI211_X1 U13951 ( .C1(n13549), .C2(n13093), .A(n11404), .B(n11403), .ZN(
        n11405) );
  OAI21_X1 U13952 ( .B1(n11422), .B2(n13082), .A(n11405), .ZN(P2_U3208) );
  INV_X1 U13953 ( .A(n11406), .ZN(n11407) );
  NAND2_X1 U13954 ( .A1(n11407), .A2(n12358), .ZN(n11408) );
  XNOR2_X1 U13955 ( .A(n11410), .B(n12159), .ZN(n11530) );
  XNOR2_X1 U13956 ( .A(n11530), .B(n12357), .ZN(n11411) );
  OAI211_X1 U13957 ( .C1(n11412), .C2(n11411), .A(n11533), .B(n12337), .ZN(
        n11418) );
  INV_X1 U13958 ( .A(n12356), .ZN(n12191) );
  OAI22_X1 U13959 ( .A1(n11413), .A2(n12340), .B1(n12191), .B2(n12327), .ZN(
        n11414) );
  AOI211_X1 U13960 ( .C1(n11416), .C2(n12330), .A(n11415), .B(n11414), .ZN(
        n11417) );
  OAI211_X1 U13961 ( .C1(n11419), .C2(n12339), .A(n11418), .B(n11417), .ZN(
        P3_U3161) );
  AOI22_X1 U13962 ( .A1(n13078), .A2(n13106), .B1(n13046), .B2(n13105), .ZN(
        n11421) );
  OAI211_X1 U13963 ( .C1(n11463), .C2(n13091), .A(n11421), .B(n11420), .ZN(
        n11428) );
  INV_X1 U13964 ( .A(n11422), .ZN(n11426) );
  INV_X1 U13965 ( .A(n13075), .ZN(n13084) );
  AOI22_X1 U13966 ( .A1(n11423), .A2(n13085), .B1(n13084), .B2(n13106), .ZN(
        n11425) );
  NOR3_X1 U13967 ( .A1(n11426), .A2(n11425), .A3(n11424), .ZN(n11427) );
  AOI211_X1 U13968 ( .C1(n12092), .C2(n13093), .A(n11428), .B(n11427), .ZN(
        n11429) );
  OAI21_X1 U13969 ( .B1(n11430), .B2(n13082), .A(n11429), .ZN(P2_U3196) );
  AOI21_X1 U13970 ( .B1(n11434), .B2(P2_REG1_REG_16__SCAN_IN), .A(n11431), 
        .ZN(n11433) );
  XNOR2_X1 U13971 ( .A(n13166), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11432) );
  NOR2_X1 U13972 ( .A1(n11433), .A2(n11432), .ZN(n13165) );
  AOI211_X1 U13973 ( .C1(n11433), .C2(n11432), .A(n14844), .B(n13165), .ZN(
        n11446) );
  INV_X1 U13974 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n11444) );
  AND2_X1 U13975 ( .A1(n11434), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11438) );
  AOI21_X1 U13976 ( .B1(n13159), .B2(P2_REG2_REG_17__SCAN_IN), .A(n11438), 
        .ZN(n11435) );
  OAI21_X1 U13977 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n13159), .A(n11435), 
        .ZN(n11439) );
  NAND2_X1 U13978 ( .A1(n13166), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11437) );
  INV_X1 U13979 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13160) );
  NAND2_X1 U13980 ( .A1(n13159), .A2(n13160), .ZN(n11436) );
  OAI211_X1 U13981 ( .C1(n11440), .C2(n11438), .A(n11437), .B(n11436), .ZN(
        n13158) );
  OAI211_X1 U13982 ( .C1(n11440), .C2(n11439), .A(n13158), .B(n14838), .ZN(
        n11443) );
  AND2_X1 U13983 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11441) );
  AOI21_X1 U13984 ( .B1(n14840), .B2(n13166), .A(n11441), .ZN(n11442) );
  OAI211_X1 U13985 ( .C1(n14848), .C2(n11444), .A(n11443), .B(n11442), .ZN(
        n11445) );
  OR2_X1 U13986 ( .A1(n11446), .A2(n11445), .ZN(P2_U3231) );
  INV_X1 U13987 ( .A(n11447), .ZN(n11448) );
  OAI222_X1 U13988 ( .A1(P3_U3151), .A2(n11450), .B1(n14376), .B2(n11449), 
        .C1(n14378), .C2(n11448), .ZN(P3_U3269) );
  NAND2_X1 U13989 ( .A1(n11452), .A2(n11451), .ZN(n11454) );
  NAND2_X1 U13990 ( .A1(n13549), .A2(n13106), .ZN(n11453) );
  XNOR2_X1 U13991 ( .A(n12094), .B(n11458), .ZN(n14498) );
  NAND2_X1 U13992 ( .A1(n13549), .A2(n11455), .ZN(n11456) );
  INV_X1 U13993 ( .A(n11458), .ZN(n11459) );
  OAI211_X1 U13994 ( .C1(n11460), .C2(n11459), .A(n14882), .B(n12061), .ZN(
        n11462) );
  AOI22_X1 U13995 ( .A1(n13444), .A2(n13106), .B1(n13105), .B2(n13441), .ZN(
        n11461) );
  OAI211_X1 U13996 ( .C1(n14498), .C2(n14922), .A(n11462), .B(n11461), .ZN(
        n14501) );
  NAND2_X1 U13997 ( .A1(n14501), .A2(n13402), .ZN(n11469) );
  OAI22_X1 U13998 ( .A1(n13402), .A2(n11464), .B1(n11463), .B2(n14881), .ZN(
        n11467) );
  INV_X1 U13999 ( .A(n12092), .ZN(n14500) );
  OAI211_X1 U14000 ( .C1(n11465), .C2(n14500), .A(n13215), .B(n13447), .ZN(
        n14499) );
  NOR2_X1 U14001 ( .A1(n14499), .A2(n14868), .ZN(n11466) );
  AOI211_X1 U14002 ( .C1(n13433), .C2(n12092), .A(n11467), .B(n11466), .ZN(
        n11468) );
  OAI211_X1 U14003 ( .C1(n14498), .C2(n11470), .A(n11469), .B(n11468), .ZN(
        P2_U3253) );
  INV_X1 U14004 ( .A(n14382), .ZN(n12365) );
  NAND2_X1 U14005 ( .A1(n11478), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n11471) );
  AOI21_X1 U14006 ( .B1(n7882), .B2(n11473), .A(n12361), .ZN(n11489) );
  AOI21_X1 U14007 ( .B1(n11475), .B2(n11478), .A(n11474), .ZN(n11477) );
  MUX2_X1 U14008 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n11248), .Z(n12364) );
  XNOR2_X1 U14009 ( .A(n12364), .B(n12365), .ZN(n11476) );
  NAND2_X1 U14010 ( .A1(n11477), .A2(n11476), .ZN(n12372) );
  OAI21_X1 U14011 ( .B1(n11477), .B2(n11476), .A(n12372), .ZN(n11487) );
  INV_X1 U14012 ( .A(n11478), .ZN(n11480) );
  OAI21_X1 U14013 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11481), .A(n12376), 
        .ZN(n11482) );
  NAND2_X1 U14014 ( .A1(n11482), .A2(n15007), .ZN(n11485) );
  NOR2_X1 U14015 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11483), .ZN(n12287) );
  AOI21_X1 U14016 ( .B1(n14995), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12287), 
        .ZN(n11484) );
  OAI211_X1 U14017 ( .C1(n14989), .C2(n14382), .A(n11485), .B(n11484), .ZN(
        n11486) );
  AOI21_X1 U14018 ( .B1(n11487), .B2(n15015), .A(n11486), .ZN(n11488) );
  OAI21_X1 U14019 ( .B1(n11489), .B2(n15001), .A(n11488), .ZN(P3_U3195) );
  INV_X1 U14020 ( .A(n11490), .ZN(n11492) );
  OAI222_X1 U14021 ( .A1(n14378), .A2(n11492), .B1(n14376), .B2(n11491), .C1(
        P3_U3151), .C2(n11248), .ZN(P3_U3268) );
  OAI222_X1 U14022 ( .A1(n13588), .A2(n11494), .B1(P2_U3088), .B2(n9693), .C1(
        n13590), .C2(n11493), .ZN(P2_U3305) );
  XNOR2_X1 U14023 ( .A(n11495), .B(n12002), .ZN(n11497) );
  OAI22_X1 U14024 ( .A1(n11496), .A2(n14127), .B1(n13850), .B2(n14617), .ZN(
        n11578) );
  AOI21_X1 U14025 ( .B1(n11497), .B2(n14403), .A(n11578), .ZN(n14549) );
  XNOR2_X1 U14026 ( .A(n11498), .B(n12002), .ZN(n14552) );
  INV_X1 U14027 ( .A(n11897), .ZN(n14550) );
  INV_X1 U14028 ( .A(n14413), .ZN(n11499) );
  OAI211_X1 U14029 ( .C1(n14550), .C2(n11499), .A(n14725), .B(n14225), .ZN(
        n14548) );
  OAI22_X1 U14030 ( .A1(n14231), .A2(n11500), .B1(n11581), .B2(n14229), .ZN(
        n11501) );
  AOI21_X1 U14031 ( .B1(n11897), .B2(n14646), .A(n11501), .ZN(n11502) );
  OAI21_X1 U14032 ( .B1(n14548), .B2(n14216), .A(n11502), .ZN(n11503) );
  AOI21_X1 U14033 ( .B1(n14552), .B2(n14634), .A(n11503), .ZN(n11504) );
  OAI21_X1 U14034 ( .B1(n14625), .B2(n14549), .A(n11504), .ZN(P1_U3280) );
  NAND2_X1 U14035 ( .A1(n11507), .A2(n14341), .ZN(n11505) );
  OAI211_X1 U14036 ( .C1(n11506), .C2(n14353), .A(n11505), .B(n12043), .ZN(
        P1_U3332) );
  NAND2_X1 U14037 ( .A1(n11507), .A2(n13577), .ZN(n11509) );
  OAI211_X1 U14038 ( .C1(n11510), .C2(n13588), .A(n11509), .B(n11508), .ZN(
        P2_U3304) );
  NOR2_X1 U14039 ( .A1(n11512), .A2(n11511), .ZN(n11513) );
  XNOR2_X1 U14040 ( .A(n11513), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14041 ( .A1(n11514), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U14042 ( .A1(n11516), .A2(n11515), .ZN(n11517) );
  NAND2_X1 U14043 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  XOR2_X1 U14044 ( .A(n11519), .B(P1_REG2_REG_19__SCAN_IN), .Z(n11523) );
  INV_X1 U14045 ( .A(n11523), .ZN(n11520) );
  NAND2_X1 U14046 ( .A1(n11520), .A2(n13976), .ZN(n11521) );
  OAI211_X1 U14047 ( .C1(n11524), .C2(n13926), .A(n11521), .B(n14602), .ZN(
        n11522) );
  INV_X1 U14048 ( .A(n11522), .ZN(n11527) );
  AOI22_X1 U14049 ( .A1(n11524), .A2(n14607), .B1(n11523), .B2(n13976), .ZN(
        n11526) );
  MUX2_X1 U14050 ( .A(n11527), .B(n11526), .S(n11525), .Z(n11528) );
  NAND2_X1 U14051 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13742)
         );
  OAI211_X1 U14052 ( .C1(n7687), .C2(n14611), .A(n11528), .B(n13742), .ZN(
        P1_U3262) );
  XNOR2_X1 U14053 ( .A(n11529), .B(n10597), .ZN(n12126) );
  XNOR2_X1 U14054 ( .A(n12126), .B(n12356), .ZN(n11536) );
  INV_X1 U14055 ( .A(n11530), .ZN(n11531) );
  NAND2_X1 U14056 ( .A1(n11531), .A2(n12357), .ZN(n11532) );
  INV_X1 U14057 ( .A(n12128), .ZN(n11534) );
  AOI21_X1 U14058 ( .B1(n11536), .B2(n11535), .A(n11534), .ZN(n11545) );
  NOR2_X1 U14059 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11537), .ZN(n14994) );
  INV_X1 U14060 ( .A(n14467), .ZN(n11538) );
  OAI22_X1 U14061 ( .A1(n11539), .A2(n12340), .B1(n11538), .B2(n12327), .ZN(
        n11540) );
  AOI211_X1 U14062 ( .C1(n11541), .C2(n12330), .A(n14994), .B(n11540), .ZN(
        n11544) );
  NAND2_X1 U14063 ( .A1(n12324), .A2(n11542), .ZN(n11543) );
  OAI211_X1 U14064 ( .C1(n11545), .C2(n12332), .A(n11544), .B(n11543), .ZN(
        P3_U3171) );
  INV_X1 U14065 ( .A(n11546), .ZN(n11549) );
  INV_X1 U14066 ( .A(n11547), .ZN(n11548) );
  OAI22_X1 U14067 ( .A1(n14554), .A2(n13752), .B1(n11552), .B2(n13749), .ZN(
        n11557) );
  NAND2_X1 U14068 ( .A1(n11882), .A2(n13699), .ZN(n11554) );
  NAND2_X1 U14069 ( .A1(n14406), .A2(n13608), .ZN(n11553) );
  NAND2_X1 U14070 ( .A1(n11554), .A2(n11553), .ZN(n11555) );
  XNOR2_X1 U14071 ( .A(n11555), .B(n13750), .ZN(n11556) );
  XOR2_X1 U14072 ( .A(n11557), .B(n11556), .Z(n14524) );
  INV_X1 U14073 ( .A(n11556), .ZN(n11559) );
  INV_X1 U14074 ( .A(n11557), .ZN(n11558) );
  NAND2_X1 U14075 ( .A1(n11559), .A2(n11558), .ZN(n11564) );
  AND2_X1 U14076 ( .A1(n14522), .A2(n11564), .ZN(n11566) );
  NAND2_X1 U14077 ( .A1(n14410), .A2(n13699), .ZN(n11561) );
  NAND2_X1 U14078 ( .A1(n14527), .A2(n13700), .ZN(n11560) );
  NAND2_X1 U14079 ( .A1(n11561), .A2(n11560), .ZN(n11562) );
  XNOR2_X1 U14080 ( .A(n11562), .B(n10692), .ZN(n11573) );
  AND2_X1 U14081 ( .A1(n14527), .A2(n13704), .ZN(n11563) );
  XNOR2_X1 U14082 ( .A(n11573), .B(n11575), .ZN(n11565) );
  OAI211_X1 U14083 ( .C1(n11566), .C2(n11565), .A(n14532), .B(n11574), .ZN(
        n11572) );
  NOR2_X1 U14084 ( .A1(n15303), .A2(n14408), .ZN(n11570) );
  OAI22_X1 U14085 ( .A1(n14510), .A2(n11568), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11567), .ZN(n11569) );
  AOI211_X1 U14086 ( .C1(n14526), .C2(n14406), .A(n11570), .B(n11569), .ZN(
        n11571) );
  OAI211_X1 U14087 ( .C1(n7185), .C2(n14530), .A(n11572), .B(n11571), .ZN(
        P1_U3224) );
  AND2_X1 U14088 ( .A1(n14405), .A2(n13704), .ZN(n11576) );
  AOI22_X1 U14089 ( .A1(n11897), .A2(n13699), .B1(n13608), .B2(n14405), .ZN(
        n11577) );
  XNOR2_X1 U14090 ( .A(n11577), .B(n13750), .ZN(n13603) );
  XOR2_X1 U14091 ( .A(n13602), .B(n13603), .Z(n13606) );
  XNOR2_X1 U14092 ( .A(n13607), .B(n13606), .ZN(n11584) );
  NAND2_X1 U14093 ( .A1(n11578), .A2(n15299), .ZN(n11580) );
  OAI211_X1 U14094 ( .C1(n15303), .C2(n11581), .A(n11580), .B(n11579), .ZN(
        n11582) );
  AOI21_X1 U14095 ( .B1(n11897), .B2(n15311), .A(n11582), .ZN(n11583) );
  OAI21_X1 U14096 ( .B1(n11584), .B2(n15306), .A(n11583), .ZN(P1_U3234) );
  INV_X1 U14097 ( .A(n11806), .ZN(n12125) );
  OAI222_X1 U14098 ( .A1(n13588), .A2(n11588), .B1(n13590), .B2(n11587), .C1(
        n11586), .C2(P2_U3088), .ZN(P2_U3307) );
  INV_X1 U14099 ( .A(n11589), .ZN(n13580) );
  OAI222_X1 U14100 ( .A1(n14353), .A2(n11590), .B1(n11585), .B2(n13580), .C1(
        P1_U3086), .C2(n6440), .ZN(P1_U3328) );
  INV_X1 U14101 ( .A(n11591), .ZN(n11799) );
  OAI222_X1 U14102 ( .A1(n11585), .A2(n11799), .B1(n11592), .B2(P1_U3086), 
        .C1(n11597), .C2(n14353), .ZN(P1_U3326) );
  INV_X1 U14103 ( .A(n11781), .ZN(n11753) );
  INV_X1 U14104 ( .A(n11594), .ZN(n11595) );
  NAND2_X1 U14105 ( .A1(n11596), .A2(n11595), .ZN(n11599) );
  NAND2_X1 U14106 ( .A1(n11597), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11598) );
  XNOR2_X1 U14107 ( .A(n12124), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11600) );
  XNOR2_X1 U14108 ( .A(n11613), .B(n11600), .ZN(n12857) );
  NAND2_X1 U14109 ( .A1(n12857), .A2(n11616), .ZN(n11602) );
  OR2_X1 U14110 ( .A1(n6441), .A2(n12859), .ZN(n11601) );
  INV_X1 U14111 ( .A(n14478), .ZN(n11623) );
  INV_X1 U14112 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n11607) );
  NAND2_X1 U14113 ( .A1(n11603), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n11606) );
  INV_X1 U14114 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12466) );
  OR2_X1 U14115 ( .A1(n11604), .A2(n12466), .ZN(n11605) );
  OAI211_X1 U14116 ( .C1(n11608), .C2(n11607), .A(n11606), .B(n11605), .ZN(
        n11609) );
  INV_X1 U14117 ( .A(n11609), .ZN(n11610) );
  AND2_X1 U14118 ( .A1(n11807), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n11612) );
  XNOR2_X1 U14119 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11614) );
  XNOR2_X1 U14120 ( .A(n11615), .B(n11614), .ZN(n12855) );
  NAND2_X1 U14121 ( .A1(n12855), .A2(n11616), .ZN(n11618) );
  OR2_X1 U14122 ( .A1(n6441), .A2(n12852), .ZN(n11617) );
  NAND2_X1 U14123 ( .A1(n11618), .A2(n11617), .ZN(n12461) );
  INV_X1 U14124 ( .A(n12348), .ZN(n11619) );
  NAND2_X1 U14125 ( .A1(n14478), .A2(n11619), .ZN(n11621) );
  AND2_X1 U14126 ( .A1(n11621), .A2(n11620), .ZN(n11622) );
  OAI21_X1 U14127 ( .B1(n11623), .B2(n12463), .A(n11784), .ZN(n11625) );
  INV_X1 U14128 ( .A(n12461), .ZN(n12785) );
  OAI22_X1 U14129 ( .A1(n11626), .A2(n11625), .B1(n12785), .B2(n11783), .ZN(
        n11627) );
  INV_X1 U14130 ( .A(n11628), .ZN(n11791) );
  MUX2_X1 U14131 ( .A(n11739), .B(n11740), .S(n11754), .Z(n11746) );
  XNOR2_X1 U14132 ( .A(n11629), .B(n11754), .ZN(n11736) );
  NAND2_X1 U14133 ( .A1(n11644), .A2(n11630), .ZN(n11635) );
  MUX2_X1 U14134 ( .A(n11632), .B(n11642), .S(n11748), .Z(n11631) );
  NAND2_X1 U14135 ( .A1(n11762), .A2(n11631), .ZN(n11641) );
  AND3_X1 U14136 ( .A1(n11632), .A2(n11637), .A3(n11793), .ZN(n11636) );
  OAI211_X1 U14137 ( .C1(n11641), .C2(n11636), .A(n11633), .B(n11645), .ZN(
        n11634) );
  MUX2_X1 U14138 ( .A(n11635), .B(n11634), .S(n11748), .Z(n11648) );
  INV_X1 U14139 ( .A(n11636), .ZN(n11638) );
  NAND2_X1 U14140 ( .A1(n11638), .A2(n11637), .ZN(n11640) );
  MUX2_X1 U14141 ( .A(n12777), .B(n11640), .S(n11639), .Z(n11643) );
  AOI21_X1 U14142 ( .B1(n11643), .B2(n11642), .A(n11641), .ZN(n11647) );
  MUX2_X1 U14143 ( .A(n11645), .B(n11644), .S(n11748), .Z(n11646) );
  OAI211_X1 U14144 ( .C1(n11648), .C2(n11647), .A(n11759), .B(n11646), .ZN(
        n11652) );
  MUX2_X1 U14145 ( .A(n11650), .B(n11649), .S(n11748), .Z(n11651) );
  AND3_X1 U14146 ( .A1(n11652), .A2(n15028), .A3(n11651), .ZN(n11656) );
  AOI21_X1 U14147 ( .B1(n11661), .B2(n11653), .A(n11754), .ZN(n11662) );
  AOI21_X1 U14148 ( .B1(n11657), .B2(n11654), .A(n11748), .ZN(n11655) );
  NOR3_X1 U14149 ( .A1(n11656), .A2(n11662), .A3(n11655), .ZN(n11667) );
  INV_X1 U14150 ( .A(n11657), .ZN(n11659) );
  AOI21_X1 U14151 ( .B1(n11659), .B2(n11748), .A(n11658), .ZN(n11660) );
  OAI21_X1 U14152 ( .B1(n11662), .B2(n11661), .A(n11660), .ZN(n11666) );
  MUX2_X1 U14153 ( .A(n11664), .B(n11663), .S(n11748), .Z(n11665) );
  OAI211_X1 U14154 ( .C1(n11667), .C2(n11666), .A(n11761), .B(n11665), .ZN(
        n11671) );
  MUX2_X1 U14155 ( .A(n11669), .B(n11668), .S(n11754), .Z(n11670) );
  NAND3_X1 U14156 ( .A1(n11671), .A2(n11760), .A3(n11670), .ZN(n11676) );
  MUX2_X1 U14157 ( .A(n11673), .B(n11672), .S(n11748), .Z(n11675) );
  AOI21_X1 U14158 ( .B1(n11676), .B2(n11675), .A(n11674), .ZN(n11682) );
  INV_X1 U14159 ( .A(n11677), .ZN(n11680) );
  INV_X1 U14160 ( .A(n11678), .ZN(n11679) );
  MUX2_X1 U14161 ( .A(n11680), .B(n11679), .S(n11754), .Z(n11681) );
  NOR3_X1 U14162 ( .A1(n11682), .A2(n11681), .A3(n14471), .ZN(n11691) );
  NAND2_X1 U14163 ( .A1(n11688), .A2(n11683), .ZN(n11686) );
  NAND2_X1 U14164 ( .A1(n11687), .A2(n11684), .ZN(n11685) );
  MUX2_X1 U14165 ( .A(n11686), .B(n11685), .S(n11754), .Z(n11690) );
  INV_X1 U14166 ( .A(n12671), .ZN(n12668) );
  MUX2_X1 U14167 ( .A(n11688), .B(n11687), .S(n11748), .Z(n11689) );
  OAI211_X1 U14168 ( .C1(n11691), .C2(n11690), .A(n12668), .B(n11689), .ZN(
        n11701) );
  INV_X1 U14169 ( .A(n11693), .ZN(n11694) );
  MUX2_X1 U14170 ( .A(n7004), .B(n11694), .S(n11754), .Z(n11695) );
  NOR3_X1 U14171 ( .A1(n12644), .A2(n11695), .A3(n12657), .ZN(n11700) );
  OAI211_X1 U14172 ( .C1(n12644), .C2(n11698), .A(n11697), .B(n11696), .ZN(
        n11699) );
  AOI22_X1 U14173 ( .A1(n11701), .A2(n11700), .B1(n11754), .B2(n11699), .ZN(
        n11708) );
  INV_X1 U14174 ( .A(n11702), .ZN(n11707) );
  INV_X1 U14175 ( .A(n11704), .ZN(n11705) );
  AOI211_X1 U14176 ( .C1(n12641), .C2(n7001), .A(n11705), .B(n11707), .ZN(
        n11706) );
  OAI22_X1 U14177 ( .A1(n11708), .A2(n11707), .B1(n11706), .B2(n11754), .ZN(
        n11710) );
  INV_X1 U14178 ( .A(n12831), .ZN(n12635) );
  NAND3_X1 U14179 ( .A1(n12635), .A2(n11748), .A3(n12646), .ZN(n11709) );
  AOI211_X1 U14180 ( .C1(n11710), .C2(n11709), .A(n12613), .B(n7296), .ZN(
        n11722) );
  INV_X1 U14181 ( .A(n11714), .ZN(n11713) );
  OAI211_X1 U14182 ( .C1(n11713), .C2(n11712), .A(n11718), .B(n11711), .ZN(
        n11717) );
  OAI211_X1 U14183 ( .C1(n7296), .C2(n11715), .A(n11719), .B(n11714), .ZN(
        n11716) );
  MUX2_X1 U14184 ( .A(n11717), .B(n11716), .S(n11754), .Z(n11721) );
  MUX2_X1 U14185 ( .A(n11719), .B(n11718), .S(n11754), .Z(n11720) );
  OAI211_X1 U14186 ( .C1(n11722), .C2(n11721), .A(n12581), .B(n11720), .ZN(
        n11726) );
  NAND2_X1 U14187 ( .A1(n12815), .A2(n12563), .ZN(n11724) );
  MUX2_X1 U14188 ( .A(n11724), .B(n11723), .S(n11748), .Z(n11725) );
  NAND3_X1 U14189 ( .A1(n11726), .A2(n12561), .A3(n11725), .ZN(n11730) );
  MUX2_X1 U14190 ( .A(n11728), .B(n11727), .S(n11754), .Z(n11729) );
  NAND3_X1 U14191 ( .A1(n11730), .A2(n12551), .A3(n11729), .ZN(n11734) );
  MUX2_X1 U14192 ( .A(n11732), .B(n11731), .S(n11748), .Z(n11733) );
  AND3_X1 U14193 ( .A1(n11734), .A2(n11775), .A3(n11733), .ZN(n11735) );
  MUX2_X1 U14194 ( .A(n11736), .B(n11735), .S(n11777), .Z(n11738) );
  NOR3_X1 U14195 ( .A1(n12521), .A2(n11775), .A3(n11754), .ZN(n11737) );
  NOR3_X1 U14196 ( .A1(n11738), .A2(n12503), .A3(n11737), .ZN(n11741) );
  NAND2_X1 U14197 ( .A1(n12476), .A2(n12491), .ZN(n11779) );
  OAI22_X1 U14198 ( .A1(n11741), .A2(n11779), .B1(n11748), .B2(n11742), .ZN(
        n11744) );
  NAND4_X1 U14199 ( .A1(n11742), .A2(n12519), .A3(n12511), .A4(n11754), .ZN(
        n11743) );
  NAND3_X1 U14200 ( .A1(n11749), .A2(n11748), .A3(n11747), .ZN(n11750) );
  NAND4_X1 U14201 ( .A1(n11761), .A2(n11760), .A3(n15028), .A4(n11759), .ZN(
        n11766) );
  NAND3_X1 U14202 ( .A1(n11764), .A2(n11763), .A3(n11762), .ZN(n11765) );
  NOR2_X1 U14203 ( .A1(n11766), .A2(n11765), .ZN(n11771) );
  INV_X1 U14204 ( .A(n14471), .ZN(n14466) );
  INV_X1 U14205 ( .A(n10546), .ZN(n11768) );
  AND4_X1 U14206 ( .A1(n15055), .A2(n11769), .A3(n11768), .A4(n11767), .ZN(
        n11770) );
  NAND4_X1 U14207 ( .A1(n11771), .A2(n14466), .A3(n12683), .A4(n11770), .ZN(
        n11772) );
  NOR4_X1 U14208 ( .A1(n11772), .A2(n12644), .A3(n12657), .A4(n12671), .ZN(
        n11773) );
  NAND4_X1 U14209 ( .A1(n12601), .A2(n12610), .A3(n12631), .A4(n11773), .ZN(
        n11774) );
  NOR4_X1 U14210 ( .A1(n7307), .A2(n12572), .A3(n7644), .A4(n11774), .ZN(
        n11776) );
  NAND4_X1 U14211 ( .A1(n11777), .A2(n12551), .A3(n11776), .A4(n11775), .ZN(
        n11778) );
  NOR4_X1 U14212 ( .A1(n11780), .A2(n11779), .A3(n12503), .A4(n11778), .ZN(
        n11782) );
  NAND4_X1 U14213 ( .A1(n11784), .A2(n11783), .A3(n11782), .A4(n11781), .ZN(
        n11786) );
  XNOR2_X1 U14214 ( .A(n11786), .B(n11785), .ZN(n11789) );
  INV_X1 U14215 ( .A(n11787), .ZN(n11788) );
  NOR3_X1 U14216 ( .A1(n15048), .A2(n8191), .A3(n11792), .ZN(n11795) );
  OAI21_X1 U14217 ( .B1(n11796), .B2(n11793), .A(P3_B_REG_SCAN_IN), .ZN(n11794) );
  OAI22_X1 U14218 ( .A1(n11797), .A2(n11796), .B1(n11795), .B2(n11794), .ZN(
        P3_U3296) );
  OAI222_X1 U14219 ( .A1(P2_U3088), .A2(n8466), .B1(n13590), .B2(n11799), .C1(
        n11798), .C2(n13588), .ZN(P2_U3298) );
  INV_X1 U14220 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n11800) );
  OR2_X1 U14221 ( .A1(n9254), .A2(n11800), .ZN(n11805) );
  INV_X1 U14222 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n11801) );
  OR2_X1 U14223 ( .A1(n11802), .A2(n11801), .ZN(n11804) );
  AND3_X1 U14224 ( .A1(n11805), .A2(n11804), .A3(n11803), .ZN(n13982) );
  INV_X1 U14225 ( .A(n13982), .ZN(n13856) );
  OAI21_X1 U14226 ( .B1(n13856), .B2(n11981), .A(n13857), .ZN(n11812) );
  NAND2_X1 U14227 ( .A1(n11806), .A2(n11980), .ZN(n11809) );
  OR2_X1 U14228 ( .A1(n11978), .A2(n11807), .ZN(n11808) );
  INV_X1 U14229 ( .A(n14357), .ZN(n11982) );
  NAND2_X1 U14230 ( .A1(n11982), .A2(n14230), .ZN(n11810) );
  MUX2_X1 U14231 ( .A(n11812), .B(n14243), .S(n11903), .Z(n11977) );
  NAND2_X1 U14232 ( .A1(n13860), .A2(n11903), .ZN(n11813) );
  MUX2_X1 U14233 ( .A(n13862), .B(n14283), .S(n6435), .Z(n11938) );
  NAND3_X1 U14234 ( .A1(n14306), .A2(n7100), .A3(n11903), .ZN(n11816) );
  OAI21_X1 U14235 ( .B1(n11817), .B2(n11903), .A(n11816), .ZN(n11818) );
  INV_X1 U14236 ( .A(n11818), .ZN(n11928) );
  NAND2_X1 U14237 ( .A1(n11820), .A2(n11824), .ZN(n11821) );
  MUX2_X1 U14238 ( .A(n11822), .B(n11821), .S(n11903), .Z(n11831) );
  AND2_X1 U14239 ( .A1(n11823), .A2(n11988), .ZN(n11830) );
  INV_X1 U14240 ( .A(n11824), .ZN(n11827) );
  INV_X1 U14241 ( .A(n11825), .ZN(n11826) );
  INV_X1 U14242 ( .A(n11828), .ZN(n11829) );
  OAI21_X1 U14243 ( .B1(n11831), .B2(n11830), .A(n11829), .ZN(n11836) );
  MUX2_X1 U14244 ( .A(n13872), .B(n11832), .S(n11903), .Z(n11835) );
  MUX2_X1 U14245 ( .A(n14692), .B(n11833), .S(n11903), .Z(n11834) );
  OAI21_X1 U14246 ( .B1(n11836), .B2(n11835), .A(n11834), .ZN(n11838) );
  NAND2_X1 U14247 ( .A1(n11836), .A2(n11835), .ZN(n11837) );
  NAND2_X1 U14248 ( .A1(n6435), .A2(n11839), .ZN(n11842) );
  NAND2_X1 U14249 ( .A1(n11903), .A2(n11840), .ZN(n11841) );
  MUX2_X1 U14250 ( .A(n11842), .B(n11841), .S(n13871), .Z(n11843) );
  MUX2_X1 U14251 ( .A(n13870), .B(n14700), .S(n11903), .Z(n11844) );
  INV_X1 U14252 ( .A(n11844), .ZN(n11846) );
  MUX2_X1 U14253 ( .A(n13870), .B(n14700), .S(n6435), .Z(n11845) );
  MUX2_X1 U14254 ( .A(n14708), .B(n13869), .S(n11903), .Z(n11849) );
  NAND2_X1 U14255 ( .A1(n11850), .A2(n11849), .ZN(n11848) );
  MUX2_X1 U14256 ( .A(n14708), .B(n13869), .S(n6435), .Z(n11847) );
  NAND2_X1 U14257 ( .A1(n11848), .A2(n11847), .ZN(n11852) );
  MUX2_X1 U14258 ( .A(n14647), .B(n13868), .S(n6435), .Z(n11855) );
  NAND2_X1 U14259 ( .A1(n11856), .A2(n11855), .ZN(n11854) );
  MUX2_X1 U14260 ( .A(n14647), .B(n13868), .S(n11903), .Z(n11853) );
  NAND2_X1 U14261 ( .A1(n11854), .A2(n11853), .ZN(n11858) );
  MUX2_X1 U14262 ( .A(n14620), .B(n14724), .S(n6435), .Z(n11861) );
  NAND2_X1 U14263 ( .A1(n14620), .A2(n6435), .ZN(n11862) );
  NAND2_X1 U14264 ( .A1(n14724), .A2(n11903), .ZN(n11865) );
  NAND3_X1 U14265 ( .A1(n11861), .A2(n11862), .A3(n11865), .ZN(n11857) );
  MUX2_X1 U14266 ( .A(n13867), .B(n15310), .S(n11903), .Z(n11860) );
  NAND2_X1 U14267 ( .A1(n11860), .A2(n11859), .ZN(n11871) );
  INV_X1 U14268 ( .A(n11861), .ZN(n11867) );
  INV_X1 U14269 ( .A(n11862), .ZN(n11863) );
  NAND3_X1 U14270 ( .A1(n11867), .A2(n11864), .A3(n11863), .ZN(n11870) );
  INV_X1 U14271 ( .A(n11865), .ZN(n11866) );
  NAND3_X1 U14272 ( .A1(n11868), .A2(n11867), .A3(n11866), .ZN(n11869) );
  AND3_X1 U14273 ( .A1(n11871), .A2(n11870), .A3(n11869), .ZN(n11872) );
  MUX2_X1 U14274 ( .A(n14618), .B(n11873), .S(n6435), .Z(n11875) );
  MUX2_X1 U14275 ( .A(n13866), .B(n7189), .S(n11903), .Z(n11874) );
  MUX2_X1 U14276 ( .A(n14525), .B(n14741), .S(n11903), .Z(n11878) );
  NAND2_X1 U14277 ( .A1(n11879), .A2(n11878), .ZN(n11877) );
  MUX2_X1 U14278 ( .A(n14525), .B(n14741), .S(n6435), .Z(n11876) );
  NAND2_X1 U14279 ( .A1(n11877), .A2(n11876), .ZN(n11881) );
  MUX2_X1 U14280 ( .A(n14406), .B(n11882), .S(n6435), .Z(n11884) );
  MUX2_X1 U14281 ( .A(n14406), .B(n11882), .S(n11903), .Z(n11883) );
  MUX2_X1 U14282 ( .A(n14527), .B(n14410), .S(n11903), .Z(n11888) );
  NAND2_X1 U14283 ( .A1(n11887), .A2(n11888), .ZN(n11886) );
  MUX2_X1 U14284 ( .A(n14527), .B(n14410), .S(n6435), .Z(n11885) );
  NAND2_X1 U14285 ( .A1(n11886), .A2(n11885), .ZN(n11892) );
  INV_X1 U14286 ( .A(n11887), .ZN(n11890) );
  INV_X1 U14287 ( .A(n11888), .ZN(n11889) );
  NAND2_X1 U14288 ( .A1(n11890), .A2(n11889), .ZN(n11891) );
  MUX2_X1 U14289 ( .A(n14405), .B(n11897), .S(n6435), .Z(n11896) );
  OR2_X1 U14290 ( .A1(n14219), .A2(n11896), .ZN(n11895) );
  AND2_X1 U14291 ( .A1(n11904), .A2(n11893), .ZN(n11894) );
  AND2_X1 U14292 ( .A1(n11901), .A2(n11897), .ZN(n11898) );
  NAND2_X1 U14293 ( .A1(n11901), .A2(n11900), .ZN(n11902) );
  OR2_X1 U14294 ( .A1(n11904), .A2(n11903), .ZN(n11912) );
  MUX2_X1 U14295 ( .A(n14182), .B(n14518), .S(n6435), .Z(n11920) );
  NAND2_X1 U14296 ( .A1(n11920), .A2(n14195), .ZN(n11905) );
  NAND2_X1 U14297 ( .A1(n13851), .A2(n6435), .ZN(n11907) );
  AOI21_X1 U14298 ( .B1(n11905), .B2(n11907), .A(n14311), .ZN(n11911) );
  NAND2_X1 U14299 ( .A1(n11920), .A2(n14511), .ZN(n11906) );
  OR2_X1 U14300 ( .A1(n14518), .A2(n6435), .ZN(n11913) );
  AOI21_X1 U14301 ( .B1(n11906), .B2(n11913), .A(n7184), .ZN(n11910) );
  NAND2_X1 U14302 ( .A1(n14195), .A2(n11903), .ZN(n11914) );
  OR2_X1 U14303 ( .A1(n14518), .A2(n11914), .ZN(n11909) );
  INV_X1 U14304 ( .A(n11907), .ZN(n11917) );
  NAND2_X1 U14305 ( .A1(n11917), .A2(n14511), .ZN(n11908) );
  NAND2_X1 U14306 ( .A1(n11909), .A2(n11908), .ZN(n11919) );
  INV_X1 U14307 ( .A(n11913), .ZN(n11916) );
  INV_X1 U14308 ( .A(n11914), .ZN(n11915) );
  AOI21_X1 U14309 ( .B1(n11920), .B2(n11916), .A(n11915), .ZN(n11923) );
  NAND2_X1 U14310 ( .A1(n11920), .A2(n11917), .ZN(n11918) );
  OAI21_X1 U14311 ( .B1(n14195), .B2(n11903), .A(n11918), .ZN(n11921) );
  AOI22_X1 U14312 ( .A1(n11921), .A2(n7184), .B1(n11920), .B2(n11919), .ZN(
        n11922) );
  OAI211_X1 U14313 ( .C1(n11923), .C2(n7184), .A(n14160), .B(n11922), .ZN(
        n11924) );
  MUX2_X1 U14314 ( .A(n11926), .B(n11925), .S(n6435), .Z(n11927) );
  MUX2_X1 U14315 ( .A(n13649), .B(n13650), .S(n6435), .Z(n11930) );
  MUX2_X1 U14316 ( .A(n14144), .B(n14293), .S(n11903), .Z(n11929) );
  NAND2_X1 U14317 ( .A1(n11931), .A2(n11930), .ZN(n11932) );
  MUX2_X1 U14318 ( .A(n13863), .B(n14288), .S(n11903), .Z(n11935) );
  MUX2_X1 U14319 ( .A(n13863), .B(n14288), .S(n6435), .Z(n11934) );
  MUX2_X1 U14320 ( .A(n13862), .B(n14283), .S(n11903), .Z(n11936) );
  MUX2_X1 U14321 ( .A(n13861), .B(n14089), .S(n11903), .Z(n11941) );
  MUX2_X1 U14322 ( .A(n13861), .B(n14089), .S(n6435), .Z(n11939) );
  NAND2_X1 U14323 ( .A1(n11940), .A2(n11939), .ZN(n11944) );
  NAND2_X1 U14324 ( .A1(n11944), .A2(n11943), .ZN(n11946) );
  MUX2_X1 U14325 ( .A(n14274), .B(n13860), .S(n6435), .Z(n11945) );
  MUX2_X1 U14326 ( .A(n14029), .B(n14269), .S(n11903), .Z(n11950) );
  MUX2_X1 U14327 ( .A(n14029), .B(n14269), .S(n6435), .Z(n11948) );
  INV_X1 U14328 ( .A(n11950), .ZN(n11951) );
  MUX2_X1 U14329 ( .A(n13859), .B(n14264), .S(n6435), .Z(n11955) );
  NAND2_X1 U14330 ( .A1(n11954), .A2(n11955), .ZN(n11953) );
  MUX2_X1 U14331 ( .A(n14264), .B(n13859), .S(n6435), .Z(n11952) );
  NAND2_X1 U14332 ( .A1(n11953), .A2(n11952), .ZN(n11959) );
  INV_X1 U14333 ( .A(n11955), .ZN(n11956) );
  NAND2_X1 U14334 ( .A1(n11957), .A2(n11956), .ZN(n11958) );
  MUX2_X1 U14335 ( .A(n14030), .B(n14022), .S(n11903), .Z(n11961) );
  MUX2_X1 U14336 ( .A(n14030), .B(n14022), .S(n6435), .Z(n11960) );
  INV_X1 U14337 ( .A(n11961), .ZN(n11962) );
  MUX2_X1 U14338 ( .A(n13858), .B(n14252), .S(n6435), .Z(n11965) );
  MUX2_X1 U14339 ( .A(n13858), .B(n14252), .S(n11903), .Z(n11963) );
  MUX2_X1 U14340 ( .A(n14247), .B(n13996), .S(n6435), .Z(n11966) );
  MUX2_X1 U14341 ( .A(n13996), .B(n14247), .S(n6435), .Z(n11967) );
  INV_X1 U14342 ( .A(n11968), .ZN(n11969) );
  OAI22_X1 U14343 ( .A1(n13982), .A2(n6435), .B1(n6895), .B2(n11969), .ZN(
        n11971) );
  AOI22_X1 U14344 ( .A1(n13991), .A2(n6435), .B1(n13857), .B2(n11971), .ZN(
        n11973) );
  INV_X1 U14345 ( .A(n11972), .ZN(n11975) );
  INV_X1 U14346 ( .A(n11973), .ZN(n11974) );
  INV_X1 U14347 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14337) );
  NOR2_X1 U14348 ( .A1(n11978), .A2(n14337), .ZN(n11979) );
  XNOR2_X1 U14349 ( .A(n14240), .B(n13856), .ZN(n12014) );
  NAND2_X1 U14350 ( .A1(n11982), .A2(n11981), .ZN(n11983) );
  NAND2_X1 U14351 ( .A1(n11984), .A2(n11983), .ZN(n11986) );
  NAND2_X1 U14352 ( .A1(n11986), .A2(n11985), .ZN(n12020) );
  XNOR2_X1 U14353 ( .A(n14243), .B(n13857), .ZN(n12016) );
  INV_X1 U14354 ( .A(n14160), .ZN(n14157) );
  INV_X1 U14355 ( .A(n14615), .ZN(n14628) );
  NAND4_X1 U14356 ( .A1(n11989), .A2(n10748), .A3(n11988), .A4(n11987), .ZN(
        n11992) );
  NOR3_X1 U14357 ( .A1(n11992), .A2(n11991), .A3(n11990), .ZN(n11994) );
  NAND3_X1 U14358 ( .A1(n11995), .A2(n11994), .A3(n11993), .ZN(n11996) );
  NOR2_X1 U14359 ( .A1(n14628), .A2(n11996), .ZN(n11999) );
  NAND4_X1 U14360 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12001) );
  OR4_X1 U14361 ( .A1(n14219), .A2(n12003), .A3(n12002), .A4(n12001), .ZN(
        n12005) );
  OR4_X1 U14362 ( .A1(n12005), .A2(n14172), .A3(n12004), .A4(n14208), .ZN(
        n12006) );
  OR4_X1 U14363 ( .A1(n14126), .A2(n14157), .A3(n14147), .A4(n12006), .ZN(
        n12007) );
  NOR2_X1 U14364 ( .A1(n14111), .A2(n12007), .ZN(n12008) );
  NAND4_X1 U14365 ( .A1(n12009), .A2(n14103), .A3(n12008), .A4(n14084), .ZN(
        n12010) );
  NOR2_X1 U14366 ( .A1(n14032), .A2(n12010), .ZN(n12012) );
  NAND4_X1 U14367 ( .A1(n13994), .A2(n12012), .A3(n12011), .A4(n14045), .ZN(
        n12013) );
  XNOR2_X1 U14368 ( .A(n12017), .B(n14230), .ZN(n12030) );
  NAND2_X1 U14369 ( .A1(n12019), .A2(n12018), .ZN(n12029) );
  INV_X1 U14370 ( .A(n12020), .ZN(n12025) );
  NAND2_X1 U14371 ( .A1(n13982), .A2(n11903), .ZN(n12033) );
  NAND2_X1 U14372 ( .A1(n12020), .A2(n12029), .ZN(n12035) );
  OAI21_X1 U14373 ( .B1(n13856), .B2(n12035), .A(n12033), .ZN(n12021) );
  OAI21_X1 U14374 ( .B1(n12025), .B2(n12033), .A(n12021), .ZN(n12027) );
  NAND2_X1 U14375 ( .A1(n13856), .A2(n6435), .ZN(n12032) );
  INV_X1 U14376 ( .A(n12035), .ZN(n12022) );
  NAND2_X1 U14377 ( .A1(n13856), .A2(n12022), .ZN(n12023) );
  NAND2_X1 U14378 ( .A1(n12032), .A2(n12023), .ZN(n12024) );
  OAI21_X1 U14379 ( .B1(n12032), .B2(n12025), .A(n12024), .ZN(n12026) );
  MUX2_X1 U14380 ( .A(n12027), .B(n12026), .S(n14240), .Z(n12028) );
  OAI21_X1 U14381 ( .B1(n12030), .B2(n12029), .A(n12028), .ZN(n12031) );
  INV_X1 U14382 ( .A(n12031), .ZN(n12038) );
  INV_X1 U14383 ( .A(n12032), .ZN(n12036) );
  NOR2_X1 U14384 ( .A1(n14240), .A2(n12033), .ZN(n12034) );
  AOI211_X1 U14385 ( .C1(n14240), .C2(n12036), .A(n12035), .B(n12034), .ZN(
        n12037) );
  NAND3_X1 U14386 ( .A1(n12040), .A2(n12039), .A3(n14619), .ZN(n12041) );
  OAI211_X1 U14387 ( .C1(n14357), .C2(n12043), .A(n12041), .B(P1_B_REG_SCAN_IN), .ZN(n12042) );
  OR2_X1 U14388 ( .A1(n15031), .A2(n15090), .ZN(n12045) );
  NOR2_X1 U14389 ( .A1(n12046), .A2(n15083), .ZN(n12464) );
  AOI21_X1 U14390 ( .B1(n15093), .B2(P3_REG2_REG_29__SCAN_IN), .A(n12464), 
        .ZN(n12047) );
  OAI21_X1 U14391 ( .B1(n12048), .B2(n12691), .A(n12047), .ZN(n12049) );
  AOI21_X1 U14392 ( .B1(n12050), .B2(n15059), .A(n12049), .ZN(n12051) );
  OAI21_X1 U14393 ( .B1(n12044), .B2(n15093), .A(n12051), .ZN(P3_U3204) );
  MUX2_X1 U14394 ( .A(n12053), .B(n12052), .S(n15149), .Z(n12054) );
  OAI21_X1 U14395 ( .B1(n12055), .B2(n12769), .A(n12054), .ZN(P3_U3459) );
  INV_X1 U14396 ( .A(n12056), .ZN(n14345) );
  OAI222_X1 U14397 ( .A1(n13588), .A2(n12057), .B1(n13590), .B2(n14345), .C1(
        P2_U3088), .C2(n9159), .ZN(P2_U3299) );
  OR2_X1 U14398 ( .A1(n12092), .A2(n12059), .ZN(n12060) );
  NAND2_X1 U14399 ( .A1(n12061), .A2(n12060), .ZN(n13440) );
  INV_X1 U14400 ( .A(n13439), .ZN(n13451) );
  OR2_X1 U14401 ( .A1(n13543), .A2(n13421), .ZN(n12062) );
  INV_X1 U14402 ( .A(n13434), .ZN(n14494) );
  AND2_X1 U14403 ( .A1(n13538), .A2(n13423), .ZN(n12065) );
  INV_X1 U14404 ( .A(n13388), .ZN(n13395) );
  OR2_X2 U14405 ( .A1(n13394), .A2(n13395), .ZN(n13392) );
  INV_X1 U14406 ( .A(n13103), .ZN(n13006) );
  NAND2_X1 U14407 ( .A1(n13533), .A2(n13006), .ZN(n12066) );
  NAND2_X2 U14408 ( .A1(n13392), .A2(n12066), .ZN(n13373) );
  INV_X1 U14409 ( .A(n13102), .ZN(n12068) );
  OR2_X1 U14410 ( .A1(n13527), .A2(n12068), .ZN(n12067) );
  NAND2_X1 U14411 ( .A1(n13527), .A2(n12068), .ZN(n12069) );
  AND2_X1 U14412 ( .A1(n13522), .A2(n13349), .ZN(n12070) );
  OR2_X1 U14413 ( .A1(n13522), .A2(n13349), .ZN(n12071) );
  INV_X1 U14414 ( .A(n13100), .ZN(n13337) );
  OR2_X1 U14415 ( .A1(n13516), .A2(n13337), .ZN(n12072) );
  OR2_X1 U14416 ( .A1(n13325), .A2(n13336), .ZN(n12075) );
  NAND2_X1 U14417 ( .A1(n13325), .A2(n13336), .ZN(n12076) );
  NAND2_X1 U14418 ( .A1(n12077), .A2(n12076), .ZN(n13297) );
  INV_X1 U14419 ( .A(n13310), .ZN(n13296) );
  INV_X1 U14420 ( .A(n13098), .ZN(n12078) );
  OR2_X1 U14421 ( .A1(n13498), .A2(n12078), .ZN(n12079) );
  NAND2_X1 U14422 ( .A1(n13256), .A2(n13257), .ZN(n13255) );
  INV_X1 U14423 ( .A(n13241), .ZN(n13073) );
  NAND2_X1 U14424 ( .A1(n13472), .A2(n13073), .ZN(n13208) );
  AOI21_X1 U14425 ( .B1(n12086), .B2(P2_B_REG_SCAN_IN), .A(n14885), .ZN(n13195) );
  INV_X1 U14426 ( .A(n13465), .ZN(n13213) );
  INV_X1 U14427 ( .A(n13527), .ZN(n13382) );
  INV_X1 U14428 ( .A(n13462), .ZN(n12091) );
  AOI22_X1 U14429 ( .A1(n12089), .A2(n14865), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13456), .ZN(n12090) );
  OAI21_X1 U14430 ( .B1(n12091), .B2(n14874), .A(n12090), .ZN(n12120) );
  AND2_X1 U14431 ( .A1(n12092), .A2(n13445), .ZN(n12093) );
  NOR2_X1 U14432 ( .A1(n13543), .A2(n13105), .ZN(n12095) );
  NAND2_X1 U14433 ( .A1(n13543), .A2(n13105), .ZN(n12096) );
  AND2_X1 U14434 ( .A1(n13434), .A2(n13442), .ZN(n12098) );
  OR2_X1 U14435 ( .A1(n13434), .A2(n13442), .ZN(n12097) );
  OR2_X1 U14436 ( .A1(n13538), .A2(n13104), .ZN(n12099) );
  NAND2_X1 U14437 ( .A1(n13363), .A2(n13364), .ZN(n13362) );
  OR2_X1 U14438 ( .A1(n13522), .A2(n13101), .ZN(n12103) );
  OR2_X1 U14439 ( .A1(n13516), .A2(n13100), .ZN(n12104) );
  NOR2_X1 U14440 ( .A1(n13511), .A2(n13099), .ZN(n12105) );
  NAND2_X1 U14441 ( .A1(n13511), .A2(n13099), .ZN(n12106) );
  AND2_X1 U14442 ( .A1(n13325), .A2(n13300), .ZN(n12107) );
  NAND2_X1 U14443 ( .A1(n13498), .A2(n13098), .ZN(n12108) );
  OR2_X1 U14444 ( .A1(n13492), .A2(n13301), .ZN(n12109) );
  NAND2_X1 U14445 ( .A1(n13292), .A2(n12109), .ZN(n12111) );
  NAND2_X1 U14446 ( .A1(n13492), .A2(n13301), .ZN(n12110) );
  NAND2_X1 U14447 ( .A1(n13279), .A2(n13278), .ZN(n12113) );
  NAND2_X1 U14448 ( .A1(n13487), .A2(n13258), .ZN(n12112) );
  AND2_X1 U14449 ( .A1(n13482), .A2(n13240), .ZN(n12114) );
  NAND2_X1 U14450 ( .A1(n13477), .A2(n13259), .ZN(n12115) );
  INV_X1 U14451 ( .A(n13472), .ZN(n13234) );
  NAND2_X1 U14452 ( .A1(n13465), .A2(n13227), .ZN(n12116) );
  NAND2_X1 U14453 ( .A1(n12117), .A2(n12116), .ZN(n12119) );
  INV_X1 U14454 ( .A(n12121), .ZN(n12123) );
  OAI222_X1 U14455 ( .A1(n8191), .A2(P3_U3151), .B1(n14378), .B2(n12123), .C1(
        n12122), .C2(n14376), .ZN(P3_U3267) );
  OAI222_X1 U14456 ( .A1(n8467), .A2(P2_U3088), .B1(n13590), .B2(n12125), .C1(
        n12124), .C2(n13588), .ZN(P2_U3297) );
  XNOR2_X1 U14457 ( .A(n12482), .B(n10597), .ZN(n12205) );
  OR2_X1 U14458 ( .A1(n12356), .A2(n12126), .ZN(n12127) );
  XNOR2_X1 U14459 ( .A(n12129), .B(n12159), .ZN(n12130) );
  XNOR2_X1 U14460 ( .A(n12130), .B(n14467), .ZN(n12190) );
  INV_X1 U14461 ( .A(n12130), .ZN(n12131) );
  NAND2_X1 U14462 ( .A1(n12131), .A2(n14467), .ZN(n12132) );
  XNOR2_X1 U14463 ( .A(n12302), .B(n10597), .ZN(n12225) );
  INV_X1 U14464 ( .A(n14468), .ZN(n12228) );
  XNOR2_X1 U14465 ( .A(n14479), .B(n12159), .ZN(n12229) );
  AOI22_X1 U14466 ( .A1(n12309), .A2(n12225), .B1(n12228), .B2(n12229), .ZN(
        n12133) );
  OR2_X1 U14467 ( .A1(n12309), .A2(n12225), .ZN(n12134) );
  INV_X1 U14468 ( .A(n12134), .ZN(n12137) );
  NAND2_X1 U14469 ( .A1(n12134), .A2(n12228), .ZN(n12136) );
  INV_X1 U14470 ( .A(n12229), .ZN(n12135) );
  AOI22_X1 U14471 ( .A1(n12137), .A2(n14468), .B1(n12136), .B2(n12135), .ZN(
        n12138) );
  XNOR2_X1 U14472 ( .A(n12845), .B(n12159), .ZN(n12139) );
  INV_X1 U14473 ( .A(n12687), .ZN(n12179) );
  NAND2_X1 U14474 ( .A1(n12139), .A2(n12179), .ZN(n12283) );
  INV_X1 U14475 ( .A(n12139), .ZN(n12140) );
  NAND2_X1 U14476 ( .A1(n12140), .A2(n12687), .ZN(n12284) );
  XNOR2_X1 U14477 ( .A(n12841), .B(n10597), .ZN(n12142) );
  XNOR2_X1 U14478 ( .A(n12142), .B(n12341), .ZN(n12177) );
  NAND2_X1 U14479 ( .A1(n12142), .A2(n12673), .ZN(n12143) );
  XNOR2_X1 U14480 ( .A(n12837), .B(n10597), .ZN(n12334) );
  XNOR2_X1 U14481 ( .A(n12831), .B(n10597), .ZN(n12144) );
  NAND2_X1 U14482 ( .A1(n12144), .A2(n12615), .ZN(n12246) );
  INV_X1 U14483 ( .A(n12144), .ZN(n12145) );
  NAND2_X1 U14484 ( .A1(n12145), .A2(n12646), .ZN(n12247) );
  XNOR2_X1 U14485 ( .A(n12828), .B(n10597), .ZN(n12146) );
  XNOR2_X1 U14486 ( .A(n12146), .B(n12603), .ZN(n12257) );
  NAND2_X1 U14487 ( .A1(n12146), .A2(n12628), .ZN(n12147) );
  XNOR2_X1 U14488 ( .A(n12313), .B(n10597), .ZN(n12148) );
  XNOR2_X1 U14489 ( .A(n12148), .B(n12589), .ZN(n12315) );
  INV_X1 U14490 ( .A(n12148), .ZN(n12149) );
  NAND2_X1 U14491 ( .A1(n12149), .A2(n12589), .ZN(n12150) );
  NAND2_X1 U14492 ( .A1(n12314), .A2(n12150), .ZN(n12200) );
  XNOR2_X1 U14493 ( .A(n12197), .B(n10597), .ZN(n12151) );
  XNOR2_X1 U14494 ( .A(n12151), .B(n12355), .ZN(n12199) );
  INV_X1 U14495 ( .A(n12151), .ZN(n12152) );
  NAND2_X1 U14496 ( .A1(n12152), .A2(n12355), .ZN(n12153) );
  XNOR2_X1 U14497 ( .A(n12815), .B(n10597), .ZN(n12154) );
  XNOR2_X1 U14498 ( .A(n12154), .B(n12590), .ZN(n12275) );
  INV_X1 U14499 ( .A(n12154), .ZN(n12155) );
  NAND2_X1 U14500 ( .A1(n12155), .A2(n12590), .ZN(n12156) );
  XNOR2_X1 U14501 ( .A(n12565), .B(n10597), .ZN(n12157) );
  XNOR2_X1 U14502 ( .A(n12157), .B(n12574), .ZN(n12219) );
  NAND2_X1 U14503 ( .A1(n12157), .A2(n12574), .ZN(n12158) );
  XNOR2_X1 U14504 ( .A(n12298), .B(n12159), .ZN(n12160) );
  INV_X1 U14505 ( .A(n12160), .ZN(n12161) );
  AND2_X1 U14506 ( .A1(n12162), .A2(n12161), .ZN(n12163) );
  XNOR2_X1 U14507 ( .A(n12525), .B(n10597), .ZN(n12266) );
  XNOR2_X1 U14508 ( .A(n12540), .B(n10597), .ZN(n12164) );
  OAI22_X1 U14509 ( .A1(n12266), .A2(n12536), .B1(n12549), .B2(n12164), .ZN(
        n12168) );
  NAND3_X1 U14510 ( .A1(n12164), .A2(n12549), .A3(n12536), .ZN(n12167) );
  INV_X1 U14511 ( .A(n12164), .ZN(n12263) );
  OAI21_X1 U14512 ( .B1(n12263), .B2(n12265), .A(n12351), .ZN(n12165) );
  NAND2_X1 U14513 ( .A1(n12266), .A2(n12165), .ZN(n12166) );
  XNOR2_X1 U14514 ( .A(n12511), .B(n10597), .ZN(n12169) );
  XNOR2_X1 U14515 ( .A(n12169), .B(n12489), .ZN(n12240) );
  XNOR2_X1 U14516 ( .A(n12496), .B(n10597), .ZN(n12170) );
  XNOR2_X1 U14517 ( .A(n12170), .B(n12507), .ZN(n12322) );
  AOI22_X1 U14518 ( .A1(n12350), .A2(n12323), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12172) );
  NAND2_X1 U14519 ( .A1(n12483), .A2(n12324), .ZN(n12171) );
  OAI211_X1 U14520 ( .C1(n12478), .C2(n12327), .A(n12172), .B(n12171), .ZN(
        n12173) );
  AOI21_X1 U14521 ( .B1(n12482), .B2(n12330), .A(n12173), .ZN(n12174) );
  OAI21_X1 U14522 ( .B1(n12175), .B2(n12332), .A(n12174), .ZN(P3_U3154) );
  OAI211_X1 U14523 ( .C1(n12178), .C2(n12177), .A(n12176), .B(n12337), .ZN(
        n12183) );
  NOR2_X1 U14524 ( .A1(n12339), .A2(n12662), .ZN(n12181) );
  NAND2_X1 U14525 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12381)
         );
  OAI21_X1 U14526 ( .B1(n12179), .B2(n12340), .A(n12381), .ZN(n12180) );
  AOI211_X1 U14527 ( .C1(n12344), .C2(n12659), .A(n12181), .B(n12180), .ZN(
        n12182) );
  OAI211_X1 U14528 ( .C1(n12347), .C2(n12841), .A(n12183), .B(n12182), .ZN(
        P3_U3155) );
  AOI22_X1 U14529 ( .A1(n12351), .A2(n12344), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12185) );
  NAND2_X1 U14530 ( .A1(n12324), .A2(n12541), .ZN(n12184) );
  OAI211_X1 U14531 ( .C1(n12564), .C2(n12340), .A(n12185), .B(n12184), .ZN(
        n12186) );
  AOI21_X1 U14532 ( .B1(n12540), .B2(n12330), .A(n12186), .ZN(n12187) );
  OAI21_X1 U14533 ( .B1(n12188), .B2(n12332), .A(n12187), .ZN(P3_U3156) );
  OAI211_X1 U14534 ( .C1(n6585), .C2(n12190), .A(n12189), .B(n12337), .ZN(
        n12195) );
  AND2_X1 U14535 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n15006) );
  OAI22_X1 U14536 ( .A1(n12191), .A2(n12340), .B1(n12309), .B2(n12327), .ZN(
        n12192) );
  AOI211_X1 U14537 ( .C1(n12193), .C2(n12330), .A(n15006), .B(n12192), .ZN(
        n12194) );
  OAI211_X1 U14538 ( .C1(n12196), .C2(n12339), .A(n12195), .B(n12194), .ZN(
        P3_U3157) );
  INV_X1 U14539 ( .A(n12197), .ZN(n12820) );
  OAI211_X1 U14540 ( .C1(n12200), .C2(n12199), .A(n12198), .B(n12337), .ZN(
        n12204) );
  NAND2_X1 U14541 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12458)
         );
  OAI21_X1 U14542 ( .B1(n12563), .B2(n12327), .A(n12458), .ZN(n12202) );
  NOR2_X1 U14543 ( .A1(n12339), .A2(n12593), .ZN(n12201) );
  AOI211_X1 U14544 ( .C1(n12323), .C2(n12589), .A(n12202), .B(n12201), .ZN(
        n12203) );
  OAI211_X1 U14545 ( .C1(n12820), .C2(n12347), .A(n12204), .B(n12203), .ZN(
        P3_U3159) );
  XNOR2_X1 U14546 ( .A(n12206), .B(n10597), .ZN(n12207) );
  INV_X1 U14547 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12208) );
  OAI22_X1 U14548 ( .A1(n12328), .A2(n12340), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12208), .ZN(n12212) );
  INV_X1 U14549 ( .A(n12468), .ZN(n12209) );
  OAI22_X1 U14550 ( .A1(n12210), .A2(n12327), .B1(n12209), .B2(n12339), .ZN(
        n12211) );
  AOI211_X1 U14551 ( .C1(n12213), .C2(n12330), .A(n12212), .B(n12211), .ZN(
        n12214) );
  OAI21_X1 U14552 ( .B1(n12215), .B2(n12332), .A(n12214), .ZN(P3_U3160) );
  INV_X1 U14553 ( .A(n12216), .ZN(n12217) );
  AOI21_X1 U14554 ( .B1(n12219), .B2(n12218), .A(n12217), .ZN(n12224) );
  AOI22_X1 U14555 ( .A1(n12590), .A2(n12323), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12221) );
  NAND2_X1 U14556 ( .A1(n12324), .A2(n12566), .ZN(n12220) );
  OAI211_X1 U14557 ( .C1(n12564), .C2(n12327), .A(n12221), .B(n12220), .ZN(
        n12222) );
  AOI21_X1 U14558 ( .B1(n12565), .B2(n12330), .A(n12222), .ZN(n12223) );
  OAI21_X1 U14559 ( .B1(n12224), .B2(n12332), .A(n12223), .ZN(P3_U3163) );
  INV_X1 U14560 ( .A(n12225), .ZN(n12226) );
  XOR2_X1 U14561 ( .A(n12225), .B(n12227), .Z(n12308) );
  NOR2_X1 U14562 ( .A1(n12308), .A2(n12309), .ZN(n12307) );
  AOI21_X1 U14563 ( .B1(n12227), .B2(n12226), .A(n12307), .ZN(n12231) );
  XNOR2_X1 U14564 ( .A(n12229), .B(n12228), .ZN(n12230) );
  XNOR2_X1 U14565 ( .A(n12231), .B(n12230), .ZN(n12238) );
  NOR2_X1 U14566 ( .A1(n12339), .A2(n12692), .ZN(n12235) );
  AOI21_X1 U14567 ( .B1(n12344), .B2(n12687), .A(n12232), .ZN(n12233) );
  OAI21_X1 U14568 ( .B1(n12309), .B2(n12340), .A(n12233), .ZN(n12234) );
  AOI211_X1 U14569 ( .C1(n12236), .C2(n12330), .A(n12235), .B(n12234), .ZN(
        n12237) );
  OAI21_X1 U14570 ( .B1(n12238), .B2(n12332), .A(n12237), .ZN(P3_U3164) );
  XOR2_X1 U14571 ( .A(n12240), .B(n12239), .Z(n12245) );
  AOI22_X1 U14572 ( .A1(n12351), .A2(n12323), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12242) );
  NAND2_X1 U14573 ( .A1(n12512), .A2(n12324), .ZN(n12241) );
  OAI211_X1 U14574 ( .C1(n12507), .C2(n12327), .A(n12242), .B(n12241), .ZN(
        n12243) );
  AOI21_X1 U14575 ( .B1(n12511), .B2(n12330), .A(n12243), .ZN(n12244) );
  OAI21_X1 U14576 ( .B1(n12245), .B2(n12332), .A(n12244), .ZN(P3_U3165) );
  NAND2_X1 U14577 ( .A1(n12247), .A2(n12246), .ZN(n12249) );
  XOR2_X1 U14578 ( .A(n12249), .B(n12248), .Z(n12255) );
  NAND2_X1 U14579 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12424)
         );
  OAI21_X1 U14580 ( .B1(n12250), .B2(n12340), .A(n12424), .ZN(n12251) );
  AOI21_X1 U14581 ( .B1(n12344), .B2(n12628), .A(n12251), .ZN(n12252) );
  OAI21_X1 U14582 ( .B1(n12636), .B2(n12339), .A(n12252), .ZN(n12253) );
  AOI21_X1 U14583 ( .B1(n12831), .B2(n12330), .A(n12253), .ZN(n12254) );
  OAI21_X1 U14584 ( .B1(n12255), .B2(n12332), .A(n12254), .ZN(P3_U3166) );
  OAI211_X1 U14585 ( .C1(n12258), .C2(n12257), .A(n12256), .B(n12337), .ZN(
        n12262) );
  NAND2_X1 U14586 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14436)
         );
  OAI21_X1 U14587 ( .B1(n12618), .B2(n12327), .A(n14436), .ZN(n12260) );
  NOR2_X1 U14588 ( .A1(n12339), .A2(n12619), .ZN(n12259) );
  AOI211_X1 U14589 ( .C1(n12323), .C2(n12646), .A(n12260), .B(n12259), .ZN(
        n12261) );
  OAI211_X1 U14590 ( .C1(n12347), .C2(n12828), .A(n12262), .B(n12261), .ZN(
        P3_U3168) );
  XNOR2_X1 U14591 ( .A(n12266), .B(n12536), .ZN(n12267) );
  XNOR2_X1 U14592 ( .A(n12268), .B(n12267), .ZN(n12273) );
  AOI22_X1 U14593 ( .A1(n12489), .A2(n12344), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12270) );
  NAND2_X1 U14594 ( .A1(n12324), .A2(n12526), .ZN(n12269) );
  OAI211_X1 U14595 ( .C1(n12549), .C2(n12340), .A(n12270), .B(n12269), .ZN(
        n12271) );
  AOI21_X1 U14596 ( .B1(n12525), .B2(n12330), .A(n12271), .ZN(n12272) );
  OAI21_X1 U14597 ( .B1(n12273), .B2(n12332), .A(n12272), .ZN(P3_U3169) );
  INV_X1 U14598 ( .A(n12815), .ZN(n12282) );
  OAI211_X1 U14599 ( .C1(n12276), .C2(n12275), .A(n12274), .B(n12337), .ZN(
        n12281) );
  INV_X1 U14600 ( .A(n12578), .ZN(n12279) );
  AOI22_X1 U14601 ( .A1(n12354), .A2(n12344), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12277) );
  OAI21_X1 U14602 ( .B1(n12604), .B2(n12340), .A(n12277), .ZN(n12278) );
  AOI21_X1 U14603 ( .B1(n12279), .B2(n12324), .A(n12278), .ZN(n12280) );
  OAI211_X1 U14604 ( .C1(n12282), .C2(n12347), .A(n12281), .B(n12280), .ZN(
        P3_U3173) );
  NAND2_X1 U14605 ( .A1(n12284), .A2(n12283), .ZN(n12286) );
  XOR2_X1 U14606 ( .A(n12286), .B(n12285), .Z(n12293) );
  AOI21_X1 U14607 ( .B1(n12344), .B2(n12673), .A(n12287), .ZN(n12289) );
  NAND2_X1 U14608 ( .A1(n12323), .A2(n14468), .ZN(n12288) );
  OAI211_X1 U14609 ( .C1(n12339), .C2(n12676), .A(n12289), .B(n12288), .ZN(
        n12290) );
  AOI21_X1 U14610 ( .B1(n12291), .B2(n12330), .A(n12290), .ZN(n12292) );
  OAI21_X1 U14611 ( .B1(n12293), .B2(n12332), .A(n12292), .ZN(P3_U3174) );
  XNOR2_X1 U14612 ( .A(n12294), .B(n12353), .ZN(n12301) );
  INV_X1 U14613 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n12295) );
  OAI22_X1 U14614 ( .A1(n12574), .A2(n12340), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12295), .ZN(n12297) );
  NOR2_X1 U14615 ( .A1(n12549), .A2(n12327), .ZN(n12296) );
  AOI211_X1 U14616 ( .C1(n12552), .C2(n12324), .A(n12297), .B(n12296), .ZN(
        n12300) );
  NAND2_X1 U14617 ( .A1(n12298), .A2(n12330), .ZN(n12299) );
  OAI211_X1 U14618 ( .C1(n12301), .C2(n12332), .A(n12300), .B(n12299), .ZN(
        P3_U3175) );
  NAND2_X1 U14619 ( .A1(n12323), .A2(n14467), .ZN(n12306) );
  NAND2_X1 U14620 ( .A1(n12344), .A2(n14468), .ZN(n12305) );
  NAND2_X1 U14621 ( .A1(n12330), .A2(n12302), .ZN(n12304) );
  NAND4_X1 U14622 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12311) );
  AOI211_X1 U14623 ( .C1(n12309), .C2(n12308), .A(n12332), .B(n12307), .ZN(
        n12310) );
  AOI211_X1 U14624 ( .C1(n14470), .C2(n12324), .A(n12311), .B(n12310), .ZN(
        n12312) );
  INV_X1 U14625 ( .A(n12312), .ZN(P3_U3176) );
  INV_X1 U14626 ( .A(n12313), .ZN(n12824) );
  OAI211_X1 U14627 ( .C1(n12316), .C2(n12315), .A(n12314), .B(n12337), .ZN(
        n12321) );
  INV_X1 U14628 ( .A(n12317), .ZN(n12605) );
  AND2_X1 U14629 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14451) );
  AOI21_X1 U14630 ( .B1(n12355), .B2(n12344), .A(n14451), .ZN(n12318) );
  OAI21_X1 U14631 ( .B1(n12603), .B2(n12340), .A(n12318), .ZN(n12319) );
  AOI21_X1 U14632 ( .B1(n12605), .B2(n12324), .A(n12319), .ZN(n12320) );
  OAI211_X1 U14633 ( .C1(n12824), .C2(n12347), .A(n12321), .B(n12320), .ZN(
        P3_U3178) );
  AOI22_X1 U14634 ( .A1(n12489), .A2(n12323), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12326) );
  NAND2_X1 U14635 ( .A1(n12497), .A2(n12324), .ZN(n12325) );
  OAI211_X1 U14636 ( .C1(n12328), .C2(n12327), .A(n12326), .B(n12325), .ZN(
        n12329) );
  AOI21_X1 U14637 ( .B1(n12496), .B2(n12330), .A(n12329), .ZN(n12331) );
  OAI21_X1 U14638 ( .B1(n12333), .B2(n12332), .A(n12331), .ZN(P3_U3180) );
  XNOR2_X1 U14639 ( .A(n12334), .B(n12659), .ZN(n12335) );
  XNOR2_X1 U14640 ( .A(n12336), .B(n12335), .ZN(n12338) );
  NAND2_X1 U14641 ( .A1(n12338), .A2(n12337), .ZN(n12346) );
  NOR2_X1 U14642 ( .A1(n12339), .A2(n12649), .ZN(n12343) );
  NAND2_X1 U14643 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12394)
         );
  OAI21_X1 U14644 ( .B1(n12341), .B2(n12340), .A(n12394), .ZN(n12342) );
  AOI211_X1 U14645 ( .C1(n12344), .C2(n12646), .A(n12343), .B(n12342), .ZN(
        n12345) );
  OAI211_X1 U14646 ( .C1(n12347), .C2(n12837), .A(n12346), .B(n12345), .ZN(
        P3_U3181) );
  MUX2_X1 U14647 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12463), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14648 ( .A(n12348), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12352), .Z(
        P3_U3521) );
  MUX2_X1 U14649 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12349), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14650 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12490), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14651 ( .A(n12350), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12352), .Z(
        P3_U3517) );
  MUX2_X1 U14652 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12489), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14653 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12351), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14654 ( .A(n12353), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12352), .Z(
        P3_U3513) );
  MUX2_X1 U14655 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12354), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14656 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12590), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14657 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12355), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14658 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12589), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14659 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12628), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14660 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12646), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14661 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12659), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14662 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12673), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14663 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12687), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14664 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n14468), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14665 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12688), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14666 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n14467), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14667 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12356), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14668 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12357), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14669 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12358), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14670 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n15029), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14671 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12359), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14672 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n15030), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14673 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15067), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14674 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12772), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14675 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n15068), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14676 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n6905), .S(P3_U3897), .Z(
        P3_U3491) );
  NOR2_X1 U14677 ( .A1(n12365), .A2(n12360), .ZN(n12362) );
  NAND2_X1 U14678 ( .A1(n12368), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12398) );
  OAI21_X1 U14679 ( .B1(n12368), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12398), 
        .ZN(n12367) );
  AOI21_X1 U14680 ( .B1(n12363), .B2(n12367), .A(n12389), .ZN(n12388) );
  INV_X1 U14681 ( .A(n12364), .ZN(n12366) );
  NAND2_X1 U14682 ( .A1(n12366), .A2(n12365), .ZN(n12371) );
  AND2_X1 U14683 ( .A1(n12372), .A2(n12371), .ZN(n12374) );
  INV_X1 U14684 ( .A(n12367), .ZN(n12370) );
  INV_X1 U14685 ( .A(n12368), .ZN(n12380) );
  NAND2_X1 U14686 ( .A1(n12368), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12397) );
  INV_X1 U14687 ( .A(n12397), .ZN(n12369) );
  AOI21_X1 U14688 ( .B1(n12380), .B2(n12763), .A(n12369), .ZN(n12378) );
  MUX2_X1 U14689 ( .A(n12370), .B(n12378), .S(n11248), .Z(n12373) );
  NAND3_X1 U14690 ( .A1(n12372), .A2(n12371), .A3(n12373), .ZN(n12400) );
  OAI211_X1 U14691 ( .C1(n12374), .C2(n12373), .A(n15015), .B(n12400), .ZN(
        n12387) );
  NAND2_X1 U14692 ( .A1(n14382), .A2(n12375), .ZN(n12377) );
  NAND2_X1 U14693 ( .A1(n12377), .A2(n12376), .ZN(n12379) );
  NAND2_X1 U14694 ( .A1(n12378), .A2(n12379), .ZN(n12392) );
  OAI21_X1 U14695 ( .B1(n12379), .B2(n12378), .A(n12392), .ZN(n12385) );
  NAND2_X1 U14696 ( .A1(n15017), .A2(n12380), .ZN(n12382) );
  OAI211_X1 U14697 ( .C1(n12383), .C2(n15024), .A(n12382), .B(n12381), .ZN(
        n12384) );
  AOI21_X1 U14698 ( .B1(n12385), .B2(n15007), .A(n12384), .ZN(n12386) );
  OAI211_X1 U14699 ( .C1(n12388), .C2(n15001), .A(n12387), .B(n12386), .ZN(
        P3_U3196) );
  INV_X1 U14700 ( .A(n14391), .ZN(n12414) );
  AOI21_X1 U14701 ( .B1(n12391), .B2(n12390), .A(n12410), .ZN(n12408) );
  NAND2_X1 U14702 ( .A1(n12397), .A2(n12392), .ZN(n12419) );
  XNOR2_X1 U14703 ( .A(n12414), .B(n12419), .ZN(n12393) );
  NAND2_X1 U14704 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12393), .ZN(n12420) );
  OAI21_X1 U14705 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12393), .A(n12420), 
        .ZN(n12406) );
  NAND2_X1 U14706 ( .A1(n15017), .A2(n12414), .ZN(n12395) );
  OAI211_X1 U14707 ( .C1(n12396), .C2(n15024), .A(n12395), .B(n12394), .ZN(
        n12405) );
  MUX2_X1 U14708 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n11248), .Z(n12402) );
  MUX2_X1 U14709 ( .A(n12398), .B(n12397), .S(n11248), .Z(n12399) );
  AOI21_X1 U14710 ( .B1(n12402), .B2(n12401), .A(n12413), .ZN(n12403) );
  NOR2_X1 U14711 ( .A1(n12403), .A2(n14991), .ZN(n12404) );
  AOI211_X1 U14712 ( .C1(n15007), .C2(n12406), .A(n12405), .B(n12404), .ZN(
        n12407) );
  OAI21_X1 U14713 ( .B1(n12408), .B2(n15001), .A(n12407), .ZN(P3_U3197) );
  AND2_X1 U14714 ( .A1(n14391), .A2(n12409), .ZN(n12411) );
  AOI22_X1 U14715 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12449), .B1(n12433), 
        .B2(n12637), .ZN(n12412) );
  AOI21_X1 U14716 ( .B1(n6546), .B2(n12412), .A(n12432), .ZN(n12431) );
  MUX2_X1 U14717 ( .A(n12637), .B(n12448), .S(n11248), .Z(n12415) );
  NOR2_X1 U14718 ( .A1(n12415), .A2(n12449), .ZN(n12440) );
  INV_X1 U14719 ( .A(n12440), .ZN(n12416) );
  NAND2_X1 U14720 ( .A1(n12415), .A2(n12449), .ZN(n12439) );
  NAND2_X1 U14721 ( .A1(n12416), .A2(n12439), .ZN(n12417) );
  XNOR2_X1 U14722 ( .A(n12441), .B(n12417), .ZN(n12418) );
  NAND2_X1 U14723 ( .A1(n12418), .A2(n15015), .ZN(n12430) );
  AOI22_X1 U14724 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12433), .B1(n12449), 
        .B2(n12448), .ZN(n12423) );
  NAND2_X1 U14725 ( .A1(n14391), .A2(n12419), .ZN(n12421) );
  NAND2_X1 U14726 ( .A1(n12421), .A2(n12420), .ZN(n12422) );
  NAND2_X1 U14727 ( .A1(n12423), .A2(n12422), .ZN(n12447) );
  OAI21_X1 U14728 ( .B1(n12423), .B2(n12422), .A(n12447), .ZN(n12428) );
  NOR2_X1 U14729 ( .A1(n14989), .A2(n12433), .ZN(n12427) );
  OAI21_X1 U14730 ( .B1(n15024), .B2(n12425), .A(n12424), .ZN(n12426) );
  AOI211_X1 U14731 ( .C1(n12428), .C2(n15007), .A(n12427), .B(n12426), .ZN(
        n12429) );
  OAI211_X1 U14732 ( .C1(n12431), .C2(n15001), .A(n12430), .B(n12429), .ZN(
        P3_U3198) );
  INV_X1 U14733 ( .A(n12450), .ZN(n14435) );
  XNOR2_X1 U14734 ( .A(n14435), .B(n12434), .ZN(n14431) );
  INV_X1 U14735 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12435) );
  NAND2_X1 U14736 ( .A1(n14449), .A2(n12435), .ZN(n12437) );
  NAND2_X1 U14737 ( .A1(n12453), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12436) );
  AND2_X1 U14738 ( .A1(n12437), .A2(n12436), .ZN(n14447) );
  XNOR2_X1 U14739 ( .A(n12459), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12444) );
  INV_X1 U14740 ( .A(n12444), .ZN(n12438) );
  MUX2_X1 U14741 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n11248), .Z(n12442) );
  OAI21_X1 U14742 ( .B1(n12441), .B2(n12440), .A(n12439), .ZN(n14440) );
  XNOR2_X1 U14743 ( .A(n12442), .B(n12450), .ZN(n14441) );
  NOR2_X1 U14744 ( .A1(n14440), .A2(n14441), .ZN(n14439) );
  AOI21_X1 U14745 ( .B1(n12442), .B2(n12450), .A(n14439), .ZN(n12443) );
  XNOR2_X1 U14746 ( .A(n12443), .B(n12453), .ZN(n14453) );
  MUX2_X1 U14747 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n11248), .Z(n14454) );
  NOR2_X1 U14748 ( .A1(n14453), .A2(n14454), .ZN(n14452) );
  AOI21_X1 U14749 ( .B1(n12443), .B2(n12453), .A(n14452), .ZN(n12446) );
  XNOR2_X1 U14750 ( .A(n12459), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12454) );
  MUX2_X1 U14751 ( .A(n12444), .B(n12454), .S(n11248), .Z(n12445) );
  NAND2_X1 U14752 ( .A1(n12450), .A2(n12451), .ZN(n12452) );
  XNOR2_X1 U14753 ( .A(n12451), .B(n14435), .ZN(n14434) );
  NAND2_X1 U14754 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14434), .ZN(n14433) );
  NAND2_X1 U14755 ( .A1(n12452), .A2(n14433), .ZN(n14457) );
  XNOR2_X1 U14756 ( .A(n12453), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U14757 ( .A1(n14457), .A2(n14456), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n14449), .ZN(n12456) );
  INV_X1 U14758 ( .A(n12454), .ZN(n12455) );
  NAND2_X1 U14759 ( .A1(n14995), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12457) );
  OAI211_X1 U14760 ( .C1(n14989), .C2(n12459), .A(n12458), .B(n12457), .ZN(
        n12460) );
  NAND2_X1 U14761 ( .A1(n12461), .A2(n14462), .ZN(n12465) );
  NAND2_X1 U14762 ( .A1(n12463), .A2(n12462), .ZN(n12783) );
  INV_X1 U14763 ( .A(n12783), .ZN(n14476) );
  AOI21_X1 U14764 ( .B1(n14476), .B2(n15091), .A(n12464), .ZN(n14464) );
  OAI211_X1 U14765 ( .C1(n15091), .C2(n12466), .A(n12465), .B(n14464), .ZN(
        P3_U3202) );
  INV_X1 U14766 ( .A(n12467), .ZN(n12473) );
  AOI22_X1 U14767 ( .A1(n12468), .A2(n15053), .B1(n15093), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12469) );
  OAI21_X1 U14768 ( .B1(n12704), .B2(n12691), .A(n12469), .ZN(n12470) );
  AOI21_X1 U14769 ( .B1(n12471), .B2(n15091), .A(n12470), .ZN(n12472) );
  OAI21_X1 U14770 ( .B1(n12473), .B2(n12697), .A(n12472), .ZN(P3_U3205) );
  XNOR2_X1 U14771 ( .A(n12474), .B(n12476), .ZN(n12481) );
  OAI21_X1 U14772 ( .B1(n12477), .B2(n12476), .A(n12475), .ZN(n12706) );
  OAI22_X1 U14773 ( .A1(n12478), .A2(n15046), .B1(n12507), .B2(n15048), .ZN(
        n12479) );
  AOI21_X1 U14774 ( .B1(n12706), .B2(n15031), .A(n12479), .ZN(n12480) );
  OAI21_X1 U14775 ( .B1(n15043), .B2(n12481), .A(n12480), .ZN(n12705) );
  INV_X1 U14776 ( .A(n12705), .ZN(n12487) );
  INV_X1 U14777 ( .A(n12482), .ZN(n12789) );
  AOI22_X1 U14778 ( .A1(n12483), .A2(n15053), .B1(n15093), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12484) );
  OAI21_X1 U14779 ( .B1(n12789), .B2(n12691), .A(n12484), .ZN(n12485) );
  AOI21_X1 U14780 ( .B1(n12706), .B2(n12544), .A(n12485), .ZN(n12486) );
  OAI21_X1 U14781 ( .B1(n12487), .B2(n15093), .A(n12486), .ZN(P3_U3206) );
  XOR2_X1 U14782 ( .A(n12491), .B(n12488), .Z(n12495) );
  AOI22_X1 U14783 ( .A1(n12490), .A2(n15066), .B1(n15069), .B2(n12489), .ZN(
        n12494) );
  XNOR2_X1 U14784 ( .A(n12492), .B(n12491), .ZN(n12710) );
  NAND2_X1 U14785 ( .A1(n12710), .A2(n15031), .ZN(n12493) );
  OAI211_X1 U14786 ( .C1(n12495), .C2(n15043), .A(n12494), .B(n12493), .ZN(
        n12709) );
  INV_X1 U14787 ( .A(n12709), .ZN(n12501) );
  INV_X1 U14788 ( .A(n12496), .ZN(n12793) );
  AOI22_X1 U14789 ( .A1(n12497), .A2(n15053), .B1(n15093), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12498) );
  OAI21_X1 U14790 ( .B1(n12793), .B2(n12691), .A(n12498), .ZN(n12499) );
  AOI21_X1 U14791 ( .B1(n12710), .B2(n12544), .A(n12499), .ZN(n12500) );
  OAI21_X1 U14792 ( .B1(n12501), .B2(n15093), .A(n12500), .ZN(P3_U3207) );
  XNOR2_X1 U14793 ( .A(n12502), .B(n12503), .ZN(n12510) );
  OAI21_X1 U14794 ( .B1(n12506), .B2(n12505), .A(n12504), .ZN(n12714) );
  OAI22_X1 U14795 ( .A1(n12507), .A2(n15046), .B1(n12536), .B2(n15048), .ZN(
        n12508) );
  AOI21_X1 U14796 ( .B1(n12714), .B2(n15031), .A(n12508), .ZN(n12509) );
  OAI21_X1 U14797 ( .B1(n15043), .B2(n12510), .A(n12509), .ZN(n12713) );
  INV_X1 U14798 ( .A(n12713), .ZN(n12516) );
  AOI22_X1 U14799 ( .A1(n12512), .A2(n15053), .B1(n15093), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12513) );
  OAI21_X1 U14800 ( .B1(n7400), .B2(n12691), .A(n12513), .ZN(n12514) );
  AOI21_X1 U14801 ( .B1(n12714), .B2(n12544), .A(n12514), .ZN(n12515) );
  OAI21_X1 U14802 ( .B1(n12516), .B2(n15093), .A(n12515), .ZN(P3_U3208) );
  XNOR2_X1 U14803 ( .A(n12517), .B(n12521), .ZN(n12518) );
  OAI222_X1 U14804 ( .A1(n15046), .A2(n12519), .B1(n15048), .B2(n12549), .C1(
        n12518), .C2(n15043), .ZN(n12717) );
  INV_X1 U14805 ( .A(n12717), .ZN(n12530) );
  INV_X1 U14806 ( .A(n12520), .ZN(n12533) );
  OAI21_X1 U14807 ( .B1(n12533), .B2(n12522), .A(n12521), .ZN(n12524) );
  NAND2_X1 U14808 ( .A1(n12524), .A2(n12523), .ZN(n12718) );
  INV_X1 U14809 ( .A(n12525), .ZN(n12800) );
  AOI22_X1 U14810 ( .A1(n15093), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12526), 
        .B2(n15053), .ZN(n12527) );
  OAI21_X1 U14811 ( .B1(n12800), .B2(n12691), .A(n12527), .ZN(n12528) );
  AOI21_X1 U14812 ( .B1(n12718), .B2(n15059), .A(n12528), .ZN(n12529) );
  OAI21_X1 U14813 ( .B1(n12530), .B2(n15093), .A(n12529), .ZN(P3_U3209) );
  XNOR2_X1 U14814 ( .A(n12531), .B(n12534), .ZN(n12539) );
  INV_X1 U14815 ( .A(n12532), .ZN(n12535) );
  AOI21_X1 U14816 ( .B1(n12535), .B2(n12534), .A(n12533), .ZN(n12722) );
  OAI22_X1 U14817 ( .A1(n12536), .A2(n15046), .B1(n12564), .B2(n15048), .ZN(
        n12537) );
  AOI21_X1 U14818 ( .B1(n12722), .B2(n15031), .A(n12537), .ZN(n12538) );
  OAI21_X1 U14819 ( .B1(n15043), .B2(n12539), .A(n12538), .ZN(n12721) );
  INV_X1 U14820 ( .A(n12721), .ZN(n12546) );
  INV_X1 U14821 ( .A(n12540), .ZN(n12804) );
  AOI22_X1 U14822 ( .A1(n15093), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15053), 
        .B2(n12541), .ZN(n12542) );
  OAI21_X1 U14823 ( .B1(n12804), .B2(n12691), .A(n12542), .ZN(n12543) );
  AOI21_X1 U14824 ( .B1(n12722), .B2(n12544), .A(n12543), .ZN(n12545) );
  OAI21_X1 U14825 ( .B1(n12546), .B2(n15093), .A(n12545), .ZN(P3_U3210) );
  XNOR2_X1 U14826 ( .A(n12547), .B(n12551), .ZN(n12548) );
  OAI222_X1 U14827 ( .A1(n15046), .A2(n12549), .B1(n15048), .B2(n12574), .C1(
        n15043), .C2(n12548), .ZN(n12725) );
  INV_X1 U14828 ( .A(n12725), .ZN(n12556) );
  XOR2_X1 U14829 ( .A(n12551), .B(n12550), .Z(n12726) );
  AOI22_X1 U14830 ( .A1(n15093), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15053), 
        .B2(n12552), .ZN(n12553) );
  OAI21_X1 U14831 ( .B1(n12808), .B2(n12691), .A(n12553), .ZN(n12554) );
  AOI21_X1 U14832 ( .B1(n12726), .B2(n15059), .A(n12554), .ZN(n12555) );
  OAI21_X1 U14833 ( .B1(n12556), .B2(n15093), .A(n12555), .ZN(P3_U3211) );
  XNOR2_X1 U14834 ( .A(n12557), .B(n7307), .ZN(n12730) );
  INV_X1 U14835 ( .A(n12730), .ZN(n12570) );
  INV_X1 U14836 ( .A(n12558), .ZN(n12559) );
  AOI21_X1 U14837 ( .B1(n12561), .B2(n12560), .A(n12559), .ZN(n12562) );
  OAI222_X1 U14838 ( .A1(n15046), .A2(n12564), .B1(n15048), .B2(n12563), .C1(
        n15043), .C2(n12562), .ZN(n12729) );
  INV_X1 U14839 ( .A(n12565), .ZN(n12812) );
  AOI22_X1 U14840 ( .A1(n15093), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15053), 
        .B2(n12566), .ZN(n12567) );
  OAI21_X1 U14841 ( .B1(n12812), .B2(n12691), .A(n12567), .ZN(n12568) );
  AOI21_X1 U14842 ( .B1(n12729), .B2(n15091), .A(n12568), .ZN(n12569) );
  OAI21_X1 U14843 ( .B1(n12570), .B2(n12697), .A(n12569), .ZN(P3_U3212) );
  OAI211_X1 U14844 ( .C1(n12573), .C2(n12572), .A(n12571), .B(n15072), .ZN(
        n12577) );
  OAI22_X1 U14845 ( .A1(n12604), .A2(n15048), .B1(n12574), .B2(n15046), .ZN(
        n12575) );
  INV_X1 U14846 ( .A(n12575), .ZN(n12576) );
  OAI22_X1 U14847 ( .A1(n15091), .A2(n12579), .B1(n12578), .B2(n15083), .ZN(
        n12584) );
  OAI21_X1 U14848 ( .B1(n12582), .B2(n12581), .A(n12580), .ZN(n12734) );
  NOR2_X1 U14849 ( .A1(n12734), .A2(n12697), .ZN(n12583) );
  AOI211_X1 U14850 ( .C1(n14462), .C2(n12815), .A(n12584), .B(n12583), .ZN(
        n12585) );
  OAI21_X1 U14851 ( .B1(n15093), .B2(n12735), .A(n12585), .ZN(P3_U3213) );
  XNOR2_X1 U14852 ( .A(n12586), .B(n7644), .ZN(n12740) );
  INV_X1 U14853 ( .A(n12740), .ZN(n12598) );
  OAI211_X1 U14854 ( .C1(n12588), .C2(n7644), .A(n15072), .B(n12587), .ZN(
        n12592) );
  AOI22_X1 U14855 ( .A1(n15066), .A2(n12590), .B1(n12589), .B2(n15069), .ZN(
        n12591) );
  NAND2_X1 U14856 ( .A1(n12592), .A2(n12591), .ZN(n12739) );
  NOR2_X1 U14857 ( .A1(n12820), .A2(n12691), .ZN(n12596) );
  OAI22_X1 U14858 ( .A1(n15091), .A2(n12594), .B1(n12593), .B2(n15083), .ZN(
        n12595) );
  AOI211_X1 U14859 ( .C1(n12739), .C2(n15091), .A(n12596), .B(n12595), .ZN(
        n12597) );
  OAI21_X1 U14860 ( .B1(n12598), .B2(n12697), .A(n12597), .ZN(P3_U3214) );
  XNOR2_X1 U14861 ( .A(n12599), .B(n12601), .ZN(n12744) );
  INV_X1 U14862 ( .A(n12744), .ZN(n12609) );
  AOI21_X1 U14863 ( .B1(n12601), .B2(n12600), .A(n6563), .ZN(n12602) );
  OAI222_X1 U14864 ( .A1(n15046), .A2(n12604), .B1(n15048), .B2(n12603), .C1(
        n15043), .C2(n12602), .ZN(n12743) );
  AOI22_X1 U14865 ( .A1(n15093), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15053), 
        .B2(n12605), .ZN(n12606) );
  OAI21_X1 U14866 ( .B1(n12824), .B2(n12691), .A(n12606), .ZN(n12607) );
  AOI21_X1 U14867 ( .B1(n12743), .B2(n15091), .A(n12607), .ZN(n12608) );
  OAI21_X1 U14868 ( .B1(n12697), .B2(n12609), .A(n12608), .ZN(P3_U3215) );
  XNOR2_X1 U14869 ( .A(n12611), .B(n12610), .ZN(n12748) );
  INV_X1 U14870 ( .A(n12748), .ZN(n12624) );
  OAI211_X1 U14871 ( .C1(n12614), .C2(n12613), .A(n12612), .B(n15072), .ZN(
        n12617) );
  OR2_X1 U14872 ( .A1(n12615), .A2(n15048), .ZN(n12616) );
  OAI211_X1 U14873 ( .C1(n12618), .C2(n15046), .A(n12617), .B(n12616), .ZN(
        n12747) );
  INV_X1 U14874 ( .A(n12619), .ZN(n12620) );
  AOI22_X1 U14875 ( .A1(n15093), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15053), 
        .B2(n12620), .ZN(n12621) );
  OAI21_X1 U14876 ( .B1(n12828), .B2(n12691), .A(n12621), .ZN(n12622) );
  AOI21_X1 U14877 ( .B1(n12747), .B2(n15091), .A(n12622), .ZN(n12623) );
  OAI21_X1 U14878 ( .B1(n12624), .B2(n12697), .A(n12623), .ZN(P3_U3216) );
  OAI211_X1 U14879 ( .C1(n12627), .C2(n12626), .A(n12625), .B(n15072), .ZN(
        n12630) );
  AOI22_X1 U14880 ( .A1(n15069), .A2(n12659), .B1(n12628), .B2(n15066), .ZN(
        n12629) );
  AND2_X1 U14881 ( .A1(n12630), .A2(n12629), .ZN(n12752) );
  OR2_X1 U14882 ( .A1(n12632), .A2(n12631), .ZN(n12633) );
  NAND2_X1 U14883 ( .A1(n12634), .A2(n12633), .ZN(n12751) );
  NOR2_X1 U14884 ( .A1(n12635), .A2(n12691), .ZN(n12639) );
  OAI22_X1 U14885 ( .A1(n15091), .A2(n12637), .B1(n12636), .B2(n15083), .ZN(
        n12638) );
  AOI211_X1 U14886 ( .C1(n12751), .C2(n15059), .A(n12639), .B(n12638), .ZN(
        n12640) );
  OAI21_X1 U14887 ( .B1(n15093), .B2(n12752), .A(n12640), .ZN(P3_U3217) );
  XNOR2_X1 U14888 ( .A(n12642), .B(n12641), .ZN(n12758) );
  INV_X1 U14889 ( .A(n12758), .ZN(n12654) );
  OAI211_X1 U14890 ( .C1(n12645), .C2(n12644), .A(n12643), .B(n15072), .ZN(
        n12648) );
  AOI22_X1 U14891 ( .A1(n12646), .A2(n15066), .B1(n15069), .B2(n12673), .ZN(
        n12647) );
  NAND2_X1 U14892 ( .A1(n12648), .A2(n12647), .ZN(n12757) );
  INV_X1 U14893 ( .A(n12649), .ZN(n12650) );
  AOI22_X1 U14894 ( .A1(n15093), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15053), 
        .B2(n12650), .ZN(n12651) );
  OAI21_X1 U14895 ( .B1(n12837), .B2(n12691), .A(n12651), .ZN(n12652) );
  AOI21_X1 U14896 ( .B1(n12757), .B2(n15091), .A(n12652), .ZN(n12653) );
  OAI21_X1 U14897 ( .B1(n12654), .B2(n12697), .A(n12653), .ZN(P3_U3218) );
  XNOR2_X1 U14898 ( .A(n12655), .B(n12657), .ZN(n12762) );
  INV_X1 U14899 ( .A(n12762), .ZN(n12667) );
  OAI211_X1 U14900 ( .C1(n12658), .C2(n12657), .A(n12656), .B(n15072), .ZN(
        n12661) );
  AOI22_X1 U14901 ( .A1(n15069), .A2(n12687), .B1(n12659), .B2(n15066), .ZN(
        n12660) );
  NAND2_X1 U14902 ( .A1(n12661), .A2(n12660), .ZN(n12761) );
  INV_X1 U14903 ( .A(n12662), .ZN(n12663) );
  AOI22_X1 U14904 ( .A1(n15093), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15053), 
        .B2(n12663), .ZN(n12664) );
  OAI21_X1 U14905 ( .B1(n12691), .B2(n12841), .A(n12664), .ZN(n12665) );
  AOI21_X1 U14906 ( .B1(n12761), .B2(n15091), .A(n12665), .ZN(n12666) );
  OAI21_X1 U14907 ( .B1(n12667), .B2(n12697), .A(n12666), .ZN(P3_U3219) );
  XNOR2_X1 U14908 ( .A(n12669), .B(n12668), .ZN(n12766) );
  INV_X1 U14909 ( .A(n12766), .ZN(n12680) );
  OAI211_X1 U14910 ( .C1(n12672), .C2(n12671), .A(n12670), .B(n15072), .ZN(
        n12675) );
  AOI22_X1 U14911 ( .A1(n15069), .A2(n14468), .B1(n12673), .B2(n15066), .ZN(
        n12674) );
  NAND2_X1 U14912 ( .A1(n12675), .A2(n12674), .ZN(n12765) );
  NOR2_X1 U14913 ( .A1(n12691), .A2(n12845), .ZN(n12678) );
  OAI22_X1 U14914 ( .A1(n15091), .A2(n7882), .B1(n12676), .B2(n15083), .ZN(
        n12677) );
  AOI211_X1 U14915 ( .C1(n12765), .C2(n15091), .A(n12678), .B(n12677), .ZN(
        n12679) );
  OAI21_X1 U14916 ( .B1(n12680), .B2(n12697), .A(n12679), .ZN(P3_U3220) );
  OAI21_X1 U14917 ( .B1(n12682), .B2(n12683), .A(n12681), .ZN(n14482) );
  INV_X1 U14918 ( .A(n14482), .ZN(n12698) );
  NAND2_X1 U14919 ( .A1(n12684), .A2(n12683), .ZN(n12685) );
  NAND3_X1 U14920 ( .A1(n12686), .A2(n15072), .A3(n12685), .ZN(n12690) );
  AOI22_X1 U14921 ( .A1(n12688), .A2(n15069), .B1(n15066), .B2(n12687), .ZN(
        n12689) );
  NAND2_X1 U14922 ( .A1(n12690), .A2(n12689), .ZN(n14480) );
  NOR2_X1 U14923 ( .A1(n12691), .A2(n14479), .ZN(n12695) );
  OAI22_X1 U14924 ( .A1(n15091), .A2(n12693), .B1(n12692), .B2(n15083), .ZN(
        n12694) );
  AOI211_X1 U14925 ( .C1(n14480), .C2(n15091), .A(n12695), .B(n12694), .ZN(
        n12696) );
  OAI21_X1 U14926 ( .B1(n12698), .B2(n12697), .A(n12696), .ZN(P3_U3221) );
  INV_X1 U14927 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n12699) );
  MUX2_X1 U14928 ( .A(n12699), .B(n12783), .S(n15149), .Z(n12700) );
  OAI21_X1 U14929 ( .B1(n12785), .B2(n12769), .A(n12700), .ZN(P3_U3490) );
  MUX2_X1 U14930 ( .A(n12702), .B(n12701), .S(n15149), .Z(n12703) );
  OAI21_X1 U14931 ( .B1(n12704), .B2(n12769), .A(n12703), .ZN(P3_U3487) );
  INV_X1 U14932 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12707) );
  AOI21_X1 U14933 ( .B1(n15132), .B2(n12706), .A(n12705), .ZN(n12786) );
  OAI21_X1 U14934 ( .B1(n12789), .B2(n12769), .A(n12708), .ZN(P3_U3486) );
  AOI21_X1 U14935 ( .B1(n15132), .B2(n12710), .A(n12709), .ZN(n12790) );
  MUX2_X1 U14936 ( .A(n12711), .B(n12790), .S(n15149), .Z(n12712) );
  OAI21_X1 U14937 ( .B1(n12793), .B2(n12769), .A(n12712), .ZN(P3_U3485) );
  INV_X1 U14938 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12715) );
  AOI21_X1 U14939 ( .B1(n15132), .B2(n12714), .A(n12713), .ZN(n12794) );
  MUX2_X1 U14940 ( .A(n12715), .B(n12794), .S(n15149), .Z(n12716) );
  OAI21_X1 U14941 ( .B1(n7400), .B2(n12769), .A(n12716), .ZN(P3_U3484) );
  INV_X1 U14942 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12719) );
  AOI21_X1 U14943 ( .B1(n15102), .B2(n12718), .A(n12717), .ZN(n12797) );
  MUX2_X1 U14944 ( .A(n12719), .B(n12797), .S(n15149), .Z(n12720) );
  OAI21_X1 U14945 ( .B1(n12800), .B2(n12769), .A(n12720), .ZN(P3_U3483) );
  INV_X1 U14946 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12723) );
  AOI21_X1 U14947 ( .B1(n15132), .B2(n12722), .A(n12721), .ZN(n12801) );
  MUX2_X1 U14948 ( .A(n12723), .B(n12801), .S(n15149), .Z(n12724) );
  OAI21_X1 U14949 ( .B1(n12804), .B2(n12769), .A(n12724), .ZN(P3_U3482) );
  INV_X1 U14950 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12727) );
  AOI21_X1 U14951 ( .B1(n15102), .B2(n12726), .A(n12725), .ZN(n12805) );
  MUX2_X1 U14952 ( .A(n12727), .B(n12805), .S(n15149), .Z(n12728) );
  OAI21_X1 U14953 ( .B1(n12808), .B2(n12769), .A(n12728), .ZN(P3_U3481) );
  AOI21_X1 U14954 ( .B1(n15102), .B2(n12730), .A(n12729), .ZN(n12809) );
  MUX2_X1 U14955 ( .A(n12731), .B(n12809), .S(n15149), .Z(n12732) );
  OAI21_X1 U14956 ( .B1(n12812), .B2(n12769), .A(n12732), .ZN(P3_U3480) );
  INV_X1 U14957 ( .A(n12769), .ZN(n12755) );
  INV_X1 U14958 ( .A(n15102), .ZN(n12733) );
  OR2_X1 U14959 ( .A1(n12734), .A2(n12733), .ZN(n12736) );
  NAND2_X1 U14960 ( .A1(n12736), .A2(n12735), .ZN(n12813) );
  MUX2_X1 U14961 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12813), .S(n15149), .Z(
        n12737) );
  AOI21_X1 U14962 ( .B1(n12755), .B2(n12815), .A(n12737), .ZN(n12738) );
  INV_X1 U14963 ( .A(n12738), .ZN(P3_U3479) );
  AOI21_X1 U14964 ( .B1(n15102), .B2(n12740), .A(n12739), .ZN(n12817) );
  MUX2_X1 U14965 ( .A(n12741), .B(n12817), .S(n15149), .Z(n12742) );
  OAI21_X1 U14966 ( .B1(n12820), .B2(n12769), .A(n12742), .ZN(P3_U3478) );
  AOI21_X1 U14967 ( .B1(n12744), .B2(n15102), .A(n12743), .ZN(n12821) );
  MUX2_X1 U14968 ( .A(n12745), .B(n12821), .S(n15149), .Z(n12746) );
  OAI21_X1 U14969 ( .B1(n12824), .B2(n12769), .A(n12746), .ZN(P3_U3477) );
  AOI21_X1 U14970 ( .B1(n12748), .B2(n15102), .A(n12747), .ZN(n12825) );
  MUX2_X1 U14971 ( .A(n12749), .B(n12825), .S(n15149), .Z(n12750) );
  OAI21_X1 U14972 ( .B1(n12769), .B2(n12828), .A(n12750), .ZN(P3_U3476) );
  NAND2_X1 U14973 ( .A1(n12751), .A2(n15102), .ZN(n12753) );
  NAND2_X1 U14974 ( .A1(n12753), .A2(n12752), .ZN(n12829) );
  MUX2_X1 U14975 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12829), .S(n15149), .Z(
        n12754) );
  AOI21_X1 U14976 ( .B1(n12755), .B2(n12831), .A(n12754), .ZN(n12756) );
  INV_X1 U14977 ( .A(n12756), .ZN(P3_U3475) );
  AOI21_X1 U14978 ( .B1(n12758), .B2(n15102), .A(n12757), .ZN(n12834) );
  MUX2_X1 U14979 ( .A(n12759), .B(n12834), .S(n15149), .Z(n12760) );
  OAI21_X1 U14980 ( .B1(n12769), .B2(n12837), .A(n12760), .ZN(P3_U3474) );
  AOI21_X1 U14981 ( .B1(n12762), .B2(n15102), .A(n12761), .ZN(n12838) );
  MUX2_X1 U14982 ( .A(n12763), .B(n12838), .S(n15149), .Z(n12764) );
  OAI21_X1 U14983 ( .B1(n12769), .B2(n12841), .A(n12764), .ZN(P3_U3473) );
  AOI21_X1 U14984 ( .B1(n12766), .B2(n15102), .A(n12765), .ZN(n12842) );
  MUX2_X1 U14985 ( .A(n12767), .B(n12842), .S(n15149), .Z(n12768) );
  OAI21_X1 U14986 ( .B1(n12769), .B2(n12845), .A(n12768), .ZN(P3_U3472) );
  XNOR2_X1 U14987 ( .A(n10546), .B(n12770), .ZN(n12776) );
  NAND2_X1 U14988 ( .A1(n6905), .A2(n15069), .ZN(n12774) );
  NAND2_X1 U14989 ( .A1(n12772), .A2(n15066), .ZN(n12773) );
  NAND2_X1 U14990 ( .A1(n12774), .A2(n12773), .ZN(n12775) );
  AOI21_X1 U14991 ( .B1(n12776), .B2(n15072), .A(n12775), .ZN(n12779) );
  XNOR2_X1 U14992 ( .A(n10546), .B(n12777), .ZN(n15089) );
  NAND2_X1 U14993 ( .A1(n15089), .A2(n15031), .ZN(n12778) );
  AND2_X1 U14994 ( .A1(n12779), .A2(n12778), .ZN(n15086) );
  NOR2_X1 U14995 ( .A1(n12780), .A2(n15111), .ZN(n15081) );
  AOI21_X1 U14996 ( .B1(n15089), .B2(n15132), .A(n15081), .ZN(n12781) );
  AND2_X1 U14997 ( .A1(n15086), .A2(n12781), .ZN(n15094) );
  INV_X1 U14998 ( .A(n15094), .ZN(n12782) );
  MUX2_X1 U14999 ( .A(n12782), .B(P3_REG1_REG_1__SCAN_IN), .S(n15147), .Z(
        P3_U3460) );
  MUX2_X1 U15000 ( .A(n11607), .B(n12783), .S(n15136), .Z(n12784) );
  OAI21_X1 U15001 ( .B1(n12785), .B2(n12846), .A(n12784), .ZN(P3_U3458) );
  INV_X1 U15002 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12787) );
  OAI21_X1 U15003 ( .B1(n12789), .B2(n12846), .A(n12788), .ZN(P3_U3454) );
  INV_X1 U15004 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12791) );
  MUX2_X1 U15005 ( .A(n12791), .B(n12790), .S(n15136), .Z(n12792) );
  OAI21_X1 U15006 ( .B1(n12793), .B2(n12846), .A(n12792), .ZN(P3_U3453) );
  INV_X1 U15007 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12795) );
  MUX2_X1 U15008 ( .A(n12795), .B(n12794), .S(n15136), .Z(n12796) );
  OAI21_X1 U15009 ( .B1(n7400), .B2(n12846), .A(n12796), .ZN(P3_U3452) );
  INV_X1 U15010 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12798) );
  MUX2_X1 U15011 ( .A(n12798), .B(n12797), .S(n15136), .Z(n12799) );
  OAI21_X1 U15012 ( .B1(n12800), .B2(n12846), .A(n12799), .ZN(P3_U3451) );
  INV_X1 U15013 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12802) );
  MUX2_X1 U15014 ( .A(n12802), .B(n12801), .S(n15136), .Z(n12803) );
  OAI21_X1 U15015 ( .B1(n12804), .B2(n12846), .A(n12803), .ZN(P3_U3450) );
  INV_X1 U15016 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12806) );
  MUX2_X1 U15017 ( .A(n12806), .B(n12805), .S(n15136), .Z(n12807) );
  OAI21_X1 U15018 ( .B1(n12808), .B2(n12846), .A(n12807), .ZN(P3_U3449) );
  MUX2_X1 U15019 ( .A(n12810), .B(n12809), .S(n15136), .Z(n12811) );
  OAI21_X1 U15020 ( .B1(n12812), .B2(n12846), .A(n12811), .ZN(P3_U3448) );
  INV_X1 U15021 ( .A(n12846), .ZN(n12832) );
  MUX2_X1 U15022 ( .A(n12813), .B(P3_REG0_REG_20__SCAN_IN), .S(n15137), .Z(
        n12814) );
  AOI21_X1 U15023 ( .B1(n12832), .B2(n12815), .A(n12814), .ZN(n12816) );
  INV_X1 U15024 ( .A(n12816), .ZN(P3_U3447) );
  INV_X1 U15025 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12818) );
  MUX2_X1 U15026 ( .A(n12818), .B(n12817), .S(n15136), .Z(n12819) );
  OAI21_X1 U15027 ( .B1(n12820), .B2(n12846), .A(n12819), .ZN(P3_U3446) );
  MUX2_X1 U15028 ( .A(n12822), .B(n12821), .S(n15136), .Z(n12823) );
  OAI21_X1 U15029 ( .B1(n12824), .B2(n12846), .A(n12823), .ZN(P3_U3444) );
  INV_X1 U15030 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12826) );
  MUX2_X1 U15031 ( .A(n12826), .B(n12825), .S(n15136), .Z(n12827) );
  OAI21_X1 U15032 ( .B1(n12846), .B2(n12828), .A(n12827), .ZN(P3_U3441) );
  MUX2_X1 U15033 ( .A(n12829), .B(P3_REG0_REG_16__SCAN_IN), .S(n15137), .Z(
        n12830) );
  AOI21_X1 U15034 ( .B1(n12832), .B2(n12831), .A(n12830), .ZN(n12833) );
  INV_X1 U15035 ( .A(n12833), .ZN(P3_U3438) );
  INV_X1 U15036 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12835) );
  MUX2_X1 U15037 ( .A(n12835), .B(n12834), .S(n15136), .Z(n12836) );
  OAI21_X1 U15038 ( .B1(n12846), .B2(n12837), .A(n12836), .ZN(P3_U3435) );
  MUX2_X1 U15039 ( .A(n12839), .B(n12838), .S(n15136), .Z(n12840) );
  OAI21_X1 U15040 ( .B1(n12846), .B2(n12841), .A(n12840), .ZN(P3_U3432) );
  INV_X1 U15041 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12843) );
  MUX2_X1 U15042 ( .A(n12843), .B(n12842), .S(n15136), .Z(n12844) );
  OAI21_X1 U15043 ( .B1(n12846), .B2(n12845), .A(n12844), .ZN(P3_U3429) );
  MUX2_X1 U15044 ( .A(n12847), .B(P3_D_REG_1__SCAN_IN), .S(n12848), .Z(
        P3_U3377) );
  MUX2_X1 U15045 ( .A(n12849), .B(P3_D_REG_0__SCAN_IN), .S(n12848), .Z(
        P3_U3376) );
  NAND3_X1 U15046 ( .A1(n12851), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12853) );
  OAI22_X1 U15047 ( .A1(n12850), .A2(n12853), .B1(n12852), .B2(n14376), .ZN(
        n12854) );
  AOI21_X1 U15048 ( .B1(n12855), .B2(n14388), .A(n12854), .ZN(n12856) );
  INV_X1 U15049 ( .A(n12856), .ZN(P3_U3264) );
  INV_X1 U15050 ( .A(n12857), .ZN(n12858) );
  OAI222_X1 U15051 ( .A1(n7678), .A2(P3_U3151), .B1(n14376), .B2(n12859), .C1(
        n14378), .C2(n12858), .ZN(P3_U3265) );
  INV_X1 U15052 ( .A(n12860), .ZN(n12861) );
  OAI222_X1 U15053 ( .A1(n14376), .A2(n12863), .B1(P3_U3151), .B2(n12862), 
        .C1(n14378), .C2(n12861), .ZN(P3_U3266) );
  NAND2_X1 U15054 ( .A1(n13259), .A2(n12864), .ZN(n12914) );
  INV_X1 U15055 ( .A(n12914), .ZN(n12917) );
  XNOR2_X1 U15056 ( .A(n13477), .B(n12966), .ZN(n12916) );
  NAND2_X1 U15057 ( .A1(n13301), .A2(n9733), .ZN(n12950) );
  INV_X1 U15058 ( .A(n12950), .ZN(n12907) );
  XNOR2_X1 U15059 ( .A(n13492), .B(n12900), .ZN(n12946) );
  INV_X1 U15060 ( .A(n12946), .ZN(n12906) );
  XNOR2_X1 U15061 ( .A(n13434), .B(n12966), .ZN(n12867) );
  NAND2_X1 U15062 ( .A1(n13442), .A2(n12864), .ZN(n12868) );
  XNOR2_X1 U15063 ( .A(n12867), .B(n12868), .ZN(n12937) );
  INV_X1 U15064 ( .A(n12867), .ZN(n12869) );
  NAND2_X1 U15065 ( .A1(n12869), .A2(n12868), .ZN(n12870) );
  XNOR2_X1 U15066 ( .A(n13538), .B(n12966), .ZN(n12873) );
  AND2_X1 U15067 ( .A1(n13104), .A2(n9733), .ZN(n12871) );
  INV_X1 U15068 ( .A(n12872), .ZN(n12874) );
  NAND2_X1 U15069 ( .A1(n12874), .A2(n12873), .ZN(n12875) );
  XNOR2_X1 U15070 ( .A(n13533), .B(n12900), .ZN(n13007) );
  NAND2_X1 U15071 ( .A1(n13103), .A2(n9733), .ZN(n12876) );
  XNOR2_X1 U15072 ( .A(n13007), .B(n12876), .ZN(n12995) );
  NAND2_X1 U15073 ( .A1(n13007), .A2(n12876), .ZN(n12877) );
  XNOR2_X1 U15074 ( .A(n13527), .B(n12966), .ZN(n12878) );
  NAND2_X1 U15075 ( .A1(n13102), .A2(n9733), .ZN(n12879) );
  XNOR2_X1 U15076 ( .A(n12878), .B(n12879), .ZN(n13005) );
  INV_X1 U15077 ( .A(n12878), .ZN(n12880) );
  NAND2_X1 U15078 ( .A1(n12880), .A2(n12879), .ZN(n12881) );
  XNOR2_X1 U15079 ( .A(n13522), .B(n12966), .ZN(n12882) );
  AND2_X1 U15080 ( .A1(n13101), .A2(n9733), .ZN(n12883) );
  NAND2_X1 U15081 ( .A1(n12882), .A2(n12883), .ZN(n12886) );
  INV_X1 U15082 ( .A(n12882), .ZN(n12957) );
  INV_X1 U15083 ( .A(n12883), .ZN(n12884) );
  NAND2_X1 U15084 ( .A1(n12957), .A2(n12884), .ZN(n12885) );
  NAND2_X1 U15085 ( .A1(n12886), .A2(n12885), .ZN(n13061) );
  XNOR2_X1 U15086 ( .A(n13516), .B(n12966), .ZN(n12888) );
  NAND2_X1 U15087 ( .A1(n13100), .A2(n9733), .ZN(n12889) );
  XNOR2_X1 U15088 ( .A(n12888), .B(n12889), .ZN(n12958) );
  AND2_X1 U15089 ( .A1(n12958), .A2(n12886), .ZN(n12887) );
  INV_X1 U15090 ( .A(n12888), .ZN(n13029) );
  NAND2_X1 U15091 ( .A1(n13029), .A2(n12889), .ZN(n12890) );
  XNOR2_X1 U15092 ( .A(n13511), .B(n12966), .ZN(n12891) );
  NAND2_X1 U15093 ( .A1(n13099), .A2(n9733), .ZN(n12892) );
  XNOR2_X1 U15094 ( .A(n12891), .B(n12892), .ZN(n13028) );
  INV_X1 U15095 ( .A(n12891), .ZN(n12893) );
  NAND2_X1 U15096 ( .A1(n12893), .A2(n12892), .ZN(n12894) );
  XNOR2_X1 U15097 ( .A(n13325), .B(n12900), .ZN(n12895) );
  NAND2_X1 U15098 ( .A1(n13300), .A2(n9733), .ZN(n12896) );
  XNOR2_X1 U15099 ( .A(n12895), .B(n12896), .ZN(n12974) );
  INV_X1 U15100 ( .A(n12895), .ZN(n12898) );
  INV_X1 U15101 ( .A(n12896), .ZN(n12897) );
  NAND2_X1 U15102 ( .A1(n12898), .A2(n12897), .ZN(n12899) );
  XNOR2_X1 U15103 ( .A(n13498), .B(n12900), .ZN(n12902) );
  AND2_X1 U15104 ( .A1(n13098), .A2(n9733), .ZN(n12901) );
  INV_X1 U15105 ( .A(n12902), .ZN(n12903) );
  NAND2_X1 U15106 ( .A1(n12904), .A2(n12903), .ZN(n12945) );
  XNOR2_X1 U15107 ( .A(n13487), .B(n12966), .ZN(n12984) );
  AND2_X1 U15108 ( .A1(n13258), .A2(n9733), .ZN(n12908) );
  NAND2_X1 U15109 ( .A1(n12984), .A2(n12908), .ZN(n12909) );
  OAI21_X1 U15110 ( .B1(n12984), .B2(n12908), .A(n12909), .ZN(n13015) );
  XNOR2_X1 U15111 ( .A(n13482), .B(n12966), .ZN(n12910) );
  AND2_X1 U15112 ( .A1(n13240), .A2(n9733), .ZN(n12911) );
  NAND2_X1 U15113 ( .A1(n12910), .A2(n12911), .ZN(n12915) );
  INV_X1 U15114 ( .A(n12910), .ZN(n13076) );
  INV_X1 U15115 ( .A(n12911), .ZN(n12912) );
  NAND2_X1 U15116 ( .A1(n13076), .A2(n12912), .ZN(n12913) );
  AND2_X1 U15117 ( .A1(n12915), .A2(n12913), .ZN(n12985) );
  XNOR2_X1 U15118 ( .A(n12916), .B(n12914), .ZN(n13077) );
  XNOR2_X1 U15119 ( .A(n13472), .B(n12966), .ZN(n12919) );
  AND2_X1 U15120 ( .A1(n13241), .A2(n9733), .ZN(n12918) );
  NAND2_X1 U15121 ( .A1(n12919), .A2(n12918), .ZN(n12963) );
  OAI21_X1 U15122 ( .B1(n12919), .B2(n12918), .A(n12963), .ZN(n12920) );
  OAI22_X1 U15123 ( .A1(n12923), .A2(n13039), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12922), .ZN(n12924) );
  AOI21_X1 U15124 ( .B1(n13231), .B2(n13070), .A(n12924), .ZN(n12925) );
  OAI21_X1 U15125 ( .B1(n12926), .B2(n13072), .A(n12925), .ZN(n12927) );
  AOI22_X1 U15126 ( .A1(n13078), .A2(n13105), .B1(n13046), .B2(n13104), .ZN(
        n12933) );
  OAI211_X1 U15127 ( .C1(n13430), .C2(n13091), .A(n12933), .B(n12932), .ZN(
        n12940) );
  NOR3_X1 U15128 ( .A1(n12934), .A2(n13421), .A3(n13075), .ZN(n12935) );
  AOI21_X1 U15129 ( .B1(n12936), .B2(n13085), .A(n12935), .ZN(n12938) );
  NOR2_X1 U15130 ( .A1(n12938), .A2(n12937), .ZN(n12939) );
  AOI211_X1 U15131 ( .C1(n13434), .C2(n13093), .A(n12940), .B(n12939), .ZN(
        n12941) );
  OAI21_X1 U15132 ( .B1(n12942), .B2(n13082), .A(n12941), .ZN(P2_U3187) );
  AOI22_X1 U15133 ( .A1(n13258), .A2(n13441), .B1(n13444), .B2(n13098), .ZN(
        n13284) );
  INV_X1 U15134 ( .A(n12943), .ZN(n13288) );
  AOI22_X1 U15135 ( .A1(n13288), .A2(n13070), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12944) );
  OAI21_X1 U15136 ( .B1(n13284), .B2(n12996), .A(n12944), .ZN(n12949) );
  NAND2_X1 U15137 ( .A1(n13036), .A2(n12945), .ZN(n12947) );
  XNOR2_X1 U15138 ( .A(n12947), .B(n12946), .ZN(n12951) );
  NOR3_X1 U15139 ( .A1(n12951), .A2(n13040), .A3(n13075), .ZN(n12948) );
  NAND3_X1 U15140 ( .A1(n12951), .A2(n13085), .A3(n12950), .ZN(n12952) );
  NAND2_X1 U15141 ( .A1(n12953), .A2(n12952), .ZN(P2_U3188) );
  OAI21_X1 U15142 ( .B1(n12958), .B2(n13059), .A(n13031), .ZN(n12954) );
  NAND2_X1 U15143 ( .A1(n12954), .A2(n13085), .ZN(n12962) );
  NAND2_X1 U15144 ( .A1(n13046), .A2(n13099), .ZN(n12955) );
  NAND2_X1 U15145 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13191)
         );
  OAI211_X1 U15146 ( .C1(n13091), .C2(n13352), .A(n12955), .B(n13191), .ZN(
        n12956) );
  AOI21_X1 U15147 ( .B1(n13516), .B2(n13093), .A(n12956), .ZN(n12961) );
  NOR3_X1 U15148 ( .A1(n12958), .A2(n12957), .A3(n13075), .ZN(n12959) );
  OAI21_X1 U15149 ( .B1(n12959), .B2(n13078), .A(n13101), .ZN(n12960) );
  NAND3_X1 U15150 ( .A1(n12962), .A2(n12961), .A3(n12960), .ZN(P2_U3191) );
  INV_X1 U15151 ( .A(n12963), .ZN(n12964) );
  NAND2_X1 U15152 ( .A1(n13227), .A2(n9733), .ZN(n12965) );
  XOR2_X1 U15153 ( .A(n12966), .B(n12965), .Z(n12967) );
  XNOR2_X1 U15154 ( .A(n13465), .B(n12967), .ZN(n12968) );
  OAI22_X1 U15155 ( .A1(n13218), .A2(n13091), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12969), .ZN(n12970) );
  AOI21_X1 U15156 ( .B1(n13046), .B2(n13209), .A(n12970), .ZN(n12971) );
  OAI21_X1 U15157 ( .B1(n13073), .B2(n13039), .A(n12971), .ZN(n12972) );
  AOI21_X1 U15158 ( .B1(n13465), .B2(n13093), .A(n12972), .ZN(n12973) );
  AOI21_X1 U15159 ( .B1(n12975), .B2(n12974), .A(n13082), .ZN(n12977) );
  NAND2_X1 U15160 ( .A1(n12977), .A2(n12976), .ZN(n12983) );
  INV_X1 U15161 ( .A(n13322), .ZN(n12981) );
  AND2_X1 U15162 ( .A1(n13099), .A2(n13444), .ZN(n12978) );
  AOI21_X1 U15163 ( .B1(n13098), .B2(n13441), .A(n12978), .ZN(n13316) );
  OAI22_X1 U15164 ( .A1(n13316), .A2(n12996), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12979), .ZN(n12980) );
  AOI21_X1 U15165 ( .B1(n12981), .B2(n13070), .A(n12980), .ZN(n12982) );
  OAI211_X1 U15166 ( .C1(n7261), .C2(n13023), .A(n12983), .B(n12982), .ZN(
        P2_U3195) );
  NAND3_X1 U15167 ( .A1(n12984), .A2(n13084), .A3(n13258), .ZN(n12988) );
  OAI21_X1 U15168 ( .B1(n6477), .B2(n12985), .A(n13085), .ZN(n12987) );
  INV_X1 U15169 ( .A(n13067), .ZN(n12986) );
  AOI21_X1 U15170 ( .B1(n12988), .B2(n12987), .A(n12986), .ZN(n12992) );
  AOI22_X1 U15171 ( .A1(n13264), .A2(n13070), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12990) );
  AOI22_X1 U15172 ( .A1(n13259), .A2(n13046), .B1(n13078), .B2(n13258), .ZN(
        n12989) );
  OAI211_X1 U15173 ( .C1(n7255), .C2(n13023), .A(n12990), .B(n12989), .ZN(
        n12991) );
  OR2_X1 U15174 ( .A1(n12992), .A2(n12991), .ZN(P2_U3197) );
  INV_X1 U15175 ( .A(n13010), .ZN(n12993) );
  AOI21_X1 U15176 ( .B1(n12995), .B2(n12994), .A(n12993), .ZN(n13000) );
  NOR2_X1 U15177 ( .A1(n13091), .A2(n13400), .ZN(n12998) );
  AOI22_X1 U15178 ( .A1(n13102), .A2(n13441), .B1(n13104), .B2(n13444), .ZN(
        n13396) );
  OAI22_X1 U15179 ( .A1(n12996), .A2(n13396), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15197), .ZN(n12997) );
  AOI211_X1 U15180 ( .C1(n13533), .C2(n13093), .A(n12998), .B(n12997), .ZN(
        n12999) );
  OAI21_X1 U15181 ( .B1(n13000), .B2(n13082), .A(n12999), .ZN(P2_U3198) );
  NAND2_X1 U15182 ( .A1(n13101), .A2(n13441), .ZN(n13002) );
  NAND2_X1 U15183 ( .A1(n13103), .A2(n13444), .ZN(n13001) );
  NAND2_X1 U15184 ( .A1(n13002), .A2(n13001), .ZN(n13374) );
  AOI22_X1 U15185 ( .A1(n13089), .A2(n13374), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13003) );
  OAI21_X1 U15186 ( .B1(n13379), .B2(n13091), .A(n13003), .ZN(n13004) );
  AOI21_X1 U15187 ( .B1(n13527), .B2(n13093), .A(n13004), .ZN(n13012) );
  INV_X1 U15188 ( .A(n13005), .ZN(n13009) );
  OAI22_X1 U15189 ( .A1(n13007), .A2(n13082), .B1(n13006), .B2(n13075), .ZN(
        n13008) );
  NAND3_X1 U15190 ( .A1(n13010), .A2(n13009), .A3(n13008), .ZN(n13011) );
  OAI211_X1 U15191 ( .C1(n13013), .C2(n13082), .A(n13012), .B(n13011), .ZN(
        P2_U3200) );
  AOI211_X1 U15192 ( .C1(n13015), .C2(n13014), .A(n13082), .B(n6477), .ZN(
        n13016) );
  INV_X1 U15193 ( .A(n13016), .ZN(n13022) );
  NAND2_X1 U15194 ( .A1(n13240), .A2(n13441), .ZN(n13018) );
  NAND2_X1 U15195 ( .A1(n13301), .A2(n13444), .ZN(n13017) );
  NAND2_X1 U15196 ( .A1(n13018), .A2(n13017), .ZN(n13271) );
  OAI22_X1 U15197 ( .A1(n13275), .A2(n13091), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13019), .ZN(n13020) );
  AOI21_X1 U15198 ( .B1(n13271), .B2(n13089), .A(n13020), .ZN(n13021) );
  OAI211_X1 U15199 ( .C1(n6888), .C2(n13023), .A(n13022), .B(n13021), .ZN(
        P2_U3201) );
  INV_X1 U15200 ( .A(n13340), .ZN(n13025) );
  OAI22_X1 U15201 ( .A1(n13091), .A2(n13025), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13024), .ZN(n13027) );
  OAI22_X1 U15202 ( .A1(n13072), .A2(n13336), .B1(n13337), .B2(n13039), .ZN(
        n13026) );
  AOI211_X1 U15203 ( .C1(n13511), .C2(n13093), .A(n13027), .B(n13026), .ZN(
        n13033) );
  OAI22_X1 U15204 ( .A1(n13029), .A2(n13082), .B1(n13337), .B2(n13075), .ZN(
        n13030) );
  NAND3_X1 U15205 ( .A1(n13031), .A2(n6640), .A3(n13030), .ZN(n13032) );
  OAI211_X1 U15206 ( .C1(n13034), .C2(n13082), .A(n13033), .B(n13032), .ZN(
        P2_U3205) );
  AOI22_X1 U15207 ( .A1(n13035), .A2(n13085), .B1(n13084), .B2(n13098), .ZN(
        n13045) );
  INV_X1 U15208 ( .A(n13036), .ZN(n13044) );
  INV_X1 U15209 ( .A(n13306), .ZN(n13038) );
  OAI22_X1 U15210 ( .A1(n13038), .A2(n13091), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13037), .ZN(n13042) );
  OAI22_X1 U15211 ( .A1(n13040), .A2(n13072), .B1(n13336), .B2(n13039), .ZN(
        n13041) );
  AOI211_X1 U15212 ( .C1(n13498), .C2(n13093), .A(n13042), .B(n13041), .ZN(
        n13043) );
  OAI21_X1 U15213 ( .B1(n13045), .B2(n13044), .A(n13043), .ZN(P2_U3207) );
  AOI22_X1 U15214 ( .A1(n13078), .A2(n13116), .B1(n13046), .B2(n13114), .ZN(
        n13055) );
  AOI22_X1 U15215 ( .A1(n13048), .A2(n13093), .B1(n13047), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n13054) );
  OAI21_X1 U15216 ( .B1(n13051), .B2(n13050), .A(n13049), .ZN(n13052) );
  NAND2_X1 U15217 ( .A1(n13052), .A2(n13085), .ZN(n13053) );
  NAND3_X1 U15218 ( .A1(n13055), .A2(n13054), .A3(n13053), .ZN(P2_U3209) );
  NAND2_X1 U15219 ( .A1(n13100), .A2(n13441), .ZN(n13057) );
  NAND2_X1 U15220 ( .A1(n13102), .A2(n13444), .ZN(n13056) );
  NAND2_X1 U15221 ( .A1(n13057), .A2(n13056), .ZN(n13360) );
  AOI22_X1 U15222 ( .A1(n13089), .A2(n13360), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13058) );
  OAI21_X1 U15223 ( .B1(n13366), .B2(n13091), .A(n13058), .ZN(n13064) );
  INV_X1 U15224 ( .A(n13059), .ZN(n13060) );
  AOI211_X1 U15225 ( .C1(n13062), .C2(n13061), .A(n13082), .B(n13060), .ZN(
        n13063) );
  AOI211_X1 U15226 ( .C1(n13522), .C2(n13093), .A(n13064), .B(n13063), .ZN(
        n13065) );
  INV_X1 U15227 ( .A(n13065), .ZN(P2_U3210) );
  OAI21_X1 U15228 ( .B1(n13077), .B2(n13067), .A(n13066), .ZN(n13068) );
  INV_X1 U15229 ( .A(n13068), .ZN(n13083) );
  INV_X1 U15230 ( .A(n13069), .ZN(n13246) );
  AOI22_X1 U15231 ( .A1(n13246), .A2(n13070), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13071) );
  OAI21_X1 U15232 ( .B1(n13073), .B2(n13072), .A(n13071), .ZN(n13074) );
  AOI21_X1 U15233 ( .B1(n13477), .B2(n13093), .A(n13074), .ZN(n13081) );
  NOR3_X1 U15234 ( .A1(n13077), .A2(n13076), .A3(n13075), .ZN(n13079) );
  OAI21_X1 U15235 ( .B1(n13079), .B2(n13078), .A(n13240), .ZN(n13080) );
  OAI211_X1 U15236 ( .C1(n13083), .C2(n13082), .A(n13081), .B(n13080), .ZN(
        P2_U3212) );
  AOI22_X1 U15237 ( .A1(n13086), .A2(n13085), .B1(n13084), .B2(n13104), .ZN(
        n13096) );
  NAND2_X1 U15238 ( .A1(n13103), .A2(n13441), .ZN(n13088) );
  NAND2_X1 U15239 ( .A1(n13442), .A2(n13444), .ZN(n13087) );
  NAND2_X1 U15240 ( .A1(n13088), .A2(n13087), .ZN(n13408) );
  AOI22_X1 U15241 ( .A1(n13089), .A2(n13408), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13090) );
  OAI21_X1 U15242 ( .B1(n13412), .B2(n13091), .A(n13090), .ZN(n13092) );
  AOI21_X1 U15243 ( .B1(n13538), .B2(n13093), .A(n13092), .ZN(n13094) );
  OAI21_X1 U15244 ( .B1(n13096), .B2(n13095), .A(n13094), .ZN(P2_U3213) );
  MUX2_X1 U15245 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13196), .S(P2_U3947), .Z(
        P2_U3562) );
  MUX2_X1 U15246 ( .A(n13097), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13117), .Z(
        P2_U3561) );
  MUX2_X1 U15247 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13209), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15248 ( .A(n13227), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13117), .Z(
        P2_U3559) );
  MUX2_X1 U15249 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13241), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15250 ( .A(n13259), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13117), .Z(
        P2_U3557) );
  MUX2_X1 U15251 ( .A(n13240), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13117), .Z(
        P2_U3556) );
  MUX2_X1 U15252 ( .A(n13258), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13117), .Z(
        P2_U3555) );
  MUX2_X1 U15253 ( .A(n13301), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13117), .Z(
        P2_U3554) );
  MUX2_X1 U15254 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13098), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15255 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13300), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15256 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13099), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15257 ( .A(n13100), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13117), .Z(
        P2_U3550) );
  MUX2_X1 U15258 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13101), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U15259 ( .A(n13102), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13117), .Z(
        P2_U3548) );
  MUX2_X1 U15260 ( .A(n13103), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13117), .Z(
        P2_U3547) );
  MUX2_X1 U15261 ( .A(n13104), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13117), .Z(
        P2_U3546) );
  MUX2_X1 U15262 ( .A(n13442), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13117), .Z(
        P2_U3545) );
  MUX2_X1 U15263 ( .A(n13105), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13117), .Z(
        P2_U3544) );
  MUX2_X1 U15264 ( .A(n13445), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13117), .Z(
        P2_U3543) );
  MUX2_X1 U15265 ( .A(n13106), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13117), .Z(
        P2_U3542) );
  MUX2_X1 U15266 ( .A(n13107), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13117), .Z(
        P2_U3541) );
  MUX2_X1 U15267 ( .A(n13108), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13117), .Z(
        P2_U3540) );
  MUX2_X1 U15268 ( .A(n13109), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13117), .Z(
        P2_U3539) );
  MUX2_X1 U15269 ( .A(n13110), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13117), .Z(
        P2_U3538) );
  MUX2_X1 U15270 ( .A(n13111), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13117), .Z(
        P2_U3537) );
  MUX2_X1 U15271 ( .A(n13112), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13117), .Z(
        P2_U3536) );
  MUX2_X1 U15272 ( .A(n13113), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13117), .Z(
        P2_U3535) );
  MUX2_X1 U15273 ( .A(n13114), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13117), .Z(
        P2_U3534) );
  MUX2_X1 U15274 ( .A(n13115), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13117), .Z(
        P2_U3533) );
  MUX2_X1 U15275 ( .A(n13116), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13117), .Z(
        P2_U3532) );
  MUX2_X1 U15276 ( .A(n13118), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13117), .Z(
        P2_U3531) );
  OAI211_X1 U15277 ( .C1(n13121), .C2(n13120), .A(n14816), .B(n13119), .ZN(
        n13131) );
  INV_X1 U15278 ( .A(n13122), .ZN(n13123) );
  AOI21_X1 U15279 ( .B1(n14840), .B2(n13124), .A(n13123), .ZN(n13130) );
  NAND2_X1 U15280 ( .A1(n14762), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n13129) );
  MUX2_X1 U15281 ( .A(n10102), .B(P2_REG2_REG_6__SCAN_IN), .S(n13124), .Z(
        n13125) );
  NAND3_X1 U15282 ( .A1(n14809), .A2(n13126), .A3(n13125), .ZN(n13127) );
  NAND3_X1 U15283 ( .A1(n14838), .A2(n13139), .A3(n13127), .ZN(n13128) );
  NAND4_X1 U15284 ( .A1(n13131), .A2(n13130), .A3(n13129), .A4(n13128), .ZN(
        P2_U3220) );
  OAI211_X1 U15285 ( .C1(n13134), .C2(n13133), .A(n14816), .B(n13132), .ZN(
        n13145) );
  AOI21_X1 U15286 ( .B1(n14840), .B2(n13136), .A(n13135), .ZN(n13144) );
  NAND2_X1 U15287 ( .A1(n14762), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n13143) );
  MUX2_X1 U15288 ( .A(n10105), .B(P2_REG2_REG_7__SCAN_IN), .S(n13136), .Z(
        n13137) );
  NAND3_X1 U15289 ( .A1(n13139), .A2(n13138), .A3(n13137), .ZN(n13140) );
  NAND3_X1 U15290 ( .A1(n14838), .A2(n13141), .A3(n13140), .ZN(n13142) );
  NAND4_X1 U15291 ( .A1(n13145), .A2(n13144), .A3(n13143), .A4(n13142), .ZN(
        P2_U3221) );
  INV_X1 U15292 ( .A(n13146), .ZN(n13149) );
  INV_X1 U15293 ( .A(n13147), .ZN(n13148) );
  OAI211_X1 U15294 ( .C1(n13149), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14816), 
        .B(n13148), .ZN(n13157) );
  AND2_X1 U15295 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13152) );
  NOR2_X1 U15296 ( .A1(n14794), .A2(n13150), .ZN(n13151) );
  AOI211_X1 U15297 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n14762), .A(n13152), 
        .B(n13151), .ZN(n13156) );
  OAI211_X1 U15298 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n13154), .A(n14838), 
        .B(n13153), .ZN(n13155) );
  NAND3_X1 U15299 ( .A1(n13157), .A2(n13156), .A3(n13155), .ZN(P2_U3229) );
  OAI21_X1 U15300 ( .B1(n13160), .B2(n13159), .A(n13158), .ZN(n13161) );
  NOR2_X1 U15301 ( .A1(n13161), .A2(n13162), .ZN(n13178) );
  AOI21_X1 U15302 ( .B1(n13162), .B2(n13161), .A(n13178), .ZN(n13163) );
  INV_X1 U15303 ( .A(n13163), .ZN(n13164) );
  NOR2_X1 U15304 ( .A1(n13164), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13179) );
  AOI21_X1 U15305 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13164), .A(n13179), 
        .ZN(n13177) );
  NOR2_X1 U15306 ( .A1(n13167), .A2(n13171), .ZN(n13181) );
  AOI21_X1 U15307 ( .B1(n13167), .B2(n13171), .A(n13181), .ZN(n13169) );
  AND2_X1 U15308 ( .A1(n13169), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13182) );
  INV_X1 U15309 ( .A(n13182), .ZN(n13168) );
  OAI211_X1 U15310 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13169), .A(n13168), 
        .B(n14816), .ZN(n13175) );
  NOR2_X1 U15311 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13170), .ZN(n13173) );
  NOR2_X1 U15312 ( .A1(n14794), .A2(n13171), .ZN(n13172) );
  AOI211_X1 U15313 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n14762), .A(n13173), 
        .B(n13172), .ZN(n13174) );
  OAI211_X1 U15314 ( .C1(n13177), .C2(n13176), .A(n13175), .B(n13174), .ZN(
        P2_U3232) );
  INV_X1 U15315 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13193) );
  NOR2_X1 U15316 ( .A1(n13179), .A2(n13178), .ZN(n13180) );
  XOR2_X1 U15317 ( .A(n13180), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13187) );
  INV_X1 U15318 ( .A(n13187), .ZN(n13185) );
  NOR2_X1 U15319 ( .A1(n13182), .A2(n13181), .ZN(n13183) );
  XNOR2_X1 U15320 ( .A(n13183), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13186) );
  OAI21_X1 U15321 ( .B1(n13186), .B2(n14844), .A(n14794), .ZN(n13184) );
  AOI21_X1 U15322 ( .B1(n14838), .B2(n13185), .A(n13184), .ZN(n13190) );
  AOI22_X1 U15323 ( .A1(n13187), .A2(n14838), .B1(n14816), .B2(n13186), .ZN(
        n13189) );
  OAI211_X1 U15324 ( .C1(n13193), .C2(n14848), .A(n13192), .B(n13191), .ZN(
        P2_U3233) );
  XNOR2_X1 U15325 ( .A(n13199), .B(n13458), .ZN(n13194) );
  NAND2_X1 U15326 ( .A1(n13194), .A2(n13215), .ZN(n13457) );
  NAND2_X1 U15327 ( .A1(n13196), .A2(n13195), .ZN(n13459) );
  NOR2_X1 U15328 ( .A1(n13459), .A2(n14890), .ZN(n13202) );
  NOR2_X1 U15329 ( .A1(n13458), .A2(n14874), .ZN(n13197) );
  AOI211_X1 U15330 ( .C1(n14890), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13202), 
        .B(n13197), .ZN(n13198) );
  OAI21_X1 U15331 ( .B1(n13457), .B2(n14868), .A(n13198), .ZN(P2_U3234) );
  OAI211_X1 U15332 ( .C1(n9125), .C2(n13200), .A(n13215), .B(n13199), .ZN(
        n13460) );
  NOR2_X1 U15333 ( .A1(n9125), .A2(n14874), .ZN(n13201) );
  AOI211_X1 U15334 ( .C1(n14890), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13202), 
        .B(n13201), .ZN(n13203) );
  OAI21_X1 U15335 ( .B1(n14868), .B2(n13460), .A(n13203), .ZN(P2_U3235) );
  XNOR2_X1 U15336 ( .A(n13204), .B(n13205), .ZN(n13470) );
  NAND2_X1 U15337 ( .A1(n13206), .A2(n14882), .ZN(n13212) );
  AOI21_X1 U15338 ( .B1(n13225), .B2(n13208), .A(n13207), .ZN(n13211) );
  AOI22_X1 U15339 ( .A1(n13241), .A2(n13444), .B1(n13209), .B2(n13441), .ZN(
        n13210) );
  OAI21_X1 U15340 ( .B1(n13212), .B2(n13211), .A(n13210), .ZN(n13467) );
  OR2_X1 U15341 ( .A1(n13213), .A2(n13230), .ZN(n13214) );
  NAND2_X1 U15342 ( .A1(n13466), .A2(n14850), .ZN(n13221) );
  OAI22_X1 U15343 ( .A1(n13218), .A2(n14881), .B1(n13217), .B2(n13402), .ZN(
        n13219) );
  AOI21_X1 U15344 ( .B1(n13465), .B2(n13433), .A(n13219), .ZN(n13220) );
  NAND2_X1 U15345 ( .A1(n13221), .A2(n13220), .ZN(n13222) );
  AOI21_X1 U15346 ( .B1(n13467), .B2(n13402), .A(n13222), .ZN(n13223) );
  OAI21_X1 U15347 ( .B1(n14871), .B2(n13470), .A(n13223), .ZN(P2_U3237) );
  XNOR2_X1 U15348 ( .A(n13226), .B(n13224), .ZN(n13475) );
  INV_X1 U15349 ( .A(n13474), .ZN(n13236) );
  NAND2_X1 U15350 ( .A1(n13472), .A2(n13243), .ZN(n13228) );
  NAND2_X1 U15351 ( .A1(n13228), .A2(n13215), .ZN(n13229) );
  NOR2_X1 U15352 ( .A1(n13230), .A2(n13229), .ZN(n13471) );
  NAND2_X1 U15353 ( .A1(n13471), .A2(n14850), .ZN(n13233) );
  AOI22_X1 U15354 ( .A1(n13231), .A2(n14865), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13456), .ZN(n13232) );
  OAI211_X1 U15355 ( .C1(n13234), .C2(n14874), .A(n13233), .B(n13232), .ZN(
        n13235) );
  AOI21_X1 U15356 ( .B1(n13236), .B2(n13402), .A(n13235), .ZN(n13237) );
  OAI21_X1 U15357 ( .B1(n13475), .B2(n14871), .A(n13237), .ZN(P2_U3238) );
  OAI21_X1 U15358 ( .B1(n13250), .B2(n13239), .A(n13238), .ZN(n13242) );
  AOI222_X1 U15359 ( .A1(n13242), .A2(n14882), .B1(n13241), .B2(n13441), .C1(
        n13240), .C2(n13444), .ZN(n13478) );
  INV_X1 U15360 ( .A(n13263), .ZN(n13245) );
  INV_X1 U15361 ( .A(n13243), .ZN(n13244) );
  AOI211_X1 U15362 ( .C1(n13477), .C2(n13245), .A(n9733), .B(n13244), .ZN(
        n13476) );
  AOI22_X1 U15363 ( .A1(n13246), .A2(n14865), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13456), .ZN(n13247) );
  OAI21_X1 U15364 ( .B1(n13248), .B2(n14874), .A(n13247), .ZN(n13252) );
  XNOR2_X1 U15365 ( .A(n13250), .B(n13249), .ZN(n13480) );
  NOR2_X1 U15366 ( .A1(n13480), .A2(n14871), .ZN(n13251) );
  AOI211_X1 U15367 ( .C1(n13476), .C2(n14850), .A(n13252), .B(n13251), .ZN(
        n13253) );
  OAI21_X1 U15368 ( .B1(n14890), .B2(n13478), .A(n13253), .ZN(P2_U3239) );
  XOR2_X1 U15369 ( .A(n13257), .B(n13254), .Z(n13485) );
  OAI21_X1 U15370 ( .B1(n13257), .B2(n13256), .A(n13255), .ZN(n13260) );
  AOI222_X1 U15371 ( .A1(n13260), .A2(n14882), .B1(n13259), .B2(n13441), .C1(
        n13258), .C2(n13444), .ZN(n13484) );
  INV_X1 U15372 ( .A(n13484), .ZN(n13268) );
  NAND2_X1 U15373 ( .A1(n13482), .A2(n13273), .ZN(n13261) );
  NAND2_X1 U15374 ( .A1(n13261), .A2(n13215), .ZN(n13262) );
  NOR2_X1 U15375 ( .A1(n13263), .A2(n13262), .ZN(n13481) );
  NAND2_X1 U15376 ( .A1(n13481), .A2(n14850), .ZN(n13266) );
  AOI22_X1 U15377 ( .A1(n13264), .A2(n14865), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13456), .ZN(n13265) );
  OAI211_X1 U15378 ( .C1(n7255), .C2(n14874), .A(n13266), .B(n13265), .ZN(
        n13267) );
  AOI21_X1 U15379 ( .B1(n13268), .B2(n13402), .A(n13267), .ZN(n13269) );
  OAI21_X1 U15380 ( .B1(n14871), .B2(n13485), .A(n13269), .ZN(P2_U3240) );
  XNOR2_X1 U15381 ( .A(n13270), .B(n13279), .ZN(n13272) );
  AOI21_X1 U15382 ( .B1(n13272), .B2(n14882), .A(n13271), .ZN(n13488) );
  INV_X1 U15383 ( .A(n13273), .ZN(n13274) );
  AOI211_X1 U15384 ( .C1(n13487), .C2(n13287), .A(n9733), .B(n13274), .ZN(
        n13486) );
  INV_X1 U15385 ( .A(n13275), .ZN(n13276) );
  AOI22_X1 U15386 ( .A1(n13276), .A2(n14865), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13456), .ZN(n13277) );
  OAI21_X1 U15387 ( .B1(n6888), .B2(n14874), .A(n13277), .ZN(n13281) );
  XNOR2_X1 U15388 ( .A(n13279), .B(n13278), .ZN(n13490) );
  NOR2_X1 U15389 ( .A1(n13490), .A2(n14871), .ZN(n13280) );
  AOI211_X1 U15390 ( .C1(n13486), .C2(n14850), .A(n13281), .B(n13280), .ZN(
        n13282) );
  OAI21_X1 U15391 ( .B1(n14890), .B2(n13488), .A(n13282), .ZN(P2_U3241) );
  XNOR2_X1 U15392 ( .A(n13283), .B(n13291), .ZN(n13286) );
  INV_X1 U15393 ( .A(n13284), .ZN(n13285) );
  AOI21_X1 U15394 ( .B1(n13286), .B2(n14882), .A(n13285), .ZN(n13493) );
  AOI211_X1 U15395 ( .C1(n13492), .C2(n13304), .A(n9733), .B(n6889), .ZN(
        n13491) );
  INV_X1 U15396 ( .A(n13492), .ZN(n13290) );
  AOI22_X1 U15397 ( .A1(n13288), .A2(n14865), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n13456), .ZN(n13289) );
  OAI21_X1 U15398 ( .B1(n13290), .B2(n14874), .A(n13289), .ZN(n13294) );
  XNOR2_X1 U15399 ( .A(n13292), .B(n13291), .ZN(n13495) );
  NOR2_X1 U15400 ( .A1(n13495), .A2(n14871), .ZN(n13293) );
  AOI211_X1 U15401 ( .C1(n13491), .C2(n14850), .A(n13294), .B(n13293), .ZN(
        n13295) );
  OAI21_X1 U15402 ( .B1(n14890), .B2(n13493), .A(n13295), .ZN(P2_U3242) );
  NAND2_X1 U15403 ( .A1(n13297), .A2(n13296), .ZN(n13298) );
  NAND3_X1 U15404 ( .A1(n13299), .A2(n14882), .A3(n13298), .ZN(n13303) );
  AOI22_X1 U15405 ( .A1(n13301), .A2(n13441), .B1(n13444), .B2(n13300), .ZN(
        n13302) );
  AOI21_X1 U15406 ( .B1(n13498), .B2(n13320), .A(n9733), .ZN(n13305) );
  NAND2_X1 U15407 ( .A1(n13305), .A2(n13304), .ZN(n13499) );
  AOI22_X1 U15408 ( .A1(n14890), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13306), 
        .B2(n14865), .ZN(n13308) );
  NAND2_X1 U15409 ( .A1(n13498), .A2(n13433), .ZN(n13307) );
  OAI211_X1 U15410 ( .C1(n13499), .C2(n14868), .A(n13308), .B(n13307), .ZN(
        n13309) );
  INV_X1 U15411 ( .A(n13309), .ZN(n13313) );
  NAND2_X1 U15412 ( .A1(n13311), .A2(n13310), .ZN(n13496) );
  NAND3_X1 U15413 ( .A1(n13497), .A2(n13496), .A3(n14859), .ZN(n13312) );
  OAI211_X1 U15414 ( .C1(n13503), .C2(n14890), .A(n13313), .B(n13312), .ZN(
        P2_U3243) );
  XNOR2_X1 U15415 ( .A(n13314), .B(n13318), .ZN(n13315) );
  NAND2_X1 U15416 ( .A1(n13315), .A2(n14882), .ZN(n13317) );
  NAND2_X1 U15417 ( .A1(n13317), .A2(n13316), .ZN(n13508) );
  INV_X1 U15418 ( .A(n13508), .ZN(n13329) );
  XNOR2_X1 U15419 ( .A(n13319), .B(n13318), .ZN(n13504) );
  AOI21_X1 U15420 ( .B1(n13325), .B2(n13338), .A(n9733), .ZN(n13321) );
  NAND2_X1 U15421 ( .A1(n13321), .A2(n13320), .ZN(n13505) );
  OAI22_X1 U15422 ( .A1(n13402), .A2(n13323), .B1(n13322), .B2(n14881), .ZN(
        n13324) );
  AOI21_X1 U15423 ( .B1(n13325), .B2(n13433), .A(n13324), .ZN(n13326) );
  OAI21_X1 U15424 ( .B1(n13505), .B2(n14868), .A(n13326), .ZN(n13327) );
  AOI21_X1 U15425 ( .B1(n13504), .B2(n14859), .A(n13327), .ZN(n13328) );
  OAI21_X1 U15426 ( .B1(n13329), .B2(n14890), .A(n13328), .ZN(P2_U3244) );
  XOR2_X1 U15427 ( .A(n13330), .B(n13334), .Z(n13513) );
  INV_X1 U15428 ( .A(n13331), .ZN(n13332) );
  AOI21_X1 U15429 ( .B1(n13334), .B2(n13333), .A(n13332), .ZN(n13335) );
  OAI222_X1 U15430 ( .A1(n13422), .A2(n13337), .B1(n14885), .B2(n13336), .C1(
        n13335), .C2(n13424), .ZN(n13509) );
  NAND2_X1 U15431 ( .A1(n13509), .A2(n13402), .ZN(n13344) );
  INV_X1 U15432 ( .A(n13338), .ZN(n13339) );
  AOI211_X1 U15433 ( .C1(n13511), .C2(n13354), .A(n9733), .B(n13339), .ZN(
        n13510) );
  AOI22_X1 U15434 ( .A1(n14890), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13340), 
        .B2(n14865), .ZN(n13341) );
  OAI21_X1 U15435 ( .B1(n7148), .B2(n14874), .A(n13341), .ZN(n13342) );
  AOI21_X1 U15436 ( .B1(n13510), .B2(n14850), .A(n13342), .ZN(n13343) );
  OAI211_X1 U15437 ( .C1(n13513), .C2(n14871), .A(n13344), .B(n13343), .ZN(
        P2_U3245) );
  XNOR2_X1 U15438 ( .A(n13345), .B(n13347), .ZN(n13519) );
  XOR2_X1 U15439 ( .A(n13347), .B(n13346), .Z(n13348) );
  NAND2_X1 U15440 ( .A1(n13348), .A2(n14882), .ZN(n13518) );
  OAI22_X1 U15441 ( .A1(n13350), .A2(n14885), .B1(n13349), .B2(n13422), .ZN(
        n13515) );
  INV_X1 U15442 ( .A(n13515), .ZN(n13351) );
  OAI211_X1 U15443 ( .C1(n14881), .C2(n13352), .A(n13518), .B(n13351), .ZN(
        n13353) );
  NAND2_X1 U15444 ( .A1(n13353), .A2(n13402), .ZN(n13358) );
  AOI211_X1 U15445 ( .C1(n13516), .C2(n13365), .A(n9733), .B(n7149), .ZN(
        n13514) );
  OAI22_X1 U15446 ( .A1(n6597), .A2(n14874), .B1(n13355), .B2(n13402), .ZN(
        n13356) );
  AOI21_X1 U15447 ( .B1(n13514), .B2(n14850), .A(n13356), .ZN(n13357) );
  OAI211_X1 U15448 ( .C1(n13519), .C2(n14871), .A(n13358), .B(n13357), .ZN(
        P2_U3246) );
  XOR2_X1 U15449 ( .A(n13359), .B(n13364), .Z(n13361) );
  AOI21_X1 U15450 ( .B1(n13361), .B2(n14882), .A(n13360), .ZN(n13524) );
  OAI21_X1 U15451 ( .B1(n13364), .B2(n13363), .A(n13362), .ZN(n13520) );
  INV_X1 U15452 ( .A(n13522), .ZN(n13370) );
  AOI211_X1 U15453 ( .C1(n13522), .C2(n13376), .A(n9733), .B(n6887), .ZN(
        n13521) );
  NAND2_X1 U15454 ( .A1(n13521), .A2(n14850), .ZN(n13369) );
  INV_X1 U15455 ( .A(n13366), .ZN(n13367) );
  AOI22_X1 U15456 ( .A1(n14890), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13367), 
        .B2(n14865), .ZN(n13368) );
  OAI211_X1 U15457 ( .C1(n13370), .C2(n14874), .A(n13369), .B(n13368), .ZN(
        n13371) );
  AOI21_X1 U15458 ( .B1(n13520), .B2(n14859), .A(n13371), .ZN(n13372) );
  OAI21_X1 U15459 ( .B1(n13524), .B2(n14890), .A(n13372), .ZN(P2_U3247) );
  XNOR2_X1 U15460 ( .A(n13373), .B(n13383), .ZN(n13375) );
  AOI21_X1 U15461 ( .B1(n13375), .B2(n14882), .A(n13374), .ZN(n13529) );
  INV_X1 U15462 ( .A(n13398), .ZN(n13378) );
  INV_X1 U15463 ( .A(n13376), .ZN(n13377) );
  AOI211_X1 U15464 ( .C1(n13527), .C2(n13378), .A(n9733), .B(n13377), .ZN(
        n13526) );
  INV_X1 U15465 ( .A(n13379), .ZN(n13380) );
  AOI22_X1 U15466 ( .A1(n14890), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13380), 
        .B2(n14865), .ZN(n13381) );
  OAI21_X1 U15467 ( .B1(n13382), .B2(n14874), .A(n13381), .ZN(n13386) );
  XOR2_X1 U15468 ( .A(n13384), .B(n13383), .Z(n13530) );
  NOR2_X1 U15469 ( .A1(n13530), .A2(n14871), .ZN(n13385) );
  AOI211_X1 U15470 ( .C1(n13526), .C2(n14850), .A(n13386), .B(n13385), .ZN(
        n13387) );
  OAI21_X1 U15471 ( .B1(n14890), .B2(n13529), .A(n13387), .ZN(P2_U3248) );
  NAND2_X1 U15472 ( .A1(n13389), .A2(n13388), .ZN(n13390) );
  NAND2_X1 U15473 ( .A1(n13391), .A2(n13390), .ZN(n13536) );
  INV_X1 U15474 ( .A(n13392), .ZN(n13393) );
  AOI21_X1 U15475 ( .B1(n13395), .B2(n13394), .A(n13393), .ZN(n13397) );
  OAI21_X1 U15476 ( .B1(n13397), .B2(n13424), .A(n13396), .ZN(n13531) );
  NAND2_X1 U15477 ( .A1(n13531), .A2(n13402), .ZN(n13406) );
  AOI211_X1 U15478 ( .C1(n13533), .C2(n13410), .A(n9733), .B(n13398), .ZN(
        n13532) );
  INV_X1 U15479 ( .A(n13533), .ZN(n13399) );
  NOR2_X1 U15480 ( .A1(n13399), .A2(n14874), .ZN(n13404) );
  OAI22_X1 U15481 ( .A1(n13402), .A2(n13401), .B1(n13400), .B2(n14881), .ZN(
        n13403) );
  AOI211_X1 U15482 ( .C1(n13532), .C2(n14850), .A(n13404), .B(n13403), .ZN(
        n13405) );
  OAI211_X1 U15483 ( .C1(n14871), .C2(n13536), .A(n13406), .B(n13405), .ZN(
        P2_U3249) );
  XOR2_X1 U15484 ( .A(n13407), .B(n13415), .Z(n13409) );
  AOI21_X1 U15485 ( .B1(n13409), .B2(n14882), .A(n13408), .ZN(n13540) );
  INV_X1 U15486 ( .A(n13410), .ZN(n13411) );
  AOI211_X1 U15487 ( .C1(n13538), .C2(n13429), .A(n9733), .B(n13411), .ZN(
        n13537) );
  INV_X1 U15488 ( .A(n13412), .ZN(n13413) );
  AOI22_X1 U15489 ( .A1(n14890), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13413), 
        .B2(n14865), .ZN(n13414) );
  OAI21_X1 U15490 ( .B1(n7143), .B2(n14874), .A(n13414), .ZN(n13418) );
  XOR2_X1 U15491 ( .A(n13416), .B(n13415), .Z(n13541) );
  NOR2_X1 U15492 ( .A1(n13541), .A2(n14871), .ZN(n13417) );
  AOI211_X1 U15493 ( .C1(n13537), .C2(n14850), .A(n13418), .B(n13417), .ZN(
        n13419) );
  OAI21_X1 U15494 ( .B1(n14890), .B2(n13540), .A(n13419), .ZN(P2_U3250) );
  XNOR2_X1 U15495 ( .A(n13420), .B(n13426), .ZN(n13425) );
  OAI222_X1 U15496 ( .A1(n13425), .A2(n13424), .B1(n14885), .B2(n13423), .C1(
        n13422), .C2(n13421), .ZN(n14495) );
  INV_X1 U15497 ( .A(n14495), .ZN(n13438) );
  XNOR2_X1 U15498 ( .A(n13427), .B(n13426), .ZN(n14497) );
  INV_X1 U15499 ( .A(n13428), .ZN(n13446) );
  OAI211_X1 U15500 ( .C1(n14494), .C2(n13446), .A(n13215), .B(n13429), .ZN(
        n14493) );
  OAI22_X1 U15501 ( .A1(n13402), .A2(n13431), .B1(n13430), .B2(n14881), .ZN(
        n13432) );
  AOI21_X1 U15502 ( .B1(n13434), .B2(n13433), .A(n13432), .ZN(n13435) );
  OAI21_X1 U15503 ( .B1(n14493), .B2(n14868), .A(n13435), .ZN(n13436) );
  AOI21_X1 U15504 ( .B1(n14497), .B2(n14859), .A(n13436), .ZN(n13437) );
  OAI21_X1 U15505 ( .B1(n13438), .B2(n13456), .A(n13437), .ZN(P2_U3251) );
  XNOR2_X1 U15506 ( .A(n13440), .B(n13439), .ZN(n13443) );
  AOI222_X1 U15507 ( .A1(n13445), .A2(n13444), .B1(n14882), .B2(n13443), .C1(
        n13442), .C2(n13441), .ZN(n13545) );
  AOI211_X1 U15508 ( .C1(n13543), .C2(n13447), .A(n9733), .B(n13446), .ZN(
        n13542) );
  INV_X1 U15509 ( .A(n13448), .ZN(n13449) );
  AOI22_X1 U15510 ( .A1(n14890), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n13449), 
        .B2(n14865), .ZN(n13450) );
  OAI21_X1 U15511 ( .B1(n6590), .B2(n14874), .A(n13450), .ZN(n13454) );
  XNOR2_X1 U15512 ( .A(n13452), .B(n13451), .ZN(n13546) );
  NOR2_X1 U15513 ( .A1(n13546), .A2(n14871), .ZN(n13453) );
  AOI211_X1 U15514 ( .C1(n13542), .C2(n14850), .A(n13454), .B(n13453), .ZN(
        n13455) );
  OAI21_X1 U15515 ( .B1(n13545), .B2(n13456), .A(n13455), .ZN(P2_U3252) );
  OAI211_X1 U15516 ( .C1(n13458), .C2(n14953), .A(n13457), .B(n13459), .ZN(
        n13554) );
  MUX2_X1 U15517 ( .A(n13554), .B(P2_REG1_REG_31__SCAN_IN), .S(n14971), .Z(
        P2_U3530) );
  OAI211_X1 U15518 ( .C1(n9125), .C2(n14953), .A(n13460), .B(n13459), .ZN(
        n13555) );
  MUX2_X1 U15519 ( .A(n13555), .B(P2_REG1_REG_30__SCAN_IN), .S(n14971), .Z(
        P2_U3529) );
  AOI21_X1 U15520 ( .B1(n14930), .B2(n13462), .A(n13461), .ZN(n13463) );
  INV_X1 U15521 ( .A(n13466), .ZN(n13469) );
  INV_X1 U15522 ( .A(n13467), .ZN(n13468) );
  MUX2_X1 U15523 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13556), .S(n14974), .Z(
        P2_U3527) );
  AOI21_X1 U15524 ( .B1(n14930), .B2(n13472), .A(n13471), .ZN(n13473) );
  OAI211_X1 U15525 ( .C1(n14934), .C2(n13475), .A(n13474), .B(n13473), .ZN(
        n13557) );
  MUX2_X1 U15526 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13557), .S(n14974), .Z(
        P2_U3526) );
  AOI21_X1 U15527 ( .B1(n14930), .B2(n13477), .A(n13476), .ZN(n13479) );
  MUX2_X1 U15528 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13558), .S(n14974), .Z(
        P2_U3525) );
  AOI21_X1 U15529 ( .B1(n14930), .B2(n13482), .A(n13481), .ZN(n13483) );
  OAI211_X1 U15530 ( .C1(n14934), .C2(n13485), .A(n13484), .B(n13483), .ZN(
        n13559) );
  MUX2_X1 U15531 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13559), .S(n14974), .Z(
        P2_U3524) );
  AOI21_X1 U15532 ( .B1(n14930), .B2(n13487), .A(n13486), .ZN(n13489) );
  OAI211_X1 U15533 ( .C1(n14934), .C2(n13490), .A(n13489), .B(n13488), .ZN(
        n13560) );
  MUX2_X1 U15534 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13560), .S(n14974), .Z(
        P2_U3523) );
  AOI21_X1 U15535 ( .B1(n14930), .B2(n13492), .A(n13491), .ZN(n13494) );
  OAI211_X1 U15536 ( .C1(n14934), .C2(n13495), .A(n13494), .B(n13493), .ZN(
        n13561) );
  MUX2_X1 U15537 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13561), .S(n14974), .Z(
        P2_U3522) );
  NAND3_X1 U15538 ( .A1(n13497), .A2(n13496), .A3(n14918), .ZN(n13501) );
  NAND2_X1 U15539 ( .A1(n13498), .A2(n14930), .ZN(n13500) );
  NAND2_X1 U15540 ( .A1(n13503), .A2(n13502), .ZN(n13562) );
  MUX2_X1 U15541 ( .A(n13562), .B(P2_REG1_REG_22__SCAN_IN), .S(n14971), .Z(
        P2_U3521) );
  NAND2_X1 U15542 ( .A1(n13504), .A2(n14918), .ZN(n13506) );
  OAI211_X1 U15543 ( .C1(n7261), .C2(n14953), .A(n13506), .B(n13505), .ZN(
        n13507) );
  MUX2_X1 U15544 ( .A(n13563), .B(P2_REG1_REG_21__SCAN_IN), .S(n14971), .Z(
        P2_U3520) );
  AOI211_X1 U15545 ( .C1(n14930), .C2(n13511), .A(n13510), .B(n13509), .ZN(
        n13512) );
  OAI21_X1 U15546 ( .B1(n14934), .B2(n13513), .A(n13512), .ZN(n13564) );
  MUX2_X1 U15547 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13564), .S(n14974), .Z(
        P2_U3519) );
  AOI211_X1 U15548 ( .C1(n14930), .C2(n13516), .A(n13515), .B(n13514), .ZN(
        n13517) );
  OAI211_X1 U15549 ( .C1(n14934), .C2(n13519), .A(n13518), .B(n13517), .ZN(
        n13565) );
  MUX2_X1 U15550 ( .A(n13565), .B(P2_REG1_REG_19__SCAN_IN), .S(n14971), .Z(
        P2_U3518) );
  INV_X1 U15551 ( .A(n13520), .ZN(n13525) );
  AOI21_X1 U15552 ( .B1(n14930), .B2(n13522), .A(n13521), .ZN(n13523) );
  OAI211_X1 U15553 ( .C1(n14934), .C2(n13525), .A(n13524), .B(n13523), .ZN(
        n13566) );
  MUX2_X1 U15554 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13566), .S(n14974), .Z(
        P2_U3517) );
  AOI21_X1 U15555 ( .B1(n14930), .B2(n13527), .A(n13526), .ZN(n13528) );
  OAI211_X1 U15556 ( .C1(n14934), .C2(n13530), .A(n13529), .B(n13528), .ZN(
        n13567) );
  MUX2_X1 U15557 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13567), .S(n14974), .Z(
        P2_U3516) );
  INV_X1 U15558 ( .A(n13531), .ZN(n13535) );
  AOI21_X1 U15559 ( .B1(n14930), .B2(n13533), .A(n13532), .ZN(n13534) );
  OAI211_X1 U15560 ( .C1(n14934), .C2(n13536), .A(n13535), .B(n13534), .ZN(
        n13568) );
  MUX2_X1 U15561 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13568), .S(n14974), .Z(
        P2_U3515) );
  AOI21_X1 U15562 ( .B1(n14930), .B2(n13538), .A(n13537), .ZN(n13539) );
  OAI211_X1 U15563 ( .C1(n14934), .C2(n13541), .A(n13540), .B(n13539), .ZN(
        n13569) );
  MUX2_X1 U15564 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13569), .S(n14974), .Z(
        P2_U3514) );
  AOI21_X1 U15565 ( .B1(n14930), .B2(n13543), .A(n13542), .ZN(n13544) );
  OAI211_X1 U15566 ( .C1(n14934), .C2(n13546), .A(n13545), .B(n13544), .ZN(
        n13570) );
  MUX2_X1 U15567 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13570), .S(n14974), .Z(
        P2_U3512) );
  INV_X1 U15568 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n13553) );
  AOI211_X1 U15569 ( .C1(n14930), .C2(n13549), .A(n13548), .B(n13547), .ZN(
        n13550) );
  OAI21_X1 U15570 ( .B1(n14934), .B2(n13551), .A(n13550), .ZN(n13571) );
  NAND2_X1 U15571 ( .A1(n13571), .A2(n14974), .ZN(n13552) );
  OAI21_X1 U15572 ( .B1(n14974), .B2(n13553), .A(n13552), .ZN(P2_U3510) );
  MUX2_X1 U15573 ( .A(n13554), .B(P2_REG0_REG_31__SCAN_IN), .S(n14958), .Z(
        P2_U3498) );
  MUX2_X1 U15574 ( .A(n13555), .B(P2_REG0_REG_30__SCAN_IN), .S(n14958), .Z(
        P2_U3497) );
  MUX2_X1 U15575 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13556), .S(n14959), .Z(
        P2_U3495) );
  MUX2_X1 U15576 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13557), .S(n14959), .Z(
        P2_U3494) );
  MUX2_X1 U15577 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13559), .S(n14959), .Z(
        P2_U3492) );
  MUX2_X1 U15578 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13560), .S(n14959), .Z(
        P2_U3491) );
  MUX2_X1 U15579 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13561), .S(n14959), .Z(
        P2_U3490) );
  MUX2_X1 U15580 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13562), .S(n14959), .Z(
        P2_U3489) );
  MUX2_X1 U15581 ( .A(n13563), .B(P2_REG0_REG_21__SCAN_IN), .S(n14958), .Z(
        P2_U3488) );
  MUX2_X1 U15582 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13564), .S(n14959), .Z(
        P2_U3487) );
  MUX2_X1 U15583 ( .A(n13565), .B(P2_REG0_REG_19__SCAN_IN), .S(n14958), .Z(
        P2_U3486) );
  MUX2_X1 U15584 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13566), .S(n14959), .Z(
        P2_U3484) );
  MUX2_X1 U15585 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13567), .S(n14959), .Z(
        P2_U3481) );
  MUX2_X1 U15586 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13568), .S(n14959), .Z(
        P2_U3478) );
  MUX2_X1 U15587 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13569), .S(n14959), .Z(
        P2_U3475) );
  MUX2_X1 U15588 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13570), .S(n14959), .Z(
        P2_U3469) );
  NAND2_X1 U15589 ( .A1(n13571), .A2(n14959), .ZN(n13572) );
  OAI21_X1 U15590 ( .B1(n14959), .B2(n8702), .A(n13572), .ZN(P2_U3463) );
  NAND3_X1 U15591 ( .A1(n13574), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13575) );
  OAI22_X1 U15592 ( .A1(n13573), .A2(n13575), .B1(n15195), .B2(n13588), .ZN(
        n13576) );
  AOI21_X1 U15593 ( .B1(n14342), .B2(n13577), .A(n13576), .ZN(n13578) );
  INV_X1 U15594 ( .A(n13578), .ZN(P2_U3296) );
  OAI222_X1 U15595 ( .A1(n13588), .A2(n13581), .B1(n13590), .B2(n13580), .C1(
        P2_U3088), .C2(n13579), .ZN(P2_U3300) );
  OAI222_X1 U15596 ( .A1(P2_U3088), .A2(n13583), .B1(n13590), .B2(n14349), 
        .C1(n13582), .C2(n13588), .ZN(P2_U3301) );
  INV_X1 U15597 ( .A(n13584), .ZN(n14352) );
  OAI222_X1 U15598 ( .A1(n13588), .A2(n13586), .B1(n13590), .B2(n14352), .C1(
        P2_U3088), .C2(n13585), .ZN(P2_U3302) );
  INV_X1 U15599 ( .A(n13587), .ZN(n14356) );
  OAI222_X1 U15600 ( .A1(P2_U3088), .A2(n13591), .B1(n13590), .B2(n14356), 
        .C1(n13589), .C2(n13588), .ZN(P2_U3303) );
  INV_X1 U15601 ( .A(n13593), .ZN(n13594) );
  MUX2_X1 U15602 ( .A(n13594), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15603 ( .A1(n14022), .A2(n13699), .ZN(n13596) );
  NAND2_X1 U15604 ( .A1(n14030), .A2(n13608), .ZN(n13595) );
  NAND2_X1 U15605 ( .A1(n13596), .A2(n13595), .ZN(n13597) );
  XNOR2_X1 U15606 ( .A(n13597), .B(n13750), .ZN(n13601) );
  NAND2_X1 U15607 ( .A1(n14022), .A2(n13608), .ZN(n13599) );
  NAND2_X1 U15608 ( .A1(n14030), .A2(n13704), .ZN(n13598) );
  NAND2_X1 U15609 ( .A1(n13599), .A2(n13598), .ZN(n13600) );
  NOR2_X1 U15610 ( .A1(n13601), .A2(n13600), .ZN(n13747) );
  AOI21_X1 U15611 ( .B1(n13601), .B2(n13600), .A(n13747), .ZN(n13712) );
  INV_X1 U15612 ( .A(n13602), .ZN(n13605) );
  INV_X1 U15613 ( .A(n13603), .ZN(n13604) );
  AOI22_X1 U15614 ( .A1(n14233), .A2(n13699), .B1(n13608), .B2(n13865), .ZN(
        n13609) );
  XOR2_X1 U15615 ( .A(n13750), .B(n13609), .Z(n13611) );
  INV_X1 U15616 ( .A(n14233), .ZN(n14545) );
  OAI22_X1 U15617 ( .A1(n14545), .A2(n13752), .B1(n13850), .B2(n13749), .ZN(
        n13610) );
  NOR2_X1 U15618 ( .A1(n13611), .A2(n13610), .ZN(n13612) );
  AOI21_X1 U15619 ( .B1(n13611), .B2(n13610), .A(n13612), .ZN(n13720) );
  INV_X1 U15620 ( .A(n13612), .ZN(n13613) );
  NAND2_X1 U15621 ( .A1(n14214), .A2(n13699), .ZN(n13615) );
  OR2_X1 U15622 ( .A1(n14508), .A2(n13752), .ZN(n13614) );
  NAND2_X1 U15623 ( .A1(n13615), .A2(n13614), .ZN(n13616) );
  XNOR2_X1 U15624 ( .A(n13616), .B(n6937), .ZN(n13618) );
  AOI22_X1 U15625 ( .A1(n14214), .A2(n13608), .B1(n13704), .B2(n14222), .ZN(
        n13848) );
  NAND2_X1 U15626 ( .A1(n14518), .A2(n13699), .ZN(n13620) );
  NAND2_X1 U15627 ( .A1(n14182), .A2(n13700), .ZN(n13619) );
  NAND2_X1 U15628 ( .A1(n13620), .A2(n13619), .ZN(n13621) );
  XNOR2_X1 U15629 ( .A(n13621), .B(n6937), .ZN(n13624) );
  AND2_X1 U15630 ( .A1(n14182), .A2(n13704), .ZN(n13622) );
  NAND2_X1 U15631 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  OAI21_X1 U15632 ( .B1(n13624), .B2(n13623), .A(n13625), .ZN(n14514) );
  INV_X1 U15633 ( .A(n13625), .ZN(n13795) );
  OAI22_X1 U15634 ( .A1(n14311), .A2(n13754), .B1(n14511), .B2(n13752), .ZN(
        n13626) );
  XNOR2_X1 U15635 ( .A(n13626), .B(n6937), .ZN(n13629) );
  OR2_X1 U15636 ( .A1(n14311), .A2(n13752), .ZN(n13628) );
  NAND2_X1 U15637 ( .A1(n14195), .A2(n13704), .ZN(n13627) );
  AND2_X1 U15638 ( .A1(n13628), .A2(n13627), .ZN(n13630) );
  NAND2_X1 U15639 ( .A1(n13629), .A2(n13630), .ZN(n13634) );
  INV_X1 U15640 ( .A(n13629), .ZN(n13632) );
  INV_X1 U15641 ( .A(n13630), .ZN(n13631) );
  NAND2_X1 U15642 ( .A1(n13632), .A2(n13631), .ZN(n13633) );
  AND2_X1 U15643 ( .A1(n13634), .A2(n13633), .ZN(n13794) );
  NAND2_X1 U15644 ( .A1(n13793), .A2(n13634), .ZN(n13828) );
  NAND2_X1 U15645 ( .A1(n14306), .A2(n13699), .ZN(n13636) );
  NAND2_X1 U15646 ( .A1(n14183), .A2(n13608), .ZN(n13635) );
  NAND2_X1 U15647 ( .A1(n13636), .A2(n13635), .ZN(n13637) );
  XNOR2_X1 U15648 ( .A(n13637), .B(n13750), .ZN(n13644) );
  AOI22_X1 U15649 ( .A1(n14306), .A2(n13608), .B1(n13704), .B2(n14183), .ZN(
        n13642) );
  XNOR2_X1 U15650 ( .A(n13644), .B(n13642), .ZN(n13829) );
  NAND2_X1 U15651 ( .A1(n13828), .A2(n13829), .ZN(n13827) );
  NAND2_X1 U15652 ( .A1(n14299), .A2(n13699), .ZN(n13639) );
  OR2_X1 U15653 ( .A1(n14164), .A2(n13752), .ZN(n13638) );
  NAND2_X1 U15654 ( .A1(n13639), .A2(n13638), .ZN(n13640) );
  XNOR2_X1 U15655 ( .A(n13640), .B(n6937), .ZN(n13647) );
  NOR2_X1 U15656 ( .A1(n14164), .A2(n13749), .ZN(n13641) );
  XNOR2_X1 U15657 ( .A(n13647), .B(n13646), .ZN(n13737) );
  INV_X1 U15658 ( .A(n13642), .ZN(n13643) );
  NOR2_X1 U15659 ( .A1(n13644), .A2(n13643), .ZN(n13738) );
  NOR2_X1 U15660 ( .A1(n13737), .A2(n13738), .ZN(n13645) );
  OR2_X1 U15661 ( .A1(n13647), .A2(n13646), .ZN(n13648) );
  OAI22_X1 U15662 ( .A1(n13650), .A2(n13752), .B1(n13649), .B2(n13749), .ZN(
        n13652) );
  OAI22_X1 U15663 ( .A1(n13650), .A2(n13754), .B1(n13649), .B2(n13752), .ZN(
        n13651) );
  XNOR2_X1 U15664 ( .A(n13651), .B(n13750), .ZN(n13653) );
  XOR2_X1 U15665 ( .A(n13652), .B(n13653), .Z(n13811) );
  NAND2_X1 U15666 ( .A1(n13653), .A2(n13652), .ZN(n13654) );
  NAND2_X1 U15667 ( .A1(n14288), .A2(n13699), .ZN(n13657) );
  NAND2_X1 U15668 ( .A1(n13863), .A2(n13700), .ZN(n13656) );
  NAND2_X1 U15669 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  XNOR2_X1 U15670 ( .A(n13658), .B(n6937), .ZN(n13661) );
  AND2_X1 U15671 ( .A1(n13863), .A2(n13704), .ZN(n13659) );
  NAND2_X1 U15672 ( .A1(n13661), .A2(n13660), .ZN(n13662) );
  OAI21_X1 U15673 ( .B1(n13661), .B2(n13660), .A(n13662), .ZN(n13774) );
  NAND2_X1 U15674 ( .A1(n14283), .A2(n13699), .ZN(n13664) );
  NAND2_X1 U15675 ( .A1(n13862), .A2(n13700), .ZN(n13663) );
  NAND2_X1 U15676 ( .A1(n13664), .A2(n13663), .ZN(n13665) );
  XNOR2_X1 U15677 ( .A(n13665), .B(n13750), .ZN(n13669) );
  NAND2_X1 U15678 ( .A1(n14283), .A2(n13700), .ZN(n13667) );
  NAND2_X1 U15679 ( .A1(n13862), .A2(n13704), .ZN(n13666) );
  NAND2_X1 U15680 ( .A1(n13667), .A2(n13666), .ZN(n13668) );
  NOR2_X1 U15681 ( .A1(n13669), .A2(n13668), .ZN(n13670) );
  AOI21_X1 U15682 ( .B1(n13669), .B2(n13668), .A(n13670), .ZN(n13820) );
  INV_X1 U15683 ( .A(n13670), .ZN(n13671) );
  NAND2_X1 U15684 ( .A1(n14089), .A2(n13699), .ZN(n13673) );
  NAND2_X1 U15685 ( .A1(n13861), .A2(n13700), .ZN(n13672) );
  NAND2_X1 U15686 ( .A1(n13673), .A2(n13672), .ZN(n13674) );
  XNOR2_X1 U15687 ( .A(n13674), .B(n13750), .ZN(n13678) );
  NAND2_X1 U15688 ( .A1(n14089), .A2(n13700), .ZN(n13676) );
  NAND2_X1 U15689 ( .A1(n13861), .A2(n13704), .ZN(n13675) );
  NAND2_X1 U15690 ( .A1(n13676), .A2(n13675), .ZN(n13677) );
  NOR2_X1 U15691 ( .A1(n13678), .A2(n13677), .ZN(n13679) );
  AOI21_X1 U15692 ( .B1(n13678), .B2(n13677), .A(n13679), .ZN(n13729) );
  NAND2_X1 U15693 ( .A1(n13728), .A2(n13729), .ZN(n13727) );
  INV_X1 U15694 ( .A(n13679), .ZN(n13680) );
  NAND2_X1 U15695 ( .A1(n14274), .A2(n13699), .ZN(n13682) );
  NAND2_X1 U15696 ( .A1(n13860), .A2(n13700), .ZN(n13681) );
  NAND2_X1 U15697 ( .A1(n13682), .A2(n13681), .ZN(n13683) );
  XNOR2_X1 U15698 ( .A(n13683), .B(n13750), .ZN(n13687) );
  NAND2_X1 U15699 ( .A1(n14274), .A2(n13700), .ZN(n13685) );
  NAND2_X1 U15700 ( .A1(n13860), .A2(n13704), .ZN(n13684) );
  NAND2_X1 U15701 ( .A1(n13685), .A2(n13684), .ZN(n13686) );
  NOR2_X1 U15702 ( .A1(n13687), .A2(n13686), .ZN(n13688) );
  AOI21_X1 U15703 ( .B1(n13687), .B2(n13686), .A(n13688), .ZN(n13805) );
  NAND2_X1 U15704 ( .A1(n13804), .A2(n13805), .ZN(n13803) );
  INV_X1 U15705 ( .A(n13688), .ZN(n13689) );
  NAND2_X1 U15706 ( .A1(n13803), .A2(n13689), .ZN(n13784) );
  NAND2_X1 U15707 ( .A1(n14269), .A2(n13699), .ZN(n13691) );
  NAND2_X1 U15708 ( .A1(n14029), .A2(n13700), .ZN(n13690) );
  NAND2_X1 U15709 ( .A1(n13691), .A2(n13690), .ZN(n13692) );
  XNOR2_X1 U15710 ( .A(n13692), .B(n13750), .ZN(n13696) );
  NAND2_X1 U15711 ( .A1(n14269), .A2(n13700), .ZN(n13694) );
  NAND2_X1 U15712 ( .A1(n14029), .A2(n13704), .ZN(n13693) );
  NAND2_X1 U15713 ( .A1(n13694), .A2(n13693), .ZN(n13695) );
  NOR2_X1 U15714 ( .A1(n13696), .A2(n13695), .ZN(n13697) );
  AOI21_X1 U15715 ( .B1(n13696), .B2(n13695), .A(n13697), .ZN(n13785) );
  NAND2_X1 U15716 ( .A1(n13784), .A2(n13785), .ZN(n13783) );
  INV_X1 U15717 ( .A(n13697), .ZN(n13698) );
  NAND2_X1 U15718 ( .A1(n14264), .A2(n13699), .ZN(n13702) );
  NAND2_X1 U15719 ( .A1(n13859), .A2(n13700), .ZN(n13701) );
  NAND2_X1 U15720 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  XNOR2_X1 U15721 ( .A(n13703), .B(n13750), .ZN(n13708) );
  NAND2_X1 U15722 ( .A1(n14264), .A2(n13608), .ZN(n13706) );
  NAND2_X1 U15723 ( .A1(n13859), .A2(n13704), .ZN(n13705) );
  NAND2_X1 U15724 ( .A1(n13706), .A2(n13705), .ZN(n13707) );
  NOR2_X1 U15725 ( .A1(n13708), .A2(n13707), .ZN(n13709) );
  AOI21_X1 U15726 ( .B1(n13708), .B2(n13707), .A(n13709), .ZN(n13838) );
  INV_X1 U15727 ( .A(n13709), .ZN(n13710) );
  OAI21_X1 U15728 ( .B1(n13712), .B2(n13711), .A(n13748), .ZN(n13713) );
  INV_X1 U15729 ( .A(n13713), .ZN(n13717) );
  OAI22_X1 U15730 ( .A1(n13786), .A2(n14127), .B1(n13753), .B2(n14617), .ZN(
        n14013) );
  AOI22_X1 U15731 ( .A1(n14013), .A2(n15299), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13714) );
  OAI21_X1 U15732 ( .B1(n15303), .B2(n14020), .A(n13714), .ZN(n13715) );
  AOI21_X1 U15733 ( .B1(n14022), .B2(n15311), .A(n13715), .ZN(n13716) );
  OAI21_X1 U15734 ( .B1(n13717), .B2(n15306), .A(n13716), .ZN(P1_U3214) );
  OAI21_X1 U15735 ( .B1(n13720), .B2(n13719), .A(n13718), .ZN(n13721) );
  NAND2_X1 U15736 ( .A1(n13721), .A2(n14532), .ZN(n13726) );
  NOR2_X1 U15737 ( .A1(n15303), .A2(n14228), .ZN(n13724) );
  OAI21_X1 U15738 ( .B1(n14510), .B2(n14508), .A(n13722), .ZN(n13723) );
  AOI211_X1 U15739 ( .C1(n14526), .C2(n14405), .A(n13724), .B(n13723), .ZN(
        n13725) );
  OAI211_X1 U15740 ( .C1(n14545), .C2(n14530), .A(n13726), .B(n13725), .ZN(
        P1_U3215) );
  OAI21_X1 U15741 ( .B1(n13729), .B2(n13728), .A(n13727), .ZN(n13735) );
  NAND2_X1 U15742 ( .A1(n14089), .A2(n14723), .ZN(n14281) );
  NOR2_X1 U15743 ( .A1(n14281), .A2(n13730), .ZN(n13734) );
  INV_X1 U15744 ( .A(n13862), .ZN(n13731) );
  INV_X1 U15745 ( .A(n13860), .ZN(n13787) );
  OAI22_X1 U15746 ( .A1(n13731), .A2(n14127), .B1(n13787), .B2(n14617), .ZN(
        n14079) );
  AOI22_X1 U15747 ( .A1(n14079), .A2(n15299), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13732) );
  OAI21_X1 U15748 ( .B1(n15303), .B2(n14087), .A(n13732), .ZN(n13733) );
  AOI211_X1 U15749 ( .C1(n13735), .C2(n14532), .A(n13734), .B(n13733), .ZN(
        n13736) );
  INV_X1 U15750 ( .A(n13736), .ZN(P1_U3216) );
  INV_X1 U15751 ( .A(n14299), .ZN(n14153) );
  INV_X1 U15752 ( .A(n13827), .ZN(n13739) );
  OAI21_X1 U15753 ( .B1(n13739), .B2(n13738), .A(n13737), .ZN(n13741) );
  NAND3_X1 U15754 ( .A1(n13741), .A2(n14532), .A3(n13740), .ZN(n13746) );
  NAND2_X1 U15755 ( .A1(n14144), .A2(n14528), .ZN(n13743) );
  OAI211_X1 U15756 ( .C1(n14509), .C2(n7100), .A(n13743), .B(n13742), .ZN(
        n13744) );
  AOI21_X1 U15757 ( .B1(n14150), .B2(n13843), .A(n13744), .ZN(n13745) );
  OAI211_X1 U15758 ( .C1(n14153), .C2(n14530), .A(n13746), .B(n13745), .ZN(
        P1_U3219) );
  OAI22_X1 U15759 ( .A1(n14006), .A2(n13752), .B1(n13753), .B2(n13749), .ZN(
        n13751) );
  XNOR2_X1 U15760 ( .A(n13751), .B(n13750), .ZN(n13756) );
  OAI22_X1 U15761 ( .A1(n14006), .A2(n13754), .B1(n13753), .B2(n13752), .ZN(
        n13755) );
  XNOR2_X1 U15762 ( .A(n13758), .B(n13757), .ZN(n13763) );
  AOI22_X1 U15763 ( .A1(n14526), .A2(n14030), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13760) );
  NAND2_X1 U15764 ( .A1(n14528), .A2(n13996), .ZN(n13759) );
  OAI211_X1 U15765 ( .C1(n15303), .C2(n14003), .A(n13760), .B(n13759), .ZN(
        n13761) );
  AOI21_X1 U15766 ( .B1(n14252), .B2(n15311), .A(n13761), .ZN(n13762) );
  OAI21_X1 U15767 ( .B1(n13763), .B2(n15306), .A(n13762), .ZN(P1_U3220) );
  OAI21_X1 U15768 ( .B1(n13766), .B2(n13765), .A(n13764), .ZN(n13767) );
  NAND2_X1 U15769 ( .A1(n13767), .A2(n14532), .ZN(n13771) );
  AOI22_X1 U15770 ( .A1(n14526), .A2(n13874), .B1(n14528), .B2(n13872), .ZN(
        n13770) );
  AOI22_X1 U15771 ( .A1(n15311), .A2(n9212), .B1(n13768), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n13769) );
  NAND3_X1 U15772 ( .A1(n13771), .A2(n13770), .A3(n13769), .ZN(P1_U3222) );
  INV_X1 U15773 ( .A(n13772), .ZN(n13773) );
  AOI21_X1 U15774 ( .B1(n13775), .B2(n13774), .A(n13773), .ZN(n13782) );
  INV_X1 U15775 ( .A(n14115), .ZN(n13779) );
  NAND2_X1 U15776 ( .A1(n14144), .A2(n14619), .ZN(n13777) );
  NAND2_X1 U15777 ( .A1(n13862), .A2(n14404), .ZN(n13776) );
  NAND2_X1 U15778 ( .A1(n13777), .A2(n13776), .ZN(n14112) );
  AOI22_X1 U15779 ( .A1(n14112), .A2(n15299), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13778) );
  OAI21_X1 U15780 ( .B1(n15303), .B2(n13779), .A(n13778), .ZN(n13780) );
  AOI21_X1 U15781 ( .B1(n14288), .B2(n15311), .A(n13780), .ZN(n13781) );
  OAI21_X1 U15782 ( .B1(n13782), .B2(n15306), .A(n13781), .ZN(P1_U3223) );
  OAI21_X1 U15783 ( .B1(n13785), .B2(n13784), .A(n13783), .ZN(n13791) );
  NAND2_X1 U15784 ( .A1(n14269), .A2(n15311), .ZN(n13789) );
  OAI22_X1 U15785 ( .A1(n13787), .A2(n14127), .B1(n13786), .B2(n14617), .ZN(
        n14047) );
  AOI22_X1 U15786 ( .A1(n14047), .A2(n15299), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13788) );
  OAI211_X1 U15787 ( .C1(n15303), .C2(n14049), .A(n13789), .B(n13788), .ZN(
        n13790) );
  AOI21_X1 U15788 ( .B1(n13791), .B2(n14532), .A(n13790), .ZN(n13792) );
  INV_X1 U15789 ( .A(n13792), .ZN(P1_U3225) );
  INV_X1 U15790 ( .A(n13793), .ZN(n13797) );
  NOR3_X1 U15791 ( .A1(n14512), .A2(n13795), .A3(n13794), .ZN(n13796) );
  OAI21_X1 U15792 ( .B1(n13797), .B2(n13796), .A(n14532), .ZN(n13802) );
  NOR2_X1 U15793 ( .A1(n15303), .A2(n14175), .ZN(n13800) );
  OAI21_X1 U15794 ( .B1(n14510), .B2(n7100), .A(n13798), .ZN(n13799) );
  AOI211_X1 U15795 ( .C1(n14526), .C2(n14182), .A(n13800), .B(n13799), .ZN(
        n13801) );
  OAI211_X1 U15796 ( .C1(n14311), .C2(n14530), .A(n13802), .B(n13801), .ZN(
        P1_U3228) );
  OAI21_X1 U15797 ( .B1(n13805), .B2(n13804), .A(n13803), .ZN(n13809) );
  NAND2_X1 U15798 ( .A1(n14274), .A2(n15311), .ZN(n13807) );
  INV_X1 U15799 ( .A(n14029), .ZN(n13841) );
  OAI22_X1 U15800 ( .A1(n13821), .A2(n14127), .B1(n13841), .B2(n14617), .ZN(
        n14062) );
  AOI22_X1 U15801 ( .A1(n14062), .A2(n15299), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13806) );
  OAI211_X1 U15802 ( .C1(n15303), .C2(n14069), .A(n13807), .B(n13806), .ZN(
        n13808) );
  AOI21_X1 U15803 ( .B1(n13809), .B2(n14532), .A(n13808), .ZN(n13810) );
  INV_X1 U15804 ( .A(n13810), .ZN(P1_U3229) );
  XNOR2_X1 U15805 ( .A(n13812), .B(n13811), .ZN(n13817) );
  AOI22_X1 U15806 ( .A1(n13863), .A2(n14528), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13814) );
  NAND2_X1 U15807 ( .A1(n13864), .A2(n14526), .ZN(n13813) );
  OAI211_X1 U15808 ( .C1(n15303), .C2(n14131), .A(n13814), .B(n13813), .ZN(
        n13815) );
  AOI21_X1 U15809 ( .B1(n14293), .B2(n15311), .A(n13815), .ZN(n13816) );
  OAI21_X1 U15810 ( .B1(n13817), .B2(n15306), .A(n13816), .ZN(P1_U3233) );
  OAI21_X1 U15811 ( .B1(n13820), .B2(n13819), .A(n13818), .ZN(n13825) );
  NAND2_X1 U15812 ( .A1(n14283), .A2(n15311), .ZN(n13823) );
  OAI22_X1 U15813 ( .A1(n14128), .A2(n14127), .B1(n13821), .B2(n14617), .ZN(
        n14104) );
  AOI22_X1 U15814 ( .A1(n14104), .A2(n15299), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13822) );
  OAI211_X1 U15815 ( .C1(n15303), .C2(n14097), .A(n13823), .B(n13822), .ZN(
        n13824) );
  AOI21_X1 U15816 ( .B1(n13825), .B2(n14532), .A(n13824), .ZN(n13826) );
  INV_X1 U15817 ( .A(n13826), .ZN(P1_U3235) );
  OAI21_X1 U15818 ( .B1(n13829), .B2(n13828), .A(n13827), .ZN(n13830) );
  NAND2_X1 U15819 ( .A1(n13830), .A2(n14532), .ZN(n13835) );
  NAND2_X1 U15820 ( .A1(n13864), .A2(n14528), .ZN(n13832) );
  OAI211_X1 U15821 ( .C1(n14509), .C2(n14511), .A(n13832), .B(n13831), .ZN(
        n13833) );
  AOI21_X1 U15822 ( .B1(n14167), .B2(n13843), .A(n13833), .ZN(n13834) );
  OAI211_X1 U15823 ( .C1(n7101), .C2(n14530), .A(n13835), .B(n13834), .ZN(
        P1_U3238) );
  OAI21_X1 U15824 ( .B1(n13838), .B2(n13837), .A(n13836), .ZN(n13839) );
  NAND2_X1 U15825 ( .A1(n13839), .A2(n14532), .ZN(n13846) );
  INV_X1 U15826 ( .A(n14035), .ZN(n13844) );
  AOI22_X1 U15827 ( .A1(n14528), .A2(n14030), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13840) );
  OAI21_X1 U15828 ( .B1(n13841), .B2(n14509), .A(n13840), .ZN(n13842) );
  AOI21_X1 U15829 ( .B1(n13844), .B2(n13843), .A(n13842), .ZN(n13845) );
  OAI211_X1 U15830 ( .C1(n13847), .C2(n14530), .A(n13846), .B(n13845), .ZN(
        P1_U3240) );
  XNOR2_X1 U15831 ( .A(n13849), .B(n13848), .ZN(n13855) );
  OAI22_X1 U15832 ( .A1(n13851), .A2(n14617), .B1(n13850), .B2(n14127), .ZN(
        n14204) );
  NAND2_X1 U15833 ( .A1(n14204), .A2(n15299), .ZN(n13852) );
  NAND2_X1 U15834 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14609)
         );
  OAI211_X1 U15835 ( .C1(n15303), .C2(n14211), .A(n13852), .B(n14609), .ZN(
        n13853) );
  AOI21_X1 U15836 ( .B1(n14214), .B2(n15311), .A(n13853), .ZN(n13854) );
  OAI21_X1 U15837 ( .B1(n13855), .B2(n15306), .A(n13854), .ZN(P1_U3241) );
  MUX2_X1 U15838 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13856), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15839 ( .A(n13857), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13878), .Z(
        P1_U3590) );
  MUX2_X1 U15840 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13996), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15841 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13858), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15842 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14030), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15843 ( .A(n13859), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13878), .Z(
        P1_U3586) );
  MUX2_X1 U15844 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14029), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15845 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13860), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15846 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13861), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15847 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13862), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15848 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13863), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15849 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14144), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15850 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13864), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15851 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14183), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15852 ( .A(n14195), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13878), .Z(
        P1_U3577) );
  MUX2_X1 U15853 ( .A(n14182), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13878), .Z(
        P1_U3576) );
  MUX2_X1 U15854 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14222), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15855 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13865), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15856 ( .A(n14405), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13878), .Z(
        P1_U3573) );
  MUX2_X1 U15857 ( .A(n14527), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13878), .Z(
        P1_U3572) );
  MUX2_X1 U15858 ( .A(n14406), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13878), .Z(
        P1_U3571) );
  MUX2_X1 U15859 ( .A(n14525), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13878), .Z(
        P1_U3570) );
  MUX2_X1 U15860 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13866), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15861 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13867), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15862 ( .A(n14620), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13878), .Z(
        P1_U3567) );
  MUX2_X1 U15863 ( .A(n13868), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13878), .Z(
        P1_U3566) );
  MUX2_X1 U15864 ( .A(n13869), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13878), .Z(
        P1_U3565) );
  MUX2_X1 U15865 ( .A(n13870), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13878), .Z(
        P1_U3564) );
  MUX2_X1 U15866 ( .A(n13871), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13878), .Z(
        P1_U3563) );
  MUX2_X1 U15867 ( .A(n13872), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13878), .Z(
        P1_U3562) );
  MUX2_X1 U15868 ( .A(n6936), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13878), .Z(
        P1_U3561) );
  MUX2_X1 U15869 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13874), .S(P1_U4016), .Z(
        P1_U3560) );
  MUX2_X1 U15870 ( .A(n13876), .B(n13875), .S(n6440), .Z(n13881) );
  OAI21_X1 U15871 ( .B1(n6440), .B2(P1_REG2_REG_0__SCAN_IN), .A(n13877), .ZN(
        n14591) );
  AOI21_X1 U15872 ( .B1(n13879), .B2(n14591), .A(n13878), .ZN(n13880) );
  OAI21_X1 U15873 ( .B1(n13881), .B2(n14344), .A(n13880), .ZN(n13933) );
  INV_X1 U15874 ( .A(n13890), .ZN(n13885) );
  OAI22_X1 U15875 ( .A1(n14611), .A2(n13883), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13882), .ZN(n13884) );
  AOI21_X1 U15876 ( .B1(n13885), .B2(n13964), .A(n13884), .ZN(n13897) );
  MUX2_X1 U15877 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9934), .S(n13890), .Z(
        n13886) );
  NAND3_X1 U15878 ( .A1(n13888), .A2(n13887), .A3(n13886), .ZN(n13889) );
  NAND3_X1 U15879 ( .A1(n14607), .A2(n13910), .A3(n13889), .ZN(n13896) );
  MUX2_X1 U15880 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9960), .S(n13890), .Z(
        n13891) );
  NAND3_X1 U15881 ( .A1(n13893), .A2(n13892), .A3(n13891), .ZN(n13894) );
  NAND3_X1 U15882 ( .A1(n13976), .A2(n13904), .A3(n13894), .ZN(n13895) );
  NAND4_X1 U15883 ( .A1(n13933), .A2(n13897), .A3(n13896), .A4(n13895), .ZN(
        P1_U3245) );
  INV_X1 U15884 ( .A(n13906), .ZN(n13901) );
  INV_X1 U15885 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n13899) );
  OAI21_X1 U15886 ( .B1(n14611), .B2(n13899), .A(n13898), .ZN(n13900) );
  AOI21_X1 U15887 ( .B1(n13901), .B2(n13964), .A(n13900), .ZN(n13914) );
  MUX2_X1 U15888 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10742), .S(n13906), .Z(
        n13902) );
  NAND3_X1 U15889 ( .A1(n13904), .A2(n13903), .A3(n13902), .ZN(n13905) );
  NAND3_X1 U15890 ( .A1(n13976), .A2(n13921), .A3(n13905), .ZN(n13913) );
  MUX2_X1 U15891 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n13907), .S(n13906), .Z(
        n13908) );
  NAND3_X1 U15892 ( .A1(n13910), .A2(n13909), .A3(n13908), .ZN(n13911) );
  NAND3_X1 U15893 ( .A1(n14607), .A2(n13916), .A3(n13911), .ZN(n13912) );
  NAND3_X1 U15894 ( .A1(n13914), .A2(n13913), .A3(n13912), .ZN(P1_U3246) );
  NAND2_X1 U15895 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n14594), .ZN(n13932) );
  MUX2_X1 U15896 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9928), .S(n13928), .Z(
        n13917) );
  NAND3_X1 U15897 ( .A1(n13917), .A2(n13916), .A3(n13915), .ZN(n13918) );
  NAND2_X1 U15898 ( .A1(n13919), .A2(n13918), .ZN(n13925) );
  MUX2_X1 U15899 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9954), .S(n13928), .Z(
        n13922) );
  NAND3_X1 U15900 ( .A1(n13922), .A2(n13921), .A3(n13920), .ZN(n13923) );
  NAND2_X1 U15901 ( .A1(n13944), .A2(n13923), .ZN(n13924) );
  OAI22_X1 U15902 ( .A1(n13926), .A2(n13925), .B1(n14604), .B2(n13924), .ZN(
        n13930) );
  OAI21_X1 U15903 ( .B1(n14602), .B2(n13928), .A(n13927), .ZN(n13929) );
  NOR2_X1 U15904 ( .A1(n13930), .A2(n13929), .ZN(n13931) );
  NAND3_X1 U15905 ( .A1(n13933), .A2(n13932), .A3(n13931), .ZN(P1_U3247) );
  OAI21_X1 U15906 ( .B1(n14611), .B2(n13935), .A(n13934), .ZN(n13936) );
  AOI21_X1 U15907 ( .B1(n13941), .B2(n13964), .A(n13936), .ZN(n13948) );
  OAI21_X1 U15908 ( .B1(n13939), .B2(n13938), .A(n13937), .ZN(n13940) );
  NAND2_X1 U15909 ( .A1(n14607), .A2(n13940), .ZN(n13947) );
  MUX2_X1 U15910 ( .A(n10643), .B(P1_REG2_REG_5__SCAN_IN), .S(n13941), .Z(
        n13942) );
  NAND3_X1 U15911 ( .A1(n13944), .A2(n13943), .A3(n13942), .ZN(n13945) );
  NAND3_X1 U15912 ( .A1(n13976), .A2(n13953), .A3(n13945), .ZN(n13946) );
  NAND3_X1 U15913 ( .A1(n13948), .A2(n13947), .A3(n13946), .ZN(P1_U3248) );
  NOR2_X1 U15914 ( .A1(n14602), .A2(n13951), .ZN(n13949) );
  AOI211_X1 U15915 ( .C1(n14594), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n13950), .B(
        n13949), .ZN(n13960) );
  MUX2_X1 U15916 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9968), .S(n13951), .Z(
        n13954) );
  NAND3_X1 U15917 ( .A1(n13954), .A2(n13953), .A3(n13952), .ZN(n13955) );
  NAND3_X1 U15918 ( .A1(n13976), .A2(n13973), .A3(n13955), .ZN(n13959) );
  OAI211_X1 U15919 ( .C1(n13957), .C2(n13956), .A(n14607), .B(n13967), .ZN(
        n13958) );
  NAND3_X1 U15920 ( .A1(n13960), .A2(n13959), .A3(n13958), .ZN(P1_U3249) );
  OAI21_X1 U15921 ( .B1(n14611), .B2(n13962), .A(n13961), .ZN(n13963) );
  AOI21_X1 U15922 ( .B1(n13970), .B2(n13964), .A(n13963), .ZN(n13979) );
  MUX2_X1 U15923 ( .A(n9942), .B(P1_REG1_REG_7__SCAN_IN), .S(n13970), .Z(
        n13965) );
  NAND3_X1 U15924 ( .A1(n13967), .A2(n13966), .A3(n13965), .ZN(n13968) );
  NAND3_X1 U15925 ( .A1(n14607), .A2(n13969), .A3(n13968), .ZN(n13978) );
  MUX2_X1 U15926 ( .A(n10805), .B(P1_REG2_REG_7__SCAN_IN), .S(n13970), .Z(
        n13971) );
  NAND3_X1 U15927 ( .A1(n13973), .A2(n13972), .A3(n13971), .ZN(n13974) );
  NAND3_X1 U15928 ( .A1(n13976), .A2(n13975), .A3(n13974), .ZN(n13977) );
  NAND3_X1 U15929 ( .A1(n13979), .A2(n13978), .A3(n13977), .ZN(P1_U3250) );
  XOR2_X1 U15930 ( .A(n14240), .B(n13986), .Z(n13980) );
  NAND2_X1 U15931 ( .A1(n13980), .A2(n14725), .ZN(n14239) );
  OR2_X1 U15932 ( .A1(n13982), .A2(n13981), .ZN(n14241) );
  NOR2_X1 U15933 ( .A1(n14625), .A2(n14241), .ZN(n13990) );
  NOR2_X1 U15934 ( .A1(n14240), .A2(n14190), .ZN(n13983) );
  AOI211_X1 U15935 ( .C1(n14625), .C2(P1_REG2_REG_31__SCAN_IN), .A(n13990), 
        .B(n13983), .ZN(n13984) );
  OAI21_X1 U15936 ( .B1(n14239), .B2(n14216), .A(n13984), .ZN(P1_U3263) );
  INV_X1 U15937 ( .A(n13985), .ZN(n13988) );
  INV_X1 U15938 ( .A(n13986), .ZN(n13987) );
  OAI211_X1 U15939 ( .C1(n14243), .C2(n13988), .A(n13987), .B(n14725), .ZN(
        n14242) );
  AND2_X1 U15940 ( .A1(n14656), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13989) );
  NOR2_X1 U15941 ( .A1(n13990), .A2(n13989), .ZN(n13993) );
  NAND2_X1 U15942 ( .A1(n13991), .A2(n14646), .ZN(n13992) );
  OAI211_X1 U15943 ( .C1(n14242), .C2(n14216), .A(n13993), .B(n13992), .ZN(
        P1_U3264) );
  XNOR2_X1 U15944 ( .A(n13995), .B(n13994), .ZN(n14000) );
  NAND2_X1 U15945 ( .A1(n13996), .A2(n14404), .ZN(n13998) );
  INV_X1 U15946 ( .A(n14001), .ZN(n14002) );
  AOI21_X1 U15947 ( .B1(n14252), .B2(n7182), .A(n14002), .ZN(n14253) );
  INV_X1 U15948 ( .A(n14003), .ZN(n14004) );
  AOI22_X1 U15949 ( .A1(n14625), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14004), 
        .B2(n14645), .ZN(n14005) );
  OAI21_X1 U15950 ( .B1(n14006), .B2(n14190), .A(n14005), .ZN(n14007) );
  AOI21_X1 U15951 ( .B1(n14253), .B2(n14652), .A(n14007), .ZN(n14011) );
  NAND3_X1 U15952 ( .A1(n14251), .A2(n14634), .A3(n14250), .ZN(n14010) );
  OAI211_X1 U15953 ( .C1(n14257), .C2(n14656), .A(n14011), .B(n14010), .ZN(
        P1_U3265) );
  XNOR2_X1 U15954 ( .A(n14012), .B(n9548), .ZN(n14014) );
  AOI21_X1 U15955 ( .B1(n14014), .B2(n14403), .A(n14013), .ZN(n14262) );
  OAI21_X1 U15956 ( .B1(n14016), .B2(n9548), .A(n14015), .ZN(n14260) );
  AND2_X1 U15957 ( .A1(n14022), .A2(n14038), .ZN(n14017) );
  OR2_X1 U15958 ( .A1(n14018), .A2(n14017), .ZN(n14258) );
  NAND2_X1 U15959 ( .A1(n14625), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n14019) );
  OAI21_X1 U15960 ( .B1(n14229), .B2(n14020), .A(n14019), .ZN(n14021) );
  AOI21_X1 U15961 ( .B1(n14022), .B2(n14646), .A(n14021), .ZN(n14023) );
  OAI21_X1 U15962 ( .B1(n14258), .B2(n14024), .A(n14023), .ZN(n14025) );
  AOI21_X1 U15963 ( .B1(n14260), .B2(n14634), .A(n14025), .ZN(n14026) );
  OAI21_X1 U15964 ( .B1(n14262), .B2(n14656), .A(n14026), .ZN(P1_U3266) );
  OAI21_X1 U15965 ( .B1(n14033), .B2(n14032), .A(n14031), .ZN(n14267) );
  NAND2_X1 U15966 ( .A1(n14625), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n14034) );
  OAI21_X1 U15967 ( .B1(n14229), .B2(n14035), .A(n14034), .ZN(n14036) );
  AOI21_X1 U15968 ( .B1(n14264), .B2(n14646), .A(n14036), .ZN(n14041) );
  INV_X1 U15969 ( .A(n14055), .ZN(n14037) );
  AOI21_X1 U15970 ( .B1(n14037), .B2(n14264), .A(n14715), .ZN(n14039) );
  AND2_X1 U15971 ( .A1(n14039), .A2(n14038), .ZN(n14263) );
  NAND2_X1 U15972 ( .A1(n14263), .A2(n14633), .ZN(n14040) );
  OAI211_X1 U15973 ( .C1(n14267), .C2(n14202), .A(n14041), .B(n14040), .ZN(
        n14042) );
  INV_X1 U15974 ( .A(n14042), .ZN(n14043) );
  OAI21_X1 U15975 ( .B1(n14266), .B2(n14656), .A(n14043), .ZN(P1_U3267) );
  OAI21_X1 U15976 ( .B1(n14046), .B2(n14045), .A(n14044), .ZN(n14048) );
  AOI21_X1 U15977 ( .B1(n14048), .B2(n14403), .A(n14047), .ZN(n14271) );
  OAI21_X1 U15978 ( .B1(n14049), .B2(n14229), .A(n14271), .ZN(n14059) );
  OAI21_X1 U15979 ( .B1(n14052), .B2(n14051), .A(n14050), .ZN(n14272) );
  AOI22_X1 U15980 ( .A1(n14269), .A2(n14646), .B1(n14625), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n14057) );
  NAND2_X1 U15981 ( .A1(n14269), .A2(n14073), .ZN(n14053) );
  NAND2_X1 U15982 ( .A1(n14053), .A2(n14725), .ZN(n14054) );
  NOR2_X1 U15983 ( .A1(n14055), .A2(n14054), .ZN(n14268) );
  NAND2_X1 U15984 ( .A1(n14268), .A2(n14633), .ZN(n14056) );
  OAI211_X1 U15985 ( .C1(n14272), .C2(n14202), .A(n14057), .B(n14056), .ZN(
        n14058) );
  AOI21_X1 U15986 ( .B1(n14059), .B2(n14231), .A(n14058), .ZN(n14060) );
  INV_X1 U15987 ( .A(n14060), .ZN(P1_U3268) );
  XNOR2_X1 U15988 ( .A(n14061), .B(n14065), .ZN(n14063) );
  AOI21_X1 U15989 ( .B1(n14063), .B2(n14403), .A(n14062), .ZN(n14276) );
  OAI21_X1 U15990 ( .B1(n14066), .B2(n14065), .A(n14064), .ZN(n14067) );
  INV_X1 U15991 ( .A(n14067), .ZN(n14277) );
  NAND2_X1 U15992 ( .A1(n14625), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n14068) );
  OAI21_X1 U15993 ( .B1(n14229), .B2(n14069), .A(n14068), .ZN(n14070) );
  AOI21_X1 U15994 ( .B1(n14274), .B2(n14646), .A(n14070), .ZN(n14075) );
  INV_X1 U15995 ( .A(n14071), .ZN(n14081) );
  AOI21_X1 U15996 ( .B1(n14274), .B2(n14081), .A(n14715), .ZN(n14072) );
  AND2_X1 U15997 ( .A1(n14073), .A2(n14072), .ZN(n14273) );
  NAND2_X1 U15998 ( .A1(n14273), .A2(n14633), .ZN(n14074) );
  OAI211_X1 U15999 ( .C1(n14277), .C2(n14202), .A(n14075), .B(n14074), .ZN(
        n14076) );
  INV_X1 U16000 ( .A(n14076), .ZN(n14077) );
  OAI21_X1 U16001 ( .B1(n14276), .B2(n14656), .A(n14077), .ZN(P1_U3269) );
  XNOR2_X1 U16002 ( .A(n14078), .B(n14084), .ZN(n14080) );
  AOI21_X1 U16003 ( .B1(n14080), .B2(n14403), .A(n14079), .ZN(n14282) );
  AOI21_X1 U16004 ( .B1(n14089), .B2(n14095), .A(n14715), .ZN(n14082) );
  NAND2_X1 U16005 ( .A1(n14082), .A2(n14081), .ZN(n14279) );
  NAND2_X1 U16006 ( .A1(n14085), .A2(n14084), .ZN(n14278) );
  NAND3_X1 U16007 ( .A1(n7429), .A2(n14278), .A3(n14634), .ZN(n14091) );
  NAND2_X1 U16008 ( .A1(n14625), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14086) );
  OAI21_X1 U16009 ( .B1(n14229), .B2(n14087), .A(n14086), .ZN(n14088) );
  AOI21_X1 U16010 ( .B1(n14089), .B2(n14646), .A(n14088), .ZN(n14090) );
  OAI211_X1 U16011 ( .C1(n14279), .C2(n14216), .A(n14091), .B(n14090), .ZN(
        n14092) );
  INV_X1 U16012 ( .A(n14092), .ZN(n14093) );
  OAI21_X1 U16013 ( .B1(n14282), .B2(n14656), .A(n14093), .ZN(P1_U3270) );
  XNOR2_X1 U16014 ( .A(n14094), .B(n14103), .ZN(n14287) );
  INV_X1 U16015 ( .A(n14095), .ZN(n14096) );
  AOI21_X1 U16016 ( .B1(n14283), .B2(n14114), .A(n14096), .ZN(n14284) );
  INV_X1 U16017 ( .A(n14097), .ZN(n14098) );
  AOI22_X1 U16018 ( .A1(n14625), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14098), 
        .B2(n14645), .ZN(n14099) );
  OAI21_X1 U16019 ( .B1(n14100), .B2(n14190), .A(n14099), .ZN(n14107) );
  OAI21_X1 U16020 ( .B1(n14103), .B2(n14102), .A(n14101), .ZN(n14105) );
  AOI21_X1 U16021 ( .B1(n14105), .B2(n14403), .A(n14104), .ZN(n14286) );
  NOR2_X1 U16022 ( .A1(n14286), .A2(n14656), .ZN(n14106) );
  AOI211_X1 U16023 ( .C1(n14284), .C2(n14652), .A(n14107), .B(n14106), .ZN(
        n14108) );
  OAI21_X1 U16024 ( .B1(n14287), .B2(n14202), .A(n14108), .ZN(P1_U3271) );
  AOI211_X1 U16025 ( .C1(n14111), .C2(n14110), .A(n14639), .B(n14109), .ZN(
        n14113) );
  NOR2_X1 U16026 ( .A1(n14113), .A2(n14112), .ZN(n14291) );
  AOI21_X1 U16027 ( .B1(n14288), .B2(n14136), .A(n7177), .ZN(n14289) );
  AOI22_X1 U16028 ( .A1(n14115), .A2(n14645), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n14625), .ZN(n14116) );
  OAI21_X1 U16029 ( .B1(n14117), .B2(n14190), .A(n14116), .ZN(n14123) );
  INV_X1 U16030 ( .A(n14118), .ZN(n14119) );
  AOI21_X1 U16031 ( .B1(n14121), .B2(n14120), .A(n14119), .ZN(n14292) );
  NOR2_X1 U16032 ( .A1(n14292), .A2(n14202), .ZN(n14122) );
  AOI211_X1 U16033 ( .C1(n14289), .C2(n14652), .A(n14123), .B(n14122), .ZN(
        n14124) );
  OAI21_X1 U16034 ( .B1(n14291), .B2(n14656), .A(n14124), .ZN(P1_U3272) );
  AOI211_X1 U16035 ( .C1(n14126), .C2(n14125), .A(n14639), .B(n6503), .ZN(
        n14130) );
  OAI22_X1 U16036 ( .A1(n14128), .A2(n14617), .B1(n14164), .B2(n14127), .ZN(
        n14129) );
  NOR2_X1 U16037 ( .A1(n14130), .A2(n14129), .ZN(n14298) );
  OAI21_X1 U16038 ( .B1(n14131), .B2(n14229), .A(n14298), .ZN(n14132) );
  NAND2_X1 U16039 ( .A1(n14132), .A2(n14231), .ZN(n14142) );
  AOI22_X1 U16040 ( .A1(n14293), .A2(n14646), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n14656), .ZN(n14141) );
  NAND2_X1 U16041 ( .A1(n14135), .A2(n14134), .ZN(n14295) );
  NAND3_X1 U16042 ( .A1(n14133), .A2(n14295), .A3(n14634), .ZN(n14140) );
  INV_X1 U16043 ( .A(n14149), .ZN(n14138) );
  INV_X1 U16044 ( .A(n14136), .ZN(n14137) );
  AOI21_X1 U16045 ( .B1(n14293), .B2(n14138), .A(n14137), .ZN(n14294) );
  NAND2_X1 U16046 ( .A1(n14294), .A2(n14652), .ZN(n14139) );
  NAND4_X1 U16047 ( .A1(n14142), .A2(n14141), .A3(n14140), .A4(n14139), .ZN(
        P1_U3273) );
  XNOR2_X1 U16048 ( .A(n14143), .B(n14147), .ZN(n14145) );
  AOI222_X1 U16049 ( .A1(n14403), .A2(n14145), .B1(n14144), .B2(n14404), .C1(
        n14183), .C2(n14619), .ZN(n14302) );
  XOR2_X1 U16050 ( .A(n14147), .B(n14146), .Z(n14303) );
  INV_X1 U16051 ( .A(n14303), .ZN(n14155) );
  AND2_X1 U16052 ( .A1(n14299), .A2(n14165), .ZN(n14148) );
  NOR2_X1 U16053 ( .A1(n14149), .A2(n14148), .ZN(n14300) );
  NAND2_X1 U16054 ( .A1(n14300), .A2(n14652), .ZN(n14152) );
  AOI22_X1 U16055 ( .A1(n14625), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14150), 
        .B2(n14645), .ZN(n14151) );
  OAI211_X1 U16056 ( .C1(n14153), .C2(n14190), .A(n14152), .B(n14151), .ZN(
        n14154) );
  AOI21_X1 U16057 ( .B1(n14155), .B2(n14634), .A(n14154), .ZN(n14156) );
  OAI21_X1 U16058 ( .B1(n14625), .B2(n14302), .A(n14156), .ZN(P1_U3274) );
  XNOR2_X1 U16059 ( .A(n14158), .B(n14157), .ZN(n14308) );
  OAI211_X1 U16060 ( .C1(n14161), .C2(n14160), .A(n14159), .B(n14403), .ZN(
        n14163) );
  NAND2_X1 U16061 ( .A1(n14195), .A2(n14619), .ZN(n14162) );
  OAI211_X1 U16062 ( .C1(n14164), .C2(n14617), .A(n14163), .B(n14162), .ZN(
        n14304) );
  INV_X1 U16063 ( .A(n14165), .ZN(n14166) );
  AOI211_X1 U16064 ( .C1(n14306), .C2(n14174), .A(n14715), .B(n14166), .ZN(
        n14305) );
  NAND2_X1 U16065 ( .A1(n14305), .A2(n14633), .ZN(n14169) );
  AOI22_X1 U16066 ( .A1(n14625), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14167), 
        .B2(n14645), .ZN(n14168) );
  OAI211_X1 U16067 ( .C1(n7101), .C2(n14190), .A(n14169), .B(n14168), .ZN(
        n14170) );
  AOI21_X1 U16068 ( .B1(n14304), .B2(n14231), .A(n14170), .ZN(n14171) );
  OAI21_X1 U16069 ( .B1(n14202), .B2(n14308), .A(n14171), .ZN(P1_U3275) );
  XNOR2_X1 U16070 ( .A(n14173), .B(n14172), .ZN(n14315) );
  OAI211_X1 U16071 ( .C1(n6554), .C2(n14311), .A(n14174), .B(n14725), .ZN(
        n14310) );
  OAI22_X1 U16072 ( .A1(n14231), .A2(n14176), .B1(n14175), .B2(n14229), .ZN(
        n14177) );
  AOI21_X1 U16073 ( .B1(n7184), .B2(n14646), .A(n14177), .ZN(n14178) );
  OAI21_X1 U16074 ( .B1(n14310), .B2(n14216), .A(n14178), .ZN(n14185) );
  OAI211_X1 U16075 ( .C1(n14181), .C2(n14180), .A(n14403), .B(n14179), .ZN(
        n14312) );
  AOI22_X1 U16076 ( .A1(n14183), .A2(n14404), .B1(n14182), .B2(n14619), .ZN(
        n14309) );
  AOI21_X1 U16077 ( .B1(n14312), .B2(n14309), .A(n14625), .ZN(n14184) );
  AOI211_X1 U16078 ( .C1(n14315), .C2(n14634), .A(n14185), .B(n14184), .ZN(
        n14186) );
  INV_X1 U16079 ( .A(n14186), .ZN(P1_U3276) );
  XNOR2_X1 U16080 ( .A(n14187), .B(n14193), .ZN(n14320) );
  AND2_X1 U16081 ( .A1(n14210), .A2(n14518), .ZN(n14188) );
  NOR2_X1 U16082 ( .A1(n6554), .A2(n14188), .ZN(n14317) );
  INV_X1 U16083 ( .A(n14518), .ZN(n14191) );
  OAI22_X1 U16084 ( .A1(n14191), .A2(n14190), .B1(n14189), .B2(n14231), .ZN(
        n14200) );
  OAI21_X1 U16085 ( .B1(n14194), .B2(n14193), .A(n14192), .ZN(n14196) );
  AOI222_X1 U16086 ( .A1(n14403), .A2(n14196), .B1(n14195), .B2(n14404), .C1(
        n14222), .C2(n14619), .ZN(n14319) );
  NAND2_X1 U16087 ( .A1(n14645), .A2(n14197), .ZN(n14198) );
  AOI21_X1 U16088 ( .B1(n14319), .B2(n14198), .A(n14656), .ZN(n14199) );
  AOI211_X1 U16089 ( .C1(n14317), .C2(n14652), .A(n14200), .B(n14199), .ZN(
        n14201) );
  OAI21_X1 U16090 ( .B1(n14202), .B2(n14320), .A(n14201), .ZN(P1_U3277) );
  AOI21_X1 U16091 ( .B1(n14203), .B2(n14208), .A(n14639), .ZN(n14206) );
  AOI21_X1 U16092 ( .B1(n14206), .B2(n14205), .A(n14204), .ZN(n14538) );
  OAI21_X1 U16093 ( .B1(n6567), .B2(n14208), .A(n14207), .ZN(n14540) );
  OAI211_X1 U16094 ( .C1(n9633), .C2(n14209), .A(n14725), .B(n14210), .ZN(
        n14537) );
  OAI22_X1 U16095 ( .A1(n14231), .A2(n14212), .B1(n14211), .B2(n14229), .ZN(
        n14213) );
  AOI21_X1 U16096 ( .B1(n14214), .B2(n14646), .A(n14213), .ZN(n14215) );
  OAI21_X1 U16097 ( .B1(n14537), .B2(n14216), .A(n14215), .ZN(n14217) );
  AOI21_X1 U16098 ( .B1(n14540), .B2(n14634), .A(n14217), .ZN(n14218) );
  OAI21_X1 U16099 ( .B1(n14625), .B2(n14538), .A(n14218), .ZN(P1_U3278) );
  XNOR2_X1 U16100 ( .A(n14220), .B(n14219), .ZN(n14221) );
  NAND2_X1 U16101 ( .A1(n14221), .A2(n14403), .ZN(n14224) );
  AOI22_X1 U16102 ( .A1(n14222), .A2(n14404), .B1(n14619), .B2(n14405), .ZN(
        n14223) );
  NAND2_X1 U16103 ( .A1(n14224), .A2(n14223), .ZN(n14546) );
  INV_X1 U16104 ( .A(n14225), .ZN(n14227) );
  OAI211_X1 U16105 ( .C1(n14545), .C2(n14227), .A(n14725), .B(n14226), .ZN(
        n14543) );
  OAI22_X1 U16106 ( .A1(n14543), .A2(n14230), .B1(n14229), .B2(n14228), .ZN(
        n14232) );
  OAI21_X1 U16107 ( .B1(n14546), .B2(n14232), .A(n14231), .ZN(n14238) );
  AOI22_X1 U16108 ( .A1(n14233), .A2(n14646), .B1(n14625), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n14237) );
  NAND2_X1 U16109 ( .A1(n14234), .A2(n14235), .ZN(n14541) );
  NAND3_X1 U16110 ( .A1(n14542), .A2(n14541), .A3(n14634), .ZN(n14236) );
  NAND3_X1 U16111 ( .A1(n14238), .A2(n14237), .A3(n14236), .ZN(P1_U3279) );
  OAI211_X1 U16112 ( .C1(n14240), .C2(n14743), .A(n14239), .B(n14241), .ZN(
        n14321) );
  MUX2_X1 U16113 ( .A(n14321), .B(P1_REG1_REG_31__SCAN_IN), .S(n14759), .Z(
        P1_U3559) );
  OAI211_X1 U16114 ( .C1(n14243), .C2(n14743), .A(n14242), .B(n14241), .ZN(
        n14322) );
  MUX2_X1 U16115 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14322), .S(n14761), .Z(
        P1_U3558) );
  AOI211_X1 U16116 ( .C1(n14247), .C2(n14723), .A(n14246), .B(n14245), .ZN(
        n14248) );
  NAND3_X1 U16117 ( .A1(n14251), .A2(n14250), .A3(n14748), .ZN(n14255) );
  AOI22_X1 U16118 ( .A1(n14253), .A2(n14725), .B1(n14252), .B2(n14723), .ZN(
        n14254) );
  MUX2_X1 U16119 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14323), .S(n14761), .Z(
        P1_U3556) );
  OAI22_X1 U16120 ( .A1(n14258), .A2(n14715), .B1(n7181), .B2(n14743), .ZN(
        n14259) );
  AOI21_X1 U16121 ( .B1(n14260), .B2(n14748), .A(n14259), .ZN(n14261) );
  NAND2_X1 U16122 ( .A1(n14262), .A2(n14261), .ZN(n14324) );
  MUX2_X1 U16123 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14324), .S(n14761), .Z(
        P1_U3555) );
  AOI21_X1 U16124 ( .B1(n14264), .B2(n14723), .A(n14263), .ZN(n14265) );
  OAI211_X1 U16125 ( .C1(n14703), .C2(n14267), .A(n14266), .B(n14265), .ZN(
        n14325) );
  MUX2_X1 U16126 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14325), .S(n14761), .Z(
        P1_U3554) );
  AOI21_X1 U16127 ( .B1(n14269), .B2(n14723), .A(n14268), .ZN(n14270) );
  OAI211_X1 U16128 ( .C1(n14703), .C2(n14272), .A(n14271), .B(n14270), .ZN(
        n14326) );
  MUX2_X1 U16129 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14326), .S(n14761), .Z(
        P1_U3553) );
  AOI21_X1 U16130 ( .B1(n14274), .B2(n14723), .A(n14273), .ZN(n14275) );
  OAI211_X1 U16131 ( .C1(n14703), .C2(n14277), .A(n14276), .B(n14275), .ZN(
        n14327) );
  MUX2_X1 U16132 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14327), .S(n14761), .Z(
        P1_U3552) );
  NAND3_X1 U16133 ( .A1(n7429), .A2(n14748), .A3(n14278), .ZN(n14280) );
  NAND4_X1 U16134 ( .A1(n14282), .A2(n14281), .A3(n14280), .A4(n14279), .ZN(
        n14328) );
  MUX2_X1 U16135 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14328), .S(n14761), .Z(
        P1_U3551) );
  AOI22_X1 U16136 ( .A1(n14284), .A2(n14725), .B1(n14283), .B2(n14723), .ZN(
        n14285) );
  OAI211_X1 U16137 ( .C1(n14703), .C2(n14287), .A(n14286), .B(n14285), .ZN(
        n14329) );
  MUX2_X1 U16138 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14329), .S(n14761), .Z(
        P1_U3550) );
  AOI22_X1 U16139 ( .A1(n14289), .A2(n14725), .B1(n14288), .B2(n14723), .ZN(
        n14290) );
  OAI211_X1 U16140 ( .C1(n14703), .C2(n14292), .A(n14291), .B(n14290), .ZN(
        n14330) );
  MUX2_X1 U16141 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14330), .S(n14761), .Z(
        P1_U3549) );
  AOI22_X1 U16142 ( .A1(n14294), .A2(n14725), .B1(n14293), .B2(n14723), .ZN(
        n14297) );
  NAND3_X1 U16143 ( .A1(n14133), .A2(n14295), .A3(n14748), .ZN(n14296) );
  NAND3_X1 U16144 ( .A1(n14298), .A2(n14297), .A3(n14296), .ZN(n14331) );
  MUX2_X1 U16145 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14331), .S(n14761), .Z(
        P1_U3548) );
  AOI22_X1 U16146 ( .A1(n14300), .A2(n14725), .B1(n14299), .B2(n14723), .ZN(
        n14301) );
  OAI211_X1 U16147 ( .C1(n14703), .C2(n14303), .A(n14302), .B(n14301), .ZN(
        n14332) );
  MUX2_X1 U16148 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14332), .S(n14761), .Z(
        P1_U3547) );
  AOI211_X1 U16149 ( .C1(n14306), .C2(n14723), .A(n14305), .B(n14304), .ZN(
        n14307) );
  OAI21_X1 U16150 ( .B1(n14703), .B2(n14308), .A(n14307), .ZN(n14333) );
  MUX2_X1 U16151 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14333), .S(n14761), .Z(
        P1_U3546) );
  OAI211_X1 U16152 ( .C1(n14311), .C2(n14743), .A(n14310), .B(n14309), .ZN(
        n14314) );
  INV_X1 U16153 ( .A(n14312), .ZN(n14313) );
  AOI211_X1 U16154 ( .C1(n14315), .C2(n14748), .A(n14314), .B(n14313), .ZN(
        n14316) );
  INV_X1 U16155 ( .A(n14316), .ZN(n14334) );
  MUX2_X1 U16156 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14334), .S(n14761), .Z(
        P1_U3545) );
  AOI22_X1 U16157 ( .A1(n14317), .A2(n14725), .B1(n14518), .B2(n14723), .ZN(
        n14318) );
  OAI211_X1 U16158 ( .C1(n14703), .C2(n14320), .A(n14319), .B(n14318), .ZN(
        n14335) );
  MUX2_X1 U16159 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14335), .S(n14761), .Z(
        P1_U3544) );
  MUX2_X1 U16160 ( .A(n14321), .B(P1_REG0_REG_31__SCAN_IN), .S(n14749), .Z(
        P1_U3527) );
  MUX2_X1 U16161 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14322), .S(n14751), .Z(
        P1_U3526) );
  MUX2_X1 U16162 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14323), .S(n14751), .Z(
        P1_U3524) );
  MUX2_X1 U16163 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14324), .S(n14751), .Z(
        P1_U3523) );
  MUX2_X1 U16164 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14325), .S(n14751), .Z(
        P1_U3522) );
  MUX2_X1 U16165 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14326), .S(n14751), .Z(
        P1_U3521) );
  MUX2_X1 U16166 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14327), .S(n14751), .Z(
        P1_U3520) );
  MUX2_X1 U16167 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14328), .S(n14751), .Z(
        P1_U3519) );
  MUX2_X1 U16168 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14329), .S(n14751), .Z(
        P1_U3518) );
  MUX2_X1 U16169 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14330), .S(n14751), .Z(
        P1_U3517) );
  MUX2_X1 U16170 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14331), .S(n14751), .Z(
        P1_U3516) );
  MUX2_X1 U16171 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14332), .S(n14751), .Z(
        P1_U3515) );
  MUX2_X1 U16172 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14333), .S(n14751), .Z(
        P1_U3513) );
  MUX2_X1 U16173 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14334), .S(n14751), .Z(
        P1_U3510) );
  MUX2_X1 U16174 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14335), .S(n14751), .Z(
        P1_U3507) );
  INV_X1 U16175 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14336) );
  NAND3_X1 U16176 ( .A1(n14336), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n14338) );
  OAI22_X1 U16177 ( .A1(n14339), .A2(n14338), .B1(n14337), .B2(n14353), .ZN(
        n14340) );
  AOI21_X1 U16178 ( .B1(n14342), .B2(n14341), .A(n14340), .ZN(n14343) );
  INV_X1 U16179 ( .A(n14343), .ZN(P1_U3324) );
  OAI222_X1 U16180 ( .A1(n14353), .A2(n14346), .B1(n11585), .B2(n14345), .C1(
        P1_U3086), .C2(n14344), .ZN(P1_U3327) );
  OAI222_X1 U16181 ( .A1(n11585), .A2(n14349), .B1(P1_U3086), .B2(n14348), 
        .C1(n14347), .C2(n14353), .ZN(P1_U3329) );
  INV_X1 U16182 ( .A(n14350), .ZN(n14351) );
  OAI222_X1 U16183 ( .A1(n14353), .A2(n15215), .B1(n11585), .B2(n14352), .C1(
        n14351), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI222_X1 U16184 ( .A1(n11585), .A2(n14356), .B1(P1_U3086), .B2(n14355), 
        .C1(n14354), .C2(n14353), .ZN(P1_U3331) );
  MUX2_X1 U16185 ( .A(n14358), .B(n14357), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16186 ( .A(n14359), .ZN(n14360) );
  MUX2_X1 U16187 ( .A(n14360), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U16188 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14364) );
  OAI21_X1 U16189 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14364), 
        .ZN(U28) );
  AOI21_X1 U16190 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14365) );
  OAI21_X1 U16191 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14365), 
        .ZN(U29) );
  INV_X1 U16192 ( .A(n14366), .ZN(n14370) );
  INV_X1 U16193 ( .A(n15325), .ZN(n14369) );
  AOI21_X1 U16194 ( .B1(n14367), .B2(n14370), .A(P2_ADDR_REG_2__SCAN_IN), .ZN(
        n14368) );
  AOI21_X1 U16195 ( .B1(n14370), .B2(n14369), .A(n14368), .ZN(SUB_1596_U61) );
  AOI22_X1 U16196 ( .A1(n14371), .A2(n14388), .B1(SI_9_), .B2(n14387), .ZN(
        n14372) );
  OAI21_X1 U16197 ( .B1(P3_U3151), .B2(n14990), .A(n14372), .ZN(P3_U3286) );
  AOI22_X1 U16198 ( .A1(n14373), .A2(n14388), .B1(SI_11_), .B2(n14387), .ZN(
        n14374) );
  OAI21_X1 U16199 ( .B1(P3_U3151), .B2(n14375), .A(n14374), .ZN(P3_U3284) );
  OAI22_X1 U16200 ( .A1(n14379), .A2(n14378), .B1(n14377), .B2(n14376), .ZN(
        n14380) );
  INV_X1 U16201 ( .A(n14380), .ZN(n14381) );
  OAI21_X1 U16202 ( .B1(P3_U3151), .B2(n14382), .A(n14381), .ZN(P3_U3282) );
  AOI21_X1 U16203 ( .B1(n14385), .B2(n14384), .A(n14383), .ZN(SUB_1596_U57) );
  INV_X1 U16204 ( .A(n14386), .ZN(n14389) );
  AOI22_X1 U16205 ( .A1(n14389), .A2(n14388), .B1(SI_15_), .B2(n14387), .ZN(
        n14390) );
  OAI21_X1 U16206 ( .B1(P3_U3151), .B2(n14391), .A(n14390), .ZN(P3_U3280) );
  OAI21_X1 U16207 ( .B1(n14393), .B2(n14828), .A(n14392), .ZN(SUB_1596_U55) );
  AOI21_X1 U16208 ( .B1(n14849), .B2(n14395), .A(n14394), .ZN(SUB_1596_U54) );
  AOI21_X1 U16209 ( .B1(n14398), .B2(n14397), .A(n14396), .ZN(SUB_1596_U70) );
  XNOR2_X1 U16210 ( .A(n14399), .B(n14400), .ZN(n14422) );
  XNOR2_X1 U16211 ( .A(n14401), .B(n14400), .ZN(n14402) );
  AOI222_X1 U16212 ( .A1(n14406), .A2(n14619), .B1(n14405), .B2(n14404), .C1(
        n14403), .C2(n14402), .ZN(n14420) );
  INV_X1 U16213 ( .A(n14420), .ZN(n14407) );
  AOI21_X1 U16214 ( .B1(n14733), .B2(n14422), .A(n14407), .ZN(n14418) );
  INV_X1 U16215 ( .A(n14408), .ZN(n14409) );
  AOI222_X1 U16216 ( .A1(n14410), .A2(n14646), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14656), .C1(n14645), .C2(n14409), .ZN(n14417) );
  INV_X1 U16217 ( .A(n14411), .ZN(n14653) );
  INV_X1 U16218 ( .A(n14412), .ZN(n14414) );
  OAI211_X1 U16219 ( .C1(n14414), .C2(n7185), .A(n14725), .B(n14413), .ZN(
        n14419) );
  INV_X1 U16220 ( .A(n14419), .ZN(n14415) );
  AOI22_X1 U16221 ( .A1(n14422), .A2(n14653), .B1(n14633), .B2(n14415), .ZN(
        n14416) );
  OAI211_X1 U16222 ( .C1(n14656), .C2(n14418), .A(n14417), .B(n14416), .ZN(
        P1_U3281) );
  OAI211_X1 U16223 ( .C1(n7185), .C2(n14743), .A(n14420), .B(n14419), .ZN(
        n14421) );
  AOI21_X1 U16224 ( .B1(n14422), .B2(n14748), .A(n14421), .ZN(n14425) );
  INV_X1 U16225 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14423) );
  AOI22_X1 U16226 ( .A1(n14751), .A2(n14425), .B1(n14423), .B2(n14749), .ZN(
        P1_U3495) );
  AOI22_X1 U16227 ( .A1(n14761), .A2(n14425), .B1(n14424), .B2(n14759), .ZN(
        P1_U3540) );
  AOI21_X1 U16228 ( .B1(n14428), .B2(n14427), .A(n14426), .ZN(n14429) );
  XOR2_X1 U16229 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14429), .Z(SUB_1596_U63)
         );
  AOI21_X1 U16230 ( .B1(n14432), .B2(n14431), .A(n14430), .ZN(n14446) );
  OAI21_X1 U16231 ( .B1(n14434), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14433), 
        .ZN(n14444) );
  NAND2_X1 U16232 ( .A1(n15017), .A2(n14435), .ZN(n14437) );
  OAI211_X1 U16233 ( .C1(n14438), .C2(n15024), .A(n14437), .B(n14436), .ZN(
        n14443) );
  AOI211_X1 U16234 ( .C1(n14441), .C2(n14440), .A(n14991), .B(n14439), .ZN(
        n14442) );
  AOI211_X1 U16235 ( .C1(n15007), .C2(n14444), .A(n14443), .B(n14442), .ZN(
        n14445) );
  OAI21_X1 U16236 ( .B1(n14446), .B2(n15001), .A(n14445), .ZN(P3_U3199) );
  NOR2_X1 U16237 ( .A1(n14989), .A2(n14449), .ZN(n14450) );
  AOI211_X1 U16238 ( .C1(n14995), .C2(P3_ADDR_REG_18__SCAN_IN), .A(n14451), 
        .B(n14450), .ZN(n14461) );
  AOI21_X1 U16239 ( .B1(n14454), .B2(n14453), .A(n14452), .ZN(n14455) );
  INV_X1 U16240 ( .A(n14455), .ZN(n14459) );
  XNOR2_X1 U16241 ( .A(n14457), .B(n14456), .ZN(n14458) );
  AOI22_X1 U16242 ( .A1(n14459), .A2(n15015), .B1(n15007), .B2(n14458), .ZN(
        n14460) );
  AOI22_X1 U16243 ( .A1(n14478), .A2(n14462), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15093), .ZN(n14463) );
  NAND2_X1 U16244 ( .A1(n14464), .A2(n14463), .ZN(P3_U3203) );
  XNOR2_X1 U16245 ( .A(n14465), .B(n14466), .ZN(n14469) );
  AOI222_X1 U16246 ( .A1(n15072), .A2(n14469), .B1(n14468), .B2(n15066), .C1(
        n14467), .C2(n15069), .ZN(n14483) );
  AOI22_X1 U16247 ( .A1(n15053), .A2(n14470), .B1(P3_REG2_REG_11__SCAN_IN), 
        .B2(n15093), .ZN(n14475) );
  XNOR2_X1 U16248 ( .A(n14472), .B(n14471), .ZN(n14486) );
  NOR2_X1 U16249 ( .A1(n14473), .A2(n15111), .ZN(n14485) );
  AOI22_X1 U16250 ( .A1(n14486), .A2(n15059), .B1(n15058), .B2(n14485), .ZN(
        n14474) );
  OAI211_X1 U16251 ( .C1(n15093), .C2(n14483), .A(n14475), .B(n14474), .ZN(
        P3_U3222) );
  AOI21_X1 U16252 ( .B1(n14478), .B2(n14477), .A(n14476), .ZN(n14487) );
  AOI22_X1 U16253 ( .A1(n15149), .A2(n14487), .B1(n15240), .B2(n15147), .ZN(
        P3_U3489) );
  NOR2_X1 U16254 ( .A1(n14479), .A2(n15111), .ZN(n14481) );
  AOI211_X1 U16255 ( .C1(n14482), .C2(n15102), .A(n14481), .B(n14480), .ZN(
        n14489) );
  AOI22_X1 U16256 ( .A1(n15149), .A2(n14489), .B1(n11257), .B2(n15147), .ZN(
        P3_U3471) );
  INV_X1 U16257 ( .A(n14483), .ZN(n14484) );
  AOI211_X1 U16258 ( .C1(n15102), .C2(n14486), .A(n14485), .B(n14484), .ZN(
        n14491) );
  AOI22_X1 U16259 ( .A1(n15149), .A2(n14491), .B1(n7845), .B2(n15147), .ZN(
        P3_U3470) );
  INV_X1 U16260 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U16261 ( .A1(n15137), .A2(n14488), .B1(n14487), .B2(n15136), .ZN(
        P3_U3457) );
  INV_X1 U16262 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14490) );
  AOI22_X1 U16263 ( .A1(n15137), .A2(n14490), .B1(n14489), .B2(n15136), .ZN(
        P3_U3426) );
  INV_X1 U16264 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U16265 ( .A1(n15137), .A2(n14492), .B1(n14491), .B2(n15136), .ZN(
        P3_U3423) );
  OAI21_X1 U16266 ( .B1(n14494), .B2(n14953), .A(n14493), .ZN(n14496) );
  AOI211_X1 U16267 ( .C1(n14918), .C2(n14497), .A(n14496), .B(n14495), .ZN(
        n14505) );
  AOI22_X1 U16268 ( .A1(n14974), .A2(n14505), .B1(n10628), .B2(n14971), .ZN(
        P2_U3513) );
  INV_X1 U16269 ( .A(n14923), .ZN(n14957) );
  INV_X1 U16270 ( .A(n14498), .ZN(n14503) );
  OAI21_X1 U16271 ( .B1(n14500), .B2(n14953), .A(n14499), .ZN(n14502) );
  AOI211_X1 U16272 ( .C1(n14957), .C2(n14503), .A(n14502), .B(n14501), .ZN(
        n14507) );
  AOI22_X1 U16273 ( .A1(n14974), .A2(n14507), .B1(n10206), .B2(n14971), .ZN(
        P2_U3511) );
  INV_X1 U16274 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14504) );
  AOI22_X1 U16275 ( .A1(n14959), .A2(n14505), .B1(n14504), .B2(n14958), .ZN(
        P2_U3472) );
  INV_X1 U16276 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U16277 ( .A1(n14959), .A2(n14507), .B1(n14506), .B2(n14958), .ZN(
        P2_U3466) );
  OAI22_X1 U16278 ( .A1(n14511), .A2(n14510), .B1(n14509), .B2(n14508), .ZN(
        n14517) );
  AOI21_X1 U16279 ( .B1(n14514), .B2(n14513), .A(n14512), .ZN(n14515) );
  NOR2_X1 U16280 ( .A1(n14515), .A2(n15306), .ZN(n14516) );
  AOI211_X1 U16281 ( .C1(n15311), .C2(n14518), .A(n14517), .B(n14516), .ZN(
        n14520) );
  OAI211_X1 U16282 ( .C1(n15303), .C2(n14521), .A(n14520), .B(n14519), .ZN(
        P1_U3226) );
  OAI21_X1 U16283 ( .B1(n14524), .B2(n14523), .A(n14522), .ZN(n14533) );
  AOI22_X1 U16284 ( .A1(n14528), .A2(n14527), .B1(n14526), .B2(n14525), .ZN(
        n14529) );
  OAI21_X1 U16285 ( .B1(n14554), .B2(n14530), .A(n14529), .ZN(n14531) );
  AOI21_X1 U16286 ( .B1(n14533), .B2(n14532), .A(n14531), .ZN(n14535) );
  OAI211_X1 U16287 ( .C1(n15303), .C2(n14536), .A(n14535), .B(n14534), .ZN(
        P1_U3236) );
  OAI211_X1 U16288 ( .C1(n9633), .C2(n14743), .A(n14538), .B(n14537), .ZN(
        n14539) );
  AOI21_X1 U16289 ( .B1(n14540), .B2(n14748), .A(n14539), .ZN(n14559) );
  AOI22_X1 U16290 ( .A1(n14761), .A2(n14559), .B1(n9395), .B2(n14759), .ZN(
        P1_U3543) );
  NAND3_X1 U16291 ( .A1(n14542), .A2(n14541), .A3(n14748), .ZN(n14544) );
  OAI211_X1 U16292 ( .C1(n14545), .C2(n14743), .A(n14544), .B(n14543), .ZN(
        n14547) );
  NOR2_X1 U16293 ( .A1(n14547), .A2(n14546), .ZN(n14561) );
  AOI22_X1 U16294 ( .A1(n14761), .A2(n14561), .B1(n10710), .B2(n14759), .ZN(
        P1_U3542) );
  OAI211_X1 U16295 ( .C1(n14550), .C2(n14743), .A(n14549), .B(n14548), .ZN(
        n14551) );
  AOI21_X1 U16296 ( .B1(n14552), .B2(n14748), .A(n14551), .ZN(n14563) );
  AOI22_X1 U16297 ( .A1(n14761), .A2(n14563), .B1(n9366), .B2(n14759), .ZN(
        P1_U3541) );
  OAI21_X1 U16298 ( .B1(n14554), .B2(n14743), .A(n14553), .ZN(n14556) );
  AOI211_X1 U16299 ( .C1(n14557), .C2(n14748), .A(n14556), .B(n14555), .ZN(
        n14565) );
  AOI22_X1 U16300 ( .A1(n14761), .A2(n14565), .B1(n10034), .B2(n14759), .ZN(
        P1_U3539) );
  INV_X1 U16301 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14558) );
  AOI22_X1 U16302 ( .A1(n14751), .A2(n14559), .B1(n14558), .B2(n14749), .ZN(
        P1_U3504) );
  INV_X1 U16303 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14560) );
  AOI22_X1 U16304 ( .A1(n14751), .A2(n14561), .B1(n14560), .B2(n14749), .ZN(
        P1_U3501) );
  INV_X1 U16305 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14562) );
  AOI22_X1 U16306 ( .A1(n14751), .A2(n14563), .B1(n14562), .B2(n14749), .ZN(
        P1_U3498) );
  INV_X1 U16307 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14564) );
  AOI22_X1 U16308 ( .A1(n14751), .A2(n14565), .B1(n14564), .B2(n14749), .ZN(
        P1_U3492) );
  AOI21_X1 U16309 ( .B1(n14568), .B2(n14567), .A(n14566), .ZN(n14569) );
  XOR2_X1 U16310 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14569), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16311 ( .B1(n14571), .B2(n14570), .A(n6573), .ZN(n14572) );
  XOR2_X1 U16312 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14572), .Z(SUB_1596_U68)
         );
  OAI21_X1 U16313 ( .B1(n14575), .B2(n14574), .A(n14573), .ZN(n14576) );
  XNOR2_X1 U16314 ( .A(n14576), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16315 ( .B1(n14579), .B2(n14578), .A(n14577), .ZN(n14580) );
  XNOR2_X1 U16316 ( .A(n14580), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16317 ( .A1(n14585), .A2(n14584), .B1(n14585), .B2(n14583), .C1(
        n14582), .C2(n14581), .ZN(SUB_1596_U65) );
  INV_X1 U16318 ( .A(n14588), .ZN(n14587) );
  OAI222_X1 U16319 ( .A1(n14590), .A2(n14589), .B1(n14590), .B2(n14588), .C1(
        n14587), .C2(n14586), .ZN(SUB_1596_U64) );
  AOI21_X1 U16320 ( .B1(n6440), .B2(n14592), .A(n14591), .ZN(n14593) );
  XNOR2_X1 U16321 ( .A(n14593), .B(P1_IR_REG_0__SCAN_IN), .ZN(n14597) );
  AOI22_X1 U16322 ( .A1(n14594), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14595) );
  OAI21_X1 U16323 ( .B1(n14597), .B2(n14596), .A(n14595), .ZN(P1_U3243) );
  INV_X1 U16324 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14612) );
  OAI21_X1 U16325 ( .B1(n14599), .B2(n9395), .A(n14598), .ZN(n14608) );
  AOI21_X1 U16326 ( .B1(n14601), .B2(P1_REG2_REG_15__SCAN_IN), .A(n14600), 
        .ZN(n14605) );
  OAI22_X1 U16327 ( .A1(n14605), .A2(n14604), .B1(n14603), .B2(n14602), .ZN(
        n14606) );
  AOI21_X1 U16328 ( .B1(n14608), .B2(n14607), .A(n14606), .ZN(n14610) );
  OAI211_X1 U16329 ( .C1(n14612), .C2(n14611), .A(n14610), .B(n14609), .ZN(
        P1_U3258) );
  INV_X1 U16330 ( .A(n14613), .ZN(n14614) );
  NOR2_X1 U16331 ( .A1(n14615), .A2(n14614), .ZN(n14616) );
  AOI21_X1 U16332 ( .B1(n10801), .B2(n14616), .A(n14639), .ZN(n14623) );
  OR2_X1 U16333 ( .A1(n14618), .A2(n14617), .ZN(n14622) );
  NAND2_X1 U16334 ( .A1(n14620), .A2(n14619), .ZN(n14621) );
  NAND2_X1 U16335 ( .A1(n14622), .A2(n14621), .ZN(n15300) );
  AOI21_X1 U16336 ( .B1(n14624), .B2(n14623), .A(n15300), .ZN(n14736) );
  INV_X1 U16337 ( .A(n15302), .ZN(n14626) );
  AOI222_X1 U16338 ( .A1(n15310), .A2(n14646), .B1(n14626), .B2(n14645), .C1(
        P1_REG2_REG_8__SCAN_IN), .C2(n14625), .ZN(n14636) );
  XNOR2_X1 U16339 ( .A(n14627), .B(n14628), .ZN(n14739) );
  INV_X1 U16340 ( .A(n14629), .ZN(n14630) );
  OAI211_X1 U16341 ( .C1(n14737), .C2(n14631), .A(n14630), .B(n14725), .ZN(
        n14735) );
  INV_X1 U16342 ( .A(n14735), .ZN(n14632) );
  AOI22_X1 U16343 ( .A1(n14739), .A2(n14634), .B1(n14633), .B2(n14632), .ZN(
        n14635) );
  OAI211_X1 U16344 ( .C1(n14656), .C2(n14736), .A(n14636), .B(n14635), .ZN(
        P1_U3285) );
  XNOR2_X1 U16345 ( .A(n14637), .B(n6438), .ZN(n14720) );
  XNOR2_X1 U16346 ( .A(n14638), .B(n6438), .ZN(n14640) );
  NOR2_X1 U16347 ( .A1(n14640), .A2(n14639), .ZN(n14641) );
  AOI211_X1 U16348 ( .C1(n14733), .C2(n14720), .A(n14642), .B(n14641), .ZN(
        n14717) );
  INV_X1 U16349 ( .A(n14643), .ZN(n14644) );
  AOI222_X1 U16350 ( .A1(n14647), .A2(n14646), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n14656), .C1(n14645), .C2(n14644), .ZN(n14655) );
  INV_X1 U16351 ( .A(n14647), .ZN(n14649) );
  OAI21_X1 U16352 ( .B1(n14650), .B2(n14649), .A(n14648), .ZN(n14716) );
  INV_X1 U16353 ( .A(n14716), .ZN(n14651) );
  AOI22_X1 U16354 ( .A1(n14720), .A2(n14653), .B1(n14652), .B2(n14651), .ZN(
        n14654) );
  OAI211_X1 U16355 ( .C1(n14656), .C2(n14717), .A(n14655), .B(n14654), .ZN(
        P1_U3287) );
  NOR2_X1 U16356 ( .A1(n14684), .A2(n15214), .ZN(P1_U3294) );
  INV_X1 U16357 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14657) );
  NOR2_X1 U16358 ( .A1(n14684), .A2(n14657), .ZN(P1_U3295) );
  INV_X1 U16359 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14658) );
  NOR2_X1 U16360 ( .A1(n14684), .A2(n14658), .ZN(P1_U3296) );
  INV_X1 U16361 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14659) );
  NOR2_X1 U16362 ( .A1(n14684), .A2(n14659), .ZN(P1_U3297) );
  INV_X1 U16363 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14660) );
  NOR2_X1 U16364 ( .A1(n14684), .A2(n14660), .ZN(P1_U3298) );
  INV_X1 U16365 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14661) );
  NOR2_X1 U16366 ( .A1(n14684), .A2(n14661), .ZN(P1_U3299) );
  INV_X1 U16367 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14662) );
  NOR2_X1 U16368 ( .A1(n14684), .A2(n14662), .ZN(P1_U3300) );
  NOR2_X1 U16369 ( .A1(n14684), .A2(n15243), .ZN(P1_U3301) );
  INV_X1 U16370 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14663) );
  NOR2_X1 U16371 ( .A1(n14684), .A2(n14663), .ZN(P1_U3302) );
  INV_X1 U16372 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14664) );
  NOR2_X1 U16373 ( .A1(n14684), .A2(n14664), .ZN(P1_U3303) );
  NOR2_X1 U16374 ( .A1(n14684), .A2(n15193), .ZN(P1_U3304) );
  INV_X1 U16375 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14665) );
  NOR2_X1 U16376 ( .A1(n14684), .A2(n14665), .ZN(P1_U3305) );
  INV_X1 U16377 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14666) );
  NOR2_X1 U16378 ( .A1(n14684), .A2(n14666), .ZN(P1_U3306) );
  INV_X1 U16379 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14667) );
  NOR2_X1 U16380 ( .A1(n14684), .A2(n14667), .ZN(P1_U3307) );
  INV_X1 U16381 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14668) );
  NOR2_X1 U16382 ( .A1(n14684), .A2(n14668), .ZN(P1_U3308) );
  INV_X1 U16383 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14669) );
  NOR2_X1 U16384 ( .A1(n14684), .A2(n14669), .ZN(P1_U3309) );
  INV_X1 U16385 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14670) );
  NOR2_X1 U16386 ( .A1(n14684), .A2(n14670), .ZN(P1_U3310) );
  INV_X1 U16387 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14671) );
  NOR2_X1 U16388 ( .A1(n14684), .A2(n14671), .ZN(P1_U3311) );
  INV_X1 U16389 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14672) );
  NOR2_X1 U16390 ( .A1(n14684), .A2(n14672), .ZN(P1_U3312) );
  INV_X1 U16391 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14673) );
  NOR2_X1 U16392 ( .A1(n14684), .A2(n14673), .ZN(P1_U3313) );
  INV_X1 U16393 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14674) );
  NOR2_X1 U16394 ( .A1(n14684), .A2(n14674), .ZN(P1_U3314) );
  INV_X1 U16395 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14675) );
  NOR2_X1 U16396 ( .A1(n14684), .A2(n14675), .ZN(P1_U3315) );
  INV_X1 U16397 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14676) );
  NOR2_X1 U16398 ( .A1(n14684), .A2(n14676), .ZN(P1_U3316) );
  INV_X1 U16399 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14677) );
  NOR2_X1 U16400 ( .A1(n14684), .A2(n14677), .ZN(P1_U3317) );
  INV_X1 U16401 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14678) );
  NOR2_X1 U16402 ( .A1(n14684), .A2(n14678), .ZN(P1_U3318) );
  INV_X1 U16403 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14679) );
  NOR2_X1 U16404 ( .A1(n14684), .A2(n14679), .ZN(P1_U3319) );
  INV_X1 U16405 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14680) );
  NOR2_X1 U16406 ( .A1(n14684), .A2(n14680), .ZN(P1_U3320) );
  INV_X1 U16407 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14681) );
  NOR2_X1 U16408 ( .A1(n14684), .A2(n14681), .ZN(P1_U3321) );
  INV_X1 U16409 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14682) );
  NOR2_X1 U16410 ( .A1(n14684), .A2(n14682), .ZN(P1_U3322) );
  NOR2_X1 U16411 ( .A1(n14684), .A2(n14683), .ZN(P1_U3323) );
  INV_X1 U16412 ( .A(n14729), .ZN(n14721) );
  AOI21_X1 U16413 ( .B1(n9212), .B2(n14723), .A(n14685), .ZN(n14686) );
  OAI21_X1 U16414 ( .B1(n14715), .B2(n14687), .A(n14686), .ZN(n14689) );
  AOI211_X1 U16415 ( .C1(n14721), .C2(n14690), .A(n14689), .B(n14688), .ZN(
        n14752) );
  INV_X1 U16416 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14691) );
  AOI22_X1 U16417 ( .A1(n14751), .A2(n14752), .B1(n14691), .B2(n14749), .ZN(
        P1_U3462) );
  OAI22_X1 U16418 ( .A1(n14693), .A2(n14715), .B1(n14692), .B2(n14743), .ZN(
        n14695) );
  AOI211_X1 U16419 ( .C1(n14748), .C2(n14696), .A(n14695), .B(n14694), .ZN(
        n14753) );
  INV_X1 U16420 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14697) );
  AOI22_X1 U16421 ( .A1(n14751), .A2(n14753), .B1(n14697), .B2(n14749), .ZN(
        P1_U3465) );
  AOI211_X1 U16422 ( .C1(n14700), .C2(n14723), .A(n14699), .B(n14698), .ZN(
        n14701) );
  OAI21_X1 U16423 ( .B1(n14703), .B2(n14702), .A(n14701), .ZN(n14704) );
  INV_X1 U16424 ( .A(n14704), .ZN(n14754) );
  INV_X1 U16425 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14705) );
  AOI22_X1 U16426 ( .A1(n14751), .A2(n14754), .B1(n14705), .B2(n14749), .ZN(
        P1_U3471) );
  INV_X1 U16427 ( .A(n14710), .ZN(n14712) );
  AOI211_X1 U16428 ( .C1(n14708), .C2(n14723), .A(n14707), .B(n14706), .ZN(
        n14709) );
  OAI21_X1 U16429 ( .B1(n14710), .B2(n14729), .A(n14709), .ZN(n14711) );
  AOI21_X1 U16430 ( .B1(n14733), .B2(n14712), .A(n14711), .ZN(n14755) );
  INV_X1 U16431 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14713) );
  AOI22_X1 U16432 ( .A1(n14751), .A2(n14755), .B1(n14713), .B2(n14749), .ZN(
        P1_U3474) );
  OAI21_X1 U16433 ( .B1(n14716), .B2(n14715), .A(n14714), .ZN(n14719) );
  INV_X1 U16434 ( .A(n14717), .ZN(n14718) );
  AOI211_X1 U16435 ( .C1(n14721), .C2(n14720), .A(n14719), .B(n14718), .ZN(
        n14756) );
  INV_X1 U16436 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14722) );
  AOI22_X1 U16437 ( .A1(n14751), .A2(n14756), .B1(n14722), .B2(n14749), .ZN(
        P1_U3477) );
  INV_X1 U16438 ( .A(n14730), .ZN(n14732) );
  AOI22_X1 U16439 ( .A1(n14726), .A2(n14725), .B1(n14724), .B2(n14723), .ZN(
        n14727) );
  OAI211_X1 U16440 ( .C1(n14730), .C2(n14729), .A(n14728), .B(n14727), .ZN(
        n14731) );
  AOI21_X1 U16441 ( .B1(n14733), .B2(n14732), .A(n14731), .ZN(n14757) );
  INV_X1 U16442 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U16443 ( .A1(n14751), .A2(n14757), .B1(n14734), .B2(n14749), .ZN(
        P1_U3480) );
  OAI211_X1 U16444 ( .C1(n14737), .C2(n14743), .A(n14736), .B(n14735), .ZN(
        n14738) );
  AOI21_X1 U16445 ( .B1(n14748), .B2(n14739), .A(n14738), .ZN(n14758) );
  INV_X1 U16446 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14740) );
  AOI22_X1 U16447 ( .A1(n14751), .A2(n14758), .B1(n14740), .B2(n14749), .ZN(
        P1_U3483) );
  INV_X1 U16448 ( .A(n14741), .ZN(n14744) );
  OAI21_X1 U16449 ( .B1(n14744), .B2(n14743), .A(n14742), .ZN(n14746) );
  AOI211_X1 U16450 ( .C1(n14748), .C2(n14747), .A(n14746), .B(n14745), .ZN(
        n14760) );
  INV_X1 U16451 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14750) );
  AOI22_X1 U16452 ( .A1(n14751), .A2(n14760), .B1(n14750), .B2(n14749), .ZN(
        P1_U3489) );
  AOI22_X1 U16453 ( .A1(n14761), .A2(n14752), .B1(n9929), .B2(n14759), .ZN(
        P1_U3529) );
  AOI22_X1 U16454 ( .A1(n14761), .A2(n14753), .B1(n9934), .B2(n14759), .ZN(
        P1_U3530) );
  AOI22_X1 U16455 ( .A1(n14761), .A2(n14754), .B1(n9928), .B2(n14759), .ZN(
        P1_U3532) );
  AOI22_X1 U16456 ( .A1(n14761), .A2(n14755), .B1(n9255), .B2(n14759), .ZN(
        P1_U3533) );
  AOI22_X1 U16457 ( .A1(n14761), .A2(n14756), .B1(n9941), .B2(n14759), .ZN(
        P1_U3534) );
  AOI22_X1 U16458 ( .A1(n14761), .A2(n14757), .B1(n9942), .B2(n14759), .ZN(
        P1_U3535) );
  AOI22_X1 U16459 ( .A1(n14761), .A2(n14758), .B1(n9927), .B2(n14759), .ZN(
        P1_U3536) );
  AOI22_X1 U16460 ( .A1(n14761), .A2(n14760), .B1(n9330), .B2(n14759), .ZN(
        P1_U3538) );
  NOR2_X1 U16461 ( .A1(n14762), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16462 ( .A1(n14762), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14774) );
  OAI21_X1 U16463 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(n14767) );
  OAI22_X1 U16464 ( .A1(n14844), .A2(n14767), .B1(n14766), .B2(n14794), .ZN(
        n14768) );
  INV_X1 U16465 ( .A(n14768), .ZN(n14773) );
  OAI211_X1 U16466 ( .C1(n14771), .C2(n14770), .A(n14838), .B(n14769), .ZN(
        n14772) );
  NAND3_X1 U16467 ( .A1(n14774), .A2(n14773), .A3(n14772), .ZN(P2_U3216) );
  INV_X1 U16468 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15327) );
  INV_X1 U16469 ( .A(n14775), .ZN(n14782) );
  OAI211_X1 U16470 ( .C1(n14778), .C2(n14777), .A(n14816), .B(n14776), .ZN(
        n14779) );
  INV_X1 U16471 ( .A(n14779), .ZN(n14780) );
  AOI211_X1 U16472 ( .C1(n14840), .C2(n14782), .A(n14781), .B(n14780), .ZN(
        n14787) );
  OAI211_X1 U16473 ( .C1(n14785), .C2(n14784), .A(n14838), .B(n14783), .ZN(
        n14786) );
  OAI211_X1 U16474 ( .C1(n14848), .C2(n15327), .A(n14787), .B(n14786), .ZN(
        P2_U3217) );
  OAI211_X1 U16475 ( .C1(n14790), .C2(n14789), .A(n14816), .B(n14788), .ZN(
        n14792) );
  OAI211_X1 U16476 ( .C1(n14794), .C2(n14793), .A(n14792), .B(n14791), .ZN(
        n14795) );
  INV_X1 U16477 ( .A(n14795), .ZN(n14800) );
  OAI211_X1 U16478 ( .C1(n14798), .C2(n14797), .A(n14838), .B(n14796), .ZN(
        n14799) );
  OAI211_X1 U16479 ( .C1(n14848), .C2(n14801), .A(n14800), .B(n14799), .ZN(
        P2_U3218) );
  OAI211_X1 U16480 ( .C1(n14804), .C2(n14803), .A(n14816), .B(n14802), .ZN(
        n14805) );
  INV_X1 U16481 ( .A(n14805), .ZN(n14806) );
  AOI211_X1 U16482 ( .C1(n14840), .C2(n14808), .A(n14807), .B(n14806), .ZN(
        n14813) );
  OAI211_X1 U16483 ( .C1(n14811), .C2(n14810), .A(n14838), .B(n14809), .ZN(
        n14812) );
  OAI211_X1 U16484 ( .C1(n14848), .C2(n15318), .A(n14813), .B(n14812), .ZN(
        P2_U3219) );
  INV_X1 U16485 ( .A(n14814), .ZN(n14821) );
  OAI211_X1 U16486 ( .C1(n14818), .C2(n14817), .A(n14816), .B(n14815), .ZN(
        n14819) );
  INV_X1 U16487 ( .A(n14819), .ZN(n14820) );
  AOI211_X1 U16488 ( .C1(n14840), .C2(n14822), .A(n14821), .B(n14820), .ZN(
        n14827) );
  OAI211_X1 U16489 ( .C1(n14825), .C2(n14824), .A(n14838), .B(n14823), .ZN(
        n14826) );
  OAI211_X1 U16490 ( .C1(n14848), .C2(n14828), .A(n14827), .B(n14826), .ZN(
        P2_U3222) );
  NAND2_X1 U16491 ( .A1(n14830), .A2(n14829), .ZN(n14831) );
  AND2_X1 U16492 ( .A1(n14832), .A2(n14831), .ZN(n14843) );
  NAND2_X1 U16493 ( .A1(n14834), .A2(n14833), .ZN(n14835) );
  NAND2_X1 U16494 ( .A1(n14836), .A2(n14835), .ZN(n14837) );
  NAND2_X1 U16495 ( .A1(n14838), .A2(n14837), .ZN(n14842) );
  NAND2_X1 U16496 ( .A1(n14840), .A2(n14839), .ZN(n14841) );
  OAI211_X1 U16497 ( .C1(n14844), .C2(n14843), .A(n14842), .B(n14841), .ZN(
        n14845) );
  INV_X1 U16498 ( .A(n14845), .ZN(n14847) );
  OAI211_X1 U16499 ( .C1(n14849), .C2(n14848), .A(n14847), .B(n14846), .ZN(
        P2_U3223) );
  NAND2_X1 U16500 ( .A1(n14851), .A2(n14850), .ZN(n14855) );
  INV_X1 U16501 ( .A(n14852), .ZN(n14853) );
  AOI22_X1 U16502 ( .A1(n14890), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14853), 
        .B2(n14865), .ZN(n14854) );
  OAI211_X1 U16503 ( .C1(n14856), .C2(n14874), .A(n14855), .B(n14854), .ZN(
        n14857) );
  AOI21_X1 U16504 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14860) );
  OAI21_X1 U16505 ( .B1(n14890), .B2(n14861), .A(n14860), .ZN(P2_U3258) );
  XNOR2_X1 U16506 ( .A(n14862), .B(n10296), .ZN(n14864) );
  AOI21_X1 U16507 ( .B1(n14864), .B2(n14882), .A(n14863), .ZN(n14907) );
  AOI22_X1 U16508 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(n14890), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n14865), .ZN(n14877) );
  OAI211_X1 U16509 ( .C1(n14906), .C2(n14867), .A(n13215), .B(n14866), .ZN(
        n14905) );
  OR2_X1 U16510 ( .A1(n14868), .A2(n14905), .ZN(n14873) );
  INV_X1 U16511 ( .A(n14869), .ZN(n14870) );
  XNOR2_X1 U16512 ( .A(n10296), .B(n14870), .ZN(n14904) );
  OR2_X1 U16513 ( .A1(n14871), .A2(n14904), .ZN(n14872) );
  OAI211_X1 U16514 ( .C1(n14874), .C2(n14906), .A(n14873), .B(n14872), .ZN(
        n14875) );
  INV_X1 U16515 ( .A(n14875), .ZN(n14876) );
  OAI211_X1 U16516 ( .C1(n14890), .C2(n14907), .A(n14877), .B(n14876), .ZN(
        P2_U3264) );
  NAND2_X1 U16517 ( .A1(n14879), .A2(n14878), .ZN(n14899) );
  OAI22_X1 U16518 ( .A1(n14881), .A2(n8495), .B1(n14880), .B2(n14899), .ZN(
        n14887) );
  OAI21_X1 U16519 ( .B1(n14883), .B2(n14882), .A(n14902), .ZN(n14884) );
  OAI21_X1 U16520 ( .B1(n14886), .B2(n14885), .A(n14884), .ZN(n14900) );
  AOI211_X1 U16521 ( .C1(n14888), .C2(n14902), .A(n14887), .B(n14900), .ZN(
        n14889) );
  AOI22_X1 U16522 ( .A1(n14890), .A2(n10199), .B1(n14889), .B2(n13402), .ZN(
        P2_U3265) );
  INV_X1 U16523 ( .A(n14895), .ZN(n14897) );
  AND2_X1 U16524 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14893), .ZN(P2_U3266) );
  AND2_X1 U16525 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14893), .ZN(P2_U3267) );
  AND2_X1 U16526 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14893), .ZN(P2_U3268) );
  AND2_X1 U16527 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14893), .ZN(P2_U3269) );
  AND2_X1 U16528 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14893), .ZN(P2_U3270) );
  NOR2_X1 U16529 ( .A1(n14892), .A2(n15210), .ZN(P2_U3271) );
  AND2_X1 U16530 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14893), .ZN(P2_U3272) );
  AND2_X1 U16531 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14893), .ZN(P2_U3273) );
  AND2_X1 U16532 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14893), .ZN(P2_U3274) );
  AND2_X1 U16533 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14893), .ZN(P2_U3275) );
  NOR2_X1 U16534 ( .A1(n14892), .A2(n15246), .ZN(P2_U3276) );
  AND2_X1 U16535 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14893), .ZN(P2_U3277) );
  AND2_X1 U16536 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14893), .ZN(P2_U3278) );
  INV_X1 U16537 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15266) );
  NOR2_X1 U16538 ( .A1(n14892), .A2(n15266), .ZN(P2_U3279) );
  NOR2_X1 U16539 ( .A1(n14892), .A2(n15183), .ZN(P2_U3280) );
  AND2_X1 U16540 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14893), .ZN(P2_U3281) );
  AND2_X1 U16541 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14893), .ZN(P2_U3282) );
  NOR2_X1 U16542 ( .A1(n14892), .A2(n15268), .ZN(P2_U3283) );
  AND2_X1 U16543 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14893), .ZN(P2_U3284) );
  AND2_X1 U16544 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14893), .ZN(P2_U3285) );
  AND2_X1 U16545 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14893), .ZN(P2_U3286) );
  AND2_X1 U16546 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14893), .ZN(P2_U3287) );
  AND2_X1 U16547 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14893), .ZN(P2_U3288) );
  AND2_X1 U16548 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14893), .ZN(P2_U3289) );
  AND2_X1 U16549 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14893), .ZN(P2_U3290) );
  AND2_X1 U16550 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14893), .ZN(P2_U3291) );
  AND2_X1 U16551 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14893), .ZN(P2_U3292) );
  AND2_X1 U16552 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14893), .ZN(P2_U3293) );
  AND2_X1 U16553 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14893), .ZN(P2_U3294) );
  AND2_X1 U16554 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14893), .ZN(P2_U3295) );
  AOI22_X1 U16555 ( .A1(n14895), .A2(n14894), .B1(n15212), .B2(n14897), .ZN(
        P2_U3416) );
  AOI21_X1 U16556 ( .B1(n14898), .B2(n14897), .A(n14896), .ZN(P2_U3417) );
  INV_X1 U16557 ( .A(n14899), .ZN(n14901) );
  AOI211_X1 U16558 ( .C1(n14957), .C2(n14902), .A(n14901), .B(n14900), .ZN(
        n14961) );
  INV_X1 U16559 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14903) );
  AOI22_X1 U16560 ( .A1(n14959), .A2(n14961), .B1(n14903), .B2(n14958), .ZN(
        P2_U3430) );
  INV_X1 U16561 ( .A(n14904), .ZN(n14910) );
  OAI21_X1 U16562 ( .B1(n14906), .B2(n14953), .A(n14905), .ZN(n14909) );
  INV_X1 U16563 ( .A(n14907), .ZN(n14908) );
  AOI211_X1 U16564 ( .C1(n14910), .C2(n14918), .A(n14909), .B(n14908), .ZN(
        n14962) );
  INV_X1 U16565 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15192) );
  AOI22_X1 U16566 ( .A1(n14959), .A2(n14962), .B1(n15192), .B2(n14958), .ZN(
        P2_U3433) );
  AOI22_X1 U16567 ( .A1(n14959), .A2(n14911), .B1(n8508), .B2(n14958), .ZN(
        P2_U3436) );
  INV_X1 U16568 ( .A(n14912), .ZN(n14919) );
  OAI21_X1 U16569 ( .B1(n14914), .B2(n14953), .A(n14913), .ZN(n14917) );
  INV_X1 U16570 ( .A(n14915), .ZN(n14916) );
  AOI211_X1 U16571 ( .C1(n14919), .C2(n14918), .A(n14917), .B(n14916), .ZN(
        n14963) );
  INV_X1 U16572 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14920) );
  AOI22_X1 U16573 ( .A1(n14959), .A2(n14963), .B1(n14920), .B2(n14958), .ZN(
        P2_U3439) );
  AOI21_X1 U16574 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14929) );
  INV_X1 U16575 ( .A(n14924), .ZN(n14925) );
  OAI211_X1 U16576 ( .C1(n14927), .C2(n14953), .A(n14926), .B(n14925), .ZN(
        n14928) );
  NOR2_X1 U16577 ( .A1(n14929), .A2(n14928), .ZN(n14965) );
  AOI22_X1 U16578 ( .A1(n14959), .A2(n14965), .B1(n8553), .B2(n14958), .ZN(
        P2_U3442) );
  AND2_X1 U16579 ( .A1(n14931), .A2(n14930), .ZN(n14932) );
  NOR2_X1 U16580 ( .A1(n14933), .A2(n14932), .ZN(n14937) );
  OR2_X1 U16581 ( .A1(n14935), .A2(n14934), .ZN(n14936) );
  AND3_X1 U16582 ( .A1(n14938), .A2(n14937), .A3(n14936), .ZN(n14966) );
  INV_X1 U16583 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14939) );
  AOI22_X1 U16584 ( .A1(n14959), .A2(n14966), .B1(n14939), .B2(n14958), .ZN(
        P2_U3445) );
  OAI21_X1 U16585 ( .B1(n14941), .B2(n14953), .A(n14940), .ZN(n14943) );
  AOI211_X1 U16586 ( .C1(n14957), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        n14968) );
  INV_X1 U16587 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14945) );
  AOI22_X1 U16588 ( .A1(n14959), .A2(n14968), .B1(n14945), .B2(n14958), .ZN(
        P2_U3448) );
  INV_X1 U16589 ( .A(n14946), .ZN(n14951) );
  OAI21_X1 U16590 ( .B1(n14948), .B2(n14953), .A(n14947), .ZN(n14950) );
  AOI211_X1 U16591 ( .C1(n14957), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14970) );
  AOI22_X1 U16592 ( .A1(n14959), .A2(n14970), .B1(n8639), .B2(n14958), .ZN(
        P2_U3454) );
  OAI21_X1 U16593 ( .B1(n7141), .B2(n14953), .A(n14952), .ZN(n14955) );
  AOI211_X1 U16594 ( .C1(n14957), .C2(n14956), .A(n14955), .B(n14954), .ZN(
        n14973) );
  AOI22_X1 U16595 ( .A1(n14959), .A2(n14973), .B1(n8682), .B2(n14958), .ZN(
        P2_U3460) );
  AOI22_X1 U16596 ( .A1(n14974), .A2(n14961), .B1(n14960), .B2(n14971), .ZN(
        P2_U3499) );
  AOI22_X1 U16597 ( .A1(n14974), .A2(n14962), .B1(n8478), .B2(n14971), .ZN(
        P2_U3500) );
  AOI22_X1 U16598 ( .A1(n14974), .A2(n14963), .B1(n10084), .B2(n14971), .ZN(
        P2_U3502) );
  INV_X1 U16599 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n14964) );
  AOI22_X1 U16600 ( .A1(n14974), .A2(n14965), .B1(n14964), .B2(n14971), .ZN(
        P2_U3503) );
  AOI22_X1 U16601 ( .A1(n14974), .A2(n14966), .B1(n10087), .B2(n14971), .ZN(
        P2_U3504) );
  AOI22_X1 U16602 ( .A1(n14974), .A2(n14968), .B1(n14967), .B2(n14971), .ZN(
        P2_U3505) );
  AOI22_X1 U16603 ( .A1(n14974), .A2(n14970), .B1(n14969), .B2(n14971), .ZN(
        P2_U3507) );
  INV_X1 U16604 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U16605 ( .A1(n14974), .A2(n14973), .B1(n14972), .B2(n14971), .ZN(
        P2_U3509) );
  NOR2_X1 U16606 ( .A1(P3_U3897), .A2(n14995), .ZN(P3_U3150) );
  AOI22_X1 U16607 ( .A1(n15017), .A2(P3_IR_REG_0__SCAN_IN), .B1(n14995), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n14981) );
  NOR2_X1 U16608 ( .A1(n14975), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14978) );
  NAND3_X1 U16609 ( .A1(n15001), .A2(n14976), .A3(n14991), .ZN(n14977) );
  OAI21_X1 U16610 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n14980) );
  OAI211_X1 U16611 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n7694), .A(n14981), .B(
        n14980), .ZN(P3_U3182) );
  AOI21_X1 U16612 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n15002) );
  INV_X1 U16613 ( .A(n15013), .ZN(n14988) );
  AOI21_X1 U16614 ( .B1(n14986), .B2(n15012), .A(n14985), .ZN(n14987) );
  AOI21_X1 U16615 ( .B1(n14988), .B2(n15012), .A(n14987), .ZN(n14992) );
  OAI22_X1 U16616 ( .A1(n14992), .A2(n14991), .B1(n14990), .B2(n14989), .ZN(
        n14993) );
  AOI211_X1 U16617 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14995), .A(n14994), .B(
        n14993), .ZN(n15000) );
  OAI21_X1 U16618 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14997), .A(n14996), .ZN(
        n14998) );
  NAND2_X1 U16619 ( .A1(n14998), .A2(n15007), .ZN(n14999) );
  OAI211_X1 U16620 ( .C1(n15002), .C2(n15001), .A(n15000), .B(n14999), .ZN(
        P3_U3191) );
  OAI21_X1 U16621 ( .B1(n15005), .B2(n15004), .A(n15003), .ZN(n15008) );
  AOI21_X1 U16622 ( .B1(n15008), .B2(n15007), .A(n15006), .ZN(n15022) );
  OAI21_X1 U16623 ( .B1(n6857), .B2(n6856), .A(n15010), .ZN(n15020) );
  NAND3_X1 U16624 ( .A1(n15013), .A2(n15012), .A3(n15011), .ZN(n15014) );
  NAND2_X1 U16625 ( .A1(n6582), .A2(n15014), .ZN(n15016) );
  AOI222_X1 U16626 ( .A1(n15020), .A2(n15019), .B1(n15018), .B2(n15017), .C1(
        n15016), .C2(n15015), .ZN(n15021) );
  OAI211_X1 U16627 ( .C1(n15024), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        P3_U3192) );
  OAI21_X1 U16628 ( .B1(n15026), .B2(n15028), .A(n15025), .ZN(n15110) );
  AOI21_X1 U16629 ( .B1(n15028), .B2(n11305), .A(n15027), .ZN(n15034) );
  AOI22_X1 U16630 ( .A1(n15069), .A2(n15030), .B1(n15029), .B2(n15066), .ZN(
        n15033) );
  NAND2_X1 U16631 ( .A1(n15110), .A2(n15031), .ZN(n15032) );
  OAI211_X1 U16632 ( .C1(n15034), .C2(n15043), .A(n15033), .B(n15032), .ZN(
        n15108) );
  AOI21_X1 U16633 ( .B1(n15090), .B2(n15110), .A(n15108), .ZN(n15038) );
  NOR2_X1 U16634 ( .A1(n15035), .A2(n15111), .ZN(n15109) );
  AOI22_X1 U16635 ( .A1(n15058), .A2(n15109), .B1(n15053), .B2(n15036), .ZN(
        n15037) );
  OAI221_X1 U16636 ( .B1(n15093), .B2(n15038), .C1(n15091), .C2(n7745), .A(
        n15037), .ZN(P3_U3228) );
  INV_X1 U16637 ( .A(n15039), .ZN(n15045) );
  AOI21_X1 U16638 ( .B1(n15040), .B2(n15042), .A(n15041), .ZN(n15044) );
  NOR3_X1 U16639 ( .A1(n15045), .A2(n15044), .A3(n15043), .ZN(n15051) );
  OAI22_X1 U16640 ( .A1(n15049), .A2(n15048), .B1(n15047), .B2(n15046), .ZN(
        n15050) );
  NOR2_X1 U16641 ( .A1(n15051), .A2(n15050), .ZN(n15098) );
  AOI22_X1 U16642 ( .A1(n15053), .A2(n15052), .B1(P3_REG2_REG_3__SCAN_IN), 
        .B2(n15093), .ZN(n15061) );
  OAI21_X1 U16643 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(n15101) );
  NOR2_X1 U16644 ( .A1(n15057), .A2(n15111), .ZN(n15100) );
  AOI22_X1 U16645 ( .A1(n15101), .A2(n15059), .B1(n15058), .B2(n15100), .ZN(
        n15060) );
  OAI211_X1 U16646 ( .C1(n15093), .C2(n15098), .A(n15061), .B(n15060), .ZN(
        P3_U3230) );
  XNOR2_X1 U16647 ( .A(n15070), .B(n15062), .ZN(n15077) );
  INV_X1 U16648 ( .A(n15077), .ZN(n15097) );
  NOR2_X1 U16649 ( .A1(n15063), .A2(n15111), .ZN(n15096) );
  INV_X1 U16650 ( .A(n15096), .ZN(n15065) );
  OAI22_X1 U16651 ( .A1(n15065), .A2(n15084), .B1(n15064), .B2(n15083), .ZN(
        n15078) );
  AOI22_X1 U16652 ( .A1(n15069), .A2(n15068), .B1(n15067), .B2(n15066), .ZN(
        n15075) );
  OAI21_X1 U16653 ( .B1(n15071), .B2(n15070), .A(n15040), .ZN(n15073) );
  NAND2_X1 U16654 ( .A1(n15073), .A2(n15072), .ZN(n15074) );
  OAI211_X1 U16655 ( .C1(n15077), .C2(n15076), .A(n15075), .B(n15074), .ZN(
        n15095) );
  AOI211_X1 U16656 ( .C1(n15090), .C2(n15097), .A(n15078), .B(n15095), .ZN(
        n15079) );
  AOI22_X1 U16657 ( .A1(n15093), .A2(n15080), .B1(n15079), .B2(n15091), .ZN(
        P3_U3231) );
  INV_X1 U16658 ( .A(n15081), .ZN(n15085) );
  OAI22_X1 U16659 ( .A1(n15085), .A2(n15084), .B1(n15083), .B2(n15082), .ZN(
        n15088) );
  INV_X1 U16660 ( .A(n15086), .ZN(n15087) );
  AOI211_X1 U16661 ( .C1(n15090), .C2(n15089), .A(n15088), .B(n15087), .ZN(
        n15092) );
  AOI22_X1 U16662 ( .A1(n15093), .A2(n7702), .B1(n15092), .B2(n15091), .ZN(
        P3_U3232) );
  AOI22_X1 U16663 ( .A1(n15137), .A2(n7703), .B1(n15094), .B2(n15136), .ZN(
        P3_U3393) );
  AOI211_X1 U16664 ( .C1(n15097), .C2(n15132), .A(n15096), .B(n15095), .ZN(
        n15138) );
  AOI22_X1 U16665 ( .A1(n15137), .A2(n7679), .B1(n15138), .B2(n15136), .ZN(
        P3_U3396) );
  INV_X1 U16666 ( .A(n15098), .ZN(n15099) );
  AOI211_X1 U16667 ( .C1(n15102), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        n15139) );
  AOI22_X1 U16668 ( .A1(n15137), .A2(n7714), .B1(n15139), .B2(n15136), .ZN(
        P3_U3399) );
  INV_X1 U16669 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15107) );
  NOR2_X1 U16670 ( .A1(n15103), .A2(n15111), .ZN(n15105) );
  AOI211_X1 U16671 ( .C1(n15106), .C2(n15132), .A(n15105), .B(n15104), .ZN(
        n15140) );
  AOI22_X1 U16672 ( .A1(n15137), .A2(n15107), .B1(n15140), .B2(n15136), .ZN(
        P3_U3402) );
  AOI211_X1 U16673 ( .C1(n15132), .C2(n15110), .A(n15109), .B(n15108), .ZN(
        n15141) );
  AOI22_X1 U16674 ( .A1(n15137), .A2(n7749), .B1(n15141), .B2(n15136), .ZN(
        P3_U3405) );
  NOR2_X1 U16675 ( .A1(n15112), .A2(n15111), .ZN(n15114) );
  AOI211_X1 U16676 ( .C1(n15115), .C2(n15132), .A(n15114), .B(n15113), .ZN(
        n15142) );
  AOI22_X1 U16677 ( .A1(n15137), .A2(n7765), .B1(n15142), .B2(n15136), .ZN(
        P3_U3408) );
  INV_X1 U16678 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15120) );
  INV_X1 U16679 ( .A(n15116), .ZN(n15117) );
  AOI211_X1 U16680 ( .C1(n15119), .C2(n15132), .A(n15118), .B(n15117), .ZN(
        n15143) );
  AOI22_X1 U16681 ( .A1(n15137), .A2(n15120), .B1(n15143), .B2(n15136), .ZN(
        P3_U3411) );
  INV_X1 U16682 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15125) );
  AOI21_X1 U16683 ( .B1(n15122), .B2(n15132), .A(n15121), .ZN(n15123) );
  AND2_X1 U16684 ( .A1(n15124), .A2(n15123), .ZN(n15144) );
  AOI22_X1 U16685 ( .A1(n15137), .A2(n15125), .B1(n15144), .B2(n15136), .ZN(
        P3_U3414) );
  INV_X1 U16686 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15130) );
  AOI21_X1 U16687 ( .B1(n15127), .B2(n15132), .A(n15126), .ZN(n15128) );
  AND2_X1 U16688 ( .A1(n15129), .A2(n15128), .ZN(n15146) );
  AOI22_X1 U16689 ( .A1(n15137), .A2(n15130), .B1(n15146), .B2(n15136), .ZN(
        P3_U3417) );
  AOI21_X1 U16690 ( .B1(n15133), .B2(n15132), .A(n15131), .ZN(n15134) );
  AND2_X1 U16691 ( .A1(n15135), .A2(n15134), .ZN(n15148) );
  AOI22_X1 U16692 ( .A1(n15137), .A2(n7829), .B1(n15148), .B2(n15136), .ZN(
        P3_U3420) );
  AOI22_X1 U16693 ( .A1(n15149), .A2(n15138), .B1(n10263), .B2(n15147), .ZN(
        P3_U3461) );
  INV_X1 U16694 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15199) );
  AOI22_X1 U16695 ( .A1(n15149), .A2(n15139), .B1(n15199), .B2(n15147), .ZN(
        P3_U3462) );
  AOI22_X1 U16696 ( .A1(n15149), .A2(n15140), .B1(n7728), .B2(n15147), .ZN(
        P3_U3463) );
  INV_X1 U16697 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15281) );
  AOI22_X1 U16698 ( .A1(n15149), .A2(n15141), .B1(n15281), .B2(n15147), .ZN(
        P3_U3464) );
  AOI22_X1 U16699 ( .A1(n15149), .A2(n15142), .B1(n7762), .B2(n15147), .ZN(
        P3_U3465) );
  AOI22_X1 U16700 ( .A1(n15149), .A2(n15143), .B1(n7782), .B2(n15147), .ZN(
        P3_U3466) );
  AOI22_X1 U16701 ( .A1(n15149), .A2(n15144), .B1(n7796), .B2(n15147), .ZN(
        P3_U3467) );
  AOI22_X1 U16702 ( .A1(n15149), .A2(n15146), .B1(n15145), .B2(n15147), .ZN(
        P3_U3468) );
  AOI22_X1 U16703 ( .A1(n15149), .A2(n15148), .B1(n11070), .B2(n15147), .ZN(
        P3_U3469) );
  NOR2_X1 U16704 ( .A1(keyinput31), .A2(keyinput12), .ZN(n15150) );
  NAND3_X1 U16705 ( .A1(keyinput37), .A2(keyinput36), .A3(n15150), .ZN(n15156)
         );
  NAND3_X1 U16706 ( .A1(keyinput0), .A2(keyinput2), .A3(keyinput49), .ZN(
        n15155) );
  NOR3_X1 U16707 ( .A1(keyinput15), .A2(keyinput22), .A3(keyinput6), .ZN(
        n15153) );
  INV_X1 U16708 ( .A(keyinput53), .ZN(n15151) );
  NOR3_X1 U16709 ( .A1(keyinput57), .A2(keyinput32), .A3(n15151), .ZN(n15152)
         );
  NAND4_X1 U16710 ( .A1(keyinput33), .A2(n15153), .A3(keyinput51), .A4(n15152), 
        .ZN(n15154) );
  NOR4_X1 U16711 ( .A1(keyinput19), .A2(n15156), .A3(n15155), .A4(n15154), 
        .ZN(n15297) );
  NAND4_X1 U16712 ( .A1(keyinput39), .A2(keyinput58), .A3(keyinput40), .A4(
        keyinput13), .ZN(n15177) );
  NOR3_X1 U16713 ( .A1(keyinput10), .A2(keyinput17), .A3(keyinput50), .ZN(
        n15161) );
  INV_X1 U16714 ( .A(keyinput5), .ZN(n15157) );
  NOR4_X1 U16715 ( .A1(keyinput60), .A2(keyinput43), .A3(keyinput59), .A4(
        n15157), .ZN(n15160) );
  NAND2_X1 U16716 ( .A1(keyinput24), .A2(keyinput16), .ZN(n15158) );
  NOR3_X1 U16717 ( .A1(keyinput38), .A2(keyinput47), .A3(n15158), .ZN(n15159)
         );
  NAND4_X1 U16718 ( .A1(keyinput30), .A2(n15161), .A3(n15160), .A4(n15159), 
        .ZN(n15176) );
  NAND2_X1 U16719 ( .A1(keyinput1), .A2(keyinput41), .ZN(n15162) );
  NOR3_X1 U16720 ( .A1(keyinput4), .A2(keyinput9), .A3(n15162), .ZN(n15167) );
  NOR3_X1 U16721 ( .A1(keyinput26), .A2(keyinput20), .A3(keyinput62), .ZN(
        n15166) );
  NAND3_X1 U16722 ( .A1(keyinput28), .A2(keyinput48), .A3(keyinput18), .ZN(
        n15164) );
  NAND3_X1 U16723 ( .A1(keyinput27), .A2(keyinput45), .A3(keyinput44), .ZN(
        n15163) );
  NOR4_X1 U16724 ( .A1(keyinput46), .A2(keyinput42), .A3(n15164), .A4(n15163), 
        .ZN(n15165) );
  NAND4_X1 U16725 ( .A1(n15167), .A2(keyinput14), .A3(n15166), .A4(n15165), 
        .ZN(n15175) );
  NAND2_X1 U16726 ( .A1(keyinput55), .A2(keyinput35), .ZN(n15168) );
  NOR3_X1 U16727 ( .A1(keyinput25), .A2(keyinput34), .A3(n15168), .ZN(n15173)
         );
  NOR3_X1 U16728 ( .A1(keyinput3), .A2(keyinput52), .A3(keyinput11), .ZN(
        n15172) );
  NAND3_X1 U16729 ( .A1(keyinput54), .A2(keyinput56), .A3(keyinput7), .ZN(
        n15170) );
  NAND3_X1 U16730 ( .A1(keyinput21), .A2(keyinput29), .A3(keyinput63), .ZN(
        n15169) );
  NOR4_X1 U16731 ( .A1(keyinput23), .A2(keyinput8), .A3(n15170), .A4(n15169), 
        .ZN(n15171) );
  NAND4_X1 U16732 ( .A1(n15173), .A2(keyinput61), .A3(n15172), .A4(n15171), 
        .ZN(n15174) );
  NOR4_X1 U16733 ( .A1(n15177), .A2(n15176), .A3(n15175), .A4(n15174), .ZN(
        n15296) );
  INV_X1 U16734 ( .A(keyinput10), .ZN(n15179) );
  AOI22_X1 U16735 ( .A1(n15180), .A2(keyinput17), .B1(P3_DATAO_REG_23__SCAN_IN), .B2(n15179), .ZN(n15178) );
  OAI221_X1 U16736 ( .B1(n15180), .B2(keyinput17), .C1(n15179), .C2(
        P3_DATAO_REG_23__SCAN_IN), .A(n15178), .ZN(n15190) );
  INV_X1 U16737 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n15182) );
  AOI22_X1 U16738 ( .A1(n15183), .A2(keyinput43), .B1(keyinput59), .B2(n15182), 
        .ZN(n15181) );
  OAI221_X1 U16739 ( .B1(n15183), .B2(keyinput43), .C1(n15182), .C2(keyinput59), .A(n15181), .ZN(n15189) );
  XNOR2_X1 U16740 ( .A(P1_REG1_REG_28__SCAN_IN), .B(keyinput50), .ZN(n15187)
         );
  XNOR2_X1 U16741 ( .A(P3_IR_REG_26__SCAN_IN), .B(keyinput30), .ZN(n15186) );
  XNOR2_X1 U16742 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput5), .ZN(n15185)
         );
  XNOR2_X1 U16743 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput60), .ZN(n15184) );
  NAND4_X1 U16744 ( .A1(n15187), .A2(n15186), .A3(n15185), .A4(n15184), .ZN(
        n15188) );
  NOR3_X1 U16745 ( .A1(n15190), .A2(n15189), .A3(n15188), .ZN(n15238) );
  AOI22_X1 U16746 ( .A1(n15193), .A2(keyinput39), .B1(n15192), .B2(keyinput58), 
        .ZN(n15191) );
  OAI221_X1 U16747 ( .B1(n15193), .B2(keyinput39), .C1(n15192), .C2(keyinput58), .A(n15191), .ZN(n15205) );
  AOI22_X1 U16748 ( .A1(n8088), .A2(keyinput16), .B1(keyinput38), .B2(n15195), 
        .ZN(n15194) );
  OAI221_X1 U16749 ( .B1(n8088), .B2(keyinput16), .C1(n15195), .C2(keyinput38), 
        .A(n15194), .ZN(n15204) );
  AOI22_X1 U16750 ( .A1(n15198), .A2(keyinput40), .B1(n15197), .B2(keyinput13), 
        .ZN(n15196) );
  OAI221_X1 U16751 ( .B1(n15198), .B2(keyinput40), .C1(n15197), .C2(keyinput13), .A(n15196), .ZN(n15203) );
  XOR2_X1 U16752 ( .A(n15199), .B(keyinput24), .Z(n15201) );
  XNOR2_X1 U16753 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput47), .ZN(n15200) );
  NAND2_X1 U16754 ( .A1(n15201), .A2(n15200), .ZN(n15202) );
  NOR4_X1 U16755 ( .A1(n15205), .A2(n15204), .A3(n15203), .A4(n15202), .ZN(
        n15237) );
  AOI22_X1 U16756 ( .A1(n15207), .A2(keyinput41), .B1(n10199), .B2(keyinput4), 
        .ZN(n15206) );
  OAI221_X1 U16757 ( .B1(n15207), .B2(keyinput41), .C1(n10199), .C2(keyinput4), 
        .A(n15206), .ZN(n15219) );
  AOI22_X1 U16758 ( .A1(n15210), .A2(keyinput1), .B1(keyinput9), .B2(n15209), 
        .ZN(n15208) );
  OAI221_X1 U16759 ( .B1(n15210), .B2(keyinput1), .C1(n15209), .C2(keyinput9), 
        .A(n15208), .ZN(n15218) );
  AOI22_X1 U16760 ( .A1(n11070), .A2(keyinput28), .B1(keyinput48), .B2(n15212), 
        .ZN(n15211) );
  OAI221_X1 U16761 ( .B1(n11070), .B2(keyinput28), .C1(n15212), .C2(keyinput48), .A(n15211), .ZN(n15217) );
  AOI22_X1 U16762 ( .A1(n15215), .A2(keyinput46), .B1(keyinput18), .B2(n15214), 
        .ZN(n15213) );
  OAI221_X1 U16763 ( .B1(n15215), .B2(keyinput46), .C1(n15214), .C2(keyinput18), .A(n15213), .ZN(n15216) );
  NOR4_X1 U16764 ( .A1(n15219), .A2(n15218), .A3(n15217), .A4(n15216), .ZN(
        n15236) );
  AOI22_X1 U16765 ( .A1(n15222), .A2(keyinput27), .B1(keyinput42), .B2(n15221), 
        .ZN(n15220) );
  OAI221_X1 U16766 ( .B1(n15222), .B2(keyinput27), .C1(n15221), .C2(keyinput42), .A(n15220), .ZN(n15223) );
  INV_X1 U16767 ( .A(n15223), .ZN(n15234) );
  XNOR2_X1 U16768 ( .A(P2_REG1_REG_15__SCAN_IN), .B(keyinput62), .ZN(n15226)
         );
  XNOR2_X1 U16769 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput20), .ZN(n15225) );
  XNOR2_X1 U16770 ( .A(keyinput26), .B(P3_REG0_REG_7__SCAN_IN), .ZN(n15224) );
  AND3_X1 U16771 ( .A1(n15226), .A2(n15225), .A3(n15224), .ZN(n15233) );
  INV_X1 U16772 ( .A(keyinput44), .ZN(n15227) );
  XNOR2_X1 U16773 ( .A(n15228), .B(n15227), .ZN(n15232) );
  XNOR2_X1 U16774 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput45), .ZN(n15230) );
  XNOR2_X1 U16775 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput14), .ZN(n15229) );
  AND2_X1 U16776 ( .A1(n15230), .A2(n15229), .ZN(n15231) );
  AND4_X1 U16777 ( .A1(n15234), .A2(n15233), .A3(n15232), .A4(n15231), .ZN(
        n15235) );
  NAND4_X1 U16778 ( .A1(n15238), .A2(n15237), .A3(n15236), .A4(n15235), .ZN(
        n15295) );
  AOI22_X1 U16779 ( .A1(n9974), .A2(keyinput29), .B1(n15240), .B2(keyinput63), 
        .ZN(n15239) );
  OAI221_X1 U16780 ( .B1(n9974), .B2(keyinput29), .C1(n15240), .C2(keyinput63), 
        .A(n15239), .ZN(n15252) );
  AOI22_X1 U16781 ( .A1(n15243), .A2(keyinput21), .B1(n15242), .B2(keyinput8), 
        .ZN(n15241) );
  OAI221_X1 U16782 ( .B1(n15243), .B2(keyinput21), .C1(n15242), .C2(keyinput8), 
        .A(n15241), .ZN(n15251) );
  INV_X1 U16783 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15245) );
  AOI22_X1 U16784 ( .A1(n15246), .A2(keyinput52), .B1(keyinput11), .B2(n15245), 
        .ZN(n15244) );
  OAI221_X1 U16785 ( .B1(n15246), .B2(keyinput52), .C1(n15245), .C2(keyinput11), .A(n15244), .ZN(n15250) );
  AOI22_X1 U16786 ( .A1(n15248), .A2(keyinput61), .B1(keyinput3), .B2(n9954), 
        .ZN(n15247) );
  OAI221_X1 U16787 ( .B1(n15248), .B2(keyinput61), .C1(n9954), .C2(keyinput3), 
        .A(n15247), .ZN(n15249) );
  NOR4_X1 U16788 ( .A1(n15252), .A2(n15251), .A3(n15250), .A4(n15249), .ZN(
        n15293) );
  AOI22_X1 U16789 ( .A1(n11444), .A2(keyinput54), .B1(n15254), .B2(keyinput56), 
        .ZN(n15253) );
  OAI221_X1 U16790 ( .B1(n11444), .B2(keyinput54), .C1(n15254), .C2(keyinput56), .A(n15253), .ZN(n15264) );
  AOI22_X1 U16791 ( .A1(n15257), .A2(keyinput35), .B1(n15256), .B2(keyinput55), 
        .ZN(n15255) );
  OAI221_X1 U16792 ( .B1(n15257), .B2(keyinput35), .C1(n15256), .C2(keyinput55), .A(n15255), .ZN(n15263) );
  XOR2_X1 U16793 ( .A(n9102), .B(keyinput23), .Z(n15261) );
  XNOR2_X1 U16794 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput7), .ZN(n15260) );
  XNOR2_X1 U16795 ( .A(P3_B_REG_SCAN_IN), .B(keyinput34), .ZN(n15259) );
  XNOR2_X1 U16796 ( .A(P3_IR_REG_23__SCAN_IN), .B(keyinput25), .ZN(n15258) );
  NAND4_X1 U16797 ( .A1(n15261), .A2(n15260), .A3(n15259), .A4(n15258), .ZN(
        n15262) );
  NOR3_X1 U16798 ( .A1(n15264), .A2(n15263), .A3(n15262), .ZN(n15292) );
  AOI22_X1 U16799 ( .A1(n15266), .A2(keyinput2), .B1(n8118), .B2(keyinput49), 
        .ZN(n15265) );
  OAI221_X1 U16800 ( .B1(n15266), .B2(keyinput2), .C1(n8118), .C2(keyinput49), 
        .A(n15265), .ZN(n15276) );
  AOI22_X1 U16801 ( .A1(n11257), .A2(keyinput57), .B1(keyinput51), .B2(n15268), 
        .ZN(n15267) );
  OAI221_X1 U16802 ( .B1(n11257), .B2(keyinput57), .C1(n15268), .C2(keyinput51), .A(n15267), .ZN(n15275) );
  AOI22_X1 U16803 ( .A1(n10951), .A2(keyinput53), .B1(n15270), .B2(keyinput32), 
        .ZN(n15269) );
  OAI221_X1 U16804 ( .B1(n10951), .B2(keyinput53), .C1(n15270), .C2(keyinput32), .A(n15269), .ZN(n15274) );
  XNOR2_X1 U16805 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput0), .ZN(n15272) );
  XNOR2_X1 U16806 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(keyinput19), .ZN(n15271)
         );
  NAND2_X1 U16807 ( .A1(n15272), .A2(n15271), .ZN(n15273) );
  NOR4_X1 U16808 ( .A1(n15276), .A2(n15275), .A3(n15274), .A4(n15273), .ZN(
        n15291) );
  AOI22_X1 U16809 ( .A1(n12579), .A2(keyinput37), .B1(keyinput31), .B2(n15278), 
        .ZN(n15277) );
  OAI221_X1 U16810 ( .B1(n12579), .B2(keyinput37), .C1(n15278), .C2(keyinput31), .A(n15277), .ZN(n15289) );
  INV_X1 U16811 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n15280) );
  AOI22_X1 U16812 ( .A1(n15281), .A2(keyinput22), .B1(keyinput6), .B2(n15280), 
        .ZN(n15279) );
  OAI221_X1 U16813 ( .B1(n15281), .B2(keyinput22), .C1(n15280), .C2(keyinput6), 
        .A(n15279), .ZN(n15288) );
  AOI22_X1 U16814 ( .A1(n7672), .A2(keyinput15), .B1(keyinput33), .B2(n15283), 
        .ZN(n15282) );
  OAI221_X1 U16815 ( .B1(n7672), .B2(keyinput15), .C1(n15283), .C2(keyinput33), 
        .A(n15282), .ZN(n15287) );
  XNOR2_X1 U16816 ( .A(P2_REG1_REG_29__SCAN_IN), .B(keyinput12), .ZN(n15285)
         );
  XNOR2_X1 U16817 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput36), .ZN(n15284)
         );
  NAND2_X1 U16818 ( .A1(n15285), .A2(n15284), .ZN(n15286) );
  NOR4_X1 U16819 ( .A1(n15289), .A2(n15288), .A3(n15287), .A4(n15286), .ZN(
        n15290) );
  NAND4_X1 U16820 ( .A1(n15293), .A2(n15292), .A3(n15291), .A4(n15290), .ZN(
        n15294) );
  AOI211_X1 U16821 ( .C1(n15297), .C2(n15296), .A(n15295), .B(n15294), .ZN(
        n15313) );
  AOI22_X1 U16822 ( .A1(n15300), .A2(n15299), .B1(P1_U3086), .B2(
        P1_REG3_REG_8__SCAN_IN), .ZN(n15301) );
  OAI21_X1 U16823 ( .B1(n15303), .B2(n15302), .A(n15301), .ZN(n15309) );
  AOI21_X1 U16824 ( .B1(n15305), .B2(n15304), .A(n6559), .ZN(n15307) );
  NOR2_X1 U16825 ( .A1(n15307), .A2(n15306), .ZN(n15308) );
  AOI211_X1 U16826 ( .C1(n15311), .C2(n15310), .A(n15309), .B(n15308), .ZN(
        n15312) );
  XNOR2_X1 U16827 ( .A(n15313), .B(n15312), .ZN(P1_U3221) );
  OAI21_X1 U16828 ( .B1(n15316), .B2(n15315), .A(n15314), .ZN(SUB_1596_U59) );
  OAI21_X1 U16829 ( .B1(n15319), .B2(n15318), .A(n15317), .ZN(SUB_1596_U58) );
  XOR2_X1 U16830 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15320), .Z(SUB_1596_U53) );
  AOI21_X1 U16831 ( .B1(n15323), .B2(n15322), .A(n15321), .ZN(SUB_1596_U56) );
  AOI21_X1 U16832 ( .B1(n15326), .B2(n15325), .A(n15324), .ZN(n15328) );
  XNOR2_X1 U16833 ( .A(n15328), .B(n15327), .ZN(SUB_1596_U60) );
  AOI21_X1 U16834 ( .B1(n15331), .B2(n15330), .A(n15329), .ZN(SUB_1596_U5) );
  NAND2_X1 U7244 ( .A1(n7266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8464) );
  CLKBUF_X3 U7224 ( .A(n7772), .Z(n6441) );
  OR2_X1 U7239 ( .A1(n15067), .A2(n15057), .ZN(n11644) );
  INV_X2 U7246 ( .A(n13215), .ZN(n12864) );
  NAND2_X2 U7269 ( .A1(n8191), .A2(n8192), .ZN(n10176) );
  AND2_X1 U7279 ( .A1(n11472), .A2(n11471), .ZN(n12360) );
  INV_X2 U7400 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U7473 ( .A1(n13255), .A2(n12081), .ZN(n13239) );
  INV_X2 U8552 ( .A(n9733), .ZN(n13215) );
  CLKBUF_X1 U9441 ( .A(n10143), .Z(n14725) );
endmodule

