

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, 
        P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN, 
        P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN, 
        P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN, 
        P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN, 
        P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN, 
        P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN, 
        P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN, 
        P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN, 
        P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN, 
        P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN,
         P3_REG3_REG_7__SCAN_IN, P3_REG3_REG_27__SCAN_IN,
         P3_REG3_REG_14__SCAN_IN, P3_REG3_REG_23__SCAN_IN,
         P3_REG3_REG_10__SCAN_IN, P3_REG3_REG_3__SCAN_IN,
         P3_REG3_REG_19__SCAN_IN, P3_REG3_REG_28__SCAN_IN,
         P3_REG3_REG_8__SCAN_IN, P3_REG3_REG_1__SCAN_IN,
         P3_REG3_REG_21__SCAN_IN, P3_REG3_REG_12__SCAN_IN,
         P3_REG3_REG_25__SCAN_IN, P3_REG3_REG_16__SCAN_IN,
         P3_REG3_REG_5__SCAN_IN, P3_REG3_REG_17__SCAN_IN,
         P3_REG3_REG_24__SCAN_IN, P3_REG3_REG_4__SCAN_IN,
         P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
         P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
         P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
         P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
         P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
         P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
         P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN,
         P3_ADDR_REG_3__SCAN_IN, P3_ADDR_REG_4__SCAN_IN,
         P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
         P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN,
         P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
         P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
         P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
         P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
         P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
         P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
         P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
         P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
         P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
         P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
         P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
         P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
         P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
         P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
         P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
         P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
         P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
         P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
         P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
         P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
         P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
         P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
         P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
         P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN,
         P3_REG0_REG_3__SCAN_IN, P3_REG0_REG_4__SCAN_IN,
         P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
         P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN,
         P3_REG0_REG_9__SCAN_IN, P3_REG0_REG_10__SCAN_IN,
         P3_REG0_REG_11__SCAN_IN, P3_REG0_REG_12__SCAN_IN,
         P3_REG0_REG_13__SCAN_IN, P3_REG0_REG_14__SCAN_IN,
         P3_REG0_REG_15__SCAN_IN, P3_REG0_REG_16__SCAN_IN,
         P3_REG0_REG_17__SCAN_IN, P3_REG0_REG_18__SCAN_IN,
         P3_REG0_REG_19__SCAN_IN, P3_REG0_REG_20__SCAN_IN,
         P3_REG0_REG_21__SCAN_IN, P3_REG0_REG_22__SCAN_IN,
         P3_REG0_REG_23__SCAN_IN, P3_REG0_REG_24__SCAN_IN,
         P3_REG0_REG_25__SCAN_IN, P3_REG0_REG_26__SCAN_IN,
         P3_REG0_REG_27__SCAN_IN, P3_REG0_REG_28__SCAN_IN,
         P3_REG0_REG_29__SCAN_IN, P3_REG0_REG_30__SCAN_IN,
         P3_REG0_REG_31__SCAN_IN, P3_REG1_REG_0__SCAN_IN,
         P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
         P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN,
         P3_REG1_REG_5__SCAN_IN, P3_REG1_REG_6__SCAN_IN,
         P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
         P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
         P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
         P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
         P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
         P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
         P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
         P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
         P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
         P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
         P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
         P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
         P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
         P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN,
         P3_REG2_REG_3__SCAN_IN, P3_REG2_REG_4__SCAN_IN,
         P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
         P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN,
         P3_REG2_REG_9__SCAN_IN, P3_REG2_REG_10__SCAN_IN,
         P3_REG2_REG_11__SCAN_IN, P3_REG2_REG_12__SCAN_IN,
         P3_REG2_REG_13__SCAN_IN, P3_REG2_REG_14__SCAN_IN,
         P3_REG2_REG_15__SCAN_IN, P3_REG2_REG_16__SCAN_IN,
         P3_REG2_REG_17__SCAN_IN, P3_REG2_REG_18__SCAN_IN,
         P3_REG2_REG_19__SCAN_IN, P3_REG2_REG_20__SCAN_IN,
         P3_REG2_REG_21__SCAN_IN, P3_REG2_REG_22__SCAN_IN,
         P3_REG2_REG_23__SCAN_IN, P3_REG2_REG_24__SCAN_IN,
         P3_REG2_REG_25__SCAN_IN, P3_REG2_REG_26__SCAN_IN,
         P3_REG2_REG_27__SCAN_IN, P3_REG2_REG_28__SCAN_IN,
         P3_REG2_REG_29__SCAN_IN, P3_REG2_REG_30__SCAN_IN,
         P3_REG2_REG_31__SCAN_IN, P3_ADDR_REG_19__SCAN_IN,
         P3_ADDR_REG_18__SCAN_IN, P3_ADDR_REG_17__SCAN_IN,
         P3_ADDR_REG_16__SCAN_IN, P3_ADDR_REG_15__SCAN_IN,
         P3_ADDR_REG_14__SCAN_IN, P3_ADDR_REG_13__SCAN_IN,
         P3_ADDR_REG_12__SCAN_IN, P3_ADDR_REG_11__SCAN_IN,
         P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14473, n14474, n14475,
         n14476, n14477, n14478, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15070,
         n15071, n15072, n15073, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013;

  NAND2_X1 U7279 ( .A1(n14286), .A2(n14272), .ZN(n14274) );
  INV_X4 U7280 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  CLKBUF_X1 U7281 ( .A(n8669), .Z(n7186) );
  AOI21_X1 U7282 ( .B1(n7898), .B2(n7900), .A(n7216), .ZN(n7896) );
  NAND2_X1 U7283 ( .A1(n7697), .A2(n7695), .ZN(n7404) );
  AND2_X1 U7284 ( .A1(n11760), .A2(n11920), .ZN(n15933) );
  AND2_X1 U7285 ( .A1(n11572), .A2(n15830), .ZN(n11599) );
  OR2_X1 U7286 ( .A1(n11687), .A2(n14787), .ZN(n11136) );
  NOR2_X1 U7287 ( .A1(n11332), .A2(n14776), .ZN(n11688) );
  OR2_X1 U7288 ( .A1(n11331), .A2(n14769), .ZN(n11332) );
  CLKBUF_X2 U7289 ( .A(n8292), .Z(n13033) );
  NAND2_X1 U7290 ( .A1(n10505), .A2(n12638), .ZN(n8499) );
  NAND2_X1 U7291 ( .A1(n9996), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9998) );
  CLKBUF_X2 U7292 ( .A(n14941), .Z(n7414) );
  CLKBUF_X1 U7293 ( .A(n9003), .Z(n8906) );
  NAND2_X2 U7294 ( .A1(n13978), .A2(n13158), .ZN(n8292) );
  NAND2_X2 U7295 ( .A1(n11277), .A2(n11276), .ZN(n15848) );
  BUF_X2 U7296 ( .A(n7378), .Z(n14944) );
  BUF_X2 U7297 ( .A(n10336), .Z(n14947) );
  AND3_X1 U7298 ( .A1(n10308), .A2(n10309), .A3(n10307), .ZN(n10771) );
  NAND2_X1 U7300 ( .A1(n7202), .A2(n10304), .ZN(n10336) );
  NAND2_X1 U7301 ( .A1(n7201), .A2(n12638), .ZN(n14929) );
  NAND2_X1 U7302 ( .A1(n14756), .A2(n8110), .ZN(n14988) );
  XNOR2_X1 U7303 ( .A(n10111), .B(n10110), .ZN(n14940) );
  NAND2_X1 U7304 ( .A1(n10109), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U7305 ( .A1(n10135), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10137) );
  NAND2_X1 U7306 ( .A1(n15479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10132) );
  NOR2_X1 U7307 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9979) );
  NOR2_X1 U7308 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9978) );
  NAND2_X1 U7309 ( .A1(n7178), .A2(n8114), .ZN(n14848) );
  NAND3_X1 U7310 ( .A1(n7354), .A2(n7317), .A3(n7353), .ZN(n7178) );
  NAND2_X1 U7311 ( .A1(n7179), .A2(n8116), .ZN(n14885) );
  NAND3_X1 U7312 ( .A1(n7356), .A2(n7314), .A3(n7355), .ZN(n7179) );
  NAND2_X1 U7313 ( .A1(n7987), .A2(n12352), .ZN(n7986) );
  NAND3_X1 U7314 ( .A1(n10146), .A2(n9987), .A3(n7233), .ZN(n8102) );
  NAND2_X1 U7315 ( .A1(n7180), .A2(n8119), .ZN(n14799) );
  NAND3_X1 U7316 ( .A1(n7400), .A2(n7274), .A3(n7399), .ZN(n7180) );
  NAND2_X1 U7317 ( .A1(n9036), .A2(n8775), .ZN(n7620) );
  NAND2_X2 U7318 ( .A1(n8773), .A2(n8772), .ZN(n9036) );
  AND2_X2 U7319 ( .A1(n12776), .A2(n10912), .ZN(n14605) );
  AND2_X2 U7320 ( .A1(n14604), .A2(n10919), .ZN(n10995) );
  NAND2_X1 U7321 ( .A1(n10123), .A2(n7199), .ZN(n7201) );
  XNOR2_X2 U7322 ( .A(n10114), .B(n10113), .ZN(n7199) );
  OR2_X2 U7323 ( .A1(n11720), .A2(n15872), .ZN(n11721) );
  NOR2_X2 U7324 ( .A1(n12212), .A2(n14845), .ZN(n7618) );
  NOR2_X2 U7325 ( .A1(n12021), .A2(n15967), .ZN(n12191) );
  OR2_X2 U7326 ( .A1(n15297), .A2(n15414), .ZN(n15282) );
  AOI22_X1 U7327 ( .A1(n14920), .A2(n14919), .B1(n14918), .B2(n14917), .ZN(
        n7181) );
  AOI22_X1 U7328 ( .A1(n14920), .A2(n14919), .B1(n14918), .B2(n14917), .ZN(
        n15031) );
  INV_X1 U7329 ( .A(n12641), .ZN(n7182) );
  INV_X1 U7330 ( .A(n9012), .ZN(n9213) );
  AND4_X1 U7331 ( .A1(n14774), .A2(n14775), .A3(n14773), .A4(n14772), .ZN(
        n7183) );
  INV_X2 U7332 ( .A(n9475), .ZN(n7188) );
  OR2_X1 U7333 ( .A1(n14191), .A2(n7583), .ZN(n14170) );
  INV_X1 U7334 ( .A(n12116), .ZN(n7540) );
  INV_X1 U7335 ( .A(n12641), .ZN(n12596) );
  OR2_X1 U7336 ( .A1(n15663), .A2(n15660), .ZN(n7709) );
  INV_X1 U7337 ( .A(n9749), .ZN(n9812) );
  INV_X1 U7338 ( .A(n8544), .ZN(n13030) );
  INV_X1 U7339 ( .A(n9321), .ZN(n9331) );
  INV_X1 U7340 ( .A(n11081), .ZN(n9019) );
  NOR2_X1 U7341 ( .A1(n7225), .A2(n7819), .ZN(n7818) );
  INV_X2 U7342 ( .A(n11286), .ZN(n14572) );
  XNOR2_X1 U7343 ( .A(n15300), .B(n14705), .ZN(n15295) );
  AND3_X1 U7344 ( .A1(n10810), .A2(n10809), .A3(n10808), .ZN(n15790) );
  OR2_X1 U7345 ( .A1(n15055), .A2(n10528), .ZN(n14759) );
  AOI21_X1 U7346 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n9881), .A(n9880), .ZN(
        n9939) );
  AOI22_X1 U7347 ( .A1(n9939), .A2(n9883), .B1(P1_ADDR_REG_11__SCAN_IN), .B2(
        n9882), .ZN(n9941) );
  NAND2_X2 U7348 ( .A1(n8669), .A2(n8670), .ZN(n10505) );
  INV_X1 U7349 ( .A(n14079), .ZN(n11064) );
  INV_X1 U7350 ( .A(n10844), .ZN(n14054) );
  NOR2_X1 U7351 ( .A1(n9033), .A2(n9032), .ZN(n10377) );
  MUX2_X1 U7352 ( .A(n14584), .B(n10756), .S(n10755), .Z(n10769) );
  AND4_X1 U7353 ( .A1(n10837), .A2(n10836), .A3(n10835), .A4(n10834), .ZN(
        n11564) );
  XNOR2_X1 U7354 ( .A(n8767), .B(n10051), .ZN(n9010) );
  NAND2_X1 U7355 ( .A1(n15627), .A2(n15625), .ZN(n15631) );
  AND2_X1 U7356 ( .A1(n7711), .A2(n7239), .ZN(n15664) );
  MUX2_X1 U7357 ( .A(n13846), .B(n13914), .S(n15997), .Z(n13847) );
  INV_X1 U7358 ( .A(n10595), .ZN(n10673) );
  INV_X1 U7359 ( .A(n11403), .ZN(n10885) );
  XNOR2_X1 U7360 ( .A(n8900), .B(n8899), .ZN(n13152) );
  CLKBUF_X3 U7361 ( .A(n7199), .Z(n7200) );
  OR2_X1 U7362 ( .A1(n14928), .A2(n10320), .ZN(n7184) );
  AND2_X1 U7363 ( .A1(n8127), .A2(n8128), .ZN(n7185) );
  NOR2_X2 U7364 ( .A1(n15172), .A2(n15146), .ZN(n15155) );
  INV_X1 U7365 ( .A(n14765), .ZN(n14767) );
  INV_X1 U7366 ( .A(n10484), .ZN(n10528) );
  NAND2_X2 U7367 ( .A1(n8686), .A2(n8685), .ZN(n12534) );
  OAI21_X2 U7368 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n9918), .A(n15604), .ZN(
        n9919) );
  OAI21_X2 U7369 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(n11864), .A(n8206), .ZN(
        n8207) );
  NAND4_X2 U7370 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), .ZN(n14080)
         );
  NAND2_X2 U7371 ( .A1(n9349), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9352) );
  NOR3_X2 U7372 ( .A1(n13076), .A2(n12875), .A3(n13690), .ZN(n12884) );
  NOR2_X2 U7373 ( .A1(n12096), .A2(n12097), .ZN(n12366) );
  OAI22_X2 U7374 ( .A1(n15577), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12103), 
        .B2(n12095), .ZN(n12096) );
  OAI21_X2 U7375 ( .B1(n14715), .B2(n14714), .A(n14713), .ZN(n14712) );
  AOI21_X2 U7376 ( .B1(n14660), .B2(n14672), .A(n14671), .ZN(n14715) );
  XNOR2_X2 U7377 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8273) );
  XNOR2_X1 U7378 ( .A(n8218), .B(n8217), .ZN(n8669) );
  AND2_X4 U7380 ( .A1(n8173), .A2(n8172), .ZN(n8654) );
  XNOR2_X2 U7381 ( .A(n7784), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8172) );
  XNOR2_X2 U7382 ( .A(n9001), .B(n9000), .ZN(n9362) );
  NOR2_X2 U7383 ( .A1(n9862), .A2(n9863), .ZN(n9864) );
  NAND2_X2 U7384 ( .A1(n8994), .A2(n8048), .ZN(n9450) );
  NAND2_X2 U7385 ( .A1(n7526), .A2(n7525), .ZN(n8790) );
  AOI211_X1 U7386 ( .C1(n14815), .C2(n14751), .A(n11824), .B(n11823), .ZN(
        n11825) );
  XNOR2_X2 U7387 ( .A(n15445), .B(n15038), .ZN(n14968) );
  AOI21_X1 U7388 ( .B1(n15664), .B2(n15663), .A(n15662), .ZN(n15665) );
  AOI21_X2 U7389 ( .B1(n11923), .B2(n7675), .A(n7672), .ZN(n12377) );
  OAI21_X2 U7390 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(n11773), .A(n8205), .ZN(
        n8537) );
  NAND2_X2 U7391 ( .A1(n9148), .A2(n9147), .ZN(n11881) );
  NAND2_X2 U7392 ( .A1(n12624), .A2(n12623), .ZN(n15300) );
  XNOR2_X1 U7393 ( .A(n11474), .B(n11064), .ZN(n10441) );
  OAI21_X2 U7394 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(n11863), .A(n8208), .ZN(
        n8574) );
  AOI21_X2 U7395 ( .B1(n14089), .B2(n14088), .A(n14087), .ZN(n14103) );
  AOI21_X2 U7396 ( .B1(n12367), .B2(P2_REG2_REG_13__SCAN_IN), .A(n12366), .ZN(
        n14089) );
  NAND2_X2 U7397 ( .A1(n12599), .A2(n12598), .ZN(n15333) );
  XNOR2_X2 U7398 ( .A(n9998), .B(n9997), .ZN(n10281) );
  NOR2_X2 U7399 ( .A1(n9923), .A2(n15611), .ZN(n9926) );
  XNOR2_X2 U7400 ( .A(n8220), .B(n8219), .ZN(n8670) );
  NOR2_X2 U7401 ( .A1(n15614), .A2(n9928), .ZN(n15667) );
  NOR2_X2 U7402 ( .A1(n15616), .A2(n15615), .ZN(n15614) );
  NAND2_X1 U7403 ( .A1(n14028), .A2(n14027), .ZN(n14026) );
  AOI21_X1 U7404 ( .B1(n13996), .B2(n13995), .A(n12817), .ZN(n14028) );
  NAND2_X1 U7405 ( .A1(n15656), .A2(n15654), .ZN(n15661) );
  NOR2_X1 U7406 ( .A1(n9949), .A2(n9950), .ZN(n15655) );
  NAND2_X1 U7407 ( .A1(n9229), .A2(n9228), .ZN(n14418) );
  AOI21_X1 U7408 ( .B1(n13580), .B2(n13579), .A(n13578), .ZN(n13600) );
  OR3_X1 U7409 ( .A1(n9486), .A2(n9489), .A3(n8084), .ZN(n8082) );
  NAND2_X1 U7410 ( .A1(n11585), .A2(n11584), .ZN(n15872) );
  AND2_X1 U7411 ( .A1(n7691), .A2(n7693), .ZN(n9931) );
  INV_X2 U7412 ( .A(n9812), .ZN(n9806) );
  INV_X1 U7413 ( .A(n15790), .ZN(n14783) );
  INV_X2 U7414 ( .A(n9464), .ZN(n11189) );
  BUF_X4 U7415 ( .A(n9475), .Z(n9549) );
  INV_X2 U7416 ( .A(n14628), .ZN(n14584) );
  BUF_X1 U7417 ( .A(n9001), .Z(n11213) );
  CLKBUF_X2 U7418 ( .A(n8270), .Z(n8528) );
  INV_X1 U7419 ( .A(n11208), .ZN(n8303) );
  OAI211_X1 U7420 ( .C1(n10054), .C2(n10505), .A(n8287), .B(n8286), .ZN(n12895) );
  BUF_X4 U7421 ( .A(n12704), .Z(n7189) );
  XNOR2_X1 U7422 ( .A(n9010), .B(n9011), .ZN(n10324) );
  CLKBUF_X2 U7423 ( .A(n9042), .Z(n9168) );
  NAND2_X2 U7424 ( .A1(n11868), .A2(n9720), .ZN(n11173) );
  NAND2_X1 U7425 ( .A1(n7200), .A2(n10123), .ZN(n12641) );
  BUF_X1 U7426 ( .A(n9361), .Z(n12145) );
  XNOR2_X1 U7427 ( .A(n9346), .B(P2_IR_REG_19__SCAN_IN), .ZN(n14140) );
  XNOR2_X1 U7428 ( .A(n7574), .B(n8877), .ZN(n12489) );
  INV_X1 U7429 ( .A(n8763), .ZN(n8995) );
  NOR2_X1 U7430 ( .A1(n9013), .A2(n7573), .ZN(n8871) );
  NAND2_X1 U7431 ( .A1(n10043), .A2(n9983), .ZN(n10046) );
  INV_X2 U7432 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8708) );
  INV_X1 U7433 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n9961) );
  OAI21_X1 U7434 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9716) );
  AND2_X1 U7435 ( .A1(n15917), .A2(n13845), .ZN(n7670) );
  OR2_X1 U7436 ( .A1(n9600), .A2(n9599), .ZN(n9609) );
  AND2_X1 U7437 ( .A1(n14169), .A2(n14168), .ZN(n14375) );
  AND2_X1 U7438 ( .A1(n7883), .A2(n7340), .ZN(n13987) );
  AOI21_X1 U7439 ( .B1(n9405), .B2(n14358), .A(n9404), .ZN(n12869) );
  AOI21_X1 U7440 ( .B1(n7408), .B2(n14358), .A(n7405), .ZN(n14388) );
  NAND2_X1 U7441 ( .A1(n7905), .A2(n7903), .ZN(n14379) );
  XNOR2_X1 U7442 ( .A(n7195), .B(n7196), .ZN(n9964) );
  AOI21_X1 U7443 ( .B1(n14734), .B2(n15387), .A(n15189), .ZN(n15179) );
  NAND2_X1 U7444 ( .A1(n7701), .A2(n7703), .ZN(n7195) );
  OR2_X1 U7445 ( .A1(n15661), .A2(n15660), .ZN(n7711) );
  AND2_X1 U7446 ( .A1(n14235), .A2(n7943), .ZN(n14218) );
  NAND2_X1 U7447 ( .A1(n9343), .A2(n9342), .ZN(n12860) );
  NOR2_X1 U7448 ( .A1(n9571), .A2(n9570), .ZN(n7375) );
  AND2_X1 U7449 ( .A1(n15274), .A2(n12727), .ZN(n8149) );
  OAI21_X1 U7450 ( .B1(n8063), .B2(n9560), .A(n8062), .ZN(n9569) );
  OR2_X1 U7451 ( .A1(n8647), .A2(n13663), .ZN(n12879) );
  NAND2_X1 U7452 ( .A1(n12452), .A2(n12451), .ZN(n12737) );
  AOI21_X1 U7453 ( .B1(n7951), .B2(n7950), .A(n7287), .ZN(n7949) );
  NAND2_X1 U7454 ( .A1(n8637), .A2(n8636), .ZN(n8699) );
  NAND2_X1 U7455 ( .A1(n13984), .A2(n10505), .ZN(n13927) );
  NAND2_X1 U7456 ( .A1(n9275), .A2(n9274), .ZN(n14403) );
  OR2_X1 U7457 ( .A1(n14123), .A2(n14122), .ZN(n14141) );
  NOR2_X1 U7458 ( .A1(n9946), .A2(n9947), .ZN(n15646) );
  XNOR2_X1 U7459 ( .A(n9273), .B(n9272), .ZN(n12650) );
  NAND2_X1 U7460 ( .A1(n15638), .A2(n9945), .ZN(n15642) );
  NAND2_X1 U7461 ( .A1(n12010), .A2(n12009), .ZN(n12195) );
  NAND2_X1 U7462 ( .A1(n9382), .A2(n7365), .ZN(n12392) );
  XNOR2_X1 U7463 ( .A(n9268), .B(n9252), .ZN(n12639) );
  NAND2_X1 U7464 ( .A1(n12611), .A2(n12610), .ZN(n15425) );
  INV_X1 U7465 ( .A(n7387), .ZN(n8607) );
  NAND2_X1 U7466 ( .A1(n12593), .A2(n12592), .ZN(n15436) );
  NOR2_X1 U7467 ( .A1(n8211), .A2(n8210), .ZN(n8562) );
  NAND2_X1 U7468 ( .A1(n12177), .A2(n12176), .ZN(n15982) );
  NAND2_X1 U7469 ( .A1(n8946), .A2(n8945), .ZN(n14444) );
  NAND2_X1 U7470 ( .A1(n8937), .A2(n8936), .ZN(n14438) );
  NAND2_X1 U7471 ( .A1(n8965), .A2(n8964), .ZN(n12126) );
  NAND2_X2 U7472 ( .A1(n12008), .A2(n12007), .ZN(n15967) );
  AND2_X1 U7473 ( .A1(n7433), .A2(n7432), .ZN(n9125) );
  AOI21_X1 U7474 ( .B1(n11377), .B2(n9378), .A(n8136), .ZN(n11339) );
  OAI21_X1 U7475 ( .B1(n11010), .B2(n7875), .A(n7874), .ZN(n11778) );
  NAND2_X1 U7476 ( .A1(n11974), .A2(n11973), .ZN(n14828) );
  NAND2_X1 U7477 ( .A1(n7363), .A2(n9156), .ZN(n8807) );
  NAND2_X1 U7478 ( .A1(n7893), .A2(n7251), .ZN(n15838) );
  XNOR2_X1 U7479 ( .A(n9128), .B(n9127), .ZN(n11742) );
  NAND2_X1 U7480 ( .A1(n8038), .A2(n8039), .ZN(n9157) );
  NAND2_X1 U7481 ( .A1(n14311), .A2(n11176), .ZN(n14349) );
  NOR2_X1 U7482 ( .A1(n9902), .A2(n9901), .ZN(n9880) );
  NAND2_X1 U7483 ( .A1(n9099), .A2(n9098), .ZN(n11389) );
  XNOR2_X1 U7484 ( .A(n9931), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15619) );
  XNOR2_X1 U7485 ( .A(n9112), .B(n9111), .ZN(n11587) );
  NAND2_X2 U7486 ( .A1(n10899), .A2(n15804), .ZN(n15810) );
  NAND2_X1 U7487 ( .A1(n11295), .A2(n11294), .ZN(n14796) );
  AOI22_X1 U7488 ( .A1(n12294), .A2(n12293), .B1(n12292), .B2(n12291), .ZN(
        n15705) );
  XNOR2_X1 U7489 ( .A(n9094), .B(n9095), .ZN(n11274) );
  AND2_X2 U7490 ( .A1(n15165), .A2(n15755), .ZN(n15946) );
  OAI22_X1 U7491 ( .A1(n15688), .A2(n15687), .B1(n11544), .B2(n11553), .ZN(
        n12294) );
  OAI21_X1 U7492 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n10392), .A(n9878), .ZN(
        n9904) );
  OAI21_X1 U7493 ( .B1(n7850), .B2(n7556), .A(n7554), .ZN(n8196) );
  NAND2_X1 U7494 ( .A1(n7619), .A2(n8784), .ZN(n9082) );
  INV_X2 U7495 ( .A(n14572), .ZN(n14587) );
  NAND2_X1 U7496 ( .A1(n7620), .A2(n8781), .ZN(n9066) );
  NAND2_X1 U7497 ( .A1(n7746), .A2(n7745), .ZN(n13487) );
  NAND2_X1 U7498 ( .A1(n9034), .A2(n7930), .ZN(n9464) );
  AND2_X1 U7499 ( .A1(n8278), .A2(n8277), .ZN(n7746) );
  NAND4_X2 U7500 ( .A1(n8311), .A2(n8310), .A3(n8309), .A4(n8308), .ZN(n13485)
         );
  AND4_X1 U7501 ( .A1(n8283), .A2(n8282), .A3(n8281), .A4(n8280), .ZN(n12896)
         );
  NAND4_X1 U7502 ( .A1(n8296), .A2(n8295), .A3(n8294), .A4(n8293), .ZN(n13486)
         );
  NAND4_X1 U7503 ( .A1(n9046), .A2(n9045), .A3(n9044), .A4(n9043), .ZN(n14079)
         );
  INV_X2 U7504 ( .A(n9529), .ZN(n9475) );
  NAND3_X2 U7505 ( .A1(n10001), .A2(n10002), .A3(n10294), .ZN(n10468) );
  CLKBUF_X1 U7506 ( .A(n8906), .Z(n9332) );
  AND2_X1 U7507 ( .A1(n11862), .A2(n12145), .ZN(n10163) );
  NAND2_X2 U7508 ( .A1(n13158), .A2(n8173), .ZN(n8544) );
  BUF_X2 U7509 ( .A(n9028), .Z(n9629) );
  NAND2_X1 U7510 ( .A1(n10276), .A2(n10109), .ZN(n14935) );
  NAND2_X1 U7511 ( .A1(n7804), .A2(n7803), .ZN(n12163) );
  INV_X1 U7512 ( .A(n8173), .ZN(n13978) );
  MUX2_X1 U7513 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10275), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n10276) );
  NOR2_X1 U7514 ( .A1(n9866), .A2(n9867), .ZN(n9908) );
  INV_X1 U7515 ( .A(n10281), .ZN(n10001) );
  OR2_X1 U7516 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  XNOR2_X1 U7517 ( .A(n10000), .B(P1_IR_REG_24__SCAN_IN), .ZN(n10294) );
  XNOR2_X1 U7518 ( .A(n8171), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8173) );
  INV_X2 U7519 ( .A(n10977), .ZN(n13087) );
  NAND2_X1 U7520 ( .A1(n10226), .A2(n10316), .ZN(n9643) );
  AND2_X1 U7521 ( .A1(n13152), .A2(n12548), .ZN(n9042) );
  INV_X2 U7522 ( .A(n10226), .ZN(n9212) );
  INV_X1 U7523 ( .A(n14140), .ZN(n9722) );
  INV_X1 U7524 ( .A(n14940), .ZN(n14757) );
  INV_X2 U7525 ( .A(n13973), .ZN(n13157) );
  OAI21_X1 U7526 ( .B1(n9999), .B2(P1_IR_REG_24__SCAN_IN), .A(n7295), .ZN(
        n7803) );
  AOI21_X1 U7527 ( .B1(n7544), .B2(n7547), .A(n7341), .ZN(n7543) );
  NAND2_X1 U7528 ( .A1(n10277), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U7529 ( .A1(n8100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10117) );
  NAND2_X1 U7530 ( .A1(n7608), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10114) );
  OR2_X1 U7531 ( .A1(n14471), .A2(n8875), .ZN(n8900) );
  INV_X4 U7532 ( .A(n12638), .ZN(n10316) );
  OAI21_X1 U7533 ( .B1(n8715), .B2(P3_IR_REG_27__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8218) );
  OR2_X1 U7534 ( .A1(n10106), .A2(n11229), .ZN(n10108) );
  NAND2_X1 U7535 ( .A1(n8876), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7574) );
  CLKBUF_X1 U7536 ( .A(n7782), .Z(n7480) );
  NAND2_X1 U7537 ( .A1(n7592), .A2(n7591), .ZN(n10272) );
  AND2_X1 U7538 ( .A1(n10130), .A2(n7410), .ZN(n10133) );
  AND2_X1 U7539 ( .A1(n8159), .A2(n8141), .ZN(n7782) );
  AND4_X2 U7540 ( .A1(n8871), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n8067)
         );
  AND4_X1 U7541 ( .A1(n8874), .A2(n8873), .A3(n9348), .A4(n8872), .ZN(n8132)
         );
  AND2_X1 U7542 ( .A1(n10112), .A2(n9997), .ZN(n10130) );
  XNOR2_X1 U7543 ( .A(n7714), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n9911) );
  AND2_X1 U7544 ( .A1(n9994), .A2(n9993), .ZN(n10112) );
  AND2_X1 U7545 ( .A1(n8161), .A2(n8160), .ZN(n7483) );
  AND3_X1 U7546 ( .A1(n8868), .A2(n8867), .A3(n8866), .ZN(n8930) );
  AND4_X1 U7547 ( .A1(n9347), .A2(n9187), .A3(n9434), .A4(n9428), .ZN(n8874)
         );
  AND3_X1 U7548 ( .A1(n8974), .A2(n9113), .A3(n9129), .ZN(n8929) );
  AND2_X1 U7549 ( .A1(n8870), .A2(n8869), .ZN(n8931) );
  NOR2_X1 U7550 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n8164) );
  INV_X1 U7551 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8513) );
  INV_X1 U7552 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10092) );
  INV_X4 U7553 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7554 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8165) );
  INV_X1 U7555 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10417) );
  INV_X1 U7556 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9014) );
  INV_X1 U7557 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9915) );
  NOR2_X1 U7558 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n9992) );
  INV_X1 U7559 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n11227) );
  INV_X1 U7560 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n11231) );
  NOR2_X1 U7561 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n9985) );
  INV_X1 U7562 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10107) );
  INV_X1 U7563 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8224) );
  NOR2_X2 U7564 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n10043) );
  INV_X1 U7565 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9428) );
  NOR2_X1 U7566 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8867) );
  NOR2_X1 U7567 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8868) );
  INV_X1 U7568 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9434) );
  INV_X1 U7569 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8933) );
  NOR2_X1 U7570 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n9348) );
  INV_X1 U7571 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8899) );
  INV_X1 U7572 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8974) );
  INV_X1 U7573 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9347) );
  INV_X1 U7574 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9113) );
  INV_X1 U7575 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U7576 ( .A1(n8127), .A2(n7193), .ZN(n7190) );
  AND2_X1 U7577 ( .A1(n7190), .A2(n7191), .ZN(n14906) );
  OR2_X1 U7578 ( .A1(n7192), .A2(n14903), .ZN(n7191) );
  INV_X1 U7579 ( .A(n14902), .ZN(n7192) );
  AND2_X1 U7580 ( .A1(n8128), .A2(n14902), .ZN(n7193) );
  NAND2_X1 U7581 ( .A1(n14853), .A2(n14852), .ZN(n14856) );
  NOR2_X2 U7582 ( .A1(n12057), .A2(n12126), .ZN(n11956) );
  NAND2_X2 U7583 ( .A1(n14209), .A2(n14194), .ZN(n14191) );
  NOR2_X2 U7584 ( .A1(n11382), .A2(n12854), .ZN(n7584) );
  NAND2_X1 U7585 ( .A1(n9366), .A2(n9365), .ZN(n10538) );
  AOI21_X1 U7586 ( .B1(n9390), .B2(n9389), .A(n9388), .ZN(n14237) );
  AOI21_X2 U7587 ( .B1(n12392), .B2(n12396), .A(n7364), .ZN(n12468) );
  NOR2_X2 U7588 ( .A1(n15632), .A2(n15631), .ZN(n15630) );
  AOI21_X2 U7589 ( .B1(P3_ADDR_REG_4__SCAN_IN), .B2(n9869), .A(n9868), .ZN(
        n9924) );
  OAI22_X1 U7590 ( .A1(n9873), .A2(n9929), .B1(P3_ADDR_REG_6__SCAN_IN), .B2(
        n9872), .ZN(n9874) );
  OAI21_X1 U7591 ( .B1(n8367), .B2(n8186), .A(n8187), .ZN(n7194) );
  OAI21_X1 U7592 ( .B1(n8367), .B2(n8186), .A(n8187), .ZN(n8264) );
  XNOR2_X1 U7593 ( .A(n8196), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8437) );
  NAND2_X1 U7594 ( .A1(n13693), .A2(n12887), .ZN(n13076) );
  OR2_X2 U7595 ( .A1(n13085), .A2(n13084), .ZN(n7249) );
  XOR2_X1 U7596 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n7196) );
  NAND2_X1 U7597 ( .A1(n8273), .A2(n8285), .ZN(n8178) );
  NAND2_X1 U7598 ( .A1(n14605), .A2(n14606), .ZN(n14604) );
  NAND2_X2 U7599 ( .A1(n14652), .A2(n14653), .ZN(n14651) );
  NOR2_X2 U7600 ( .A1(n9936), .A2(n9937), .ZN(n15626) );
  OR2_X1 U7601 ( .A1(n7197), .A2(n14769), .ZN(n7413) );
  NOR2_X1 U7602 ( .A1(n14770), .A2(n14814), .ZN(n7197) );
  INV_X1 U7603 ( .A(n11700), .ZN(n7198) );
  NAND2_X1 U7604 ( .A1(n12228), .A2(n7799), .ZN(n12275) );
  AOI21_X1 U7605 ( .B1(n9559), .B2(n9558), .A(n9557), .ZN(n9560) );
  INV_X1 U7606 ( .A(n15053), .ZN(n14607) );
  OR2_X1 U7607 ( .A1(n12705), .A2(n11734), .ZN(n10332) );
  BUF_X4 U7608 ( .A(n12692), .Z(n12705) );
  OR2_X2 U7609 ( .A1(n14755), .A2(n15140), .ZN(n14756) );
  INV_X1 U7610 ( .A(n13159), .ZN(n10298) );
  NAND4_X2 U7611 ( .A1(n10323), .A2(n7184), .A3(n10322), .A4(n10321), .ZN(
        n15053) );
  NOR2_X2 U7612 ( .A1(n13103), .A2(n7389), .ZN(n12816) );
  NOR3_X2 U7613 ( .A1(n13095), .A2(n12811), .A3(n14009), .ZN(n13103) );
  NAND2_X1 U7614 ( .A1(n11073), .A2(n10952), .ZN(n11010) );
  OAI211_X2 U7615 ( .C1(n7518), .C2(n11875), .A(n11803), .B(n7517), .ZN(n11893) );
  INV_X1 U7616 ( .A(n14581), .ZN(n14627) );
  INV_X1 U7617 ( .A(n14563), .ZN(n14626) );
  CLKBUF_X3 U7618 ( .A(n14814), .Z(n14991) );
  NAND2_X2 U7619 ( .A1(n7393), .A2(n8109), .ZN(n14814) );
  NOR2_X2 U7620 ( .A1(n11879), .A2(n11509), .ZN(n11846) );
  INV_X2 U7621 ( .A(n14814), .ZN(n14941) );
  INV_X1 U7622 ( .A(n14814), .ZN(n14992) );
  AND2_X1 U7623 ( .A1(n9361), .A2(n14140), .ZN(n9452) );
  NAND2_X2 U7624 ( .A1(n10298), .A2(n10297), .ZN(n12704) );
  AOI21_X2 U7625 ( .B1(n14693), .B2(n7810), .A(n7808), .ZN(n7807) );
  AOI21_X2 U7626 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(n9938), .A(n15630), .ZN(
        n15636) );
  NAND2_X1 U7627 ( .A1(n7199), .A2(n10123), .ZN(n7202) );
  OR2_X1 U7628 ( .A1(n11700), .A2(n8131), .ZN(n10109) );
  NOR2_X1 U7629 ( .A1(n11700), .A2(n7291), .ZN(n10106) );
  XNOR2_X2 U7630 ( .A(n7575), .B(n8898), .ZN(n9400) );
  NOR2_X2 U7631 ( .A1(n11136), .A2(n15813), .ZN(n11572) );
  AND2_X2 U7632 ( .A1(n15257), .A2(n12667), .ZN(n15246) );
  NOR2_X2 U7633 ( .A1(n15409), .A2(n15282), .ZN(n15257) );
  NOR2_X2 U7634 ( .A1(n15327), .A2(n15425), .ZN(n15311) );
  NAND2_X1 U7635 ( .A1(n13978), .A2(n8172), .ZN(n8270) );
  INV_X2 U7636 ( .A(n13002), .ZN(n13012) );
  OAI21_X1 U7637 ( .B1(n7227), .B2(n7900), .A(n9251), .ZN(n7899) );
  OR2_X1 U7638 ( .A1(n14413), .A2(n14251), .ZN(n9251) );
  INV_X1 U7639 ( .A(n7901), .ZN(n7900) );
  INV_X1 U7640 ( .A(n11841), .ZN(n7919) );
  INV_X1 U7641 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8866) );
  OR2_X1 U7642 ( .A1(n9419), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9433) );
  OR2_X1 U7643 ( .A1(n9158), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9160) );
  INV_X1 U7644 ( .A(n9004), .ZN(n9321) );
  XNOR2_X1 U7645 ( .A(n7628), .B(n15140), .ZN(n14987) );
  AOI21_X1 U7646 ( .B1(n12937), .B2(n12936), .A(n12935), .ZN(n12942) );
  INV_X1 U7647 ( .A(n13076), .ZN(n13004) );
  OR2_X1 U7648 ( .A1(n13873), .A2(n13763), .ZN(n12992) );
  NAND2_X1 U7649 ( .A1(n7639), .A2(n7638), .ZN(n8860) );
  AOI21_X1 U7650 ( .B1(n7640), .B2(n9299), .A(n7347), .ZN(n7638) );
  NAND2_X1 U7651 ( .A1(n8820), .A2(n13405), .ZN(n8823) );
  NAND2_X1 U7652 ( .A1(n7461), .A2(n7458), .ZN(n7460) );
  NOR2_X1 U7653 ( .A1(n9797), .A2(n7459), .ZN(n7458) );
  INV_X1 U7654 ( .A(n9796), .ZN(n7459) );
  NAND2_X1 U7655 ( .A1(n7457), .A2(n7455), .ZN(n9799) );
  AOI21_X1 U7656 ( .B1(n13176), .B2(n9796), .A(n7456), .ZN(n7455) );
  INV_X1 U7657 ( .A(n9785), .ZN(n7492) );
  NOR2_X1 U7658 ( .A1(n13631), .A2(n7752), .ZN(n13630) );
  OR2_X1 U7659 ( .A1(n8699), .A2(n13675), .ZN(n12877) );
  OR2_X1 U7660 ( .A1(n13784), .A2(n13800), .ZN(n12983) );
  INV_X1 U7661 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8710) );
  INV_X1 U7662 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7484) );
  INV_X1 U7663 ( .A(n7555), .ZN(n7554) );
  OAI21_X1 U7664 ( .B1(n7849), .B2(n7556), .A(n8195), .ZN(n7555) );
  INV_X1 U7665 ( .A(n8194), .ZN(n7854) );
  INV_X1 U7666 ( .A(n7853), .ZN(n7852) );
  OAI21_X1 U7667 ( .B1(n8405), .B2(n7854), .A(n8417), .ZN(n7853) );
  OR2_X1 U7668 ( .A1(n14407), .A2(n14396), .ZN(n7579) );
  NAND2_X1 U7669 ( .A1(n14217), .A2(n14220), .ZN(n14216) );
  NAND3_X1 U7670 ( .A1(n8067), .A2(n8066), .A3(n8132), .ZN(n8901) );
  AND2_X1 U7671 ( .A1(n8877), .A2(n8898), .ZN(n8066) );
  INV_X1 U7672 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8898) );
  AND2_X1 U7673 ( .A1(n9354), .A2(n9353), .ZN(n9357) );
  INV_X1 U7674 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9354) );
  INV_X1 U7675 ( .A(n12649), .ZN(n7506) );
  OR2_X1 U7676 ( .A1(n15224), .A2(n8105), .ZN(n8104) );
  INV_X1 U7677 ( .A(n12668), .ZN(n8105) );
  NAND2_X1 U7678 ( .A1(n15254), .A2(n7981), .ZN(n7984) );
  NOR2_X1 U7679 ( .A1(n7982), .A2(n15240), .ZN(n7981) );
  INV_X1 U7680 ( .A(n12729), .ZN(n7982) );
  NOR2_X1 U7681 ( .A1(n8108), .A2(n8107), .ZN(n8106) );
  INV_X1 U7682 ( .A(n15240), .ZN(n8107) );
  INV_X1 U7683 ( .A(n12653), .ZN(n8108) );
  NAND2_X1 U7684 ( .A1(n8149), .A2(n12728), .ZN(n15254) );
  AND2_X1 U7685 ( .A1(n12594), .A2(n12589), .ZN(n8094) );
  INV_X1 U7686 ( .A(n15340), .ZN(n12594) );
  NAND2_X1 U7687 ( .A1(n11580), .A2(n7977), .ZN(n7976) );
  NOR2_X1 U7688 ( .A1(n11654), .A2(n7978), .ZN(n7977) );
  INV_X1 U7689 ( .A(n11579), .ZN(n7978) );
  NAND2_X1 U7690 ( .A1(n7651), .A2(n7649), .ZN(n9287) );
  AOI21_X1 U7691 ( .B1(n7653), .B2(n7655), .A(n7650), .ZN(n7649) );
  INV_X1 U7692 ( .A(n8847), .ZN(n7650) );
  NAND2_X1 U7693 ( .A1(n7411), .A2(n7277), .ZN(n9183) );
  NAND2_X1 U7694 ( .A1(n8807), .A2(n7625), .ZN(n7411) );
  NAND2_X1 U7695 ( .A1(n7625), .A2(n7627), .ZN(n7623) );
  NAND2_X1 U7696 ( .A1(n8032), .A2(n8811), .ZN(n8939) );
  NAND2_X1 U7697 ( .A1(n9112), .A2(n8792), .ZN(n8795) );
  INV_X1 U7698 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U7699 ( .A1(n8004), .A2(n8007), .ZN(n8003) );
  INV_X1 U7700 ( .A(n8005), .ZN(n8004) );
  INV_X1 U7701 ( .A(n9759), .ZN(n7477) );
  INV_X1 U7702 ( .A(n7231), .ZN(n7471) );
  NAND2_X1 U7703 ( .A1(n11239), .A2(n11238), .ZN(n11237) );
  NAND2_X1 U7704 ( .A1(n7559), .A2(n13014), .ZN(n7362) );
  NAND2_X1 U7705 ( .A1(n7742), .A2(n13595), .ZN(n7741) );
  AND2_X1 U7706 ( .A1(n13043), .A2(n13040), .ZN(n13051) );
  NAND2_X1 U7707 ( .A1(n7688), .A2(n8553), .ZN(n13754) );
  NAND2_X1 U7708 ( .A1(n13774), .A2(n8552), .ZN(n7688) );
  NOR2_X1 U7709 ( .A1(n13818), .A2(n12972), .ZN(n7682) );
  AOI21_X1 U7710 ( .B1(n7660), .B2(n7662), .A(n13070), .ZN(n7658) );
  OAI21_X1 U7711 ( .B1(n12254), .B2(n8409), .A(n12943), .ZN(n12382) );
  NAND2_X1 U7712 ( .A1(n11926), .A2(n8682), .ZN(n12044) );
  AOI21_X1 U7713 ( .B1(n13054), .B2(n7769), .A(n7768), .ZN(n7767) );
  INV_X1 U7714 ( .A(n12924), .ZN(n7768) );
  INV_X1 U7715 ( .A(n12919), .ZN(n7769) );
  INV_X1 U7716 ( .A(n13610), .ZN(n8706) );
  NAND2_X1 U7717 ( .A1(n10895), .A2(n10894), .ZN(n10899) );
  NAND2_X1 U7718 ( .A1(n8226), .A2(n8225), .ZN(n13638) );
  INV_X1 U7719 ( .A(n13756), .ZN(n13831) );
  INV_X1 U7720 ( .A(n13026), .ZN(n13021) );
  INV_X1 U7721 ( .A(n8499), .ZN(n13028) );
  OR2_X1 U7722 ( .A1(n13012), .A2(n9841), .ZN(n13833) );
  NAND2_X1 U7723 ( .A1(n13967), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U7724 ( .A1(n8170), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8171) );
  INV_X1 U7725 ( .A(n7496), .ZN(n7493) );
  NAND2_X1 U7726 ( .A1(n8469), .A2(n8470), .ZN(n8201) );
  NAND2_X1 U7727 ( .A1(n8406), .A2(n7852), .ZN(n7850) );
  XNOR2_X1 U7728 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8326) );
  NAND2_X1 U7729 ( .A1(n8061), .A2(n10009), .ZN(n8058) );
  INV_X1 U7730 ( .A(n8904), .ZN(n9633) );
  NOR2_X1 U7731 ( .A1(n13152), .A2(n8905), .ZN(n9005) );
  AND2_X1 U7732 ( .A1(n8903), .A2(n8905), .ZN(n9004) );
  INV_X1 U7733 ( .A(n8067), .ZN(n9211) );
  OAI22_X1 U7734 ( .A1(n14201), .A2(n14205), .B1(n14213), .B2(n14221), .ZN(
        n14189) );
  OAI22_X1 U7735 ( .A1(n14295), .A2(n7428), .B1(n7279), .B2(n7427), .ZN(n14242) );
  INV_X1 U7736 ( .A(n7431), .ZN(n7427) );
  NAND2_X1 U7737 ( .A1(n7896), .A2(n7431), .ZN(n7428) );
  AND2_X1 U7738 ( .A1(n14407), .A2(n14009), .ZN(n9388) );
  NAND2_X1 U7739 ( .A1(n14257), .A2(n14065), .ZN(n9389) );
  NAND2_X1 U7740 ( .A1(n14323), .A2(n9200), .ZN(n14296) );
  OR2_X1 U7741 ( .A1(n14428), .A2(n14356), .ZN(n9200) );
  OAI21_X1 U7742 ( .B1(n14339), .B2(n14351), .A(n7426), .ZN(n14325) );
  OR2_X1 U7743 ( .A1(n14433), .A2(n14068), .ZN(n7426) );
  AND2_X1 U7744 ( .A1(n14318), .A2(n7246), .ZN(n7937) );
  OR2_X1 U7745 ( .A1(n14438), .A2(n12394), .ZN(n9383) );
  NOR2_X1 U7746 ( .A1(n7895), .A2(n9553), .ZN(n7364) );
  NAND2_X1 U7747 ( .A1(n7912), .A2(n7911), .ZN(n11952) );
  NAND2_X1 U7748 ( .A1(n7915), .A2(n7237), .ZN(n7911) );
  NAND2_X1 U7749 ( .A1(n7919), .A2(n9141), .ZN(n7916) );
  NAND2_X1 U7750 ( .A1(n7935), .A2(n7934), .ZN(n11513) );
  AOI21_X1 U7751 ( .B1(n11342), .B2(n7203), .A(n7281), .ZN(n7934) );
  NAND2_X1 U7752 ( .A1(n9372), .A2(n9371), .ZN(n10778) );
  NAND2_X1 U7753 ( .A1(n7376), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U7754 ( .A1(n8067), .A2(n7258), .ZN(n7376) );
  AND2_X1 U7755 ( .A1(n9161), .A2(n9160), .ZN(n12367) );
  XNOR2_X1 U7756 ( .A(n11300), .B(n11299), .ZN(n11416) );
  AND2_X1 U7757 ( .A1(n7820), .A2(n7234), .ZN(n7819) );
  INV_X1 U7758 ( .A(n7823), .ZN(n7821) );
  AND2_X1 U7759 ( .A1(n14624), .A2(n7795), .ZN(n7794) );
  NAND2_X1 U7760 ( .A1(n7796), .A2(n14730), .ZN(n7795) );
  INV_X1 U7761 ( .A(n14728), .ZN(n7796) );
  OAI21_X1 U7762 ( .B1(n15000), .B2(n7644), .A(n7294), .ZN(n8015) );
  OR2_X1 U7763 ( .A1(n15009), .A2(n15013), .ZN(n7644) );
  INV_X1 U7764 ( .A(n14924), .ZN(n12686) );
  INV_X1 U7765 ( .A(n14928), .ZN(n12711) );
  INV_X1 U7766 ( .A(n15176), .ZN(n15196) );
  NAND2_X1 U7767 ( .A1(n12667), .A2(n14599), .ZN(n7983) );
  NAND2_X1 U7768 ( .A1(n7512), .A2(n7511), .ZN(n12607) );
  AND2_X1 U7769 ( .A1(n7513), .A2(n15324), .ZN(n7511) );
  NAND2_X1 U7770 ( .A1(n12720), .A2(n12719), .ZN(n15338) );
  NOR2_X1 U7771 ( .A1(n7263), .A2(n10829), .ZN(n8090) );
  INV_X1 U7772 ( .A(n15195), .ZN(n15342) );
  NAND2_X1 U7773 ( .A1(n10349), .A2(n10348), .ZN(n15988) );
  AND2_X1 U7774 ( .A1(n10468), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10119) );
  NAND2_X1 U7775 ( .A1(n12588), .A2(n12587), .ZN(n15387) );
  NAND2_X1 U7776 ( .A1(n15648), .A2(n15649), .ZN(n15645) );
  MUX2_X1 U7777 ( .A(n14776), .B(n15052), .S(n14941), .Z(n14780) );
  NAND2_X1 U7778 ( .A1(n9450), .A2(n9529), .ZN(n9454) );
  NAND2_X1 U7779 ( .A1(n8070), .A2(n9482), .ZN(n8069) );
  NOR2_X1 U7780 ( .A1(n9471), .A2(n9468), .ZN(n9469) );
  OR2_X1 U7781 ( .A1(n9492), .A2(n9493), .ZN(n8083) );
  NOR2_X1 U7782 ( .A1(n8086), .A2(n8085), .ZN(n8084) );
  INV_X1 U7783 ( .A(n7310), .ZN(n8078) );
  NAND2_X1 U7784 ( .A1(n8064), .A2(n8065), .ZN(n9559) );
  NAND2_X1 U7785 ( .A1(n9554), .A2(n7254), .ZN(n8065) );
  INV_X1 U7786 ( .A(n9577), .ZN(n7374) );
  INV_X1 U7787 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9977) );
  INV_X1 U7788 ( .A(n7529), .ZN(n7528) );
  OAI21_X1 U7789 ( .B1(n8785), .B2(n7530), .A(n8788), .ZN(n7529) );
  INV_X1 U7790 ( .A(n8787), .ZN(n7530) );
  NOR2_X1 U7791 ( .A1(n7754), .A2(n7751), .ZN(n7750) );
  NAND2_X1 U7792 ( .A1(n7752), .A2(n12882), .ZN(n7751) );
  NAND2_X1 U7793 ( .A1(n13487), .A2(n11217), .ZN(n12894) );
  INV_X1 U7794 ( .A(n9133), .ZN(n7539) );
  NOR2_X1 U7795 ( .A1(n15275), .A2(n7508), .ZN(n7507) );
  INV_X1 U7796 ( .A(n12636), .ZN(n7508) );
  INV_X1 U7797 ( .A(n8841), .ZN(n7655) );
  NAND2_X1 U7798 ( .A1(n8816), .A2(n13409), .ZN(n8819) );
  AOI21_X1 U7799 ( .B1(n8033), .B2(n8035), .A(n8031), .ZN(n8030) );
  INV_X1 U7800 ( .A(n8815), .ZN(n8031) );
  INV_X1 U7801 ( .A(n8799), .ZN(n8041) );
  NAND2_X1 U7802 ( .A1(n9758), .A2(n13482), .ZN(n8007) );
  INV_X1 U7803 ( .A(n11932), .ZN(n7474) );
  AND2_X1 U7804 ( .A1(n10622), .A2(n10598), .ZN(n7723) );
  INV_X1 U7805 ( .A(n10598), .ZN(n7720) );
  NOR2_X1 U7806 ( .A1(n10987), .A2(n7335), .ZN(n11545) );
  NOR2_X1 U7807 ( .A1(n15694), .A2(n7732), .ZN(n12280) );
  NOR2_X1 U7808 ( .A1(n15686), .A2(n7733), .ZN(n7732) );
  AOI21_X1 U7809 ( .B1(n12302), .B2(P3_REG1_REG_12__SCAN_IN), .A(n15714), .ZN(
        n12284) );
  AOI21_X1 U7810 ( .B1(n13065), .B2(n8453), .A(n7664), .ZN(n7663) );
  NAND2_X1 U7811 ( .A1(n8409), .A2(n7674), .ZN(n7673) );
  INV_X1 U7812 ( .A(n7676), .ZN(n7674) );
  NAND2_X1 U7813 ( .A1(n7680), .A2(n7678), .ZN(n7677) );
  NAND2_X1 U7814 ( .A1(n12931), .A2(n7681), .ZN(n7678) );
  INV_X1 U7815 ( .A(n13055), .ZN(n8353) );
  OR2_X1 U7816 ( .A1(n13485), .A2(n15782), .ZN(n12893) );
  NAND2_X1 U7817 ( .A1(n11149), .A2(n12897), .ZN(n7684) );
  OR2_X1 U7818 ( .A1(n8488), .A2(n13457), .ZN(n8281) );
  NAND2_X1 U7819 ( .A1(n7776), .A2(n7774), .ZN(n7773) );
  AND2_X1 U7820 ( .A1(n8747), .A2(n13092), .ZN(n13002) );
  INV_X1 U7821 ( .A(n7863), .ZN(n7862) );
  OAI21_X1 U7822 ( .B1(n8622), .B2(n7864), .A(n8633), .ZN(n7863) );
  INV_X1 U7823 ( .A(n8214), .ZN(n7864) );
  AND2_X1 U7824 ( .A1(n8519), .A2(n8539), .ZN(n7496) );
  OR2_X1 U7825 ( .A1(n8458), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8516) );
  INV_X1 U7826 ( .A(n8423), .ZN(n7556) );
  INV_X1 U7827 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U7828 ( .A1(n7538), .A2(n9643), .ZN(n7534) );
  NAND2_X1 U7829 ( .A1(n7539), .A2(n7540), .ZN(n7537) );
  NOR2_X1 U7830 ( .A1(n12116), .A2(n9643), .ZN(n7535) );
  NAND2_X1 U7831 ( .A1(n9690), .A2(n9660), .ZN(n9679) );
  NAND2_X1 U7832 ( .A1(n9638), .A2(n9694), .ZN(n9699) );
  OR2_X1 U7833 ( .A1(n14365), .A2(n14153), .ZN(n9638) );
  AOI21_X1 U7834 ( .B1(n7928), .B2(n14185), .A(n7926), .ZN(n7925) );
  INV_X1 U7835 ( .A(n9394), .ZN(n7926) );
  NAND2_X1 U7836 ( .A1(n8891), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n9276) );
  INV_X1 U7837 ( .A(n9260), .ZN(n8891) );
  NAND2_X1 U7838 ( .A1(n14407), .A2(n14065), .ZN(n7431) );
  NOR2_X1 U7839 ( .A1(n9385), .A2(n7940), .ZN(n7939) );
  AND2_X1 U7840 ( .A1(n14433), .A2(n14321), .ZN(n9385) );
  INV_X1 U7841 ( .A(n8143), .ZN(n7940) );
  INV_X1 U7842 ( .A(n9553), .ZN(n7894) );
  OR2_X1 U7843 ( .A1(n11507), .A2(n9141), .ZN(n7913) );
  INV_X1 U7844 ( .A(n11290), .ZN(n7836) );
  OR2_X1 U7845 ( .A1(n14928), .A2(n10467), .ZN(n10312) );
  NOR2_X1 U7846 ( .A1(n15324), .A2(n7971), .ZN(n7970) );
  INV_X1 U7847 ( .A(n12722), .ZN(n7971) );
  NOR2_X1 U7848 ( .A1(n12209), .A2(n7989), .ZN(n7988) );
  INV_X1 U7849 ( .A(n12179), .ZN(n7989) );
  OAI21_X1 U7850 ( .B1(n11969), .B2(n7958), .A(n14964), .ZN(n7957) );
  AND2_X1 U7851 ( .A1(n11592), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11603) );
  NOR2_X1 U7852 ( .A1(n11567), .A2(n11564), .ZN(n7962) );
  INV_X1 U7853 ( .A(n11127), .ZN(n7964) );
  AND2_X1 U7854 ( .A1(n7961), .A2(n10829), .ZN(n7960) );
  INV_X1 U7855 ( .A(n7962), .ZN(n7961) );
  INV_X1 U7856 ( .A(n11130), .ZN(n7500) );
  NAND2_X1 U7857 ( .A1(n14607), .A2(n15775), .ZN(n10329) );
  OR2_X2 U7858 ( .A1(n15054), .A2(n10771), .ZN(n14765) );
  NAND2_X2 U7859 ( .A1(n14757), .A2(n14935), .ZN(n14758) );
  NAND2_X1 U7860 ( .A1(n15263), .A2(n15262), .ZN(n15261) );
  INV_X1 U7861 ( .A(n14960), .ZN(n7979) );
  AND2_X1 U7862 ( .A1(n7187), .A2(n10342), .ZN(n10462) );
  INV_X1 U7863 ( .A(n11321), .ZN(n14951) );
  INV_X1 U7864 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9994) );
  INV_X1 U7865 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9993) );
  CLKBUF_X1 U7866 ( .A(n10134), .Z(n9995) );
  NAND2_X1 U7867 ( .A1(n8017), .A2(n8850), .ZN(n9300) );
  NAND2_X1 U7868 ( .A1(n9287), .A2(n8849), .ZN(n8017) );
  NOR2_X1 U7869 ( .A1(n8842), .A2(n7657), .ZN(n7656) );
  INV_X1 U7870 ( .A(n8837), .ZN(n7657) );
  NAND2_X1 U7871 ( .A1(n9992), .A2(n7396), .ZN(n8131) );
  XNOR2_X1 U7872 ( .A(n9204), .B(n13291), .ZN(n9201) );
  AND2_X1 U7873 ( .A1(n8823), .A2(n8822), .ZN(n9182) );
  INV_X1 U7874 ( .A(n8030), .ZN(n7627) );
  INV_X1 U7875 ( .A(n8811), .ZN(n8035) );
  INV_X1 U7876 ( .A(n9157), .ZN(n7363) );
  NOR2_X1 U7877 ( .A1(n9127), .A2(n8044), .ZN(n8043) );
  INV_X1 U7878 ( .A(n8794), .ZN(n8044) );
  INV_X1 U7879 ( .A(n8972), .ZN(n8016) );
  INV_X1 U7880 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7714) );
  XNOR2_X1 U7881 ( .A(n9864), .B(n9865), .ZN(n9910) );
  NAND2_X1 U7882 ( .A1(n7241), .A2(n7331), .ZN(n8001) );
  AND2_X1 U7883 ( .A1(n12246), .A2(n12243), .ZN(n9762) );
  OR2_X1 U7884 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  INV_X1 U7885 ( .A(n11427), .ZN(n7472) );
  AND2_X1 U7886 ( .A1(n8003), .A2(n7474), .ZN(n7473) );
  AND2_X1 U7887 ( .A1(n9965), .A2(n9809), .ZN(n13184) );
  AND2_X1 U7888 ( .A1(n9801), .A2(n9800), .ZN(n13205) );
  AND2_X1 U7889 ( .A1(n7454), .A2(n7453), .ZN(n11239) );
  NAND2_X1 U7890 ( .A1(n9752), .A2(n13485), .ZN(n7453) );
  INV_X1 U7891 ( .A(n7464), .ZN(n7463) );
  INV_X1 U7892 ( .A(n12409), .ZN(n7991) );
  INV_X1 U7893 ( .A(n7996), .ZN(n7995) );
  AOI21_X1 U7894 ( .B1(n12317), .B2(n7997), .A(n9771), .ZN(n7996) );
  INV_X1 U7895 ( .A(n9765), .ZN(n7997) );
  NAND2_X1 U7896 ( .A1(n9799), .A2(n7460), .ZN(n13224) );
  OR2_X1 U7897 ( .A1(n13224), .A2(n13743), .ZN(n13225) );
  NAND2_X1 U7898 ( .A1(n7204), .A2(n9744), .ZN(n9746) );
  AND2_X1 U7899 ( .A1(n7492), .A2(n12481), .ZN(n7491) );
  INV_X1 U7900 ( .A(n9787), .ZN(n7488) );
  NAND2_X1 U7901 ( .A1(n7492), .A2(n7284), .ZN(n7490) );
  NOR2_X1 U7902 ( .A1(n11854), .A2(n8006), .ZN(n8005) );
  INV_X1 U7903 ( .A(n9757), .ZN(n8006) );
  NAND2_X1 U7904 ( .A1(n11427), .A2(n11428), .ZN(n11426) );
  OR2_X1 U7905 ( .A1(n13012), .A2(n9732), .ZN(n10890) );
  OR2_X1 U7906 ( .A1(n12873), .A2(n8737), .ZN(n10004) );
  NAND2_X1 U7907 ( .A1(n10707), .A2(n7268), .ZN(n10735) );
  XNOR2_X1 U7908 ( .A(n11545), .B(n11541), .ZN(n11546) );
  OR2_X1 U7909 ( .A1(n11549), .A2(n11538), .ZN(n7731) );
  NAND2_X1 U7910 ( .A1(n12285), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7735) );
  NOR2_X1 U7911 ( .A1(n12284), .A2(n7566), .ZN(n12286) );
  NAND2_X1 U7912 ( .A1(n15707), .A2(n12307), .ZN(n12308) );
  AOI21_X1 U7913 ( .B1(n13536), .B2(n13535), .A(n13534), .ZN(n13538) );
  OR2_X1 U7914 ( .A1(n7756), .A2(n13075), .ZN(n7755) );
  AOI22_X1 U7915 ( .A1(n13660), .A2(n8646), .B1(n8699), .B2(n13651), .ZN(
        n13650) );
  AOI21_X1 U7916 ( .B1(n13664), .B2(n13665), .A(n8700), .ZN(n13647) );
  AND3_X1 U7917 ( .A1(n8551), .A2(n8550), .A3(n8549), .ZN(n13800) );
  INV_X1 U7918 ( .A(n13260), .ZN(n13834) );
  NAND2_X1 U7919 ( .A1(n8494), .A2(n8493), .ZN(n13826) );
  AOI21_X1 U7920 ( .B1(n7762), .B2(n12952), .A(n12961), .ZN(n7759) );
  INV_X1 U7921 ( .A(n7763), .ZN(n7762) );
  OAI21_X1 U7922 ( .B1(n12044), .B2(n8683), .A(n12939), .ZN(n12254) );
  AOI21_X1 U7923 ( .B1(n7767), .B2(n11669), .A(n7766), .ZN(n7765) );
  OR2_X1 U7924 ( .A1(n8355), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8357) );
  AND2_X1 U7925 ( .A1(n8744), .A2(n8743), .ZN(n10895) );
  NAND2_X1 U7926 ( .A1(n13862), .A2(n8695), .ZN(n13689) );
  INV_X1 U7927 ( .A(n13742), .ZN(n13835) );
  AND2_X1 U7928 ( .A1(n12919), .A2(n12920), .ZN(n13055) );
  NAND2_X1 U7929 ( .A1(n11500), .A2(n13055), .ZN(n11502) );
  OR2_X1 U7930 ( .A1(n13083), .A2(n9734), .ZN(n13756) );
  OR2_X1 U7931 ( .A1(n8747), .A2(n13092), .ZN(n15912) );
  NAND2_X1 U7932 ( .A1(n13023), .A2(n13024), .ZN(n7869) );
  AND2_X1 U7933 ( .A1(n8217), .A2(n8219), .ZN(n7686) );
  INV_X1 U7934 ( .A(n13020), .ZN(n13023) );
  AOI21_X1 U7935 ( .B1(n13018), .B2(n13019), .A(n7843), .ZN(n13020) );
  AND2_X1 U7936 ( .A1(n14946), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7843) );
  NAND2_X1 U7937 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7848), .ZN(n7847) );
  INV_X1 U7938 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8217) );
  INV_X1 U7939 ( .A(n8670), .ZN(n10977) );
  NAND2_X1 U7940 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n12670), .ZN(n8214) );
  AND4_X1 U7941 ( .A1(n8167), .A2(n8665), .A3(n8710), .A4(n8010), .ZN(n8168)
         );
  NOR2_X1 U7942 ( .A1(n8607), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8212) );
  AND2_X1 U7943 ( .A1(n8441), .A2(n8008), .ZN(n8740) );
  AND2_X1 U7944 ( .A1(n8012), .A2(n8009), .ZN(n8008) );
  AND2_X1 U7945 ( .A1(n8665), .A2(n8010), .ZN(n8009) );
  NOR2_X1 U7946 ( .A1(n8574), .A2(n8573), .ZN(n8211) );
  OR2_X1 U7947 ( .A1(n8554), .A2(n12609), .ZN(n7870) );
  XNOR2_X1 U7948 ( .A(n8207), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n8554) );
  AND2_X1 U7949 ( .A1(n7545), .A2(n7871), .ZN(n7544) );
  NAND2_X1 U7950 ( .A1(n7337), .A2(n8204), .ZN(n7871) );
  NAND2_X1 U7951 ( .A1(n7330), .A2(n7546), .ZN(n7545) );
  INV_X1 U7952 ( .A(n7330), .ZN(n7547) );
  NAND2_X1 U7953 ( .A1(n8201), .A2(n8200), .ZN(n8485) );
  OAI21_X1 U7954 ( .B1(n8437), .B2(n7842), .A(n7839), .ZN(n8199) );
  AOI21_X1 U7955 ( .B1(n7852), .B2(n7854), .A(n7293), .ZN(n7849) );
  NAND2_X1 U7956 ( .A1(n8193), .A2(n8192), .ZN(n8406) );
  XNOR2_X1 U7957 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n8249) );
  XNOR2_X1 U7958 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8340) );
  XNOR2_X1 U7959 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8314) );
  XNOR2_X1 U7960 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8299) );
  NAND2_X1 U7961 ( .A1(n8178), .A2(n8177), .ZN(n8300) );
  OR2_X1 U7962 ( .A1(n8297), .A2(n8708), .ZN(n8298) );
  NOR3_X1 U7963 ( .A1(n12391), .A2(n12158), .A3(n12161), .ZN(n9976) );
  NAND2_X1 U7964 ( .A1(n8892), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9290) );
  INV_X1 U7965 ( .A(n9276), .ZN(n8892) );
  NOR2_X1 U7966 ( .A1(n7890), .A2(n7889), .ZN(n7888) );
  INV_X1 U7967 ( .A(n12499), .ZN(n7889) );
  AND2_X1 U7968 ( .A1(n13139), .A2(n11795), .ZN(n11796) );
  NAND2_X1 U7969 ( .A1(n7531), .A2(n7252), .ZN(n7883) );
  OAI21_X1 U7970 ( .B1(n10272), .B2(n10218), .A(n7419), .ZN(n10262) );
  NAND2_X1 U7971 ( .A1(n10272), .A2(n10218), .ZN(n7419) );
  NOR2_X1 U7972 ( .A1(n12099), .A2(n7599), .ZN(n15579) );
  AND2_X1 U7973 ( .A1(n12100), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7599) );
  NAND2_X1 U7974 ( .A1(n14109), .A2(n7417), .ZN(n14116) );
  NOR2_X1 U7975 ( .A1(n7349), .A2(n7418), .ZN(n7417) );
  NOR2_X1 U7976 ( .A1(n14127), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U7977 ( .A1(n7910), .A2(n9312), .ZN(n7906) );
  INV_X1 U7978 ( .A(n7908), .ZN(n7907) );
  OAI21_X1 U7979 ( .B1(n14205), .B2(n7909), .A(n9329), .ZN(n7908) );
  OR2_X1 U7980 ( .A1(n7579), .A2(n14392), .ZN(n7578) );
  NAND2_X1 U7981 ( .A1(n14190), .A2(n14355), .ZN(n7407) );
  OR2_X1 U7982 ( .A1(n14396), .A2(n14064), .ZN(n9298) );
  INV_X1 U7983 ( .A(n9709), .ZN(n14205) );
  OAI21_X1 U7984 ( .B1(n14237), .B2(n7942), .A(n7941), .ZN(n7945) );
  INV_X1 U7985 ( .A(n7943), .ZN(n7942) );
  AOI21_X1 U7986 ( .B1(n14241), .B2(n7943), .A(n9391), .ZN(n7941) );
  NAND2_X1 U7987 ( .A1(n14237), .A2(n14236), .ZN(n14235) );
  NAND2_X1 U7988 ( .A1(n7206), .A2(n7243), .ZN(n7901) );
  NAND2_X1 U7989 ( .A1(n7952), .A2(n7208), .ZN(n7951) );
  INV_X1 U7990 ( .A(n14300), .ZN(n7952) );
  NAND2_X1 U7991 ( .A1(n7300), .A2(n7208), .ZN(n7950) );
  NAND2_X1 U7992 ( .A1(n14296), .A2(n14300), .ZN(n14295) );
  NAND2_X1 U7993 ( .A1(n7586), .A2(n7585), .ZN(n14306) );
  INV_X1 U7994 ( .A(n14424), .ZN(n7585) );
  OR2_X1 U7995 ( .A1(n14299), .A2(n14300), .ZN(n7953) );
  OR2_X1 U7996 ( .A1(n12473), .A2(n14354), .ZN(n8143) );
  NAND2_X1 U7997 ( .A1(n14340), .A2(n14350), .ZN(n14341) );
  NAND2_X1 U7998 ( .A1(n12474), .A2(n7260), .ZN(n14339) );
  NOR2_X1 U7999 ( .A1(n12396), .A2(n7448), .ZN(n7446) );
  OR2_X1 U8000 ( .A1(n12126), .A2(n12393), .ZN(n7365) );
  OR2_X1 U8001 ( .A1(n9381), .A2(n14070), .ZN(n8144) );
  NAND2_X1 U8002 ( .A1(n11952), .A2(n11951), .ZN(n11950) );
  NAND2_X1 U8003 ( .A1(n11508), .A2(n7211), .ZN(n7918) );
  NAND2_X1 U8004 ( .A1(n7299), .A2(n7916), .ZN(n7915) );
  INV_X1 U8005 ( .A(n12052), .ZN(n7917) );
  OAI21_X1 U8006 ( .B1(n11339), .B2(n11342), .A(n7936), .ZN(n11354) );
  AND2_X1 U8007 ( .A1(n11340), .A2(n11342), .ZN(n9110) );
  INV_X1 U8008 ( .A(n9701), .ZN(n11386) );
  XNOR2_X1 U8009 ( .A(n15840), .B(n11011), .ZN(n9093) );
  NAND2_X1 U8010 ( .A1(n11454), .A2(n11463), .ZN(n7893) );
  INV_X1 U8011 ( .A(n9093), .ZN(n11202) );
  NAND2_X1 U8012 ( .A1(n11466), .A2(n9375), .ZN(n11194) );
  INV_X1 U8013 ( .A(n14322), .ZN(n14355) );
  NAND2_X1 U8014 ( .A1(n9369), .A2(n9368), .ZN(n10442) );
  NAND2_X1 U8015 ( .A1(n10542), .A2(n10855), .ZN(n10783) );
  OR2_X1 U8016 ( .A1(n11172), .A2(n11171), .ZN(n11185) );
  NAND2_X1 U8017 ( .A1(n9645), .A2(n9644), .ZN(n14369) );
  NAND2_X1 U8018 ( .A1(n9316), .A2(n9315), .ZN(n14386) );
  OR2_X1 U8019 ( .A1(n9430), .A2(n12391), .ZN(n9441) );
  XNOR2_X1 U8020 ( .A(n8902), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8905) );
  NAND2_X1 U8021 ( .A1(n7954), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U8022 ( .A1(n9422), .A2(n9421), .ZN(n9427) );
  OAI21_X1 U8023 ( .B1(n9433), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9425) );
  XNOR2_X1 U8024 ( .A(n9435), .B(n9434), .ZN(n10224) );
  NAND2_X1 U8025 ( .A1(n8985), .A2(n10417), .ZN(n9013) );
  AOI21_X1 U8026 ( .B1(n7794), .B2(n7797), .A(n7297), .ZN(n7793) );
  INV_X1 U8027 ( .A(n14730), .ZN(n7797) );
  OAI22_X1 U8028 ( .A1(n11416), .A2(n7835), .B1(n11301), .B2(n11302), .ZN(
        n7834) );
  INV_X1 U8029 ( .A(n11289), .ZN(n7835) );
  NAND2_X1 U8030 ( .A1(n12207), .A2(n12206), .ZN(n14845) );
  NAND2_X1 U8031 ( .A1(n11639), .A2(n11640), .ZN(n7837) );
  AND2_X1 U8032 ( .A1(n7235), .A2(n7837), .ZN(n7828) );
  NOR2_X1 U8033 ( .A1(n7834), .A2(n11304), .ZN(n7832) );
  INV_X1 U8034 ( .A(n14540), .ZN(n7813) );
  AND2_X1 U8035 ( .A1(n14547), .A2(n7811), .ZN(n7810) );
  AND2_X1 U8036 ( .A1(n14701), .A2(n14702), .ZN(n14547) );
  NAND2_X1 U8037 ( .A1(n7812), .A2(n14540), .ZN(n7811) );
  INV_X1 U8038 ( .A(n14532), .ZN(n7812) );
  AOI21_X1 U8039 ( .B1(n11909), .B2(n11908), .A(n7800), .ZN(n11910) );
  AND2_X1 U8040 ( .A1(n11906), .A2(n11907), .ZN(n7800) );
  NAND2_X1 U8041 ( .A1(n12777), .A2(n12778), .ZN(n12776) );
  AOI21_X1 U8042 ( .B1(n7818), .B2(n12425), .A(n7816), .ZN(n7815) );
  AND4_X1 U8043 ( .A1(n11983), .A2(n11982), .A3(n11981), .A4(n11980), .ZN(
        n12268) );
  NOR2_X1 U8044 ( .A1(n8022), .A2(n14929), .ZN(n8019) );
  NOR2_X1 U8045 ( .A1(n8023), .A2(n8025), .ZN(n8022) );
  INV_X1 U8046 ( .A(n8026), .ZN(n8023) );
  NAND2_X1 U8047 ( .A1(n8026), .A2(n8028), .ZN(n8024) );
  NAND2_X1 U8048 ( .A1(n14932), .A2(n14931), .ZN(n15146) );
  OR2_X1 U8049 ( .A1(n14930), .A2(n14929), .ZN(n14932) );
  NOR2_X1 U8050 ( .A1(n15378), .A2(n7610), .ZN(n7609) );
  INV_X1 U8051 ( .A(n7611), .ZN(n7610) );
  AOI21_X1 U8052 ( .B1(n7505), .B2(n7506), .A(n8103), .ZN(n7502) );
  AND2_X1 U8053 ( .A1(n15224), .A2(n7983), .ZN(n7980) );
  NAND2_X1 U8054 ( .A1(n15261), .A2(n8106), .ZN(n15239) );
  CLKBUF_X1 U8055 ( .A(n15254), .Z(n7412) );
  NAND2_X1 U8056 ( .A1(n15276), .A2(n15275), .ZN(n15274) );
  NAND2_X1 U8057 ( .A1(n15305), .A2(n12620), .ZN(n15288) );
  NAND2_X1 U8058 ( .A1(n7975), .A2(n7974), .ZN(n7973) );
  NAND2_X1 U8059 ( .A1(n12723), .A2(n7970), .ZN(n7969) );
  AOI21_X1 U8060 ( .B1(n8094), .B2(n12347), .A(n7282), .ZN(n7513) );
  OR2_X1 U8061 ( .A1(n12333), .A2(n7514), .ZN(n7512) );
  INV_X1 U8062 ( .A(n8094), .ZN(n7514) );
  AOI21_X1 U8063 ( .B1(n12030), .B2(n7253), .A(n7985), .ZN(n12720) );
  NAND2_X1 U8064 ( .A1(n12351), .A2(n7986), .ZN(n7985) );
  OR2_X1 U8065 ( .A1(n15982), .A2(n15040), .ZN(n12346) );
  NAND2_X1 U8066 ( .A1(n15974), .A2(n7988), .ZN(n12354) );
  AND2_X1 U8067 ( .A1(n11997), .A2(n11746), .ZN(n14962) );
  NOR2_X1 U8068 ( .A1(n7226), .A2(n8098), .ZN(n8097) );
  INV_X1 U8069 ( .A(n11621), .ZN(n8098) );
  XNOR2_X1 U8070 ( .A(n14796), .B(n11617), .ZN(n14958) );
  NAND2_X1 U8071 ( .A1(n11685), .A2(n10811), .ZN(n10821) );
  NAND2_X1 U8072 ( .A1(n10821), .A2(n10829), .ZN(n11128) );
  AND2_X1 U8073 ( .A1(n14755), .A2(n14940), .ZN(n11263) );
  AOI211_X1 U8074 ( .C1(n15372), .C2(n15981), .A(n15371), .B(n15370), .ZN(
        n15373) );
  NAND2_X1 U8075 ( .A1(n15182), .A2(n15988), .ZN(n15376) );
  AND2_X1 U8076 ( .A1(n10820), .A2(n10819), .ZN(n11129) );
  NAND2_X1 U8077 ( .A1(n11328), .A2(n15875), .ZN(n15973) );
  AND2_X1 U8078 ( .A1(n11263), .A2(n7187), .ZN(n15932) );
  OR2_X1 U8079 ( .A1(n10479), .A2(P1_U3086), .ZN(n15012) );
  NOR2_X1 U8080 ( .A1(n10282), .A2(n10281), .ZN(n15472) );
  NAND2_X1 U8081 ( .A1(n7633), .A2(n7632), .ZN(n9640) );
  AOI21_X1 U8082 ( .B1(n7635), .B2(n7637), .A(n7346), .ZN(n7632) );
  OR2_X1 U8083 ( .A1(n9640), .A2(n9639), .ZN(n9642) );
  XNOR2_X1 U8084 ( .A(n9622), .B(n9621), .ZN(n14945) );
  NAND2_X1 U8085 ( .A1(n7634), .A2(n9341), .ZN(n9622) );
  NAND2_X1 U8086 ( .A1(n9995), .A2(n10112), .ZN(n9996) );
  INV_X1 U8087 ( .A(n9996), .ZN(n7806) );
  NOR2_X1 U8088 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n7805) );
  INV_X1 U8089 ( .A(n9995), .ZN(n9999) );
  NAND2_X1 U8090 ( .A1(n7648), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U8091 ( .A1(n9961), .A2(n7647), .ZN(n8045) );
  XNOR2_X1 U8092 ( .A(n9911), .B(n7403), .ZN(n9912) );
  INV_X1 U8093 ( .A(n9914), .ZN(n7403) );
  XNOR2_X1 U8094 ( .A(n9910), .B(n7694), .ZN(n9921) );
  AOI22_X1 U8095 ( .A1(n9924), .A2(n9871), .B1(P1_ADDR_REG_5__SCAN_IN), .B2(
        n9870), .ZN(n9929) );
  AND2_X1 U8096 ( .A1(n9933), .A2(n15617), .ZN(n9934) );
  AND2_X1 U8097 ( .A1(n7689), .A2(n15641), .ZN(n9946) );
  OAI21_X1 U8098 ( .B1(n15642), .B2(n15643), .A(n7690), .ZN(n7689) );
  AND4_X1 U8099 ( .A1(n8532), .A2(n8531), .A3(n8530), .A4(n8529), .ZN(n13808)
         );
  OAI22_X1 U8100 ( .A1(n12570), .A2(n12571), .B1(n13808), .B2(n9788), .ZN(
        n13169) );
  NAND2_X1 U8101 ( .A1(n8543), .A2(n8542), .ZN(n13784) );
  XNOR2_X1 U8102 ( .A(n7479), .B(n9749), .ZN(n10685) );
  XNOR2_X1 U8103 ( .A(n10572), .B(n9748), .ZN(n7479) );
  AND2_X1 U8104 ( .A1(n8584), .A2(n8583), .ZN(n13710) );
  AND4_X1 U8105 ( .A1(n8248), .A2(n8247), .A3(n8246), .A4(n8245), .ZN(n12892)
         );
  INV_X1 U8106 ( .A(n13487), .ZN(n10572) );
  INV_X1 U8107 ( .A(n13879), .ZN(n13219) );
  AND4_X1 U8108 ( .A1(n8399), .A2(n8398), .A3(n8397), .A4(n8396), .ZN(n12379)
         );
  AND2_X1 U8109 ( .A1(n8421), .A2(n8420), .ZN(n12324) );
  INV_X1 U8110 ( .A(n13691), .ZN(n13662) );
  AOI21_X1 U8111 ( .B1(n13085), .B2(n9732), .A(n7280), .ZN(n7386) );
  XNOR2_X1 U8112 ( .A(n8271), .B(n7572), .ZN(n10524) );
  NAND2_X1 U8113 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7572) );
  XNOR2_X1 U8114 ( .A(n12308), .B(n7566), .ZN(n13490) );
  NAND2_X1 U8115 ( .A1(n13490), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n13489) );
  OR2_X1 U8116 ( .A1(n13529), .A2(n13530), .ZN(n7717) );
  INV_X1 U8117 ( .A(n7565), .ZN(n13543) );
  INV_X1 U8118 ( .A(n7563), .ZN(n13563) );
  AND2_X1 U8119 ( .A1(n7717), .A2(n7716), .ZN(n13552) );
  INV_X1 U8120 ( .A(n13531), .ZN(n7716) );
  XNOR2_X1 U8121 ( .A(n13570), .B(n7561), .ZN(n13553) );
  INV_X1 U8122 ( .A(n13612), .ZN(n7567) );
  NAND2_X1 U8123 ( .A1(n7380), .A2(n7379), .ZN(n7737) );
  NAND2_X1 U8124 ( .A1(n7741), .A2(n13597), .ZN(n7379) );
  OR2_X1 U8125 ( .A1(n7741), .A2(n7739), .ZN(n7380) );
  OR2_X1 U8126 ( .A1(n7741), .A2(n13601), .ZN(n7740) );
  AOI21_X1 U8127 ( .B1(n13974), .B2(n13028), .A(n13027), .ZN(n16003) );
  NOR2_X1 U8128 ( .A1(n8675), .A2(n8674), .ZN(n8676) );
  NAND2_X1 U8129 ( .A1(n8589), .A2(n8588), .ZN(n13873) );
  NAND2_X1 U8130 ( .A1(n11146), .A2(n8706), .ZN(n13084) );
  AND3_X1 U8131 ( .A1(n8331), .A2(n8330), .A3(n8329), .ZN(n11255) );
  NOR2_X1 U8132 ( .A1(n13622), .A2(n8707), .ZN(n9742) );
  AND2_X1 U8133 ( .A1(n13627), .A2(n15917), .ZN(n8707) );
  AND2_X1 U8134 ( .A1(n8429), .A2(n8428), .ZN(n12566) );
  NAND2_X1 U8135 ( .A1(n16000), .A2(n15865), .ZN(n13960) );
  NAND2_X1 U8136 ( .A1(n7883), .A2(n7884), .ZN(n13985) );
  AOI21_X1 U8137 ( .B1(n7884), .B2(n7882), .A(n12835), .ZN(n7881) );
  INV_X1 U8138 ( .A(n7252), .ZN(n7882) );
  NAND2_X1 U8139 ( .A1(n8980), .A2(n8979), .ZN(n12854) );
  AOI21_X1 U8140 ( .B1(n12737), .B2(n12499), .A(n12738), .ZN(n12746) );
  NAND2_X1 U8141 ( .A1(n9163), .A2(n9162), .ZN(n12134) );
  NAND2_X1 U8142 ( .A1(n7541), .A2(n9133), .ZN(n11879) );
  AND2_X1 U8143 ( .A1(n8051), .A2(n8050), .ZN(n8056) );
  NOR2_X1 U8144 ( .A1(n12202), .A2(n9722), .ZN(n8050) );
  NAND2_X1 U8145 ( .A1(n7219), .A2(n8058), .ZN(n8051) );
  INV_X1 U8146 ( .A(n8058), .ZN(n8057) );
  OAI21_X1 U8147 ( .B1(n9724), .B2(n12202), .A(n9729), .ZN(n8054) );
  NAND2_X1 U8148 ( .A1(n9311), .A2(n9310), .ZN(n14221) );
  NAND2_X1 U8149 ( .A1(n9250), .A2(n9249), .ZN(n14251) );
  NAND2_X1 U8150 ( .A1(n9199), .A2(n9198), .ZN(n14356) );
  INV_X1 U8151 ( .A(n7597), .ZN(n15562) );
  OAI22_X1 U8152 ( .A1(n7435), .A2(n9395), .B1(n9712), .B2(n7207), .ZN(n7434)
         );
  OR2_X1 U8153 ( .A1(n14379), .A2(n7321), .ZN(n7439) );
  AND2_X1 U8154 ( .A1(n14379), .A2(n7440), .ZN(n14164) );
  NAND2_X1 U8155 ( .A1(n7929), .A2(n7928), .ZN(n14166) );
  NAND2_X1 U8156 ( .A1(n7369), .A2(n12836), .ZN(n7368) );
  NAND2_X1 U8157 ( .A1(n8880), .A2(n8879), .ZN(n14373) );
  NAND2_X1 U8158 ( .A1(n9240), .A2(n9239), .ZN(n14413) );
  NAND2_X1 U8159 ( .A1(n10011), .A2(n14445), .ZN(n14308) );
  INV_X1 U8160 ( .A(n12163), .ZN(n10002) );
  AND4_X1 U8161 ( .A1(n12696), .A2(n12695), .A3(n12694), .A4(n12693), .ZN(
        n15194) );
  NAND2_X1 U8162 ( .A1(n11815), .A2(n7801), .ZN(n11909) );
  NAND2_X1 U8163 ( .A1(n11814), .A2(n7802), .ZN(n7801) );
  INV_X1 U8164 ( .A(n11816), .ZN(n7802) );
  INV_X1 U8165 ( .A(n11129), .ZN(n14787) );
  AND4_X1 U8166 ( .A1(n12680), .A2(n12679), .A3(n12678), .A4(n12677), .ZN(
        n14733) );
  NAND2_X1 U8167 ( .A1(n12684), .A2(n12683), .ZN(n15392) );
  AND2_X1 U8168 ( .A1(n8015), .A2(n7643), .ZN(n14994) );
  INV_X1 U8169 ( .A(n15023), .ZN(n7643) );
  INV_X1 U8170 ( .A(n14705), .ZN(n15272) );
  AOI21_X1 U8171 ( .B1(n12718), .B2(n15988), .A(n12717), .ZN(n15384) );
  NAND2_X1 U8172 ( .A1(n12657), .A2(n12656), .ZN(n15250) );
  NAND2_X1 U8173 ( .A1(n11132), .A2(n14953), .ZN(n11568) );
  XNOR2_X1 U8174 ( .A(n9912), .B(n9913), .ZN(n15673) );
  OR2_X1 U8175 ( .A1(n15667), .A2(n15668), .ZN(n7693) );
  NAND2_X1 U8176 ( .A1(n7416), .A2(n7415), .ZN(n15622) );
  INV_X1 U8177 ( .A(n9935), .ZN(n7415) );
  INV_X1 U8178 ( .A(n9934), .ZN(n7416) );
  OR2_X1 U8179 ( .A1(n15636), .A2(n15635), .ZN(n7697) );
  XNOR2_X1 U8180 ( .A(n7404), .B(n9943), .ZN(n15640) );
  NAND2_X1 U8181 ( .A1(n15640), .A2(n15639), .ZN(n15638) );
  INV_X1 U8182 ( .A(n15652), .ZN(n7401) );
  NAND2_X1 U8183 ( .A1(n14794), .A2(n8120), .ZN(n8119) );
  NAND2_X1 U8184 ( .A1(n14805), .A2(n14807), .ZN(n8130) );
  NAND2_X1 U8185 ( .A1(n14816), .A2(n8113), .ZN(n8112) );
  NAND2_X1 U8186 ( .A1(n9479), .A2(n8072), .ZN(n8071) );
  INV_X1 U8187 ( .A(n9482), .ZN(n8072) );
  NAND2_X1 U8188 ( .A1(n8126), .A2(n14826), .ZN(n8125) );
  NAND2_X1 U8189 ( .A1(n9504), .A2(n7310), .ZN(n8075) );
  AND2_X1 U8190 ( .A1(n8078), .A2(n8077), .ZN(n8076) );
  NAND2_X1 U8191 ( .A1(n14843), .A2(n8115), .ZN(n8114) );
  NAND2_X1 U8192 ( .A1(n7229), .A2(n8089), .ZN(n8088) );
  NAND2_X1 U8193 ( .A1(n8123), .A2(n14862), .ZN(n8122) );
  NAND2_X1 U8194 ( .A1(n8073), .A2(n7220), .ZN(n7372) );
  NAND2_X1 U8195 ( .A1(n9564), .A2(n7334), .ZN(n8062) );
  OAI21_X1 U8196 ( .B1(n9559), .B2(n9558), .A(n7262), .ZN(n8063) );
  NAND2_X1 U8197 ( .A1(n8117), .A2(n14878), .ZN(n8116) );
  NAND2_X1 U8198 ( .A1(n8081), .A2(n7333), .ZN(n8080) );
  AOI21_X1 U8199 ( .B1(n12890), .B2(n12889), .A(n13075), .ZN(n13006) );
  NAND2_X1 U8200 ( .A1(n14901), .A2(n14899), .ZN(n8128) );
  NOR2_X1 U8201 ( .A1(n8855), .A2(n7641), .ZN(n7640) );
  INV_X1 U8202 ( .A(n8854), .ZN(n7641) );
  NAND2_X1 U8203 ( .A1(n8778), .A2(n9051), .ZN(n8776) );
  OR2_X1 U8204 ( .A1(n9813), .A2(n9966), .ZN(n9815) );
  INV_X1 U8205 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8800) );
  INV_X1 U8206 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U8207 ( .A1(n9408), .A2(n14183), .ZN(n7583) );
  INV_X1 U8208 ( .A(n7654), .ZN(n7653) );
  OAI21_X1 U8209 ( .B1(n7656), .B2(n7655), .A(n8844), .ZN(n7654) );
  AOI21_X1 U8210 ( .B1(n8030), .B2(n8034), .A(n7626), .ZN(n7625) );
  INV_X1 U8211 ( .A(n8927), .ZN(n7626) );
  NOR2_X1 U8212 ( .A1(n8961), .A2(n8037), .ZN(n8036) );
  INV_X1 U8213 ( .A(n8806), .ZN(n8037) );
  AOI21_X1 U8214 ( .B1(n7528), .B2(n7530), .A(n7292), .ZN(n7525) );
  INV_X1 U8215 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n9865) );
  OAI21_X1 U8216 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n9890), .A(n9889), .ZN(
        n9892) );
  OR2_X1 U8217 ( .A1(n7212), .A2(n7476), .ZN(n7470) );
  OAI21_X1 U8218 ( .B1(n8003), .B2(n7470), .A(n7465), .ZN(n7464) );
  INV_X1 U8219 ( .A(n7466), .ZN(n7465) );
  OAI21_X1 U8220 ( .B1(n7470), .B2(n7474), .A(n7469), .ZN(n7466) );
  OR2_X1 U8221 ( .A1(n7476), .A2(n12082), .ZN(n7469) );
  AND2_X1 U8222 ( .A1(n8505), .A2(n13360), .ZN(n8524) );
  NOR2_X1 U8223 ( .A1(n13013), .A2(n13002), .ZN(n13014) );
  OR2_X1 U8224 ( .A1(n7749), .A2(n13647), .ZN(n7747) );
  AOI21_X1 U8225 ( .B1(n7750), .B2(n13649), .A(n7289), .ZN(n7748) );
  NAND2_X1 U8226 ( .A1(n10656), .A2(n10598), .ZN(n7718) );
  NAND2_X1 U8227 ( .A1(n7723), .A2(n10656), .ZN(n7726) );
  AND2_X1 U8228 ( .A1(n7563), .A2(n7562), .ZN(n13585) );
  NAND2_X1 U8229 ( .A1(n13564), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7562) );
  INV_X1 U8230 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n13446) );
  NOR2_X1 U8231 ( .A1(n8638), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8227) );
  AND2_X1 U8232 ( .A1(n8577), .A2(n13227), .ZN(n8565) );
  OAI21_X1 U8233 ( .B1(n12549), .B2(n12952), .A(n13065), .ZN(n7763) );
  NAND2_X1 U8234 ( .A1(n7679), .A2(n7681), .ZN(n7676) );
  OAI21_X1 U8235 ( .B1(n8562), .B2(n8561), .A(n7557), .ZN(n7387) );
  NAND2_X1 U8236 ( .A1(n10754), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7557) );
  INV_X1 U8237 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8665) );
  INV_X1 U8238 ( .A(n8202), .ZN(n7872) );
  INV_X1 U8239 ( .A(n8200), .ZN(n7546) );
  INV_X1 U8240 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U8241 ( .A1(n7551), .A2(n8326), .ZN(n7550) );
  INV_X1 U8242 ( .A(n8181), .ZN(n7551) );
  OR2_X1 U8243 ( .A1(n12504), .A2(n12503), .ZN(n7890) );
  NAND2_X1 U8244 ( .A1(n14006), .A2(n7515), .ZN(n12813) );
  NAND2_X1 U8245 ( .A1(n12809), .A2(n7516), .ZN(n7515) );
  INV_X1 U8246 ( .A(n12810), .ZN(n7516) );
  NOR2_X1 U8247 ( .A1(n7583), .A2(n12860), .ZN(n7582) );
  OR2_X1 U8248 ( .A1(n14373), .A2(n13988), .ZN(n9394) );
  AND2_X1 U8249 ( .A1(n7946), .A2(n7944), .ZN(n7943) );
  INV_X1 U8250 ( .A(n14220), .ZN(n7944) );
  OR2_X1 U8251 ( .A1(n14403), .A2(n14032), .ZN(n7946) );
  OR2_X1 U8252 ( .A1(n14403), .A2(n14252), .ZN(n9284) );
  NAND2_X1 U8253 ( .A1(n7896), .A2(n7899), .ZN(n7430) );
  INV_X1 U8254 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9164) );
  INV_X1 U8255 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9149) );
  OR2_X1 U8256 ( .A1(n9150), .A2(n9149), .ZN(n9165) );
  NAND2_X1 U8257 ( .A1(n11513), .A2(n11512), .ZN(n7933) );
  NAND2_X1 U8258 ( .A1(n8885), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9150) );
  INV_X1 U8259 ( .A(n9135), .ZN(n8885) );
  NAND2_X1 U8260 ( .A1(n12854), .A2(n14074), .ZN(n7432) );
  OR2_X1 U8261 ( .A1(n12854), .A2(n12795), .ZN(n7936) );
  INV_X1 U8262 ( .A(n14413), .ZN(n14272) );
  AND2_X1 U8263 ( .A1(n9348), .A2(n9347), .ZN(n9353) );
  OR2_X1 U8264 ( .A1(n9096), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8978) );
  AND2_X1 U8265 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n12581), .ZN(n12659) );
  INV_X1 U8266 ( .A(n14484), .ZN(n7816) );
  XNOR2_X1 U8267 ( .A(n15146), .B(n15164), .ZN(n7630) );
  NOR2_X1 U8268 ( .A1(n14976), .A2(n14977), .ZN(n7629) );
  NOR2_X1 U8269 ( .A1(n7612), .A2(n15387), .ZN(n7611) );
  INV_X1 U8270 ( .A(n7613), .ZN(n7612) );
  AND2_X1 U8271 ( .A1(n7509), .A2(n7247), .ZN(n7505) );
  AND2_X1 U8272 ( .A1(n15262), .A2(n7510), .ZN(n7509) );
  INV_X1 U8273 ( .A(n8104), .ZN(n7510) );
  NOR2_X1 U8274 ( .A1(n15392), .A2(n15232), .ZN(n7613) );
  INV_X1 U8275 ( .A(n12626), .ZN(n12644) );
  INV_X1 U8276 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n12214) );
  INV_X1 U8277 ( .A(n7988), .ZN(n7987) );
  INV_X1 U8278 ( .A(n12211), .ZN(n8095) );
  INV_X1 U8279 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11985) );
  NOR2_X1 U8280 ( .A1(n11986), .A2(n11985), .ZN(n12011) );
  OR2_X1 U8281 ( .A1(n11977), .A2(n11976), .ZN(n11986) );
  INV_X1 U8282 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11306) );
  NOR2_X1 U8283 ( .A1(n11307), .A2(n11306), .ZN(n11592) );
  INV_X1 U8284 ( .A(n14954), .ZN(n8092) );
  NAND2_X1 U8285 ( .A1(n7504), .A2(n12649), .ZN(n15263) );
  NAND2_X1 U8286 ( .A1(n12637), .A2(n7507), .ZN(n7504) );
  INV_X1 U8287 ( .A(n7636), .ZN(n7635) );
  OAI21_X1 U8288 ( .B1(n9339), .B2(n7637), .A(n9621), .ZN(n7636) );
  INV_X1 U8289 ( .A(n9341), .ZN(n7637) );
  NAND2_X1 U8290 ( .A1(n8862), .A2(n8861), .ZN(n9340) );
  OR2_X1 U8291 ( .A1(n8860), .A2(n8859), .ZN(n8861) );
  XNOR2_X1 U8292 ( .A(n8860), .B(n8858), .ZN(n8913) );
  INV_X1 U8293 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9981) );
  INV_X1 U8294 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9984) );
  AOI21_X1 U8295 ( .B1(n8146), .B2(n8041), .A(n8040), .ZN(n8039) );
  INV_X1 U8296 ( .A(n8804), .ZN(n8040) );
  XNOR2_X1 U8297 ( .A(n8777), .B(n7622), .ZN(n9048) );
  NAND4_X1 U8298 ( .A1(n9961), .A2(n8224), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U8299 ( .A1(n9859), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7713) );
  INV_X1 U8300 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n9861) );
  NOR2_X1 U8301 ( .A1(n9877), .A2(n9876), .ZN(n9905) );
  NOR2_X1 U8302 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9932), .ZN(n9876) );
  AOI21_X1 U8303 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(n9886), .A(n9885), .ZN(
        n9898) );
  AND2_X1 U8304 ( .A1(n9900), .A2(n9899), .ZN(n9885) );
  INV_X1 U8305 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n13378) );
  INV_X1 U8306 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n13454) );
  NAND2_X1 U8307 ( .A1(n9810), .A2(n13184), .ZN(n13186) );
  NAND2_X1 U8308 ( .A1(n8000), .A2(n8001), .ZN(n13206) );
  OR2_X1 U8309 ( .A1(n8557), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8590) );
  AND2_X1 U8310 ( .A1(n8742), .A2(n8741), .ZN(n10504) );
  OR2_X1 U8311 ( .A1(n8544), .A2(n8269), .ZN(n8277) );
  AND2_X1 U8312 ( .A1(n8275), .A2(n8276), .ZN(n7745) );
  NAND2_X1 U8313 ( .A1(n8654), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8276) );
  OR2_X1 U8314 ( .A1(n8270), .A2(n11221), .ZN(n8275) );
  INV_X1 U8315 ( .A(n7727), .ZN(n7724) );
  NAND2_X1 U8316 ( .A1(n7726), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7725) );
  XNOR2_X1 U8317 ( .A(n10588), .B(n10622), .ZN(n10613) );
  INV_X1 U8318 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U8319 ( .A1(n7720), .A2(n10599), .ZN(n7719) );
  NOR2_X1 U8320 ( .A1(n10599), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7722) );
  OR2_X1 U8321 ( .A1(n7723), .A2(n8306), .ZN(n7721) );
  NAND2_X1 U8322 ( .A1(n7729), .A2(n10644), .ZN(n7728) );
  NAND2_X1 U8323 ( .A1(n10736), .A2(n10737), .ZN(n10738) );
  INV_X1 U8324 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n13448) );
  AOI21_X1 U8325 ( .B1(n7423), .B2(P3_REG1_REG_9__SCAN_IN), .A(n7218), .ZN(
        n15696) );
  AND2_X1 U8326 ( .A1(n7731), .A2(n7730), .ZN(n15716) );
  NAND2_X1 U8327 ( .A1(n12282), .A2(n12303), .ZN(n7730) );
  NOR2_X1 U8328 ( .A1(n12286), .A2(n7735), .ZN(n13495) );
  NAND2_X1 U8329 ( .A1(n7736), .A2(n12285), .ZN(n13496) );
  INV_X1 U8330 ( .A(n12286), .ZN(n7736) );
  OR2_X1 U8331 ( .A1(n13507), .A2(n13506), .ZN(n13508) );
  AND2_X1 U8332 ( .A1(n13512), .A2(n13525), .ZN(n7392) );
  NOR2_X1 U8333 ( .A1(n13520), .A2(n7221), .ZN(n13539) );
  NAND2_X1 U8334 ( .A1(n13508), .A2(n13536), .ZN(n13528) );
  NAND2_X1 U8335 ( .A1(n7565), .A2(n7564), .ZN(n7563) );
  INV_X1 U8336 ( .A(n13542), .ZN(n7564) );
  OR2_X1 U8337 ( .A1(n13539), .A2(n13540), .ZN(n7565) );
  NOR2_X1 U8338 ( .A1(n13552), .A2(n7715), .ZN(n13570) );
  NOR2_X1 U8339 ( .A1(n13541), .A2(n13903), .ZN(n7715) );
  XNOR2_X1 U8340 ( .A(n13585), .B(n7561), .ZN(n13565) );
  NOR2_X1 U8341 ( .A1(n13814), .A2(n13565), .ZN(n13586) );
  NOR2_X1 U8342 ( .A1(n7743), .A2(n13601), .ZN(n7739) );
  INV_X1 U8343 ( .A(n13573), .ZN(n7743) );
  AOI21_X1 U8344 ( .B1(n13652), .B2(n13638), .A(n13630), .ZN(n8659) );
  NAND2_X1 U8345 ( .A1(n13673), .A2(n8142), .ZN(n13660) );
  AND2_X1 U8346 ( .A1(n8645), .A2(n8644), .ZN(n13675) );
  OR2_X1 U8347 ( .A1(n13671), .A2(n13684), .ZN(n13673) );
  NAND2_X1 U8348 ( .A1(n8565), .A2(n13378), .ZN(n8612) );
  OR2_X1 U8349 ( .A1(n8612), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8626) );
  AND2_X1 U8350 ( .A1(n13755), .A2(n13703), .ZN(n13740) );
  OR2_X1 U8351 ( .A1(n13754), .A2(n13765), .ZN(n13755) );
  OR2_X1 U8352 ( .A1(n8475), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8506) );
  NAND2_X1 U8353 ( .A1(n7771), .A2(n7774), .ZN(n13819) );
  NAND2_X1 U8354 ( .A1(n12534), .A2(n7775), .ZN(n7771) );
  AOI21_X1 U8355 ( .B1(n7663), .B2(n7661), .A(n7283), .ZN(n7660) );
  INV_X1 U8356 ( .A(n8453), .ZN(n7661) );
  INV_X1 U8357 ( .A(n7663), .ZN(n7662) );
  OR2_X1 U8358 ( .A1(n8410), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8430) );
  AND4_X1 U8359 ( .A1(n8435), .A2(n8434), .A3(n8433), .A4(n8432), .ZN(n12380)
         );
  AND2_X1 U8360 ( .A1(n8409), .A2(n7677), .ZN(n7675) );
  NAND2_X1 U8361 ( .A1(n7673), .A2(n7266), .ZN(n7672) );
  AND2_X1 U8362 ( .A1(n12950), .A2(n12947), .ZN(n13061) );
  AND2_X1 U8363 ( .A1(n12943), .A2(n12944), .ZN(n13062) );
  NAND2_X1 U8364 ( .A1(n7671), .A2(n7676), .ZN(n12255) );
  NAND2_X1 U8365 ( .A1(n11923), .A2(n7677), .ZN(n7671) );
  AND2_X1 U8366 ( .A1(n11496), .A2(n8354), .ZN(n11670) );
  NAND2_X1 U8367 ( .A1(n11249), .A2(n8332), .ZN(n11494) );
  NAND2_X1 U8368 ( .A1(n7684), .A2(n8304), .ZN(n11442) );
  AND2_X1 U8369 ( .A1(n8304), .A2(n8680), .ZN(n7683) );
  OR2_X1 U8370 ( .A1(n8292), .A2(n8279), .ZN(n8283) );
  NAND2_X1 U8371 ( .A1(n13029), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8282) );
  INV_X1 U8372 ( .A(n7756), .ZN(n13639) );
  OAI21_X1 U8373 ( .B1(n13754), .B2(n8600), .A(n8606), .ZN(n13692) );
  OR2_X1 U8374 ( .A1(n13729), .A2(n13728), .ZN(n13731) );
  NAND2_X1 U8375 ( .A1(n8576), .A2(n8575), .ZN(n13870) );
  NAND2_X1 U8376 ( .A1(n7777), .A2(n7774), .ZN(n7770) );
  AND2_X1 U8377 ( .A1(n8692), .A2(n7773), .ZN(n7772) );
  NAND2_X1 U8378 ( .A1(n12550), .A2(n12549), .ZN(n7761) );
  AND3_X1 U8379 ( .A1(n8391), .A2(n8390), .A3(n8389), .ZN(n15866) );
  NAND2_X1 U8380 ( .A1(n11928), .A2(n11927), .ZN(n11926) );
  INV_X1 U8381 ( .A(n13833), .ZN(n13759) );
  INV_X1 U8382 ( .A(n15912), .ZN(n15865) );
  AND2_X1 U8383 ( .A1(n10004), .A2(n13966), .ZN(n10898) );
  INV_X1 U8384 ( .A(n10504), .ZN(n9830) );
  NAND2_X1 U8385 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n7868), .ZN(n7867) );
  NAND2_X1 U8386 ( .A1(n7846), .A2(n7844), .ZN(n13018) );
  NAND2_X1 U8387 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n7845), .ZN(n7844) );
  NAND2_X1 U8388 ( .A1(n8648), .A2(n8649), .ZN(n7846) );
  AOI21_X1 U8389 ( .B1(n7862), .B2(n7864), .A(n7351), .ZN(n7859) );
  NAND2_X1 U8390 ( .A1(n7870), .A2(n7250), .ZN(n8208) );
  NAND2_X1 U8391 ( .A1(n8441), .A2(n8011), .ZN(n8738) );
  AND2_X1 U8392 ( .A1(n8012), .A2(n8665), .ZN(n8011) );
  OAI21_X1 U8393 ( .B1(n8516), .B2(n7494), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8660) );
  INV_X1 U8394 ( .A(n8515), .ZN(n7495) );
  INV_X1 U8395 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8514) );
  AND2_X1 U8396 ( .A1(n7482), .A2(n7483), .ZN(n7481) );
  AND3_X1 U8397 ( .A1(n7485), .A2(n7484), .A3(n8163), .ZN(n7482) );
  AOI21_X1 U8398 ( .B1(n7554), .B2(n7556), .A(P2_DATAO_REG_13__SCAN_IN), .ZN(
        n7553) );
  AND2_X1 U8399 ( .A1(n10099), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8186) );
  XNOR2_X1 U8400 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8262) );
  OR2_X1 U8401 ( .A1(n9165), .A2(n9164), .ZN(n9167) );
  INV_X1 U8402 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9118) );
  OR2_X1 U8403 ( .A1(n9119), .A2(n9118), .ZN(n9135) );
  INV_X1 U8404 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8923) );
  AND2_X1 U8405 ( .A1(n7210), .A2(n13117), .ZN(n7521) );
  OR2_X1 U8406 ( .A1(n8949), .A2(n8923), .ZN(n9174) );
  AND2_X1 U8407 ( .A1(n12813), .A2(n12812), .ZN(n7389) );
  NAND2_X1 U8408 ( .A1(n8884), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9119) );
  INV_X1 U8409 ( .A(n9102), .ZN(n8884) );
  NAND2_X1 U8410 ( .A1(n7887), .A2(n12738), .ZN(n7886) );
  INV_X1 U8411 ( .A(n7890), .ZN(n7887) );
  INV_X1 U8412 ( .A(n7538), .ZN(n7536) );
  NAND2_X1 U8413 ( .A1(n11794), .A2(n11793), .ZN(n13138) );
  INV_X1 U8414 ( .A(n11875), .ZN(n11794) );
  NAND2_X1 U8415 ( .A1(n7879), .A2(n7878), .ZN(n11008) );
  INV_X1 U8416 ( .A(n11010), .ZN(n7879) );
  NAND2_X1 U8417 ( .A1(n8886), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8955) );
  INV_X1 U8418 ( .A(n9167), .ZN(n8886) );
  NAND2_X1 U8419 ( .A1(n8887), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8949) );
  INV_X1 U8420 ( .A(n8955), .ZN(n8887) );
  INV_X1 U8421 ( .A(n8061), .ZN(n8059) );
  INV_X1 U8422 ( .A(n9679), .ZN(n9675) );
  OR3_X1 U8423 ( .A1(n9679), .A2(n9678), .A3(n9677), .ZN(n9692) );
  AOI21_X1 U8424 ( .B1(n10232), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10261), .ZN(
        n10252) );
  OR2_X1 U8425 ( .A1(n15529), .A2(n15528), .ZN(n7590) );
  OR2_X1 U8426 ( .A1(n15540), .A2(n15539), .ZN(n7588) );
  NOR2_X1 U8427 ( .A1(n11109), .A2(n7601), .ZN(n11113) );
  AND2_X1 U8428 ( .A1(n11110), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7601) );
  NAND2_X1 U8429 ( .A1(n11113), .A2(n11112), .ZN(n11528) );
  NAND2_X1 U8430 ( .A1(n15579), .A2(n15580), .ZN(n15578) );
  NOR2_X1 U8431 ( .A1(n14083), .A2(n7598), .ZN(n14098) );
  AND2_X1 U8432 ( .A1(n14084), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7598) );
  OR2_X1 U8433 ( .A1(n15564), .A2(n15563), .ZN(n7597) );
  NAND2_X1 U8434 ( .A1(n7597), .A2(n7596), .ZN(n7595) );
  NAND2_X1 U8435 ( .A1(n15567), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7596) );
  AND2_X1 U8436 ( .A1(n7595), .A2(n14122), .ZN(n14135) );
  NOR2_X1 U8437 ( .A1(n14191), .A2(n7580), .ZN(n14158) );
  INV_X1 U8438 ( .A(n7582), .ZN(n7580) );
  OR2_X1 U8439 ( .A1(n14191), .A2(n7581), .ZN(n14157) );
  NAND2_X1 U8440 ( .A1(n14159), .A2(n7582), .ZN(n7581) );
  OAI21_X1 U8441 ( .B1(n9395), .B2(n7925), .A(n7922), .ZN(n7921) );
  NAND2_X1 U8442 ( .A1(n7925), .A2(n7923), .ZN(n7922) );
  NAND2_X1 U8443 ( .A1(n9712), .A2(n7927), .ZN(n7923) );
  NAND2_X1 U8444 ( .A1(n7928), .A2(n9395), .ZN(n7924) );
  NOR2_X1 U8445 ( .A1(n9712), .A2(n7438), .ZN(n7437) );
  INV_X1 U8446 ( .A(n7440), .ZN(n7438) );
  NOR2_X1 U8447 ( .A1(n7440), .A2(n7207), .ZN(n7435) );
  NAND2_X1 U8448 ( .A1(n14377), .A2(n14190), .ZN(n7442) );
  NOR2_X1 U8449 ( .A1(n14167), .A2(n7441), .ZN(n7440) );
  INV_X1 U8450 ( .A(n7442), .ZN(n7441) );
  NAND2_X1 U8451 ( .A1(n7929), .A2(n7236), .ZN(n7369) );
  NAND2_X1 U8452 ( .A1(n14235), .A2(n7946), .ZN(n14219) );
  NAND2_X1 U8453 ( .A1(n14242), .A2(n14241), .ZN(n14240) );
  NAND2_X1 U8454 ( .A1(n8889), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9243) );
  INV_X1 U8455 ( .A(n9217), .ZN(n8889) );
  NAND2_X1 U8456 ( .A1(n14325), .A2(n14324), .ZN(n14323) );
  AND2_X1 U8457 ( .A1(n7938), .A2(n7246), .ZN(n14319) );
  NAND2_X1 U8458 ( .A1(n7444), .A2(n7228), .ZN(n7443) );
  INV_X1 U8459 ( .A(n7446), .ZN(n7444) );
  OR2_X1 U8460 ( .A1(n12134), .A2(n9379), .ZN(n9380) );
  OR2_X1 U8461 ( .A1(n12059), .A2(n12134), .ZN(n12057) );
  NAND2_X1 U8462 ( .A1(n13145), .A2(n11846), .ZN(n12059) );
  NAND2_X1 U8463 ( .A1(n7933), .A2(n7932), .ZN(n11840) );
  AND2_X1 U8464 ( .A1(n11841), .A2(n7244), .ZN(n7932) );
  AND2_X1 U8465 ( .A1(n7933), .A2(n7244), .ZN(n11842) );
  NAND2_X1 U8466 ( .A1(n7584), .A2(n15904), .ZN(n11509) );
  OR2_X1 U8467 ( .A1(n9100), .A2(n10963), .ZN(n9102) );
  INV_X1 U8468 ( .A(n11463), .ZN(n7366) );
  NAND2_X1 U8469 ( .A1(n9041), .A2(n9040), .ZN(n11474) );
  NAND2_X1 U8470 ( .A1(n10536), .A2(n10537), .ZN(n10535) );
  AND2_X1 U8471 ( .A1(n9396), .A2(n9647), .ZN(n14298) );
  INV_X1 U8472 ( .A(n10495), .ZN(n7576) );
  XNOR2_X1 U8473 ( .A(n14081), .B(n9019), .ZN(n10447) );
  INV_X1 U8474 ( .A(n10447), .ZN(n10450) );
  NAND2_X1 U8475 ( .A1(n7892), .A2(n13125), .ZN(n10487) );
  INV_X1 U8476 ( .A(n9362), .ZN(n7892) );
  OR2_X1 U8477 ( .A1(n9437), .A2(n9401), .ZN(n14322) );
  NAND2_X1 U8478 ( .A1(n14204), .A2(n9312), .ZN(n14196) );
  NAND2_X1 U8479 ( .A1(n9302), .A2(n9301), .ZN(n14392) );
  NAND2_X1 U8480 ( .A1(n9190), .A2(n9189), .ZN(n14428) );
  NAND2_X1 U8481 ( .A1(n10163), .A2(n11868), .ZN(n15821) );
  NOR2_X1 U8482 ( .A1(n9012), .A2(n8180), .ZN(n7931) );
  INV_X1 U8483 ( .A(n15821), .ZN(n14445) );
  INV_X1 U8484 ( .A(n9444), .ZN(n14449) );
  INV_X1 U8485 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U8486 ( .A1(n9420), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9422) );
  INV_X1 U8487 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9421) );
  INV_X1 U8488 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9424) );
  XNOR2_X1 U8489 ( .A(n9359), .B(n9358), .ZN(n9361) );
  NAND2_X1 U8490 ( .A1(n9419), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9359) );
  INV_X1 U8491 ( .A(n9253), .ZN(n9254) );
  XNOR2_X1 U8492 ( .A(n9132), .B(P2_IR_REG_11__SCAN_IN), .ZN(n12100) );
  OR2_X1 U8493 ( .A1(n9053), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9068) );
  OR2_X1 U8494 ( .A1(n9037), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9053) );
  NOR2_X1 U8495 ( .A1(n9029), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9032) );
  OR2_X1 U8496 ( .A1(n9013), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U8497 ( .A1(n7825), .A2(n7824), .ZN(n7823) );
  INV_X1 U8498 ( .A(n12424), .ZN(n7824) );
  INV_X1 U8499 ( .A(n12423), .ZN(n7825) );
  INV_X1 U8500 ( .A(n12643), .ZN(n10748) );
  AND2_X1 U8501 ( .A1(n7786), .A2(n7785), .ZN(n10910) );
  NAND2_X1 U8502 ( .A1(n14563), .A2(n7377), .ZN(n7786) );
  NAND2_X1 U8503 ( .A1(n11286), .A2(n14769), .ZN(n7785) );
  AND2_X1 U8504 ( .A1(n12600), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n12612) );
  NAND2_X1 U8505 ( .A1(n11291), .A2(n7235), .ZN(n7833) );
  AND2_X1 U8506 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n10812) );
  NOR2_X1 U8507 ( .A1(n10995), .A2(n10997), .ZN(n10999) );
  XNOR2_X1 U8508 ( .A(n10909), .B(n10910), .ZN(n12778) );
  INV_X1 U8509 ( .A(n12705), .ZN(n14923) );
  AND4_X1 U8510 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11817) );
  NAND4_X1 U8511 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n15055) );
  OR2_X1 U8512 ( .A1(n12704), .A2(n15754), .ZN(n10313) );
  NAND2_X1 U8513 ( .A1(n14924), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n10310) );
  OR2_X1 U8514 ( .A1(n10397), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n10565) );
  OR2_X1 U8515 ( .A1(n11160), .A2(n11159), .ZN(n11157) );
  AND2_X1 U8516 ( .A1(n12674), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12687) );
  NAND2_X1 U8517 ( .A1(n15246), .A2(n7613), .ZN(n15208) );
  NAND2_X1 U8518 ( .A1(n15246), .A2(n15398), .ZN(n15227) );
  NAND2_X1 U8519 ( .A1(n12625), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12626) );
  INV_X1 U8520 ( .A(n7966), .ZN(n7965) );
  OAI21_X1 U8521 ( .B1(n7970), .B2(n7968), .A(n12725), .ZN(n7966) );
  NAND2_X1 U8522 ( .A1(n7969), .A2(n7967), .ZN(n15308) );
  NAND2_X1 U8523 ( .A1(n7616), .A2(n7615), .ZN(n15356) );
  INV_X1 U8524 ( .A(n15355), .ZN(n7616) );
  NAND2_X1 U8525 ( .A1(n7614), .A2(n7975), .ZN(n15327) );
  INV_X1 U8526 ( .A(n15356), .ZN(n7614) );
  NOR2_X1 U8527 ( .A1(n12215), .A2(n12214), .ZN(n12337) );
  AND2_X1 U8528 ( .A1(n12337), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n12600) );
  NAND2_X1 U8529 ( .A1(n12590), .A2(n8094), .ZN(n15348) );
  NAND2_X1 U8530 ( .A1(n12590), .A2(n12589), .ZN(n15341) );
  NAND2_X1 U8531 ( .A1(n7618), .A2(n7617), .ZN(n15355) );
  NAND2_X1 U8532 ( .A1(n12333), .A2(n14968), .ZN(n12590) );
  INV_X1 U8533 ( .A(n7618), .ZN(n12335) );
  INV_X1 U8534 ( .A(n7957), .ZN(n7956) );
  NAND2_X1 U8535 ( .A1(n15933), .A2(n15934), .ZN(n15931) );
  NAND2_X1 U8536 ( .A1(n7607), .A2(n7606), .ZN(n12021) );
  INV_X1 U8537 ( .A(n15931), .ZN(n7607) );
  NAND2_X1 U8538 ( .A1(n11603), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11750) );
  INV_X1 U8539 ( .A(n11964), .ZN(n15930) );
  NAND2_X1 U8540 ( .A1(n15930), .A2(n11969), .ZN(n15929) );
  NOR2_X1 U8541 ( .A1(n11721), .A2(n14815), .ZN(n11760) );
  NAND2_X1 U8542 ( .A1(n11717), .A2(n11586), .ZN(n11764) );
  NAND2_X1 U8543 ( .A1(n11599), .A2(n11662), .ZN(n11720) );
  INV_X1 U8544 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n11278) );
  OR2_X1 U8545 ( .A1(n11279), .A2(n11278), .ZN(n11307) );
  NAND2_X1 U8546 ( .A1(n11580), .A2(n11579), .ZN(n11652) );
  NAND2_X1 U8547 ( .A1(n7959), .A2(n7261), .ZN(n11578) );
  AOI21_X1 U8548 ( .B1(n11564), .B2(n11567), .A(n7964), .ZN(n7963) );
  AOI21_X1 U8549 ( .B1(n14953), .B2(n7500), .A(n7286), .ZN(n7499) );
  INV_X1 U8550 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10831) );
  NOR2_X1 U8551 ( .A1(n10832), .A2(n10831), .ZN(n11037) );
  NAND2_X1 U8552 ( .A1(n11131), .A2(n11130), .ZN(n11132) );
  AND3_X1 U8553 ( .A1(n10340), .A2(n10339), .A3(n10338), .ZN(n10825) );
  NAND2_X1 U8554 ( .A1(n10065), .A2(n7378), .ZN(n10340) );
  NAND2_X1 U8555 ( .A1(n10328), .A2(n10329), .ZN(n11321) );
  NAND2_X1 U8556 ( .A1(n7976), .A2(n11581), .ZN(n11719) );
  AND2_X1 U8557 ( .A1(n11263), .A2(n10362), .ZN(n15981) );
  INV_X1 U8558 ( .A(n15973), .ZN(n15985) );
  AND2_X1 U8559 ( .A1(n10131), .A2(n10113), .ZN(n7410) );
  AND2_X1 U8560 ( .A1(n9626), .A2(n8028), .ZN(n8025) );
  NAND2_X1 U8561 ( .A1(n8027), .A2(n9628), .ZN(n8026) );
  INV_X1 U8562 ( .A(n9626), .ZN(n8027) );
  INV_X1 U8563 ( .A(n9628), .ZN(n8028) );
  XNOR2_X1 U8564 ( .A(n9340), .B(n9339), .ZN(n12698) );
  INV_X1 U8565 ( .A(n11700), .ZN(n7498) );
  XNOR2_X1 U8566 ( .A(n8914), .B(SI_27_), .ZN(n12586) );
  INV_X1 U8567 ( .A(n8913), .ZN(n8914) );
  INV_X1 U8568 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U8569 ( .A1(n7642), .A2(n8854), .ZN(n9314) );
  OR2_X1 U8570 ( .A1(n9300), .A2(n9299), .ZN(n7642) );
  NAND2_X1 U8571 ( .A1(n7652), .A2(n8841), .ZN(n9268) );
  NAND2_X1 U8572 ( .A1(n8838), .A2(n8837), .ZN(n9238) );
  XNOR2_X1 U8573 ( .A(n9210), .B(n9209), .ZN(n12595) );
  AOI21_X1 U8574 ( .B1(n8807), .B2(n8033), .A(n7627), .ZN(n7624) );
  NAND2_X1 U8575 ( .A1(n8029), .A2(n8033), .ZN(n8941) );
  OR2_X1 U8576 ( .A1(n8807), .A2(n8035), .ZN(n8029) );
  NAND2_X1 U8577 ( .A1(n8807), .A2(n8806), .ZN(n8962) );
  NAND2_X1 U8578 ( .A1(n8042), .A2(n8799), .ZN(n9142) );
  NAND2_X1 U8579 ( .A1(n8795), .A2(n8043), .ZN(n8042) );
  NAND2_X1 U8580 ( .A1(n7527), .A2(n8787), .ZN(n9094) );
  NAND2_X1 U8581 ( .A1(n9082), .A2(n8785), .ZN(n7527) );
  XNOR2_X1 U8582 ( .A(n9036), .B(n7621), .ZN(n10806) );
  INV_X1 U8583 ( .A(n9048), .ZN(n7621) );
  INV_X1 U8584 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10067) );
  NAND2_X1 U8585 ( .A1(n7692), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7691) );
  AND2_X1 U8586 ( .A1(n15620), .A2(n15622), .ZN(n9936) );
  OAI21_X1 U8587 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n15110), .A(n9879), .ZN(
        n9902) );
  AOI21_X1 U8588 ( .B1(n10702), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n9884), .ZN(
        n9900) );
  AND2_X1 U8589 ( .A1(n9942), .A2(n9941), .ZN(n9884) );
  NAND2_X1 U8590 ( .A1(n7699), .A2(n7698), .ZN(n9949) );
  NAND2_X1 U8591 ( .A1(n7700), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7699) );
  AND2_X1 U8592 ( .A1(n15663), .A2(n7239), .ZN(n7707) );
  AND2_X1 U8593 ( .A1(n7709), .A2(n7706), .ZN(n7705) );
  OR2_X1 U8594 ( .A1(n15660), .A2(n7710), .ZN(n7706) );
  AND4_X1 U8595 ( .A1(n8362), .A2(n8361), .A3(n8360), .A4(n8359), .ZN(n11935)
         );
  NAND2_X1 U8596 ( .A1(n7475), .A2(n8003), .ZN(n11933) );
  NAND2_X1 U8597 ( .A1(n12482), .A2(n12481), .ZN(n12480) );
  NAND2_X1 U8598 ( .A1(n8001), .A2(n13205), .ZN(n13162) );
  AND2_X1 U8599 ( .A1(n8408), .A2(n8407), .ZN(n12248) );
  NAND2_X1 U8600 ( .A1(n12244), .A2(n9762), .ZN(n12245) );
  OR2_X1 U8601 ( .A1(n11084), .A2(n11085), .ZN(n9751) );
  NAND2_X1 U8602 ( .A1(n7468), .A2(n7467), .ZN(n12083) );
  AOI21_X1 U8603 ( .B1(n7473), .B2(n7471), .A(n7212), .ZN(n7467) );
  NAND2_X1 U8604 ( .A1(n7472), .A2(n7473), .ZN(n7468) );
  AOI21_X1 U8605 ( .B1(n12244), .B2(n7209), .A(n7995), .ZN(n12411) );
  NAND2_X1 U8606 ( .A1(n8487), .A2(n8486), .ZN(n13836) );
  AND4_X1 U8607 ( .A1(n8325), .A2(n8324), .A3(n8323), .A4(n8322), .ZN(n11497)
         );
  NAND2_X1 U8608 ( .A1(n7486), .A2(n7490), .ZN(n12541) );
  NAND2_X1 U8609 ( .A1(n12482), .A2(n7491), .ZN(n7486) );
  NAND2_X1 U8610 ( .A1(n13169), .A2(n13168), .ZN(n9792) );
  OAI21_X1 U8611 ( .B1(n7994), .B2(n7992), .A(n7990), .ZN(n12459) );
  OAI21_X1 U8612 ( .B1(n7995), .B2(n7991), .A(n7993), .ZN(n7990) );
  NAND2_X1 U8613 ( .A1(n7209), .A2(n7993), .ZN(n7992) );
  AND3_X1 U8614 ( .A1(n8595), .A2(n8594), .A3(n8593), .ZN(n13763) );
  INV_X1 U8615 ( .A(n13224), .ZN(n9798) );
  NAND2_X1 U8616 ( .A1(n12245), .A2(n9765), .ZN(n12318) );
  XNOR2_X1 U8617 ( .A(n9749), .B(n9748), .ZN(n7478) );
  AOI21_X1 U8618 ( .B1(n12482), .B2(n7489), .A(n7487), .ZN(n12570) );
  OAI21_X1 U8619 ( .B1(n7490), .B2(n7488), .A(n7248), .ZN(n7487) );
  AND2_X1 U8620 ( .A1(n7491), .A2(n9787), .ZN(n7489) );
  NAND2_X1 U8621 ( .A1(n11426), .A2(n9757), .ZN(n11853) );
  OR2_X1 U8622 ( .A1(n9843), .A2(n9839), .ZN(n13247) );
  NAND2_X1 U8623 ( .A1(n9837), .A2(n9836), .ZN(n13250) );
  INV_X1 U8624 ( .A(n13222), .ZN(n13241) );
  INV_X1 U8625 ( .A(n12899), .ZN(n13092) );
  INV_X1 U8626 ( .A(n13663), .ZN(n13257) );
  INV_X1 U8627 ( .A(n13675), .ZN(n13651) );
  NAND2_X1 U8628 ( .A1(n8632), .A2(n8631), .ZN(n13691) );
  INV_X1 U8629 ( .A(n13710), .ZN(n13743) );
  INV_X1 U8630 ( .A(n13832), .ZN(n13262) );
  OR2_X1 U8631 ( .A1(n10004), .A2(n13964), .ZN(n13265) );
  INV_X1 U8632 ( .A(n11935), .ZN(n13482) );
  INV_X1 U8633 ( .A(n11497), .ZN(n13484) );
  OR2_X1 U8634 ( .A1(n8528), .A2(n8307), .ZN(n8308) );
  OR2_X1 U8635 ( .A1(n8544), .A2(n8290), .ZN(n8296) );
  NAND2_X1 U8636 ( .A1(n13029), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8293) );
  AOI22_X1 U8637 ( .A1(n10579), .A2(n15679), .B1(n10578), .B2(n10577), .ZN(
        n10669) );
  OR2_X1 U8638 ( .A1(n7725), .A2(n7724), .ZN(n10616) );
  XNOR2_X1 U8639 ( .A(n10735), .B(n10727), .ZN(n10639) );
  NAND2_X1 U8640 ( .A1(n10639), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n10736) );
  OAI22_X1 U8641 ( .A1(n10717), .A2(n10718), .B1(n10631), .B2(n10716), .ZN(
        n10729) );
  NOR2_X1 U8642 ( .A1(n10731), .A2(n7744), .ZN(n10986) );
  INV_X1 U8643 ( .A(n10647), .ZN(n7744) );
  OAI22_X1 U8644 ( .A1(n10980), .A2(n10979), .B1(n10978), .B2(n10988), .ZN(
        n11543) );
  INV_X1 U8645 ( .A(n7731), .ZN(n12281) );
  NOR2_X1 U8646 ( .A1(n7734), .A2(n12286), .ZN(n12289) );
  NAND2_X1 U8647 ( .A1(n13489), .A2(n12309), .ZN(n13510) );
  INV_X1 U8648 ( .A(n13598), .ZN(n7421) );
  AOI22_X1 U8649 ( .A1(n13022), .A2(n13028), .B1(SI_30_), .B2(n13021), .ZN(
        n15995) );
  AND2_X1 U8650 ( .A1(n7755), .A2(n13009), .ZN(n13044) );
  NAND2_X1 U8651 ( .A1(n13637), .A2(n13636), .ZN(n13844) );
  NAND2_X1 U8652 ( .A1(n8625), .A2(n8624), .ZN(n13683) );
  AND2_X1 U8653 ( .A1(n8556), .A2(n8555), .ZN(n13879) );
  NAND2_X1 U8654 ( .A1(n13826), .A2(n8495), .ZN(n13807) );
  NAND2_X1 U8655 ( .A1(n12534), .A2(n13070), .ZN(n13824) );
  NAND2_X1 U8656 ( .A1(n8474), .A2(n8473), .ZN(n13254) );
  INV_X1 U8657 ( .A(n12324), .ZN(n15913) );
  INV_X1 U8658 ( .A(n12248), .ZN(n15885) );
  NAND2_X1 U8659 ( .A1(n11923), .A2(n12931), .ZN(n12041) );
  OAI21_X1 U8660 ( .B1(n11502), .B2(n11669), .A(n7767), .ZN(n11828) );
  NAND2_X1 U8661 ( .A1(n11667), .A2(n13054), .ZN(n11666) );
  NAND2_X1 U8662 ( .A1(n11502), .A2(n12919), .ZN(n11667) );
  NAND2_X1 U8663 ( .A1(n10896), .A2(n11680), .ZN(n15806) );
  INV_X1 U8664 ( .A(n15804), .ZN(n13802) );
  INV_X1 U8665 ( .A(n13638), .ZN(n13916) );
  AND3_X1 U8666 ( .A1(n8352), .A2(n8351), .A3(n8350), .ZN(n11811) );
  INV_X1 U8667 ( .A(n13905), .ZN(n16005) );
  NAND2_X1 U8668 ( .A1(n15997), .A2(n15865), .ZN(n13905) );
  NOR2_X1 U8669 ( .A1(n13916), .A2(n13960), .ZN(n7668) );
  INV_X1 U8670 ( .A(n8699), .ZN(n13921) );
  NAND2_X1 U8671 ( .A1(n8564), .A2(n8563), .ZN(n13933) );
  AND3_X1 U8672 ( .A1(n8255), .A2(n8254), .A3(n8253), .ZN(n12891) );
  INV_X1 U8673 ( .A(n11255), .ZN(n11436) );
  OR2_X1 U8674 ( .A1(n8499), .A2(n10050), .ZN(n8302) );
  INV_X1 U8675 ( .A(n13966), .ZN(n13964) );
  AND2_X1 U8676 ( .A1(n9830), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13966) );
  XNOR2_X1 U8677 ( .A(n7866), .B(n7865), .ZN(n13974) );
  INV_X1 U8678 ( .A(n13025), .ZN(n7865) );
  NAND2_X1 U8679 ( .A1(n7869), .A2(n7867), .ZN(n7866) );
  AND2_X1 U8680 ( .A1(n7686), .A2(n8169), .ZN(n7685) );
  XNOR2_X1 U8681 ( .A(n13023), .B(n13024), .ZN(n13156) );
  INV_X1 U8682 ( .A(SI_27_), .ZN(n13385) );
  NAND2_X1 U8683 ( .A1(n7861), .A2(n8214), .ZN(n8635) );
  NAND2_X1 U8684 ( .A1(n8715), .A2(n8714), .ZN(n12873) );
  OR2_X1 U8685 ( .A1(n8740), .A2(n8708), .ZN(n8709) );
  INV_X1 U8686 ( .A(SI_23_), .ZN(n13390) );
  INV_X1 U8687 ( .A(n8747), .ZN(n12898) );
  AND2_X1 U8688 ( .A1(n7870), .A2(n7222), .ZN(n8587) );
  INV_X1 U8689 ( .A(SI_20_), .ZN(n13381) );
  XNOR2_X1 U8690 ( .A(n8663), .B(n8662), .ZN(n11146) );
  INV_X1 U8691 ( .A(SI_19_), .ZN(n13403) );
  NAND2_X1 U8692 ( .A1(n8540), .A2(n8661), .ZN(n13610) );
  OAI21_X1 U8693 ( .B1(n8201), .B2(n7547), .A(n7544), .ZN(n8512) );
  INV_X1 U8694 ( .A(SI_18_), .ZN(n13291) );
  INV_X1 U8695 ( .A(SI_17_), .ZN(n13405) );
  NAND2_X1 U8696 ( .A1(n7873), .A2(n8202), .ZN(n8498) );
  NAND2_X1 U8697 ( .A1(n8485), .A2(n8483), .ZN(n7873) );
  INV_X1 U8698 ( .A(SI_15_), .ZN(n13412) );
  INV_X1 U8699 ( .A(SI_14_), .ZN(n13272) );
  INV_X1 U8700 ( .A(SI_13_), .ZN(n13299) );
  INV_X1 U8701 ( .A(SI_12_), .ZN(n13414) );
  NAND2_X1 U8702 ( .A1(n7850), .A2(n7849), .ZN(n8424) );
  NAND2_X1 U8703 ( .A1(n8406), .A2(n8405), .ZN(n7851) );
  INV_X1 U8704 ( .A(n10733), .ZN(n10988) );
  NAND2_X1 U8705 ( .A1(n7549), .A2(n8181), .ZN(n8327) );
  INV_X1 U8706 ( .A(n10622), .ZN(n10599) );
  NAND2_X1 U8707 ( .A1(n11292), .A2(n9629), .ZN(n7449) );
  XNOR2_X1 U8708 ( .A(n12816), .B(n12814), .ZN(n13996) );
  NAND2_X1 U8709 ( .A1(n11083), .A2(n10028), .ZN(n10036) );
  AOI21_X1 U8710 ( .B1(n7876), .B2(n7877), .A(n7348), .ZN(n7874) );
  INV_X1 U8711 ( .A(n7876), .ZN(n7875) );
  INV_X1 U8712 ( .A(n10958), .ZN(n7877) );
  NAND2_X1 U8713 ( .A1(n11008), .A2(n10958), .ZN(n11100) );
  AND2_X1 U8714 ( .A1(n7885), .A2(n7213), .ZN(n14008) );
  INV_X1 U8715 ( .A(n14015), .ZN(n12826) );
  NAND2_X1 U8716 ( .A1(n9186), .A2(n9185), .ZN(n14433) );
  NAND2_X1 U8717 ( .A1(n9289), .A2(n9288), .ZN(n14396) );
  NAND2_X1 U8718 ( .A1(n7886), .A2(n7885), .ZN(n12808) );
  XNOR2_X1 U8719 ( .A(n14424), .B(n12116), .ZN(n12500) );
  OR2_X1 U8720 ( .A1(n11796), .A2(n7238), .ZN(n7517) );
  NAND2_X1 U8721 ( .A1(n11793), .A2(n7519), .ZN(n7518) );
  INV_X1 U8722 ( .A(n7238), .ZN(n7519) );
  INV_X1 U8723 ( .A(n14252), .ZN(n14032) );
  OR2_X1 U8724 ( .A1(n10034), .A2(n10013), .ZN(n14002) );
  AND2_X1 U8725 ( .A1(n10881), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14046) );
  INV_X1 U8726 ( .A(n12450), .ZN(n12451) );
  INV_X1 U8727 ( .A(n7883), .ZN(n14055) );
  NAND2_X1 U8728 ( .A1(n10012), .A2(n14308), .ZN(n14035) );
  NAND2_X1 U8729 ( .A1(n9267), .A2(n9266), .ZN(n14065) );
  NAND2_X1 U8730 ( .A1(n9042), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U8731 ( .A1(n9004), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8994) );
  NOR2_X1 U8732 ( .A1(n10373), .A2(n10372), .ZN(n10371) );
  AOI21_X1 U8733 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n10377), .A(n10371), .ZN(
        n10231) );
  NOR2_X1 U8734 ( .A1(n10231), .A2(n10230), .ZN(n10861) );
  INV_X1 U8735 ( .A(n7590), .ZN(n15527) );
  AND2_X1 U8736 ( .A1(n7590), .A2(n7589), .ZN(n15540) );
  NAND2_X1 U8737 ( .A1(n15535), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7589) );
  INV_X1 U8738 ( .A(n7588), .ZN(n15538) );
  AND2_X1 U8739 ( .A1(n7588), .A2(n7587), .ZN(n15551) );
  NAND2_X1 U8740 ( .A1(n15546), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7587) );
  NOR2_X1 U8741 ( .A1(n10873), .A2(n10872), .ZN(n11109) );
  NOR2_X1 U8742 ( .A1(n15549), .A2(n7602), .ZN(n10873) );
  AND2_X1 U8743 ( .A1(n15557), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7602) );
  NOR2_X1 U8744 ( .A1(n11533), .A2(n11532), .ZN(n12099) );
  NOR2_X1 U8745 ( .A1(n15587), .A2(n7600), .ZN(n11533) );
  AND2_X1 U8746 ( .A1(n15597), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7600) );
  NOR2_X1 U8747 ( .A1(n12362), .A2(n7343), .ZN(n12363) );
  NOR2_X1 U8748 ( .A1(n12363), .A2(n12364), .ZN(n14083) );
  XNOR2_X1 U8749 ( .A(n14098), .B(n14097), .ZN(n14086) );
  NAND2_X1 U8750 ( .A1(n14116), .A2(n7350), .ZN(n15570) );
  NOR2_X1 U8751 ( .A1(n14135), .A2(n7594), .ZN(n14128) );
  NOR2_X1 U8752 ( .A1(n7595), .A2(n14122), .ZN(n7594) );
  OR2_X1 U8753 ( .A1(n10239), .A2(n10238), .ZN(n15588) );
  INV_X1 U8754 ( .A(n14145), .ZN(n7391) );
  NAND2_X1 U8755 ( .A1(n9632), .A2(n9631), .ZN(n14365) );
  INV_X1 U8756 ( .A(n14369), .ZN(n14159) );
  AND2_X1 U8757 ( .A1(n8895), .A2(n8894), .ZN(n12862) );
  AND2_X1 U8758 ( .A1(n14185), .A2(n7904), .ZN(n7903) );
  NAND2_X1 U8759 ( .A1(n7205), .A2(n7906), .ZN(n7904) );
  NAND2_X1 U8760 ( .A1(n7902), .A2(n7205), .ZN(n14186) );
  OR2_X1 U8761 ( .A1(n14206), .A2(n7906), .ZN(n7902) );
  NAND2_X1 U8762 ( .A1(n7407), .A2(n7406), .ZN(n7405) );
  XNOR2_X1 U8763 ( .A(n14189), .B(n14195), .ZN(n7408) );
  NAND2_X1 U8764 ( .A1(n14221), .A2(n14353), .ZN(n7406) );
  AND2_X1 U8765 ( .A1(n9318), .A2(n9305), .ZN(n14210) );
  AND2_X1 U8766 ( .A1(n14239), .A2(n14238), .ZN(n14405) );
  NAND2_X1 U8767 ( .A1(n7429), .A2(n7896), .ZN(n14259) );
  NAND2_X1 U8768 ( .A1(n14295), .A2(n7898), .ZN(n7429) );
  NAND2_X1 U8769 ( .A1(n7897), .A2(n7901), .ZN(n14267) );
  NAND2_X1 U8770 ( .A1(n14295), .A2(n7227), .ZN(n7897) );
  NAND2_X1 U8771 ( .A1(n7948), .A2(n7950), .ZN(n14263) );
  OR2_X1 U8772 ( .A1(n14299), .A2(n7951), .ZN(n7948) );
  NAND2_X1 U8773 ( .A1(n14295), .A2(n9225), .ZN(n14283) );
  AND2_X1 U8774 ( .A1(n7953), .A2(n7223), .ZN(n14279) );
  NAND2_X1 U8775 ( .A1(n9384), .A2(n8143), .ZN(n14352) );
  NAND2_X1 U8776 ( .A1(n11950), .A2(n7447), .ZN(n12395) );
  NOR2_X1 U8777 ( .A1(n7914), .A2(n7915), .ZN(n12049) );
  INV_X1 U8778 ( .A(n7918), .ZN(n7914) );
  AOI21_X1 U8779 ( .B1(n11507), .B2(n11508), .A(n9141), .ZN(n11839) );
  NAND2_X1 U8780 ( .A1(n7345), .A2(n7433), .ZN(n11375) );
  NAND2_X1 U8781 ( .A1(n7893), .A2(n9080), .ZN(n11203) );
  NAND2_X1 U8782 ( .A1(n14311), .A2(n11174), .ZN(n14231) );
  INV_X1 U8783 ( .A(n14349), .ZN(n14271) );
  INV_X1 U8784 ( .A(n7425), .ZN(n7424) );
  OAI21_X1 U8785 ( .B1(n9441), .B2(P2_D_REG_1__SCAN_IN), .A(n9438), .ZN(n15519) );
  AND2_X1 U8786 ( .A1(n10224), .A2(n9436), .ZN(n15526) );
  OAI21_X1 U8787 ( .B1(n9441), .B2(P2_D_REG_0__SCAN_IN), .A(n9440), .ZN(n15525) );
  XNOR2_X1 U8788 ( .A(n9429), .B(n9428), .ZN(n12391) );
  NAND2_X1 U8789 ( .A1(n9427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U8790 ( .A1(n9427), .A2(n9423), .ZN(n12161) );
  OR2_X1 U8791 ( .A1(n9422), .A2(n9421), .ZN(n9423) );
  XNOR2_X1 U8792 ( .A(n9425), .B(n9424), .ZN(n12158) );
  INV_X1 U8793 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11863) );
  INV_X1 U8794 ( .A(n9720), .ZN(n11862) );
  INV_X1 U8795 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11869) );
  INV_X1 U8796 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11864) );
  INV_X1 U8797 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11773) );
  INV_X1 U8798 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n11407) );
  INV_X1 U8799 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11226) );
  INV_X1 U8800 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11126) );
  INV_X1 U8801 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11018) );
  INV_X1 U8802 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10610) );
  INV_X1 U8803 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10424) );
  INV_X1 U8804 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10099) );
  INV_X1 U8805 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10087) );
  AND2_X1 U8806 ( .A1(n9013), .A2(n7593), .ZN(n7592) );
  NAND2_X1 U8807 ( .A1(n8985), .A2(n8875), .ZN(n7593) );
  XNOR2_X1 U8809 ( .A(n9990), .B(n9989), .ZN(n10293) );
  INV_X1 U8810 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9989) );
  OAI21_X1 U8811 ( .B1(n9988), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9990) );
  AOI21_X1 U8812 ( .B1(n11291), .B2(n11290), .A(n11289), .ZN(n11417) );
  NAND2_X1 U8813 ( .A1(n7826), .A2(n7823), .ZN(n12427) );
  OR2_X1 U8814 ( .A1(n12426), .A2(n12425), .ZN(n7826) );
  NAND2_X1 U8815 ( .A1(n12274), .A2(n7820), .ZN(n7814) );
  NAND2_X1 U8816 ( .A1(n14558), .A2(n7809), .ZN(n7808) );
  NAND2_X1 U8817 ( .A1(n7810), .A2(n7813), .ZN(n7809) );
  AND2_X1 U8818 ( .A1(n14596), .A2(n14597), .ZN(n14558) );
  NAND2_X1 U8819 ( .A1(n7793), .A2(n14632), .ZN(n7792) );
  OAI22_X1 U8820 ( .A1(n7789), .A2(n7788), .B1(n7798), .B2(n7793), .ZN(n7787)
         );
  INV_X1 U8821 ( .A(n7793), .ZN(n7788) );
  NOR2_X1 U8822 ( .A1(n7798), .A2(n7794), .ZN(n7789) );
  AND4_X1 U8823 ( .A1(n11042), .A2(n11041), .A3(n11040), .A4(n11039), .ZN(
        n11617) );
  NAND2_X1 U8824 ( .A1(n7833), .A2(n7831), .ZN(n11303) );
  INV_X1 U8825 ( .A(n7834), .ZN(n7831) );
  INV_X1 U8826 ( .A(n10769), .ZN(n10765) );
  OR2_X1 U8827 ( .A1(n12229), .A2(n12230), .ZN(n7799) );
  OR2_X1 U8828 ( .A1(n7832), .A2(n7830), .ZN(n7829) );
  INV_X1 U8829 ( .A(n7837), .ZN(n7830) );
  NAND2_X1 U8830 ( .A1(n14693), .A2(n14532), .ZN(n14690) );
  NOR2_X1 U8831 ( .A1(n12274), .A2(n7234), .ZN(n12426) );
  NAND2_X1 U8832 ( .A1(n14690), .A2(n14540), .ZN(n14703) );
  OAI21_X1 U8833 ( .B1(n14693), .B2(n7813), .A(n7810), .ZN(n14700) );
  OR2_X1 U8834 ( .A1(n14665), .A2(n15195), .ZN(n14747) );
  AOI21_X2 U8835 ( .B1(n11027), .B2(n11026), .A(n11025), .ZN(n11291) );
  OR2_X1 U8836 ( .A1(n14665), .A2(n15345), .ZN(n14743) );
  AND2_X1 U8837 ( .A1(n14645), .A2(n15981), .ZN(n14751) );
  INV_X1 U8838 ( .A(n14733), .ZN(n15241) );
  OR2_X1 U8839 ( .A1(n14928), .A2(n10299), .ZN(n10300) );
  OR2_X1 U8840 ( .A1(n12704), .A2(n11265), .ZN(n10303) );
  OAI211_X1 U8841 ( .C1(n9642), .C2(n8020), .A(n8018), .B(n14934), .ZN(n15153)
         );
  NAND2_X1 U8842 ( .A1(n8024), .A2(n14944), .ZN(n8020) );
  NAND2_X1 U8843 ( .A1(n9642), .A2(n8019), .ZN(n8018) );
  INV_X1 U8844 ( .A(n15146), .ZN(n15368) );
  NAND2_X1 U8845 ( .A1(n14949), .A2(n14948), .ZN(n15372) );
  AOI211_X1 U8846 ( .C1(n15385), .C2(n15880), .A(n15198), .B(n15197), .ZN(
        n15389) );
  AND2_X1 U8847 ( .A1(n7984), .A2(n7983), .ZN(n15225) );
  NAND2_X1 U8848 ( .A1(n15239), .A2(n12668), .ZN(n15222) );
  NAND2_X1 U8849 ( .A1(n7412), .A2(n12729), .ZN(n15236) );
  INV_X1 U8850 ( .A(n14880), .ZN(n15414) );
  NAND2_X1 U8851 ( .A1(n12637), .A2(n12636), .ZN(n15270) );
  NAND2_X1 U8852 ( .A1(n12607), .A2(n12606), .ZN(n15307) );
  NAND2_X1 U8853 ( .A1(n12723), .A2(n12722), .ZN(n15325) );
  NAND2_X1 U8854 ( .A1(n7512), .A2(n7513), .ZN(n15323) );
  NAND2_X1 U8855 ( .A1(n8096), .A2(n12211), .ZN(n12327) );
  NAND2_X1 U8856 ( .A1(n15974), .A2(n12179), .ZN(n12181) );
  NAND2_X1 U8857 ( .A1(n12030), .A2(n12029), .ZN(n15974) );
  INV_X1 U8858 ( .A(n14962), .ZN(n11767) );
  NAND2_X1 U8859 ( .A1(n11623), .A2(n7271), .ZN(n15895) );
  INV_X1 U8860 ( .A(n14959), .ZN(n11624) );
  NAND2_X1 U8861 ( .A1(n11623), .A2(n11622), .ZN(n11625) );
  NAND2_X1 U8862 ( .A1(n8099), .A2(n11621), .ZN(n11714) );
  INV_X1 U8863 ( .A(n15358), .ZN(n15951) );
  NAND2_X1 U8864 ( .A1(n11128), .A2(n11127), .ZN(n11565) );
  NAND2_X1 U8865 ( .A1(n15792), .A2(n10828), .ZN(n10830) );
  NAND2_X1 U8866 ( .A1(n8093), .A2(n14954), .ZN(n15792) );
  INV_X1 U8867 ( .A(n11695), .ZN(n8093) );
  NAND2_X1 U8868 ( .A1(n15760), .A2(n10342), .ZN(n15358) );
  INV_X2 U8869 ( .A(n10825), .ZN(n14776) );
  INV_X1 U8870 ( .A(n15285), .ZN(n15952) );
  AND2_X1 U8871 ( .A1(n15760), .A2(n11264), .ZN(n15947) );
  INV_X1 U8872 ( .A(n15991), .ZN(n15990) );
  NAND2_X1 U8873 ( .A1(n15367), .A2(n7604), .ZN(n7603) );
  INV_X1 U8874 ( .A(n7605), .ZN(n7604) );
  OAI21_X1 U8875 ( .B1(n15368), .B2(n15970), .A(n15366), .ZN(n7605) );
  NAND2_X1 U8876 ( .A1(n7371), .A2(n7370), .ZN(n15457) );
  NAND2_X1 U8877 ( .A1(n15369), .A2(n15973), .ZN(n7371) );
  AND2_X1 U8878 ( .A1(n15376), .A2(n15375), .ZN(n7370) );
  AND2_X1 U8879 ( .A1(n15374), .A2(n15373), .ZN(n15375) );
  AND2_X1 U8880 ( .A1(n15382), .A2(n15381), .ZN(n15383) );
  AND2_X1 U8881 ( .A1(n15380), .A2(n15379), .ZN(n15381) );
  AND2_X2 U8882 ( .A1(n10367), .A2(n10366), .ZN(n15994) );
  INV_X1 U8883 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n15475) );
  OAI211_X1 U8884 ( .C1(n9642), .C2(n8028), .A(n8026), .B(n8021), .ZN(n15482)
         );
  NAND2_X1 U8885 ( .A1(n9642), .A2(n8025), .ZN(n8021) );
  NAND2_X1 U8886 ( .A1(n9642), .A2(n9641), .ZN(n14930) );
  BUF_X1 U8887 ( .A(n10123), .Z(n7409) );
  NOR2_X1 U8888 ( .A1(n7806), .A2(n7805), .ZN(n7804) );
  OR2_X1 U8889 ( .A1(n10293), .A2(P1_U3086), .ZN(n15013) );
  INV_X1 U8890 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n10110) );
  INV_X1 U8891 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12622) );
  NAND2_X1 U8892 ( .A1(n7395), .A2(n10273), .ZN(n10274) );
  INV_X1 U8893 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12609) );
  INV_X1 U8894 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n11236) );
  INV_X1 U8895 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11124) );
  INV_X1 U8896 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11024) );
  INV_X1 U8897 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10198) );
  INV_X1 U8898 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10162) );
  INV_X1 U8899 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10148) );
  INV_X1 U8900 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10102) );
  AND2_X1 U8901 ( .A1(n10094), .A2(n10103), .ZN(n10818) );
  INV_X1 U8902 ( .A(n10065), .ZN(n10335) );
  INV_X1 U8903 ( .A(n10318), .ZN(n7357) );
  NOR2_X1 U8904 ( .A1(n15671), .A2(n9916), .ZN(n15606) );
  XNOR2_X1 U8905 ( .A(n9920), .B(n9921), .ZN(n15610) );
  NAND2_X1 U8906 ( .A1(n9936), .A2(n9937), .ZN(n15628) );
  NAND2_X1 U8907 ( .A1(n15628), .A2(n15629), .ZN(n15625) );
  INV_X1 U8908 ( .A(n7404), .ZN(n9944) );
  NAND2_X1 U8909 ( .A1(n9946), .A2(n9947), .ZN(n15648) );
  AND2_X1 U8910 ( .A1(n7704), .A2(n7708), .ZN(n7703) );
  OR2_X1 U8911 ( .A1(n15661), .A2(n7705), .ZN(n7701) );
  OR2_X1 U8912 ( .A1(n7707), .A2(n7710), .ZN(n7704) );
  INV_X1 U8913 ( .A(n7717), .ZN(n13532) );
  NAND2_X1 U8914 ( .A1(n7569), .A2(n15711), .ZN(n7568) );
  INV_X1 U8915 ( .A(n9740), .ZN(n9741) );
  OAI21_X1 U8916 ( .B1(n13625), .B2(n13960), .A(n9739), .ZN(n9740) );
  NAND2_X1 U8917 ( .A1(n7669), .A2(n7666), .ZN(P3_U3455) );
  NOR2_X1 U8918 ( .A1(n7668), .A2(n7667), .ZN(n7666) );
  OR2_X1 U8919 ( .A1(n13914), .A2(n16008), .ZN(n7669) );
  NOR2_X1 U8920 ( .A1(n16000), .A2(n13915), .ZN(n7667) );
  NAND2_X1 U8921 ( .A1(n8060), .A2(n9719), .ZN(n8055) );
  AOI21_X1 U8922 ( .B1(n8056), .B2(n8057), .A(n8054), .ZN(n8053) );
  INV_X1 U8923 ( .A(n15027), .ZN(n8013) );
  NOR2_X1 U8924 ( .A1(n15028), .A2(n7267), .ZN(n8014) );
  INV_X1 U8925 ( .A(n7693), .ZN(n15666) );
  INV_X1 U8926 ( .A(n15622), .ZN(n15621) );
  INV_X1 U8927 ( .A(n7697), .ZN(n15634) );
  INV_X1 U8928 ( .A(n7698), .ZN(n15650) );
  CLKBUF_X3 U8929 ( .A(n7188), .Z(n9662) );
  AND2_X1 U8930 ( .A1(n7290), .A2(n7936), .ZN(n7203) );
  AND2_X1 U8931 ( .A1(n12898), .A2(n9733), .ZN(n7204) );
  OR2_X1 U8932 ( .A1(n7907), .A2(n9328), .ZN(n7205) );
  OR2_X1 U8933 ( .A1(n14418), .A2(n14066), .ZN(n7206) );
  AND2_X1 U8934 ( .A1(n9408), .A2(n13988), .ZN(n7207) );
  INV_X1 U8935 ( .A(n12926), .ZN(n7766) );
  NAND2_X1 U8936 ( .A1(n14418), .A2(n14302), .ZN(n7208) );
  AND2_X1 U8937 ( .A1(n12317), .A2(n9762), .ZN(n7209) );
  INV_X1 U8938 ( .A(n12724), .ZN(n7972) );
  AND2_X1 U8939 ( .A1(n12440), .A2(n12439), .ZN(n7210) );
  INV_X1 U8940 ( .A(n13075), .ZN(n7752) );
  XNOR2_X1 U8941 ( .A(n12854), .B(n12795), .ZN(n11342) );
  AND2_X1 U8942 ( .A1(n7919), .A2(n7913), .ZN(n7211) );
  AND2_X1 U8943 ( .A1(n7477), .A2(n13481), .ZN(n7212) );
  NAND2_X1 U8944 ( .A1(n9117), .A2(n9116), .ZN(n12797) );
  INV_X1 U8945 ( .A(n12425), .ZN(n7820) );
  AND2_X1 U8946 ( .A1(n7886), .A2(n7269), .ZN(n7213) );
  OR2_X1 U8947 ( .A1(n8688), .A2(n13829), .ZN(n7214) );
  OR3_X1 U8948 ( .A1(n14274), .A2(n14407), .A3(n14403), .ZN(n7215) );
  INV_X1 U8949 ( .A(n11856), .ZN(n13483) );
  AND4_X1 U8950 ( .A1(n8339), .A2(n8338), .A3(n8337), .A4(n8336), .ZN(n11856)
         );
  INV_X1 U8951 ( .A(n11009), .ZN(n7878) );
  AND2_X1 U8952 ( .A1(n13790), .A2(n12977), .ZN(n13818) );
  NOR2_X1 U8953 ( .A1(n14272), .A2(n12505), .ZN(n7216) );
  NAND2_X1 U8954 ( .A1(n7375), .A2(n7374), .ZN(n7217) );
  INV_X1 U8955 ( .A(n9504), .ZN(n8077) );
  AND2_X1 U8956 ( .A1(n11547), .A2(n11554), .ZN(n7218) );
  AND2_X1 U8957 ( .A1(n8059), .A2(n9717), .ZN(n7219) );
  INV_X1 U8958 ( .A(n9406), .ZN(n7895) );
  AND2_X1 U8959 ( .A1(n9540), .A2(n9539), .ZN(n7220) );
  INV_X1 U8960 ( .A(n7187), .ZN(n8111) );
  INV_X1 U8961 ( .A(n13067), .ZN(n7664) );
  INV_X1 U8962 ( .A(n12952), .ZN(n12948) );
  AND2_X1 U8963 ( .A1(n12566), .A2(n12380), .ZN(n12952) );
  INV_X1 U8964 ( .A(n12832), .ZN(n12811) );
  NAND2_X2 U8965 ( .A1(n10163), .A2(n7891), .ZN(n12832) );
  OR2_X1 U8966 ( .A1(n13540), .A2(n7392), .ZN(n7221) );
  XNOR2_X1 U8967 ( .A(n8709), .B(P3_IR_REG_24__SCAN_IN), .ZN(n8719) );
  OR2_X1 U8968 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8207), .ZN(n7222) );
  XNOR2_X1 U8969 ( .A(n8660), .B(P3_IR_REG_21__SCAN_IN), .ZN(n8747) );
  INV_X1 U8970 ( .A(n7480), .ZN(n8251) );
  NAND2_X1 U8971 ( .A1(n7585), .A2(n14067), .ZN(n7223) );
  AND2_X1 U8972 ( .A1(n15246), .A2(n7611), .ZN(n7224) );
  AND2_X1 U8973 ( .A1(n12924), .A2(n12923), .ZN(n13054) );
  OR2_X1 U8974 ( .A1(n12428), .A2(n7821), .ZN(n7225) );
  NOR2_X1 U8975 ( .A1(n15872), .A2(n11821), .ZN(n7226) );
  INV_X1 U8976 ( .A(n15378), .ZN(n15177) );
  NAND2_X1 U8977 ( .A1(n12700), .A2(n12699), .ZN(n15378) );
  AND2_X1 U8978 ( .A1(n9225), .A2(n7206), .ZN(n7227) );
  OR2_X1 U8979 ( .A1(n7895), .A2(n7894), .ZN(n7228) );
  AND2_X1 U8980 ( .A1(n9524), .A2(n9523), .ZN(n7229) );
  NAND3_X1 U8981 ( .A1(n9018), .A2(n9017), .A3(n8145), .ZN(n11081) );
  NOR2_X1 U8982 ( .A1(n12999), .A2(n13718), .ZN(n7230) );
  AND2_X1 U8983 ( .A1(n11428), .A2(n8007), .ZN(n7231) );
  INV_X1 U8984 ( .A(n15003), .ZN(n7631) );
  NAND2_X1 U8985 ( .A1(n8520), .A2(n8519), .ZN(n7232) );
  AND4_X1 U8986 ( .A1(n9992), .A2(n9991), .A3(n7396), .A4(n10107), .ZN(n7233)
         );
  AND2_X1 U8987 ( .A1(n12232), .A2(n12233), .ZN(n7234) );
  OR2_X1 U8988 ( .A1(n13638), .A2(n9970), .ZN(n13009) );
  NOR2_X1 U8989 ( .A1(n11416), .A2(n7836), .ZN(n7235) );
  OR2_X1 U8990 ( .A1(n14183), .A2(n14190), .ZN(n7236) );
  NAND2_X1 U8991 ( .A1(n12062), .A2(n9379), .ZN(n7237) );
  AND2_X1 U8992 ( .A1(n11798), .A2(n11797), .ZN(n7238) );
  NAND2_X1 U8993 ( .A1(n9951), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7239) );
  NAND2_X1 U8994 ( .A1(n7851), .A2(n8194), .ZN(n8416) );
  INV_X1 U8995 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8363) );
  INV_X1 U8996 ( .A(n7968), .ZN(n7967) );
  NAND2_X1 U8997 ( .A1(n7972), .A2(n7973), .ZN(n7968) );
  OR2_X1 U8998 ( .A1(n13145), .A2(n9530), .ZN(n7240) );
  AND2_X1 U8999 ( .A1(n13225), .A2(n9799), .ZN(n7241) );
  NAND2_X1 U9000 ( .A1(n8916), .A2(n8915), .ZN(n14377) );
  INV_X1 U9001 ( .A(n14377), .ZN(n14183) );
  OR2_X1 U9002 ( .A1(n15995), .A2(n13256), .ZN(n7242) );
  INV_X1 U9003 ( .A(n11779), .ZN(n12116) );
  AND2_X1 U9004 ( .A1(n14418), .A2(n14066), .ZN(n7243) );
  NAND2_X1 U9005 ( .A1(n11879), .A2(n12794), .ZN(n7244) );
  OR2_X1 U9006 ( .A1(n14191), .A2(n14377), .ZN(n7245) );
  NAND2_X1 U9007 ( .A1(n14350), .A2(n14068), .ZN(n7246) );
  INV_X1 U9008 ( .A(n14844), .ZN(n8115) );
  INV_X1 U9009 ( .A(n14795), .ZN(n8120) );
  OR2_X1 U9010 ( .A1(n7507), .A2(n7506), .ZN(n7247) );
  OR2_X1 U9011 ( .A1(n12539), .A2(n13834), .ZN(n7248) );
  INV_X1 U9012 ( .A(n14632), .ZN(n7798) );
  INV_X1 U9013 ( .A(n14929), .ZN(n7378) );
  INV_X1 U9014 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8877) );
  INV_X1 U9015 ( .A(n8034), .ZN(n8033) );
  OAI21_X1 U9016 ( .B1(n8036), .B2(n8035), .A(n8938), .ZN(n8034) );
  AND2_X1 U9017 ( .A1(n7222), .A2(n8585), .ZN(n7250) );
  AND2_X1 U9018 ( .A1(n9093), .A2(n9080), .ZN(n7251) );
  NOR2_X1 U9019 ( .A1(n14043), .A2(n12829), .ZN(n7252) );
  AND2_X1 U9020 ( .A1(n12352), .A2(n12029), .ZN(n7253) );
  AND2_X1 U9021 ( .A1(n9551), .A2(n9550), .ZN(n7254) );
  OR2_X1 U9022 ( .A1(n14786), .A2(n14785), .ZN(n7255) );
  AND2_X1 U9023 ( .A1(n8179), .A2(n8177), .ZN(n7256) );
  OR2_X1 U9024 ( .A1(n14333), .A2(n14356), .ZN(n7257) );
  NOR2_X1 U9025 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7258) );
  OR2_X1 U9026 ( .A1(n9125), .A2(n15904), .ZN(n7259) );
  OR2_X1 U9027 ( .A1(n12473), .A2(n12394), .ZN(n7260) );
  OR2_X1 U9028 ( .A1(n7963), .A2(n7962), .ZN(n7261) );
  OR2_X1 U9029 ( .A1(n14392), .A2(n14221), .ZN(n9312) );
  OR2_X1 U9030 ( .A1(n9564), .A2(n7334), .ZN(n7262) );
  INV_X1 U9031 ( .A(n7899), .ZN(n7898) );
  INV_X1 U9032 ( .A(n7577), .ZN(n14225) );
  NOR3_X1 U9033 ( .A1(n14274), .A2(n14403), .A3(n7579), .ZN(n7577) );
  AND2_X1 U9034 ( .A1(n8092), .A2(n10828), .ZN(n7263) );
  AND2_X1 U9035 ( .A1(n9042), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7264) );
  INV_X1 U9036 ( .A(n15232), .ZN(n15398) );
  NAND2_X1 U9037 ( .A1(n12672), .A2(n12671), .ZN(n15232) );
  AND2_X1 U9038 ( .A1(n13005), .A2(n13006), .ZN(n7265) );
  INV_X1 U9039 ( .A(n7531), .ZN(n14042) );
  NAND2_X1 U9040 ( .A1(n12827), .A2(n12826), .ZN(n7531) );
  INV_X1 U9041 ( .A(n14827), .ZN(n8126) );
  OR2_X1 U9042 ( .A1(n12379), .A2(n15885), .ZN(n7266) );
  AND2_X1 U9043 ( .A1(n8015), .A2(n15029), .ZN(n7267) );
  INV_X1 U9044 ( .A(n14863), .ZN(n8123) );
  OR2_X1 U9045 ( .A1(n10638), .A2(n15809), .ZN(n7268) );
  INV_X1 U9046 ( .A(n14879), .ZN(n8117) );
  NAND2_X1 U9047 ( .A1(n12807), .A2(n12806), .ZN(n7269) );
  NAND2_X1 U9048 ( .A1(n13823), .A2(n8687), .ZN(n7270) );
  AND2_X1 U9049 ( .A1(n11624), .A2(n11622), .ZN(n7271) );
  OR2_X1 U9050 ( .A1(n9510), .A2(n9509), .ZN(n7272) );
  XOR2_X1 U9051 ( .A(n8719), .B(P3_B_REG_SCAN_IN), .Z(n7273) );
  INV_X1 U9052 ( .A(n7448), .ZN(n7447) );
  OR2_X1 U9053 ( .A1(n8120), .A2(n14794), .ZN(n7274) );
  OR2_X1 U9054 ( .A1(n14805), .A2(n14807), .ZN(n7275) );
  AND2_X1 U9055 ( .A1(n11950), .A2(n7446), .ZN(n7276) );
  NAND2_X1 U9056 ( .A1(n7214), .A2(n7270), .ZN(n7774) );
  AND2_X1 U9057 ( .A1(n7623), .A2(n8819), .ZN(n7277) );
  AND2_X1 U9058 ( .A1(n7478), .A2(n10572), .ZN(n7278) );
  NAND2_X1 U9059 ( .A1(n8067), .A2(n9187), .ZN(n9355) );
  AND2_X1 U9060 ( .A1(n14258), .A2(n7430), .ZN(n7279) );
  NOR2_X1 U9061 ( .A1(n14274), .A2(n14407), .ZN(n14243) );
  AND2_X1 U9062 ( .A1(n13082), .A2(n7204), .ZN(n7280) );
  NOR2_X1 U9063 ( .A1(n15904), .A2(n14073), .ZN(n7281) );
  NOR2_X1 U9064 ( .A1(n15436), .A2(n14676), .ZN(n7282) );
  NOR2_X1 U9065 ( .A1(n13913), .A2(n13248), .ZN(n7283) );
  INV_X1 U9066 ( .A(n9479), .ZN(n8070) );
  INV_X1 U9067 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9187) );
  INV_X1 U9068 ( .A(n9328), .ZN(n7910) );
  NOR2_X1 U9069 ( .A1(n14386), .A2(n14063), .ZN(n9328) );
  NAND2_X1 U9070 ( .A1(n9786), .A2(n9779), .ZN(n7284) );
  NAND2_X1 U9071 ( .A1(n13043), .A2(n13009), .ZN(n7285) );
  AND2_X1 U9072 ( .A1(n11567), .A2(n15049), .ZN(n7286) );
  NOR2_X1 U9073 ( .A1(n14272), .A2(n14251), .ZN(n7287) );
  NAND3_X1 U9074 ( .A1(n7480), .A2(n7783), .A3(n8012), .ZN(n7288) );
  AND2_X1 U9075 ( .A1(n7757), .A2(n7285), .ZN(n7289) );
  OR2_X1 U9076 ( .A1(n12797), .A2(n12851), .ZN(n7290) );
  OR2_X1 U9077 ( .A1(n8131), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n7291) );
  AND2_X1 U9078 ( .A1(n8789), .A2(SI_8_), .ZN(n7292) );
  AND2_X1 U9079 ( .A1(n10422), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7293) );
  INV_X1 U9080 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U9081 ( .A1(n15016), .A2(n15015), .ZN(n7294) );
  AND2_X1 U9082 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n7295) );
  AND2_X1 U9083 ( .A1(n7228), .A2(n11951), .ZN(n7296) );
  OAI21_X1 U9084 ( .B1(n8106), .B2(n8104), .A(n8138), .ZN(n8103) );
  AND2_X1 U9085 ( .A1(n14623), .A2(n14622), .ZN(n7297) );
  INV_X1 U9086 ( .A(n7680), .ZN(n7679) );
  OAI21_X1 U9087 ( .B1(n12931), .B2(n7681), .A(n15866), .ZN(n7680) );
  INV_X1 U9088 ( .A(n7928), .ZN(n7927) );
  AND2_X1 U9089 ( .A1(n7236), .A2(n14167), .ZN(n7928) );
  AND2_X1 U9090 ( .A1(n10966), .A2(n10960), .ZN(n7298) );
  AND2_X1 U9091 ( .A1(n7240), .A2(n7917), .ZN(n7299) );
  NAND2_X1 U9092 ( .A1(n7223), .A2(n9386), .ZN(n7300) );
  INV_X1 U9093 ( .A(n7776), .ZN(n7775) );
  NAND2_X1 U9094 ( .A1(n7214), .A2(n13070), .ZN(n7776) );
  INV_X1 U9095 ( .A(n9541), .ZN(n8073) );
  AND2_X1 U9096 ( .A1(n7925), .A2(n9712), .ZN(n7301) );
  AND2_X1 U9097 ( .A1(n12606), .A2(n12724), .ZN(n7302) );
  OR2_X1 U9098 ( .A1(n9554), .A2(n7254), .ZN(n7303) );
  INV_X1 U9099 ( .A(n13649), .ZN(n7560) );
  NAND2_X1 U9100 ( .A1(n13009), .A2(n13010), .ZN(n13075) );
  OR2_X1 U9101 ( .A1(n13870), .A2(n13743), .ZN(n7304) );
  AND2_X1 U9102 ( .A1(n8043), .A2(n8146), .ZN(n7305) );
  AND2_X1 U9103 ( .A1(n7798), .A2(n7794), .ZN(n7306) );
  NOR2_X1 U9104 ( .A1(n12349), .A2(n8095), .ZN(n7307) );
  AND2_X1 U9105 ( .A1(n12443), .A2(n12442), .ZN(n7308) );
  INV_X1 U9106 ( .A(n10634), .ZN(n10799) );
  AND2_X1 U9107 ( .A1(n8349), .A2(n8364), .ZN(n10634) );
  INV_X1 U9108 ( .A(n11970), .ZN(n7958) );
  AND2_X1 U9109 ( .A1(n7979), .A2(n11581), .ZN(n7309) );
  AND2_X1 U9110 ( .A1(n9502), .A2(n9501), .ZN(n7310) );
  OR2_X1 U9111 ( .A1(n14901), .A2(n14899), .ZN(n7311) );
  OR2_X1 U9112 ( .A1(n8126), .A2(n14826), .ZN(n7312) );
  AND2_X1 U9113 ( .A1(n15261), .A2(n12653), .ZN(n7313) );
  OR2_X1 U9114 ( .A1(n8117), .A2(n14878), .ZN(n7314) );
  AND2_X1 U9115 ( .A1(n8353), .A2(n8332), .ZN(n7315) );
  OR2_X1 U9116 ( .A1(n14862), .A2(n8123), .ZN(n7316) );
  OR2_X1 U9117 ( .A1(n8115), .A2(n14843), .ZN(n7317) );
  AND2_X1 U9118 ( .A1(n7571), .A2(n7567), .ZN(n7318) );
  INV_X1 U9119 ( .A(n13073), .ZN(n13745) );
  AND2_X1 U9120 ( .A1(n12992), .A2(n13717), .ZN(n13073) );
  OR2_X1 U9121 ( .A1(n8113), .A2(n14816), .ZN(n7319) );
  OR2_X1 U9122 ( .A1(n7229), .A2(n8089), .ZN(n7320) );
  OR2_X1 U9123 ( .A1(n9395), .A2(n7207), .ZN(n7321) );
  OR2_X1 U9124 ( .A1(n8081), .A2(n7333), .ZN(n7322) );
  AND2_X1 U9125 ( .A1(n10033), .A2(n10028), .ZN(n7323) );
  AND2_X1 U9126 ( .A1(n7233), .A2(n10130), .ZN(n7324) );
  AND2_X1 U9127 ( .A1(n7550), .A2(n8182), .ZN(n7325) );
  AND2_X1 U9128 ( .A1(n13986), .A2(n7340), .ZN(n7884) );
  INV_X1 U9129 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n10113) );
  INV_X1 U9130 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8219) );
  NOR2_X1 U9131 ( .A1(n7471), .A2(n7470), .ZN(n7326) );
  OR2_X1 U9132 ( .A1(n8073), .A2(n7220), .ZN(n7327) );
  INV_X1 U9133 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8010) );
  INV_X1 U9134 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8985) );
  OR2_X1 U9135 ( .A1(n13930), .A2(n13929), .ZN(P3_U3451) );
  OR2_X1 U9136 ( .A1(n13861), .A2(n13860), .ZN(P3_U3483) );
  INV_X1 U9137 ( .A(n13065), .ZN(n7665) );
  NAND2_X1 U9138 ( .A1(n14762), .A2(n14765), .ZN(n10525) );
  AND4_X1 U9139 ( .A1(n8379), .A2(n8378), .A3(n8377), .A4(n8376), .ZN(n12256)
         );
  INV_X1 U9140 ( .A(n12256), .ZN(n7681) );
  NAND2_X1 U9141 ( .A1(n12737), .A2(n7888), .ZN(n7885) );
  INV_X1 U9142 ( .A(n9168), .ZN(n9637) );
  AND2_X1 U9143 ( .A1(n8717), .A2(n8716), .ZN(n8722) );
  AND2_X1 U9144 ( .A1(n12480), .A2(n9779), .ZN(n13193) );
  INV_X1 U9145 ( .A(n15333), .ZN(n7975) );
  AND2_X1 U9146 ( .A1(n7480), .A2(n7783), .ZN(n8441) );
  NAND2_X1 U9147 ( .A1(n12117), .A2(n12120), .ZN(n12441) );
  NAND2_X1 U9148 ( .A1(n13138), .A2(n11796), .ZN(n11801) );
  AND2_X1 U9149 ( .A1(n8483), .A2(n8204), .ZN(n7330) );
  NAND2_X1 U9150 ( .A1(n12381), .A2(n12950), .ZN(n12550) );
  NAND2_X1 U9151 ( .A1(n15929), .A2(n11970), .ZN(n12026) );
  NAND2_X1 U9152 ( .A1(n7761), .A2(n12948), .ZN(n12514) );
  XOR2_X1 U9153 ( .A(n13933), .B(n9806), .Z(n7331) );
  NAND2_X1 U9154 ( .A1(n8404), .A2(n8425), .ZN(n11553) );
  NAND2_X1 U9155 ( .A1(n7480), .A2(n7481), .ZN(n8458) );
  AND2_X1 U9156 ( .A1(n8383), .A2(n8386), .ZN(n7485) );
  INV_X1 U9157 ( .A(n9797), .ZN(n7456) );
  NAND2_X1 U9158 ( .A1(n8922), .A2(n8921), .ZN(n14190) );
  NOR2_X1 U9159 ( .A1(n13743), .A2(n7331), .ZN(n7332) );
  AND2_X1 U9160 ( .A1(n9581), .A2(n9580), .ZN(n7333) );
  AND2_X1 U9161 ( .A1(n9562), .A2(n9561), .ZN(n7334) );
  NAND2_X1 U9162 ( .A1(n12893), .A2(n12911), .ZN(n8680) );
  AND2_X1 U9163 ( .A1(n10988), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7335) );
  AND2_X1 U9164 ( .A1(n7969), .A2(n7973), .ZN(n7336) );
  INV_X1 U9165 ( .A(n7586), .ZN(n14329) );
  NOR2_X1 U9166 ( .A1(n14341), .A2(n14428), .ZN(n7586) );
  OR2_X1 U9167 ( .A1(n8496), .A2(n7872), .ZN(n7337) );
  NOR2_X1 U9168 ( .A1(n9968), .A2(n9816), .ZN(n7338) );
  AND2_X1 U9169 ( .A1(n7818), .A2(n7814), .ZN(n7339) );
  NAND2_X1 U9170 ( .A1(n12831), .A2(n12830), .ZN(n7340) );
  INV_X1 U9171 ( .A(n14828), .ZN(n7606) );
  INV_X1 U9172 ( .A(n13501), .ZN(n7566) );
  XOR2_X1 U9173 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .Z(n7341) );
  NAND2_X1 U9174 ( .A1(n8002), .A2(n8721), .ZN(n9743) );
  OAI21_X1 U9175 ( .B1(n11131), .B2(n7501), .A(n7499), .ZN(n11616) );
  INV_X1 U9176 ( .A(n15445), .ZN(n7617) );
  INV_X1 U9177 ( .A(n15436), .ZN(n7615) );
  AND2_X1 U9178 ( .A1(n8572), .A2(n8571), .ZN(n13727) );
  NAND2_X1 U9179 ( .A1(n8090), .A2(n8091), .ZN(n11131) );
  AND2_X1 U9180 ( .A1(n11426), .A2(n8005), .ZN(n7342) );
  AND2_X1 U9181 ( .A1(n12367), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7343) );
  AND2_X1 U9182 ( .A1(n7832), .A2(n7833), .ZN(n7344) );
  OR2_X1 U9183 ( .A1(n11343), .A2(n11342), .ZN(n7345) );
  AND2_X1 U9184 ( .A1(n9624), .A2(n13977), .ZN(n7346) );
  AND2_X1 U9185 ( .A1(n8857), .A2(SI_26_), .ZN(n7347) );
  OR2_X1 U9186 ( .A1(n11086), .A2(n9751), .ZN(n7454) );
  INV_X1 U9187 ( .A(n13727), .ZN(n13690) );
  INV_X1 U9188 ( .A(n13579), .ZN(n7561) );
  NAND2_X2 U9189 ( .A1(n9360), .A2(n9722), .ZN(n10019) );
  INV_X1 U9190 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7845) );
  INV_X1 U9191 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7848) );
  AND2_X1 U9192 ( .A1(n9452), .A2(n11868), .ZN(n9444) );
  INV_X1 U9193 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U9194 ( .A1(n12894), .A2(n12902), .ZN(n8678) );
  INV_X1 U9195 ( .A(n13541), .ZN(n13564) );
  XOR2_X1 U9196 ( .A(n11775), .B(n11776), .Z(n7348) );
  AND2_X1 U9197 ( .A1(n14127), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7349) );
  INV_X1 U9198 ( .A(n12408), .ZN(n7993) );
  OR2_X1 U9199 ( .A1(n14117), .A2(n14118), .ZN(n7350) );
  AND2_X1 U9200 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n12682), .ZN(n7351) );
  INV_X1 U9201 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12490) );
  INV_X1 U9202 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8878) );
  AND2_X1 U9203 ( .A1(n7743), .A2(n13601), .ZN(n7352) );
  NAND2_X1 U9204 ( .A1(n7718), .A2(n10599), .ZN(n7727) );
  NOR2_X1 U9205 ( .A1(n8901), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n14471) );
  INV_X1 U9206 ( .A(n12202), .ZN(n8060) );
  INV_X1 U9207 ( .A(SI_4_), .ZN(n7622) );
  INV_X1 U9208 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7841) );
  INV_X1 U9209 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7694) );
  INV_X1 U9210 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U9211 ( .A1(n14842), .A2(n14841), .ZN(n7353) );
  NAND2_X1 U9212 ( .A1(n14838), .A2(n14837), .ZN(n7354) );
  NAND2_X1 U9213 ( .A1(n14877), .A2(n14876), .ZN(n7355) );
  NAND2_X1 U9214 ( .A1(n14873), .A2(n14872), .ZN(n7356) );
  NOR2_X1 U9215 ( .A1(n7358), .A2(n7357), .ZN(n15485) );
  INV_X1 U9216 ( .A(n10317), .ZN(n7358) );
  INV_X1 U9217 ( .A(n14988), .ZN(n7394) );
  INV_X2 U9218 ( .A(n8995), .ZN(n12638) );
  AOI21_X1 U9219 ( .B1(n14913), .B2(n14912), .A(n14911), .ZN(n14914) );
  NAND2_X1 U9220 ( .A1(n7388), .A2(n7255), .ZN(n14790) );
  NAND2_X1 U9221 ( .A1(n7360), .A2(n8112), .ZN(n14820) );
  NAND2_X1 U9222 ( .A1(n8121), .A2(n8122), .ZN(n14866) );
  NAND2_X1 U9223 ( .A1(n14779), .A2(n14780), .ZN(n14778) );
  NAND4_X1 U9224 ( .A1(n14774), .A2(n14775), .A3(n14773), .A4(n14772), .ZN(
        n14779) );
  NAND2_X1 U9225 ( .A1(n14866), .A2(n14867), .ZN(n14865) );
  NAND2_X1 U9226 ( .A1(n14799), .A2(n14800), .ZN(n14798) );
  NAND2_X1 U9227 ( .A1(n14820), .A2(n14821), .ZN(n14819) );
  NAND2_X1 U9228 ( .A1(n14790), .A2(n14791), .ZN(n14789) );
  XNOR2_X1 U9229 ( .A(n9082), .B(n9081), .ZN(n11292) );
  AOI21_X2 U9230 ( .B1(n14739), .B2(n14740), .A(n7359), .ZN(n14661) );
  NAND2_X1 U9231 ( .A1(n14570), .A2(n14681), .ZN(n14683) );
  NOR2_X2 U9232 ( .A1(n12275), .A2(n12276), .ZN(n12274) );
  AND2_X1 U9233 ( .A1(n14492), .A2(n14491), .ZN(n7359) );
  AND2_X4 U9234 ( .A1(n14581), .A2(n11729), .ZN(n14563) );
  INV_X1 U9235 ( .A(n10768), .ZN(n10766) );
  NAND2_X1 U9236 ( .A1(n14726), .A2(n14730), .ZN(n14625) );
  NAND2_X1 U9237 ( .A1(n14712), .A2(n14521), .ZN(n14612) );
  NAND3_X1 U9238 ( .A1(n7398), .A2(n7319), .A3(n7397), .ZN(n7360) );
  NAND2_X1 U9239 ( .A1(n7394), .A2(n7187), .ZN(n7393) );
  NAND2_X1 U9240 ( .A1(n7361), .A2(n7265), .ZN(n13008) );
  OR2_X1 U9241 ( .A1(n13007), .A2(n13012), .ZN(n7361) );
  MUX2_X1 U9242 ( .A(n10524), .B(n10042), .S(n10505), .Z(n11217) );
  INV_X1 U9243 ( .A(n7779), .ZN(n12900) );
  AOI21_X1 U9244 ( .B1(n12914), .B2(n13002), .A(n12913), .ZN(n12918) );
  OAI21_X1 U9245 ( .B1(n12907), .B2(n12906), .A(n12905), .ZN(n12912) );
  NOR3_X1 U9246 ( .A1(n12996), .A2(n13728), .A3(n12995), .ZN(n13001) );
  AOI22_X1 U9247 ( .A1(n12960), .A2(n13065), .B1(n12959), .B2(n12958), .ZN(
        n12966) );
  AOI211_X1 U9248 ( .C1(n12975), .C2(n12974), .A(n13795), .B(n12973), .ZN(
        n12987) );
  AND3_X1 U9249 ( .A1(n7362), .A2(n7242), .A3(n13017), .ZN(n13038) );
  NAND2_X1 U9250 ( .A1(n12476), .A2(n12475), .ZN(n12474) );
  NAND2_X1 U9251 ( .A1(n10438), .A2(n9047), .ZN(n10776) );
  NAND2_X1 U9252 ( .A1(n7385), .A2(n13086), .ZN(n13094) );
  NAND2_X1 U9253 ( .A1(n9110), .A2(n11341), .ZN(n7433) );
  OAI21_X1 U9254 ( .B1(n14376), .B2(n14442), .A(n14374), .ZN(n7425) );
  NAND2_X1 U9255 ( .A1(n8765), .A2(n8766), .ZN(n8767) );
  NAND2_X1 U9256 ( .A1(n8824), .A2(n8823), .ZN(n9204) );
  NAND2_X1 U9257 ( .A1(n8838), .A2(n7656), .ZN(n7652) );
  NAND2_X1 U9258 ( .A1(n7503), .A2(n7502), .ZN(n15215) );
  NAND2_X1 U9259 ( .A1(n7367), .A2(n7366), .ZN(n11466) );
  INV_X1 U9260 ( .A(n11464), .ZN(n7367) );
  NAND3_X1 U9261 ( .A1(n14166), .A2(n7368), .A3(n14358), .ZN(n14169) );
  NAND2_X1 U9262 ( .A1(n7938), .A2(n7937), .ZN(n14317) );
  NAND2_X1 U9263 ( .A1(n14299), .A2(n7950), .ZN(n7947) );
  NAND3_X1 U9264 ( .A1(n9579), .A2(n7217), .A3(n7322), .ZN(n8079) );
  OR3_X2 U9265 ( .A1(n9497), .A2(n9500), .A3(n8076), .ZN(n8074) );
  NAND2_X1 U9266 ( .A1(n8082), .A2(n8083), .ZN(n9499) );
  NAND2_X1 U9267 ( .A1(n7373), .A2(n7372), .ZN(n9547) );
  NAND2_X1 U9268 ( .A1(n9593), .A2(n9592), .ZN(n9598) );
  NAND3_X1 U9269 ( .A1(n9538), .A2(n9537), .A3(n7327), .ZN(n7373) );
  OAI22_X1 U9270 ( .A1(n9609), .A2(n9608), .B1(n9614), .B2(n9613), .ZN(n9620)
         );
  INV_X1 U9271 ( .A(n7375), .ZN(n9578) );
  NAND3_X1 U9272 ( .A1(n9548), .A2(n8152), .A3(n7303), .ZN(n8064) );
  NAND2_X2 U9273 ( .A1(n9444), .A2(n9720), .ZN(n9529) );
  NAND2_X1 U9274 ( .A1(n7984), .A2(n7980), .ZN(n15223) );
  INV_X1 U9275 ( .A(n7624), .ZN(n8928) );
  AOI21_X1 U9276 ( .B1(n15176), .B2(n15378), .A(n15161), .ZN(n15162) );
  AOI22_X1 U9277 ( .A1(n15207), .A2(n15206), .B1(n15035), .B2(n15392), .ZN(
        n15188) );
  OAI211_X1 U9278 ( .C1(n9716), .C2(n8055), .A(n8053), .B(n8052), .ZN(P2_U3328) );
  NOR2_X2 U9279 ( .A1(n13641), .A2(n13640), .ZN(n13845) );
  NAND2_X1 U9280 ( .A1(n7758), .A2(n13073), .ZN(n13748) );
  NAND2_X1 U9281 ( .A1(n11248), .A2(n11247), .ZN(n11246) );
  NOR2_X1 U9282 ( .A1(n13844), .A2(n7670), .ZN(n13914) );
  INV_X2 U9283 ( .A(n8292), .ZN(n8305) );
  NAND2_X2 U9284 ( .A1(n14924), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n10302) );
  INV_X1 U9285 ( .A(n14817), .ZN(n8113) );
  NAND2_X2 U9286 ( .A1(n13159), .A2(n10297), .ZN(n14928) );
  CLKBUF_X1 U9287 ( .A(n15053), .Z(n7377) );
  XNOR2_X1 U9288 ( .A(n9027), .B(n9026), .ZN(n10065) );
  NAND2_X1 U9289 ( .A1(n11447), .A2(n12893), .ZN(n11248) );
  NAND2_X1 U9290 ( .A1(n7422), .A2(n10634), .ZN(n7729) );
  NOR2_X1 U9291 ( .A1(n12289), .A2(n12288), .ZN(n13507) );
  INV_X1 U9292 ( .A(n11546), .ZN(n7423) );
  NAND2_X1 U9293 ( .A1(n13572), .A2(n7743), .ZN(n7742) );
  OAI211_X1 U9294 ( .C1(n13614), .C2(n15718), .A(n7568), .B(n7318), .ZN(
        P3_U3201) );
  OR2_X1 U9295 ( .A1(n10336), .A2(n10325), .ZN(n10326) );
  INV_X1 U9296 ( .A(n14759), .ZN(n14763) );
  CLKBUF_X2 U9297 ( .A(n15055), .Z(n7381) );
  NAND3_X1 U9298 ( .A1(n7382), .A2(n14782), .A3(n14954), .ZN(n7388) );
  NAND2_X1 U9299 ( .A1(n14778), .A2(n14777), .ZN(n7382) );
  NAND3_X1 U9300 ( .A1(n7780), .A2(n7386), .A3(n7249), .ZN(n7385) );
  NAND2_X1 U9301 ( .A1(n8215), .A2(n7847), .ZN(n8648) );
  NAND2_X1 U9302 ( .A1(n7558), .A2(n8189), .ZN(n8250) );
  NAND2_X1 U9303 ( .A1(n7860), .A2(n7859), .ZN(n8238) );
  INV_X1 U9304 ( .A(n7757), .ZN(n7754) );
  INV_X1 U9305 ( .A(n7750), .ZN(n7749) );
  NAND2_X1 U9306 ( .A1(n7498), .A2(n7324), .ZN(n7608) );
  NAND2_X1 U9307 ( .A1(n15623), .A2(n15624), .ZN(n15620) );
  XNOR2_X1 U9308 ( .A(n9908), .B(n9907), .ZN(n9909) );
  NAND2_X2 U9309 ( .A1(n14317), .A2(n7257), .ZN(n14299) );
  NAND2_X1 U9310 ( .A1(n15651), .A2(n15652), .ZN(n7700) );
  NAND2_X1 U9311 ( .A1(n15645), .A2(n15647), .ZN(n15651) );
  NAND2_X1 U9312 ( .A1(n14375), .A2(n7424), .ZN(n14456) );
  XNOR2_X2 U9313 ( .A(n8790), .B(SI_9_), .ZN(n8973) );
  INV_X1 U9314 ( .A(n7945), .ZN(n14201) );
  NAND3_X1 U9315 ( .A1(n7885), .A2(n14007), .A3(n7213), .ZN(n14006) );
  NAND2_X1 U9316 ( .A1(n8769), .A2(n8768), .ZN(n9027) );
  NAND2_X1 U9317 ( .A1(n7198), .A2(n7396), .ZN(n10277) );
  NAND2_X2 U9318 ( .A1(n14651), .A2(n14580), .ZN(n14727) );
  INV_X1 U9319 ( .A(n7818), .ZN(n7817) );
  INV_X1 U9320 ( .A(n7822), .ZN(n14492) );
  NAND2_X1 U9321 ( .A1(n14105), .A2(n14106), .ZN(n14109) );
  NOR2_X1 U9322 ( .A1(n14125), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n14143) );
  AOI21_X1 U9323 ( .B1(n7390), .B2(n15583), .A(n14149), .ZN(n14150) );
  XNOR2_X1 U9324 ( .A(n14144), .B(n7391), .ZN(n7390) );
  AOI21_X1 U9325 ( .B1(n15557), .B2(P2_REG2_REG_7__SCAN_IN), .A(n15552), .ZN(
        n10866) );
  AOI21_X1 U9326 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n15535), .A(n15530), .ZN(
        n15543) );
  AOI21_X1 U9327 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n15597), .A(n15591), .ZN(
        n11524) );
  NAND2_X1 U9328 ( .A1(n9934), .A2(n9935), .ZN(n15623) );
  NAND2_X1 U9329 ( .A1(n10134), .A2(n8135), .ZN(n15479) );
  NAND2_X1 U9330 ( .A1(n15708), .A2(n15709), .ZN(n15707) );
  AOI21_X1 U9331 ( .B1(n14910), .B2(n14909), .A(n14908), .ZN(n14911) );
  NOR2_X1 U9332 ( .A1(n13606), .A2(n13605), .ZN(n7570) );
  XNOR2_X1 U9333 ( .A(n7570), .B(n13607), .ZN(n7569) );
  AOI21_X2 U9334 ( .B1(n15775), .B2(n15053), .A(n14992), .ZN(n14768) );
  INV_X1 U9335 ( .A(n10277), .ZN(n7395) );
  INV_X1 U9336 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7396) );
  NAND3_X1 U9337 ( .A1(n14898), .A2(n14897), .A3(n7311), .ZN(n8127) );
  NAND3_X1 U9338 ( .A1(n14861), .A2(n14860), .A3(n7316), .ZN(n8121) );
  NAND2_X1 U9339 ( .A1(n14813), .A2(n14812), .ZN(n7397) );
  NAND2_X1 U9340 ( .A1(n14809), .A2(n14808), .ZN(n7398) );
  NAND3_X1 U9341 ( .A1(n14825), .A2(n14824), .A3(n7312), .ZN(n8124) );
  NAND2_X1 U9342 ( .A1(n14793), .A2(n14792), .ZN(n7399) );
  NAND2_X1 U9343 ( .A1(n14789), .A2(n14788), .ZN(n7400) );
  MUX2_X1 U9344 ( .A(n12956), .B(n12955), .S(n13012), .Z(n12960) );
  AOI211_X1 U9345 ( .C1(n12899), .C2(n12903), .A(n12898), .B(n12897), .ZN(
        n12901) );
  INV_X1 U9346 ( .A(n15651), .ZN(n7402) );
  NAND2_X1 U9347 ( .A1(n7402), .A2(n7401), .ZN(n7698) );
  NAND2_X1 U9348 ( .A1(n13003), .A2(n13004), .ZN(n13005) );
  NAND2_X1 U9349 ( .A1(n9949), .A2(n9950), .ZN(n15657) );
  OAI21_X1 U9350 ( .B1(n9911), .B2(n9914), .A(n7713), .ZN(n7712) );
  NAND2_X1 U9351 ( .A1(n7696), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7695) );
  NAND4_X1 U9352 ( .A1(n7782), .A2(n7783), .A3(n8012), .A4(n8168), .ZN(n8715)
         );
  NOR2_X1 U9353 ( .A1(n15606), .A2(n15605), .ZN(n9918) );
  AOI22_X1 U9354 ( .A1(n11543), .A2(n11542), .B1(n11541), .B2(n11540), .ZN(
        n15688) );
  AOI22_X1 U9355 ( .A1(n10611), .A2(n10612), .B1(n10622), .B2(n10582), .ZN(
        n10628) );
  XOR2_X1 U9356 ( .A(n13536), .B(n13533), .Z(n13522) );
  INV_X1 U9357 ( .A(n14250), .ZN(n9390) );
  NAND2_X1 U9358 ( .A1(n13613), .A2(n15712), .ZN(n7571) );
  AOI21_X1 U9359 ( .B1(n13518), .B2(n13517), .A(n13516), .ZN(n13533) );
  OR2_X1 U9360 ( .A1(n14929), .A2(n10324), .ZN(n10327) );
  OAI211_X4 U9361 ( .C1(n12641), .C2(n15079), .A(n10327), .B(n10326), .ZN(
        n14769) );
  INV_X1 U9362 ( .A(n15053), .ZN(n14770) );
  NAND2_X1 U9363 ( .A1(n11448), .A2(n13052), .ZN(n11447) );
  INV_X1 U9364 ( .A(n7755), .ZN(n13640) );
  NAND2_X1 U9365 ( .A1(n9066), .A2(n8782), .ZN(n7619) );
  OAI21_X1 U9366 ( .B1(n12723), .B2(n7968), .A(n7965), .ZN(n15294) );
  NAND2_X1 U9367 ( .A1(n7413), .A2(n14771), .ZN(n14772) );
  INV_X1 U9368 ( .A(n8102), .ZN(n10134) );
  NAND2_X1 U9369 ( .A1(n15636), .A2(n15635), .ZN(n7696) );
  NAND2_X1 U9370 ( .A1(n15667), .A2(n15668), .ZN(n7692) );
  INV_X1 U9371 ( .A(n7712), .ZN(n9860) );
  NAND2_X1 U9372 ( .A1(n7702), .A2(n7708), .ZN(n15662) );
  NAND2_X1 U9373 ( .A1(n10648), .A2(n10734), .ZN(n10647) );
  NAND2_X1 U9374 ( .A1(n12284), .A2(n7566), .ZN(n12285) );
  NOR2_X1 U9375 ( .A1(n15716), .A2(n15715), .ZN(n15714) );
  INV_X1 U9376 ( .A(n10643), .ZN(n7422) );
  XNOR2_X1 U9377 ( .A(n12280), .B(n12292), .ZN(n11549) );
  NAND2_X1 U9378 ( .A1(n14090), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n14105) );
  XNOR2_X1 U9379 ( .A(n14103), .B(n14097), .ZN(n14090) );
  AOI21_X1 U9380 ( .B1(n7421), .B2(n7420), .A(n15681), .ZN(n13583) );
  NAND2_X1 U9381 ( .A1(n13581), .A2(n13582), .ZN(n7420) );
  NOR2_X1 U9382 ( .A1(n13509), .A2(n13519), .ZN(n13529) );
  NOR2_X1 U9383 ( .A1(n13574), .A2(n13573), .ZN(n13596) );
  OAI21_X1 U9384 ( .B1(n10778), .B2(n9373), .A(n9374), .ZN(n11464) );
  AOI21_X1 U9385 ( .B1(n11194), .B2(n9377), .A(n9376), .ZN(n11377) );
  NAND2_X2 U9386 ( .A1(n9393), .A2(n9392), .ZN(n14178) );
  NAND2_X1 U9387 ( .A1(n7779), .A2(n7778), .ZN(n11448) );
  NAND2_X1 U9388 ( .A1(n7753), .A2(n12882), .ZN(n7756) );
  NAND2_X1 U9389 ( .A1(n13689), .A2(n12874), .ZN(n8696) );
  INV_X1 U9390 ( .A(n8678), .ZN(n8679) );
  INV_X1 U9391 ( .A(n13746), .ZN(n7758) );
  NAND2_X1 U9392 ( .A1(n7760), .A2(n7759), .ZN(n12493) );
  NAND2_X1 U9393 ( .A1(n13766), .A2(n13765), .ZN(n13764) );
  NAND2_X1 U9394 ( .A1(n15608), .A2(n9922), .ZN(n15612) );
  NAND2_X1 U9395 ( .A1(n15610), .A2(n15609), .ZN(n15608) );
  NAND2_X1 U9396 ( .A1(n14379), .A2(n7437), .ZN(n7436) );
  NAND2_X1 U9397 ( .A1(n14379), .A2(n7442), .ZN(n14165) );
  NAND3_X1 U9398 ( .A1(n7439), .A2(n7436), .A3(n7434), .ZN(n12867) );
  NAND2_X1 U9399 ( .A1(n11952), .A2(n7296), .ZN(n7445) );
  NAND2_X1 U9400 ( .A1(n7445), .A2(n7443), .ZN(n12476) );
  NOR2_X1 U9401 ( .A1(n9381), .A2(n12393), .ZN(n7448) );
  NAND2_X2 U9402 ( .A1(n7449), .A2(n9085), .ZN(n15840) );
  NAND2_X1 U9403 ( .A1(n7450), .A2(n9975), .ZN(P3_U3154) );
  NAND2_X1 U9404 ( .A1(n7451), .A2(n13241), .ZN(n7450) );
  NAND2_X1 U9405 ( .A1(n7452), .A2(n9967), .ZN(n7451) );
  NAND2_X1 U9406 ( .A1(n13232), .A2(n7338), .ZN(n7452) );
  NOR2_X1 U9407 ( .A1(n10971), .A2(n10970), .ZN(n11086) );
  OR2_X1 U9408 ( .A1(n13175), .A2(n13176), .ZN(n7461) );
  NAND2_X1 U9409 ( .A1(n13175), .A2(n9796), .ZN(n7457) );
  NAND3_X1 U9410 ( .A1(n7460), .A2(n9799), .A3(n7332), .ZN(n9801) );
  NAND2_X1 U9411 ( .A1(n7326), .A2(n11427), .ZN(n7462) );
  NAND2_X1 U9412 ( .A1(n7462), .A2(n7463), .ZN(n12165) );
  NAND2_X1 U9413 ( .A1(n11427), .A2(n7231), .ZN(n7475) );
  AND2_X1 U9414 ( .A1(n9760), .A2(n13480), .ZN(n7476) );
  NOR2_X1 U9415 ( .A1(n10686), .A2(n10685), .ZN(n10684) );
  AND3_X1 U9416 ( .A1(n7483), .A2(n7485), .A3(n7484), .ZN(n7783) );
  NAND3_X1 U9417 ( .A1(n7485), .A2(n8160), .A3(n8161), .ZN(n8162) );
  NOR2_X1 U9418 ( .A1(n8516), .A2(n8515), .ZN(n8520) );
  OR3_X1 U9419 ( .A1(n8516), .A2(n7493), .A3(n8515), .ZN(n8661) );
  NAND3_X1 U9420 ( .A1(n7495), .A2(n7496), .A3(n8662), .ZN(n7494) );
  NOR2_X2 U9421 ( .A1(n9986), .A2(n10046), .ZN(n10146) );
  CLKBUF_X1 U9422 ( .A(n10146), .Z(n7497) );
  NAND2_X1 U9423 ( .A1(n9987), .A2(n10146), .ZN(n11700) );
  INV_X1 U9424 ( .A(n14769), .ZN(n15775) );
  INV_X1 U9425 ( .A(n14953), .ZN(n7501) );
  NAND2_X1 U9426 ( .A1(n12637), .A2(n7505), .ZN(n7503) );
  NAND2_X1 U9427 ( .A1(n15895), .A2(n11741), .ZN(n11747) );
  NAND4_X1 U9428 ( .A1(n8221), .A2(n8223), .A3(n8222), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7646) );
  INV_X2 U9429 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8222) );
  INV_X2 U9430 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U9431 ( .A1(n11893), .A2(n11892), .ZN(n11894) );
  NAND2_X1 U9432 ( .A1(n7522), .A2(n7520), .ZN(n12444) );
  AOI21_X1 U9433 ( .B1(n7524), .B2(n7521), .A(n7308), .ZN(n7520) );
  NAND2_X1 U9434 ( .A1(n12117), .A2(n7523), .ZN(n7522) );
  AND2_X1 U9435 ( .A1(n7524), .A2(n13117), .ZN(n7523) );
  OAI21_X1 U9436 ( .B1(n12117), .B2(n7210), .A(n7523), .ZN(n13105) );
  OR2_X1 U9437 ( .A1(n12120), .A2(n7210), .ZN(n7524) );
  NAND2_X1 U9438 ( .A1(n9082), .A2(n7528), .ZN(n7526) );
  NAND2_X1 U9439 ( .A1(n11742), .A2(n7535), .ZN(n7532) );
  NAND2_X1 U9440 ( .A1(n11742), .A2(n9629), .ZN(n7541) );
  INV_X1 U9441 ( .A(n11791), .ZN(n13136) );
  OAI211_X1 U9442 ( .C1(n11742), .C2(n7536), .A(n7533), .B(n7532), .ZN(n11791)
         );
  AND2_X1 U9443 ( .A1(n7534), .A2(n7537), .ZN(n7533) );
  NOR2_X1 U9444 ( .A1(n7539), .A2(n7540), .ZN(n7538) );
  NAND2_X1 U9445 ( .A1(n8201), .A2(n7544), .ZN(n7542) );
  NAND2_X1 U9446 ( .A1(n7542), .A2(n7543), .ZN(n8205) );
  NAND2_X1 U9447 ( .A1(n7548), .A2(n7325), .ZN(n8341) );
  NAND4_X1 U9448 ( .A1(n7856), .A2(n7857), .A3(n8314), .A4(n8326), .ZN(n7548)
         );
  NAND3_X1 U9449 ( .A1(n7856), .A2(n7857), .A3(n8314), .ZN(n7549) );
  NAND2_X1 U9450 ( .A1(n7850), .A2(n7554), .ZN(n7552) );
  NAND2_X1 U9451 ( .A1(n7552), .A2(n7553), .ZN(n8197) );
  NAND2_X1 U9452 ( .A1(n8264), .A2(n8262), .ZN(n7558) );
  NAND2_X1 U9453 ( .A1(n8185), .A2(n8184), .ZN(n8367) );
  NAND2_X1 U9454 ( .A1(n13011), .A2(n13010), .ZN(n7559) );
  AND3_X2 U9455 ( .A1(n7560), .A2(n13684), .A3(n13665), .ZN(n12887) );
  NAND3_X1 U9456 ( .A1(n9014), .A2(n8933), .A3(n8047), .ZN(n7573) );
  NAND2_X2 U9457 ( .A1(n10226), .A2(n12638), .ZN(n9012) );
  NAND2_X2 U9458 ( .A1(n9400), .A2(n12489), .ZN(n10226) );
  OR2_X2 U9459 ( .A1(n10783), .A2(n10947), .ZN(n11456) );
  NOR2_X2 U9460 ( .A1(n10543), .A2(n9464), .ZN(n10542) );
  NAND2_X1 U9461 ( .A1(n7576), .A2(n9019), .ZN(n10543) );
  NOR3_X4 U9462 ( .A1(n14274), .A2(n14403), .A3(n7578), .ZN(n14209) );
  NOR2_X2 U9463 ( .A1(n12470), .A2(n14438), .ZN(n14340) );
  MUX2_X1 U9464 ( .A(n10502), .B(P2_REG1_REG_1__SCAN_IN), .S(n10272), .Z(
        n10264) );
  NAND3_X1 U9465 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n7591) );
  MUX2_X1 U9466 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n7603), .S(n15991), .Z(
        P1_U3558) );
  MUX2_X1 U9467 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n7603), .S(n15994), .Z(
        P1_U3526) );
  NAND2_X1 U9468 ( .A1(n15246), .A2(n7609), .ZN(n15171) );
  NAND3_X1 U9469 ( .A1(n7631), .A2(n7630), .A3(n7629), .ZN(n7628) );
  NAND2_X1 U9470 ( .A1(n9340), .A2(n7635), .ZN(n7633) );
  NAND2_X1 U9471 ( .A1(n9340), .A2(n9339), .ZN(n7634) );
  NAND2_X1 U9472 ( .A1(n9300), .A2(n7640), .ZN(n7639) );
  NAND2_X2 U9473 ( .A1(n7645), .A2(n7646), .ZN(n8763) );
  NAND3_X1 U9474 ( .A1(n8224), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7647) );
  NAND3_X1 U9475 ( .A1(n8223), .A2(n8221), .A3(n8222), .ZN(n7648) );
  NAND2_X1 U9476 ( .A1(n8838), .A2(n7653), .ZN(n7651) );
  OAI21_X1 U9477 ( .B1(n12515), .B2(n7662), .A(n7660), .ZN(n12532) );
  NAND2_X1 U9478 ( .A1(n7659), .A2(n7658), .ZN(n8482) );
  NAND2_X1 U9479 ( .A1(n12515), .A2(n7660), .ZN(n7659) );
  OAI21_X1 U9480 ( .B1(n12515), .B2(n13065), .A(n8453), .ZN(n12491) );
  NAND2_X1 U9481 ( .A1(n13826), .A2(n7682), .ZN(n13811) );
  NAND2_X1 U9482 ( .A1(n7684), .A2(n7683), .ZN(n11444) );
  NAND2_X1 U9483 ( .A1(n11249), .A2(n7315), .ZN(n11496) );
  INV_X1 U9484 ( .A(n8715), .ZN(n7687) );
  NAND2_X1 U9485 ( .A1(n7687), .A2(n7686), .ZN(n8170) );
  NAND2_X1 U9486 ( .A1(n7687), .A2(n7685), .ZN(n13967) );
  NAND2_X1 U9487 ( .A1(n15642), .A2(n15643), .ZN(n15641) );
  INV_X1 U9488 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7690) );
  OR2_X1 U9489 ( .A1(n15661), .A2(n7709), .ZN(n7702) );
  OR2_X1 U9490 ( .A1(n7239), .A2(n15663), .ZN(n7708) );
  INV_X1 U9491 ( .A(n7711), .ZN(n15659) );
  INV_X1 U9492 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7710) );
  OAI211_X1 U9493 ( .C1(n10656), .C2(n7722), .A(n7721), .B(n7719), .ZN(n10600)
         );
  NAND2_X1 U9494 ( .A1(n7727), .A2(n7726), .ZN(n10614) );
  NAND3_X1 U9495 ( .A1(n7729), .A2(n10644), .A3(P3_REG1_REG_5__SCAN_IN), .ZN(
        n10796) );
  NAND2_X1 U9496 ( .A1(n7728), .A2(n11810), .ZN(n10795) );
  INV_X1 U9497 ( .A(n7735), .ZN(n7734) );
  NAND2_X1 U9498 ( .A1(n13571), .A2(n7352), .ZN(n7738) );
  OAI211_X1 U9499 ( .C1(n13571), .C2(n7740), .A(n7738), .B(n7737), .ZN(n13614)
         );
  NOR2_X1 U9500 ( .A1(n13571), .A2(n13572), .ZN(n13574) );
  NAND3_X1 U9501 ( .A1(n7745), .A2(n7746), .A3(n9748), .ZN(n12902) );
  NAND2_X1 U9502 ( .A1(n13647), .A2(n7560), .ZN(n7753) );
  NAND2_X1 U9503 ( .A1(n7747), .A2(n7748), .ZN(n13047) );
  NOR2_X2 U9504 ( .A1(n13049), .A2(n13042), .ZN(n7757) );
  AOI21_X2 U9505 ( .B1(n13748), .B2(n8694), .A(n7230), .ZN(n13862) );
  NAND2_X1 U9506 ( .A1(n12550), .A2(n7762), .ZN(n7760) );
  NAND2_X1 U9507 ( .A1(n11502), .A2(n7767), .ZN(n7764) );
  NAND2_X1 U9508 ( .A1(n7764), .A2(n7765), .ZN(n11827) );
  OAI22_X1 U9509 ( .A1(n12534), .A2(n7770), .B1(n8139), .B2(n7772), .ZN(n13766) );
  INV_X1 U9510 ( .A(n8139), .ZN(n7777) );
  NAND2_X1 U9511 ( .A1(n11147), .A2(n13057), .ZN(n7779) );
  INV_X1 U9512 ( .A(n12904), .ZN(n7778) );
  NAND2_X1 U9513 ( .A1(n7781), .A2(n13083), .ZN(n7780) );
  XNOR2_X1 U9514 ( .A(n13048), .B(n13610), .ZN(n7781) );
  NOR2_X1 U9515 ( .A1(n8251), .A2(n8162), .ZN(n8438) );
  NOR2_X1 U9517 ( .A1(n13047), .A2(n13046), .ZN(n13048) );
  NAND2_X1 U9518 ( .A1(n11827), .A2(n12929), .ZN(n11928) );
  NAND2_X1 U9519 ( .A1(n8679), .A2(n8148), .ZN(n11223) );
  NAND2_X1 U9520 ( .A1(n8696), .A2(n12886), .ZN(n13686) );
  XNOR2_X2 U9521 ( .A(n8298), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10595) );
  OAI21_X1 U9522 ( .B1(n8677), .B2(n13831), .A(n8676), .ZN(n13622) );
  INV_X1 U9523 ( .A(n13630), .ZN(n13633) );
  NAND2_X1 U9524 ( .A1(n13633), .A2(n13632), .ZN(n13637) );
  NAND2_X1 U9525 ( .A1(n14727), .A2(n14728), .ZN(n14726) );
  NAND3_X1 U9526 ( .A1(n7791), .A2(n7790), .A3(n7787), .ZN(n14639) );
  NAND2_X1 U9527 ( .A1(n14727), .A2(n7306), .ZN(n7790) );
  OR2_X1 U9528 ( .A1(n14727), .A2(n7792), .ZN(n7791) );
  NAND2_X1 U9529 ( .A1(n11910), .A2(n11911), .ZN(n12228) );
  INV_X1 U9530 ( .A(n7807), .ZN(n14595) );
  OAI21_X1 U9531 ( .B1(n12274), .B2(n7817), .A(n7815), .ZN(n7822) );
  NAND2_X1 U9532 ( .A1(n7828), .A2(n11291), .ZN(n7827) );
  NAND2_X1 U9533 ( .A1(n7827), .A2(n7829), .ZN(n11646) );
  NAND2_X1 U9534 ( .A1(n7838), .A2(n8197), .ZN(n8454) );
  NAND2_X1 U9535 ( .A1(n8437), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7838) );
  AOI21_X1 U9536 ( .B1(n8197), .B2(n7841), .A(n7840), .ZN(n7839) );
  INV_X1 U9537 ( .A(n8455), .ZN(n7840) );
  INV_X1 U9538 ( .A(n8197), .ZN(n7842) );
  INV_X1 U9539 ( .A(n8299), .ZN(n7855) );
  NAND2_X1 U9540 ( .A1(n7855), .A2(n8179), .ZN(n7856) );
  NAND2_X1 U9541 ( .A1(n8178), .A2(n7256), .ZN(n7857) );
  NAND2_X1 U9542 ( .A1(n7858), .A2(n8179), .ZN(n8315) );
  NAND2_X1 U9543 ( .A1(n8300), .A2(n8299), .ZN(n7858) );
  NAND2_X1 U9544 ( .A1(n8621), .A2(n8622), .ZN(n7861) );
  NAND2_X1 U9545 ( .A1(n8621), .A2(n7862), .ZN(n7860) );
  NAND2_X1 U9546 ( .A1(n11083), .A2(n7323), .ZN(n10851) );
  NAND2_X1 U9547 ( .A1(n10024), .A2(n11076), .ZN(n11083) );
  AOI21_X1 U9548 ( .B1(n10958), .B2(n11009), .A(n7298), .ZN(n7876) );
  NAND2_X1 U9549 ( .A1(n14042), .A2(n7884), .ZN(n7880) );
  NAND2_X1 U9550 ( .A1(n7880), .A2(n7881), .ZN(n12839) );
  AND2_X1 U9551 ( .A1(n11868), .A2(n9722), .ZN(n7891) );
  OAI211_X1 U9552 ( .C1(n10226), .C2(n10272), .A(n8990), .B(n8991), .ZN(n9001)
         );
  NAND2_X1 U9553 ( .A1(n8067), .A2(n8132), .ZN(n8876) );
  NAND2_X1 U9554 ( .A1(n14206), .A2(n7205), .ZN(n7905) );
  INV_X1 U9555 ( .A(n9312), .ZN(n7909) );
  NAND2_X1 U9556 ( .A1(n14206), .A2(n14205), .ZN(n14204) );
  NAND3_X1 U9557 ( .A1(n11508), .A2(n7237), .A3(n7211), .ZN(n7912) );
  NAND3_X1 U9558 ( .A1(n7918), .A2(n7240), .A3(n7916), .ZN(n12050) );
  NAND2_X1 U9559 ( .A1(n14178), .A2(n7301), .ZN(n7920) );
  NAND2_X1 U9560 ( .A1(n14178), .A2(n14177), .ZN(n7929) );
  OAI211_X1 U9561 ( .C1(n14178), .C2(n7924), .A(n7921), .B(n7920), .ZN(n9405)
         );
  AOI21_X1 U9562 ( .B1(n9212), .B2(n10377), .A(n7931), .ZN(n7930) );
  NAND2_X1 U9563 ( .A1(n11339), .A2(n7203), .ZN(n7935) );
  NAND2_X1 U9564 ( .A1(n9384), .A2(n7939), .ZN(n7938) );
  NAND2_X1 U9565 ( .A1(n7947), .A2(n7949), .ZN(n9387) );
  INV_X1 U9566 ( .A(n7953), .ZN(n14297) );
  NAND3_X1 U9567 ( .A1(n8067), .A2(n8132), .A3(n8877), .ZN(n7954) );
  NOR2_X2 U9568 ( .A1(n11121), .A2(n9982), .ZN(n9987) );
  NAND4_X1 U9569 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), .ZN(n11121)
         );
  NAND2_X1 U9570 ( .A1(n7955), .A2(n7956), .ZN(n12028) );
  NAND2_X1 U9571 ( .A1(n11964), .A2(n11970), .ZN(n7955) );
  NAND2_X1 U9572 ( .A1(n10821), .A2(n7960), .ZN(n7959) );
  INV_X1 U9573 ( .A(n15343), .ZN(n7974) );
  NAND2_X1 U9574 ( .A1(n7976), .A2(n7309), .ZN(n11717) );
  INV_X1 U9575 ( .A(n7984), .ZN(n15237) );
  INV_X1 U9576 ( .A(n12244), .ZN(n7994) );
  NAND3_X1 U9577 ( .A1(n7241), .A2(n13205), .A3(n7331), .ZN(n7999) );
  NAND3_X1 U9578 ( .A1(n7999), .A2(n7998), .A3(n9805), .ZN(n13182) );
  NAND2_X1 U9579 ( .A1(n13205), .A2(n13690), .ZN(n7998) );
  AND2_X1 U9580 ( .A1(n13205), .A2(n13727), .ZN(n8000) );
  INV_X1 U9581 ( .A(n9743), .ZN(n9744) );
  NAND3_X1 U9582 ( .A1(n8717), .A2(n8718), .A3(n8716), .ZN(n8002) );
  NOR2_X2 U9583 ( .A1(n8147), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8012) );
  NAND4_X1 U9584 ( .A1(n15033), .A2(n15032), .A3(n8014), .A4(n8013), .ZN(
        P1_U3242) );
  OAI21_X2 U9585 ( .B1(n8973), .B2(n8016), .A(n8791), .ZN(n9112) );
  NAND2_X1 U9586 ( .A1(n8807), .A2(n8036), .ZN(n8032) );
  NAND2_X1 U9587 ( .A1(n8795), .A2(n7305), .ZN(n8038) );
  NAND2_X1 U9588 ( .A1(n8795), .A2(n8794), .ZN(n9128) );
  NAND3_X1 U9589 ( .A1(n8046), .A2(n8045), .A3(n8759), .ZN(n10318) );
  MUX2_X1 U9590 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9030), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9031) );
  NOR2_X1 U9591 ( .A1(n8049), .A2(n7264), .ZN(n8048) );
  NAND2_X1 U9592 ( .A1(n8993), .A2(n8992), .ZN(n8049) );
  NAND2_X1 U9593 ( .A1(n9716), .A2(n8056), .ZN(n8052) );
  AND2_X1 U9594 ( .A1(n9721), .A2(n11862), .ZN(n8061) );
  NAND2_X1 U9595 ( .A1(n8068), .A2(n8071), .ZN(n9488) );
  NAND3_X1 U9596 ( .A1(n9480), .A2(n9481), .A3(n8069), .ZN(n8068) );
  AOI21_X1 U9597 ( .B1(n9547), .B2(n9546), .A(n9544), .ZN(n9545) );
  NAND2_X1 U9598 ( .A1(n8074), .A2(n8075), .ZN(n9510) );
  NAND2_X1 U9599 ( .A1(n8079), .A2(n8080), .ZN(n9588) );
  INV_X1 U9600 ( .A(n9582), .ZN(n8081) );
  INV_X1 U9601 ( .A(n9493), .ZN(n8085) );
  INV_X1 U9602 ( .A(n9492), .ZN(n8086) );
  NAND2_X1 U9603 ( .A1(n8087), .A2(n8088), .ZN(n9533) );
  NAND3_X1 U9604 ( .A1(n9522), .A2(n7320), .A3(n9521), .ZN(n8087) );
  INV_X1 U9605 ( .A(n9525), .ZN(n8089) );
  NAND2_X1 U9606 ( .A1(n11695), .A2(n10828), .ZN(n8091) );
  NAND2_X1 U9607 ( .A1(n12210), .A2(n12209), .ZN(n8096) );
  NAND2_X1 U9608 ( .A1(n8096), .A2(n7307), .ZN(n12329) );
  NAND2_X1 U9609 ( .A1(n11653), .A2(n11654), .ZN(n8099) );
  NAND2_X1 U9610 ( .A1(n8099), .A2(n8097), .ZN(n11623) );
  NAND2_X1 U9611 ( .A1(n12607), .A2(n7302), .ZN(n15305) );
  INV_X1 U9612 ( .A(n8102), .ZN(n8101) );
  NAND2_X1 U9613 ( .A1(n8101), .A2(n10116), .ZN(n8100) );
  NAND2_X1 U9614 ( .A1(n14988), .A2(n14757), .ZN(n8109) );
  NAND2_X1 U9615 ( .A1(n14755), .A2(n15140), .ZN(n8110) );
  INV_X1 U9616 ( .A(n15140), .ZN(n10342) );
  INV_X1 U9617 ( .A(n14755), .ZN(n10343) );
  NAND2_X1 U9618 ( .A1(n8124), .A2(n8125), .ZN(n14831) );
  NAND3_X1 U9619 ( .A1(n14804), .A2(n14803), .A3(n7275), .ZN(n8129) );
  NAND2_X1 U9620 ( .A1(n8129), .A2(n8130), .ZN(n14810) );
  NAND2_X1 U9621 ( .A1(n15384), .A2(n15383), .ZN(n15458) );
  XNOR2_X1 U9622 ( .A(n8635), .B(n8634), .ZN(n12870) );
  AND2_X1 U9623 ( .A1(n8982), .A2(n8981), .ZN(n8134) );
  NAND2_X1 U9624 ( .A1(n9410), .A2(n8151), .ZN(n9855) );
  NAND2_X1 U9625 ( .A1(n10525), .A2(n10527), .ZN(n10526) );
  NAND2_X1 U9626 ( .A1(n9126), .A2(n7259), .ZN(n11508) );
  NAND2_X1 U9627 ( .A1(n8666), .A2(n8738), .ZN(n12899) );
  AND2_X1 U9628 ( .A1(n9676), .A2(n8140), .ZN(n9698) );
  AND2_X1 U9629 ( .A1(n10505), .A2(n10515), .ZN(n9838) );
  OAI211_X1 U9630 ( .C1(n9463), .C2(n9462), .A(n9461), .B(n9460), .ZN(n9474)
         );
  OAI222_X1 U9631 ( .A1(n14477), .A2(n14930), .B1(P2_U3088), .B2(n13152), .C1(
        n13151), .C2(n13150), .ZN(P2_U3297) );
  OAI21_X1 U9632 ( .B1(n15313), .B2(n7189), .A(n12618), .ZN(n15290) );
  NAND4_X4 U9633 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n15052) );
  OR2_X1 U9634 ( .A1(n7189), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10331) );
  INV_X1 U9635 ( .A(n14359), .ZN(n14311) );
  AND2_X2 U9636 ( .A1(n11185), .A2(n14308), .ZN(n14359) );
  AND2_X1 U9637 ( .A1(n13638), .A2(n13218), .ZN(n8133) );
  INV_X1 U9638 ( .A(n16000), .ZN(n16008) );
  INV_X2 U9639 ( .A(n15810), .ZN(n15802) );
  XNOR2_X1 U9640 ( .A(n8711), .B(P3_IR_REG_25__SCAN_IN), .ZN(n8736) );
  AND4_X1 U9641 ( .A1(n8452), .A2(n8451), .A3(n8450), .A4(n8449), .ZN(n12957)
         );
  INV_X1 U9642 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10754) );
  AND2_X1 U9643 ( .A1(n10133), .A2(n10136), .ZN(n8135) );
  INV_X1 U9644 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10136) );
  AND2_X1 U9645 ( .A1(n15857), .A2(n14075), .ZN(n8136) );
  AND2_X1 U9646 ( .A1(n9473), .A2(n9472), .ZN(n8137) );
  OR2_X1 U9647 ( .A1(n15398), .A2(n15241), .ZN(n8138) );
  NOR2_X1 U9648 ( .A1(n8691), .A2(n13778), .ZN(n8139) );
  AND2_X1 U9649 ( .A1(n9675), .A2(n9674), .ZN(n8140) );
  AND4_X1 U9650 ( .A1(n8343), .A2(n8158), .A3(n8347), .A4(n8363), .ZN(n8141)
         );
  OR2_X1 U9651 ( .A1(n14937), .A2(n7409), .ZN(n15345) );
  OR2_X1 U9652 ( .A1(n13925), .A2(n13662), .ZN(n8142) );
  OR2_X1 U9653 ( .A1(n10226), .A2(n10260), .ZN(n8145) );
  AND2_X1 U9654 ( .A1(n8804), .A2(n8803), .ZN(n8146) );
  NAND4_X1 U9655 ( .A1(n8166), .A2(n8165), .A3(n8164), .A4(n8513), .ZN(n8147)
         );
  INV_X1 U9656 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12162) );
  INV_X1 U9657 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12682) );
  INV_X1 U9658 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12389) );
  INV_X1 U9659 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12670) );
  INV_X1 U9660 ( .A(n14403), .ZN(n9407) );
  INV_X1 U9661 ( .A(n14067), .ZN(n9224) );
  INV_X1 U9662 ( .A(n15841), .ZN(n15903) );
  NAND2_X1 U9663 ( .A1(n9236), .A2(n9235), .ZN(n14066) );
  INV_X1 U9664 ( .A(n12999), .ZN(n13719) );
  AND2_X1 U9665 ( .A1(n12896), .A2(n12895), .ZN(n8148) );
  INV_X1 U9666 ( .A(n12818), .ZN(n11779) );
  INV_X1 U9667 ( .A(n14063), .ZN(n14019) );
  NAND2_X1 U9668 ( .A1(n9327), .A2(n9326), .ZN(n14063) );
  NAND2_X1 U9669 ( .A1(n9854), .A2(n9853), .ZN(n15908) );
  OR2_X1 U9670 ( .A1(n14922), .A2(n14921), .ZN(n8150) );
  AND2_X1 U9671 ( .A1(n12869), .A2(n9409), .ZN(n8151) );
  INV_X1 U9672 ( .A(n14386), .ZN(n14194) );
  OR2_X1 U9673 ( .A1(n9547), .A2(n9546), .ZN(n8152) );
  NAND2_X1 U9674 ( .A1(n9529), .A2(n11403), .ZN(n9448) );
  NAND2_X1 U9675 ( .A1(n9449), .A2(n9448), .ZN(n9451) );
  OAI21_X1 U9676 ( .B1(n9454), .B2(n11403), .A(n9453), .ZN(n9457) );
  OR2_X1 U9677 ( .A1(n9455), .A2(n9456), .ZN(n9473) );
  AOI21_X1 U9678 ( .B1(n9470), .B2(n9474), .A(n9469), .ZN(n9480) );
  OAI21_X1 U9679 ( .B1(n11064), .B2(n9529), .A(n9478), .ZN(n9479) );
  INV_X1 U9680 ( .A(n14806), .ZN(n14807) );
  OAI21_X1 U9681 ( .B1(n12852), .B2(n9529), .A(n9503), .ZN(n9504) );
  OAI21_X1 U9682 ( .B1(n12851), .B2(n9529), .A(n9514), .ZN(n9515) );
  NAND2_X1 U9683 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  INV_X1 U9684 ( .A(n9534), .ZN(n9535) );
  INV_X1 U9685 ( .A(n12893), .ZN(n12914) );
  INV_X1 U9686 ( .A(n12888), .ZN(n12889) );
  INV_X1 U9687 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U9688 ( .A1(n13016), .A2(n13002), .ZN(n13017) );
  INV_X1 U9689 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13344) );
  INV_X1 U9690 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10131) );
  NOR2_X1 U9691 ( .A1(n8590), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8577) );
  INV_X1 U9692 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13379) );
  NOR2_X1 U9693 ( .A1(n8506), .A2(n8155), .ZN(n8505) );
  NOR2_X1 U9694 ( .A1(n8447), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8446) );
  INV_X1 U9695 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8169) );
  INV_X1 U9696 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8383) );
  NOR2_X1 U9697 ( .A1(n9304), .A2(n14020), .ZN(n9303) );
  INV_X1 U9698 ( .A(n9174), .ZN(n8888) );
  NAND2_X1 U9699 ( .A1(n9005), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8981) );
  INV_X1 U9700 ( .A(n9643), .ZN(n9028) );
  INV_X1 U9701 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11976) );
  AND2_X1 U9702 ( .A1(n12659), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n12674) );
  INV_X1 U9703 ( .A(n15250), .ZN(n12667) );
  INV_X1 U9704 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11749) );
  INV_X1 U9705 ( .A(n12957), .ZN(n9776) );
  INV_X1 U9706 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U9707 ( .A1(n8524), .A2(n13446), .ZN(n8557) );
  INV_X1 U9708 ( .A(n9763), .ZN(n9764) );
  OR2_X1 U9709 ( .A1(n8229), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8653) );
  AOI21_X1 U9710 ( .B1(n13631), .B2(n7752), .A(n13831), .ZN(n13632) );
  OAI22_X1 U9711 ( .A1(n13692), .A2(n8620), .B1(n13699), .B2(n13708), .ZN(
        n13671) );
  OR2_X1 U9712 ( .A1(n8430), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8447) );
  NOR2_X1 U9713 ( .A1(n13625), .A2(n13905), .ZN(n8755) );
  INV_X1 U9714 ( .A(n9838), .ZN(n9841) );
  AND2_X1 U9715 ( .A1(n12146), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8210) );
  INV_X1 U9716 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8519) );
  INV_X1 U9717 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8188) );
  INV_X1 U9718 ( .A(n10035), .ZN(n10033) );
  NAND2_X1 U9719 ( .A1(n9303), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9320) );
  OR2_X1 U9720 ( .A1(n9290), .A2(n14029), .ZN(n9304) );
  OR2_X1 U9721 ( .A1(n9243), .A2(n8890), .ZN(n9260) );
  NAND2_X1 U9722 ( .A1(n8888), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9192) );
  AND2_X1 U9723 ( .A1(n14396), .A2(n14018), .ZN(n9391) );
  INV_X1 U9724 ( .A(n14243), .ZN(n14254) );
  INV_X1 U9725 ( .A(n14444), .ZN(n9406) );
  AND2_X1 U9726 ( .A1(n11288), .A2(n11287), .ZN(n11289) );
  INV_X1 U9727 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U9728 ( .A1(n12644), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12643) );
  NAND2_X1 U9729 ( .A1(n12667), .A2(n15036), .ZN(n12668) );
  NAND2_X1 U9730 ( .A1(n10748), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12660) );
  OR2_X1 U9731 ( .A1(n11750), .A2(n11749), .ZN(n11977) );
  INV_X1 U9732 ( .A(n15928), .ZN(n11969) );
  INV_X1 U9733 ( .A(SI_22_), .ZN(n9252) );
  AND2_X1 U9734 ( .A1(n8815), .A2(n8814), .ZN(n8938) );
  INV_X1 U9735 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9983) );
  INV_X1 U9736 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U9737 ( .A1(n9775), .A2(n9776), .ZN(n9777) );
  NOR2_X1 U9738 ( .A1(n8357), .A2(n8153), .ZN(n8242) );
  OR2_X1 U9739 ( .A1(n8626), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8638) );
  AND2_X1 U9740 ( .A1(n8242), .A2(n8154), .ZN(n8373) );
  NAND2_X1 U9741 ( .A1(n9764), .A2(n13479), .ZN(n9765) );
  OR2_X1 U9742 ( .A1(n9843), .A2(n9842), .ZN(n13236) );
  INV_X1 U9743 ( .A(n10505), .ZN(n8541) );
  AND4_X1 U9744 ( .A1(n8415), .A2(n8414), .A3(n8413), .A4(n8412), .ZN(n12552)
         );
  INV_X1 U9745 ( .A(n13635), .ZN(n13636) );
  OR2_X1 U9746 ( .A1(n16000), .A2(n9738), .ZN(n9739) );
  AND2_X1 U9747 ( .A1(n12989), .A2(n12988), .ZN(n13765) );
  AND2_X1 U9748 ( .A1(n12948), .A2(n12953), .ZN(n12549) );
  INV_X1 U9749 ( .A(n8680), .ZN(n13052) );
  INV_X1 U9750 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8539) );
  AND2_X1 U9751 ( .A1(n8387), .A2(n8386), .ZN(n8403) );
  INV_X1 U9752 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10963) );
  OR2_X1 U9753 ( .A1(n9192), .A2(n9191), .ZN(n9217) );
  INV_X1 U9754 ( .A(n12145), .ZN(n9726) );
  INV_X1 U9755 ( .A(n10243), .ZN(n10242) );
  AND2_X1 U9756 ( .A1(n10242), .A2(n12512), .ZN(n10237) );
  INV_X1 U9757 ( .A(n14062), .ZN(n13988) );
  INV_X1 U9758 ( .A(n14064), .ZN(n14018) );
  INV_X1 U9759 ( .A(n11956), .ZN(n12401) );
  OR2_X1 U9760 ( .A1(n9437), .A2(n9400), .ZN(n14320) );
  INV_X1 U9761 ( .A(n9708), .ZN(n14258) );
  INV_X1 U9762 ( .A(n12797), .ZN(n15904) );
  AND2_X1 U9763 ( .A1(n12161), .A2(n9426), .ZN(n9430) );
  INV_X1 U9764 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9358) );
  OR2_X1 U9765 ( .A1(n12183), .A2(n12182), .ZN(n12215) );
  AND2_X1 U9766 ( .A1(n14692), .A2(n14691), .ZN(n14532) );
  AND2_X1 U9767 ( .A1(n14640), .A2(n14641), .ZN(n14540) );
  NAND2_X1 U9768 ( .A1(n10935), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14746) );
  OR2_X1 U9769 ( .A1(n7189), .A2(n15229), .ZN(n12678) );
  AND2_X1 U9770 ( .A1(n12612), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n12625) );
  INV_X1 U9771 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10392) );
  OR2_X1 U9772 ( .A1(n11164), .A2(n11163), .ZN(n11161) );
  INV_X1 U9773 ( .A(n14975), .ZN(n12710) );
  INV_X1 U9774 ( .A(n15262), .ZN(n12728) );
  INV_X1 U9775 ( .A(n14966), .ZN(n12029) );
  INV_X1 U9776 ( .A(n15947), .ZN(n15317) );
  OAI21_X1 U9777 ( .B1(n10295), .B2(P1_D_REG_0__SCAN_IN), .A(n15474), .ZN(
        n11258) );
  OR2_X1 U9778 ( .A1(n14937), .A2(n15072), .ZN(n15195) );
  INV_X1 U9779 ( .A(n10280), .ZN(n10282) );
  AND2_X1 U9780 ( .A1(n9341), .A2(n8865), .ZN(n9339) );
  AND2_X1 U9781 ( .A1(n8837), .A2(n8836), .ZN(n9226) );
  AND2_X1 U9782 ( .A1(n8819), .A2(n8818), .ZN(n8927) );
  AOI21_X1 U9783 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n9888), .A(n9887), .ZN(
        n9895) );
  INV_X1 U9784 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n13329) );
  INV_X1 U9785 ( .A(n13236), .ZN(n13245) );
  AND2_X1 U9786 ( .A1(n9849), .A2(n9848), .ZN(n13218) );
  AND2_X1 U9787 ( .A1(n8235), .A2(n8234), .ZN(n13663) );
  AND4_X1 U9788 ( .A1(n8480), .A2(n8479), .A3(n8478), .A4(n8477), .ZN(n13832)
         );
  INV_X1 U9789 ( .A(n12552), .ZN(n13266) );
  INV_X1 U9790 ( .A(n15718), .ZN(n15675) );
  INV_X1 U9791 ( .A(n15677), .ZN(n15711) );
  INV_X1 U9792 ( .A(n13611), .ZN(n15704) );
  NAND2_X1 U9793 ( .A1(n10898), .A2(n10897), .ZN(n15804) );
  AND2_X1 U9794 ( .A1(n15810), .A2(n15800), .ZN(n13820) );
  AND3_X1 U9795 ( .A1(n8268), .A2(n8267), .A3(n8266), .ZN(n11836) );
  OR2_X1 U9796 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  OR2_X1 U9797 ( .A1(n15769), .A2(n15889), .ZN(n15917) );
  NAND2_X1 U9798 ( .A1(n8705), .A2(n8745), .ZN(n15769) );
  INV_X1 U9799 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8662) );
  NOR2_X1 U9800 ( .A1(n8388), .A2(n8403), .ZN(n11541) );
  INV_X1 U9801 ( .A(n14050), .ZN(n13142) );
  OR2_X1 U9802 ( .A1(n14002), .A2(n14322), .ZN(n14050) );
  OR2_X1 U9803 ( .A1(n14045), .A2(n9321), .ZN(n9327) );
  INV_X1 U9804 ( .A(n14148), .ZN(n15598) );
  AND2_X1 U9805 ( .A1(n10237), .A2(n10238), .ZN(n15583) );
  INV_X1 U9806 ( .A(n12836), .ZN(n14167) );
  NAND2_X1 U9807 ( .A1(n9283), .A2(n9282), .ZN(n14252) );
  INV_X1 U9808 ( .A(n14320), .ZN(n14353) );
  INV_X1 U9809 ( .A(n14308), .ZN(n14345) );
  NAND2_X1 U9810 ( .A1(n14231), .A2(n11175), .ZN(n14292) );
  INV_X1 U9811 ( .A(n15860), .ZN(n14442) );
  AND3_X1 U9812 ( .A1(n10006), .A2(n9439), .A3(n15519), .ZN(n9854) );
  AND2_X1 U9813 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10016), .ZN(n9436) );
  INV_X1 U9814 ( .A(n14753), .ZN(n14716) );
  INV_X1 U9815 ( .A(n14943), .ZN(n15151) );
  AND4_X1 U9816 ( .A1(n12585), .A2(n12584), .A3(n12583), .A4(n12582), .ZN(
        n14734) );
  AND2_X1 U9817 ( .A1(n12634), .A2(n12633), .ZN(n14705) );
  AND4_X1 U9818 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n14748) );
  AND4_X1 U9819 ( .A1(n11608), .A2(n11607), .A3(n11606), .A4(n11605), .ZN(
        n12269) );
  INV_X1 U9820 ( .A(n15135), .ZN(n15739) );
  INV_X1 U9821 ( .A(n15087), .ZN(n15730) );
  AND2_X1 U9822 ( .A1(n10176), .A2(n7409), .ZN(n15741) );
  OAI21_X1 U9823 ( .B1(n14734), .B2(n15345), .A(n12716), .ZN(n12717) );
  INV_X1 U9824 ( .A(n15345), .ZN(n15289) );
  AND2_X1 U9825 ( .A1(n14628), .A2(n10344), .ZN(n11566) );
  INV_X1 U9826 ( .A(n15981), .ZN(n15970) );
  INV_X1 U9827 ( .A(n15988), .ZN(n15959) );
  INV_X1 U9828 ( .A(n11328), .ZN(n15880) );
  AND3_X1 U9829 ( .A1(n10482), .A2(n10472), .A3(n11259), .ZN(n10367) );
  NAND2_X1 U9830 ( .A1(n10293), .A2(n10119), .ZN(n15471) );
  INV_X1 U9831 ( .A(n9919), .ZN(n9920) );
  AND2_X1 U9832 ( .A1(n10511), .A2(n10510), .ZN(n15702) );
  NOR2_X1 U9833 ( .A1(n9850), .A2(n8133), .ZN(n9851) );
  NAND2_X1 U9834 ( .A1(n9828), .A2(n10898), .ZN(n13222) );
  INV_X1 U9835 ( .A(n13250), .ZN(n13200) );
  AND2_X1 U9836 ( .A1(n13037), .A2(n8658), .ZN(n13634) );
  INV_X1 U9837 ( .A(n13800), .ZN(n13760) );
  INV_X1 U9838 ( .A(n12380), .ZN(n13264) );
  INV_X1 U9839 ( .A(n15712), .ZN(n15681) );
  OR2_X1 U9840 ( .A1(n10516), .A2(n10515), .ZN(n15677) );
  OR2_X1 U9841 ( .A1(n10516), .A2(n10977), .ZN(n15718) );
  NOR2_X1 U9842 ( .A1(n8755), .A2(n8757), .ZN(n8758) );
  INV_X1 U9843 ( .A(n15997), .ZN(n16004) );
  AND2_X2 U9844 ( .A1(n10895), .A2(n8753), .ZN(n15997) );
  INV_X1 U9845 ( .A(n13683), .ZN(n13925) );
  INV_X1 U9846 ( .A(n12519), .ZN(n12531) );
  AND3_X1 U9847 ( .A1(n15869), .A2(n15868), .A3(n15867), .ZN(n15871) );
  AND2_X2 U9848 ( .A1(n9737), .A2(n10898), .ZN(n16000) );
  OR2_X1 U9849 ( .A1(n8722), .A2(n13964), .ZN(n12578) );
  AND2_X1 U9850 ( .A1(n8725), .A2(n8724), .ZN(n13965) );
  INV_X1 U9851 ( .A(SI_16_), .ZN(n13409) );
  INV_X1 U9852 ( .A(SI_11_), .ZN(n13419) );
  INV_X1 U9853 ( .A(n14035), .ZN(n14044) );
  NAND2_X1 U9854 ( .A1(n8912), .A2(n8911), .ZN(n14062) );
  NAND2_X1 U9855 ( .A1(n9297), .A2(n9296), .ZN(n14064) );
  INV_X1 U9856 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10152) );
  OR2_X1 U9857 ( .A1(n15575), .A2(P2_U3088), .ZN(n14148) );
  INV_X1 U9858 ( .A(n15522), .ZN(n15601) );
  INV_X1 U9859 ( .A(n14292), .ZN(n14364) );
  INV_X1 U9860 ( .A(n14311), .ZN(n14347) );
  NAND2_X1 U9861 ( .A1(n15909), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9442) );
  INV_X2 U9862 ( .A(n15909), .ZN(n14469) );
  NAND2_X1 U9863 ( .A1(n9854), .A2(n15525), .ZN(n15909) );
  OR2_X1 U9864 ( .A1(n15523), .A2(n15520), .ZN(n15521) );
  INV_X1 U9865 ( .A(n14104), .ZN(n14097) );
  INV_X1 U9866 ( .A(n15922), .ZN(n11920) );
  OR2_X1 U9867 ( .A1(n10483), .A2(n10476), .ZN(n14753) );
  INV_X1 U9868 ( .A(n14734), .ZN(n15217) );
  OAI21_X1 U9869 ( .B1(n15329), .B2(n7189), .A(n12605), .ZN(n15343) );
  INV_X1 U9870 ( .A(n11564), .ZN(n15049) );
  OR2_X1 U9871 ( .A1(n10179), .A2(n15149), .ZN(n15135) );
  OR2_X1 U9872 ( .A1(n10180), .A2(n7409), .ZN(n15087) );
  NAND2_X1 U9873 ( .A1(n15760), .A2(n11566), .ZN(n15285) );
  AND2_X2 U9874 ( .A1(n10367), .A2(n10296), .ZN(n15991) );
  OR2_X1 U9875 ( .A1(n15441), .A2(n15440), .ZN(n15468) );
  AND2_X1 U9876 ( .A1(n15925), .A2(n15924), .ZN(n15927) );
  INV_X1 U9877 ( .A(n15994), .ZN(n15992) );
  NOR2_X1 U9878 ( .A1(n15472), .A2(n15471), .ZN(n15502) );
  CLKBUF_X1 U9879 ( .A(n15502), .Z(n15517) );
  INV_X1 U9880 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n11411) );
  INV_X1 U9881 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10422) );
  INV_X2 U9882 ( .A(n13265), .ZN(P3_U3897) );
  OAI21_X1 U9883 ( .B1(n9742), .B2(n16004), .A(n8758), .ZN(P3_U3488) );
  OAI21_X1 U9884 ( .B1(n9742), .B2(n16008), .A(n9741), .ZN(P3_U3456) );
  AND2_X1 U9885 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10223), .ZN(P2_U3947) );
  XNOR2_X1 U9886 ( .A(n9964), .B(n9963), .ZN(SUB_1596_U4) );
  NOR2_X1 U9887 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8319) );
  INV_X1 U9888 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10794) );
  NAND2_X1 U9889 ( .A1(n8319), .A2(n10794), .ZN(n8355) );
  NAND2_X1 U9890 ( .A1(n13454), .A2(n13329), .ZN(n8153) );
  NAND2_X1 U9891 ( .A1(n8373), .A2(n13448), .ZN(n8410) );
  NAND2_X1 U9892 ( .A1(n8446), .A2(n13379), .ZN(n8475) );
  INV_X1 U9893 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13370) );
  NAND2_X1 U9894 ( .A1(n13370), .A2(n13344), .ZN(n8155) );
  INV_X1 U9895 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n13360) );
  INV_X1 U9896 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n13227) );
  INV_X1 U9897 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U9898 ( .A1(n8227), .A2(n9969), .ZN(n8229) );
  NAND2_X1 U9899 ( .A1(n8229), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U9900 ( .A1(n8653), .A2(n8156), .ZN(n13642) );
  NOR2_X2 U9901 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8297) );
  NAND2_X1 U9902 ( .A1(n8297), .A2(n8157), .ZN(n8312) );
  INV_X1 U9903 ( .A(n8312), .ZN(n8159) );
  NOR2_X2 U9904 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8161) );
  NOR2_X2 U9905 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8160) );
  NOR2_X1 U9906 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8166) );
  NOR2_X1 U9907 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n8167) );
  INV_X1 U9908 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13915) );
  NAND2_X1 U9909 ( .A1(n13029), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U9910 ( .A1(n13030), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8174) );
  OAI211_X1 U9911 ( .C1(n13915), .C2(n13033), .A(n8175), .B(n8174), .ZN(n8176)
         );
  AOI21_X1 U9912 ( .B1(n13642), .B2(n8654), .A(n8176), .ZN(n9970) );
  INV_X1 U9913 ( .A(n9970), .ZN(n13652) );
  AOI22_X1 U9914 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n12490), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n7848), .ZN(n8236) );
  INV_X1 U9915 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U9916 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11864), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n11866), .ZN(n8535) );
  INV_X1 U9917 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8996) );
  AND2_X1 U9918 ( .A1(n8996), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8285) );
  INV_X1 U9919 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10048) );
  NAND2_X1 U9920 ( .A1(n10048), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8177) );
  INV_X1 U9921 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U9922 ( .A1(n10049), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8179) );
  INV_X1 U9923 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U9924 ( .A1(n8180), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U9925 ( .A1(n10087), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U9926 ( .A1(n8341), .A2(n8340), .ZN(n8185) );
  INV_X1 U9927 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U9928 ( .A1(n8183), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U9929 ( .A1(n10102), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U9930 ( .A1(n8188), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U9931 ( .A1(n8250), .A2(n8249), .ZN(n8191) );
  NAND2_X1 U9932 ( .A1(n10148), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U9933 ( .A1(n8191), .A2(n8190), .ZN(n8380) );
  XNOR2_X1 U9934 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8381) );
  NAND2_X1 U9935 ( .A1(n8380), .A2(n8381), .ZN(n8193) );
  NAND2_X1 U9936 ( .A1(n10162), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8192) );
  XNOR2_X1 U9937 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8405) );
  NAND2_X1 U9938 ( .A1(n10198), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8194) );
  XNOR2_X1 U9939 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8417) );
  XNOR2_X1 U9940 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8423) );
  NAND2_X1 U9941 ( .A1(n8800), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8195) );
  XNOR2_X1 U9942 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8455) );
  NAND2_X1 U9943 ( .A1(n11024), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U9944 ( .A1(n8199), .A2(n8198), .ZN(n8469) );
  XNOR2_X1 U9945 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8470) );
  NAND2_X1 U9946 ( .A1(n11124), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8200) );
  XNOR2_X1 U9947 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n8483) );
  NAND2_X1 U9948 ( .A1(n11236), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U9949 ( .A1(n11407), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8204) );
  NAND2_X1 U9950 ( .A1(n11411), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U9951 ( .A1(n8204), .A2(n8203), .ZN(n8496) );
  NAND2_X1 U9952 ( .A1(n8535), .A2(n8537), .ZN(n8206) );
  AOI22_X1 U9953 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11863), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n12622), .ZN(n8585) );
  INV_X1 U9954 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12146) );
  INV_X1 U9955 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8209) );
  AOI22_X1 U9956 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(P1_DATAO_REG_22__SCAN_IN), .B1(n12146), .B2(n8209), .ZN(n8573) );
  INV_X1 U9957 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U9958 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P1_DATAO_REG_23__SCAN_IN), .B1(n10754), .B2(n10568), .ZN(n8561) );
  NAND2_X1 U9959 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8607), .ZN(n8213) );
  AOI21_X2 U9960 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(n8213), .A(n8212), .ZN(
        n8621) );
  AOI22_X1 U9961 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n12162), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n12670), .ZN(n8622) );
  AOI22_X1 U9962 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n12389), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n12682), .ZN(n8633) );
  NAND2_X1 U9963 ( .A1(n8236), .A2(n8238), .ZN(n8215) );
  AOI22_X1 U9964 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n8878), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n7845), .ZN(n8649) );
  INV_X1 U9965 ( .A(n8649), .ZN(n8216) );
  XNOR2_X1 U9966 ( .A(n8648), .B(n8216), .ZN(n13980) );
  NAND2_X1 U9967 ( .A1(n8715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8220) );
  INV_X1 U9968 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U9969 ( .A1(n13980), .A2(n13028), .ZN(n8226) );
  INV_X4 U9970 ( .A(n8763), .ZN(n10304) );
  NAND2_X4 U9971 ( .A1(n10505), .A2(n10304), .ZN(n13026) );
  INV_X1 U9972 ( .A(SI_28_), .ZN(n13982) );
  OR2_X1 U9973 ( .A1(n13026), .A2(n13982), .ZN(n8225) );
  INV_X1 U9974 ( .A(n8227), .ZN(n8640) );
  NAND2_X1 U9975 ( .A1(n8640), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U9976 ( .A1(n8229), .A2(n8228), .ZN(n13654) );
  NAND2_X1 U9977 ( .A1(n13654), .A2(n8654), .ZN(n8235) );
  INV_X1 U9978 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U9979 ( .A1(n13029), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U9980 ( .A1(n13030), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8230) );
  OAI211_X1 U9981 ( .C1(n8232), .C2(n13033), .A(n8231), .B(n8230), .ZN(n8233)
         );
  INV_X1 U9982 ( .A(n8233), .ZN(n8234) );
  INV_X1 U9983 ( .A(n8236), .ZN(n8237) );
  XNOR2_X1 U9984 ( .A(n8238), .B(n8237), .ZN(n12466) );
  NAND2_X1 U9985 ( .A1(n12466), .A2(n13028), .ZN(n8240) );
  OR2_X1 U9986 ( .A1(n13026), .A2(n13385), .ZN(n8239) );
  NAND2_X2 U9987 ( .A1(n8240), .A2(n8239), .ZN(n8647) );
  NAND2_X1 U9988 ( .A1(n13030), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8248) );
  INV_X1 U9989 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8241) );
  OR2_X1 U9990 ( .A1(n13033), .A2(n8241), .ZN(n8247) );
  INV_X2 U9991 ( .A(n8654), .ZN(n8488) );
  INV_X1 U9992 ( .A(n8242), .ZN(n8374) );
  OAI21_X1 U9993 ( .B1(n8357), .B2(P3_REG3_REG_7__SCAN_IN), .A(
        P3_REG3_REG_8__SCAN_IN), .ZN(n8243) );
  AND2_X1 U9994 ( .A1(n8374), .A2(n8243), .ZN(n12090) );
  OR2_X1 U9995 ( .A1(n8488), .A2(n12090), .ZN(n8246) );
  INV_X1 U9996 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n8244) );
  OR2_X1 U9997 ( .A1(n8528), .A2(n8244), .ZN(n8245) );
  XNOR2_X1 U9998 ( .A(n8250), .B(n8249), .ZN(n10071) );
  OR2_X1 U9999 ( .A1(n8499), .A2(n10071), .ZN(n8255) );
  INV_X1 U10000 ( .A(SI_8_), .ZN(n10070) );
  OR2_X1 U10001 ( .A1(n13026), .A2(n10070), .ZN(n8254) );
  NOR2_X1 U10002 ( .A1(n8251), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8384) );
  OR2_X1 U10003 ( .A1(n8384), .A2(n8708), .ZN(n8252) );
  XNOR2_X1 U10004 ( .A(n8252), .B(P3_IR_REG_8__SCAN_IN), .ZN(n10733) );
  OR2_X1 U10005 ( .A1(n10505), .A2(n10988), .ZN(n8253) );
  NAND2_X1 U10006 ( .A1(n12892), .A2(n12891), .ZN(n12931) );
  INV_X1 U10007 ( .A(n12892), .ZN(n13480) );
  INV_X1 U10008 ( .A(n12891), .ZN(n8681) );
  NAND2_X1 U10009 ( .A1(n13480), .A2(n8681), .ZN(n12936) );
  NAND2_X1 U10010 ( .A1(n12931), .A2(n12936), .ZN(n11927) );
  INV_X1 U10011 ( .A(n11927), .ZN(n13059) );
  NAND2_X1 U10012 ( .A1(n8305), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8261) );
  INV_X1 U10013 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8256) );
  OR2_X1 U10014 ( .A1(n8528), .A2(n8256), .ZN(n8260) );
  INV_X1 U10015 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8257) );
  OR2_X1 U10016 ( .A1(n8544), .A2(n8257), .ZN(n8259) );
  XNOR2_X1 U10017 ( .A(n8357), .B(n13329), .ZN(n12035) );
  OR2_X1 U10018 ( .A1(n8488), .A2(n12035), .ZN(n8258) );
  NAND4_X1 U10019 ( .A1(n8261), .A2(n8260), .A3(n8259), .A4(n8258), .ZN(n13481) );
  INV_X1 U10020 ( .A(n8262), .ZN(n8263) );
  XNOR2_X1 U10021 ( .A(n7194), .B(n8263), .ZN(n10075) );
  OR2_X1 U10022 ( .A1(n8499), .A2(n10075), .ZN(n8268) );
  OR2_X1 U10023 ( .A1(n13026), .A2(SI_7_), .ZN(n8267) );
  NAND2_X1 U10024 ( .A1(n8251), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8265) );
  XNOR2_X1 U10025 ( .A(n8265), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10727) );
  OR2_X1 U10026 ( .A1(n10505), .A2(n10727), .ZN(n8266) );
  NAND2_X1 U10027 ( .A1(n13481), .A2(n11836), .ZN(n11921) );
  AND2_X1 U10028 ( .A1(n13059), .A2(n11921), .ZN(n8371) );
  NAND2_X1 U10029 ( .A1(n8305), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8278) );
  INV_X1 U10030 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8269) );
  INV_X1 U10031 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10513) );
  INV_X1 U10032 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11221) );
  INV_X1 U10033 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8271) );
  INV_X1 U10034 ( .A(n8285), .ZN(n8272) );
  XNOR2_X1 U10035 ( .A(n8273), .B(n8272), .ZN(n8274) );
  INV_X1 U10036 ( .A(SI_1_), .ZN(n8986) );
  MUX2_X1 U10037 ( .A(n8274), .B(n8986), .S(n10316), .Z(n10042) );
  INV_X1 U10038 ( .A(n11217), .ZN(n9748) );
  INV_X1 U10039 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8279) );
  INV_X1 U10040 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10901) );
  INV_X1 U10041 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n13457) );
  INV_X1 U10042 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10888) );
  OR2_X1 U10043 ( .A1(n8544), .A2(n10888), .ZN(n8280) );
  INV_X1 U10044 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10054) );
  INV_X1 U10045 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10314) );
  AND2_X1 U10046 ( .A1(n10314), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8284) );
  NOR2_X1 U10047 ( .A1(n8285), .A2(n8284), .ZN(n10053) );
  OR2_X1 U10048 ( .A1(n8499), .A2(n10053), .ZN(n8287) );
  INV_X1 U10049 ( .A(SI_0_), .ZN(n10315) );
  OR2_X1 U10050 ( .A1(n13026), .A2(n10315), .ZN(n8286) );
  INV_X1 U10051 ( .A(n12895), .ZN(n10571) );
  OR2_X1 U10052 ( .A1(n12896), .A2(n10571), .ZN(n11218) );
  NAND2_X1 U10053 ( .A1(n8678), .A2(n11218), .ZN(n8289) );
  NAND2_X1 U10054 ( .A1(n10572), .A2(n11217), .ZN(n8288) );
  NAND2_X1 U10055 ( .A1(n8289), .A2(n8288), .ZN(n11149) );
  INV_X1 U10056 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n8290) );
  INV_X1 U10057 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10660) );
  OR2_X1 U10058 ( .A1(n8488), .A2(n10660), .ZN(n8295) );
  INV_X1 U10059 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8291) );
  OR2_X1 U10060 ( .A1(n8292), .A2(n8291), .ZN(n8294) );
  INV_X1 U10061 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10584) );
  XNOR2_X1 U10062 ( .A(n8300), .B(n8299), .ZN(n10050) );
  OR2_X1 U10063 ( .A1(n13026), .A2(SI_2_), .ZN(n8301) );
  OAI211_X1 U10064 ( .C1(n10595), .C2(n10505), .A(n8302), .B(n8301), .ZN(
        n11208) );
  XNOR2_X1 U10065 ( .A(n8303), .B(n13486), .ZN(n13057) );
  INV_X1 U10066 ( .A(n13057), .ZN(n12897) );
  INV_X1 U10067 ( .A(n13486), .ZN(n12909) );
  NAND2_X1 U10068 ( .A1(n12909), .A2(n11208), .ZN(n8304) );
  NAND2_X1 U10069 ( .A1(n8305), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8311) );
  INV_X1 U10070 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n8306) );
  OR2_X1 U10071 ( .A1(n8544), .A2(n8306), .ZN(n8310) );
  OR2_X1 U10072 ( .A1(n8488), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8309) );
  INV_X1 U10073 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U10074 ( .A1(n8312), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8313) );
  XNOR2_X1 U10075 ( .A(n8313), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10622) );
  XNOR2_X1 U10076 ( .A(n8315), .B(n8314), .ZN(n10060) );
  OR2_X1 U10077 ( .A1(n8499), .A2(n10060), .ZN(n8317) );
  OR2_X1 U10078 ( .A1(n13026), .A2(SI_3_), .ZN(n8316) );
  OAI211_X1 U10079 ( .C1(n10622), .C2(n10505), .A(n8317), .B(n8316), .ZN(
        n15782) );
  NAND2_X1 U10080 ( .A1(n13485), .A2(n15782), .ZN(n12911) );
  INV_X1 U10081 ( .A(n15782), .ZN(n11449) );
  NAND2_X1 U10082 ( .A1(n13485), .A2(n11449), .ZN(n8318) );
  NAND2_X1 U10083 ( .A1(n11444), .A2(n8318), .ZN(n11250) );
  NAND2_X1 U10084 ( .A1(n13030), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8325) );
  INV_X1 U10085 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10583) );
  OR2_X1 U10086 ( .A1(n8528), .A2(n10583), .ZN(n8324) );
  INV_X1 U10087 ( .A(n8319), .ZN(n8333) );
  NAND2_X1 U10088 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8320) );
  AND2_X1 U10089 ( .A1(n8333), .A2(n8320), .ZN(n11435) );
  OR2_X1 U10090 ( .A1(n8488), .A2(n11435), .ZN(n8323) );
  INV_X1 U10091 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8321) );
  OR2_X1 U10092 ( .A1(n13033), .A2(n8321), .ZN(n8322) );
  OR2_X1 U10093 ( .A1(n13026), .A2(SI_4_), .ZN(n8331) );
  XNOR2_X1 U10094 ( .A(n8327), .B(n8326), .ZN(n10079) );
  OR2_X1 U10095 ( .A1(n8499), .A2(n10079), .ZN(n8330) );
  OR2_X1 U10096 ( .A1(n8312), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n8342) );
  NAND2_X1 U10097 ( .A1(n8342), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8328) );
  XNOR2_X1 U10098 ( .A(n8328), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10640) );
  OR2_X1 U10099 ( .A1(n10505), .A2(n10640), .ZN(n8329) );
  NAND2_X1 U10100 ( .A1(n11497), .A2(n11255), .ZN(n12916) );
  NAND2_X1 U10101 ( .A1(n13484), .A2(n11436), .ZN(n12915) );
  NAND2_X1 U10102 ( .A1(n12916), .A2(n12915), .ZN(n13053) );
  NAND2_X1 U10103 ( .A1(n11250), .A2(n13053), .ZN(n11249) );
  OR2_X1 U10104 ( .A1(n11497), .A2(n11436), .ZN(n8332) );
  NAND2_X1 U10105 ( .A1(n13029), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8339) );
  INV_X1 U10106 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11810) );
  OR2_X1 U10107 ( .A1(n8544), .A2(n11810), .ZN(n8338) );
  NAND2_X1 U10108 ( .A1(n8333), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8334) );
  AND2_X1 U10109 ( .A1(n8355), .A2(n8334), .ZN(n11940) );
  OR2_X1 U10110 ( .A1(n8488), .A2(n11940), .ZN(n8337) );
  INV_X1 U10111 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8335) );
  OR2_X1 U10112 ( .A1(n13033), .A2(n8335), .ZN(n8336) );
  OR2_X1 U10113 ( .A1(n13026), .A2(SI_5_), .ZN(n8352) );
  XNOR2_X1 U10114 ( .A(n8341), .B(n8340), .ZN(n10057) );
  OR2_X1 U10115 ( .A1(n8499), .A2(n10057), .ZN(n8351) );
  INV_X1 U10116 ( .A(n8342), .ZN(n8344) );
  NAND2_X1 U10117 ( .A1(n8344), .A2(n8343), .ZN(n8346) );
  NAND2_X1 U10118 ( .A1(n8346), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8345) );
  MUX2_X1 U10119 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8345), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8349) );
  INV_X1 U10120 ( .A(n8346), .ZN(n8348) );
  NAND2_X1 U10121 ( .A1(n8348), .A2(n8347), .ZN(n8364) );
  OR2_X1 U10122 ( .A1(n10505), .A2(n10634), .ZN(n8350) );
  NAND2_X1 U10123 ( .A1(n11856), .A2(n11811), .ZN(n12919) );
  INV_X1 U10124 ( .A(n11811), .ZN(n11941) );
  NAND2_X1 U10125 ( .A1(n13483), .A2(n11941), .ZN(n12920) );
  NAND2_X1 U10126 ( .A1(n11856), .A2(n11941), .ZN(n8354) );
  NAND2_X1 U10127 ( .A1(n13030), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8362) );
  OR2_X1 U10128 ( .A1(n8528), .A2(n15809), .ZN(n8361) );
  NAND2_X1 U10129 ( .A1(n8355), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8356) );
  AND2_X1 U10130 ( .A1(n8357), .A2(n8356), .ZN(n15803) );
  OR2_X1 U10131 ( .A1(n8488), .A2(n15803), .ZN(n8360) );
  INV_X1 U10132 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8358) );
  OR2_X1 U10133 ( .A1(n13033), .A2(n8358), .ZN(n8359) );
  NAND2_X1 U10134 ( .A1(n8364), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8365) );
  XNOR2_X1 U10135 ( .A(n8363), .B(n8365), .ZN(n10716) );
  XNOR2_X1 U10136 ( .A(n10099), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8366) );
  XNOR2_X1 U10137 ( .A(n8367), .B(n8366), .ZN(n10056) );
  OR2_X1 U10138 ( .A1(n8499), .A2(n10056), .ZN(n8369) );
  INV_X1 U10139 ( .A(SI_6_), .ZN(n10055) );
  OR2_X1 U10140 ( .A1(n13026), .A2(n10055), .ZN(n8368) );
  OAI211_X1 U10141 ( .C1(n10505), .C2(n10716), .A(n8369), .B(n8368), .ZN(
        n11675) );
  NAND2_X1 U10142 ( .A1(n11935), .A2(n11675), .ZN(n12924) );
  INV_X1 U10143 ( .A(n11675), .ZN(n15805) );
  NAND2_X1 U10144 ( .A1(n13482), .A2(n15805), .ZN(n12923) );
  INV_X1 U10145 ( .A(n13054), .ZN(n11669) );
  NAND2_X1 U10146 ( .A1(n11670), .A2(n11669), .ZN(n11668) );
  OR2_X1 U10147 ( .A1(n11935), .A2(n15805), .ZN(n8370) );
  NAND2_X1 U10148 ( .A1(n11668), .A2(n8370), .ZN(n11829) );
  XNOR2_X1 U10149 ( .A(n13481), .B(n11836), .ZN(n12926) );
  NAND2_X1 U10150 ( .A1(n11829), .A2(n7766), .ZN(n11922) );
  NAND2_X1 U10151 ( .A1(n8371), .A2(n11922), .ZN(n11923) );
  NAND2_X1 U10152 ( .A1(n8305), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8379) );
  INV_X1 U10153 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n8372) );
  OR2_X1 U10154 ( .A1(n8544), .A2(n8372), .ZN(n8378) );
  INV_X1 U10155 ( .A(n8373), .ZN(n8393) );
  NAND2_X1 U10156 ( .A1(n8374), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8375) );
  AND2_X1 U10157 ( .A1(n8393), .A2(n8375), .ZN(n12173) );
  OR2_X1 U10158 ( .A1(n8488), .A2(n12173), .ZN(n8377) );
  INV_X1 U10159 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12045) );
  OR2_X1 U10160 ( .A1(n8528), .A2(n12045), .ZN(n8376) );
  INV_X1 U10161 ( .A(n8381), .ZN(n8382) );
  XNOR2_X1 U10162 ( .A(n8380), .B(n8382), .ZN(n10072) );
  OR2_X1 U10163 ( .A1(n8499), .A2(n10072), .ZN(n8391) );
  OR2_X1 U10164 ( .A1(n13026), .A2(SI_9_), .ZN(n8390) );
  AND2_X1 U10165 ( .A1(n8384), .A2(n8383), .ZN(n8387) );
  NOR2_X1 U10166 ( .A1(n8387), .A2(n8708), .ZN(n8385) );
  MUX2_X1 U10167 ( .A(n8708), .B(n8385), .S(P3_IR_REG_9__SCAN_IN), .Z(n8388)
         );
  OR2_X1 U10168 ( .A1(n10505), .A2(n11541), .ZN(n8389) );
  NAND2_X1 U10169 ( .A1(n13030), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8399) );
  INV_X1 U10170 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n8392) );
  OR2_X1 U10171 ( .A1(n8528), .A2(n8392), .ZN(n8398) );
  NAND2_X1 U10172 ( .A1(n8393), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8394) );
  AND2_X1 U10173 ( .A1(n8410), .A2(n8394), .ZN(n12260) );
  OR2_X1 U10174 ( .A1(n8488), .A2(n12260), .ZN(n8397) );
  INV_X1 U10175 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8395) );
  OR2_X1 U10176 ( .A1(n13033), .A2(n8395), .ZN(n8396) );
  INV_X1 U10177 ( .A(SI_10_), .ZN(n13304) );
  NOR2_X1 U10178 ( .A1(n8403), .A2(n8708), .ZN(n8400) );
  MUX2_X1 U10179 ( .A(n8708), .B(n8400), .S(P3_IR_REG_10__SCAN_IN), .Z(n8401)
         );
  INV_X1 U10180 ( .A(n8401), .ZN(n8404) );
  INV_X1 U10181 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10182 ( .A1(n8403), .A2(n8402), .ZN(n8425) );
  AOI22_X1 U10183 ( .A1(n13021), .A2(n13304), .B1(n8541), .B2(n11553), .ZN(
        n8408) );
  XNOR2_X1 U10184 ( .A(n8406), .B(n8405), .ZN(n10069) );
  NAND2_X1 U10185 ( .A1(n10069), .A2(n13028), .ZN(n8407) );
  NAND2_X1 U10186 ( .A1(n12379), .A2(n12248), .ZN(n12943) );
  INV_X1 U10187 ( .A(n12379), .ZN(n13479) );
  NAND2_X1 U10188 ( .A1(n13479), .A2(n15885), .ZN(n12944) );
  INV_X1 U10189 ( .A(n13062), .ZN(n8409) );
  NAND2_X1 U10190 ( .A1(n8305), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8415) );
  INV_X1 U10191 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11538) );
  OR2_X1 U10192 ( .A1(n8544), .A2(n11538), .ZN(n8414) );
  INV_X1 U10193 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12384) );
  OR2_X1 U10194 ( .A1(n8528), .A2(n12384), .ZN(n8413) );
  NAND2_X1 U10195 ( .A1(n8410), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8411) );
  AND2_X1 U10196 ( .A1(n8430), .A2(n8411), .ZN(n12383) );
  OR2_X1 U10197 ( .A1(n8488), .A2(n12383), .ZN(n8412) );
  XNOR2_X1 U10198 ( .A(n8416), .B(n8417), .ZN(n10078) );
  NAND2_X1 U10199 ( .A1(n10078), .A2(n13028), .ZN(n8421) );
  NAND2_X1 U10200 ( .A1(n8425), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8419) );
  INV_X1 U10201 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8418) );
  XNOR2_X1 U10202 ( .A(n8419), .B(n8418), .ZN(n12303) );
  AOI22_X1 U10203 ( .A1(n13021), .A2(n13419), .B1(n8541), .B2(n12303), .ZN(
        n8420) );
  NAND2_X1 U10204 ( .A1(n13266), .A2(n12324), .ZN(n9768) );
  NAND2_X1 U10205 ( .A1(n12377), .A2(n9768), .ZN(n8422) );
  NAND2_X1 U10206 ( .A1(n15913), .A2(n12552), .ZN(n9766) );
  NAND2_X1 U10207 ( .A1(n8422), .A2(n9766), .ZN(n12551) );
  XNOR2_X1 U10208 ( .A(n8424), .B(n8423), .ZN(n10089) );
  NAND2_X1 U10209 ( .A1(n10089), .A2(n13028), .ZN(n8429) );
  OAI21_X1 U10210 ( .B1(n8425), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8427) );
  INV_X1 U10211 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8426) );
  XNOR2_X1 U10212 ( .A(n8427), .B(n8426), .ZN(n12302) );
  AOI22_X1 U10213 ( .A1(n13021), .A2(n13414), .B1(n8541), .B2(n12302), .ZN(
        n8428) );
  NAND2_X1 U10214 ( .A1(n13030), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8435) );
  INV_X1 U10215 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12559) );
  OR2_X1 U10216 ( .A1(n8528), .A2(n12559), .ZN(n8434) );
  NAND2_X1 U10217 ( .A1(n8430), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8431) );
  AND2_X1 U10218 ( .A1(n8447), .A2(n8431), .ZN(n12560) );
  OR2_X1 U10219 ( .A1(n8488), .A2(n12560), .ZN(n8433) );
  INV_X1 U10220 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n12565) );
  OR2_X1 U10221 ( .A1(n13033), .A2(n12565), .ZN(n8432) );
  NAND2_X1 U10222 ( .A1(n12566), .A2(n13264), .ZN(n9772) );
  NAND2_X1 U10223 ( .A1(n12551), .A2(n9772), .ZN(n8436) );
  OR2_X1 U10224 ( .A1(n12566), .A2(n13264), .ZN(n9773) );
  NAND2_X1 U10225 ( .A1(n8436), .A2(n9773), .ZN(n12515) );
  XNOR2_X1 U10226 ( .A(n8437), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U10227 ( .A1(n10143), .A2(n13028), .ZN(n8445) );
  NOR2_X1 U10228 ( .A1(n8438), .A2(n8708), .ZN(n8439) );
  MUX2_X1 U10229 ( .A(n8708), .B(n8439), .S(P3_IR_REG_13__SCAN_IN), .Z(n8440)
         );
  INV_X1 U10230 ( .A(n8440), .ZN(n8443) );
  INV_X1 U10231 ( .A(n8441), .ZN(n8442) );
  NAND2_X1 U10232 ( .A1(n8443), .A2(n8442), .ZN(n13501) );
  AOI22_X1 U10233 ( .A1(n13021), .A2(n13299), .B1(n8541), .B2(n13501), .ZN(
        n8444) );
  NAND2_X1 U10234 ( .A1(n8445), .A2(n8444), .ZN(n12958) );
  NAND2_X1 U10235 ( .A1(n8305), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8452) );
  INV_X1 U10236 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12526) );
  OR2_X1 U10237 ( .A1(n8528), .A2(n12526), .ZN(n8451) );
  INV_X1 U10238 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12290) );
  OR2_X1 U10239 ( .A1(n8544), .A2(n12290), .ZN(n8450) );
  INV_X1 U10240 ( .A(n8446), .ZN(n8463) );
  NAND2_X1 U10241 ( .A1(n8447), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8448) );
  AND2_X1 U10242 ( .A1(n8463), .A2(n8448), .ZN(n12460) );
  OR2_X1 U10243 ( .A1(n8488), .A2(n12460), .ZN(n8449) );
  XNOR2_X1 U10244 ( .A(n12958), .B(n12957), .ZN(n13065) );
  OR2_X1 U10245 ( .A1(n12958), .A2(n12957), .ZN(n8453) );
  XNOR2_X1 U10246 ( .A(n8454), .B(n8455), .ZN(n10153) );
  NAND2_X1 U10247 ( .A1(n10153), .A2(n13028), .ZN(n8461) );
  NOR2_X1 U10248 ( .A1(n8441), .A2(n8708), .ZN(n8456) );
  MUX2_X1 U10249 ( .A(n8708), .B(n8456), .S(P3_IR_REG_14__SCAN_IN), .Z(n8457)
         );
  INV_X1 U10250 ( .A(n8457), .ZN(n8459) );
  NAND2_X1 U10251 ( .A1(n8459), .A2(n8458), .ZN(n13517) );
  AOI22_X1 U10252 ( .A1(n13021), .A2(n13272), .B1(n8541), .B2(n13517), .ZN(
        n8460) );
  NAND2_X1 U10253 ( .A1(n8461), .A2(n8460), .ZN(n13913) );
  NAND2_X1 U10254 ( .A1(n13030), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8468) );
  INV_X1 U10255 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n8462) );
  OR2_X1 U10256 ( .A1(n13033), .A2(n8462), .ZN(n8467) );
  NAND2_X1 U10257 ( .A1(n8463), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8464) );
  AND2_X1 U10258 ( .A1(n8475), .A2(n8464), .ZN(n12483) );
  OR2_X1 U10259 ( .A1(n8488), .A2(n12483), .ZN(n8466) );
  INV_X1 U10260 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12310) );
  OR2_X1 U10261 ( .A1(n8528), .A2(n12310), .ZN(n8465) );
  NAND4_X1 U10262 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(n13263) );
  NOR2_X1 U10263 ( .A1(n13913), .A2(n13263), .ZN(n12962) );
  INV_X1 U10264 ( .A(n12962), .ZN(n8685) );
  NAND2_X1 U10265 ( .A1(n13913), .A2(n13263), .ZN(n12963) );
  NAND2_X1 U10266 ( .A1(n8685), .A2(n12963), .ZN(n13067) );
  INV_X1 U10267 ( .A(n13263), .ZN(n13248) );
  XNOR2_X1 U10268 ( .A(n8469), .B(n8470), .ZN(n10154) );
  NAND2_X1 U10269 ( .A1(n10154), .A2(n13028), .ZN(n8474) );
  NAND2_X1 U10270 ( .A1(n8458), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8472) );
  INV_X1 U10271 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8471) );
  XNOR2_X1 U10272 ( .A(n8472), .B(n8471), .ZN(n13536) );
  AOI22_X1 U10273 ( .A1(n13021), .A2(n13412), .B1(n8541), .B2(n13536), .ZN(
        n8473) );
  NAND2_X1 U10274 ( .A1(n8305), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8480) );
  INV_X1 U10275 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13519) );
  OR2_X1 U10276 ( .A1(n8544), .A2(n13519), .ZN(n8479) );
  NAND2_X1 U10277 ( .A1(n8475), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8476) );
  AND2_X1 U10278 ( .A1(n8506), .A2(n8476), .ZN(n12535) );
  OR2_X1 U10279 ( .A1(n8488), .A2(n12535), .ZN(n8478) );
  INV_X1 U10280 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13520) );
  OR2_X1 U10281 ( .A1(n8528), .A2(n13520), .ZN(n8477) );
  XNOR2_X1 U10282 ( .A(n13254), .B(n13832), .ZN(n13070) );
  OR2_X1 U10283 ( .A1(n13254), .A2(n13832), .ZN(n8481) );
  NAND2_X1 U10284 ( .A1(n8482), .A2(n8481), .ZN(n13828) );
  INV_X1 U10285 ( .A(n13828), .ZN(n8494) );
  INV_X1 U10286 ( .A(n8483), .ZN(n8484) );
  XNOR2_X1 U10287 ( .A(n8485), .B(n8484), .ZN(n10195) );
  NAND2_X1 U10288 ( .A1(n10195), .A2(n13028), .ZN(n8487) );
  NAND2_X1 U10289 ( .A1(n8516), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8500) );
  XNOR2_X1 U10290 ( .A(n8500), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U10291 ( .A1(n13021), .A2(SI_16_), .B1(n8541), .B2(n13541), .ZN(
        n8486) );
  NAND2_X1 U10292 ( .A1(n8305), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8492) );
  INV_X1 U10293 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13838) );
  OR2_X1 U10294 ( .A1(n8528), .A2(n13838), .ZN(n8491) );
  INV_X1 U10295 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13903) );
  OR2_X1 U10296 ( .A1(n8544), .A2(n13903), .ZN(n8490) );
  XNOR2_X1 U10297 ( .A(n8506), .B(n13370), .ZN(n13837) );
  OR2_X1 U10298 ( .A1(n8488), .A2(n13837), .ZN(n8489) );
  NAND4_X1 U10299 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n13261) );
  NOR2_X1 U10300 ( .A1(n13836), .A2(n13261), .ZN(n12972) );
  INV_X1 U10301 ( .A(n12972), .ZN(n8495) );
  NAND2_X1 U10302 ( .A1(n13836), .A2(n13261), .ZN(n12970) );
  NAND2_X1 U10303 ( .A1(n8495), .A2(n12970), .ZN(n13829) );
  INV_X1 U10304 ( .A(n13829), .ZN(n8493) );
  INV_X1 U10305 ( .A(n8496), .ZN(n8497) );
  XNOR2_X1 U10306 ( .A(n8498), .B(n8497), .ZN(n10217) );
  NAND2_X1 U10307 ( .A1(n10217), .A2(n13028), .ZN(n8504) );
  NAND2_X1 U10308 ( .A1(n8500), .A2(n8514), .ZN(n8501) );
  NAND2_X1 U10309 ( .A1(n8501), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8502) );
  XNOR2_X1 U10310 ( .A(n8502), .B(n8513), .ZN(n13579) );
  AOI22_X1 U10311 ( .A1(n13021), .A2(n13405), .B1(n8541), .B2(n13579), .ZN(
        n8503) );
  NAND2_X1 U10312 ( .A1(n8504), .A2(n8503), .ZN(n13900) );
  NAND2_X1 U10313 ( .A1(n8305), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8511) );
  INV_X1 U10314 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13554) );
  OR2_X1 U10315 ( .A1(n8544), .A2(n13554), .ZN(n8510) );
  INV_X1 U10316 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13814) );
  OR2_X1 U10317 ( .A1(n8528), .A2(n13814), .ZN(n8509) );
  INV_X1 U10318 ( .A(n8505), .ZN(n8525) );
  OAI21_X1 U10319 ( .B1(n8506), .B2(P3_REG3_REG_16__SCAN_IN), .A(
        P3_REG3_REG_17__SCAN_IN), .ZN(n8507) );
  AND2_X1 U10320 ( .A1(n8525), .A2(n8507), .ZN(n13813) );
  OR2_X1 U10321 ( .A1(n8488), .A2(n13813), .ZN(n8508) );
  NAND4_X1 U10322 ( .A1(n8511), .A2(n8510), .A3(n8509), .A4(n8508), .ZN(n13260) );
  OR2_X1 U10323 ( .A1(n13900), .A2(n13260), .ZN(n13790) );
  NAND2_X1 U10324 ( .A1(n13900), .A2(n13260), .ZN(n12977) );
  XNOR2_X1 U10325 ( .A(n8512), .B(n7341), .ZN(n10569) );
  NAND2_X1 U10326 ( .A1(n10569), .A2(n13028), .ZN(n8523) );
  NAND2_X1 U10327 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  INV_X1 U10328 ( .A(n8520), .ZN(n8517) );
  NAND2_X1 U10329 ( .A1(n8517), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8518) );
  MUX2_X1 U10330 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8518), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8521) );
  AND2_X1 U10331 ( .A1(n8521), .A2(n7232), .ZN(n13599) );
  AOI22_X1 U10332 ( .A1(n13021), .A2(SI_18_), .B1(n8541), .B2(n13599), .ZN(
        n8522) );
  NAND2_X1 U10333 ( .A1(n8523), .A2(n8522), .ZN(n12573) );
  INV_X1 U10334 ( .A(n8524), .ZN(n8547) );
  NAND2_X1 U10335 ( .A1(n8525), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U10336 ( .A1(n8547), .A2(n8526), .ZN(n13801) );
  NAND2_X1 U10337 ( .A1(n8654), .A2(n13801), .ZN(n8532) );
  INV_X1 U10338 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13895) );
  OR2_X1 U10339 ( .A1(n8544), .A2(n13895), .ZN(n8531) );
  INV_X1 U10340 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n8527) );
  OR2_X1 U10341 ( .A1(n8528), .A2(n8527), .ZN(n8530) );
  INV_X1 U10342 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13953) );
  OR2_X1 U10343 ( .A1(n13033), .A2(n13953), .ZN(n8529) );
  OR2_X1 U10344 ( .A1(n12573), .A2(n13808), .ZN(n12976) );
  NAND2_X1 U10345 ( .A1(n12573), .A2(n13808), .ZN(n12979) );
  NAND2_X1 U10346 ( .A1(n12976), .A2(n12979), .ZN(n13795) );
  OR2_X1 U10347 ( .A1(n13900), .A2(n13834), .ZN(n13796) );
  AND2_X1 U10348 ( .A1(n13795), .A2(n13796), .ZN(n8533) );
  NAND2_X1 U10349 ( .A1(n13811), .A2(n8533), .ZN(n13794) );
  INV_X1 U10350 ( .A(n13808), .ZN(n13259) );
  OR2_X1 U10351 ( .A1(n12573), .A2(n13259), .ZN(n8534) );
  NAND2_X1 U10352 ( .A1(n13794), .A2(n8534), .ZN(n13774) );
  INV_X1 U10353 ( .A(n8535), .ZN(n8536) );
  XNOR2_X1 U10354 ( .A(n8537), .B(n8536), .ZN(n10842) );
  NAND2_X1 U10355 ( .A1(n10842), .A2(n13028), .ZN(n8543) );
  NAND2_X1 U10356 ( .A1(n7232), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8538) );
  MUX2_X1 U10357 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8538), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8540) );
  AOI22_X1 U10358 ( .A1(n13021), .A2(SI_19_), .B1(n8706), .B2(n8541), .ZN(
        n8542) );
  INV_X1 U10359 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13891) );
  OR2_X1 U10360 ( .A1(n8544), .A2(n13891), .ZN(n8546) );
  INV_X1 U10361 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13949) );
  OR2_X1 U10362 ( .A1(n13033), .A2(n13949), .ZN(n8545) );
  AND2_X1 U10363 ( .A1(n8546), .A2(n8545), .ZN(n8551) );
  NAND2_X1 U10364 ( .A1(n8547), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10365 ( .A1(n8557), .A2(n8548), .ZN(n13785) );
  NAND2_X1 U10366 ( .A1(n13785), .A2(n8654), .ZN(n8550) );
  NAND2_X1 U10367 ( .A1(n13029), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10368 ( .A1(n13784), .A2(n13760), .ZN(n8552) );
  OR2_X1 U10369 ( .A1(n13784), .A2(n13760), .ZN(n8553) );
  XNOR2_X1 U10370 ( .A(n8554), .B(n12609), .ZN(n11144) );
  NAND2_X1 U10371 ( .A1(n11144), .A2(n13028), .ZN(n8556) );
  OR2_X1 U10372 ( .A1(n13026), .A2(n13381), .ZN(n8555) );
  INV_X1 U10373 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13943) );
  NAND2_X1 U10374 ( .A1(n8557), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10375 ( .A1(n8590), .A2(n8558), .ZN(n13768) );
  NAND2_X1 U10376 ( .A1(n13768), .A2(n8654), .ZN(n8560) );
  AOI22_X1 U10377 ( .A1(n13029), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n13030), 
        .B2(P3_REG1_REG_20__SCAN_IN), .ZN(n8559) );
  OAI211_X1 U10378 ( .C1(n13033), .C2(n13943), .A(n8560), .B(n8559), .ZN(
        n13741) );
  NAND2_X1 U10379 ( .A1(n13879), .A2(n13741), .ZN(n12989) );
  INV_X1 U10380 ( .A(n13741), .ZN(n13776) );
  NAND2_X1 U10381 ( .A1(n13219), .A2(n13776), .ZN(n12988) );
  XNOR2_X1 U10382 ( .A(n8562), .B(n8561), .ZN(n11739) );
  NAND2_X1 U10383 ( .A1(n11739), .A2(n13028), .ZN(n8564) );
  OR2_X1 U10384 ( .A1(n13026), .A2(n13390), .ZN(n8563) );
  INV_X1 U10385 ( .A(n8565), .ZN(n8579) );
  NAND2_X1 U10386 ( .A1(n8579), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10387 ( .A1(n8612), .A2(n8566), .ZN(n13713) );
  NAND2_X1 U10388 ( .A1(n13713), .A2(n8654), .ZN(n8572) );
  INV_X1 U10389 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10390 ( .A1(n13030), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U10391 ( .A1(n13029), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8567) );
  OAI211_X1 U10392 ( .C1(n8569), .C2(n13033), .A(n8568), .B(n8567), .ZN(n8570)
         );
  INV_X1 U10393 ( .A(n8570), .ZN(n8571) );
  NAND2_X1 U10394 ( .A1(n13933), .A2(n13690), .ZN(n8602) );
  INV_X1 U10395 ( .A(n8602), .ZN(n8599) );
  XNOR2_X1 U10396 ( .A(n13933), .B(n13727), .ZN(n12999) );
  XNOR2_X1 U10397 ( .A(n8574), .B(n8573), .ZN(n11424) );
  NAND2_X1 U10398 ( .A1(n11424), .A2(n13028), .ZN(n8576) );
  OR2_X1 U10399 ( .A1(n13026), .A2(n9252), .ZN(n8575) );
  INV_X1 U10400 ( .A(n8577), .ZN(n8592) );
  NAND2_X1 U10401 ( .A1(n8592), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U10402 ( .A1(n8579), .A2(n8578), .ZN(n13732) );
  NAND2_X1 U10403 ( .A1(n13732), .A2(n8654), .ZN(n8584) );
  INV_X1 U10404 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13936) );
  NAND2_X1 U10405 ( .A1(n13030), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U10406 ( .A1(n13029), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8580) );
  OAI211_X1 U10407 ( .C1(n13033), .C2(n13936), .A(n8581), .B(n8580), .ZN(n8582) );
  INV_X1 U10408 ( .A(n8582), .ZN(n8583) );
  NAND2_X1 U10409 ( .A1(n13870), .A2(n13743), .ZN(n8601) );
  INV_X1 U10410 ( .A(n8601), .ZN(n8597) );
  INV_X1 U10411 ( .A(n8585), .ZN(n8586) );
  XNOR2_X1 U10412 ( .A(n8587), .B(n8586), .ZN(n11317) );
  NAND2_X1 U10413 ( .A1(n11317), .A2(n13028), .ZN(n8589) );
  INV_X1 U10414 ( .A(SI_21_), .ZN(n13398) );
  OR2_X1 U10415 ( .A1(n13026), .A2(n13398), .ZN(n8588) );
  NAND2_X1 U10416 ( .A1(n8590), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U10417 ( .A1(n8592), .A2(n8591), .ZN(n13749) );
  NAND2_X1 U10418 ( .A1(n13749), .A2(n8654), .ZN(n8595) );
  AOI22_X1 U10419 ( .A1(n13029), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13030), 
        .B2(P3_REG1_REG_21__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10420 ( .A1(n8305), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8593) );
  INV_X1 U10421 ( .A(n13763), .ZN(n13258) );
  OR2_X1 U10422 ( .A1(n13873), .A2(n13258), .ZN(n13723) );
  AND2_X1 U10423 ( .A1(n7304), .A2(n13723), .ZN(n8596) );
  OR2_X1 U10424 ( .A1(n8597), .A2(n8596), .ZN(n13705) );
  AND2_X1 U10425 ( .A1(n12999), .A2(n13705), .ZN(n8598) );
  NOR2_X1 U10426 ( .A1(n8599), .A2(n8598), .ZN(n8605) );
  OR2_X1 U10427 ( .A1(n13765), .A2(n8605), .ZN(n8600) );
  NAND2_X1 U10428 ( .A1(n13873), .A2(n13763), .ZN(n13717) );
  AND2_X1 U10429 ( .A1(n13745), .A2(n8601), .ZN(n13704) );
  AND2_X1 U10430 ( .A1(n13704), .A2(n8602), .ZN(n8603) );
  NAND2_X1 U10431 ( .A1(n13219), .A2(n13741), .ZN(n13703) );
  AND2_X1 U10432 ( .A1(n8603), .A2(n13703), .ZN(n8604) );
  OR2_X1 U10433 ( .A1(n8605), .A2(n8604), .ZN(n8606) );
  XOR2_X1 U10434 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n8607), .Z(n8609) );
  NOR2_X1 U10435 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n8609), .ZN(n8608) );
  AOI21_X1 U10436 ( .B1(n8609), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8608), .ZN(
        n8610) );
  INV_X1 U10437 ( .A(n8610), .ZN(n8611) );
  MUX2_X1 U10438 ( .A(SI_24_), .B(n8611), .S(n12638), .Z(n13984) );
  NAND2_X1 U10439 ( .A1(n8612), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U10440 ( .A1(n8626), .A2(n8613), .ZN(n13698) );
  NAND2_X1 U10441 ( .A1(n13698), .A2(n8654), .ZN(n8619) );
  INV_X1 U10442 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U10443 ( .A1(n13029), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U10444 ( .A1(n13030), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8614) );
  OAI211_X1 U10445 ( .C1(n8616), .C2(n13033), .A(n8615), .B(n8614), .ZN(n8617)
         );
  INV_X1 U10446 ( .A(n8617), .ZN(n8618) );
  NAND2_X1 U10447 ( .A1(n8619), .A2(n8618), .ZN(n13708) );
  INV_X1 U10448 ( .A(n13708), .ZN(n13674) );
  NOR2_X1 U10449 ( .A1(n13927), .A2(n13674), .ZN(n8620) );
  INV_X1 U10450 ( .A(n13927), .ZN(n13699) );
  INV_X1 U10451 ( .A(n8622), .ZN(n8623) );
  XNOR2_X1 U10452 ( .A(n8621), .B(n8623), .ZN(n12264) );
  NAND2_X1 U10453 ( .A1(n12264), .A2(n13028), .ZN(n8625) );
  INV_X1 U10454 ( .A(SI_25_), .ZN(n12266) );
  OR2_X1 U10455 ( .A1(n13026), .A2(n12266), .ZN(n8624) );
  NAND2_X1 U10456 ( .A1(n8626), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U10457 ( .A1(n8638), .A2(n8627), .ZN(n13679) );
  NAND2_X1 U10458 ( .A1(n13679), .A2(n8654), .ZN(n8632) );
  INV_X1 U10459 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13922) );
  NAND2_X1 U10460 ( .A1(n13029), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U10461 ( .A1(n13030), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8628) );
  OAI211_X1 U10462 ( .C1(n13922), .C2(n13033), .A(n8629), .B(n8628), .ZN(n8630) );
  INV_X1 U10463 ( .A(n8630), .ZN(n8631) );
  XNOR2_X1 U10464 ( .A(n13683), .B(n13691), .ZN(n13684) );
  INV_X1 U10465 ( .A(n8633), .ZN(n8634) );
  NAND2_X1 U10466 ( .A1(n12870), .A2(n13028), .ZN(n8637) );
  INV_X1 U10467 ( .A(SI_26_), .ZN(n12872) );
  OR2_X1 U10468 ( .A1(n13026), .A2(n12872), .ZN(n8636) );
  NAND2_X1 U10469 ( .A1(n8638), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8639) );
  NAND2_X1 U10470 ( .A1(n8640), .A2(n8639), .ZN(n13666) );
  NAND2_X1 U10471 ( .A1(n13666), .A2(n8654), .ZN(n8645) );
  INV_X1 U10472 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13919) );
  NAND2_X1 U10473 ( .A1(n13029), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8642) );
  NAND2_X1 U10474 ( .A1(n13030), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8641) );
  OAI211_X1 U10475 ( .C1(n13919), .C2(n13033), .A(n8642), .B(n8641), .ZN(n8643) );
  INV_X1 U10476 ( .A(n8643), .ZN(n8644) );
  NAND2_X1 U10477 ( .A1(n13921), .A2(n13675), .ZN(n8646) );
  NAND2_X1 U10478 ( .A1(n8647), .A2(n13663), .ZN(n12882) );
  NAND2_X2 U10479 ( .A1(n12879), .A2(n12882), .ZN(n13649) );
  NAND2_X1 U10480 ( .A1(n13650), .A2(n13649), .ZN(n13648) );
  OAI21_X1 U10481 ( .B1(n13257), .B2(n8647), .A(n13648), .ZN(n13631) );
  NAND2_X1 U10482 ( .A1(n13638), .A2(n9970), .ZN(n13010) );
  INV_X1 U10483 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14946) );
  INV_X1 U10484 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12547) );
  OAI22_X1 U10485 ( .A1(n14946), .A2(n12547), .B1(P1_DATAO_REG_29__SCAN_IN), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13019) );
  INV_X1 U10486 ( .A(n13019), .ZN(n8650) );
  XNOR2_X1 U10487 ( .A(n13018), .B(n8650), .ZN(n13976) );
  NAND2_X1 U10488 ( .A1(n13976), .A2(n13028), .ZN(n8652) );
  INV_X1 U10489 ( .A(SI_29_), .ZN(n13977) );
  OR2_X1 U10490 ( .A1(n13026), .A2(n13977), .ZN(n8651) );
  NAND2_X1 U10491 ( .A1(n8652), .A2(n8651), .ZN(n8754) );
  INV_X1 U10492 ( .A(n8653), .ZN(n13615) );
  NAND2_X1 U10493 ( .A1(n13615), .A2(n8654), .ZN(n13037) );
  INV_X1 U10494 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9738) );
  NAND2_X1 U10495 ( .A1(n13030), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U10496 ( .A1(n13029), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8655) );
  OAI211_X1 U10497 ( .C1(n9738), .C2(n13033), .A(n8656), .B(n8655), .ZN(n8657)
         );
  INV_X1 U10498 ( .A(n8657), .ZN(n8658) );
  OR2_X1 U10499 ( .A1(n8754), .A2(n13634), .ZN(n13043) );
  NAND2_X1 U10500 ( .A1(n8754), .A2(n13634), .ZN(n13040) );
  XNOR2_X1 U10501 ( .A(n8659), .B(n13051), .ZN(n8677) );
  NAND2_X1 U10502 ( .A1(n8661), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8663) );
  INV_X1 U10503 ( .A(n11146), .ZN(n9733) );
  AND2_X1 U10504 ( .A1(n8747), .A2(n9733), .ZN(n13083) );
  NAND2_X1 U10505 ( .A1(n7288), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8664) );
  MUX2_X1 U10506 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8664), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8666) );
  NAND2_X1 U10507 ( .A1(n8706), .A2(n13092), .ZN(n8704) );
  INV_X1 U10508 ( .A(n8704), .ZN(n9734) );
  INV_X1 U10509 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n8668) );
  AOI22_X1 U10510 ( .A1(n13029), .A2(P3_REG2_REG_30__SCAN_IN), .B1(n13030), 
        .B2(P3_REG1_REG_30__SCAN_IN), .ZN(n8667) );
  OAI211_X1 U10511 ( .C1(n13033), .C2(n8668), .A(n13037), .B(n8667), .ZN(
        n13256) );
  INV_X1 U10512 ( .A(n13256), .ZN(n8673) );
  OR2_X1 U10513 ( .A1(n7186), .A2(n13087), .ZN(n10515) );
  NOR2_X2 U10514 ( .A1(n13012), .A2(n9838), .ZN(n13742) );
  INV_X1 U10515 ( .A(P3_B_REG_SCAN_IN), .ZN(n8671) );
  OR2_X1 U10516 ( .A1(n7186), .A2(n8671), .ZN(n8672) );
  NAND2_X1 U10517 ( .A1(n13742), .A2(n8672), .ZN(n13616) );
  NOR2_X1 U10518 ( .A1(n8673), .A2(n13616), .ZN(n8675) );
  NOR2_X1 U10519 ( .A1(n9970), .A2(n13833), .ZN(n8674) );
  NAND2_X1 U10520 ( .A1(n11223), .A2(n12902), .ZN(n11147) );
  NOR2_X1 U10521 ( .A1(n13486), .A2(n11208), .ZN(n12904) );
  INV_X1 U10522 ( .A(n13053), .ZN(n11247) );
  NAND2_X1 U10523 ( .A1(n11246), .A2(n12916), .ZN(n11500) );
  INV_X1 U10524 ( .A(n13481), .ZN(n12085) );
  NAND2_X1 U10525 ( .A1(n12085), .A2(n11836), .ZN(n12929) );
  NAND2_X1 U10526 ( .A1(n12892), .A2(n8681), .ZN(n8682) );
  NAND2_X1 U10527 ( .A1(n12256), .A2(n15866), .ZN(n12938) );
  INV_X1 U10528 ( .A(n12938), .ZN(n8683) );
  INV_X1 U10529 ( .A(n15866), .ZN(n12168) );
  NAND2_X1 U10530 ( .A1(n7681), .A2(n12168), .ZN(n12939) );
  NAND2_X1 U10531 ( .A1(n12324), .A2(n12552), .ZN(n12950) );
  NAND2_X1 U10532 ( .A1(n15913), .A2(n13266), .ZN(n12947) );
  NAND2_X1 U10533 ( .A1(n12382), .A2(n13061), .ZN(n12381) );
  INV_X1 U10534 ( .A(n12566), .ZN(n8684) );
  NAND2_X1 U10535 ( .A1(n8684), .A2(n13264), .ZN(n12953) );
  NOR2_X1 U10536 ( .A1(n12958), .A2(n9776), .ZN(n12961) );
  NAND2_X1 U10537 ( .A1(n12493), .A2(n7664), .ZN(n8686) );
  NOR2_X1 U10538 ( .A1(n13254), .A2(n13262), .ZN(n12967) );
  INV_X1 U10539 ( .A(n12967), .ZN(n13823) );
  INV_X1 U10540 ( .A(n13261), .ZN(n13809) );
  NAND2_X1 U10541 ( .A1(n13836), .A2(n13809), .ZN(n8687) );
  INV_X1 U10542 ( .A(n8687), .ZN(n8688) );
  AND2_X1 U10543 ( .A1(n13818), .A2(n12976), .ZN(n13777) );
  AND2_X1 U10544 ( .A1(n13777), .A2(n12983), .ZN(n8692) );
  INV_X1 U10545 ( .A(n12983), .ZN(n8691) );
  NAND2_X1 U10546 ( .A1(n13784), .A2(n13800), .ZN(n12984) );
  NAND2_X1 U10547 ( .A1(n12983), .A2(n12984), .ZN(n13781) );
  INV_X1 U10548 ( .A(n13781), .ZN(n8690) );
  INV_X1 U10549 ( .A(n12976), .ZN(n12980) );
  AND2_X1 U10550 ( .A1(n13790), .A2(n12979), .ZN(n8689) );
  OR2_X1 U10551 ( .A1(n12980), .A2(n8689), .ZN(n13779) );
  AND2_X1 U10552 ( .A1(n8690), .A2(n13779), .ZN(n13778) );
  NAND2_X1 U10553 ( .A1(n13764), .A2(n12989), .ZN(n13746) );
  XNOR2_X1 U10554 ( .A(n13870), .B(n13710), .ZN(n13728) );
  NOR2_X1 U10555 ( .A1(n13728), .A2(n12999), .ZN(n8693) );
  AND2_X1 U10556 ( .A1(n8693), .A2(n13717), .ZN(n8694) );
  NOR2_X1 U10557 ( .A1(n13870), .A2(n13710), .ZN(n12997) );
  INV_X1 U10558 ( .A(n12997), .ZN(n13718) );
  INV_X1 U10559 ( .A(n13933), .ZN(n12875) );
  NAND2_X1 U10560 ( .A1(n12875), .A2(n13690), .ZN(n8695) );
  NOR2_X1 U10561 ( .A1(n13927), .A2(n13708), .ZN(n12883) );
  INV_X1 U10562 ( .A(n12883), .ZN(n12874) );
  NAND2_X1 U10563 ( .A1(n13927), .A2(n13708), .ZN(n12886) );
  NAND2_X1 U10564 ( .A1(n13686), .A2(n13684), .ZN(n8698) );
  OR2_X1 U10565 ( .A1(n13683), .A2(n13662), .ZN(n8697) );
  NAND2_X1 U10566 ( .A1(n8698), .A2(n8697), .ZN(n13664) );
  NAND2_X1 U10567 ( .A1(n8699), .A2(n13675), .ZN(n12876) );
  AND2_X2 U10568 ( .A1(n12877), .A2(n12876), .ZN(n13665) );
  INV_X1 U10569 ( .A(n12877), .ZN(n8700) );
  XNOR2_X1 U10570 ( .A(n13044), .B(n13051), .ZN(n13627) );
  OR2_X1 U10571 ( .A1(n9733), .A2(n8747), .ZN(n8748) );
  XNOR2_X1 U10572 ( .A(n8748), .B(n13092), .ZN(n8702) );
  OR2_X1 U10573 ( .A1(n8706), .A2(n8747), .ZN(n8701) );
  NAND2_X1 U10574 ( .A1(n8702), .A2(n8701), .ZN(n9831) );
  NAND2_X1 U10575 ( .A1(n11146), .A2(n13610), .ZN(n13039) );
  INV_X1 U10576 ( .A(n13039), .ZN(n9732) );
  AND2_X1 U10577 ( .A1(n15912), .A2(n9732), .ZN(n8703) );
  NAND2_X1 U10578 ( .A1(n9831), .A2(n8703), .ZN(n8705) );
  NAND2_X1 U10579 ( .A1(n13039), .A2(n8704), .ZN(n8749) );
  OR2_X1 U10580 ( .A1(n8749), .A2(n12899), .ZN(n8745) );
  NOR2_X1 U10581 ( .A1(n13084), .A2(n13092), .ZN(n15889) );
  NAND2_X1 U10582 ( .A1(n8740), .A2(n8710), .ZN(n8712) );
  NAND2_X1 U10583 ( .A1(n8712), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8711) );
  NAND2_X1 U10584 ( .A1(n7273), .A2(n12267), .ZN(n8717) );
  OAI21_X1 U10585 ( .B1(n8712), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8713) );
  MUX2_X1 U10586 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8713), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8714) );
  INV_X1 U10587 ( .A(n12873), .ZN(n8716) );
  INV_X1 U10588 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8718) );
  INV_X1 U10589 ( .A(n8719), .ZN(n8720) );
  NAND2_X1 U10590 ( .A1(n12873), .A2(n8720), .ZN(n8721) );
  INV_X1 U10591 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U10592 ( .A1(n8722), .A2(n8723), .ZN(n8725) );
  INV_X1 U10593 ( .A(n8736), .ZN(n12267) );
  NAND2_X1 U10594 ( .A1(n12873), .A2(n12267), .ZN(n8724) );
  XNOR2_X1 U10595 ( .A(n9743), .B(n13965), .ZN(n8744) );
  NOR2_X1 U10596 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n8729) );
  NOR4_X1 U10597 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8728) );
  NOR4_X1 U10598 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8727) );
  NOR4_X1 U10599 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8726) );
  NAND4_X1 U10600 ( .A1(n8729), .A2(n8728), .A3(n8727), .A4(n8726), .ZN(n8735)
         );
  NOR4_X1 U10601 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8733) );
  NOR4_X1 U10602 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8732) );
  NOR4_X1 U10603 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n8731) );
  NOR4_X1 U10604 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n8730) );
  NAND4_X1 U10605 ( .A1(n8733), .A2(n8732), .A3(n8731), .A4(n8730), .ZN(n8734)
         );
  OAI21_X1 U10606 ( .B1(n8735), .B2(n8734), .A(n8722), .ZN(n9731) );
  NAND2_X1 U10607 ( .A1(n8736), .A2(n8719), .ZN(n8737) );
  NAND2_X1 U10608 ( .A1(n8738), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8739) );
  MUX2_X1 U10609 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8739), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8742) );
  INV_X1 U10610 ( .A(n8740), .ZN(n8741) );
  AND2_X1 U10611 ( .A1(n9731), .A2(n10898), .ZN(n8743) );
  NAND2_X1 U10612 ( .A1(n8745), .A2(n13012), .ZN(n10892) );
  NAND2_X1 U10613 ( .A1(n10892), .A2(n10890), .ZN(n8746) );
  NAND2_X1 U10614 ( .A1(n13965), .A2(n8746), .ZN(n8752) );
  INV_X1 U10615 ( .A(n13965), .ZN(n9730) );
  AOI22_X1 U10616 ( .A1(n12898), .A2(n8749), .B1(n8748), .B2(n12899), .ZN(
        n8750) );
  NAND2_X1 U10617 ( .A1(n9730), .A2(n8750), .ZN(n8751) );
  AND2_X1 U10618 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  INV_X1 U10619 ( .A(n8754), .ZN(n13625) );
  INV_X1 U10620 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8756) );
  NOR2_X1 U10621 ( .A1(n15997), .A2(n8756), .ZN(n8757) );
  AND2_X1 U10622 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8759) );
  AND2_X1 U10623 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U10624 ( .A1(n8995), .A2(n8760), .ZN(n8998) );
  NAND2_X1 U10625 ( .A1(n10318), .A2(n8998), .ZN(n8987) );
  INV_X1 U10626 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U10627 ( .A1(n8995), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8761) );
  OAI211_X1 U10628 ( .C1(n8995), .C2(n10305), .A(n8761), .B(n8986), .ZN(n8762)
         );
  NAND2_X1 U10629 ( .A1(n8987), .A2(n8762), .ZN(n8766) );
  OR2_X1 U10630 ( .A1(n8763), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8764) );
  OAI211_X1 U10631 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n10304), .A(n8764), .B(
        SI_1_), .ZN(n8765) );
  INV_X1 U10632 ( .A(SI_2_), .ZN(n10051) );
  MUX2_X1 U10633 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n10304), .Z(n9011) );
  NAND2_X1 U10634 ( .A1(n9010), .A2(n9011), .ZN(n8769) );
  NAND2_X1 U10635 ( .A1(n8767), .A2(SI_2_), .ZN(n8768) );
  MUX2_X1 U10636 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n10304), .Z(n8771) );
  XNOR2_X1 U10637 ( .A(n8771), .B(SI_3_), .ZN(n9026) );
  INV_X1 U10638 ( .A(n9026), .ZN(n8770) );
  NAND2_X1 U10639 ( .A1(n9027), .A2(n8770), .ZN(n8773) );
  NAND2_X1 U10640 ( .A1(n8771), .A2(SI_3_), .ZN(n8772) );
  MUX2_X1 U10641 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n10304), .Z(n8774) );
  NAND2_X1 U10642 ( .A1(n8774), .A2(SI_5_), .ZN(n8778) );
  XNOR2_X1 U10643 ( .A(n8774), .B(SI_5_), .ZN(n9051) );
  MUX2_X1 U10644 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n10304), .Z(n8777) );
  AND2_X1 U10645 ( .A1(n8776), .A2(n9048), .ZN(n8775) );
  INV_X1 U10646 ( .A(n8776), .ZN(n8780) );
  NAND2_X1 U10647 ( .A1(n8777), .A2(SI_4_), .ZN(n9049) );
  AND2_X1 U10648 ( .A1(n9049), .A2(n8778), .ZN(n8779) );
  MUX2_X1 U10649 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10304), .Z(n8783) );
  XNOR2_X1 U10650 ( .A(n8783), .B(SI_6_), .ZN(n9067) );
  INV_X1 U10651 ( .A(n9067), .ZN(n8782) );
  NAND2_X1 U10652 ( .A1(n8783), .A2(SI_6_), .ZN(n8784) );
  MUX2_X1 U10653 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10304), .Z(n8786) );
  XNOR2_X1 U10654 ( .A(n8786), .B(SI_7_), .ZN(n9081) );
  INV_X1 U10655 ( .A(n9081), .ZN(n8785) );
  NAND2_X1 U10656 ( .A1(n8786), .A2(SI_7_), .ZN(n8787) );
  MUX2_X1 U10657 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10304), .Z(n8789) );
  XNOR2_X1 U10658 ( .A(n8789), .B(SI_8_), .ZN(n9095) );
  INV_X1 U10659 ( .A(n9095), .ZN(n8788) );
  MUX2_X1 U10660 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10304), .Z(n8972) );
  NAND2_X1 U10661 ( .A1(n8790), .A2(SI_9_), .ZN(n8791) );
  MUX2_X1 U10662 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10304), .Z(n8793) );
  XNOR2_X1 U10663 ( .A(n8793), .B(SI_10_), .ZN(n9111) );
  INV_X1 U10664 ( .A(n9111), .ZN(n8792) );
  NAND2_X1 U10665 ( .A1(n8793), .A2(SI_10_), .ZN(n8794) );
  MUX2_X1 U10666 ( .A(n10422), .B(n10424), .S(n10304), .Z(n8796) );
  NAND2_X1 U10667 ( .A1(n8796), .A2(n13419), .ZN(n8799) );
  INV_X1 U10668 ( .A(n8796), .ZN(n8797) );
  NAND2_X1 U10669 ( .A1(n8797), .A2(SI_11_), .ZN(n8798) );
  NAND2_X1 U10670 ( .A1(n8799), .A2(n8798), .ZN(n9127) );
  MUX2_X1 U10671 ( .A(n8800), .B(n10610), .S(n10304), .Z(n8801) );
  NAND2_X1 U10672 ( .A1(n8801), .A2(n13414), .ZN(n8804) );
  INV_X1 U10673 ( .A(n8801), .ZN(n8802) );
  NAND2_X1 U10674 ( .A1(n8802), .A2(SI_12_), .ZN(n8803) );
  MUX2_X1 U10675 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10316), .Z(n8805) );
  XNOR2_X1 U10676 ( .A(n8805), .B(n13299), .ZN(n9156) );
  NAND2_X1 U10677 ( .A1(n8805), .A2(SI_13_), .ZN(n8806) );
  MUX2_X1 U10678 ( .A(n11024), .B(n11018), .S(n10316), .Z(n8808) );
  NAND2_X1 U10679 ( .A1(n8808), .A2(n13272), .ZN(n8811) );
  INV_X1 U10680 ( .A(n8808), .ZN(n8809) );
  NAND2_X1 U10681 ( .A1(n8809), .A2(SI_14_), .ZN(n8810) );
  NAND2_X1 U10682 ( .A1(n8811), .A2(n8810), .ZN(n8961) );
  MUX2_X1 U10683 ( .A(n11124), .B(n11126), .S(n10316), .Z(n8812) );
  NAND2_X1 U10684 ( .A1(n8812), .A2(n13412), .ZN(n8815) );
  INV_X1 U10685 ( .A(n8812), .ZN(n8813) );
  NAND2_X1 U10686 ( .A1(n8813), .A2(SI_15_), .ZN(n8814) );
  MUX2_X1 U10687 ( .A(n11236), .B(n11226), .S(n10316), .Z(n8816) );
  INV_X1 U10688 ( .A(n8816), .ZN(n8817) );
  NAND2_X1 U10689 ( .A1(n8817), .A2(SI_16_), .ZN(n8818) );
  MUX2_X1 U10690 ( .A(n11411), .B(n11407), .S(n10316), .Z(n8820) );
  INV_X1 U10691 ( .A(n8820), .ZN(n8821) );
  NAND2_X1 U10692 ( .A1(n8821), .A2(SI_17_), .ZN(n8822) );
  NAND2_X1 U10693 ( .A1(n9183), .A2(n9182), .ZN(n8824) );
  MUX2_X1 U10694 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10316), .Z(n9202) );
  INV_X1 U10695 ( .A(n9202), .ZN(n8825) );
  MUX2_X1 U10696 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10316), .Z(n8828) );
  NAND2_X1 U10697 ( .A1(n8828), .A2(SI_19_), .ZN(n9208) );
  OAI21_X1 U10698 ( .B1(n13291), .B2(n8825), .A(n9208), .ZN(n8826) );
  INV_X1 U10699 ( .A(n8826), .ZN(n8827) );
  NAND2_X1 U10700 ( .A1(n9204), .A2(n8827), .ZN(n8833) );
  NOR2_X1 U10701 ( .A1(n9202), .A2(SI_18_), .ZN(n8831) );
  INV_X1 U10702 ( .A(n8828), .ZN(n8829) );
  NAND2_X1 U10703 ( .A1(n8829), .A2(n13403), .ZN(n9207) );
  INV_X1 U10704 ( .A(n9207), .ZN(n8830) );
  AOI21_X1 U10705 ( .B1(n8831), .B2(n9208), .A(n8830), .ZN(n8832) );
  NAND2_X1 U10706 ( .A1(n8833), .A2(n8832), .ZN(n9227) );
  MUX2_X1 U10707 ( .A(n12609), .B(n11869), .S(n10316), .Z(n8834) );
  NAND2_X1 U10708 ( .A1(n8834), .A2(n13381), .ZN(n8837) );
  INV_X1 U10709 ( .A(n8834), .ZN(n8835) );
  NAND2_X1 U10710 ( .A1(n8835), .A2(SI_20_), .ZN(n8836) );
  NAND2_X1 U10711 ( .A1(n9227), .A2(n9226), .ZN(n8838) );
  MUX2_X1 U10712 ( .A(n12622), .B(n11863), .S(n10316), .Z(n8839) );
  XNOR2_X1 U10713 ( .A(n8839), .B(SI_21_), .ZN(n9237) );
  INV_X1 U10714 ( .A(n9237), .ZN(n8842) );
  INV_X1 U10715 ( .A(n8839), .ZN(n8840) );
  NAND2_X1 U10716 ( .A1(n8840), .A2(SI_21_), .ZN(n8841) );
  MUX2_X1 U10717 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10316), .Z(n9253) );
  MUX2_X1 U10718 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10316), .Z(n9271) );
  INV_X1 U10719 ( .A(n9271), .ZN(n8843) );
  AOI22_X1 U10720 ( .A1(n9254), .A2(n9252), .B1(n8843), .B2(n13390), .ZN(n8844) );
  OAI21_X1 U10721 ( .B1(n9254), .B2(n9252), .A(n13390), .ZN(n8846) );
  AND2_X1 U10722 ( .A1(SI_22_), .A2(SI_23_), .ZN(n8845) );
  AOI22_X1 U10723 ( .A1(n8846), .A2(n9271), .B1(n9253), .B2(n8845), .ZN(n8847)
         );
  MUX2_X1 U10724 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10316), .Z(n9285) );
  INV_X1 U10725 ( .A(n9285), .ZN(n8848) );
  INV_X1 U10726 ( .A(SI_24_), .ZN(n13391) );
  NAND2_X1 U10727 ( .A1(n8848), .A2(n13391), .ZN(n8849) );
  NAND2_X1 U10728 ( .A1(n9285), .A2(SI_24_), .ZN(n8850) );
  MUX2_X1 U10729 ( .A(n12670), .B(n12162), .S(n10316), .Z(n8851) );
  NAND2_X1 U10730 ( .A1(n8851), .A2(n12266), .ZN(n8854) );
  INV_X1 U10731 ( .A(n8851), .ZN(n8852) );
  NAND2_X1 U10732 ( .A1(n8852), .A2(SI_25_), .ZN(n8853) );
  NAND2_X1 U10733 ( .A1(n8854), .A2(n8853), .ZN(n9299) );
  MUX2_X1 U10734 ( .A(n12682), .B(n12389), .S(n10316), .Z(n8856) );
  XNOR2_X1 U10735 ( .A(n8856), .B(SI_26_), .ZN(n9313) );
  INV_X1 U10736 ( .A(n9313), .ZN(n8855) );
  INV_X1 U10737 ( .A(n8856), .ZN(n8857) );
  MUX2_X1 U10738 ( .A(n7848), .B(n12490), .S(n10316), .Z(n8858) );
  NAND2_X1 U10739 ( .A1(n8913), .A2(n13385), .ZN(n8862) );
  INV_X1 U10740 ( .A(n8858), .ZN(n8859) );
  MUX2_X1 U10741 ( .A(n7845), .B(n8878), .S(n10316), .Z(n8863) );
  NAND2_X1 U10742 ( .A1(n8863), .A2(n13982), .ZN(n9341) );
  INV_X1 U10743 ( .A(n8863), .ZN(n8864) );
  NAND2_X1 U10744 ( .A1(n8864), .A2(SI_28_), .ZN(n8865) );
  NOR2_X1 U10745 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n8870) );
  NOR2_X1 U10746 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), 
        .ZN(n8869) );
  NOR2_X1 U10747 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n8873) );
  NOR2_X1 U10748 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8872) );
  INV_X1 U10749 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U10750 ( .A1(n12698), .A2(n9629), .ZN(n8880) );
  OR2_X1 U10751 ( .A1(n9012), .A2(n8878), .ZN(n8879) );
  INV_X1 U10752 ( .A(n14373), .ZN(n9408) );
  NAND2_X1 U10753 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9058) );
  INV_X1 U10754 ( .A(n9058), .ZN(n8881) );
  NAND2_X1 U10755 ( .A1(n8881), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9073) );
  INV_X1 U10756 ( .A(n9073), .ZN(n8882) );
  NAND2_X1 U10757 ( .A1(n8882), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9087) );
  INV_X1 U10758 ( .A(n9087), .ZN(n8883) );
  NAND2_X1 U10759 ( .A1(n8883), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9100) );
  INV_X1 U10760 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U10761 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n8890) );
  INV_X1 U10762 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n14029) );
  INV_X1 U10763 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n14020) );
  INV_X1 U10764 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13989) );
  INV_X1 U10765 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8893) );
  OAI21_X1 U10766 ( .B1(n9320), .B2(n13989), .A(n8893), .ZN(n8897) );
  INV_X1 U10767 ( .A(n9320), .ZN(n8895) );
  AND2_X1 U10768 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8894) );
  INV_X1 U10769 ( .A(n12862), .ZN(n8896) );
  NAND2_X1 U10770 ( .A1(n8897), .A2(n8896), .ZN(n14173) );
  INV_X1 U10771 ( .A(n13152), .ZN(n8903) );
  NAND2_X1 U10772 ( .A1(n8901), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8902) );
  OR2_X1 U10773 ( .A1(n14173), .A2(n9321), .ZN(n8912) );
  INV_X1 U10774 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8909) );
  INV_X1 U10775 ( .A(n8905), .ZN(n12548) );
  INV_X1 U10776 ( .A(n9005), .ZN(n8904) );
  INV_X2 U10777 ( .A(n8904), .ZN(n9230) );
  NAND2_X1 U10778 ( .A1(n9230), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8908) );
  AND2_X2 U10779 ( .A1(n13152), .A2(n8905), .ZN(n9003) );
  NAND2_X1 U10780 ( .A1(n9332), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8907) );
  OAI211_X1 U10781 ( .C1(n8909), .C2(n9637), .A(n8908), .B(n8907), .ZN(n8910)
         );
  INV_X1 U10782 ( .A(n8910), .ZN(n8911) );
  NAND2_X1 U10783 ( .A1(n12586), .A2(n9629), .ZN(n8916) );
  OR2_X1 U10784 ( .A1(n9012), .A2(n12490), .ZN(n8915) );
  XNOR2_X1 U10785 ( .A(n9320), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14181) );
  NAND2_X1 U10786 ( .A1(n14181), .A2(n9331), .ZN(n8922) );
  INV_X1 U10787 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U10788 ( .A1(n9633), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U10789 ( .A1(n9332), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8917) );
  OAI211_X1 U10790 ( .C1(n8919), .C2(n9637), .A(n8918), .B(n8917), .ZN(n8920)
         );
  INV_X1 U10791 ( .A(n8920), .ZN(n8921) );
  INV_X1 U10792 ( .A(n14190), .ZN(n14051) );
  NAND2_X1 U10793 ( .A1(n8949), .A2(n8923), .ZN(n8924) );
  NAND2_X1 U10794 ( .A1(n9174), .A2(n8924), .ZN(n13115) );
  AOI22_X1 U10795 ( .A1(n9633), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9332), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n8926) );
  NAND2_X1 U10796 ( .A1(n9168), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8925) );
  OAI211_X1 U10797 ( .C1(n13115), .C2(n9321), .A(n8926), .B(n8925), .ZN(n14354) );
  INV_X1 U10798 ( .A(n14354), .ZN(n12394) );
  XNOR2_X1 U10799 ( .A(n8928), .B(n8927), .ZN(n12204) );
  NAND2_X1 U10800 ( .A1(n12204), .A2(n9629), .ZN(n8937) );
  AND2_X1 U10801 ( .A1(n8930), .A2(n8929), .ZN(n8942) );
  NAND3_X1 U10802 ( .A1(n9032), .A2(n8942), .A3(n8931), .ZN(n8932) );
  NAND2_X1 U10803 ( .A1(n8932), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8934) );
  MUX2_X1 U10804 ( .A(n8934), .B(P2_IR_REG_31__SCAN_IN), .S(n8933), .Z(n8935)
         );
  AND2_X1 U10805 ( .A1(n9211), .A2(n8935), .ZN(n14127) );
  AOI22_X1 U10806 ( .A1(n9213), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9212), 
        .B2(n14127), .ZN(n8936) );
  INV_X1 U10807 ( .A(n14438), .ZN(n12473) );
  OR2_X1 U10808 ( .A1(n8939), .A2(n8938), .ZN(n8940) );
  NAND2_X1 U10809 ( .A1(n8941), .A2(n8940), .ZN(n12174) );
  NAND2_X1 U10810 ( .A1(n12174), .A2(n9629), .ZN(n8946) );
  AND2_X1 U10811 ( .A1(n9032), .A2(n8942), .ZN(n9143) );
  INV_X1 U10812 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8943) );
  NAND2_X1 U10813 ( .A1(n9143), .A2(n8943), .ZN(n9158) );
  OAI21_X1 U10814 ( .B1(n9160), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8944) );
  XNOR2_X1 U10815 ( .A(n8944), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U10816 ( .A1(n9213), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n14104), 
        .B2(n9212), .ZN(n8945) );
  INV_X1 U10817 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8952) );
  INV_X1 U10818 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U10819 ( .A1(n8955), .A2(n8947), .ZN(n8948) );
  NAND2_X1 U10820 ( .A1(n8949), .A2(n8948), .ZN(n12402) );
  OR2_X1 U10821 ( .A1(n12402), .A2(n9321), .ZN(n8951) );
  AOI22_X1 U10822 ( .A1(n9633), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9332), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n8950) );
  OAI211_X1 U10823 ( .C1(n9637), .C2(n8952), .A(n8951), .B(n8950), .ZN(n14069)
         );
  INV_X1 U10824 ( .A(n14069), .ZN(n9553) );
  INV_X1 U10825 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8960) );
  INV_X1 U10826 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U10827 ( .A1(n9167), .A2(n8953), .ZN(n8954) );
  NAND2_X1 U10828 ( .A1(n8955), .A2(n8954), .ZN(n11954) );
  OR2_X1 U10829 ( .A1(n11954), .A2(n9321), .ZN(n8959) );
  NAND2_X1 U10830 ( .A1(n8906), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U10831 ( .A1(n9230), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8956) );
  AND2_X1 U10832 ( .A1(n8957), .A2(n8956), .ZN(n8958) );
  OAI211_X1 U10833 ( .C1(n9637), .C2(n8960), .A(n8959), .B(n8958), .ZN(n14070)
         );
  INV_X1 U10834 ( .A(n14070), .ZN(n12393) );
  XNOR2_X1 U10835 ( .A(n8962), .B(n8961), .ZN(n12005) );
  NAND2_X1 U10836 ( .A1(n12005), .A2(n9629), .ZN(n8965) );
  NAND2_X1 U10837 ( .A1(n9160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8963) );
  XNOR2_X1 U10838 ( .A(n8963), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U10839 ( .A1(n9213), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9212), 
        .B2(n14084), .ZN(n8964) );
  INV_X1 U10840 ( .A(n12126), .ZN(n9381) );
  NAND2_X1 U10841 ( .A1(n9003), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U10842 ( .A1(n9633), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8970) );
  INV_X1 U10843 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U10844 ( .A1(n9102), .A2(n8966), .ZN(n8967) );
  AND2_X1 U10845 ( .A1(n9119), .A2(n8967), .ZN(n12850) );
  NAND2_X1 U10846 ( .A1(n9331), .A2(n12850), .ZN(n8969) );
  NAND2_X1 U10847 ( .A1(n9168), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8968) );
  NAND4_X1 U10848 ( .A1(n8971), .A2(n8970), .A3(n8969), .A4(n8968), .ZN(n14074) );
  XNOR2_X1 U10849 ( .A(n8973), .B(n8972), .ZN(n11582) );
  NAND2_X1 U10850 ( .A1(n11582), .A2(n9629), .ZN(n8980) );
  INV_X1 U10851 ( .A(n9032), .ZN(n9037) );
  INV_X1 U10852 ( .A(n9068), .ZN(n8975) );
  NAND2_X1 U10853 ( .A1(n8975), .A2(n8974), .ZN(n9083) );
  INV_X1 U10854 ( .A(n9083), .ZN(n8977) );
  INV_X1 U10855 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8976) );
  NAND2_X1 U10856 ( .A1(n8977), .A2(n8976), .ZN(n9096) );
  NAND2_X1 U10857 ( .A1(n8978), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9114) );
  XNOR2_X1 U10858 ( .A(n9114), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U10859 ( .A1(n11529), .A2(n9212), .B1(n9213), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U10860 ( .A1(n9003), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U10861 ( .A1(n9004), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8983) );
  NAND3_X2 U10862 ( .A1(n8134), .A2(n8984), .A3(n8983), .ZN(n9000) );
  XNOR2_X1 U10863 ( .A(n8987), .B(n8986), .ZN(n8989) );
  MUX2_X1 U10864 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n10304), .Z(n8988) );
  XNOR2_X1 U10865 ( .A(n8989), .B(n8988), .ZN(n10306) );
  OR2_X1 U10866 ( .A1(n9643), .A2(n10306), .ZN(n8991) );
  OR2_X1 U10867 ( .A1(n9012), .A2(n10048), .ZN(n8990) );
  NAND2_X1 U10868 ( .A1(n9003), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U10869 ( .A1(n9005), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U10870 ( .A1(n10316), .A2(SI_0_), .ZN(n8997) );
  NAND2_X1 U10871 ( .A1(n8997), .A2(n8996), .ZN(n8999) );
  AND2_X1 U10872 ( .A1(n8999), .A2(n8998), .ZN(n14480) );
  MUX2_X1 U10873 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14480), .S(n10226), .Z(n11403) );
  NAND2_X1 U10874 ( .A1(n9450), .A2(n11403), .ZN(n13125) );
  INV_X1 U10875 ( .A(n9000), .ZN(n9363) );
  INV_X1 U10876 ( .A(n11213), .ZN(n13127) );
  NAND2_X1 U10877 ( .A1(n9363), .A2(n13127), .ZN(n9002) );
  NAND2_X1 U10878 ( .A1(n10487), .A2(n9002), .ZN(n10448) );
  NAND2_X1 U10879 ( .A1(n9003), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U10880 ( .A1(n9004), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U10881 ( .A1(n9042), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U10882 ( .A1(n9005), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9006) );
  NAND4_X1 U10883 ( .A1(n9009), .A2(n9008), .A3(n9007), .A4(n9006), .ZN(n14081) );
  OR2_X1 U10884 ( .A1(n10324), .A2(n9643), .ZN(n9018) );
  OR2_X1 U10885 ( .A1(n9012), .A2(n10049), .ZN(n9017) );
  NAND2_X1 U10886 ( .A1(n9013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9015) );
  MUX2_X1 U10887 ( .A(n9015), .B(P2_IR_REG_31__SCAN_IN), .S(n9014), .Z(n9016)
         );
  NAND2_X1 U10888 ( .A1(n9016), .A2(n9029), .ZN(n10260) );
  NAND2_X1 U10889 ( .A1(n10448), .A2(n10447), .ZN(n10446) );
  INV_X1 U10890 ( .A(n14081), .ZN(n13128) );
  NAND2_X1 U10891 ( .A1(n13128), .A2(n9019), .ZN(n9020) );
  NAND2_X1 U10892 ( .A1(n10446), .A2(n9020), .ZN(n10536) );
  NAND2_X1 U10893 ( .A1(n8906), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9025) );
  INV_X1 U10894 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9021) );
  NAND2_X1 U10895 ( .A1(n9004), .A2(n9021), .ZN(n9024) );
  NAND2_X1 U10896 ( .A1(n9168), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U10897 ( .A1(n9230), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U10898 ( .A1(n10065), .A2(n9028), .ZN(n9034) );
  NAND2_X1 U10899 ( .A1(n9029), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9030) );
  INV_X1 U10900 ( .A(n9031), .ZN(n9033) );
  XNOR2_X1 U10901 ( .A(n14080), .B(n11189), .ZN(n10537) );
  INV_X1 U10902 ( .A(n14080), .ZN(n10845) );
  NAND2_X1 U10903 ( .A1(n10845), .A2(n11189), .ZN(n9035) );
  NAND2_X1 U10904 ( .A1(n10535), .A2(n9035), .ZN(n10439) );
  NAND2_X1 U10905 ( .A1(n10806), .A2(n9028), .ZN(n9041) );
  NAND2_X1 U10906 ( .A1(n9037), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9038) );
  MUX2_X1 U10907 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9038), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9039) );
  AND2_X1 U10908 ( .A1(n9039), .A2(n9053), .ZN(n10868) );
  AOI22_X1 U10909 ( .A1(n9213), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9212), .B2(
        n10868), .ZN(n9040) );
  NAND2_X1 U10910 ( .A1(n9230), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U10911 ( .A1(n9003), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9045) );
  OAI21_X1 U10912 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9058), .ZN(n10854) );
  INV_X1 U10913 ( .A(n10854), .ZN(n11473) );
  NAND2_X1 U10914 ( .A1(n9004), .A2(n11473), .ZN(n9044) );
  NAND2_X1 U10915 ( .A1(n9042), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U10916 ( .A1(n10439), .A2(n10441), .ZN(n10438) );
  OR2_X1 U10917 ( .A1(n14079), .A2(n11474), .ZN(n9047) );
  NAND2_X1 U10918 ( .A1(n9036), .A2(n9048), .ZN(n9050) );
  NAND2_X1 U10919 ( .A1(n9050), .A2(n9049), .ZN(n9052) );
  XNOR2_X1 U10920 ( .A(n9052), .B(n9051), .ZN(n10817) );
  NAND2_X1 U10921 ( .A1(n10817), .A2(n9629), .ZN(n9056) );
  NAND2_X1 U10922 ( .A1(n9053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9054) );
  XNOR2_X1 U10923 ( .A(n9054), .B(P2_IR_REG_5__SCAN_IN), .ZN(n15535) );
  AOI22_X1 U10924 ( .A1(n9213), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9212), .B2(
        n15535), .ZN(n9055) );
  NAND2_X1 U10925 ( .A1(n9056), .A2(n9055), .ZN(n10947) );
  INV_X1 U10926 ( .A(n10947), .ZN(n11367) );
  NAND2_X1 U10927 ( .A1(n9003), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9063) );
  NAND2_X1 U10928 ( .A1(n9230), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9062) );
  INV_X1 U10929 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U10930 ( .A1(n9058), .A2(n9057), .ZN(n9059) );
  AND2_X1 U10931 ( .A1(n9073), .A2(n9059), .ZN(n11363) );
  NAND2_X1 U10932 ( .A1(n9331), .A2(n11363), .ZN(n9061) );
  NAND2_X1 U10933 ( .A1(n9168), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9060) );
  NAND4_X1 U10934 ( .A1(n9063), .A2(n9062), .A3(n9061), .A4(n9060), .ZN(n14078) );
  INV_X1 U10935 ( .A(n14078), .ZN(n11013) );
  OAI21_X1 U10936 ( .B1(n10776), .B2(n11367), .A(n11013), .ZN(n9065) );
  NAND2_X1 U10937 ( .A1(n10776), .A2(n11367), .ZN(n9064) );
  NAND2_X1 U10938 ( .A1(n9065), .A2(n9064), .ZN(n11454) );
  XNOR2_X1 U10939 ( .A(n9066), .B(n9067), .ZN(n11028) );
  NAND2_X1 U10940 ( .A1(n11028), .A2(n9629), .ZN(n9071) );
  NAND2_X1 U10941 ( .A1(n9068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9069) );
  XNOR2_X1 U10942 ( .A(n9069), .B(P2_IR_REG_6__SCAN_IN), .ZN(n15546) );
  AOI22_X1 U10943 ( .A1(n9213), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9212), .B2(
        n15546), .ZN(n9070) );
  NAND2_X1 U10944 ( .A1(n9071), .A2(n9070), .ZN(n11455) );
  NAND2_X1 U10945 ( .A1(n9230), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U10946 ( .A1(n8906), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9077) );
  INV_X1 U10947 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U10948 ( .A1(n9073), .A2(n9072), .ZN(n9074) );
  AND2_X1 U10949 ( .A1(n9087), .A2(n9074), .ZN(n11460) );
  NAND2_X1 U10950 ( .A1(n9331), .A2(n11460), .ZN(n9076) );
  NAND2_X1 U10951 ( .A1(n9168), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9075) );
  NAND4_X1 U10952 ( .A1(n9078), .A2(n9077), .A3(n9076), .A4(n9075), .ZN(n14077) );
  INV_X1 U10953 ( .A(n14077), .ZN(n11092) );
  NAND2_X1 U10954 ( .A1(n11455), .A2(n11092), .ZN(n9375) );
  OR2_X1 U10955 ( .A1(n11455), .A2(n11092), .ZN(n9079) );
  NAND2_X1 U10956 ( .A1(n9375), .A2(n9079), .ZN(n11463) );
  OR2_X1 U10957 ( .A1(n11455), .A2(n14077), .ZN(n9080) );
  NAND2_X1 U10958 ( .A1(n9083), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9084) );
  XNOR2_X1 U10959 ( .A(n9084), .B(P2_IR_REG_7__SCAN_IN), .ZN(n15557) );
  AOI22_X1 U10960 ( .A1(n9213), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9212), .B2(
        n15557), .ZN(n9085) );
  NAND2_X1 U10961 ( .A1(n8906), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U10962 ( .A1(n9168), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9091) );
  INV_X1 U10963 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U10964 ( .A1(n9087), .A2(n9086), .ZN(n9088) );
  AND2_X1 U10965 ( .A1(n9100), .A2(n9088), .ZN(n11198) );
  NAND2_X1 U10966 ( .A1(n9331), .A2(n11198), .ZN(n9090) );
  NAND2_X1 U10967 ( .A1(n9230), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9089) );
  NAND4_X1 U10968 ( .A1(n9092), .A2(n9091), .A3(n9090), .A4(n9089), .ZN(n14076) );
  NAND2_X1 U10969 ( .A1(n15840), .A2(n14076), .ZN(n11384) );
  NAND2_X1 U10970 ( .A1(n11274), .A2(n9629), .ZN(n9099) );
  NAND2_X1 U10971 ( .A1(n9096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9097) );
  XNOR2_X1 U10972 ( .A(n9097), .B(P2_IR_REG_8__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U10973 ( .A1(n9213), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11110), 
        .B2(n9212), .ZN(n9098) );
  NAND2_X1 U10974 ( .A1(n9230), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9106) );
  NAND2_X1 U10975 ( .A1(n8906), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U10976 ( .A1(n9100), .A2(n10963), .ZN(n9101) );
  AND2_X1 U10977 ( .A1(n9102), .A2(n9101), .ZN(n11381) );
  NAND2_X1 U10978 ( .A1(n9331), .A2(n11381), .ZN(n9104) );
  NAND2_X1 U10979 ( .A1(n9168), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9103) );
  NAND4_X1 U10980 ( .A1(n9106), .A2(n9105), .A3(n9104), .A4(n9103), .ZN(n14075) );
  NAND2_X1 U10981 ( .A1(n11389), .A2(n14075), .ZN(n9108) );
  AND2_X1 U10982 ( .A1(n11384), .A2(n9108), .ZN(n9107) );
  NAND2_X1 U10983 ( .A1(n15838), .A2(n9107), .ZN(n11341) );
  INV_X1 U10984 ( .A(n9108), .ZN(n9109) );
  XNOR2_X1 U10985 ( .A(n11389), .B(n14075), .ZN(n9701) );
  OR2_X1 U10986 ( .A1(n9109), .A2(n11386), .ZN(n11340) );
  INV_X1 U10987 ( .A(n14074), .ZN(n12795) );
  INV_X1 U10988 ( .A(n9125), .ZN(n11352) );
  NAND2_X1 U10989 ( .A1(n11587), .A2(n9629), .ZN(n9117) );
  NAND2_X1 U10990 ( .A1(n9114), .A2(n9113), .ZN(n9115) );
  NAND2_X1 U10991 ( .A1(n9115), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9130) );
  XNOR2_X1 U10992 ( .A(n9130), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15597) );
  AOI22_X1 U10993 ( .A1(n15597), .A2(n9212), .B1(n9213), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U10994 ( .A1(n8906), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U10995 ( .A1(n9168), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9123) );
  NAND2_X1 U10996 ( .A1(n9119), .A2(n9118), .ZN(n9120) );
  AND2_X1 U10997 ( .A1(n9135), .A2(n9120), .ZN(n12793) );
  NAND2_X1 U10998 ( .A1(n9331), .A2(n12793), .ZN(n9122) );
  NAND2_X1 U10999 ( .A1(n9230), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9121) );
  NAND4_X1 U11000 ( .A1(n9124), .A2(n9123), .A3(n9122), .A4(n9121), .ZN(n14073) );
  OAI21_X1 U11001 ( .B1(n11352), .B2(n12797), .A(n14073), .ZN(n9126) );
  NAND2_X1 U11002 ( .A1(n9130), .A2(n9129), .ZN(n9131) );
  NAND2_X1 U11003 ( .A1(n9131), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9132) );
  AOI22_X1 U11004 ( .A1(n12100), .A2(n9212), .B1(n9213), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n9133) );
  NAND2_X1 U11005 ( .A1(n9633), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9140) );
  NAND2_X1 U11006 ( .A1(n8906), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9139) );
  INV_X1 U11007 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9134) );
  NAND2_X1 U11008 ( .A1(n9135), .A2(n9134), .ZN(n9136) );
  AND2_X1 U11009 ( .A1(n9150), .A2(n9136), .ZN(n11870) );
  NAND2_X1 U11010 ( .A1(n9331), .A2(n11870), .ZN(n9138) );
  NAND2_X1 U11011 ( .A1(n9168), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9137) );
  NAND4_X1 U11012 ( .A1(n9140), .A2(n9139), .A3(n9138), .A4(n9137), .ZN(n14072) );
  INV_X1 U11013 ( .A(n14072), .ZN(n12794) );
  XNOR2_X1 U11014 ( .A(n11879), .B(n12794), .ZN(n11507) );
  AND2_X1 U11015 ( .A1(n11879), .A2(n14072), .ZN(n9141) );
  XNOR2_X1 U11016 ( .A(n9142), .B(n8146), .ZN(n11965) );
  NAND2_X1 U11017 ( .A1(n11965), .A2(n9629), .ZN(n9148) );
  INV_X1 U11018 ( .A(n9143), .ZN(n9144) );
  NAND2_X1 U11019 ( .A1(n9144), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9145) );
  MUX2_X1 U11020 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9145), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9146) );
  NAND2_X1 U11021 ( .A1(n9146), .A2(n9158), .ZN(n15574) );
  INV_X1 U11022 ( .A(n15574), .ZN(n12103) );
  AOI22_X1 U11023 ( .A1(n9213), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9212), 
        .B2(n12103), .ZN(n9147) );
  NAND2_X1 U11024 ( .A1(n9230), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9155) );
  NAND2_X1 U11025 ( .A1(n8906), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9154) );
  NAND2_X1 U11026 ( .A1(n9150), .A2(n9149), .ZN(n9151) );
  AND2_X1 U11027 ( .A1(n9165), .A2(n9151), .ZN(n13140) );
  NAND2_X1 U11028 ( .A1(n9331), .A2(n13140), .ZN(n9153) );
  NAND2_X1 U11029 ( .A1(n9168), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9152) );
  NAND4_X1 U11030 ( .A1(n9155), .A2(n9154), .A3(n9153), .A4(n9152), .ZN(n14071) );
  XNOR2_X1 U11031 ( .A(n11881), .B(n14071), .ZN(n11841) );
  INV_X1 U11032 ( .A(n14071), .ZN(n9530) );
  INV_X1 U11033 ( .A(n11881), .ZN(n13145) );
  XNOR2_X1 U11034 ( .A(n9157), .B(n9156), .ZN(n11971) );
  NAND2_X1 U11035 ( .A1(n11971), .A2(n9629), .ZN(n9163) );
  NAND2_X1 U11036 ( .A1(n9158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9159) );
  MUX2_X1 U11037 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9159), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9161) );
  AOI22_X1 U11038 ( .A1(n9213), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9212), 
        .B2(n12367), .ZN(n9162) );
  NAND2_X1 U11039 ( .A1(n9165), .A2(n9164), .ZN(n9166) );
  AND2_X1 U11040 ( .A1(n9167), .A2(n9166), .ZN(n12060) );
  NAND2_X1 U11041 ( .A1(n12060), .A2(n9331), .ZN(n9172) );
  NAND2_X1 U11042 ( .A1(n9230), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9171) );
  NAND2_X1 U11043 ( .A1(n8906), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U11044 ( .A1(n9168), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9169) );
  NAND4_X1 U11045 ( .A1(n9172), .A2(n9171), .A3(n9170), .A4(n9169), .ZN(n13141) );
  XNOR2_X1 U11046 ( .A(n12134), .B(n13141), .ZN(n12052) );
  INV_X1 U11047 ( .A(n12134), .ZN(n12062) );
  INV_X1 U11048 ( .A(n13141), .ZN(n9379) );
  XNOR2_X1 U11049 ( .A(n12126), .B(n12393), .ZN(n11951) );
  XNOR2_X1 U11050 ( .A(n14444), .B(n14069), .ZN(n12396) );
  XNOR2_X1 U11051 ( .A(n14438), .B(n12394), .ZN(n12475) );
  INV_X1 U11052 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U11053 ( .A1(n9174), .A2(n9173), .ZN(n9175) );
  NAND2_X1 U11054 ( .A1(n9192), .A2(n9175), .ZN(n14344) );
  OR2_X1 U11055 ( .A1(n14344), .A2(n9321), .ZN(n9181) );
  INV_X1 U11056 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U11057 ( .A1(n9332), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U11058 ( .A1(n9168), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9176) );
  OAI211_X1 U11059 ( .C1(n9178), .C2(n8904), .A(n9177), .B(n9176), .ZN(n9179)
         );
  INV_X1 U11060 ( .A(n9179), .ZN(n9180) );
  NAND2_X1 U11061 ( .A1(n9181), .A2(n9180), .ZN(n14068) );
  XNOR2_X1 U11062 ( .A(n9183), .B(n9182), .ZN(n12330) );
  NAND2_X1 U11063 ( .A1(n12330), .A2(n9629), .ZN(n9186) );
  NAND2_X1 U11064 ( .A1(n9211), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9184) );
  XNOR2_X1 U11065 ( .A(n9184), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15567) );
  AOI22_X1 U11066 ( .A1(n9213), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9212), 
        .B2(n15567), .ZN(n9185) );
  XOR2_X1 U11067 ( .A(n14068), .B(n14433), .Z(n14338) );
  INV_X1 U11068 ( .A(n14338), .ZN(n14351) );
  XNOR2_X1 U11069 ( .A(n9201), .B(n9202), .ZN(n12591) );
  NAND2_X1 U11070 ( .A1(n12591), .A2(n9629), .ZN(n9190) );
  NAND2_X1 U11071 ( .A1(n9355), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9188) );
  XNOR2_X1 U11072 ( .A(n9188), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U11073 ( .A1(n9213), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9212), 
        .B2(n14122), .ZN(n9189) );
  NAND2_X1 U11074 ( .A1(n9192), .A2(n9191), .ZN(n9193) );
  AND2_X1 U11075 ( .A1(n9217), .A2(n9193), .ZN(n14330) );
  NAND2_X1 U11076 ( .A1(n14330), .A2(n9331), .ZN(n9199) );
  INV_X1 U11077 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U11078 ( .A1(n9332), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U11079 ( .A1(n9230), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9194) );
  OAI211_X1 U11080 ( .C1(n9637), .C2(n9196), .A(n9195), .B(n9194), .ZN(n9197)
         );
  INV_X1 U11081 ( .A(n9197), .ZN(n9198) );
  XNOR2_X1 U11082 ( .A(n14428), .B(n14356), .ZN(n14318) );
  INV_X1 U11083 ( .A(n14318), .ZN(n14324) );
  INV_X1 U11084 ( .A(n9201), .ZN(n9203) );
  NAND2_X1 U11085 ( .A1(n9203), .A2(n9202), .ZN(n9206) );
  OR2_X1 U11086 ( .A1(n9204), .A2(n13291), .ZN(n9205) );
  NAND2_X1 U11087 ( .A1(n9206), .A2(n9205), .ZN(n9210) );
  NAND2_X1 U11088 ( .A1(n9208), .A2(n9207), .ZN(n9209) );
  NAND2_X1 U11089 ( .A1(n12595), .A2(n9629), .ZN(n9215) );
  AOI22_X1 U11090 ( .A1(n9213), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9212), 
        .B2(n14140), .ZN(n9214) );
  NAND2_X2 U11091 ( .A1(n9215), .A2(n9214), .ZN(n14424) );
  INV_X1 U11092 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U11093 ( .A1(n9217), .A2(n9216), .ZN(n9218) );
  NAND2_X1 U11094 ( .A1(n9243), .A2(n9218), .ZN(n14309) );
  OR2_X1 U11095 ( .A1(n14309), .A2(n9321), .ZN(n9223) );
  INV_X1 U11096 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U11097 ( .A1(n9168), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11098 ( .A1(n9332), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9219) );
  OAI211_X1 U11099 ( .C1(n8904), .C2(n14310), .A(n9220), .B(n9219), .ZN(n9221)
         );
  INV_X1 U11100 ( .A(n9221), .ZN(n9222) );
  NAND2_X1 U11101 ( .A1(n9223), .A2(n9222), .ZN(n14067) );
  XNOR2_X1 U11102 ( .A(n14424), .B(n9224), .ZN(n14300) );
  NAND2_X1 U11103 ( .A1(n7585), .A2(n9224), .ZN(n9225) );
  XNOR2_X1 U11104 ( .A(n9227), .B(n9226), .ZN(n12608) );
  NAND2_X1 U11105 ( .A1(n12608), .A2(n9629), .ZN(n9229) );
  OR2_X1 U11106 ( .A1(n9012), .A2(n11869), .ZN(n9228) );
  XNOR2_X1 U11107 ( .A(n9243), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n14287) );
  NAND2_X1 U11108 ( .A1(n14287), .A2(n9331), .ZN(n9236) );
  INV_X1 U11109 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U11110 ( .A1(n9230), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U11111 ( .A1(n9332), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9231) );
  OAI211_X1 U11112 ( .C1(n9233), .C2(n9637), .A(n9232), .B(n9231), .ZN(n9234)
         );
  INV_X1 U11113 ( .A(n9234), .ZN(n9235) );
  INV_X1 U11114 ( .A(n14418), .ZN(n14290) );
  INV_X1 U11115 ( .A(n14066), .ZN(n14302) );
  XNOR2_X1 U11116 ( .A(n9238), .B(n9237), .ZN(n12621) );
  NAND2_X1 U11117 ( .A1(n12621), .A2(n9629), .ZN(n9240) );
  OR2_X1 U11118 ( .A1(n9012), .A2(n11863), .ZN(n9239) );
  INV_X1 U11119 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9242) );
  INV_X1 U11120 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9241) );
  OAI21_X1 U11121 ( .B1(n9243), .B2(n9242), .A(n9241), .ZN(n9244) );
  NAND2_X1 U11122 ( .A1(n9244), .A2(n9260), .ZN(n14269) );
  OR2_X1 U11123 ( .A1(n14269), .A2(n9321), .ZN(n9250) );
  INV_X1 U11124 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U11125 ( .A1(n9332), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U11126 ( .A1(n9633), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9245) );
  OAI211_X1 U11127 ( .C1(n9247), .C2(n9637), .A(n9246), .B(n9245), .ZN(n9248)
         );
  INV_X1 U11128 ( .A(n9248), .ZN(n9249) );
  INV_X1 U11129 ( .A(n14251), .ZN(n12505) );
  NAND2_X1 U11130 ( .A1(n12639), .A2(n9253), .ZN(n9270) );
  INV_X1 U11131 ( .A(n12639), .ZN(n9255) );
  NAND2_X1 U11132 ( .A1(n9255), .A2(n9254), .ZN(n9256) );
  NAND2_X1 U11133 ( .A1(n9270), .A2(n9256), .ZN(n12144) );
  OR2_X1 U11134 ( .A1(n12144), .A2(n9643), .ZN(n9258) );
  OR2_X1 U11135 ( .A1(n9012), .A2(n12146), .ZN(n9257) );
  NAND2_X2 U11136 ( .A1(n9258), .A2(n9257), .ZN(n14407) );
  INV_X1 U11137 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9259) );
  NAND2_X1 U11138 ( .A1(n9260), .A2(n9259), .ZN(n9261) );
  NAND2_X1 U11139 ( .A1(n9276), .A2(n9261), .ZN(n13097) );
  OR2_X1 U11140 ( .A1(n13097), .A2(n9321), .ZN(n9267) );
  INV_X1 U11141 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U11142 ( .A1(n9633), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9263) );
  NAND2_X1 U11143 ( .A1(n9332), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9262) );
  OAI211_X1 U11144 ( .C1(n9264), .C2(n9637), .A(n9263), .B(n9262), .ZN(n9265)
         );
  INV_X1 U11145 ( .A(n9265), .ZN(n9266) );
  XNOR2_X1 U11146 ( .A(n14407), .B(n14065), .ZN(n9708) );
  NAND2_X1 U11147 ( .A1(n9268), .A2(SI_22_), .ZN(n9269) );
  NAND2_X1 U11148 ( .A1(n9270), .A2(n9269), .ZN(n9273) );
  XNOR2_X1 U11149 ( .A(n9271), .B(SI_23_), .ZN(n9272) );
  NAND2_X1 U11150 ( .A1(n12650), .A2(n9629), .ZN(n9275) );
  OR2_X1 U11151 ( .A1(n9012), .A2(n10754), .ZN(n9274) );
  INV_X1 U11152 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14001) );
  NAND2_X1 U11153 ( .A1(n9276), .A2(n14001), .ZN(n9277) );
  NAND2_X1 U11154 ( .A1(n9290), .A2(n9277), .ZN(n13999) );
  OR2_X1 U11155 ( .A1(n13999), .A2(n9321), .ZN(n9283) );
  INV_X1 U11156 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9280) );
  NAND2_X1 U11157 ( .A1(n9332), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U11158 ( .A1(n9633), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9278) );
  OAI211_X1 U11159 ( .C1(n9637), .C2(n9280), .A(n9279), .B(n9278), .ZN(n9281)
         );
  INV_X1 U11160 ( .A(n9281), .ZN(n9282) );
  XNOR2_X1 U11161 ( .A(n14403), .B(n14032), .ZN(n14241) );
  NAND2_X1 U11162 ( .A1(n14240), .A2(n9284), .ZN(n14217) );
  XNOR2_X1 U11163 ( .A(n9285), .B(SI_24_), .ZN(n9286) );
  XNOR2_X1 U11164 ( .A(n9287), .B(n9286), .ZN(n12654) );
  NAND2_X1 U11165 ( .A1(n12654), .A2(n9629), .ZN(n9289) );
  INV_X1 U11166 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12160) );
  OR2_X1 U11167 ( .A1(n9012), .A2(n12160), .ZN(n9288) );
  NAND2_X1 U11168 ( .A1(n9290), .A2(n14029), .ZN(n9291) );
  NAND2_X1 U11169 ( .A1(n9304), .A2(n9291), .ZN(n14226) );
  OR2_X1 U11170 ( .A1(n14226), .A2(n9321), .ZN(n9297) );
  INV_X1 U11171 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9294) );
  NAND2_X1 U11172 ( .A1(n9633), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11173 ( .A1(n9332), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9292) );
  OAI211_X1 U11174 ( .C1(n9294), .C2(n9637), .A(n9293), .B(n9292), .ZN(n9295)
         );
  INV_X1 U11175 ( .A(n9295), .ZN(n9296) );
  XNOR2_X1 U11176 ( .A(n14396), .B(n14018), .ZN(n14220) );
  NAND2_X1 U11177 ( .A1(n14216), .A2(n9298), .ZN(n14206) );
  XNOR2_X1 U11178 ( .A(n9300), .B(n9299), .ZN(n12669) );
  NAND2_X1 U11179 ( .A1(n12669), .A2(n9629), .ZN(n9302) );
  OR2_X1 U11180 ( .A1(n9012), .A2(n12162), .ZN(n9301) );
  INV_X1 U11181 ( .A(n9303), .ZN(n9318) );
  NAND2_X1 U11182 ( .A1(n9304), .A2(n14020), .ZN(n9305) );
  NAND2_X1 U11183 ( .A1(n14210), .A2(n9331), .ZN(n9311) );
  INV_X1 U11184 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U11185 ( .A1(n9633), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U11186 ( .A1(n9332), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n9306) );
  OAI211_X1 U11187 ( .C1(n9308), .C2(n9637), .A(n9307), .B(n9306), .ZN(n9309)
         );
  INV_X1 U11188 ( .A(n9309), .ZN(n9310) );
  XNOR2_X1 U11189 ( .A(n14392), .B(n14221), .ZN(n9709) );
  XNOR2_X1 U11190 ( .A(n9314), .B(n9313), .ZN(n12681) );
  NAND2_X1 U11191 ( .A1(n12681), .A2(n9629), .ZN(n9316) );
  OR2_X1 U11192 ( .A1(n9012), .A2(n12389), .ZN(n9315) );
  INV_X1 U11193 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11194 ( .A1(n9318), .A2(n9317), .ZN(n9319) );
  NAND2_X1 U11195 ( .A1(n9320), .A2(n9319), .ZN(n14045) );
  INV_X1 U11196 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U11197 ( .A1(n9633), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U11198 ( .A1(n9332), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9322) );
  OAI211_X1 U11199 ( .C1(n9324), .C2(n9637), .A(n9323), .B(n9322), .ZN(n9325)
         );
  INV_X1 U11200 ( .A(n9325), .ZN(n9326) );
  NAND2_X1 U11201 ( .A1(n14386), .A2(n14063), .ZN(n9329) );
  XOR2_X1 U11202 ( .A(n14190), .B(n14377), .Z(n14185) );
  NAND2_X1 U11203 ( .A1(n14373), .A2(n13988), .ZN(n9330) );
  NAND2_X1 U11204 ( .A1(n9394), .A2(n9330), .ZN(n12836) );
  NAND2_X1 U11205 ( .A1(n12862), .A2(n9331), .ZN(n9338) );
  INV_X1 U11206 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9335) );
  NAND2_X1 U11207 ( .A1(n9633), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U11208 ( .A1(n9332), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9333) );
  OAI211_X1 U11209 ( .C1(n9335), .C2(n9637), .A(n9334), .B(n9333), .ZN(n9336)
         );
  INV_X1 U11210 ( .A(n9336), .ZN(n9337) );
  NAND2_X1 U11211 ( .A1(n9338), .A2(n9337), .ZN(n14061) );
  INV_X1 U11212 ( .A(n14061), .ZN(n9344) );
  MUX2_X1 U11213 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n10316), .Z(n9623) );
  XNOR2_X1 U11214 ( .A(n9623), .B(n13977), .ZN(n9621) );
  NAND2_X1 U11215 ( .A1(n14945), .A2(n9629), .ZN(n9343) );
  OR2_X1 U11216 ( .A1(n9012), .A2(n12547), .ZN(n9342) );
  XOR2_X1 U11217 ( .A(n9344), .B(n12860), .Z(n9712) );
  INV_X1 U11218 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9345) );
  AOI21_X1 U11219 ( .B1(n9346), .B2(n9345), .A(n8875), .ZN(n9351) );
  NAND2_X1 U11220 ( .A1(n9356), .A2(n9353), .ZN(n9349) );
  INV_X1 U11221 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9350) );
  MUX2_X2 U11222 ( .A(n9351), .B(n9352), .S(n9350), .Z(n11868) );
  XNOR2_X2 U11223 ( .A(n9352), .B(P2_IR_REG_21__SCAN_IN), .ZN(n9720) );
  INV_X1 U11224 ( .A(n9355), .ZN(n9356) );
  NAND2_X1 U11225 ( .A1(n9357), .A2(n9356), .ZN(n9419) );
  XNOR2_X1 U11226 ( .A(n11173), .B(n9726), .ZN(n9360) );
  NAND2_X1 U11227 ( .A1(n10019), .A2(n14449), .ZN(n15860) );
  NAND2_X1 U11228 ( .A1(n12867), .A2(n15860), .ZN(n9410) );
  INV_X1 U11229 ( .A(n14428), .ZN(n14333) );
  INV_X1 U11230 ( .A(n14433), .ZN(n14350) );
  NOR2_X1 U11231 ( .A1(n9450), .A2(n10885), .ZN(n10491) );
  NAND2_X1 U11232 ( .A1(n9362), .A2(n10491), .ZN(n10490) );
  NAND2_X1 U11233 ( .A1(n9363), .A2(n11213), .ZN(n9364) );
  NAND2_X1 U11234 ( .A1(n10490), .A2(n9364), .ZN(n10451) );
  NAND2_X1 U11235 ( .A1(n10451), .A2(n10450), .ZN(n9366) );
  NAND2_X1 U11236 ( .A1(n13128), .A2(n11081), .ZN(n9365) );
  INV_X1 U11237 ( .A(n10537), .ZN(n9367) );
  NAND2_X1 U11238 ( .A1(n10538), .A2(n9367), .ZN(n9369) );
  NAND2_X1 U11239 ( .A1(n10845), .A2(n9464), .ZN(n9368) );
  INV_X1 U11240 ( .A(n10441), .ZN(n9370) );
  NAND2_X1 U11241 ( .A1(n10442), .A2(n9370), .ZN(n9372) );
  NAND2_X1 U11242 ( .A1(n11474), .A2(n11064), .ZN(n9371) );
  AND2_X1 U11243 ( .A1(n10947), .A2(n11013), .ZN(n9373) );
  OR2_X1 U11244 ( .A1(n10947), .A2(n11013), .ZN(n9374) );
  INV_X1 U11245 ( .A(n14076), .ZN(n11011) );
  OR2_X1 U11246 ( .A1(n15840), .A2(n11011), .ZN(n9377) );
  AND2_X1 U11247 ( .A1(n15840), .A2(n11011), .ZN(n9376) );
  INV_X1 U11248 ( .A(n14075), .ZN(n12852) );
  NAND2_X1 U11249 ( .A1(n11389), .A2(n12852), .ZN(n9378) );
  INV_X1 U11250 ( .A(n11389), .ZN(n15857) );
  INV_X1 U11251 ( .A(n14073), .ZN(n12851) );
  INV_X1 U11252 ( .A(n11507), .ZN(n11512) );
  OAI21_X1 U11253 ( .B1(n9530), .B2(n11881), .A(n11840), .ZN(n12053) );
  NAND2_X1 U11254 ( .A1(n12053), .A2(n12052), .ZN(n12051) );
  NAND2_X1 U11255 ( .A1(n12051), .A2(n9380), .ZN(n11948) );
  NAND2_X1 U11256 ( .A1(n11948), .A2(n8144), .ZN(n9382) );
  NAND2_X1 U11257 ( .A1(n12468), .A2(n9383), .ZN(n9384) );
  INV_X1 U11258 ( .A(n14068), .ZN(n14321) );
  NAND2_X1 U11259 ( .A1(n14290), .A2(n14066), .ZN(n9386) );
  OAI21_X1 U11260 ( .B1(n12505), .B2(n14413), .A(n9387), .ZN(n14250) );
  INV_X1 U11261 ( .A(n14407), .ZN(n14257) );
  INV_X1 U11262 ( .A(n14065), .ZN(n14009) );
  INV_X1 U11263 ( .A(n14241), .ZN(n14236) );
  INV_X1 U11264 ( .A(n14392), .ZN(n14213) );
  XNOR2_X1 U11265 ( .A(n14386), .B(n14063), .ZN(n14195) );
  NAND2_X1 U11266 ( .A1(n14189), .A2(n14195), .ZN(n9393) );
  NAND2_X1 U11267 ( .A1(n14386), .A2(n14019), .ZN(n9392) );
  INV_X1 U11268 ( .A(n14185), .ZN(n14177) );
  INV_X1 U11269 ( .A(n9712), .ZN(n9395) );
  INV_X1 U11270 ( .A(n11868), .ZN(n10009) );
  NAND2_X1 U11271 ( .A1(n10009), .A2(n9720), .ZN(n9396) );
  NAND2_X1 U11272 ( .A1(n9726), .A2(n14140), .ZN(n9647) );
  INV_X2 U11273 ( .A(n14298), .ZN(n14358) );
  INV_X1 U11274 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9399) );
  NAND2_X1 U11275 ( .A1(n9633), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9398) );
  NAND2_X1 U11276 ( .A1(n9332), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9397) );
  OAI211_X1 U11277 ( .C1(n9637), .C2(n9399), .A(n9398), .B(n9397), .ZN(n14060)
         );
  INV_X1 U11278 ( .A(n14060), .ZN(n9650) );
  NAND2_X1 U11279 ( .A1(n9726), .A2(n9720), .ZN(n9437) );
  INV_X1 U11280 ( .A(n9400), .ZN(n9401) );
  INV_X1 U11281 ( .A(n12489), .ZN(n10238) );
  NAND2_X1 U11282 ( .A1(n10238), .A2(P2_B_REG_SCAN_IN), .ZN(n9402) );
  NAND2_X1 U11283 ( .A1(n14355), .A2(n9402), .ZN(n14152) );
  NAND2_X1 U11284 ( .A1(n14062), .A2(n14353), .ZN(n9403) );
  OAI21_X1 U11285 ( .B1(n9650), .B2(n14152), .A(n9403), .ZN(n9404) );
  NAND2_X1 U11286 ( .A1(n13127), .A2(n10885), .ZN(n10495) );
  INV_X1 U11287 ( .A(n11474), .ZN(n10855) );
  NOR2_X2 U11288 ( .A1(n11456), .A2(n11455), .ZN(n11457) );
  INV_X1 U11289 ( .A(n15840), .ZN(n11200) );
  AND2_X1 U11290 ( .A1(n11457), .A2(n11200), .ZN(n11383) );
  NAND2_X1 U11291 ( .A1(n11383), .A2(n15857), .ZN(n11382) );
  NAND2_X1 U11292 ( .A1(n11956), .A2(n9406), .ZN(n12470) );
  NOR2_X2 U11293 ( .A1(n14306), .A2(n14418), .ZN(n14286) );
  AOI21_X1 U11294 ( .B1(n12860), .B2(n14170), .A(n14158), .ZN(n12861) );
  NAND2_X1 U11295 ( .A1(n11868), .A2(n9722), .ZN(n10013) );
  AND2_X2 U11296 ( .A1(n10163), .A2(n10013), .ZN(n15841) );
  AOI22_X1 U11297 ( .A1(n12861), .A2(n14445), .B1(n15841), .B2(n12860), .ZN(
        n9409) );
  NOR4_X1 U11298 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9414) );
  NOR4_X1 U11299 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9413) );
  NOR4_X1 U11300 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9412) );
  NOR4_X1 U11301 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9411) );
  NAND4_X1 U11302 ( .A1(n9414), .A2(n9413), .A3(n9412), .A4(n9411), .ZN(n9432)
         );
  NOR2_X1 U11303 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n9418) );
  NOR4_X1 U11304 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9417) );
  NOR4_X1 U11305 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9416) );
  NOR4_X1 U11306 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n9415) );
  NAND4_X1 U11307 ( .A1(n9418), .A2(n9417), .A3(n9416), .A4(n9415), .ZN(n9431)
         );
  NAND2_X1 U11308 ( .A1(n9425), .A2(n9424), .ZN(n9420) );
  XNOR2_X1 U11309 ( .A(P2_B_REG_SCAN_IN), .B(n12158), .ZN(n9426) );
  INV_X1 U11310 ( .A(n9441), .ZN(n15520) );
  OAI21_X1 U11311 ( .B1(n9432), .B2(n9431), .A(n15520), .ZN(n10006) );
  OR2_X1 U11312 ( .A1(n15821), .A2(n9722), .ZN(n10014) );
  NAND2_X1 U11313 ( .A1(n9433), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9435) );
  INV_X1 U11314 ( .A(n9976), .ZN(n10016) );
  INV_X1 U11315 ( .A(n9437), .ZN(n10225) );
  NAND2_X1 U11316 ( .A1(n10225), .A2(n10013), .ZN(n11170) );
  AND3_X1 U11317 ( .A1(n10014), .A2(n15526), .A3(n11170), .ZN(n9439) );
  NAND2_X1 U11318 ( .A1(n12391), .A2(n12161), .ZN(n9438) );
  NAND2_X1 U11319 ( .A1(n12391), .A2(n12158), .ZN(n9440) );
  NAND2_X1 U11320 ( .A1(n9855), .A2(n14469), .ZN(n9443) );
  NAND2_X1 U11321 ( .A1(n9443), .A2(n9442), .ZN(P2_U3496) );
  NAND2_X1 U11322 ( .A1(n14080), .A2(n9529), .ZN(n9445) );
  OAI21_X1 U11323 ( .B1(n11189), .B2(n9529), .A(n9445), .ZN(n9467) );
  NAND2_X1 U11324 ( .A1(n14081), .A2(n9529), .ZN(n9447) );
  NAND2_X1 U11325 ( .A1(n9475), .A2(n11081), .ZN(n9446) );
  NAND2_X1 U11326 ( .A1(n9447), .A2(n9446), .ZN(n9455) );
  AOI22_X1 U11327 ( .A1(n14081), .A2(n9475), .B1(n11081), .B2(n9529), .ZN(
        n9456) );
  AND2_X1 U11328 ( .A1(n9467), .A2(n9473), .ZN(n9470) );
  NAND2_X1 U11329 ( .A1(n9450), .A2(n10885), .ZN(n9449) );
  NAND2_X1 U11330 ( .A1(n9451), .A2(n9454), .ZN(n9459) );
  NOR2_X1 U11331 ( .A1(n9452), .A2(n11173), .ZN(n9453) );
  AOI22_X1 U11332 ( .A1(n9475), .A2(n9000), .B1(n11213), .B2(n9529), .ZN(n9458) );
  AOI21_X1 U11333 ( .B1(n9459), .B2(n9457), .A(n9458), .ZN(n9463) );
  AOI22_X1 U11334 ( .A1(n9000), .A2(n9529), .B1(n9475), .B2(n11213), .ZN(n9462) );
  NAND2_X1 U11335 ( .A1(n9456), .A2(n9455), .ZN(n9461) );
  NAND3_X1 U11336 ( .A1(n9459), .A2(n9458), .A3(n9457), .ZN(n9460) );
  NAND2_X1 U11337 ( .A1(n14080), .A2(n9475), .ZN(n9466) );
  NAND2_X1 U11338 ( .A1(n9464), .A2(n7188), .ZN(n9465) );
  NAND2_X1 U11339 ( .A1(n9466), .A2(n9465), .ZN(n9471) );
  INV_X1 U11340 ( .A(n9467), .ZN(n9468) );
  INV_X1 U11341 ( .A(n9471), .ZN(n9472) );
  NAND2_X1 U11342 ( .A1(n9474), .A2(n8137), .ZN(n9481) );
  NAND2_X1 U11343 ( .A1(n11474), .A2(n9549), .ZN(n9477) );
  NAND2_X1 U11344 ( .A1(n14079), .A2(n7188), .ZN(n9476) );
  NAND2_X1 U11345 ( .A1(n9477), .A2(n9476), .ZN(n9482) );
  NAND2_X1 U11346 ( .A1(n11474), .A2(n7188), .ZN(n9478) );
  NAND2_X1 U11347 ( .A1(n10947), .A2(n7188), .ZN(n9484) );
  NAND2_X1 U11348 ( .A1(n14078), .A2(n9549), .ZN(n9483) );
  NAND2_X1 U11349 ( .A1(n9484), .A2(n9483), .ZN(n9487) );
  AOI22_X1 U11350 ( .A1(n10947), .A2(n9549), .B1(n14078), .B2(n7188), .ZN(
        n9485) );
  AOI21_X1 U11351 ( .B1(n9488), .B2(n9487), .A(n9485), .ZN(n9486) );
  NOR2_X1 U11352 ( .A1(n9488), .A2(n9487), .ZN(n9489) );
  NAND2_X1 U11353 ( .A1(n11455), .A2(n9549), .ZN(n9491) );
  NAND2_X1 U11354 ( .A1(n14077), .A2(n7188), .ZN(n9490) );
  NAND2_X1 U11355 ( .A1(n9491), .A2(n9490), .ZN(n9493) );
  AOI22_X1 U11356 ( .A1(n11455), .A2(n9662), .B1(n9604), .B2(n14077), .ZN(
        n9492) );
  NAND2_X1 U11357 ( .A1(n15840), .A2(n9662), .ZN(n9495) );
  NAND2_X1 U11358 ( .A1(n14076), .A2(n9549), .ZN(n9494) );
  NAND2_X1 U11359 ( .A1(n9495), .A2(n9494), .ZN(n9498) );
  AOI22_X1 U11360 ( .A1(n15840), .A2(n9549), .B1(n14076), .B2(n9662), .ZN(
        n9496) );
  AOI21_X1 U11361 ( .B1(n9499), .B2(n9498), .A(n9496), .ZN(n9497) );
  NOR2_X1 U11362 ( .A1(n9499), .A2(n9498), .ZN(n9500) );
  NAND2_X1 U11364 ( .A1(n11389), .A2(n9604), .ZN(n9502) );
  NAND2_X1 U11365 ( .A1(n14075), .A2(n9662), .ZN(n9501) );
  NAND2_X1 U11366 ( .A1(n11389), .A2(n9662), .ZN(n9503) );
  NAND2_X1 U11367 ( .A1(n12854), .A2(n9662), .ZN(n9506) );
  NAND2_X1 U11368 ( .A1(n14074), .A2(n9549), .ZN(n9505) );
  NAND2_X1 U11369 ( .A1(n9506), .A2(n9505), .ZN(n9509) );
  AOI22_X1 U11370 ( .A1(n12854), .A2(n9549), .B1(n14074), .B2(n9662), .ZN(
        n9507) );
  AOI21_X1 U11371 ( .B1(n9510), .B2(n9509), .A(n9507), .ZN(n9508) );
  INV_X1 U11372 ( .A(n9508), .ZN(n9511) );
  NAND2_X1 U11373 ( .A1(n9511), .A2(n7272), .ZN(n9517) );
  NAND2_X1 U11374 ( .A1(n12797), .A2(n9549), .ZN(n9513) );
  NAND2_X1 U11375 ( .A1(n14073), .A2(n7188), .ZN(n9512) );
  NAND2_X1 U11376 ( .A1(n9513), .A2(n9512), .ZN(n9518) );
  NAND2_X1 U11377 ( .A1(n9517), .A2(n9518), .ZN(n9516) );
  NAND2_X1 U11378 ( .A1(n12797), .A2(n9662), .ZN(n9514) );
  NAND2_X1 U11379 ( .A1(n9516), .A2(n9515), .ZN(n9522) );
  INV_X1 U11380 ( .A(n9517), .ZN(n9520) );
  INV_X1 U11381 ( .A(n9518), .ZN(n9519) );
  NAND2_X1 U11382 ( .A1(n11879), .A2(n7188), .ZN(n9524) );
  NAND2_X1 U11383 ( .A1(n14072), .A2(n9604), .ZN(n9523) );
  AOI22_X1 U11384 ( .A1(n11879), .A2(n9549), .B1(n14072), .B2(n7188), .ZN(
        n9525) );
  NAND2_X1 U11385 ( .A1(n11881), .A2(n9549), .ZN(n9527) );
  NAND2_X1 U11386 ( .A1(n14071), .A2(n7188), .ZN(n9526) );
  NAND2_X1 U11387 ( .A1(n9527), .A2(n9526), .ZN(n9534) );
  NAND2_X1 U11388 ( .A1(n9533), .A2(n9534), .ZN(n9532) );
  NAND2_X1 U11389 ( .A1(n11881), .A2(n9662), .ZN(n9528) );
  OAI21_X1 U11390 ( .B1(n9530), .B2(n9529), .A(n9528), .ZN(n9531) );
  NAND2_X1 U11391 ( .A1(n9532), .A2(n9531), .ZN(n9538) );
  INV_X1 U11392 ( .A(n9533), .ZN(n9536) );
  NAND2_X1 U11393 ( .A1(n9536), .A2(n9535), .ZN(n9537) );
  NAND2_X1 U11394 ( .A1(n12134), .A2(n9662), .ZN(n9540) );
  NAND2_X1 U11395 ( .A1(n13141), .A2(n9604), .ZN(n9539) );
  AOI22_X1 U11396 ( .A1(n12134), .A2(n9549), .B1(n13141), .B2(n7188), .ZN(
        n9541) );
  NAND2_X1 U11397 ( .A1(n12126), .A2(n9604), .ZN(n9543) );
  NAND2_X1 U11398 ( .A1(n14070), .A2(n9662), .ZN(n9542) );
  NAND2_X1 U11399 ( .A1(n9543), .A2(n9542), .ZN(n9546) );
  AOI22_X1 U11400 ( .A1(n12126), .A2(n7188), .B1(n9549), .B2(n14070), .ZN(
        n9544) );
  INV_X1 U11401 ( .A(n9545), .ZN(n9548) );
  NAND2_X1 U11402 ( .A1(n14444), .A2(n9662), .ZN(n9551) );
  NAND2_X1 U11403 ( .A1(n14069), .A2(n9549), .ZN(n9550) );
  NAND2_X1 U11404 ( .A1(n14444), .A2(n9604), .ZN(n9552) );
  OAI21_X1 U11405 ( .B1(n9553), .B2(n9549), .A(n9552), .ZN(n9554) );
  NAND2_X1 U11406 ( .A1(n14438), .A2(n9604), .ZN(n9556) );
  NAND2_X1 U11407 ( .A1(n14354), .A2(n9662), .ZN(n9555) );
  NAND2_X1 U11408 ( .A1(n9556), .A2(n9555), .ZN(n9558) );
  AOI22_X1 U11409 ( .A1(n14438), .A2(n9662), .B1(n9549), .B2(n14354), .ZN(
        n9557) );
  NAND2_X1 U11410 ( .A1(n14433), .A2(n9662), .ZN(n9562) );
  NAND2_X1 U11411 ( .A1(n14068), .A2(n9604), .ZN(n9561) );
  NAND2_X1 U11412 ( .A1(n14433), .A2(n9604), .ZN(n9563) );
  OAI21_X1 U11413 ( .B1(n14321), .B2(n9549), .A(n9563), .ZN(n9564) );
  NAND2_X1 U11414 ( .A1(n14428), .A2(n9604), .ZN(n9566) );
  NAND2_X1 U11415 ( .A1(n14356), .A2(n9662), .ZN(n9565) );
  NAND2_X1 U11416 ( .A1(n9566), .A2(n9565), .ZN(n9568) );
  AOI22_X1 U11417 ( .A1(n14428), .A2(n7188), .B1(n9549), .B2(n14356), .ZN(
        n9567) );
  AOI21_X1 U11418 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9571) );
  NOR2_X1 U11419 ( .A1(n9569), .A2(n9568), .ZN(n9570) );
  NAND2_X1 U11420 ( .A1(n14424), .A2(n7188), .ZN(n9573) );
  NAND2_X1 U11421 ( .A1(n14067), .A2(n9549), .ZN(n9572) );
  NAND2_X1 U11422 ( .A1(n9573), .A2(n9572), .ZN(n9577) );
  NAND2_X1 U11423 ( .A1(n9578), .A2(n9577), .ZN(n9576) );
  NAND2_X1 U11424 ( .A1(n14424), .A2(n9604), .ZN(n9574) );
  OAI21_X1 U11425 ( .B1(n9224), .B2(n9549), .A(n9574), .ZN(n9575) );
  NAND2_X1 U11426 ( .A1(n9576), .A2(n9575), .ZN(n9579) );
  NAND2_X1 U11427 ( .A1(n14418), .A2(n9604), .ZN(n9581) );
  NAND2_X1 U11428 ( .A1(n14066), .A2(n9662), .ZN(n9580) );
  AOI22_X1 U11429 ( .A1(n14418), .A2(n9662), .B1(n9549), .B2(n14066), .ZN(
        n9582) );
  NAND2_X1 U11430 ( .A1(n14413), .A2(n9662), .ZN(n9584) );
  NAND2_X1 U11431 ( .A1(n14251), .A2(n9549), .ZN(n9583) );
  NAND2_X1 U11432 ( .A1(n9584), .A2(n9583), .ZN(n9589) );
  NAND2_X1 U11433 ( .A1(n9588), .A2(n9589), .ZN(n9587) );
  NAND2_X1 U11434 ( .A1(n14413), .A2(n9549), .ZN(n9585) );
  OAI21_X1 U11435 ( .B1(n12505), .B2(n9549), .A(n9585), .ZN(n9586) );
  NAND2_X1 U11436 ( .A1(n9587), .A2(n9586), .ZN(n9593) );
  INV_X1 U11437 ( .A(n9588), .ZN(n9591) );
  INV_X1 U11438 ( .A(n9589), .ZN(n9590) );
  NAND2_X1 U11439 ( .A1(n9591), .A2(n9590), .ZN(n9592) );
  NAND2_X1 U11440 ( .A1(n14407), .A2(n9604), .ZN(n9595) );
  NAND2_X1 U11441 ( .A1(n14065), .A2(n7188), .ZN(n9594) );
  NAND2_X1 U11442 ( .A1(n9595), .A2(n9594), .ZN(n9597) );
  AOI22_X1 U11443 ( .A1(n14407), .A2(n9662), .B1(n9549), .B2(n14065), .ZN(
        n9596) );
  AOI21_X1 U11444 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n9600) );
  NOR2_X1 U11445 ( .A1(n9598), .A2(n9597), .ZN(n9599) );
  NAND2_X1 U11446 ( .A1(n14403), .A2(n7188), .ZN(n9602) );
  NAND2_X1 U11447 ( .A1(n14252), .A2(n9549), .ZN(n9601) );
  NAND2_X1 U11448 ( .A1(n9602), .A2(n9601), .ZN(n9608) );
  AND2_X1 U11449 ( .A1(n14064), .A2(n9662), .ZN(n9603) );
  AOI21_X1 U11450 ( .B1(n14396), .B2(n9549), .A(n9603), .ZN(n9614) );
  NAND2_X1 U11451 ( .A1(n14396), .A2(n9662), .ZN(n9606) );
  NAND2_X1 U11452 ( .A1(n14064), .A2(n9604), .ZN(n9605) );
  NAND2_X1 U11453 ( .A1(n9606), .A2(n9605), .ZN(n9613) );
  AOI22_X1 U11454 ( .A1(n14403), .A2(n9549), .B1(n14252), .B2(n7188), .ZN(
        n9607) );
  AOI21_X1 U11455 ( .B1(n9609), .B2(n9608), .A(n9607), .ZN(n9619) );
  AND2_X1 U11456 ( .A1(n14221), .A2(n7188), .ZN(n9610) );
  AOI21_X1 U11457 ( .B1(n14392), .B2(n9549), .A(n9610), .ZN(n9666) );
  NAND2_X1 U11458 ( .A1(n14392), .A2(n7188), .ZN(n9612) );
  NAND2_X1 U11459 ( .A1(n14221), .A2(n9549), .ZN(n9611) );
  NAND2_X1 U11460 ( .A1(n9612), .A2(n9611), .ZN(n9665) );
  AOI22_X1 U11461 ( .A1(n9666), .A2(n9665), .B1(n9614), .B2(n9613), .ZN(n9618)
         );
  AND2_X1 U11462 ( .A1(n14063), .A2(n9662), .ZN(n9615) );
  AOI21_X1 U11463 ( .B1(n14386), .B2(n9549), .A(n9615), .ZN(n9672) );
  NAND2_X1 U11464 ( .A1(n14386), .A2(n9662), .ZN(n9617) );
  NAND2_X1 U11465 ( .A1(n14063), .A2(n9549), .ZN(n9616) );
  NAND2_X1 U11466 ( .A1(n9617), .A2(n9616), .ZN(n9671) );
  NAND2_X1 U11467 ( .A1(n9672), .A2(n9671), .ZN(n9669) );
  OAI211_X1 U11468 ( .C1(n9620), .C2(n9619), .A(n9618), .B(n9669), .ZN(n9676)
         );
  INV_X1 U11469 ( .A(n9623), .ZN(n9624) );
  MUX2_X1 U11470 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10316), .Z(n9625) );
  NAND2_X1 U11471 ( .A1(n9625), .A2(SI_30_), .ZN(n9626) );
  OAI21_X1 U11472 ( .B1(n9625), .B2(SI_30_), .A(n9626), .ZN(n9639) );
  MUX2_X1 U11473 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10304), .Z(n9627) );
  XNOR2_X1 U11474 ( .A(n9627), .B(SI_31_), .ZN(n9628) );
  NAND2_X1 U11475 ( .A1(n15482), .A2(n9629), .ZN(n9632) );
  INV_X1 U11476 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9630) );
  OR2_X1 U11477 ( .A1(n9012), .A2(n9630), .ZN(n9631) );
  INV_X1 U11478 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U11479 ( .A1(n9633), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9635) );
  NAND2_X1 U11480 ( .A1(n9332), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9634) );
  OAI211_X1 U11481 ( .C1(n9637), .C2(n9636), .A(n9635), .B(n9634), .ZN(n14059)
         );
  INV_X1 U11482 ( .A(n14059), .ZN(n14153) );
  NAND2_X1 U11483 ( .A1(n14365), .A2(n14153), .ZN(n9694) );
  NAND2_X1 U11484 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  OR2_X1 U11485 ( .A1(n14930), .A2(n9643), .ZN(n9645) );
  INV_X1 U11486 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13151) );
  OR2_X1 U11487 ( .A1(n9012), .A2(n13151), .ZN(n9644) );
  AND2_X1 U11488 ( .A1(n14060), .A2(n9549), .ZN(n9646) );
  AOI21_X1 U11489 ( .B1(n14369), .B2(n9662), .A(n9646), .ZN(n9686) );
  NAND2_X1 U11490 ( .A1(n14369), .A2(n9549), .ZN(n9652) );
  OAI211_X1 U11491 ( .C1(n9647), .C2(n10009), .A(n9720), .B(n10013), .ZN(n9648) );
  AOI21_X1 U11492 ( .B1(n14059), .B2(n9662), .A(n9648), .ZN(n9649) );
  OR2_X1 U11493 ( .A1(n9650), .A2(n9649), .ZN(n9651) );
  NAND2_X1 U11494 ( .A1(n9652), .A2(n9651), .ZN(n9685) );
  AND2_X1 U11495 ( .A1(n14061), .A2(n9549), .ZN(n9653) );
  AOI21_X1 U11496 ( .B1(n12860), .B2(n7188), .A(n9653), .ZN(n9683) );
  NAND2_X1 U11497 ( .A1(n12860), .A2(n9549), .ZN(n9655) );
  NAND2_X1 U11498 ( .A1(n14061), .A2(n9662), .ZN(n9654) );
  NAND2_X1 U11499 ( .A1(n9655), .A2(n9654), .ZN(n9682) );
  AOI22_X1 U11500 ( .A1(n9686), .A2(n9685), .B1(n9683), .B2(n9682), .ZN(n9656)
         );
  OR2_X1 U11501 ( .A1(n9699), .A2(n9656), .ZN(n9690) );
  AND2_X1 U11502 ( .A1(n14062), .A2(n9549), .ZN(n9657) );
  AOI21_X1 U11503 ( .B1(n14373), .B2(n7188), .A(n9657), .ZN(n9681) );
  NAND2_X1 U11504 ( .A1(n14373), .A2(n9549), .ZN(n9659) );
  NAND2_X1 U11505 ( .A1(n14062), .A2(n7188), .ZN(n9658) );
  NAND2_X1 U11506 ( .A1(n9659), .A2(n9658), .ZN(n9680) );
  NAND2_X1 U11507 ( .A1(n9681), .A2(n9680), .ZN(n9660) );
  AND2_X1 U11508 ( .A1(n14190), .A2(n9604), .ZN(n9661) );
  AOI21_X1 U11509 ( .B1(n14377), .B2(n9662), .A(n9661), .ZN(n9678) );
  NAND2_X1 U11510 ( .A1(n14377), .A2(n9549), .ZN(n9664) );
  NAND2_X1 U11511 ( .A1(n14190), .A2(n7188), .ZN(n9663) );
  NAND2_X1 U11512 ( .A1(n9664), .A2(n9663), .ZN(n9677) );
  INV_X1 U11513 ( .A(n9665), .ZN(n9668) );
  INV_X1 U11514 ( .A(n9666), .ZN(n9667) );
  NAND3_X1 U11515 ( .A1(n9669), .A2(n9668), .A3(n9667), .ZN(n9670) );
  OAI21_X1 U11516 ( .B1(n9672), .B2(n9671), .A(n9670), .ZN(n9673) );
  AOI21_X1 U11517 ( .B1(n9678), .B2(n9677), .A(n9673), .ZN(n9674) );
  OAI22_X1 U11518 ( .A1(n9683), .A2(n9682), .B1(n9681), .B2(n9680), .ZN(n9684)
         );
  OR2_X1 U11519 ( .A1(n9699), .A2(n9684), .ZN(n9689) );
  INV_X1 U11520 ( .A(n9685), .ZN(n9688) );
  INV_X1 U11521 ( .A(n9686), .ZN(n9687) );
  AOI22_X1 U11522 ( .A1(n9690), .A2(n9689), .B1(n9688), .B2(n9687), .ZN(n9691)
         );
  NAND2_X1 U11523 ( .A1(n9692), .A2(n9691), .ZN(n9697) );
  NAND2_X1 U11524 ( .A1(n14059), .A2(n9475), .ZN(n9693) );
  OAI22_X1 U11525 ( .A1(n9694), .A2(n9604), .B1(n9693), .B2(n14365), .ZN(n9695) );
  INV_X1 U11526 ( .A(n9695), .ZN(n9696) );
  MUX2_X1 U11527 ( .A(n11862), .B(n12145), .S(n11868), .Z(n9717) );
  INV_X1 U11528 ( .A(n9699), .ZN(n9715) );
  XNOR2_X1 U11529 ( .A(n14413), .B(n14251), .ZN(n14266) );
  XNOR2_X1 U11530 ( .A(n12797), .B(n12851), .ZN(n11353) );
  OAI21_X1 U11531 ( .B1(n9450), .B2(n11403), .A(n13125), .ZN(n11406) );
  NAND4_X1 U11532 ( .A1(n10450), .A2(n9362), .A3(n10009), .A4(n11406), .ZN(
        n9700) );
  NOR4_X1 U11533 ( .A1(n10537), .A2(n10441), .A3(n9700), .A4(n11463), .ZN(
        n9702) );
  XNOR2_X1 U11534 ( .A(n10947), .B(n14078), .ZN(n10777) );
  NAND4_X1 U11535 ( .A1(n9702), .A2(n9701), .A3(n11202), .A4(n10777), .ZN(
        n9703) );
  NOR4_X1 U11536 ( .A1(n11507), .A2(n11353), .A3(n11342), .A4(n9703), .ZN(
        n9704) );
  NAND4_X1 U11537 ( .A1(n12396), .A2(n9704), .A3(n12052), .A4(n11841), .ZN(
        n9705) );
  NOR4_X1 U11538 ( .A1(n14338), .A2(n12475), .A3(n11951), .A4(n9705), .ZN(
        n9706) );
  XNOR2_X1 U11539 ( .A(n14418), .B(n14066), .ZN(n14282) );
  NAND4_X1 U11540 ( .A1(n14266), .A2(n14318), .A3(n9706), .A4(n14282), .ZN(
        n9707) );
  NOR3_X1 U11541 ( .A1(n14220), .A2(n14300), .A3(n9707), .ZN(n9710) );
  NAND4_X1 U11542 ( .A1(n14195), .A2(n9710), .A3(n9709), .A4(n9708), .ZN(n9711) );
  NOR4_X1 U11543 ( .A1(n14185), .A2(n12836), .A3(n14241), .A4(n9711), .ZN(
        n9714) );
  XNOR2_X1 U11544 ( .A(n14369), .B(n14060), .ZN(n9713) );
  NAND4_X1 U11545 ( .A1(n9715), .A2(n9714), .A3(n9713), .A4(n9712), .ZN(n9721)
         );
  NAND2_X1 U11546 ( .A1(n9720), .A2(n9722), .ZN(n9718) );
  OAI211_X1 U11547 ( .C1(n11173), .C2(n9726), .A(n10013), .B(n9718), .ZN(n9719) );
  NOR2_X1 U11548 ( .A1(n9721), .A2(n9720), .ZN(n9723) );
  NAND2_X1 U11549 ( .A1(n9723), .A2(n9722), .ZN(n9724) );
  INV_X1 U11550 ( .A(n10224), .ZN(n9725) );
  NAND2_X1 U11551 ( .A1(n9725), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12202) );
  INV_X1 U11552 ( .A(n15526), .ZN(n15523) );
  NOR4_X1 U11553 ( .A1(n15523), .A2(n14320), .A3(n12489), .A4(n10013), .ZN(
        n9728) );
  OAI21_X1 U11554 ( .B1(n12202), .B2(n9726), .A(P2_B_REG_SCAN_IN), .ZN(n9727)
         );
  OR2_X1 U11555 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  NAND3_X1 U11556 ( .A1(n9730), .A2(n9743), .A3(n9731), .ZN(n9843) );
  INV_X1 U11557 ( .A(n9831), .ZN(n9736) );
  NAND3_X1 U11558 ( .A1(n9744), .A2(n13965), .A3(n9731), .ZN(n9847) );
  AND2_X1 U11559 ( .A1(n13002), .A2(n9732), .ZN(n10678) );
  AND2_X1 U11560 ( .A1(n7204), .A2(n9734), .ZN(n9829) );
  NOR2_X1 U11561 ( .A1(n10678), .A2(n9829), .ZN(n9735) );
  OAI22_X1 U11562 ( .A1(n9843), .A2(n9736), .B1(n9847), .B2(n9735), .ZN(n9737)
         );
  OAI21_X1 U11563 ( .B1(n8747), .B2(n13610), .A(n11146), .ZN(n9745) );
  NAND2_X2 U11564 ( .A1(n9746), .A2(n9745), .ZN(n9749) );
  XNOR2_X1 U11565 ( .A(n12573), .B(n9749), .ZN(n9788) );
  XNOR2_X1 U11566 ( .A(n9806), .B(n15805), .ZN(n9758) );
  XNOR2_X1 U11567 ( .A(n9749), .B(n15782), .ZN(n9752) );
  XNOR2_X1 U11568 ( .A(n9752), .B(n13485), .ZN(n11084) );
  INV_X1 U11569 ( .A(n11208), .ZN(n12908) );
  XNOR2_X1 U11570 ( .A(n9749), .B(n12908), .ZN(n9750) );
  INV_X1 U11571 ( .A(n9750), .ZN(n9747) );
  NOR2_X1 U11572 ( .A1(n9747), .A2(n13486), .ZN(n11085) );
  OAI21_X1 U11573 ( .B1(n9812), .B2(n12895), .A(n11218), .ZN(n10686) );
  NOR2_X1 U11574 ( .A1(n10684), .A2(n7278), .ZN(n10971) );
  XNOR2_X1 U11575 ( .A(n9750), .B(n12909), .ZN(n10970) );
  XNOR2_X1 U11576 ( .A(n9806), .B(n11436), .ZN(n9753) );
  NOR2_X1 U11577 ( .A1(n9753), .A2(n13484), .ZN(n9754) );
  AOI21_X1 U11578 ( .B1(n13484), .B2(n9753), .A(n9754), .ZN(n11238) );
  INV_X1 U11579 ( .A(n9754), .ZN(n9755) );
  NAND2_X1 U11580 ( .A1(n11237), .A2(n9755), .ZN(n11427) );
  XNOR2_X1 U11581 ( .A(n9806), .B(n11811), .ZN(n9756) );
  XNOR2_X1 U11582 ( .A(n9756), .B(n13483), .ZN(n11428) );
  NAND2_X1 U11583 ( .A1(n9756), .A2(n11856), .ZN(n9757) );
  XNOR2_X1 U11584 ( .A(n9758), .B(n13482), .ZN(n11854) );
  XNOR2_X1 U11585 ( .A(n9806), .B(n11836), .ZN(n9759) );
  XNOR2_X1 U11586 ( .A(n9759), .B(n12085), .ZN(n11932) );
  XNOR2_X1 U11587 ( .A(n9806), .B(n12891), .ZN(n9760) );
  XNOR2_X1 U11588 ( .A(n9760), .B(n12892), .ZN(n12082) );
  XNOR2_X1 U11589 ( .A(n9806), .B(n15866), .ZN(n9761) );
  XNOR2_X1 U11590 ( .A(n9761), .B(n7681), .ZN(n12166) );
  NAND2_X1 U11591 ( .A1(n12165), .A2(n12166), .ZN(n12244) );
  XNOR2_X1 U11592 ( .A(n9806), .B(n12248), .ZN(n9763) );
  XNOR2_X1 U11593 ( .A(n9763), .B(n13479), .ZN(n12246) );
  NAND2_X1 U11594 ( .A1(n9761), .A2(n12256), .ZN(n12243) );
  AND2_X1 U11595 ( .A1(n9766), .A2(n9768), .ZN(n9767) );
  MUX2_X1 U11596 ( .A(n9767), .B(n13061), .S(n9806), .Z(n12317) );
  INV_X1 U11597 ( .A(n9768), .ZN(n9770) );
  INV_X1 U11598 ( .A(n12947), .ZN(n9769) );
  MUX2_X1 U11599 ( .A(n9770), .B(n9769), .S(n9806), .Z(n9771) );
  MUX2_X1 U11600 ( .A(n9772), .B(n12953), .S(n9806), .Z(n12409) );
  INV_X1 U11601 ( .A(n9773), .ZN(n9774) );
  MUX2_X1 U11602 ( .A(n9774), .B(n12952), .S(n9806), .Z(n12408) );
  XNOR2_X1 U11603 ( .A(n12958), .B(n9806), .ZN(n9775) );
  XNOR2_X1 U11604 ( .A(n9775), .B(n12957), .ZN(n12458) );
  NAND2_X1 U11605 ( .A1(n12459), .A2(n12458), .ZN(n12457) );
  NAND2_X1 U11606 ( .A1(n12457), .A2(n9777), .ZN(n12482) );
  XNOR2_X1 U11607 ( .A(n13913), .B(n9749), .ZN(n9778) );
  XNOR2_X1 U11608 ( .A(n9778), .B(n13248), .ZN(n12481) );
  NAND2_X1 U11609 ( .A1(n9778), .A2(n13263), .ZN(n9779) );
  XOR2_X1 U11610 ( .A(n9806), .B(n13836), .Z(n13194) );
  XNOR2_X1 U11611 ( .A(n13254), .B(n9806), .ZN(n13243) );
  AOI22_X1 U11612 ( .A1(n13194), .A2(n13261), .B1(n13262), .B2(n13243), .ZN(
        n9786) );
  INV_X1 U11613 ( .A(n13243), .ZN(n9780) );
  AND2_X1 U11614 ( .A1(n9780), .A2(n13832), .ZN(n9782) );
  INV_X1 U11615 ( .A(n9782), .ZN(n9784) );
  INV_X1 U11616 ( .A(n13194), .ZN(n9781) );
  OAI21_X1 U11617 ( .B1(n9782), .B2(n13809), .A(n9781), .ZN(n9783) );
  OAI21_X1 U11618 ( .B1(n9784), .B2(n13261), .A(n9783), .ZN(n9785) );
  XOR2_X1 U11619 ( .A(n9749), .B(n13900), .Z(n12539) );
  NAND2_X1 U11620 ( .A1(n12539), .A2(n13834), .ZN(n9787) );
  XNOR2_X1 U11621 ( .A(n9788), .B(n13808), .ZN(n12571) );
  XNOR2_X1 U11622 ( .A(n13784), .B(n9806), .ZN(n9789) );
  XNOR2_X1 U11623 ( .A(n9789), .B(n13760), .ZN(n13168) );
  INV_X1 U11624 ( .A(n9789), .ZN(n9790) );
  NAND2_X1 U11625 ( .A1(n9790), .A2(n13760), .ZN(n9791) );
  NAND2_X1 U11626 ( .A1(n9792), .A2(n9791), .ZN(n13213) );
  XNOR2_X1 U11627 ( .A(n13879), .B(n9749), .ZN(n9793) );
  XNOR2_X1 U11628 ( .A(n9793), .B(n13776), .ZN(n13214) );
  NAND2_X1 U11629 ( .A1(n13213), .A2(n13214), .ZN(n9795) );
  NAND2_X1 U11630 ( .A1(n9793), .A2(n13741), .ZN(n9794) );
  NAND2_X1 U11631 ( .A1(n9795), .A2(n9794), .ZN(n13175) );
  XNOR2_X1 U11632 ( .A(n13745), .B(n9806), .ZN(n13176) );
  MUX2_X1 U11633 ( .A(n13723), .B(n13717), .S(n9749), .Z(n9796) );
  XNOR2_X1 U11634 ( .A(n13870), .B(n9749), .ZN(n9797) );
  OR2_X1 U11635 ( .A1(n7331), .A2(n9799), .ZN(n9800) );
  XNOR2_X1 U11636 ( .A(n13927), .B(n9812), .ZN(n9802) );
  NAND2_X1 U11637 ( .A1(n9802), .A2(n13674), .ZN(n13183) );
  INV_X1 U11638 ( .A(n9802), .ZN(n9803) );
  NAND2_X1 U11639 ( .A1(n9803), .A2(n13708), .ZN(n9804) );
  NAND2_X1 U11640 ( .A1(n13183), .A2(n9804), .ZN(n13204) );
  INV_X1 U11641 ( .A(n13204), .ZN(n9805) );
  NAND2_X1 U11642 ( .A1(n13182), .A2(n13183), .ZN(n9810) );
  XNOR2_X1 U11643 ( .A(n13683), .B(n9806), .ZN(n9807) );
  NAND2_X1 U11644 ( .A1(n9807), .A2(n13662), .ZN(n9965) );
  INV_X1 U11645 ( .A(n9807), .ZN(n9808) );
  NAND2_X1 U11646 ( .A1(n9808), .A2(n13691), .ZN(n9809) );
  XNOR2_X1 U11647 ( .A(n8647), .B(n9812), .ZN(n9811) );
  NOR2_X1 U11648 ( .A1(n9811), .A2(n13257), .ZN(n9822) );
  AOI21_X1 U11649 ( .B1(n9811), .B2(n13257), .A(n9822), .ZN(n9968) );
  INV_X1 U11650 ( .A(n9968), .ZN(n9813) );
  XNOR2_X1 U11651 ( .A(n8699), .B(n9812), .ZN(n9817) );
  NOR2_X1 U11652 ( .A1(n9817), .A2(n13651), .ZN(n9816) );
  INV_X1 U11653 ( .A(n9816), .ZN(n9966) );
  AND2_X1 U11654 ( .A1(n9965), .A2(n9815), .ZN(n9814) );
  NAND2_X1 U11655 ( .A1(n13186), .A2(n9814), .ZN(n9821) );
  INV_X1 U11656 ( .A(n9815), .ZN(n9819) );
  AOI21_X1 U11657 ( .B1(n9817), .B2(n13651), .A(n9816), .ZN(n13234) );
  AND2_X1 U11658 ( .A1(n13234), .A2(n9968), .ZN(n9818) );
  NAND2_X1 U11659 ( .A1(n9821), .A2(n9820), .ZN(n9967) );
  INV_X1 U11660 ( .A(n9822), .ZN(n9823) );
  NAND2_X1 U11661 ( .A1(n9967), .A2(n9823), .ZN(n9825) );
  XNOR2_X1 U11662 ( .A(n13075), .B(n9749), .ZN(n9824) );
  XNOR2_X1 U11663 ( .A(n9825), .B(n9824), .ZN(n9852) );
  INV_X1 U11664 ( .A(n9829), .ZN(n9827) );
  NAND2_X1 U11665 ( .A1(n9831), .A2(n15912), .ZN(n9826) );
  OAI22_X1 U11666 ( .A1(n9843), .A2(n9827), .B1(n9847), .B2(n9826), .ZN(n9828)
         );
  NAND2_X1 U11667 ( .A1(n9843), .A2(n9829), .ZN(n9834) );
  AND2_X1 U11668 ( .A1(n10004), .A2(n9830), .ZN(n9833) );
  NAND2_X1 U11669 ( .A1(n9847), .A2(n9831), .ZN(n9832) );
  NAND4_X1 U11670 ( .A1(n9834), .A2(n9833), .A3(n10890), .A4(n9832), .ZN(n9835) );
  NAND2_X1 U11671 ( .A1(n9835), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9837) );
  AND2_X1 U11672 ( .A1(n10678), .A2(n10898), .ZN(n13089) );
  NAND2_X1 U11673 ( .A1(n9843), .A2(n13089), .ZN(n9836) );
  NAND2_X1 U11674 ( .A1(n13089), .A2(n9838), .ZN(n9839) );
  INV_X1 U11675 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n9840) );
  OAI22_X1 U11676 ( .A1(n13663), .A2(n13247), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9840), .ZN(n9845) );
  NAND2_X1 U11677 ( .A1(n13089), .A2(n9841), .ZN(n9842) );
  NOR2_X1 U11678 ( .A1(n13634), .A2(n13236), .ZN(n9844) );
  AOI211_X1 U11679 ( .C1(n13642), .C2(n13250), .A(n9845), .B(n9844), .ZN(n9846) );
  INV_X1 U11680 ( .A(n9846), .ZN(n9850) );
  NAND2_X1 U11681 ( .A1(n9847), .A2(n13084), .ZN(n9849) );
  AND2_X1 U11682 ( .A1(n10898), .A2(n15865), .ZN(n9848) );
  OAI21_X1 U11683 ( .B1(n9852), .B2(n13222), .A(n9851), .ZN(P3_U3160) );
  INV_X1 U11684 ( .A(n15525), .ZN(n9853) );
  NAND2_X1 U11685 ( .A1(n9855), .A2(n14451), .ZN(n9857) );
  NAND2_X1 U11686 ( .A1(n15908), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U11687 ( .A1(n9857), .A2(n9856), .ZN(P2_U3528) );
  INV_X1 U11688 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n13556) );
  INV_X1 U11689 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n9890) );
  NOR2_X1 U11690 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n9890), .ZN(n9858) );
  AOI21_X1 U11691 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(n9890), .A(n9858), .ZN(
        n9896) );
  INV_X1 U11692 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n9888) );
  INV_X1 U11693 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n9886) );
  INV_X1 U11694 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10702) );
  XNOR2_X1 U11695 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9942) );
  INV_X1 U11696 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9881) );
  INV_X1 U11697 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15110) );
  XNOR2_X1 U11698 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9903) );
  XNOR2_X1 U11699 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9906) );
  INV_X1 U11700 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n9875) );
  AND2_X1 U11701 ( .A1(n9872), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n9873) );
  INV_X1 U11702 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9859) );
  NAND2_X1 U11703 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n9915), .ZN(n9914) );
  NOR2_X1 U11704 ( .A1(n9860), .A2(n9861), .ZN(n9863) );
  XNOR2_X1 U11705 ( .A(n9861), .B(n9860), .ZN(n9917) );
  NOR2_X1 U11706 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n9917), .ZN(n9862) );
  NOR2_X1 U11707 ( .A1(n9864), .A2(n9865), .ZN(n9867) );
  NOR2_X1 U11708 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n9910), .ZN(n9866) );
  XNOR2_X1 U11709 ( .A(n9869), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U11710 ( .A1(n9908), .A2(n9907), .ZN(n9868) );
  INV_X1 U11711 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10178) );
  NAND2_X1 U11712 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n10178), .ZN(n9871) );
  INV_X1 U11713 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n9870) );
  NOR2_X1 U11714 ( .A1(n9875), .A2(n9874), .ZN(n9877) );
  XNOR2_X1 U11715 ( .A(n9875), .B(n9874), .ZN(n9932) );
  NAND2_X1 U11716 ( .A1(n9906), .A2(n9905), .ZN(n9878) );
  NAND2_X1 U11717 ( .A1(n9903), .A2(n9904), .ZN(n9879) );
  XOR2_X1 U11718 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n9901) );
  INV_X1 U11719 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10401) );
  NAND2_X1 U11720 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n10401), .ZN(n9883) );
  INV_X1 U11721 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n9882) );
  XNOR2_X1 U11722 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9899) );
  XOR2_X1 U11723 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n9897) );
  NOR2_X1 U11724 ( .A1(n9898), .A2(n9897), .ZN(n9887) );
  NAND2_X1 U11725 ( .A1(n9896), .A2(n9895), .ZN(n9889) );
  INV_X1 U11726 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9891) );
  NOR2_X1 U11727 ( .A1(n9892), .A2(n9891), .ZN(n9894) );
  XOR2_X1 U11728 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n9892), .Z(n9948) );
  NOR2_X1 U11729 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n9948), .ZN(n9893) );
  NOR2_X1 U11730 ( .A1(n9894), .A2(n9893), .ZN(n9953) );
  XOR2_X1 U11731 ( .A(n9953), .B(P1_ADDR_REG_17__SCAN_IN), .Z(n9954) );
  XNOR2_X1 U11732 ( .A(n13556), .B(n9954), .ZN(n9951) );
  XOR2_X1 U11733 ( .A(n9896), .B(n9895), .Z(n15652) );
  XOR2_X1 U11734 ( .A(n9898), .B(n9897), .Z(n9947) );
  XNOR2_X1 U11735 ( .A(n9900), .B(n9899), .ZN(n15643) );
  XOR2_X1 U11736 ( .A(n9902), .B(n9901), .Z(n15632) );
  XOR2_X1 U11737 ( .A(n9904), .B(n9903), .Z(n9937) );
  XOR2_X1 U11738 ( .A(n9906), .B(n9905), .Z(n9935) );
  AND2_X1 U11739 ( .A1(n9909), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n9923) );
  XNOR2_X1 U11740 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n9909), .ZN(n15613) );
  INV_X1 U11741 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9913) );
  NOR2_X1 U11742 ( .A1(n9912), .A2(n9913), .ZN(n9916) );
  OAI21_X1 U11743 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n9915), .A(n9914), .ZN(
        n15603) );
  NAND2_X1 U11744 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15603), .ZN(n15672) );
  NOR2_X1 U11745 ( .A1(n15673), .A2(n15672), .ZN(n15671) );
  XOR2_X1 U11746 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n9917), .Z(n15605) );
  NAND2_X1 U11747 ( .A1(n15606), .A2(n15605), .ZN(n15604) );
  NAND2_X1 U11748 ( .A1(n9921), .A2(n9919), .ZN(n9922) );
  INV_X1 U11749 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15609) );
  NOR2_X1 U11750 ( .A1(n15613), .A2(n15612), .ZN(n15611) );
  XNOR2_X1 U11751 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n9925) );
  XNOR2_X1 U11752 ( .A(n9925), .B(n9924), .ZN(n9927) );
  NOR2_X1 U11753 ( .A1(n9926), .A2(n9927), .ZN(n9928) );
  XNOR2_X1 U11754 ( .A(n9927), .B(n9926), .ZN(n15616) );
  INV_X1 U11755 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15615) );
  XNOR2_X1 U11756 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9930) );
  XOR2_X1 U11757 ( .A(n9930), .B(n9929), .Z(n15668) );
  INV_X1 U11758 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n15560) );
  NAND2_X1 U11759 ( .A1(n9931), .A2(n15560), .ZN(n9933) );
  XOR2_X1 U11760 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9932), .Z(n15618) );
  NAND2_X1 U11761 ( .A1(n15619), .A2(n15618), .ZN(n15617) );
  INV_X1 U11762 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15624) );
  INV_X1 U11763 ( .A(n15626), .ZN(n15627) );
  INV_X1 U11764 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15629) );
  NAND2_X1 U11765 ( .A1(n15632), .A2(n15631), .ZN(n9938) );
  XNOR2_X1 U11766 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9940) );
  XNOR2_X1 U11767 ( .A(n9940), .B(n9939), .ZN(n15635) );
  XOR2_X1 U11768 ( .A(n9942), .B(n9941), .Z(n9943) );
  NAND2_X1 U11769 ( .A1(n9944), .A2(n9943), .ZN(n9945) );
  INV_X1 U11770 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15639) );
  INV_X1 U11771 ( .A(n15646), .ZN(n15647) );
  INV_X1 U11772 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15649) );
  XOR2_X1 U11773 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n9948), .Z(n9950) );
  INV_X1 U11774 ( .A(n15655), .ZN(n15656) );
  INV_X1 U11775 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15658) );
  NAND2_X1 U11776 ( .A1(n15658), .A2(n15657), .ZN(n15654) );
  XNOR2_X1 U11777 ( .A(n9951), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(n15660) );
  INV_X1 U11778 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9952) );
  NOR2_X1 U11779 ( .A1(n9953), .A2(n9952), .ZN(n9956) );
  NOR2_X1 U11780 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n9954), .ZN(n9955) );
  NOR2_X1 U11781 ( .A1(n9956), .A2(n9955), .ZN(n9959) );
  INV_X1 U11782 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n13576) );
  NAND2_X1 U11783 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n13576), .ZN(n9957) );
  OAI21_X1 U11784 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n13576), .A(n9957), .ZN(
        n9958) );
  XNOR2_X1 U11785 ( .A(n9959), .B(n9958), .ZN(n15663) );
  NOR2_X1 U11786 ( .A1(n9959), .A2(n9958), .ZN(n9960) );
  AOI21_X1 U11787 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n13576), .A(n9960), .ZN(
        n9962) );
  XNOR2_X1 U11788 ( .A(n9962), .B(n9961), .ZN(n9963) );
  NAND2_X1 U11789 ( .A1(n13186), .A2(n9965), .ZN(n13233) );
  NAND2_X1 U11790 ( .A1(n13233), .A2(n13234), .ZN(n13232) );
  INV_X1 U11791 ( .A(n8647), .ZN(n13656) );
  INV_X1 U11792 ( .A(n13218), .ZN(n13255) );
  OAI22_X1 U11793 ( .A1(n13675), .A2(n13247), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9969), .ZN(n9972) );
  NOR2_X1 U11794 ( .A1(n9970), .A2(n13236), .ZN(n9971) );
  AOI211_X1 U11795 ( .C1(n13654), .C2(n13250), .A(n9972), .B(n9971), .ZN(n9973) );
  OAI21_X1 U11796 ( .B1(n13656), .B2(n13255), .A(n9973), .ZN(n9974) );
  INV_X1 U11797 ( .A(n9974), .ZN(n9975) );
  AND2_X1 U11798 ( .A1(n10224), .A2(n9976), .ZN(n10223) );
  NOR2_X1 U11799 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .ZN(n9980) );
  NAND3_X1 U11800 ( .A1(n11231), .A2(n11227), .A3(n9981), .ZN(n9982) );
  NAND4_X1 U11801 ( .A1(n9985), .A2(n9984), .A3(n10092), .A4(n10067), .ZN(
        n9986) );
  INV_X1 U11802 ( .A(n10106), .ZN(n9988) );
  NOR2_X1 U11803 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9991) );
  NAND2_X1 U11804 ( .A1(n9999), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10000) );
  NOR2_X1 U11805 ( .A1(n10468), .A2(P1_U3086), .ZN(n10003) );
  AND2_X2 U11806 ( .A1(n10293), .A2(n10003), .ZN(P1_U4016) );
  INV_X2 U11807 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U11808 ( .A(n15519), .ZN(n10007) );
  NAND2_X1 U11809 ( .A1(n10007), .A2(n10006), .ZN(n11172) );
  OR2_X1 U11810 ( .A1(n11172), .A2(n15525), .ZN(n10015) );
  INV_X1 U11811 ( .A(n10015), .ZN(n10008) );
  NAND2_X1 U11812 ( .A1(n10008), .A2(n15526), .ZN(n10034) );
  INV_X1 U11813 ( .A(n10034), .ZN(n10010) );
  AND2_X1 U11814 ( .A1(n10163), .A2(n10009), .ZN(n11176) );
  NAND2_X1 U11815 ( .A1(n10010), .A2(n11176), .ZN(n10012) );
  AND2_X1 U11816 ( .A1(n15526), .A2(n14140), .ZN(n10011) );
  OAI22_X1 U11817 ( .A1(n14044), .A2(n11189), .B1(n14050), .B2(n11064), .ZN(
        n10040) );
  OR2_X1 U11818 ( .A1(n14002), .A2(n14320), .ZN(n14031) );
  NOR2_X1 U11819 ( .A1(n14031), .A2(n13128), .ZN(n10039) );
  NAND2_X1 U11820 ( .A1(n10015), .A2(n10014), .ZN(n10018) );
  AND3_X1 U11821 ( .A1(n11170), .A2(n10224), .A3(n10016), .ZN(n10017) );
  NAND2_X1 U11822 ( .A1(n10018), .A2(n10017), .ZN(n10881) );
  INV_X1 U11823 ( .A(n14046), .ZN(n14030) );
  OAI22_X1 U11824 ( .A1(n14030), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n9021), .ZN(n10038) );
  NAND2_X1 U11825 ( .A1(n9000), .A2(n12832), .ZN(n10021) );
  NAND2_X1 U11826 ( .A1(n10019), .A2(n11173), .ZN(n12818) );
  XNOR2_X1 U11827 ( .A(n12818), .B(n11213), .ZN(n11075) );
  XNOR2_X1 U11828 ( .A(n10021), .B(n11075), .ZN(n13123) );
  INV_X1 U11829 ( .A(n13125), .ZN(n10489) );
  NAND2_X1 U11830 ( .A1(n10489), .A2(n12832), .ZN(n10880) );
  NAND2_X1 U11831 ( .A1(n11779), .A2(n10885), .ZN(n13124) );
  AND2_X1 U11832 ( .A1(n10880), .A2(n13124), .ZN(n10020) );
  NAND2_X1 U11833 ( .A1(n13123), .A2(n10020), .ZN(n13135) );
  INV_X1 U11834 ( .A(n11075), .ZN(n10022) );
  NAND2_X1 U11835 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  NAND2_X1 U11836 ( .A1(n13135), .A2(n10023), .ZN(n10024) );
  XNOR2_X1 U11837 ( .A(n12818), .B(n11081), .ZN(n10025) );
  NAND2_X1 U11838 ( .A1(n14081), .A2(n12832), .ZN(n10026) );
  XNOR2_X1 U11839 ( .A(n10025), .B(n10026), .ZN(n11076) );
  INV_X1 U11840 ( .A(n10025), .ZN(n10027) );
  NAND2_X1 U11841 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  XNOR2_X1 U11842 ( .A(n11189), .B(n12818), .ZN(n10846) );
  NAND2_X1 U11843 ( .A1(n14080), .A2(n12832), .ZN(n10029) );
  NAND2_X1 U11844 ( .A1(n10846), .A2(n10029), .ZN(n10032) );
  INV_X1 U11845 ( .A(n10846), .ZN(n10031) );
  INV_X1 U11846 ( .A(n10029), .ZN(n10030) );
  NAND2_X1 U11847 ( .A1(n10031), .A2(n10030), .ZN(n10849) );
  NAND2_X1 U11848 ( .A1(n10032), .A2(n10849), .ZN(n10035) );
  INV_X1 U11849 ( .A(n10851), .ZN(n10848) );
  OR3_X2 U11850 ( .A1(n10034), .A2(n10225), .A3(n15841), .ZN(n10844) );
  AOI211_X1 U11851 ( .C1(n10036), .C2(n10035), .A(n10848), .B(n10844), .ZN(
        n10037) );
  OR4_X1 U11852 ( .A1(n10040), .A2(n10039), .A3(n10038), .A4(n10037), .ZN(
        P2_U3190) );
  INV_X1 U11853 ( .A(n10524), .ZN(n10578) );
  NAND2_X1 U11854 ( .A1(n10578), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10041) );
  OAI21_X1 U11855 ( .B1(n10042), .B2(P3_STATE_REG_SCAN_IN), .A(n10041), .ZN(
        P3_U3294) );
  NAND2_X2 U11856 ( .A1(n10316), .A2(P1_U3086), .ZN(n15476) );
  INV_X1 U11857 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10325) );
  NOR2_X1 U11858 ( .A1(n10304), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15481) );
  INV_X2 U11859 ( .A(n15481), .ZN(n13160) );
  INV_X1 U11860 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n11229) );
  NOR2_X1 U11861 ( .A1(n10043), .A2(n11229), .ZN(n10044) );
  MUX2_X1 U11862 ( .A(n11229), .B(n10044), .S(P1_IR_REG_2__SCAN_IN), .Z(n10045) );
  INV_X1 U11863 ( .A(n10045), .ZN(n10047) );
  NAND2_X1 U11864 ( .A1(n10047), .A2(n10046), .ZN(n15079) );
  OAI222_X1 U11865 ( .A1(n15476), .A2(n10325), .B1(n13160), .B2(n10324), .C1(
        P1_U3086), .C2(n15079), .ZN(P1_U3353) );
  AND2_X1 U11866 ( .A1(n10304), .A2(P2_U3088), .ZN(n12201) );
  INV_X2 U11867 ( .A(n12201), .ZN(n14477) );
  NOR2_X1 U11868 ( .A1(n10316), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14475) );
  INV_X2 U11869 ( .A(n14475), .ZN(n13150) );
  OAI222_X1 U11870 ( .A1(n10272), .A2(P2_U3088), .B1(n14477), .B2(n10306), 
        .C1(n10048), .C2(n13150), .ZN(P2_U3326) );
  OAI222_X1 U11871 ( .A1(n13150), .A2(n10049), .B1(n14477), .B2(n10324), .C1(
        P2_U3088), .C2(n10260), .ZN(P2_U3325) );
  NOR2_X1 U11872 ( .A1(n10316), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13973) );
  INV_X1 U11873 ( .A(n10050), .ZN(n10052) );
  NAND2_X1 U11874 ( .A1(n10304), .A2(P3_U3151), .ZN(n13983) );
  OAI222_X1 U11875 ( .A1(n10673), .A2(P3_U3151), .B1(n13157), .B2(n10052), 
        .C1(n10051), .C2(n13983), .ZN(P3_U3293) );
  OAI222_X1 U11876 ( .A1(n10054), .A2(P3_U3151), .B1(n13157), .B2(n10053), 
        .C1(n10315), .C2(n13983), .ZN(P3_U3295) );
  OAI222_X1 U11877 ( .A1(n10716), .A2(P3_U3151), .B1(n13157), .B2(n10056), 
        .C1(n10055), .C2(n13983), .ZN(P3_U3289) );
  INV_X1 U11878 ( .A(n10057), .ZN(n10059) );
  INV_X1 U11879 ( .A(SI_5_), .ZN(n10058) );
  OAI222_X1 U11880 ( .A1(n10799), .A2(P3_U3151), .B1(n13157), .B2(n10059), 
        .C1(n10058), .C2(n13983), .ZN(P3_U3290) );
  INV_X1 U11881 ( .A(n10060), .ZN(n10062) );
  INV_X1 U11882 ( .A(SI_3_), .ZN(n10061) );
  OAI222_X1 U11883 ( .A1(n10599), .A2(P3_U3151), .B1(n13157), .B2(n10062), 
        .C1(n10061), .C2(n13983), .ZN(P3_U3292) );
  INV_X1 U11884 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U11885 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10063) );
  XNOR2_X1 U11886 ( .A(n10064), .B(n10063), .ZN(n15057) );
  OAI222_X1 U11887 ( .A1(n15057), .A2(P1_U3086), .B1(n13160), .B2(n10306), 
        .C1(n10305), .C2(n15476), .ZN(P1_U3354) );
  AOI22_X1 U11888 ( .A1(n10377), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n14475), .ZN(n10066) );
  OAI21_X1 U11889 ( .B1(n10335), .B2(n14477), .A(n10066), .ZN(P2_U3324) );
  INV_X1 U11890 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U11891 ( .A1(n10046), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10068) );
  XNOR2_X1 U11892 ( .A(n10068), .B(n10067), .ZN(n15096) );
  OAI222_X1 U11893 ( .A1(n15476), .A2(n10337), .B1(n13160), .B2(n10335), .C1(
        P1_U3086), .C2(n15096), .ZN(P1_U3352) );
  CLKBUF_X1 U11894 ( .A(n13983), .Z(n13969) );
  OAI222_X1 U11895 ( .A1(n13157), .A2(n10069), .B1(n13969), .B2(n13304), .C1(
        n11553), .C2(P3_U3151), .ZN(P3_U3285) );
  OAI222_X1 U11896 ( .A1(n13157), .A2(n10071), .B1(n13969), .B2(n10070), .C1(
        n10988), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U11897 ( .A(n10072), .ZN(n10074) );
  INV_X1 U11898 ( .A(SI_9_), .ZN(n10073) );
  INV_X1 U11899 ( .A(n11541), .ZN(n11554) );
  OAI222_X1 U11900 ( .A1(n13157), .A2(n10074), .B1(n13969), .B2(n10073), .C1(
        n11554), .C2(P3_U3151), .ZN(P3_U3286) );
  INV_X1 U11901 ( .A(n10075), .ZN(n10077) );
  INV_X1 U11902 ( .A(SI_7_), .ZN(n10076) );
  INV_X1 U11903 ( .A(n10727), .ZN(n10734) );
  OAI222_X1 U11904 ( .A1(n13157), .A2(n10077), .B1(n13969), .B2(n10076), .C1(
        n10734), .C2(P3_U3151), .ZN(P3_U3288) );
  OAI222_X1 U11905 ( .A1(n13157), .A2(n10078), .B1(n13969), .B2(n13419), .C1(
        n12303), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U11906 ( .A(n10640), .ZN(n10625) );
  INV_X1 U11907 ( .A(n10079), .ZN(n10080) );
  OAI222_X1 U11908 ( .A1(n10625), .A2(P3_U3151), .B1(n13157), .B2(n10080), 
        .C1(n7622), .C2(n13969), .ZN(P3_U3291) );
  INV_X1 U11909 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10807) );
  INV_X1 U11910 ( .A(n10806), .ZN(n10086) );
  OR2_X1 U11911 ( .A1(n10046), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U11912 ( .A1(n10082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10081) );
  MUX2_X1 U11913 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10081), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n10085) );
  INV_X1 U11914 ( .A(n10082), .ZN(n10084) );
  INV_X1 U11915 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U11916 ( .A1(n10084), .A2(n10083), .ZN(n10091) );
  NAND2_X1 U11917 ( .A1(n10085), .A2(n10091), .ZN(n15724) );
  OAI222_X1 U11918 ( .A1(n15476), .A2(n10807), .B1(n13160), .B2(n10086), .C1(
        P1_U3086), .C2(n15724), .ZN(P1_U3351) );
  INV_X1 U11919 ( .A(n10868), .ZN(n10246) );
  OAI222_X1 U11920 ( .A1(n13150), .A2(n10087), .B1(n14477), .B2(n10086), .C1(
        P2_U3088), .C2(n10246), .ZN(P2_U3323) );
  INV_X1 U11921 ( .A(n10817), .ZN(n10096) );
  AOI22_X1 U11922 ( .A1(n15535), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n14475), .ZN(n10088) );
  OAI21_X1 U11923 ( .B1(n10096), .B2(n14477), .A(n10088), .ZN(P2_U3322) );
  OAI222_X1 U11924 ( .A1(n13157), .A2(n10089), .B1(n13969), .B2(n13414), .C1(
        n12302), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U11925 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10097) );
  NAND2_X1 U11926 ( .A1(n10091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10090) );
  MUX2_X1 U11927 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10090), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n10094) );
  INV_X1 U11928 ( .A(n10091), .ZN(n10093) );
  NAND2_X1 U11929 ( .A1(n10093), .A2(n10092), .ZN(n10103) );
  INV_X1 U11930 ( .A(n10818), .ZN(n10095) );
  OAI222_X1 U11931 ( .A1(n15476), .A2(n10097), .B1(n13160), .B2(n10096), .C1(
        P1_U3086), .C2(n10095), .ZN(P1_U3350) );
  INV_X1 U11932 ( .A(n11028), .ZN(n10101) );
  INV_X1 U11933 ( .A(n15546), .ZN(n10098) );
  OAI222_X1 U11934 ( .A1(n13150), .A2(n10099), .B1(n14477), .B2(n10101), .C1(
        P2_U3088), .C2(n10098), .ZN(P2_U3321) );
  NAND2_X1 U11935 ( .A1(n10103), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10100) );
  XNOR2_X1 U11936 ( .A(n10100), .B(P1_IR_REG_6__SCAN_IN), .ZN(n11029) );
  INV_X1 U11937 ( .A(n11029), .ZN(n10437) );
  OAI222_X1 U11938 ( .A1(n15476), .A2(n10102), .B1(n13160), .B2(n10101), .C1(
        P1_U3086), .C2(n10437), .ZN(P1_U3349) );
  INV_X1 U11939 ( .A(n11292), .ZN(n10121) );
  OAI21_X1 U11940 ( .B1(n10103), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10104) );
  XNOR2_X1 U11941 ( .A(n10104), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11293) );
  INV_X1 U11942 ( .A(n15476), .ZN(n11702) );
  AOI22_X1 U11943 ( .A1(n11293), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n11702), .ZN(n10105) );
  OAI21_X1 U11944 ( .B1(n10121), .B2(n13160), .A(n10105), .ZN(P1_U3348) );
  XNOR2_X2 U11945 ( .A(n10108), .B(n10107), .ZN(n14755) );
  NAND2_X1 U11946 ( .A1(n10343), .A2(n14757), .ZN(n14937) );
  INV_X1 U11947 ( .A(n14937), .ZN(n10475) );
  NAND2_X1 U11948 ( .A1(n10475), .A2(n10293), .ZN(n10118) );
  INV_X1 U11949 ( .A(n10130), .ZN(n10115) );
  NOR2_X1 U11950 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(n10115), .ZN(n10116) );
  XNOR2_X2 U11951 ( .A(n10117), .B(n10131), .ZN(n10123) );
  NAND2_X1 U11952 ( .A1(n10118), .A2(n12641), .ZN(n10125) );
  NAND2_X1 U11953 ( .A1(n15013), .A2(n15471), .ZN(n10126) );
  AND2_X1 U11954 ( .A1(n10125), .A2(n10126), .ZN(n15732) );
  NOR2_X1 U11955 ( .A1(n15732), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11956 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10122) );
  INV_X1 U11957 ( .A(n15557), .ZN(n10120) );
  OAI222_X1 U11958 ( .A1(n13150), .A2(n10122), .B1(n14477), .B2(n10121), .C1(
        P2_U3088), .C2(n10120), .ZN(P2_U3320) );
  INV_X1 U11959 ( .A(n7200), .ZN(n15149) );
  INV_X1 U11960 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n15762) );
  AOI21_X1 U11961 ( .B1(n15149), .B2(n15762), .A(n7409), .ZN(n15076) );
  OAI21_X1 U11962 ( .B1(n15149), .B2(P1_REG1_REG_0__SCAN_IN), .A(n15076), .ZN(
        n10124) );
  XOR2_X1 U11963 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10124), .Z(n10129) );
  INV_X1 U11964 ( .A(n10125), .ZN(n10127) );
  NAND2_X1 U11965 ( .A1(n10127), .A2(n10126), .ZN(n10179) );
  AOI22_X1 U11966 ( .A1(n15732), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10128) );
  OAI21_X1 U11967 ( .B1(n10129), .B2(n10179), .A(n10128), .ZN(P1_U3243) );
  XNOR2_X2 U11968 ( .A(n10132), .B(n15475), .ZN(n13159) );
  NAND2_X1 U11969 ( .A1(n8101), .A2(n10133), .ZN(n10135) );
  XNOR2_X2 U11970 ( .A(n10137), .B(P1_IR_REG_29__SCAN_IN), .ZN(n10297) );
  INV_X2 U11971 ( .A(n10297), .ZN(n13153) );
  AND2_X4 U11972 ( .A1(n13159), .A2(n13153), .ZN(n14924) );
  NAND2_X1 U11973 ( .A1(n14924), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n10141) );
  INV_X1 U11974 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n10138) );
  OR2_X1 U11975 ( .A1(n14928), .A2(n10138), .ZN(n10140) );
  NAND2_X2 U11976 ( .A1(n10298), .A2(n13153), .ZN(n12692) );
  INV_X1 U11977 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n15148) );
  OR2_X1 U11978 ( .A1(n12705), .A2(n15148), .ZN(n10139) );
  AND3_X1 U11979 ( .A1(n10141), .A2(n10140), .A3(n10139), .ZN(n14943) );
  NAND2_X1 U11980 ( .A1(n15151), .A2(P1_U4016), .ZN(n10142) );
  OAI21_X1 U11981 ( .B1(P1_U4016), .B2(n9630), .A(n10142), .ZN(P1_U3591) );
  OAI222_X1 U11982 ( .A1(n13157), .A2(n10143), .B1(n13969), .B2(n13299), .C1(
        n13501), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U11983 ( .A(n11274), .ZN(n10149) );
  INV_X1 U11984 ( .A(n7497), .ZN(n11122) );
  NAND2_X1 U11985 ( .A1(n11122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10144) );
  MUX2_X1 U11986 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10144), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n10147) );
  INV_X1 U11987 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U11988 ( .A1(n7497), .A2(n10145), .ZN(n10157) );
  NAND2_X1 U11989 ( .A1(n10147), .A2(n10157), .ZN(n10402) );
  OAI222_X1 U11990 ( .A1(n15476), .A2(n10148), .B1(n13160), .B2(n10149), .C1(
        P1_U3086), .C2(n10402), .ZN(P1_U3347) );
  INV_X1 U11991 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10150) );
  INV_X1 U11992 ( .A(n11110), .ZN(n10876) );
  OAI222_X1 U11993 ( .A1(n13150), .A2(n10150), .B1(n14477), .B2(n10149), .C1(
        P2_U3088), .C2(n10876), .ZN(P2_U3319) );
  NAND2_X1 U11994 ( .A1(n13141), .A2(P2_U3947), .ZN(n10151) );
  OAI21_X1 U11995 ( .B1(n10152), .B2(P2_U3947), .A(n10151), .ZN(P2_U3544) );
  OAI222_X1 U11996 ( .A1(n13157), .A2(n10153), .B1(n13969), .B2(n13272), .C1(
        n13517), .C2(P3_U3151), .ZN(P3_U3281) );
  OAI222_X1 U11997 ( .A1(n13157), .A2(n10154), .B1(n13969), .B2(n13412), .C1(
        n13536), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U11998 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10155) );
  INV_X1 U11999 ( .A(n11582), .ZN(n10161) );
  INV_X1 U12000 ( .A(n11529), .ZN(n11117) );
  OAI222_X1 U12001 ( .A1(n13150), .A2(n10155), .B1(n14477), .B2(n10161), .C1(
        P2_U3088), .C2(n11117), .ZN(P2_U3318) );
  NAND2_X1 U12002 ( .A1(n10157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10156) );
  MUX2_X1 U12003 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10156), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n10160) );
  INV_X1 U12004 ( .A(n10157), .ZN(n10159) );
  INV_X1 U12005 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U12006 ( .A1(n10159), .A2(n10158), .ZN(n10397) );
  NAND2_X1 U12007 ( .A1(n10160), .A2(n10397), .ZN(n11583) );
  OAI222_X1 U12008 ( .A1(n15476), .A2(n10162), .B1(n13160), .B2(n10161), .C1(
        P1_U3086), .C2(n11583), .ZN(P1_U3346) );
  INV_X1 U12009 ( .A(n10163), .ZN(n10164) );
  OAI22_X1 U12010 ( .A1(n11406), .A2(n14449), .B1(n10164), .B2(n10885), .ZN(
        n10168) );
  AND2_X1 U12011 ( .A1(n10019), .A2(n14298), .ZN(n10165) );
  OR2_X1 U12012 ( .A1(n11406), .A2(n10165), .ZN(n10167) );
  NAND2_X1 U12013 ( .A1(n9000), .A2(n14355), .ZN(n10166) );
  NAND2_X1 U12014 ( .A1(n10167), .A2(n10166), .ZN(n11399) );
  NOR2_X1 U12015 ( .A1(n10168), .A2(n11399), .ZN(n15764) );
  NAND2_X1 U12016 ( .A1(n15908), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10169) );
  OAI21_X1 U12017 ( .B1(n15908), .B2(n15764), .A(n10169), .ZN(P2_U3499) );
  INV_X1 U12018 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10170) );
  MUX2_X1 U12019 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10170), .S(n10818), .Z(
        n10175) );
  INV_X1 U12020 ( .A(n15724), .ZN(n15740) );
  INV_X1 U12021 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10320) );
  MUX2_X1 U12022 ( .A(n10320), .B(P1_REG1_REG_2__SCAN_IN), .S(n15079), .Z(
        n15082) );
  INV_X1 U12023 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10299) );
  MUX2_X1 U12024 ( .A(n10299), .B(P1_REG1_REG_1__SCAN_IN), .S(n15057), .Z(
        n15062) );
  AND2_X1 U12025 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n15063) );
  NAND2_X1 U12026 ( .A1(n15062), .A2(n15063), .ZN(n15061) );
  INV_X1 U12027 ( .A(n15057), .ZN(n15064) );
  NAND2_X1 U12028 ( .A1(n15064), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U12029 ( .A1(n15061), .A2(n10171), .ZN(n15081) );
  NAND2_X1 U12030 ( .A1(n15082), .A2(n15081), .ZN(n15099) );
  OR2_X1 U12031 ( .A1(n15079), .A2(n10320), .ZN(n15098) );
  NAND2_X1 U12032 ( .A1(n15099), .A2(n15098), .ZN(n10173) );
  INV_X1 U12033 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10330) );
  MUX2_X1 U12034 ( .A(n10330), .B(P1_REG1_REG_3__SCAN_IN), .S(n15096), .Z(
        n10172) );
  NAND2_X1 U12035 ( .A1(n10173), .A2(n10172), .ZN(n15736) );
  OR2_X1 U12036 ( .A1(n15096), .A2(n10330), .ZN(n15735) );
  MUX2_X1 U12037 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10355), .S(n15724), .Z(
        n15734) );
  AOI21_X1 U12038 ( .B1(n15736), .B2(n15735), .A(n15734), .ZN(n15733) );
  AOI21_X1 U12039 ( .B1(n15740), .B2(P1_REG1_REG_4__SCAN_IN), .A(n15733), .ZN(
        n10174) );
  NAND2_X1 U12040 ( .A1(n10174), .A2(n10175), .ZN(n10202) );
  OAI21_X1 U12041 ( .B1(n10175), .B2(n10174), .A(n10202), .ZN(n10193) );
  INV_X1 U12042 ( .A(n15732), .ZN(n15145) );
  INV_X1 U12043 ( .A(n10179), .ZN(n10176) );
  NAND2_X1 U12044 ( .A1(n15741), .A2(n10818), .ZN(n10177) );
  NAND2_X1 U12045 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10934) );
  OAI211_X1 U12046 ( .C1(n10178), .C2(n15145), .A(n10177), .B(n10934), .ZN(
        n10192) );
  NOR2_X1 U12047 ( .A1(n10179), .A2(n7200), .ZN(n15139) );
  INV_X1 U12048 ( .A(n15139), .ZN(n10180) );
  XNOR2_X1 U12049 ( .A(n15079), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n15078) );
  INV_X1 U12050 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10181) );
  NAND2_X1 U12051 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n15056) );
  AOI21_X1 U12052 ( .B1(n15057), .B2(n10181), .A(n15056), .ZN(n10182) );
  OR2_X1 U12053 ( .A1(n15057), .A2(n10181), .ZN(n10183) );
  NAND2_X1 U12054 ( .A1(n10182), .A2(n10183), .ZN(n15058) );
  NAND2_X1 U12055 ( .A1(n15058), .A2(n10183), .ZN(n15077) );
  NAND2_X1 U12056 ( .A1(n15078), .A2(n15077), .ZN(n10185) );
  INV_X1 U12057 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n11330) );
  OR2_X1 U12058 ( .A1(n15079), .A2(n11330), .ZN(n10184) );
  NAND2_X1 U12059 ( .A1(n10185), .A2(n10184), .ZN(n15094) );
  INV_X1 U12060 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11734) );
  MUX2_X1 U12061 ( .A(n11734), .B(P1_REG2_REG_3__SCAN_IN), .S(n15096), .Z(
        n15095) );
  NAND2_X1 U12062 ( .A1(n15094), .A2(n15095), .ZN(n15726) );
  OR2_X1 U12063 ( .A1(n15096), .A2(n11734), .ZN(n15725) );
  NAND2_X1 U12064 ( .A1(n15726), .A2(n15725), .ZN(n10187) );
  INV_X1 U12065 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11692) );
  MUX2_X1 U12066 ( .A(n11692), .B(P1_REG2_REG_4__SCAN_IN), .S(n15724), .Z(
        n10186) );
  NAND2_X1 U12067 ( .A1(n10187), .A2(n10186), .ZN(n15729) );
  NAND2_X1 U12068 ( .A1(n15740), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10189) );
  INV_X1 U12069 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11706) );
  MUX2_X1 U12070 ( .A(n11706), .B(P1_REG2_REG_5__SCAN_IN), .S(n10818), .Z(
        n10188) );
  AOI21_X1 U12071 ( .B1(n15729), .B2(n10189), .A(n10188), .ZN(n10207) );
  AND3_X1 U12072 ( .A1(n15729), .A2(n10189), .A3(n10188), .ZN(n10190) );
  NOR3_X1 U12073 ( .A1(n15087), .A2(n10207), .A3(n10190), .ZN(n10191) );
  AOI211_X1 U12074 ( .C1(n15739), .C2(n10193), .A(n10192), .B(n10191), .ZN(
        n10194) );
  INV_X1 U12075 ( .A(n10194), .ZN(P1_U3248) );
  INV_X1 U12076 ( .A(n10195), .ZN(n10196) );
  OAI222_X1 U12077 ( .A1(n13157), .A2(n10196), .B1(n13969), .B2(n13409), .C1(
        n13564), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12078 ( .A(n11587), .ZN(n10200) );
  NAND2_X1 U12079 ( .A1(n10397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10197) );
  XNOR2_X1 U12080 ( .A(n10197), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11588) );
  INV_X1 U12081 ( .A(n11588), .ZN(n10561) );
  OAI222_X1 U12082 ( .A1(n15476), .A2(n10198), .B1(n13160), .B2(n10200), .C1(
        P1_U3086), .C2(n10561), .ZN(P1_U3345) );
  INV_X1 U12083 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10201) );
  INV_X1 U12084 ( .A(n15597), .ZN(n10199) );
  OAI222_X1 U12085 ( .A1(n13150), .A2(n10201), .B1(n14477), .B2(n10200), .C1(
        P2_U3088), .C2(n10199), .ZN(P2_U3317) );
  OAI21_X1 U12086 ( .B1(n10818), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10202), .ZN(
        n10426) );
  INV_X1 U12087 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11140) );
  MUX2_X1 U12088 ( .A(n11140), .B(P1_REG1_REG_6__SCAN_IN), .S(n11029), .Z(
        n10425) );
  OR2_X1 U12089 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  NAND2_X1 U12090 ( .A1(n11029), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10204) );
  INV_X1 U12091 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15835) );
  MUX2_X1 U12092 ( .A(n15835), .B(P1_REG1_REG_7__SCAN_IN), .S(n11293), .Z(
        n10203) );
  AOI21_X1 U12093 ( .B1(n10427), .B2(n10204), .A(n10203), .ZN(n10388) );
  NAND3_X1 U12094 ( .A1(n10427), .A2(n10204), .A3(n10203), .ZN(n10205) );
  NAND2_X1 U12095 ( .A1(n15739), .A2(n10205), .ZN(n10216) );
  INV_X1 U12096 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10206) );
  NAND2_X1 U12097 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11414) );
  OAI21_X1 U12098 ( .B1(n15145), .B2(n10206), .A(n11414), .ZN(n10214) );
  AOI21_X1 U12099 ( .B1(n10818), .B2(P1_REG2_REG_5__SCAN_IN), .A(n10207), .ZN(
        n10431) );
  INV_X1 U12100 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10208) );
  MUX2_X1 U12101 ( .A(n10208), .B(P1_REG2_REG_6__SCAN_IN), .S(n11029), .Z(
        n10430) );
  NOR2_X1 U12102 ( .A1(n10431), .A2(n10430), .ZN(n10429) );
  NOR2_X1 U12103 ( .A1(n10437), .A2(n10208), .ZN(n10210) );
  INV_X1 U12104 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11571) );
  MUX2_X1 U12105 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n11571), .S(n11293), .Z(
        n10209) );
  OAI21_X1 U12106 ( .B1(n10429), .B2(n10210), .A(n10209), .ZN(n10386) );
  INV_X1 U12107 ( .A(n10386), .ZN(n10212) );
  NOR3_X1 U12108 ( .A1(n10429), .A2(n10210), .A3(n10209), .ZN(n10211) );
  NOR3_X1 U12109 ( .A1(n10212), .A2(n10211), .A3(n15087), .ZN(n10213) );
  AOI211_X1 U12110 ( .C1(n15741), .C2(n11293), .A(n10214), .B(n10213), .ZN(
        n10215) );
  OAI21_X1 U12111 ( .B1(n10388), .B2(n10216), .A(n10215), .ZN(P1_U3250) );
  OAI222_X1 U12112 ( .A1(n13579), .A2(P3_U3151), .B1(n13157), .B2(n10217), 
        .C1(n13405), .C2(n13969), .ZN(P3_U3278) );
  INV_X1 U12113 ( .A(n10260), .ZN(n10234) );
  INV_X1 U12114 ( .A(n10272), .ZN(n10232) );
  INV_X1 U12115 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U12116 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10263) );
  NOR2_X1 U12117 ( .A1(n10262), .A2(n10263), .ZN(n10261) );
  INV_X1 U12118 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10219) );
  MUX2_X1 U12119 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10219), .S(n10260), .Z(
        n10251) );
  NOR2_X1 U12120 ( .A1(n10252), .A2(n10251), .ZN(n10250) );
  AOI21_X1 U12121 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10234), .A(n10250), .ZN(
        n10373) );
  INV_X1 U12122 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10220) );
  MUX2_X1 U12123 ( .A(n10220), .B(P2_REG2_REG_3__SCAN_IN), .S(n10377), .Z(
        n10372) );
  INV_X1 U12124 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10221) );
  MUX2_X1 U12125 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10221), .S(n10868), .Z(
        n10222) );
  INV_X1 U12126 ( .A(n10222), .ZN(n10230) );
  INV_X1 U12127 ( .A(n10223), .ZN(n10229) );
  NAND2_X1 U12128 ( .A1(n10225), .A2(n10224), .ZN(n10227) );
  NAND2_X1 U12129 ( .A1(n10227), .A2(n10226), .ZN(n10228) );
  AND2_X1 U12130 ( .A1(n10229), .A2(n10228), .ZN(n10243) );
  NOR2_X1 U12131 ( .A1(n9400), .A2(P2_U3088), .ZN(n12512) );
  INV_X1 U12132 ( .A(n15583), .ZN(n15592) );
  AOI211_X1 U12133 ( .C1(n10231), .C2(n10230), .A(n15592), .B(n10861), .ZN(
        n10249) );
  INV_X1 U12134 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10502) );
  AND3_X1 U12135 ( .A1(n10264), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG1_REG_0__SCAN_IN), .ZN(n10265) );
  AOI21_X1 U12136 ( .B1(n10232), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10265), .ZN(
        n10255) );
  INV_X1 U12137 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10233) );
  MUX2_X1 U12138 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10233), .S(n10260), .Z(
        n10254) );
  NOR2_X1 U12139 ( .A1(n10255), .A2(n10254), .ZN(n10253) );
  AOI21_X1 U12140 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n10234), .A(n10253), .ZN(
        n10376) );
  INV_X1 U12141 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10235) );
  MUX2_X1 U12142 ( .A(n10235), .B(P2_REG1_REG_3__SCAN_IN), .S(n10377), .Z(
        n10375) );
  NOR2_X1 U12143 ( .A1(n10376), .A2(n10375), .ZN(n10374) );
  AOI21_X1 U12144 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n10377), .A(n10374), .ZN(
        n10241) );
  INV_X1 U12145 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10236) );
  MUX2_X1 U12146 ( .A(n10236), .B(P2_REG1_REG_4__SCAN_IN), .S(n10868), .Z(
        n10240) );
  INV_X1 U12147 ( .A(n10237), .ZN(n10239) );
  NOR2_X1 U12148 ( .A1(n10241), .A2(n10240), .ZN(n10867) );
  AOI211_X1 U12149 ( .C1(n10241), .C2(n10240), .A(n15588), .B(n10867), .ZN(
        n10248) );
  NAND2_X1 U12150 ( .A1(n10242), .A2(n9400), .ZN(n15575) );
  AND2_X1 U12151 ( .A1(n10243), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15522) );
  NAND2_X1 U12152 ( .A1(n15522), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U12153 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10244) );
  OAI211_X1 U12154 ( .C1(n14148), .C2(n10246), .A(n10245), .B(n10244), .ZN(
        n10247) );
  OR3_X1 U12155 ( .A1(n10249), .A2(n10248), .A3(n10247), .ZN(P2_U3218) );
  AOI211_X1 U12156 ( .C1(n10252), .C2(n10251), .A(n10250), .B(n15592), .ZN(
        n10257) );
  AOI211_X1 U12157 ( .C1(n10255), .C2(n10254), .A(n10253), .B(n15588), .ZN(
        n10256) );
  NOR2_X1 U12158 ( .A1(n10257), .A2(n10256), .ZN(n10259) );
  INV_X1 U12159 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U12160 ( .A1(n15522), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(P2_U3088), 
        .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n10258) );
  OAI211_X1 U12161 ( .C1(n10260), .C2(n14148), .A(n10259), .B(n10258), .ZN(
        P2_U3216) );
  AOI211_X1 U12162 ( .C1(n10263), .C2(n10262), .A(n10261), .B(n15592), .ZN(
        n10269) );
  NAND2_X1 U12163 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10267) );
  INV_X1 U12164 ( .A(n10264), .ZN(n10266) );
  AOI211_X1 U12165 ( .C1(n10267), .C2(n10266), .A(n10265), .B(n15588), .ZN(
        n10268) );
  NOR2_X1 U12166 ( .A1(n10269), .A2(n10268), .ZN(n10271) );
  AOI22_X1 U12167 ( .A1(n15522), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(P2_U3088), 
        .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n10270) );
  OAI211_X1 U12168 ( .C1(n10272), .C2(n14148), .A(n10271), .B(n10270), .ZN(
        P2_U3215) );
  INV_X1 U12169 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U12170 ( .A1(n10274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10275) );
  XNOR2_X2 U12171 ( .A(n10278), .B(P1_IR_REG_19__SCAN_IN), .ZN(n15140) );
  NAND2_X1 U12172 ( .A1(n15932), .A2(n15140), .ZN(n10482) );
  NAND2_X1 U12173 ( .A1(n12163), .A2(P1_B_REG_SCAN_IN), .ZN(n10279) );
  MUX2_X1 U12174 ( .A(n10279), .B(P1_B_REG_SCAN_IN), .S(n10294), .Z(n10280) );
  INV_X1 U12175 ( .A(n15472), .ZN(n10295) );
  NAND2_X1 U12176 ( .A1(n10281), .A2(n12163), .ZN(n15473) );
  OAI21_X1 U12177 ( .B1(n10295), .B2(P1_D_REG_1__SCAN_IN), .A(n15473), .ZN(
        n10472) );
  NOR4_X1 U12178 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n10286) );
  NOR4_X1 U12179 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n10285) );
  NOR4_X1 U12180 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n10284) );
  NOR4_X1 U12181 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n10283) );
  NAND4_X1 U12182 ( .A1(n10286), .A2(n10285), .A3(n10284), .A4(n10283), .ZN(
        n10292) );
  NOR2_X1 U12183 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n10290) );
  NOR4_X1 U12184 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n10289) );
  NOR4_X1 U12185 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n10288) );
  NOR4_X1 U12186 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n10287) );
  NAND4_X1 U12187 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n10291) );
  OAI21_X1 U12188 ( .B1(n10292), .B2(n10291), .A(n15472), .ZN(n11259) );
  OAI211_X1 U12189 ( .C1(n14937), .C2(n10462), .A(n10293), .B(n10468), .ZN(
        n10479) );
  INV_X1 U12190 ( .A(n10294), .ZN(n12157) );
  NAND2_X1 U12191 ( .A1(n10281), .A2(n12157), .ZN(n15474) );
  NOR2_X1 U12192 ( .A1(n15012), .A2(n11258), .ZN(n10296) );
  INV_X1 U12193 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11265) );
  OR2_X1 U12194 ( .A1(n12692), .A2(n10181), .ZN(n10301) );
  NAND4_X4 U12195 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n15054) );
  OR2_X1 U12196 ( .A1(n10336), .A2(n10305), .ZN(n10309) );
  OR2_X1 U12197 ( .A1(n14929), .A2(n10306), .ZN(n10308) );
  OR2_X1 U12198 ( .A1(n7202), .A2(n15057), .ZN(n10307) );
  NAND2_X1 U12199 ( .A1(n15054), .A2(n10771), .ZN(n14762) );
  INV_X1 U12200 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n15754) );
  INV_X1 U12201 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10467) );
  OR2_X1 U12202 ( .A1(n12692), .A2(n15762), .ZN(n10311) );
  OAI21_X1 U12203 ( .B1(n10316), .B2(n10315), .A(n10314), .ZN(n10317) );
  NAND2_X1 U12205 ( .A1(n7381), .A2(n10484), .ZN(n10527) );
  INV_X1 U12206 ( .A(n10771), .ZN(n11271) );
  OR2_X1 U12207 ( .A1(n15054), .A2(n11271), .ZN(n10319) );
  NAND2_X1 U12208 ( .A1(n10526), .A2(n10319), .ZN(n11320) );
  NAND2_X1 U12209 ( .A1(n14924), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n10323) );
  OR2_X1 U12210 ( .A1(n12692), .A2(n11330), .ZN(n10322) );
  INV_X1 U12211 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11329) );
  OR2_X1 U12212 ( .A1(n12704), .A2(n11329), .ZN(n10321) );
  NAND2_X1 U12213 ( .A1(n7377), .A2(n14769), .ZN(n10328) );
  NAND2_X1 U12214 ( .A1(n11320), .A2(n14951), .ZN(n11319) );
  NAND2_X1 U12215 ( .A1(n11319), .A2(n10329), .ZN(n10341) );
  NAND2_X1 U12216 ( .A1(n14924), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n10334) );
  OR2_X1 U12217 ( .A1(n14928), .A2(n10330), .ZN(n10333) );
  OR2_X1 U12218 ( .A1(n10336), .A2(n10337), .ZN(n10339) );
  OR2_X1 U12219 ( .A1(n12641), .A2(n15096), .ZN(n10338) );
  XNOR2_X1 U12220 ( .A(n15052), .B(n10825), .ZN(n14950) );
  NAND2_X1 U12221 ( .A1(n10341), .A2(n14950), .ZN(n10805) );
  OAI21_X1 U12222 ( .B1(n10341), .B2(n14950), .A(n10805), .ZN(n11736) );
  INV_X1 U12223 ( .A(n11736), .ZN(n10364) );
  NAND2_X4 U12224 ( .A1(n14756), .A2(n14758), .ZN(n14628) );
  OR2_X1 U12225 ( .A1(n14756), .A2(n14758), .ZN(n10344) );
  NAND2_X1 U12226 ( .A1(n11566), .A2(n10342), .ZN(n11328) );
  AND2_X1 U12227 ( .A1(n7187), .A2(n15140), .ZN(n15750) );
  NAND2_X1 U12228 ( .A1(n14755), .A2(n15750), .ZN(n15875) );
  INV_X1 U12229 ( .A(n10525), .ZN(n10345) );
  NAND2_X1 U12230 ( .A1(n14763), .A2(n10345), .ZN(n10529) );
  NAND2_X1 U12231 ( .A1(n10529), .A2(n14765), .ZN(n10346) );
  NAND2_X1 U12232 ( .A1(n10346), .A2(n11321), .ZN(n11323) );
  NAND2_X1 U12233 ( .A1(n14607), .A2(n14769), .ZN(n14764) );
  NAND2_X1 U12234 ( .A1(n11323), .A2(n14764), .ZN(n10824) );
  INV_X1 U12235 ( .A(n14950), .ZN(n10347) );
  XNOR2_X1 U12236 ( .A(n10824), .B(n10347), .ZN(n10350) );
  NAND2_X1 U12237 ( .A1(n10343), .A2(n15140), .ZN(n10349) );
  NAND2_X1 U12238 ( .A1(n14757), .A2(n8111), .ZN(n10348) );
  NAND2_X1 U12239 ( .A1(n10350), .A2(n15988), .ZN(n10361) );
  NAND2_X1 U12240 ( .A1(n14924), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10359) );
  OR2_X1 U12241 ( .A1(n12692), .A2(n11692), .ZN(n10358) );
  INV_X1 U12242 ( .A(n10812), .ZN(n10354) );
  INV_X1 U12243 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10352) );
  INV_X1 U12244 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10351) );
  NAND2_X1 U12245 ( .A1(n10352), .A2(n10351), .ZN(n10353) );
  NAND2_X1 U12246 ( .A1(n10354), .A2(n10353), .ZN(n11689) );
  OR2_X1 U12247 ( .A1(n12704), .A2(n11689), .ZN(n10357) );
  INV_X1 U12248 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10355) );
  OR2_X1 U12249 ( .A1(n14928), .A2(n10355), .ZN(n10356) );
  NAND4_X1 U12250 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n15051) );
  INV_X1 U12251 ( .A(n7409), .ZN(n15072) );
  AOI22_X1 U12252 ( .A1(n15289), .A2(n7377), .B1(n15051), .B2(n15342), .ZN(
        n10360) );
  AND2_X1 U12253 ( .A1(n10361), .A2(n10360), .ZN(n11733) );
  NAND2_X1 U12254 ( .A1(n10771), .A2(n10528), .ZN(n11331) );
  AOI21_X1 U12255 ( .B1(n14776), .B2(n11332), .A(n11688), .ZN(n11731) );
  INV_X1 U12256 ( .A(n10462), .ZN(n10362) );
  AOI22_X1 U12257 ( .A1(n11731), .A2(n15932), .B1(n15981), .B2(n14776), .ZN(
        n10363) );
  OAI211_X1 U12258 ( .C1(n10364), .C2(n15985), .A(n11733), .B(n10363), .ZN(
        n10368) );
  NAND2_X1 U12259 ( .A1(n10368), .A2(n15991), .ZN(n10365) );
  OAI21_X1 U12260 ( .B1(n15991), .B2(n10330), .A(n10365), .ZN(P1_U3531) );
  INV_X1 U12261 ( .A(n11258), .ZN(n10473) );
  NOR2_X1 U12262 ( .A1(n15012), .A2(n10473), .ZN(n10366) );
  INV_X1 U12263 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10370) );
  NAND2_X1 U12264 ( .A1(n10368), .A2(n15994), .ZN(n10369) );
  OAI21_X1 U12265 ( .B1(n15994), .B2(n10370), .A(n10369), .ZN(P1_U3468) );
  AOI211_X1 U12266 ( .C1(n10373), .C2(n10372), .A(n10371), .B(n15592), .ZN(
        n10382) );
  AOI211_X1 U12267 ( .C1(n10376), .C2(n10375), .A(n15588), .B(n10374), .ZN(
        n10381) );
  NAND2_X1 U12268 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n10379) );
  NAND2_X1 U12269 ( .A1(n15598), .A2(n10377), .ZN(n10378) );
  OAI211_X1 U12270 ( .C1(n15601), .C2(n15609), .A(n10379), .B(n10378), .ZN(
        n10380) );
  OR3_X1 U12271 ( .A1(n10382), .A2(n10381), .A3(n10380), .ZN(P2_U3217) );
  NAND2_X1 U12272 ( .A1(n11293), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10385) );
  INV_X1 U12273 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10383) );
  MUX2_X1 U12274 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10383), .S(n10402), .Z(
        n10384) );
  AOI21_X1 U12275 ( .B1(n10386), .B2(n10385), .A(n10384), .ZN(n15115) );
  NAND3_X1 U12276 ( .A1(n10386), .A2(n10385), .A3(n10384), .ZN(n10387) );
  NAND2_X1 U12277 ( .A1(n10387), .A2(n15730), .ZN(n10396) );
  INV_X1 U12278 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n15853) );
  MUX2_X1 U12279 ( .A(n15853), .B(P1_REG1_REG_8__SCAN_IN), .S(n10402), .Z(
        n10390) );
  AOI21_X1 U12280 ( .B1(n11293), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10388), .ZN(
        n10389) );
  NAND2_X1 U12281 ( .A1(n10389), .A2(n10390), .ZN(n15106) );
  OAI21_X1 U12282 ( .B1(n10390), .B2(n10389), .A(n15106), .ZN(n10391) );
  NAND2_X1 U12283 ( .A1(n10391), .A2(n15739), .ZN(n10395) );
  INV_X1 U12284 ( .A(n10402), .ZN(n11275) );
  NAND2_X1 U12285 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11305) );
  OAI21_X1 U12286 ( .B1(n15145), .B2(n10392), .A(n11305), .ZN(n10393) );
  AOI21_X1 U12287 ( .B1(n11275), .B2(n15741), .A(n10393), .ZN(n10394) );
  OAI211_X1 U12288 ( .C1(n15115), .C2(n10396), .A(n10395), .B(n10394), .ZN(
        P1_U3251) );
  INV_X1 U12289 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11602) );
  NAND2_X1 U12290 ( .A1(n10565), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10398) );
  XNOR2_X1 U12291 ( .A(n10398), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11743) );
  MUX2_X1 U12292 ( .A(n11602), .B(P1_REG1_REG_11__SCAN_IN), .S(n11743), .Z(
        n10400) );
  INV_X1 U12293 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15899) );
  INV_X1 U12294 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15881) );
  NAND2_X1 U12295 ( .A1(n10402), .A2(n15853), .ZN(n15104) );
  MUX2_X1 U12296 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15881), .S(n11583), .Z(
        n15105) );
  AOI21_X1 U12297 ( .B1(n15106), .B2(n15104), .A(n15105), .ZN(n15108) );
  AOI21_X1 U12298 ( .B1(n15881), .B2(n11583), .A(n15108), .ZN(n10553) );
  MUX2_X1 U12299 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n15899), .S(n11588), .Z(
        n10552) );
  NAND2_X1 U12300 ( .A1(n10553), .A2(n10552), .ZN(n10551) );
  OAI21_X1 U12301 ( .B1(n15899), .B2(n10561), .A(n10551), .ZN(n10399) );
  NOR2_X1 U12302 ( .A1(n10399), .A2(n10400), .ZN(n10691) );
  AOI21_X1 U12303 ( .B1(n10400), .B2(n10399), .A(n10691), .ZN(n10413) );
  NAND2_X1 U12304 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11913)
         );
  OAI21_X1 U12305 ( .B1(n15145), .B2(n10401), .A(n11913), .ZN(n10411) );
  INV_X1 U12306 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10403) );
  NOR2_X1 U12307 ( .A1(n10402), .A2(n10383), .ZN(n15114) );
  MUX2_X1 U12308 ( .A(n10403), .B(P1_REG2_REG_9__SCAN_IN), .S(n11583), .Z(
        n15113) );
  OAI21_X1 U12309 ( .B1(n15115), .B2(n15114), .A(n15113), .ZN(n15117) );
  OAI21_X1 U12310 ( .B1(n10403), .B2(n11583), .A(n15117), .ZN(n10556) );
  INV_X1 U12311 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10404) );
  MUX2_X1 U12312 ( .A(n10404), .B(P1_REG2_REG_10__SCAN_IN), .S(n11588), .Z(
        n10405) );
  INV_X1 U12313 ( .A(n10405), .ZN(n10555) );
  NAND2_X1 U12314 ( .A1(n10556), .A2(n10555), .ZN(n10554) );
  NAND2_X1 U12315 ( .A1(n11588), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10408) );
  INV_X1 U12316 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10406) );
  MUX2_X1 U12317 ( .A(n10406), .B(P1_REG2_REG_11__SCAN_IN), .S(n11743), .Z(
        n10407) );
  AOI21_X1 U12318 ( .B1(n10554), .B2(n10408), .A(n10407), .ZN(n10698) );
  AND3_X1 U12319 ( .A1(n10554), .A2(n10408), .A3(n10407), .ZN(n10409) );
  NOR3_X1 U12320 ( .A1(n10698), .A2(n10409), .A3(n15087), .ZN(n10410) );
  AOI211_X1 U12321 ( .C1(n15741), .C2(n11743), .A(n10411), .B(n10410), .ZN(
        n10412) );
  OAI21_X1 U12322 ( .B1(n10413), .B2(n15135), .A(n10412), .ZN(P1_U3254) );
  INV_X1 U12323 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10414) );
  NAND2_X1 U12324 ( .A1(n15583), .A2(n10414), .ZN(n10415) );
  OAI211_X1 U12325 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15588), .A(n10415), .B(
        n14148), .ZN(n10416) );
  INV_X1 U12326 ( .A(n10416), .ZN(n10419) );
  INV_X1 U12327 ( .A(n15588), .ZN(n15581) );
  AOI22_X1 U12328 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n15581), .B1(n15583), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10418) );
  MUX2_X1 U12329 ( .A(n10419), .B(n10418), .S(n10417), .Z(n10421) );
  AOI22_X1 U12330 ( .A1(n15522), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10420) );
  NAND2_X1 U12331 ( .A1(n10421), .A2(n10420), .ZN(P2_U3214) );
  INV_X1 U12332 ( .A(n11742), .ZN(n10423) );
  INV_X1 U12333 ( .A(n11743), .ZN(n10692) );
  OAI222_X1 U12334 ( .A1(n15476), .A2(n10422), .B1(n13160), .B2(n10423), .C1(
        P1_U3086), .C2(n10692), .ZN(P1_U3344) );
  INV_X1 U12335 ( .A(n12100), .ZN(n11527) );
  OAI222_X1 U12336 ( .A1(n13150), .A2(n10424), .B1(n14477), .B2(n10423), .C1(
        P2_U3088), .C2(n11527), .ZN(P2_U3316) );
  INV_X1 U12337 ( .A(n15741), .ZN(n12771) );
  AOI21_X1 U12338 ( .B1(n10426), .B2(n10425), .A(n15135), .ZN(n10428) );
  NAND2_X1 U12339 ( .A1(n10428), .A2(n10427), .ZN(n10436) );
  NAND2_X1 U12340 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n11045) );
  AOI211_X1 U12341 ( .C1(n10431), .C2(n10430), .A(n10429), .B(n15087), .ZN(
        n10432) );
  INV_X1 U12342 ( .A(n10432), .ZN(n10433) );
  NAND2_X1 U12343 ( .A1(n11045), .A2(n10433), .ZN(n10434) );
  AOI21_X1 U12344 ( .B1(n15732), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10434), .ZN(
        n10435) );
  OAI211_X1 U12345 ( .C1(n12771), .C2(n10437), .A(n10436), .B(n10435), .ZN(
        P1_U3249) );
  OAI21_X1 U12346 ( .B1(n10439), .B2(n10441), .A(n10438), .ZN(n11481) );
  OR2_X1 U12347 ( .A1(n10542), .A2(n10855), .ZN(n10440) );
  NAND2_X1 U12348 ( .A1(n10783), .A2(n10440), .ZN(n11477) );
  OAI22_X1 U12349 ( .A1(n11477), .A2(n15821), .B1(n10855), .B2(n15903), .ZN(
        n10444) );
  XNOR2_X1 U12350 ( .A(n10442), .B(n10441), .ZN(n10443) );
  AOI22_X1 U12351 ( .A1(n14353), .A2(n14080), .B1(n14078), .B2(n14355), .ZN(
        n10853) );
  OAI21_X1 U12352 ( .B1(n10443), .B2(n14298), .A(n10853), .ZN(n11478) );
  AOI211_X1 U12353 ( .C1(n15860), .C2(n11481), .A(n10444), .B(n11478), .ZN(
        n10562) );
  NAND2_X1 U12354 ( .A1(n15908), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10445) );
  OAI21_X1 U12355 ( .B1(n10562), .B2(n15908), .A(n10445), .ZN(P2_U3503) );
  INV_X1 U12356 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10459) );
  OAI21_X1 U12357 ( .B1(n10448), .B2(n10447), .A(n10446), .ZN(n11182) );
  INV_X1 U12358 ( .A(n11182), .ZN(n10457) );
  INV_X1 U12359 ( .A(n10543), .ZN(n10449) );
  AOI211_X1 U12360 ( .C1(n11081), .C2(n10495), .A(n15821), .B(n10449), .ZN(
        n11179) );
  AOI21_X1 U12361 ( .B1(n15841), .B2(n11081), .A(n11179), .ZN(n10456) );
  XNOR2_X1 U12362 ( .A(n10451), .B(n10450), .ZN(n10455) );
  NAND2_X1 U12363 ( .A1(n9000), .A2(n14353), .ZN(n10453) );
  NAND2_X1 U12364 ( .A1(n14080), .A2(n14355), .ZN(n10452) );
  AND2_X1 U12365 ( .A1(n10453), .A2(n10452), .ZN(n11074) );
  INV_X1 U12366 ( .A(n11074), .ZN(n10454) );
  AOI21_X1 U12367 ( .B1(n10455), .B2(n14358), .A(n10454), .ZN(n11184) );
  OAI211_X1 U12368 ( .C1(n10457), .C2(n14442), .A(n10456), .B(n11184), .ZN(
        n14453) );
  NAND2_X1 U12369 ( .A1(n14453), .A2(n14469), .ZN(n10458) );
  OAI21_X1 U12370 ( .B1(n14469), .B2(n10459), .A(n10458), .ZN(P2_U3436) );
  INV_X1 U12371 ( .A(n15875), .ZN(n15779) );
  NAND2_X1 U12372 ( .A1(n7381), .A2(n10528), .ZN(n14760) );
  NAND2_X1 U12373 ( .A1(n14759), .A2(n14760), .ZN(n15758) );
  AND2_X1 U12374 ( .A1(n10484), .A2(n11263), .ZN(n15752) );
  INV_X1 U12375 ( .A(n15054), .ZN(n12780) );
  OAI21_X1 U12376 ( .B1(n15880), .B2(n15988), .A(n15758), .ZN(n10460) );
  OAI21_X1 U12377 ( .B1(n12780), .B2(n15195), .A(n10460), .ZN(n15756) );
  AOI211_X1 U12378 ( .C1(n15779), .C2(n15758), .A(n15752), .B(n15756), .ZN(
        n15749) );
  NAND2_X1 U12379 ( .A1(n15990), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10461) );
  OAI21_X1 U12380 ( .B1(n15749), .B2(n15990), .A(n10461), .ZN(P1_U3528) );
  NAND2_X1 U12381 ( .A1(n11263), .A2(n10462), .ZN(n11729) );
  AND2_X4 U12382 ( .A1(n14758), .A2(n10468), .ZN(n14581) );
  NAND2_X1 U12383 ( .A1(n7381), .A2(n14563), .ZN(n10466) );
  INV_X1 U12384 ( .A(n14758), .ZN(n10463) );
  AND2_X2 U12385 ( .A1(n10463), .A2(n10468), .ZN(n11286) );
  INV_X1 U12386 ( .A(n10468), .ZN(n10464) );
  AOI22_X1 U12387 ( .A1(n10484), .A2(n11286), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n10464), .ZN(n10465) );
  NAND2_X1 U12388 ( .A1(n10466), .A2(n10465), .ZN(n10756) );
  NAND2_X1 U12389 ( .A1(n7381), .A2(n11286), .ZN(n10471) );
  NOR2_X1 U12390 ( .A1(n10468), .A2(n10467), .ZN(n10469) );
  AOI21_X1 U12391 ( .B1(n10484), .B2(n14581), .A(n10469), .ZN(n10470) );
  NAND2_X1 U12392 ( .A1(n10471), .A2(n10470), .ZN(n10755) );
  XNOR2_X1 U12393 ( .A(n10756), .B(n10755), .ZN(n15070) );
  INV_X1 U12394 ( .A(n10472), .ZN(n11260) );
  AND3_X1 U12395 ( .A1(n10473), .A2(n11260), .A3(n11259), .ZN(n10477) );
  INV_X1 U12396 ( .A(n15471), .ZN(n10474) );
  NAND2_X1 U12397 ( .A1(n10477), .A2(n10474), .ZN(n10483) );
  OR2_X1 U12398 ( .A1(n15981), .A2(n10475), .ZN(n10476) );
  INV_X1 U12399 ( .A(n15012), .ZN(n11261) );
  NAND2_X1 U12400 ( .A1(n10477), .A2(n11261), .ZN(n14665) );
  INV_X1 U12401 ( .A(n14747), .ZN(n14644) );
  INV_X1 U12402 ( .A(n10477), .ZN(n10478) );
  NAND2_X1 U12403 ( .A1(n10478), .A2(n10482), .ZN(n10481) );
  INV_X1 U12404 ( .A(n10479), .ZN(n10480) );
  NAND2_X1 U12405 ( .A1(n10481), .A2(n10480), .ZN(n10935) );
  OR2_X1 U12406 ( .A1(n10935), .A2(P1_U3086), .ZN(n12783) );
  AOI22_X1 U12407 ( .A1(n14644), .A2(n15054), .B1(n12783), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10486) );
  OR2_X2 U12408 ( .A1(n10482), .A2(n15471), .ZN(n15755) );
  NAND2_X1 U12409 ( .A1(n10483), .A2(n15755), .ZN(n14645) );
  NAND2_X1 U12410 ( .A1(n14751), .A2(n10484), .ZN(n10485) );
  OAI211_X1 U12411 ( .C1(n15070), .C2(n14753), .A(n10486), .B(n10485), .ZN(
        P1_U3232) );
  INV_X1 U12412 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10499) );
  INV_X1 U12413 ( .A(n10487), .ZN(n10488) );
  AOI21_X1 U12414 ( .B1(n10489), .B2(n9362), .A(n10488), .ZN(n11216) );
  OAI21_X1 U12415 ( .B1(n10491), .B2(n9362), .A(n10490), .ZN(n10494) );
  INV_X1 U12416 ( .A(n9450), .ZN(n13129) );
  OAI22_X1 U12417 ( .A1(n13129), .A2(n14320), .B1(n13128), .B2(n14322), .ZN(
        n10493) );
  NOR2_X1 U12418 ( .A1(n11216), .A2(n10019), .ZN(n10492) );
  AOI211_X1 U12419 ( .C1(n14358), .C2(n10494), .A(n10493), .B(n10492), .ZN(
        n11209) );
  OAI21_X1 U12420 ( .B1(n13127), .B2(n10885), .A(n10495), .ZN(n11211) );
  INV_X1 U12421 ( .A(n11211), .ZN(n10496) );
  AOI22_X1 U12422 ( .A1(n10496), .A2(n14445), .B1(n15841), .B2(n11213), .ZN(
        n10497) );
  OAI211_X1 U12423 ( .C1(n11216), .C2(n14449), .A(n11209), .B(n10497), .ZN(
        n10500) );
  NAND2_X1 U12424 ( .A1(n10500), .A2(n14469), .ZN(n10498) );
  OAI21_X1 U12425 ( .B1(n14469), .B2(n10499), .A(n10498), .ZN(P2_U3433) );
  INV_X2 U12426 ( .A(n15908), .ZN(n14451) );
  NAND2_X1 U12427 ( .A1(n10500), .A2(n14451), .ZN(n10501) );
  OAI21_X1 U12428 ( .B1(n14451), .B2(n10502), .A(n10501), .ZN(P2_U3500) );
  INV_X1 U12429 ( .A(n10898), .ZN(n10503) );
  AND2_X1 U12430 ( .A1(n10504), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13086) );
  INV_X1 U12431 ( .A(n13086), .ZN(n13091) );
  NAND2_X1 U12432 ( .A1(n10503), .A2(n13091), .ZN(n10511) );
  OR2_X1 U12433 ( .A1(n13012), .A2(n10504), .ZN(n10506) );
  AND2_X1 U12434 ( .A1(n10506), .A2(n10505), .ZN(n10509) );
  NAND2_X1 U12435 ( .A1(n10511), .A2(n10509), .ZN(n10516) );
  MUX2_X1 U12436 ( .A(n13265), .B(n10516), .S(n7186), .Z(n13611) );
  NOR2_X1 U12437 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10888), .ZN(n15674) );
  NAND2_X1 U12438 ( .A1(n8297), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10596) );
  OAI21_X1 U12439 ( .B1(n10524), .B2(n15674), .A(n10596), .ZN(n10507) );
  OR2_X1 U12440 ( .A1(n10507), .A2(n8269), .ZN(n10597) );
  NAND2_X1 U12441 ( .A1(n10507), .A2(n8269), .ZN(n10508) );
  NAND2_X1 U12442 ( .A1(n10597), .A2(n10508), .ZN(n10520) );
  INV_X1 U12443 ( .A(n10509), .ZN(n10510) );
  NAND2_X1 U12444 ( .A1(n15702), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10512) );
  OAI21_X1 U12445 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n10513), .A(n10512), .ZN(
        n10519) );
  NOR2_X1 U12446 ( .A1(n10901), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15676) );
  NAND2_X1 U12447 ( .A1(n8297), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10585) );
  OAI21_X1 U12448 ( .B1(n10524), .B2(n15676), .A(n10585), .ZN(n10514) );
  OR2_X1 U12449 ( .A1(n10514), .A2(n11221), .ZN(n10586) );
  NAND2_X1 U12450 ( .A1(n10514), .A2(n11221), .ZN(n10517) );
  AOI21_X1 U12451 ( .B1(n10586), .B2(n10517), .A(n15677), .ZN(n10518) );
  AOI211_X1 U12452 ( .C1(n15675), .C2(n10520), .A(n10519), .B(n10518), .ZN(
        n10523) );
  MUX2_X1 U12453 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n8670), .Z(n10576) );
  XOR2_X1 U12454 ( .A(n10524), .B(n10576), .Z(n10579) );
  MUX2_X1 U12455 ( .A(n10901), .B(n10888), .S(n8670), .Z(n15680) );
  AND2_X1 U12456 ( .A1(n15680), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15679) );
  XNOR2_X1 U12457 ( .A(n10579), .B(n15679), .ZN(n10521) );
  AND2_X1 U12458 ( .A1(P3_U3897), .A2(n7186), .ZN(n15712) );
  NAND2_X1 U12459 ( .A1(n10521), .A2(n15712), .ZN(n10522) );
  OAI211_X1 U12460 ( .C1(n13611), .C2(n10524), .A(n10523), .B(n10522), .ZN(
        P3_U3183) );
  OAI21_X1 U12461 ( .B1(n10525), .B2(n10527), .A(n10526), .ZN(n11266) );
  OAI211_X1 U12462 ( .C1(n10528), .C2(n10771), .A(n15932), .B(n11331), .ZN(
        n11267) );
  OAI21_X1 U12463 ( .B1(n10771), .B2(n15970), .A(n11267), .ZN(n10533) );
  INV_X1 U12464 ( .A(n10529), .ZN(n11322) );
  AOI21_X1 U12465 ( .B1(n14759), .B2(n10525), .A(n11322), .ZN(n10532) );
  AOI22_X1 U12466 ( .A1(n15289), .A2(n7381), .B1(n7377), .B2(n15342), .ZN(
        n10531) );
  NAND2_X1 U12467 ( .A1(n11266), .A2(n15880), .ZN(n10530) );
  OAI211_X1 U12468 ( .C1(n10532), .C2(n15959), .A(n10531), .B(n10530), .ZN(
        n11262) );
  AOI211_X1 U12469 ( .C1(n15779), .C2(n11266), .A(n10533), .B(n11262), .ZN(
        n10548) );
  OR2_X1 U12470 ( .A1(n10548), .A2(n15990), .ZN(n10534) );
  OAI21_X1 U12471 ( .B1(n15991), .B2(n10299), .A(n10534), .ZN(P1_U3529) );
  INV_X1 U12472 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10547) );
  OAI21_X1 U12473 ( .B1(n10536), .B2(n10537), .A(n10535), .ZN(n11191) );
  INV_X1 U12474 ( .A(n11191), .ZN(n10545) );
  INV_X1 U12475 ( .A(n10019), .ZN(n14305) );
  OAI22_X1 U12476 ( .A1(n11064), .A2(n14322), .B1(n13128), .B2(n14320), .ZN(
        n10541) );
  XNOR2_X1 U12477 ( .A(n10538), .B(n10537), .ZN(n10539) );
  NOR2_X1 U12478 ( .A1(n10539), .A2(n14298), .ZN(n10540) );
  AOI211_X1 U12479 ( .C1(n14305), .C2(n11191), .A(n10541), .B(n10540), .ZN(
        n11193) );
  AOI21_X1 U12480 ( .B1(n9464), .B2(n10543), .A(n10542), .ZN(n11187) );
  AOI22_X1 U12481 ( .A1(n11187), .A2(n14445), .B1(n15841), .B2(n9464), .ZN(
        n10544) );
  OAI211_X1 U12482 ( .C1(n10545), .C2(n14449), .A(n11193), .B(n10544), .ZN(
        n14452) );
  NAND2_X1 U12483 ( .A1(n14452), .A2(n14469), .ZN(n10546) );
  OAI21_X1 U12484 ( .B1(n14469), .B2(n10547), .A(n10546), .ZN(P2_U3439) );
  INV_X1 U12485 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10550) );
  OR2_X1 U12486 ( .A1(n10548), .A2(n15992), .ZN(n10549) );
  OAI21_X1 U12487 ( .B1(n15994), .B2(n10550), .A(n10549), .ZN(P1_U3462) );
  OAI211_X1 U12488 ( .C1(n10553), .C2(n10552), .A(n10551), .B(n15739), .ZN(
        n10560) );
  NAND2_X1 U12489 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n11820)
         );
  OAI211_X1 U12490 ( .C1(n10556), .C2(n10555), .A(n15730), .B(n10554), .ZN(
        n10557) );
  NAND2_X1 U12491 ( .A1(n11820), .A2(n10557), .ZN(n10558) );
  AOI21_X1 U12492 ( .B1(n15732), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10558), 
        .ZN(n10559) );
  OAI211_X1 U12493 ( .C1(n12771), .C2(n10561), .A(n10560), .B(n10559), .ZN(
        P1_U3253) );
  INV_X1 U12494 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10564) );
  OR2_X1 U12495 ( .A1(n10562), .A2(n15909), .ZN(n10563) );
  OAI21_X1 U12496 ( .B1(n14469), .B2(n10564), .A(n10563), .ZN(P2_U3442) );
  INV_X1 U12497 ( .A(n11965), .ZN(n10609) );
  OAI21_X1 U12498 ( .B1(n10565), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10675) );
  XNOR2_X1 U12499 ( .A(n10675), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U12500 ( .A1(n11966), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n11702), .ZN(n10566) );
  OAI21_X1 U12501 ( .B1(n10609), .B2(n13160), .A(n10566), .ZN(P1_U3343) );
  NAND2_X1 U12502 ( .A1(n14252), .A2(P2_U3947), .ZN(n10567) );
  OAI21_X1 U12503 ( .B1(n10568), .B2(P2_U3947), .A(n10567), .ZN(P2_U3554) );
  INV_X1 U12504 ( .A(n13599), .ZN(n13588) );
  INV_X1 U12505 ( .A(n10569), .ZN(n10570) );
  OAI222_X1 U12506 ( .A1(n13588), .A2(P3_U3151), .B1(n13157), .B2(n10570), 
        .C1(n13291), .C2(n13969), .ZN(P3_U3277) );
  NAND2_X1 U12507 ( .A1(n13200), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10974) );
  INV_X1 U12508 ( .A(n10974), .ZN(n10575) );
  INV_X1 U12509 ( .A(n12896), .ZN(n13488) );
  XNOR2_X1 U12510 ( .A(n13488), .B(n10571), .ZN(n13058) );
  OAI22_X1 U12511 ( .A1(n13255), .A2(n10571), .B1(n10572), .B2(n13236), .ZN(
        n10573) );
  AOI21_X1 U12512 ( .B1(n13058), .B2(n13241), .A(n10573), .ZN(n10574) );
  OAI21_X1 U12513 ( .B1(n10575), .B2(n13457), .A(n10574), .ZN(P3_U3172) );
  MUX2_X1 U12514 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13087), .Z(n10626) );
  XOR2_X1 U12515 ( .A(n10640), .B(n10626), .Z(n10627) );
  INV_X1 U12516 ( .A(n10576), .ZN(n10577) );
  MUX2_X1 U12517 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n8670), .Z(n10580) );
  XOR2_X1 U12518 ( .A(n10595), .B(n10580), .Z(n10668) );
  OAI22_X1 U12519 ( .A1(n10669), .A2(n10668), .B1(n10580), .B2(n10673), .ZN(
        n10611) );
  MUX2_X1 U12520 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13087), .Z(n10581) );
  XNOR2_X1 U12521 ( .A(n10581), .B(n10622), .ZN(n10612) );
  INV_X1 U12522 ( .A(n10581), .ZN(n10582) );
  XOR2_X1 U12523 ( .A(n10628), .B(n10627), .Z(n10608) );
  MUX2_X1 U12524 ( .A(n10583), .B(P3_REG2_REG_4__SCAN_IN), .S(n10640), .Z(
        n10592) );
  MUX2_X1 U12525 ( .A(n10584), .B(P3_REG2_REG_2__SCAN_IN), .S(n10595), .Z(
        n10663) );
  NAND2_X1 U12526 ( .A1(n10586), .A2(n10585), .ZN(n10662) );
  NAND2_X1 U12527 ( .A1(n10663), .A2(n10662), .ZN(n10661) );
  NAND2_X1 U12528 ( .A1(n10673), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10587) );
  NAND2_X1 U12529 ( .A1(n10661), .A2(n10587), .ZN(n10588) );
  NAND2_X1 U12530 ( .A1(n10613), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10590) );
  NAND2_X1 U12531 ( .A1(n10588), .A2(n10599), .ZN(n10589) );
  NAND2_X1 U12532 ( .A1(n10590), .A2(n10589), .ZN(n10591) );
  NAND2_X1 U12533 ( .A1(n10591), .A2(n10592), .ZN(n10633) );
  OAI21_X1 U12534 ( .B1(n10592), .B2(n10591), .A(n10633), .ZN(n10593) );
  NAND2_X1 U12535 ( .A1(n15711), .A2(n10593), .ZN(n10605) );
  INV_X1 U12536 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10594) );
  MUX2_X1 U12537 ( .A(n10594), .B(P3_REG1_REG_4__SCAN_IN), .S(n10640), .Z(
        n10601) );
  MUX2_X1 U12538 ( .A(n8290), .B(P3_REG1_REG_2__SCAN_IN), .S(n10595), .Z(
        n10658) );
  NAND2_X1 U12539 ( .A1(n10597), .A2(n10596), .ZN(n10657) );
  NAND2_X1 U12540 ( .A1(n10658), .A2(n10657), .ZN(n10656) );
  NAND2_X1 U12541 ( .A1(n10673), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10598) );
  NAND2_X1 U12542 ( .A1(n10600), .A2(n10601), .ZN(n10642) );
  OAI21_X1 U12543 ( .B1(n10601), .B2(n10600), .A(n10642), .ZN(n10602) );
  NAND2_X1 U12544 ( .A1(n15675), .A2(n10602), .ZN(n10604) );
  INV_X1 U12545 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n13367) );
  NOR2_X1 U12546 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13367), .ZN(n11243) );
  AOI21_X1 U12547 ( .B1(n15702), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11243), .ZN(
        n10603) );
  NAND3_X1 U12548 ( .A1(n10605), .A2(n10604), .A3(n10603), .ZN(n10606) );
  AOI21_X1 U12549 ( .B1(n10640), .B2(n15704), .A(n10606), .ZN(n10607) );
  OAI21_X1 U12550 ( .B1(n10608), .B2(n15681), .A(n10607), .ZN(P3_U3186) );
  OAI222_X1 U12551 ( .A1(n13150), .A2(n10610), .B1(n14477), .B2(n10609), .C1(
        n15574), .C2(P2_U3088), .ZN(P2_U3315) );
  XOR2_X1 U12552 ( .A(n10612), .B(n10611), .Z(n10624) );
  XOR2_X1 U12553 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n10613), .Z(n10620) );
  NAND2_X1 U12554 ( .A1(n10614), .A2(n8306), .ZN(n10615) );
  NAND2_X1 U12555 ( .A1(n10616), .A2(n10615), .ZN(n10617) );
  NAND2_X1 U12556 ( .A1(n15675), .A2(n10617), .ZN(n10619) );
  INV_X1 U12557 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n13333) );
  NOR2_X1 U12558 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13333), .ZN(n11089) );
  AOI21_X1 U12559 ( .B1(n15702), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n11089), .ZN(
        n10618) );
  OAI211_X1 U12560 ( .C1(n10620), .C2(n15677), .A(n10619), .B(n10618), .ZN(
        n10621) );
  AOI21_X1 U12561 ( .B1(n10622), .B2(n15704), .A(n10621), .ZN(n10623) );
  OAI21_X1 U12562 ( .B1(n10624), .B2(n15681), .A(n10623), .ZN(P3_U3185) );
  MUX2_X1 U12563 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13087), .Z(n10725) );
  XNOR2_X1 U12564 ( .A(n10725), .B(n10727), .ZN(n10728) );
  OAI22_X1 U12565 ( .A1(n10628), .A2(n10627), .B1(n10626), .B2(n10625), .ZN(
        n10791) );
  MUX2_X1 U12566 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13087), .Z(n10629) );
  XNOR2_X1 U12567 ( .A(n10629), .B(n10634), .ZN(n10792) );
  INV_X1 U12568 ( .A(n10629), .ZN(n10630) );
  AOI22_X1 U12569 ( .A1(n10791), .A2(n10792), .B1(n10634), .B2(n10630), .ZN(
        n10717) );
  MUX2_X1 U12570 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13087), .Z(n10631) );
  XNOR2_X1 U12571 ( .A(n10631), .B(n10716), .ZN(n10718) );
  XOR2_X1 U12572 ( .A(n10729), .B(n10728), .Z(n10655) );
  INV_X1 U12573 ( .A(n10716), .ZN(n10638) );
  INV_X1 U12574 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15809) );
  OR2_X1 U12575 ( .A1(n10640), .A2(n10583), .ZN(n10632) );
  NAND2_X1 U12576 ( .A1(n10633), .A2(n10632), .ZN(n10635) );
  XNOR2_X1 U12577 ( .A(n10635), .B(n10634), .ZN(n10793) );
  NAND2_X1 U12578 ( .A1(n10793), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n10637) );
  NAND2_X1 U12579 ( .A1(n10635), .A2(n10799), .ZN(n10636) );
  NAND2_X1 U12580 ( .A1(n10637), .A2(n10636), .ZN(n10708) );
  MUX2_X1 U12581 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n15809), .S(n10716), .Z(
        n10709) );
  NAND2_X1 U12582 ( .A1(n10708), .A2(n10709), .ZN(n10707) );
  OAI21_X1 U12583 ( .B1(n10639), .B2(P3_REG2_REG_7__SCAN_IN), .A(n10736), .ZN(
        n10653) );
  OR2_X1 U12584 ( .A1(n10640), .A2(n10594), .ZN(n10641) );
  NAND2_X1 U12585 ( .A1(n10642), .A2(n10641), .ZN(n10643) );
  NAND2_X1 U12586 ( .A1(n10643), .A2(n10799), .ZN(n10644) );
  NAND2_X1 U12587 ( .A1(n10796), .A2(n10644), .ZN(n10711) );
  INV_X1 U12588 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10645) );
  MUX2_X1 U12589 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10645), .S(n10716), .Z(
        n10712) );
  NAND2_X1 U12590 ( .A1(n10711), .A2(n10712), .ZN(n10710) );
  NAND2_X1 U12591 ( .A1(n10716), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10646) );
  NAND2_X1 U12592 ( .A1(n10710), .A2(n10646), .ZN(n10648) );
  OAI21_X1 U12593 ( .B1(n10648), .B2(n10734), .A(n10647), .ZN(n10730) );
  XNOR2_X1 U12594 ( .A(n10730), .B(n8257), .ZN(n10649) );
  NAND2_X1 U12595 ( .A1(n10649), .A2(n15675), .ZN(n10651) );
  NOR2_X1 U12596 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13329), .ZN(n11937) );
  AOI21_X1 U12597 ( .B1(n15702), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11937), .ZN(
        n10650) );
  OAI211_X1 U12598 ( .C1(n13611), .C2(n10734), .A(n10651), .B(n10650), .ZN(
        n10652) );
  AOI21_X1 U12599 ( .B1(n15711), .B2(n10653), .A(n10652), .ZN(n10654) );
  OAI21_X1 U12600 ( .B1(n10655), .B2(n15681), .A(n10654), .ZN(P3_U3189) );
  OAI21_X1 U12601 ( .B1(n10658), .B2(n10657), .A(n10656), .ZN(n10667) );
  NAND2_X1 U12602 ( .A1(n15702), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10659) );
  OAI21_X1 U12603 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n10660), .A(n10659), .ZN(
        n10666) );
  OAI21_X1 U12604 ( .B1(n10663), .B2(n10662), .A(n10661), .ZN(n10664) );
  AND2_X1 U12605 ( .A1(n15711), .A2(n10664), .ZN(n10665) );
  AOI211_X1 U12606 ( .C1(n15675), .C2(n10667), .A(n10666), .B(n10665), .ZN(
        n10672) );
  XNOR2_X1 U12607 ( .A(n10669), .B(n10668), .ZN(n10670) );
  NAND2_X1 U12608 ( .A1(n10670), .A2(n15712), .ZN(n10671) );
  OAI211_X1 U12609 ( .C1(n13611), .C2(n10673), .A(n10672), .B(n10671), .ZN(
        P3_U3184) );
  INV_X1 U12610 ( .A(n11971), .ZN(n10724) );
  INV_X1 U12611 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U12612 ( .A1(n10675), .A2(n10674), .ZN(n10676) );
  NAND2_X1 U12613 ( .A1(n10676), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11020) );
  XNOR2_X1 U12614 ( .A(n11020), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U12615 ( .A1(n11972), .A2(P1_STATE_REG_SCAN_IN), .B1(n11702), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n10677) );
  OAI21_X1 U12616 ( .B1(n10724), .B2(n13160), .A(n10677), .ZN(P1_U3342) );
  INV_X1 U12617 ( .A(n10678), .ZN(n10679) );
  NAND3_X1 U12618 ( .A1(n13058), .A2(n10679), .A3(n15912), .ZN(n10681) );
  NAND2_X1 U12619 ( .A1(n13487), .A2(n13742), .ZN(n10680) );
  NAND2_X1 U12620 ( .A1(n10681), .A2(n10680), .ZN(n10887) );
  NOR2_X1 U12621 ( .A1(n16000), .A2(n8279), .ZN(n10682) );
  AOI21_X1 U12622 ( .B1(n16000), .B2(n10887), .A(n10682), .ZN(n10683) );
  OAI21_X1 U12623 ( .B1(n10571), .B2(n13960), .A(n10683), .ZN(P3_U3390) );
  AOI21_X1 U12624 ( .B1(n10686), .B2(n10685), .A(n10684), .ZN(n10690) );
  OAI22_X1 U12625 ( .A1(n12896), .A2(n13247), .B1(n13236), .B2(n12909), .ZN(
        n10688) );
  NOR2_X1 U12626 ( .A1(n13255), .A2(n11217), .ZN(n10687) );
  AOI211_X1 U12627 ( .C1(n10974), .C2(P3_REG3_REG_1__SCAN_IN), .A(n10688), .B(
        n10687), .ZN(n10689) );
  OAI21_X1 U12628 ( .B1(n10690), .B2(n13222), .A(n10689), .ZN(P3_U3162) );
  AOI21_X1 U12629 ( .B1(n11602), .B2(n10692), .A(n10691), .ZN(n11051) );
  XOR2_X1 U12630 ( .A(n11966), .B(n11051), .Z(n10694) );
  INV_X1 U12631 ( .A(n10694), .ZN(n10696) );
  INV_X1 U12632 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10693) );
  NAND2_X1 U12633 ( .A1(n10694), .A2(n10693), .ZN(n11050) );
  INV_X1 U12634 ( .A(n11050), .ZN(n10695) );
  AOI21_X1 U12635 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n10696), .A(n10695), 
        .ZN(n10706) );
  INV_X1 U12636 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10697) );
  MUX2_X1 U12637 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10697), .S(n11966), .Z(
        n10700) );
  AOI21_X1 U12638 ( .B1(n11743), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10698), 
        .ZN(n10699) );
  NAND2_X1 U12639 ( .A1(n10699), .A2(n10700), .ZN(n11056) );
  OAI21_X1 U12640 ( .B1(n10700), .B2(n10699), .A(n11056), .ZN(n10704) );
  NAND2_X1 U12641 ( .A1(n15741), .A2(n11966), .ZN(n10701) );
  NAND2_X1 U12642 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n12272)
         );
  OAI211_X1 U12643 ( .C1(n10702), .C2(n15145), .A(n10701), .B(n12272), .ZN(
        n10703) );
  AOI21_X1 U12644 ( .B1(n10704), .B2(n15730), .A(n10703), .ZN(n10705) );
  OAI21_X1 U12645 ( .B1(n10706), .B2(n15135), .A(n10705), .ZN(P1_U3255) );
  OAI21_X1 U12646 ( .B1(n10709), .B2(n10708), .A(n10707), .ZN(n10722) );
  INV_X1 U12647 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n13364) );
  NOR2_X1 U12648 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13364), .ZN(n11858) );
  AOI21_X1 U12649 ( .B1(n15702), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11858), .ZN(
        n10715) );
  OAI21_X1 U12650 ( .B1(n10712), .B2(n10711), .A(n10710), .ZN(n10713) );
  NAND2_X1 U12651 ( .A1(n15675), .A2(n10713), .ZN(n10714) );
  OAI211_X1 U12652 ( .C1(n13611), .C2(n10716), .A(n10715), .B(n10714), .ZN(
        n10721) );
  XOR2_X1 U12653 ( .A(n10717), .B(n10718), .Z(n10719) );
  NOR2_X1 U12654 ( .A1(n10719), .A2(n15681), .ZN(n10720) );
  AOI211_X1 U12655 ( .C1(n15711), .C2(n10722), .A(n10721), .B(n10720), .ZN(
        n10723) );
  INV_X1 U12656 ( .A(n10723), .ZN(P3_U3188) );
  INV_X1 U12657 ( .A(n12367), .ZN(n12108) );
  OAI222_X1 U12658 ( .A1(n13150), .A2(n7841), .B1(n14477), .B2(n10724), .C1(
        n12108), .C2(P2_U3088), .ZN(P2_U3314) );
  MUX2_X1 U12659 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13087), .Z(n10978) );
  XNOR2_X1 U12660 ( .A(n10978), .B(n10988), .ZN(n10979) );
  INV_X1 U12661 ( .A(n10725), .ZN(n10726) );
  AOI22_X1 U12662 ( .A1(n10729), .A2(n10728), .B1(n10727), .B2(n10726), .ZN(
        n10980) );
  XOR2_X1 U12663 ( .A(n10979), .B(n10980), .Z(n10746) );
  NOR2_X1 U12664 ( .A1(n8257), .A2(n10730), .ZN(n10731) );
  NAND2_X1 U12665 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10988), .ZN(n10732) );
  OAI21_X1 U12666 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10988), .A(n10732), .ZN(
        n10985) );
  XNOR2_X1 U12667 ( .A(n10986), .B(n10985), .ZN(n10744) );
  AOI22_X1 U12668 ( .A1(n10733), .A2(n8244), .B1(P3_REG2_REG_8__SCAN_IN), .B2(
        n10988), .ZN(n10739) );
  NAND2_X1 U12669 ( .A1(n10735), .A2(n10734), .ZN(n10737) );
  NAND2_X1 U12670 ( .A1(n10739), .A2(n10738), .ZN(n10981) );
  OAI21_X1 U12671 ( .B1(n10739), .B2(n10738), .A(n10981), .ZN(n10740) );
  NAND2_X1 U12672 ( .A1(n10740), .A2(n15711), .ZN(n10742) );
  NOR2_X1 U12673 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13454), .ZN(n12087) );
  AOI21_X1 U12674 ( .B1(n15702), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12087), .ZN(
        n10741) );
  OAI211_X1 U12675 ( .C1(n13611), .C2(n10988), .A(n10742), .B(n10741), .ZN(
        n10743) );
  AOI21_X1 U12676 ( .B1(n15675), .B2(n10744), .A(n10743), .ZN(n10745) );
  OAI21_X1 U12677 ( .B1(n10746), .B2(n15681), .A(n10745), .ZN(P3_U3190) );
  NAND2_X1 U12678 ( .A1(n12711), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n10752) );
  INV_X1 U12679 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10747) );
  OR2_X1 U12680 ( .A1(n12686), .A2(n10747), .ZN(n10751) );
  NAND2_X1 U12681 ( .A1(n10812), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10832) );
  NAND2_X1 U12682 ( .A1(n11037), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11279) );
  NAND2_X1 U12683 ( .A1(n12011), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12183) );
  OAI21_X1 U12684 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n10748), .A(n12660), 
        .ZN(n15266) );
  OR2_X1 U12685 ( .A1(n7189), .A2(n15266), .ZN(n10750) );
  INV_X1 U12686 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n15259) );
  OR2_X1 U12687 ( .A1(n12705), .A2(n15259), .ZN(n10749) );
  NAND4_X1 U12688 ( .A1(n10752), .A2(n10751), .A3(n10750), .A4(n10749), .ZN(
        n15271) );
  NAND2_X1 U12689 ( .A1(n15271), .A2(P1_U4016), .ZN(n10753) );
  OAI21_X1 U12690 ( .B1(P1_U4016), .B2(n10754), .A(n10753), .ZN(P1_U3583) );
  NAND2_X1 U12691 ( .A1(n15054), .A2(n11286), .ZN(n10758) );
  NAND2_X1 U12692 ( .A1(n11271), .A2(n14581), .ZN(n10757) );
  NAND2_X1 U12693 ( .A1(n10758), .A2(n10757), .ZN(n10759) );
  XNOR2_X1 U12694 ( .A(n10759), .B(n14584), .ZN(n10760) );
  AOI22_X1 U12695 ( .A1(n15054), .A2(n14563), .B1(n11271), .B2(n11286), .ZN(
        n10761) );
  NAND2_X1 U12696 ( .A1(n10760), .A2(n10761), .ZN(n10904) );
  INV_X1 U12697 ( .A(n10760), .ZN(n10763) );
  INV_X1 U12698 ( .A(n10761), .ZN(n10762) );
  NAND2_X1 U12699 ( .A1(n10763), .A2(n10762), .ZN(n10764) );
  NAND2_X1 U12700 ( .A1(n10904), .A2(n10764), .ZN(n10768) );
  NAND2_X1 U12701 ( .A1(n10766), .A2(n10765), .ZN(n10905) );
  INV_X1 U12702 ( .A(n10905), .ZN(n10767) );
  AOI21_X1 U12703 ( .B1(n10769), .B2(n10768), .A(n10767), .ZN(n10775) );
  INV_X1 U12704 ( .A(n7381), .ZN(n10770) );
  OAI22_X1 U12705 ( .A1(n10770), .A2(n14743), .B1(n14747), .B2(n14607), .ZN(
        n10773) );
  INV_X1 U12706 ( .A(n14751), .ZN(n14725) );
  NOR2_X1 U12707 ( .A1(n14725), .A2(n10771), .ZN(n10772) );
  AOI211_X1 U12708 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n12783), .A(n10773), .B(
        n10772), .ZN(n10774) );
  OAI21_X1 U12709 ( .B1(n10775), .B2(n14753), .A(n10774), .ZN(P1_U3222) );
  INV_X1 U12710 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10787) );
  XOR2_X1 U12711 ( .A(n10776), .B(n10777), .Z(n11369) );
  INV_X1 U12712 ( .A(n11369), .ZN(n10785) );
  XOR2_X1 U12713 ( .A(n10778), .B(n10777), .Z(n10780) );
  AOI22_X1 U12714 ( .A1(n14355), .A2(n14077), .B1(n14079), .B2(n14353), .ZN(
        n10779) );
  OAI21_X1 U12715 ( .B1(n10780), .B2(n14298), .A(n10779), .ZN(n10781) );
  AOI21_X1 U12716 ( .B1(n11369), .B2(n14305), .A(n10781), .ZN(n11371) );
  INV_X1 U12717 ( .A(n11456), .ZN(n10782) );
  AOI21_X1 U12718 ( .B1(n10947), .B2(n10783), .A(n10782), .ZN(n11364) );
  AOI22_X1 U12719 ( .A1(n11364), .A2(n14445), .B1(n15841), .B2(n10947), .ZN(
        n10784) );
  OAI211_X1 U12720 ( .C1(n14449), .C2(n10785), .A(n11371), .B(n10784), .ZN(
        n10788) );
  NAND2_X1 U12721 ( .A1(n10788), .A2(n14451), .ZN(n10786) );
  OAI21_X1 U12722 ( .B1(n14451), .B2(n10787), .A(n10786), .ZN(P2_U3504) );
  INV_X1 U12723 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10790) );
  NAND2_X1 U12724 ( .A1(n10788), .A2(n14469), .ZN(n10789) );
  OAI21_X1 U12725 ( .B1(n14469), .B2(n10790), .A(n10789), .ZN(P2_U3445) );
  XOR2_X1 U12726 ( .A(n10791), .B(n10792), .Z(n10803) );
  XNOR2_X1 U12727 ( .A(n10793), .B(P3_REG2_REG_5__SCAN_IN), .ZN(n10801) );
  NOR2_X1 U12728 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10794), .ZN(n11431) );
  AOI21_X1 U12729 ( .B1(n10796), .B2(n10795), .A(n15718), .ZN(n10797) );
  AOI211_X1 U12730 ( .C1(n15702), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n11431), .B(
        n10797), .ZN(n10798) );
  OAI21_X1 U12731 ( .B1(n10799), .B2(n13611), .A(n10798), .ZN(n10800) );
  AOI21_X1 U12732 ( .B1(n15711), .B2(n10801), .A(n10800), .ZN(n10802) );
  OAI21_X1 U12733 ( .B1(n10803), .B2(n15681), .A(n10802), .ZN(P3_U3187) );
  OR2_X1 U12734 ( .A1(n15052), .A2(n14776), .ZN(n10804) );
  NAND2_X1 U12735 ( .A1(n10805), .A2(n10804), .ZN(n11686) );
  NAND2_X1 U12736 ( .A1(n7378), .A2(n10806), .ZN(n10810) );
  OR2_X1 U12737 ( .A1(n12641), .A2(n15724), .ZN(n10809) );
  OR2_X1 U12738 ( .A1(n14947), .A2(n10807), .ZN(n10808) );
  XNOR2_X1 U12739 ( .A(n15051), .B(n15790), .ZN(n11696) );
  NAND2_X1 U12740 ( .A1(n11686), .A2(n8092), .ZN(n11685) );
  OR2_X1 U12741 ( .A1(n15051), .A2(n14783), .ZN(n10811) );
  NAND2_X1 U12742 ( .A1(n14924), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n10816) );
  OR2_X1 U12743 ( .A1(n14928), .A2(n10170), .ZN(n10815) );
  OAI21_X1 U12744 ( .B1(n10812), .B2(P1_REG3_REG_5__SCAN_IN), .A(n10832), .ZN(
        n11705) );
  OR2_X1 U12745 ( .A1(n7189), .A2(n11705), .ZN(n10814) );
  OR2_X1 U12746 ( .A1(n12705), .A2(n11706), .ZN(n10813) );
  NAND4_X1 U12747 ( .A1(n10816), .A2(n10815), .A3(n10814), .A4(n10813), .ZN(
        n15050) );
  NAND2_X1 U12748 ( .A1(n10817), .A2(n14944), .ZN(n10820) );
  INV_X2 U12749 ( .A(n14947), .ZN(n12597) );
  AOI22_X1 U12750 ( .A1(n12597), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7182), 
        .B2(n10818), .ZN(n10819) );
  XNOR2_X1 U12751 ( .A(n15050), .B(n11129), .ZN(n10829) );
  OAI21_X1 U12752 ( .B1(n10821), .B2(n10829), .A(n11128), .ZN(n11711) );
  NAND2_X1 U12753 ( .A1(n11688), .A2(n15790), .ZN(n11687) );
  INV_X1 U12754 ( .A(n15932), .ZN(n15354) );
  AOI21_X1 U12755 ( .B1(n11687), .B2(n14787), .A(n15354), .ZN(n10822) );
  NAND2_X1 U12756 ( .A1(n10822), .A2(n11136), .ZN(n11709) );
  OAI21_X1 U12757 ( .B1(n11129), .B2(n15970), .A(n11709), .ZN(n10840) );
  NAND2_X1 U12758 ( .A1(n15052), .A2(n10825), .ZN(n10823) );
  NAND2_X1 U12759 ( .A1(n10824), .A2(n10823), .ZN(n10827) );
  OR2_X1 U12760 ( .A1(n15052), .A2(n10825), .ZN(n10826) );
  NAND2_X1 U12761 ( .A1(n10827), .A2(n10826), .ZN(n11695) );
  INV_X1 U12762 ( .A(n11696), .ZN(n14954) );
  NAND2_X1 U12763 ( .A1(n15051), .A2(n15790), .ZN(n10828) );
  INV_X1 U12764 ( .A(n10829), .ZN(n14952) );
  OAI211_X1 U12765 ( .C1(n10830), .C2(n14952), .A(n11131), .B(n15988), .ZN(
        n10839) );
  NAND2_X1 U12766 ( .A1(n14924), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10837) );
  OR2_X1 U12767 ( .A1(n12705), .A2(n10208), .ZN(n10836) );
  AND2_X1 U12768 ( .A1(n10832), .A2(n10831), .ZN(n10833) );
  OR2_X1 U12769 ( .A1(n10833), .A2(n11037), .ZN(n15811) );
  OR2_X1 U12770 ( .A1(n12704), .A2(n15811), .ZN(n10835) );
  OR2_X1 U12771 ( .A1(n14928), .A2(n11140), .ZN(n10834) );
  AOI22_X1 U12772 ( .A1(n15049), .A2(n15342), .B1(n15289), .B2(n15051), .ZN(
        n10838) );
  NAND2_X1 U12773 ( .A1(n10839), .A2(n10838), .ZN(n11704) );
  AOI211_X1 U12774 ( .C1(n15973), .C2(n11711), .A(n10840), .B(n11704), .ZN(
        n10940) );
  NAND2_X1 U12775 ( .A1(n15990), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10841) );
  OAI21_X1 U12776 ( .B1(n10940), .B2(n15990), .A(n10841), .ZN(P1_U3533) );
  INV_X1 U12777 ( .A(n10842), .ZN(n10843) );
  OAI222_X1 U12778 ( .A1(n13610), .A2(P3_U3151), .B1(n13969), .B2(n13403), 
        .C1(n13157), .C2(n10843), .ZN(P3_U3276) );
  NAND2_X1 U12779 ( .A1(n14054), .A2(n12832), .ZN(n14038) );
  NOR3_X1 U12780 ( .A1(n14038), .A2(n10846), .A3(n10845), .ZN(n10847) );
  AOI21_X1 U12781 ( .B1(n14054), .B2(n10848), .A(n10847), .ZN(n10860) );
  XNOR2_X1 U12782 ( .A(n11474), .B(n12804), .ZN(n11067) );
  NAND2_X1 U12783 ( .A1(n14079), .A2(n12832), .ZN(n10943) );
  XNOR2_X1 U12784 ( .A(n11067), .B(n10943), .ZN(n10859) );
  AND2_X1 U12785 ( .A1(n10859), .A2(n10849), .ZN(n10850) );
  NAND2_X1 U12786 ( .A1(n10851), .A2(n10850), .ZN(n10946) );
  INV_X1 U12787 ( .A(n10946), .ZN(n11069) );
  INV_X1 U12788 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10852) );
  OAI22_X1 U12789 ( .A1(n14002), .A2(n10853), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10852), .ZN(n10857) );
  OAI22_X1 U12790 ( .A1(n14044), .A2(n10855), .B1(n14030), .B2(n10854), .ZN(
        n10856) );
  AOI211_X1 U12791 ( .C1(n11069), .C2(n14054), .A(n10857), .B(n10856), .ZN(
        n10858) );
  OAI21_X1 U12792 ( .B1(n10860), .B2(n10859), .A(n10858), .ZN(P2_U3202) );
  AOI21_X1 U12793 ( .B1(n10868), .B2(P2_REG2_REG_4__SCAN_IN), .A(n10861), .ZN(
        n15532) );
  XNOR2_X1 U12794 ( .A(n15535), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n15531) );
  NOR2_X1 U12795 ( .A1(n15532), .A2(n15531), .ZN(n15530) );
  INV_X1 U12796 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10862) );
  MUX2_X1 U12797 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10862), .S(n15546), .Z(
        n10863) );
  INV_X1 U12798 ( .A(n10863), .ZN(n15542) );
  NOR2_X1 U12799 ( .A1(n15543), .A2(n15542), .ZN(n15541) );
  AOI21_X1 U12800 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n15546), .A(n15541), .ZN(
        n15554) );
  XNOR2_X1 U12801 ( .A(n15557), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n15553) );
  NOR2_X1 U12802 ( .A1(n15554), .A2(n15553), .ZN(n15552) );
  INV_X1 U12803 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10864) );
  MUX2_X1 U12804 ( .A(n10864), .B(P2_REG2_REG_8__SCAN_IN), .S(n11110), .Z(
        n10865) );
  NOR2_X1 U12805 ( .A1(n10866), .A2(n10865), .ZN(n11106) );
  AOI211_X1 U12806 ( .C1(n10866), .C2(n10865), .A(n15592), .B(n11106), .ZN(
        n10879) );
  AOI21_X1 U12807 ( .B1(n10868), .B2(P2_REG1_REG_4__SCAN_IN), .A(n10867), .ZN(
        n15529) );
  XNOR2_X1 U12808 ( .A(n15535), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n15528) );
  INV_X1 U12809 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10869) );
  MUX2_X1 U12810 ( .A(n10869), .B(P2_REG1_REG_6__SCAN_IN), .S(n15546), .Z(
        n15539) );
  INV_X1 U12811 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10870) );
  MUX2_X1 U12812 ( .A(n10870), .B(P2_REG1_REG_7__SCAN_IN), .S(n15557), .Z(
        n15550) );
  NOR2_X1 U12813 ( .A1(n15551), .A2(n15550), .ZN(n15549) );
  INV_X1 U12814 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10871) );
  MUX2_X1 U12815 ( .A(n10871), .B(P2_REG1_REG_8__SCAN_IN), .S(n11110), .Z(
        n10872) );
  AOI211_X1 U12816 ( .C1(n10873), .C2(n10872), .A(n15588), .B(n11109), .ZN(
        n10878) );
  NAND2_X1 U12817 ( .A1(n15522), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10875) );
  NAND2_X1 U12818 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10874) );
  OAI211_X1 U12819 ( .C1(n14148), .C2(n10876), .A(n10875), .B(n10874), .ZN(
        n10877) );
  OR3_X1 U12820 ( .A1(n10879), .A2(n10878), .A3(n10877), .ZN(P2_U3222) );
  AOI21_X1 U12821 ( .B1(n14054), .B2(n10880), .A(n14035), .ZN(n10886) );
  NOR2_X1 U12822 ( .A1(n10881), .A2(P2_U3088), .ZN(n13126) );
  INV_X1 U12823 ( .A(n13126), .ZN(n10882) );
  AOI22_X1 U12824 ( .A1(n13142), .A2(n9000), .B1(n10882), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10884) );
  INV_X1 U12825 ( .A(n14038), .ZN(n13994) );
  NAND3_X1 U12826 ( .A1(n13994), .A2(n9450), .A3(n13125), .ZN(n10883) );
  OAI211_X1 U12827 ( .C1(n10886), .C2(n10885), .A(n10884), .B(n10883), .ZN(
        P2_U3204) );
  INV_X1 U12828 ( .A(n10887), .ZN(n10900) );
  MUX2_X1 U12829 ( .A(n10888), .B(n10900), .S(n15997), .Z(n10889) );
  OAI21_X1 U12830 ( .B1(n10571), .B2(n13905), .A(n10889), .ZN(P3_U3459) );
  INV_X1 U12831 ( .A(n10890), .ZN(n10891) );
  NOR2_X1 U12832 ( .A1(n13965), .A2(n10891), .ZN(n10893) );
  MUX2_X1 U12833 ( .A(n13965), .B(n10893), .S(n10892), .Z(n10894) );
  INV_X1 U12834 ( .A(n10899), .ZN(n10896) );
  INV_X1 U12835 ( .A(n13084), .ZN(n11222) );
  NOR2_X1 U12836 ( .A1(n15912), .A2(n11222), .ZN(n11680) );
  INV_X1 U12837 ( .A(n15806), .ZN(n13816) );
  NOR2_X1 U12838 ( .A1(n15912), .A2(n13084), .ZN(n10897) );
  AOI22_X1 U12839 ( .A1(n13816), .A2(n12895), .B1(n13802), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10903) );
  MUX2_X1 U12840 ( .A(n10901), .B(n10900), .S(n15810), .Z(n10902) );
  NAND2_X1 U12841 ( .A1(n10903), .A2(n10902), .ZN(P3_U3233) );
  NAND2_X1 U12842 ( .A1(n10905), .A2(n10904), .ZN(n12777) );
  NAND2_X1 U12843 ( .A1(n7377), .A2(n11286), .ZN(n10907) );
  NAND2_X1 U12844 ( .A1(n14769), .A2(n14581), .ZN(n10906) );
  NAND2_X1 U12845 ( .A1(n10907), .A2(n10906), .ZN(n10908) );
  XNOR2_X1 U12846 ( .A(n10908), .B(n14628), .ZN(n10909) );
  INV_X1 U12847 ( .A(n10909), .ZN(n10911) );
  NAND2_X1 U12848 ( .A1(n10911), .A2(n10910), .ZN(n10912) );
  NAND2_X1 U12849 ( .A1(n15052), .A2(n11286), .ZN(n10914) );
  NAND2_X1 U12850 ( .A1(n14776), .A2(n14581), .ZN(n10913) );
  NAND2_X1 U12851 ( .A1(n10914), .A2(n10913), .ZN(n10915) );
  XNOR2_X1 U12852 ( .A(n10915), .B(n14628), .ZN(n10916) );
  AOI22_X1 U12853 ( .A1(n15052), .A2(n14563), .B1(n14776), .B2(n14587), .ZN(
        n10917) );
  XNOR2_X1 U12854 ( .A(n10916), .B(n10917), .ZN(n14606) );
  INV_X1 U12855 ( .A(n10916), .ZN(n10918) );
  OR2_X1 U12856 ( .A1(n10918), .A2(n10917), .ZN(n10922) );
  AOI22_X1 U12857 ( .A1(n15051), .A2(n14563), .B1(n14783), .B2(n14587), .ZN(
        n10921) );
  AND2_X1 U12858 ( .A1(n10922), .A2(n10921), .ZN(n10919) );
  INV_X1 U12859 ( .A(n15051), .ZN(n14784) );
  OAI22_X1 U12860 ( .A1(n14784), .A2(n14572), .B1(n15790), .B2(n14627), .ZN(
        n10920) );
  XOR2_X1 U12861 ( .A(n14628), .B(n10920), .Z(n10997) );
  AOI21_X1 U12862 ( .B1(n14604), .B2(n10922), .A(n10921), .ZN(n10996) );
  NOR2_X2 U12863 ( .A1(n10999), .A2(n10996), .ZN(n11027) );
  NAND2_X1 U12864 ( .A1(n15050), .A2(n14587), .ZN(n10924) );
  OR2_X1 U12865 ( .A1(n11129), .A2(n14627), .ZN(n10923) );
  NAND2_X1 U12866 ( .A1(n10924), .A2(n10923), .ZN(n10925) );
  XNOR2_X1 U12867 ( .A(n10925), .B(n14584), .ZN(n10928) );
  NAND2_X1 U12868 ( .A1(n15050), .A2(n14563), .ZN(n10927) );
  OR2_X1 U12869 ( .A1(n11129), .A2(n14572), .ZN(n10926) );
  AND2_X1 U12870 ( .A1(n10927), .A2(n10926), .ZN(n10929) );
  AND2_X1 U12871 ( .A1(n10928), .A2(n10929), .ZN(n11025) );
  INV_X1 U12872 ( .A(n11025), .ZN(n10932) );
  INV_X1 U12873 ( .A(n10928), .ZN(n10931) );
  INV_X1 U12874 ( .A(n10929), .ZN(n10930) );
  NAND2_X1 U12875 ( .A1(n10931), .A2(n10930), .ZN(n11026) );
  NAND2_X1 U12876 ( .A1(n10932), .A2(n11026), .ZN(n10933) );
  XNOR2_X1 U12877 ( .A(n11027), .B(n10933), .ZN(n10939) );
  OAI21_X1 U12878 ( .B1(n14743), .B2(n14784), .A(n10934), .ZN(n10937) );
  OAI22_X1 U12879 ( .A1(n11564), .A2(n14747), .B1(n14746), .B2(n11705), .ZN(
        n10936) );
  AOI211_X1 U12880 ( .C1(n14751), .C2(n14787), .A(n10937), .B(n10936), .ZN(
        n10938) );
  OAI21_X1 U12881 ( .B1(n10939), .B2(n14753), .A(n10938), .ZN(P1_U3227) );
  INV_X1 U12882 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10942) );
  OR2_X1 U12883 ( .A1(n10940), .A2(n15992), .ZN(n10941) );
  OAI21_X1 U12884 ( .B1(n15994), .B2(n10942), .A(n10941), .ZN(P1_U3474) );
  INV_X1 U12885 ( .A(n11067), .ZN(n10944) );
  NAND2_X1 U12886 ( .A1(n10944), .A2(n10943), .ZN(n10945) );
  NAND2_X1 U12887 ( .A1(n10946), .A2(n10945), .ZN(n10948) );
  INV_X2 U12888 ( .A(n11779), .ZN(n12804) );
  XNOR2_X1 U12889 ( .A(n10947), .B(n12804), .ZN(n10949) );
  NAND2_X1 U12890 ( .A1(n14078), .A2(n12832), .ZN(n10950) );
  XNOR2_X1 U12891 ( .A(n10949), .B(n10950), .ZN(n11068) );
  NAND2_X1 U12892 ( .A1(n10948), .A2(n11068), .ZN(n11073) );
  INV_X1 U12893 ( .A(n10949), .ZN(n10951) );
  NAND2_X1 U12894 ( .A1(n10951), .A2(n10950), .ZN(n10952) );
  XNOR2_X1 U12895 ( .A(n11455), .B(n12804), .ZN(n10953) );
  AND2_X1 U12896 ( .A1(n14077), .A2(n12832), .ZN(n10954) );
  NAND2_X1 U12897 ( .A1(n10953), .A2(n10954), .ZN(n10957) );
  INV_X1 U12898 ( .A(n10953), .ZN(n11093) );
  INV_X1 U12899 ( .A(n10954), .ZN(n10955) );
  NAND2_X1 U12900 ( .A1(n11093), .A2(n10955), .ZN(n10956) );
  NAND2_X1 U12901 ( .A1(n10957), .A2(n10956), .ZN(n11009) );
  XNOR2_X1 U12902 ( .A(n15840), .B(n12804), .ZN(n10959) );
  NAND2_X1 U12903 ( .A1(n14076), .A2(n12832), .ZN(n10960) );
  XNOR2_X1 U12904 ( .A(n10959), .B(n10960), .ZN(n11104) );
  AND2_X1 U12905 ( .A1(n11104), .A2(n10957), .ZN(n10958) );
  INV_X1 U12906 ( .A(n10959), .ZN(n10966) );
  XNOR2_X1 U12907 ( .A(n11389), .B(n12804), .ZN(n11775) );
  NAND2_X1 U12908 ( .A1(n14075), .A2(n12832), .ZN(n11776) );
  NAND2_X1 U12909 ( .A1(n14074), .A2(n14355), .ZN(n10962) );
  NAND2_X1 U12910 ( .A1(n14076), .A2(n14353), .ZN(n10961) );
  AND2_X1 U12911 ( .A1(n10962), .A2(n10961), .ZN(n11379) );
  OAI22_X1 U12912 ( .A1(n14002), .A2(n11379), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10963), .ZN(n10965) );
  NOR2_X1 U12913 ( .A1(n14044), .A2(n15857), .ZN(n10964) );
  AOI211_X1 U12914 ( .C1(n14046), .C2(n11381), .A(n10965), .B(n10964), .ZN(
        n10969) );
  OAI22_X1 U12915 ( .A1(n14038), .A2(n11011), .B1(n10966), .B2(n10844), .ZN(
        n10967) );
  NAND3_X1 U12916 ( .A1(n11100), .A2(n7348), .A3(n10967), .ZN(n10968) );
  OAI211_X1 U12917 ( .C1(n10844), .C2(n11778), .A(n10969), .B(n10968), .ZN(
        P2_U3193) );
  AOI21_X1 U12918 ( .B1(n10971), .B2(n10970), .A(n11086), .ZN(n10976) );
  INV_X1 U12919 ( .A(n13247), .ZN(n13198) );
  AOI22_X1 U12920 ( .A1(n13198), .A2(n13487), .B1(n13245), .B2(n13485), .ZN(
        n10972) );
  OAI21_X1 U12921 ( .B1(n11208), .B2(n13255), .A(n10972), .ZN(n10973) );
  AOI21_X1 U12922 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10974), .A(n10973), .ZN(
        n10975) );
  OAI21_X1 U12923 ( .B1(n10976), .B2(n13222), .A(n10975), .ZN(P3_U3177) );
  MUX2_X1 U12924 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13087), .Z(n11539) );
  XNOR2_X1 U12925 ( .A(n11539), .B(n11541), .ZN(n11542) );
  XOR2_X1 U12926 ( .A(n11542), .B(n11543), .Z(n10994) );
  NAND2_X1 U12927 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10988), .ZN(n10982) );
  NAND2_X1 U12928 ( .A1(n10982), .A2(n10981), .ZN(n11555) );
  XNOR2_X1 U12929 ( .A(n11555), .B(n11541), .ZN(n10983) );
  NAND2_X1 U12930 ( .A1(P3_REG2_REG_9__SCAN_IN), .A2(n10983), .ZN(n11556) );
  OAI21_X1 U12931 ( .B1(n10983), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11556), .ZN(
        n10992) );
  NOR2_X1 U12932 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8154), .ZN(n12170) );
  AOI21_X1 U12933 ( .B1(n15702), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12170), .ZN(
        n10984) );
  OAI21_X1 U12934 ( .B1(n13611), .B2(n11554), .A(n10984), .ZN(n10991) );
  NOR2_X1 U12935 ( .A1(n10986), .A2(n10985), .ZN(n10987) );
  XOR2_X1 U12936 ( .A(n8372), .B(n11546), .Z(n10989) );
  NOR2_X1 U12937 ( .A1(n10989), .A2(n15718), .ZN(n10990) );
  AOI211_X1 U12938 ( .C1(n15711), .C2(n10992), .A(n10991), .B(n10990), .ZN(
        n10993) );
  OAI21_X1 U12939 ( .B1(n10994), .B2(n15681), .A(n10993), .ZN(P3_U3191) );
  INV_X1 U12940 ( .A(n10995), .ZN(n11001) );
  INV_X1 U12941 ( .A(n10996), .ZN(n10998) );
  AOI21_X1 U12942 ( .B1(n10999), .B2(n10998), .A(n10997), .ZN(n11000) );
  AOI21_X1 U12943 ( .B1(n11027), .B2(n11001), .A(n11000), .ZN(n11007) );
  NAND2_X1 U12944 ( .A1(n15050), .A2(n15342), .ZN(n11003) );
  NAND2_X1 U12945 ( .A1(n15052), .A2(n15289), .ZN(n11002) );
  NAND2_X1 U12946 ( .A1(n11003), .A2(n11002), .ZN(n11691) );
  INV_X1 U12947 ( .A(n14665), .ZN(n14694) );
  AOI22_X1 U12948 ( .A1(n11691), .A2(n14694), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11004) );
  OAI21_X1 U12949 ( .B1(n11689), .B2(n14746), .A(n11004), .ZN(n11005) );
  AOI21_X1 U12950 ( .B1(n14751), .B2(n14783), .A(n11005), .ZN(n11006) );
  OAI21_X1 U12951 ( .B1(n11007), .B2(n14753), .A(n11006), .ZN(P1_U3230) );
  INV_X1 U12952 ( .A(n11008), .ZN(n11095) );
  AOI211_X1 U12953 ( .C1(n11010), .C2(n11009), .A(n10844), .B(n11095), .ZN(
        n11016) );
  INV_X1 U12954 ( .A(n11455), .ZN(n15820) );
  OAI22_X1 U12955 ( .A1(n14044), .A2(n15820), .B1(n14050), .B2(n11011), .ZN(
        n11015) );
  NAND2_X1 U12956 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n15547) );
  NAND2_X1 U12957 ( .A1(n14046), .A2(n11460), .ZN(n11012) );
  OAI211_X1 U12958 ( .C1(n14031), .C2(n11013), .A(n15547), .B(n11012), .ZN(
        n11014) );
  OR3_X1 U12959 ( .A1(n11016), .A2(n11015), .A3(n11014), .ZN(P2_U3211) );
  NAND2_X1 U12960 ( .A1(n13265), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11017) );
  OAI21_X1 U12961 ( .B1(n13634), .B2(n13265), .A(n11017), .ZN(P3_U3520) );
  INV_X1 U12962 ( .A(n12005), .ZN(n11023) );
  INV_X1 U12963 ( .A(n14084), .ZN(n12376) );
  OAI222_X1 U12964 ( .A1(n13150), .A2(n11018), .B1(n14477), .B2(n11023), .C1(
        P2_U3088), .C2(n12376), .ZN(P2_U3313) );
  INV_X1 U12965 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n11019) );
  NAND2_X1 U12966 ( .A1(n11020), .A2(n11019), .ZN(n11021) );
  NAND2_X1 U12967 ( .A1(n11021), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11022) );
  XNOR2_X1 U12968 ( .A(n11022), .B(P1_IR_REG_14__SCAN_IN), .ZN(n12006) );
  INV_X1 U12969 ( .A(n12006), .ZN(n11488) );
  OAI222_X1 U12970 ( .A1(n15476), .A2(n11024), .B1(n13160), .B2(n11023), .C1(
        P1_U3086), .C2(n11488), .ZN(P1_U3341) );
  OR2_X1 U12971 ( .A1(n11564), .A2(n14626), .ZN(n11033) );
  NAND2_X1 U12972 ( .A1(n11028), .A2(n14944), .ZN(n11031) );
  AOI22_X1 U12973 ( .A1(n12597), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12596), 
        .B2(n11029), .ZN(n11030) );
  AND2_X2 U12974 ( .A1(n11031), .A2(n11030), .ZN(n11567) );
  OR2_X1 U12975 ( .A1(n11567), .A2(n14572), .ZN(n11032) );
  NAND2_X1 U12976 ( .A1(n11033), .A2(n11032), .ZN(n11288) );
  OR2_X1 U12977 ( .A1(n11567), .A2(n14627), .ZN(n11034) );
  OAI21_X1 U12978 ( .B1(n11564), .B2(n14572), .A(n11034), .ZN(n11035) );
  XNOR2_X1 U12979 ( .A(n11035), .B(n14628), .ZN(n11287) );
  XOR2_X1 U12980 ( .A(n11288), .B(n11287), .Z(n11290) );
  XNOR2_X1 U12981 ( .A(n11291), .B(n11290), .ZN(n11049) );
  INV_X2 U12982 ( .A(n11567), .ZN(n15813) );
  NAND2_X1 U12983 ( .A1(n12711), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11042) );
  INV_X1 U12984 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11036) );
  OR2_X1 U12985 ( .A1(n12686), .A2(n11036), .ZN(n11041) );
  OR2_X1 U12986 ( .A1(n11037), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11038) );
  NAND2_X1 U12987 ( .A1(n11279), .A2(n11038), .ZN(n11573) );
  OR2_X1 U12988 ( .A1(n7189), .A2(n11573), .ZN(n11040) );
  OR2_X1 U12989 ( .A1(n12705), .A2(n11571), .ZN(n11039) );
  OR2_X1 U12990 ( .A1(n11617), .A2(n15195), .ZN(n11044) );
  NAND2_X1 U12991 ( .A1(n15050), .A2(n15289), .ZN(n11043) );
  NAND2_X1 U12992 ( .A1(n11044), .A2(n11043), .ZN(n11135) );
  NAND2_X1 U12993 ( .A1(n11135), .A2(n14694), .ZN(n11046) );
  OAI211_X1 U12994 ( .C1(n14746), .C2(n15811), .A(n11046), .B(n11045), .ZN(
        n11047) );
  AOI21_X1 U12995 ( .B1(n14751), .B2(n15813), .A(n11047), .ZN(n11048) );
  OAI21_X1 U12996 ( .B1(n11049), .B2(n14753), .A(n11048), .ZN(P1_U3239) );
  OAI21_X1 U12997 ( .B1(n11966), .B2(n11051), .A(n11050), .ZN(n11160) );
  INV_X1 U12998 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15965) );
  MUX2_X1 U12999 ( .A(n15965), .B(P1_REG1_REG_13__SCAN_IN), .S(n11972), .Z(
        n11159) );
  NAND2_X1 U13000 ( .A1(n11972), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11053) );
  INV_X1 U13001 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15978) );
  MUX2_X1 U13002 ( .A(n15978), .B(P1_REG1_REG_14__SCAN_IN), .S(n12006), .Z(
        n11052) );
  AOI21_X1 U13003 ( .B1(n11157), .B2(n11053), .A(n11052), .ZN(n11483) );
  INV_X1 U13004 ( .A(n11483), .ZN(n11055) );
  NAND3_X1 U13005 ( .A1(n11157), .A2(n11053), .A3(n11052), .ZN(n11054) );
  NAND3_X1 U13006 ( .A1(n11055), .A2(n15739), .A3(n11054), .ZN(n11062) );
  NAND2_X1 U13007 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n12431)
         );
  INV_X1 U13008 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11979) );
  INV_X1 U13009 ( .A(n11972), .ZN(n11166) );
  OAI21_X1 U13010 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n11966), .A(n11056), 
        .ZN(n11164) );
  MUX2_X1 U13011 ( .A(n11979), .B(P1_REG2_REG_13__SCAN_IN), .S(n11972), .Z(
        n11163) );
  OAI21_X1 U13012 ( .B1(n11979), .B2(n11166), .A(n11161), .ZN(n11058) );
  INV_X1 U13013 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11989) );
  MUX2_X1 U13014 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11989), .S(n12006), .Z(
        n11057) );
  NAND2_X1 U13015 ( .A1(n11058), .A2(n11057), .ZN(n11487) );
  OAI211_X1 U13016 ( .C1(n11058), .C2(n11057), .A(n15730), .B(n11487), .ZN(
        n11059) );
  NAND2_X1 U13017 ( .A1(n12431), .A2(n11059), .ZN(n11060) );
  AOI21_X1 U13018 ( .B1(n15732), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n11060), 
        .ZN(n11061) );
  OAI211_X1 U13019 ( .C1(n12771), .C2(n11488), .A(n11062), .B(n11061), .ZN(
        P1_U3257) );
  INV_X1 U13020 ( .A(n11363), .ZN(n11063) );
  NAND2_X1 U13021 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n15536) );
  OAI21_X1 U13022 ( .B1(n14030), .B2(n11063), .A(n15536), .ZN(n11066) );
  OAI22_X1 U13023 ( .A1(n14044), .A2(n11367), .B1(n14031), .B2(n11064), .ZN(
        n11065) );
  AOI211_X1 U13024 ( .C1(n13142), .C2(n14077), .A(n11066), .B(n11065), .ZN(
        n11072) );
  AOI22_X1 U13025 ( .A1(n13994), .A2(n14079), .B1(n14054), .B2(n11067), .ZN(
        n11070) );
  OR3_X1 U13026 ( .A1(n11070), .A2(n11069), .A3(n11068), .ZN(n11071) );
  OAI211_X1 U13027 ( .C1(n10844), .C2(n11073), .A(n11072), .B(n11071), .ZN(
        P2_U3199) );
  OAI22_X1 U13028 ( .A1(n13126), .A2(n11177), .B1(n14002), .B2(n11074), .ZN(
        n11080) );
  AOI22_X1 U13029 ( .A1(n13994), .A2(n9000), .B1(n14054), .B2(n11075), .ZN(
        n11078) );
  INV_X1 U13030 ( .A(n13135), .ZN(n11077) );
  NOR3_X1 U13031 ( .A1(n11078), .A2(n11077), .A3(n11076), .ZN(n11079) );
  AOI211_X1 U13032 ( .C1(n11081), .C2(n14035), .A(n11080), .B(n11079), .ZN(
        n11082) );
  OAI21_X1 U13033 ( .B1(n11083), .B2(n10844), .A(n11082), .ZN(P2_U3209) );
  OAI21_X1 U13034 ( .B1(n11086), .B2(n11085), .A(n11084), .ZN(n11087) );
  NAND3_X1 U13035 ( .A1(n7454), .A2(n13241), .A3(n11087), .ZN(n11091) );
  OAI22_X1 U13036 ( .A1(n13255), .A2(n15782), .B1(n12909), .B2(n13247), .ZN(
        n11088) );
  AOI211_X1 U13037 ( .C1(n13245), .C2(n13484), .A(n11089), .B(n11088), .ZN(
        n11090) );
  OAI211_X1 U13038 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n13200), .A(n11091), .B(
        n11090), .ZN(P3_U3158) );
  NOR3_X1 U13039 ( .A1(n14038), .A2(n11093), .A3(n11092), .ZN(n11094) );
  AOI21_X1 U13040 ( .B1(n14054), .B2(n11095), .A(n11094), .ZN(n11105) );
  NAND2_X1 U13041 ( .A1(n14075), .A2(n14355), .ZN(n11097) );
  NAND2_X1 U13042 ( .A1(n14077), .A2(n14353), .ZN(n11096) );
  NAND2_X1 U13043 ( .A1(n11097), .A2(n11096), .ZN(n11195) );
  INV_X1 U13044 ( .A(n11195), .ZN(n11099) );
  NAND2_X1 U13045 ( .A1(n14046), .A2(n11198), .ZN(n11098) );
  NAND2_X1 U13046 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15558) );
  OAI211_X1 U13047 ( .C1(n14002), .C2(n11099), .A(n11098), .B(n15558), .ZN(
        n11102) );
  NOR2_X1 U13048 ( .A1(n11100), .A2(n10844), .ZN(n11101) );
  AOI211_X1 U13049 ( .C1(n15840), .C2(n14035), .A(n11102), .B(n11101), .ZN(
        n11103) );
  OAI21_X1 U13050 ( .B1(n11105), .B2(n11104), .A(n11103), .ZN(P2_U3185) );
  XOR2_X1 U13051 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11529), .Z(n11108) );
  AOI21_X1 U13052 ( .B1(n11110), .B2(P2_REG2_REG_8__SCAN_IN), .A(n11106), .ZN(
        n11107) );
  NAND2_X1 U13053 ( .A1(n11107), .A2(n11108), .ZN(n11520) );
  OAI21_X1 U13054 ( .B1(n11108), .B2(n11107), .A(n11520), .ZN(n11119) );
  INV_X1 U13055 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11111) );
  MUX2_X1 U13056 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n11111), .S(n11529), .Z(
        n11112) );
  OAI21_X1 U13057 ( .B1(n11113), .B2(n11112), .A(n11528), .ZN(n11114) );
  NAND2_X1 U13058 ( .A1(n11114), .A2(n15581), .ZN(n11116) );
  AND2_X1 U13059 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n12849) );
  AOI21_X1 U13060 ( .B1(n15522), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n12849), .ZN(
        n11115) );
  OAI211_X1 U13061 ( .C1(n14148), .C2(n11117), .A(n11116), .B(n11115), .ZN(
        n11118) );
  AOI21_X1 U13062 ( .B1(n15583), .B2(n11119), .A(n11118), .ZN(n11120) );
  INV_X1 U13063 ( .A(n11120), .ZN(P2_U3223) );
  INV_X1 U13064 ( .A(n12174), .ZN(n11125) );
  NOR2_X1 U13065 ( .A1(n11122), .A2(n11121), .ZN(n11228) );
  OR2_X1 U13066 ( .A1(n11228), .A2(n11229), .ZN(n11123) );
  XNOR2_X1 U13067 ( .A(n11123), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12175) );
  INV_X1 U13068 ( .A(n12175), .ZN(n12074) );
  OAI222_X1 U13069 ( .A1(n15476), .A2(n11124), .B1(n13160), .B2(n11125), .C1(
        P1_U3086), .C2(n12074), .ZN(P1_U3340) );
  OAI222_X1 U13070 ( .A1(n13150), .A2(n11126), .B1(n14477), .B2(n11125), .C1(
        P2_U3088), .C2(n14097), .ZN(P2_U3312) );
  XNOR2_X1 U13071 ( .A(n15813), .B(n15049), .ZN(n14953) );
  OR2_X1 U13072 ( .A1(n15050), .A2(n14787), .ZN(n11127) );
  XOR2_X1 U13073 ( .A(n14953), .B(n11565), .Z(n15816) );
  INV_X1 U13074 ( .A(n15816), .ZN(n11138) );
  NAND2_X1 U13075 ( .A1(n15050), .A2(n11129), .ZN(n11130) );
  OAI211_X1 U13076 ( .C1(n11132), .C2(n14953), .A(n11568), .B(n15988), .ZN(
        n11133) );
  INV_X1 U13077 ( .A(n11133), .ZN(n11134) );
  AOI211_X1 U13078 ( .C1(n15816), .C2(n15880), .A(n11135), .B(n11134), .ZN(
        n15819) );
  AOI211_X1 U13079 ( .C1(n15813), .C2(n11136), .A(n15354), .B(n11572), .ZN(
        n15814) );
  AOI21_X1 U13080 ( .B1(n15981), .B2(n15813), .A(n15814), .ZN(n11137) );
  OAI211_X1 U13081 ( .C1(n15875), .C2(n11138), .A(n15819), .B(n11137), .ZN(
        n11141) );
  NAND2_X1 U13082 ( .A1(n11141), .A2(n15991), .ZN(n11139) );
  OAI21_X1 U13083 ( .B1(n15991), .B2(n11140), .A(n11139), .ZN(P1_U3534) );
  INV_X1 U13084 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11143) );
  NAND2_X1 U13085 ( .A1(n11141), .A2(n15994), .ZN(n11142) );
  OAI21_X1 U13086 ( .B1(n15994), .B2(n11143), .A(n11142), .ZN(P1_U3477) );
  INV_X1 U13087 ( .A(n11144), .ZN(n11145) );
  OAI222_X1 U13088 ( .A1(n11146), .A2(P3_U3151), .B1(n13983), .B2(n13381), 
        .C1(n13157), .C2(n11145), .ZN(P3_U3275) );
  NOR2_X1 U13089 ( .A1(n11147), .A2(n13057), .ZN(n11148) );
  NOR2_X1 U13090 ( .A1(n12900), .A2(n11148), .ZN(n11153) );
  INV_X1 U13091 ( .A(n15769), .ZN(n13880) );
  AOI22_X1 U13092 ( .A1(n13759), .A2(n13487), .B1(n13485), .B2(n13742), .ZN(
        n11152) );
  XNOR2_X1 U13093 ( .A(n12897), .B(n11149), .ZN(n11150) );
  NAND2_X1 U13094 ( .A1(n11150), .A2(n13756), .ZN(n11151) );
  OAI211_X1 U13095 ( .C1(n11153), .C2(n13880), .A(n11152), .B(n11151), .ZN(
        n11678) );
  INV_X1 U13096 ( .A(n11678), .ZN(n11156) );
  INV_X1 U13097 ( .A(n11153), .ZN(n11682) );
  NAND2_X1 U13098 ( .A1(n15997), .A2(n15889), .ZN(n13885) );
  INV_X1 U13099 ( .A(n13885), .ZN(n12153) );
  OAI22_X1 U13100 ( .A1(n13905), .A2(n11208), .B1(n15997), .B2(n8290), .ZN(
        n11154) );
  AOI21_X1 U13101 ( .B1(n11682), .B2(n12153), .A(n11154), .ZN(n11155) );
  OAI21_X1 U13102 ( .B1(n11156), .B2(n16004), .A(n11155), .ZN(P3_U3461) );
  INV_X1 U13103 ( .A(n11157), .ZN(n11158) );
  AOI211_X1 U13104 ( .C1(n11160), .C2(n11159), .A(n15135), .B(n11158), .ZN(
        n11169) );
  INV_X1 U13105 ( .A(n11161), .ZN(n11162) );
  AOI211_X1 U13106 ( .C1(n11164), .C2(n11163), .A(n15087), .B(n11162), .ZN(
        n11168) );
  NAND2_X1 U13107 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12236)
         );
  NAND2_X1 U13108 ( .A1(n15732), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n11165) );
  OAI211_X1 U13109 ( .C1(n12771), .C2(n11166), .A(n12236), .B(n11165), .ZN(
        n11167) );
  OR3_X1 U13110 ( .A1(n11169), .A2(n11168), .A3(n11167), .ZN(P1_U3256) );
  NAND3_X1 U13111 ( .A1(n15525), .A2(n15526), .A3(n11170), .ZN(n11171) );
  NOR2_X1 U13112 ( .A1(n11173), .A2(n9722), .ZN(n11174) );
  NAND2_X1 U13113 ( .A1(n14311), .A2(n14305), .ZN(n11175) );
  NOR2_X1 U13114 ( .A1(n11185), .A2(n14140), .ZN(n14314) );
  OAI22_X1 U13115 ( .A1(n14311), .A2(n10219), .B1(n11177), .B2(n14308), .ZN(
        n11178) );
  AOI21_X1 U13116 ( .B1(n14314), .B2(n11179), .A(n11178), .ZN(n11180) );
  OAI21_X1 U13117 ( .B1(n9019), .B2(n14349), .A(n11180), .ZN(n11181) );
  AOI21_X1 U13118 ( .B1(n14292), .B2(n11182), .A(n11181), .ZN(n11183) );
  OAI21_X1 U13119 ( .B1(n14359), .B2(n11184), .A(n11183), .ZN(P2_U3263) );
  INV_X1 U13120 ( .A(n14231), .ZN(n14335) );
  NOR2_X2 U13121 ( .A1(n11185), .A2(n12832), .ZN(n14362) );
  OAI22_X1 U13122 ( .A1(n14311), .A2(n10220), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14308), .ZN(n11186) );
  AOI21_X1 U13123 ( .B1(n14362), .B2(n11187), .A(n11186), .ZN(n11188) );
  OAI21_X1 U13124 ( .B1(n11189), .B2(n14349), .A(n11188), .ZN(n11190) );
  AOI21_X1 U13125 ( .B1(n14335), .B2(n11191), .A(n11190), .ZN(n11192) );
  OAI21_X1 U13126 ( .B1(n14359), .B2(n11193), .A(n11192), .ZN(P2_U3262) );
  XNOR2_X1 U13127 ( .A(n11194), .B(n11202), .ZN(n11196) );
  AOI21_X1 U13128 ( .B1(n11196), .B2(n14358), .A(n11195), .ZN(n15843) );
  INV_X1 U13129 ( .A(n11457), .ZN(n11197) );
  AOI211_X1 U13130 ( .C1(n15840), .C2(n11197), .A(n15821), .B(n11383), .ZN(
        n15839) );
  AOI22_X1 U13131 ( .A1(n14359), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n11198), 
        .B2(n14345), .ZN(n11199) );
  OAI21_X1 U13132 ( .B1(n11200), .B2(n14349), .A(n11199), .ZN(n11201) );
  AOI21_X1 U13133 ( .B1(n15839), .B2(n14314), .A(n11201), .ZN(n11205) );
  NAND2_X1 U13134 ( .A1(n11203), .A2(n11202), .ZN(n15837) );
  NAND3_X1 U13135 ( .A1(n15838), .A2(n15837), .A3(n14292), .ZN(n11204) );
  OAI211_X1 U13136 ( .C1(n15843), .C2(n14359), .A(n11205), .B(n11204), .ZN(
        P2_U3258) );
  NAND2_X1 U13137 ( .A1(n11678), .A2(n16000), .ZN(n11207) );
  NAND2_X1 U13138 ( .A1(n16000), .A2(n15889), .ZN(n13946) );
  INV_X1 U13139 ( .A(n13946), .ZN(n15771) );
  AOI22_X1 U13140 ( .A1(n11682), .A2(n15771), .B1(P3_REG0_REG_2__SCAN_IN), 
        .B2(n16008), .ZN(n11206) );
  OAI211_X1 U13141 ( .C1(n13960), .C2(n11208), .A(n11207), .B(n11206), .ZN(
        P3_U3396) );
  MUX2_X1 U13142 ( .A(n10218), .B(n11209), .S(n14311), .Z(n11215) );
  INV_X1 U13143 ( .A(n14362), .ZN(n14163) );
  INV_X1 U13144 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11210) );
  OAI22_X1 U13145 ( .A1(n14163), .A2(n11211), .B1(n11210), .B2(n14308), .ZN(
        n11212) );
  AOI21_X1 U13146 ( .B1(n14271), .B2(n11213), .A(n11212), .ZN(n11214) );
  OAI211_X1 U13147 ( .C1(n11216), .C2(n14231), .A(n11215), .B(n11214), .ZN(
        P2_U3264) );
  NOR2_X1 U13148 ( .A1(n11217), .A2(n15912), .ZN(n15765) );
  XNOR2_X1 U13149 ( .A(n8679), .B(n11218), .ZN(n11219) );
  OAI222_X1 U13150 ( .A1(n13835), .A2(n12909), .B1(n13833), .B2(n12896), .C1(
        n13831), .C2(n11219), .ZN(n15766) );
  AOI21_X1 U13151 ( .B1(n15765), .B2(n13084), .A(n15766), .ZN(n11220) );
  MUX2_X1 U13152 ( .A(n11221), .B(n11220), .S(n15810), .Z(n11225) );
  AND2_X1 U13153 ( .A1(n11222), .A2(n8747), .ZN(n11681) );
  OR2_X1 U13154 ( .A1(n15769), .A2(n11681), .ZN(n15800) );
  OAI21_X1 U13155 ( .B1(n8679), .B2(n8148), .A(n11223), .ZN(n15770) );
  AOI22_X1 U13156 ( .A1(n13820), .A2(n15770), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n13802), .ZN(n11224) );
  NAND2_X1 U13157 ( .A1(n11225), .A2(n11224), .ZN(P3_U3232) );
  INV_X1 U13158 ( .A(n12204), .ZN(n11235) );
  INV_X1 U13159 ( .A(n14127), .ZN(n14117) );
  OAI222_X1 U13160 ( .A1(n13150), .A2(n11226), .B1(n14477), .B2(n11235), .C1(
        n14117), .C2(P2_U3088), .ZN(P2_U3311) );
  AND2_X1 U13161 ( .A1(n11228), .A2(n11227), .ZN(n11232) );
  NOR2_X1 U13162 ( .A1(n11232), .A2(n11229), .ZN(n11230) );
  MUX2_X1 U13163 ( .A(n11229), .B(n11230), .S(P1_IR_REG_16__SCAN_IN), .Z(
        n11234) );
  NAND2_X1 U13164 ( .A1(n11232), .A2(n11231), .ZN(n11408) );
  INV_X1 U13165 ( .A(n11408), .ZN(n11233) );
  NOR2_X1 U13166 ( .A1(n11234), .A2(n11233), .ZN(n12205) );
  INV_X1 U13167 ( .A(n12205), .ZN(n12755) );
  OAI222_X1 U13168 ( .A1(n15476), .A2(n11236), .B1(n13160), .B2(n11235), .C1(
        n12755), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI21_X1 U13169 ( .B1(n11239), .B2(n11238), .A(n11237), .ZN(n11240) );
  NAND2_X1 U13170 ( .A1(n11240), .A2(n13241), .ZN(n11245) );
  INV_X1 U13171 ( .A(n13485), .ZN(n11241) );
  OAI22_X1 U13172 ( .A1(n13255), .A2(n11436), .B1(n11241), .B2(n13247), .ZN(
        n11242) );
  AOI211_X1 U13173 ( .C1(n13245), .C2(n13483), .A(n11243), .B(n11242), .ZN(
        n11244) );
  OAI211_X1 U13174 ( .C1(n11435), .C2(n13200), .A(n11245), .B(n11244), .ZN(
        P3_U3170) );
  OAI21_X1 U13175 ( .B1(n11248), .B2(n11247), .A(n11246), .ZN(n11439) );
  OAI211_X1 U13176 ( .C1(n11250), .C2(n13053), .A(n11249), .B(n13756), .ZN(
        n11252) );
  AOI22_X1 U13177 ( .A1(n13483), .A2(n13742), .B1(n13759), .B2(n13485), .ZN(
        n11251) );
  NAND2_X1 U13178 ( .A1(n11252), .A2(n11251), .ZN(n11434) );
  AOI21_X1 U13179 ( .B1(n15917), .B2(n11439), .A(n11434), .ZN(n11257) );
  OAI22_X1 U13180 ( .A1(n13960), .A2(n11436), .B1(n16000), .B2(n8321), .ZN(
        n11253) );
  INV_X1 U13181 ( .A(n11253), .ZN(n11254) );
  OAI21_X1 U13182 ( .B1(n11257), .B2(n16008), .A(n11254), .ZN(P3_U3402) );
  AOI22_X1 U13183 ( .A1(n16005), .A2(n11255), .B1(n16004), .B2(
        P3_REG1_REG_4__SCAN_IN), .ZN(n11256) );
  OAI21_X1 U13184 ( .B1(n11257), .B2(n16004), .A(n11256), .ZN(P3_U3463) );
  NAND4_X1 U13185 ( .A1(n11261), .A2(n11260), .A3(n11259), .A4(n11258), .ZN(
        n15165) );
  INV_X1 U13186 ( .A(n11262), .ZN(n11273) );
  INV_X2 U13187 ( .A(n15946), .ZN(n15760) );
  AND2_X1 U13188 ( .A1(n11263), .A2(n8111), .ZN(n11264) );
  OAI22_X1 U13189 ( .A1(n15760), .A2(n10181), .B1(n11265), .B2(n15755), .ZN(
        n11270) );
  INV_X1 U13190 ( .A(n11266), .ZN(n11268) );
  OR2_X1 U13191 ( .A1(n14758), .A2(n10342), .ZN(n14938) );
  INV_X1 U13192 ( .A(n14938), .ZN(n15759) );
  NAND2_X1 U13193 ( .A1(n15760), .A2(n15759), .ZN(n15363) );
  OAI22_X1 U13194 ( .A1(n11268), .A2(n15363), .B1(n15358), .B2(n11267), .ZN(
        n11269) );
  AOI211_X1 U13195 ( .C1(n15947), .C2(n11271), .A(n11270), .B(n11269), .ZN(
        n11272) );
  OAI21_X1 U13196 ( .B1(n15946), .B2(n11273), .A(n11272), .ZN(P1_U3292) );
  NAND2_X1 U13197 ( .A1(n11274), .A2(n14944), .ZN(n11277) );
  AOI22_X1 U13198 ( .A1(n12597), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12596), 
        .B2(n11275), .ZN(n11276) );
  INV_X1 U13199 ( .A(n15848), .ZN(n11662) );
  NAND2_X1 U13200 ( .A1(n14924), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11284) );
  OR2_X1 U13201 ( .A1(n14928), .A2(n15853), .ZN(n11283) );
  NAND2_X1 U13202 ( .A1(n11279), .A2(n11278), .ZN(n11280) );
  NAND2_X1 U13203 ( .A1(n11307), .A2(n11280), .ZN(n11661) );
  OR2_X1 U13204 ( .A1(n7189), .A2(n11661), .ZN(n11282) );
  OR2_X1 U13205 ( .A1(n12705), .A2(n10383), .ZN(n11281) );
  NAND4_X1 U13206 ( .A1(n11284), .A2(n11283), .A3(n11282), .A4(n11281), .ZN(
        n15047) );
  INV_X1 U13207 ( .A(n15047), .ZN(n11620) );
  OAI22_X1 U13208 ( .A1(n11662), .A2(n14627), .B1(n11620), .B2(n14572), .ZN(
        n11285) );
  XNOR2_X1 U13209 ( .A(n11285), .B(n14628), .ZN(n11638) );
  OAI22_X1 U13210 ( .A1(n11662), .A2(n14572), .B1(n11620), .B2(n14626), .ZN(
        n11637) );
  XNOR2_X1 U13211 ( .A(n11638), .B(n11637), .ZN(n11304) );
  NAND2_X1 U13212 ( .A1(n11292), .A2(n14944), .ZN(n11295) );
  AOI22_X1 U13213 ( .A1(n12597), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7182), 
        .B2(n11293), .ZN(n11294) );
  INV_X1 U13214 ( .A(n14796), .ZN(n15830) );
  OAI22_X1 U13215 ( .A1(n15830), .A2(n14627), .B1(n11617), .B2(n14572), .ZN(
        n11296) );
  XNOR2_X1 U13216 ( .A(n11296), .B(n14628), .ZN(n11300) );
  NAND2_X1 U13217 ( .A1(n14796), .A2(n14587), .ZN(n11298) );
  OR2_X1 U13218 ( .A1(n11617), .A2(n14626), .ZN(n11297) );
  NAND2_X1 U13219 ( .A1(n11298), .A2(n11297), .ZN(n11299) );
  INV_X1 U13220 ( .A(n11299), .ZN(n11302) );
  INV_X1 U13221 ( .A(n11300), .ZN(n11301) );
  AOI21_X1 U13222 ( .B1(n11304), .B2(n11303), .A(n7344), .ZN(n11316) );
  OAI21_X1 U13223 ( .B1(n14743), .B2(n11617), .A(n11305), .ZN(n11314) );
  NAND2_X1 U13224 ( .A1(n14924), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11312) );
  OR2_X1 U13225 ( .A1(n14928), .A2(n15881), .ZN(n11311) );
  AND2_X1 U13226 ( .A1(n11307), .A2(n11306), .ZN(n11308) );
  OR2_X1 U13227 ( .A1(n11308), .A2(n11592), .ZN(n11723) );
  OR2_X1 U13228 ( .A1(n7189), .A2(n11723), .ZN(n11310) );
  OR2_X1 U13229 ( .A1(n12705), .A2(n10403), .ZN(n11309) );
  NAND4_X1 U13230 ( .A1(n11312), .A2(n11311), .A3(n11310), .A4(n11309), .ZN(
        n15046) );
  INV_X1 U13231 ( .A(n15046), .ZN(n11821) );
  OAI22_X1 U13232 ( .A1(n11821), .A2(n14747), .B1(n14746), .B2(n11661), .ZN(
        n11313) );
  AOI211_X1 U13233 ( .C1(n14751), .C2(n15848), .A(n11314), .B(n11313), .ZN(
        n11315) );
  OAI21_X1 U13234 ( .B1(n11316), .B2(n14753), .A(n11315), .ZN(P1_U3221) );
  INV_X1 U13235 ( .A(n11317), .ZN(n11318) );
  OAI222_X1 U13236 ( .A1(n12898), .A2(P3_U3151), .B1(n13983), .B2(n13398), 
        .C1(n13157), .C2(n11318), .ZN(P3_U3274) );
  OAI21_X1 U13237 ( .B1(n11320), .B2(n14951), .A(n11319), .ZN(n15778) );
  INV_X1 U13238 ( .A(n15778), .ZN(n11338) );
  NOR3_X1 U13239 ( .A1(n11322), .A2(n14767), .A3(n11321), .ZN(n11325) );
  INV_X1 U13240 ( .A(n11323), .ZN(n11324) );
  OAI21_X1 U13241 ( .B1(n11325), .B2(n11324), .A(n15988), .ZN(n11327) );
  AOI22_X1 U13242 ( .A1(n15342), .A2(n15052), .B1(n15054), .B2(n15289), .ZN(
        n11326) );
  OAI211_X1 U13243 ( .C1(n11338), .C2(n11328), .A(n11327), .B(n11326), .ZN(
        n15776) );
  NAND2_X1 U13244 ( .A1(n15776), .A2(n15760), .ZN(n11337) );
  OAI22_X1 U13245 ( .A1(n15760), .A2(n11330), .B1(n11329), .B2(n15755), .ZN(
        n11335) );
  AOI21_X1 U13246 ( .B1(n11331), .B2(n14769), .A(n15354), .ZN(n11333) );
  NAND2_X1 U13247 ( .A1(n11333), .A2(n11332), .ZN(n15774) );
  NOR2_X1 U13248 ( .A1(n15358), .A2(n15774), .ZN(n11334) );
  AOI211_X1 U13249 ( .C1(n15947), .C2(n14769), .A(n11335), .B(n11334), .ZN(
        n11336) );
  OAI211_X1 U13250 ( .C1(n11338), .C2(n15363), .A(n11337), .B(n11336), .ZN(
        P1_U3291) );
  XOR2_X1 U13251 ( .A(n11339), .B(n11342), .Z(n11346) );
  AND2_X1 U13252 ( .A1(n11341), .A2(n11340), .ZN(n11343) );
  AOI22_X1 U13253 ( .A1(n14353), .A2(n14075), .B1(n14073), .B2(n14355), .ZN(
        n11344) );
  OAI21_X1 U13254 ( .B1(n11375), .B2(n10019), .A(n11344), .ZN(n11345) );
  AOI21_X1 U13255 ( .B1(n11346), .B2(n14358), .A(n11345), .ZN(n11374) );
  AOI211_X1 U13256 ( .C1(n12854), .C2(n11382), .A(n15821), .B(n7584), .ZN(
        n11372) );
  INV_X1 U13257 ( .A(n12854), .ZN(n11348) );
  AOI22_X1 U13258 ( .A1(n14347), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n12850), 
        .B2(n14345), .ZN(n11347) );
  OAI21_X1 U13259 ( .B1(n11348), .B2(n14349), .A(n11347), .ZN(n11350) );
  NOR2_X1 U13260 ( .A1(n11375), .A2(n14231), .ZN(n11349) );
  AOI211_X1 U13261 ( .C1(n11372), .C2(n14314), .A(n11350), .B(n11349), .ZN(
        n11351) );
  OAI21_X1 U13262 ( .B1(n14347), .B2(n11374), .A(n11351), .ZN(P2_U3256) );
  XNOR2_X1 U13263 ( .A(n11352), .B(n11353), .ZN(n15901) );
  XNOR2_X1 U13264 ( .A(n11354), .B(n11353), .ZN(n11356) );
  OAI22_X1 U13265 ( .A1(n12795), .A2(n14320), .B1(n12794), .B2(n14322), .ZN(
        n11355) );
  AOI21_X1 U13266 ( .B1(n11356), .B2(n14358), .A(n11355), .ZN(n11357) );
  OAI21_X1 U13267 ( .B1(n15901), .B2(n10019), .A(n11357), .ZN(n15905) );
  NAND2_X1 U13268 ( .A1(n15905), .A2(n14311), .ZN(n11362) );
  OAI211_X1 U13269 ( .C1(n15904), .C2(n7584), .A(n14445), .B(n11509), .ZN(
        n15902) );
  INV_X1 U13270 ( .A(n15902), .ZN(n11360) );
  AOI22_X1 U13271 ( .A1(n14359), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12793), 
        .B2(n14345), .ZN(n11358) );
  OAI21_X1 U13272 ( .B1(n15904), .B2(n14349), .A(n11358), .ZN(n11359) );
  AOI21_X1 U13273 ( .B1(n11360), .B2(n14314), .A(n11359), .ZN(n11361) );
  OAI211_X1 U13274 ( .C1(n15901), .C2(n14231), .A(n11362), .B(n11361), .ZN(
        P2_U3255) );
  AOI22_X1 U13275 ( .A1(n14347), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n11363), 
        .B2(n14345), .ZN(n11366) );
  NAND2_X1 U13276 ( .A1(n14362), .A2(n11364), .ZN(n11365) );
  OAI211_X1 U13277 ( .C1(n11367), .C2(n14349), .A(n11366), .B(n11365), .ZN(
        n11368) );
  AOI21_X1 U13278 ( .B1(n11369), .B2(n14335), .A(n11368), .ZN(n11370) );
  OAI21_X1 U13279 ( .B1(n11371), .B2(n14359), .A(n11370), .ZN(P2_U3260) );
  AOI21_X1 U13280 ( .B1(n15841), .B2(n12854), .A(n11372), .ZN(n11373) );
  OAI211_X1 U13281 ( .C1(n14449), .C2(n11375), .A(n11374), .B(n11373), .ZN(
        n11396) );
  NAND2_X1 U13282 ( .A1(n11396), .A2(n14451), .ZN(n11376) );
  OAI21_X1 U13283 ( .B1(n14451), .B2(n11111), .A(n11376), .ZN(P2_U3508) );
  XNOR2_X1 U13284 ( .A(n11377), .B(n11386), .ZN(n11378) );
  NAND2_X1 U13285 ( .A1(n11378), .A2(n14358), .ZN(n11380) );
  NAND2_X1 U13286 ( .A1(n11380), .A2(n11379), .ZN(n15858) );
  AOI21_X1 U13287 ( .B1(n11381), .B2(n14345), .A(n15858), .ZN(n11395) );
  INV_X1 U13288 ( .A(n14314), .ZN(n11392) );
  OAI211_X1 U13289 ( .C1(n11383), .C2(n15857), .A(n14445), .B(n11382), .ZN(
        n15856) );
  NAND2_X1 U13290 ( .A1(n15838), .A2(n11384), .ZN(n11387) );
  NAND2_X1 U13291 ( .A1(n11387), .A2(n11386), .ZN(n11385) );
  OAI21_X1 U13292 ( .B1(n11387), .B2(n11386), .A(n11385), .ZN(n11388) );
  INV_X1 U13293 ( .A(n11388), .ZN(n15861) );
  NAND2_X1 U13294 ( .A1(n15861), .A2(n14292), .ZN(n11391) );
  AOI22_X1 U13295 ( .A1(n14271), .A2(n11389), .B1(n14347), .B2(
        P2_REG2_REG_8__SCAN_IN), .ZN(n11390) );
  OAI211_X1 U13296 ( .C1(n11392), .C2(n15856), .A(n11391), .B(n11390), .ZN(
        n11393) );
  INV_X1 U13297 ( .A(n11393), .ZN(n11394) );
  OAI21_X1 U13298 ( .B1(n14359), .B2(n11395), .A(n11394), .ZN(P2_U3257) );
  INV_X1 U13299 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11398) );
  NAND2_X1 U13300 ( .A1(n11396), .A2(n14469), .ZN(n11397) );
  OAI21_X1 U13301 ( .B1(n14469), .B2(n11398), .A(n11397), .ZN(P2_U3457) );
  INV_X1 U13302 ( .A(n11399), .ZN(n11401) );
  INV_X1 U13303 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11400) );
  OAI22_X1 U13304 ( .A1(n14347), .A2(n11401), .B1(n11400), .B2(n14308), .ZN(
        n11402) );
  AOI21_X1 U13305 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n14347), .A(n11402), .ZN(
        n11405) );
  OAI21_X1 U13306 ( .B1(n14271), .B2(n14362), .A(n11403), .ZN(n11404) );
  OAI211_X1 U13307 ( .C1(n14231), .C2(n11406), .A(n11405), .B(n11404), .ZN(
        P2_U3265) );
  INV_X1 U13308 ( .A(n12330), .ZN(n11410) );
  INV_X1 U13309 ( .A(n15567), .ZN(n14120) );
  OAI222_X1 U13310 ( .A1(n13150), .A2(n11407), .B1(n14477), .B2(n11410), .C1(
        n14120), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U13311 ( .A1(n11408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11409) );
  XNOR2_X1 U13312 ( .A(n11409), .B(P1_IR_REG_17__SCAN_IN), .ZN(n12757) );
  INV_X1 U13313 ( .A(n12757), .ZN(n12770) );
  OAI222_X1 U13314 ( .A1(n15476), .A2(n11411), .B1(n13160), .B2(n11410), .C1(
        n12770), .C2(P1_U3086), .ZN(P1_U3338) );
  OR2_X1 U13315 ( .A1(n11564), .A2(n15345), .ZN(n11413) );
  NAND2_X1 U13316 ( .A1(n15047), .A2(n15342), .ZN(n11412) );
  NAND2_X1 U13317 ( .A1(n11413), .A2(n11412), .ZN(n11569) );
  NAND2_X1 U13318 ( .A1(n11569), .A2(n14694), .ZN(n11415) );
  OAI211_X1 U13319 ( .C1(n14746), .C2(n11573), .A(n11415), .B(n11414), .ZN(
        n11420) );
  XNOR2_X1 U13320 ( .A(n11417), .B(n11416), .ZN(n11418) );
  NOR2_X1 U13321 ( .A1(n11418), .A2(n14753), .ZN(n11419) );
  AOI211_X1 U13322 ( .C1(n14751), .C2(n14796), .A(n11420), .B(n11419), .ZN(
        n11421) );
  INV_X1 U13323 ( .A(n11421), .ZN(P1_U3213) );
  NOR2_X1 U13324 ( .A1(n13969), .A2(SI_22_), .ZN(n11422) );
  AOI21_X1 U13325 ( .B1(n12899), .B2(P3_STATE_REG_SCAN_IN), .A(n11422), .ZN(
        n11423) );
  OAI21_X1 U13326 ( .B1(n11424), .B2(n13157), .A(n11423), .ZN(n11425) );
  INV_X1 U13327 ( .A(n11425), .ZN(P3_U3273) );
  OAI21_X1 U13328 ( .B1(n11428), .B2(n11427), .A(n11426), .ZN(n11429) );
  NAND2_X1 U13329 ( .A1(n11429), .A2(n13241), .ZN(n11433) );
  OAI22_X1 U13330 ( .A1(n13255), .A2(n11941), .B1(n11497), .B2(n13247), .ZN(
        n11430) );
  AOI211_X1 U13331 ( .C1(n13245), .C2(n13482), .A(n11431), .B(n11430), .ZN(
        n11432) );
  OAI211_X1 U13332 ( .C1(n11940), .C2(n13200), .A(n11433), .B(n11432), .ZN(
        P3_U3167) );
  INV_X1 U13333 ( .A(n11434), .ZN(n11441) );
  NOR2_X1 U13334 ( .A1(n15810), .A2(n10583), .ZN(n11438) );
  OAI22_X1 U13335 ( .A1(n15806), .A2(n11436), .B1(n11435), .B2(n15804), .ZN(
        n11437) );
  AOI211_X1 U13336 ( .C1(n11439), .C2(n13820), .A(n11438), .B(n11437), .ZN(
        n11440) );
  OAI21_X1 U13337 ( .B1(n15802), .B2(n11441), .A(n11440), .ZN(P3_U3229) );
  NAND2_X1 U13338 ( .A1(n11442), .A2(n13052), .ZN(n11443) );
  NAND3_X1 U13339 ( .A1(n11444), .A2(n13756), .A3(n11443), .ZN(n11446) );
  AOI22_X1 U13340 ( .A1(n13484), .A2(n13742), .B1(n13759), .B2(n13486), .ZN(
        n11445) );
  NAND2_X1 U13341 ( .A1(n11446), .A2(n11445), .ZN(n15783) );
  INV_X1 U13342 ( .A(n15783), .ZN(n11453) );
  OAI21_X1 U13343 ( .B1(n11448), .B2(n13052), .A(n11447), .ZN(n15785) );
  AOI22_X1 U13344 ( .A1(n13816), .A2(n11449), .B1(n13802), .B2(n13333), .ZN(
        n11450) );
  OAI21_X1 U13345 ( .B1(n8307), .B2(n15810), .A(n11450), .ZN(n11451) );
  AOI21_X1 U13346 ( .B1(n13820), .B2(n15785), .A(n11451), .ZN(n11452) );
  OAI21_X1 U13347 ( .B1(n15802), .B2(n11453), .A(n11452), .ZN(P3_U3230) );
  XNOR2_X1 U13348 ( .A(n11454), .B(n11463), .ZN(n15825) );
  AND2_X1 U13349 ( .A1(n11456), .A2(n11455), .ZN(n11458) );
  OR2_X1 U13350 ( .A1(n11458), .A2(n11457), .ZN(n15822) );
  INV_X1 U13351 ( .A(n15822), .ZN(n11459) );
  NAND2_X1 U13352 ( .A1(n14362), .A2(n11459), .ZN(n11462) );
  NAND2_X1 U13353 ( .A1(n14345), .A2(n11460), .ZN(n11461) );
  OAI211_X1 U13354 ( .C1(n14349), .C2(n15820), .A(n11462), .B(n11461), .ZN(
        n11471) );
  NAND2_X1 U13355 ( .A1(n11464), .A2(n11463), .ZN(n11465) );
  NAND2_X1 U13356 ( .A1(n11466), .A2(n11465), .ZN(n11467) );
  NAND2_X1 U13357 ( .A1(n11467), .A2(n14358), .ZN(n11469) );
  AOI22_X1 U13358 ( .A1(n14355), .A2(n14076), .B1(n14078), .B2(n14353), .ZN(
        n11468) );
  NAND2_X1 U13359 ( .A1(n11469), .A2(n11468), .ZN(n15823) );
  MUX2_X1 U13360 ( .A(n15823), .B(P2_REG2_REG_6__SCAN_IN), .S(n14359), .Z(
        n11470) );
  AOI211_X1 U13361 ( .C1(n14292), .C2(n15825), .A(n11471), .B(n11470), .ZN(
        n11472) );
  INV_X1 U13362 ( .A(n11472), .ZN(P2_U3259) );
  NAND2_X1 U13363 ( .A1(n14345), .A2(n11473), .ZN(n11476) );
  NAND2_X1 U13364 ( .A1(n14271), .A2(n11474), .ZN(n11475) );
  OAI211_X1 U13365 ( .C1(n14163), .C2(n11477), .A(n11476), .B(n11475), .ZN(
        n11480) );
  MUX2_X1 U13366 ( .A(n11478), .B(P2_REG2_REG_4__SCAN_IN), .S(n14359), .Z(
        n11479) );
  AOI211_X1 U13367 ( .C1(n14292), .C2(n11481), .A(n11480), .B(n11479), .ZN(
        n11482) );
  INV_X1 U13368 ( .A(n11482), .ZN(P2_U3261) );
  AOI21_X1 U13369 ( .B1(n12006), .B2(P1_REG1_REG_14__SCAN_IN), .A(n11483), 
        .ZN(n12075) );
  XNOR2_X1 U13370 ( .A(n12075), .B(n12074), .ZN(n11484) );
  NOR2_X1 U13371 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n11484), .ZN(n12073) );
  AOI21_X1 U13372 ( .B1(n11484), .B2(P1_REG1_REG_15__SCAN_IN), .A(n12073), 
        .ZN(n11493) );
  INV_X1 U13373 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n14741) );
  NOR2_X1 U13374 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14741), .ZN(n11486) );
  NOR2_X1 U13375 ( .A1(n12771), .A2(n12074), .ZN(n11485) );
  AOI211_X1 U13376 ( .C1(n15732), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n11486), 
        .B(n11485), .ZN(n11492) );
  OAI21_X1 U13377 ( .B1(n11989), .B2(n11488), .A(n11487), .ZN(n12066) );
  XNOR2_X1 U13378 ( .A(n12066), .B(n12175), .ZN(n11489) );
  NOR2_X1 U13379 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11489), .ZN(n12069) );
  AOI21_X1 U13380 ( .B1(n11489), .B2(P1_REG2_REG_15__SCAN_IN), .A(n12069), 
        .ZN(n11490) );
  OR2_X1 U13381 ( .A1(n11490), .A2(n15087), .ZN(n11491) );
  OAI211_X1 U13382 ( .C1(n11493), .C2(n15135), .A(n11492), .B(n11491), .ZN(
        P1_U3258) );
  NAND2_X1 U13383 ( .A1(n11494), .A2(n13055), .ZN(n11495) );
  NAND2_X1 U13384 ( .A1(n11496), .A2(n11495), .ZN(n11499) );
  OAI22_X1 U13385 ( .A1(n11935), .A2(n13835), .B1(n11497), .B2(n13833), .ZN(
        n11498) );
  AOI21_X1 U13386 ( .B1(n11499), .B2(n13756), .A(n11498), .ZN(n11504) );
  OR2_X1 U13387 ( .A1(n11500), .A2(n13055), .ZN(n11501) );
  NAND2_X1 U13388 ( .A1(n11502), .A2(n11501), .ZN(n11945) );
  NAND2_X1 U13389 ( .A1(n11945), .A2(n15769), .ZN(n11503) );
  NAND2_X1 U13390 ( .A1(n11504), .A2(n11503), .ZN(n11942) );
  INV_X1 U13391 ( .A(n11942), .ZN(n11809) );
  OAI22_X1 U13392 ( .A1(n13960), .A2(n11941), .B1(n16000), .B2(n8335), .ZN(
        n11505) );
  AOI21_X1 U13393 ( .B1(n11945), .B2(n15771), .A(n11505), .ZN(n11506) );
  OAI21_X1 U13394 ( .B1(n11809), .B2(n16008), .A(n11506), .ZN(P3_U3405) );
  XNOR2_X1 U13395 ( .A(n11508), .B(n11507), .ZN(n11632) );
  AOI211_X1 U13396 ( .C1(n11879), .C2(n11509), .A(n15821), .B(n11846), .ZN(
        n11629) );
  INV_X1 U13397 ( .A(n11879), .ZN(n11511) );
  AOI22_X1 U13398 ( .A1(n14359), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11870), 
        .B2(n14345), .ZN(n11510) );
  OAI21_X1 U13399 ( .B1(n11511), .B2(n14349), .A(n11510), .ZN(n11518) );
  XNOR2_X1 U13400 ( .A(n11513), .B(n11512), .ZN(n11516) );
  NAND2_X1 U13401 ( .A1(n14071), .A2(n14355), .ZN(n11515) );
  NAND2_X1 U13402 ( .A1(n14073), .A2(n14353), .ZN(n11514) );
  NAND2_X1 U13403 ( .A1(n11515), .A2(n11514), .ZN(n11871) );
  AOI21_X1 U13404 ( .B1(n11516), .B2(n14358), .A(n11871), .ZN(n11631) );
  NOR2_X1 U13405 ( .A1(n11631), .A2(n14347), .ZN(n11517) );
  AOI211_X1 U13406 ( .C1(n11629), .C2(n14314), .A(n11518), .B(n11517), .ZN(
        n11519) );
  OAI21_X1 U13407 ( .B1(n14364), .B2(n11632), .A(n11519), .ZN(P2_U3254) );
  OAI21_X1 U13408 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n11529), .A(n11520), .ZN(
        n15593) );
  XNOR2_X1 U13409 ( .A(n15597), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n15594) );
  NOR2_X1 U13410 ( .A1(n15593), .A2(n15594), .ZN(n15591) );
  INV_X1 U13411 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11521) );
  MUX2_X1 U13412 ( .A(n11521), .B(P2_REG2_REG_11__SCAN_IN), .S(n12100), .Z(
        n11522) );
  INV_X1 U13413 ( .A(n11522), .ZN(n11523) );
  NAND2_X1 U13414 ( .A1(n11524), .A2(n11523), .ZN(n12093) );
  OAI21_X1 U13415 ( .B1(n11524), .B2(n11523), .A(n12093), .ZN(n11536) );
  NAND2_X1 U13416 ( .A1(n15522), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n11526) );
  NAND2_X1 U13417 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11525)
         );
  OAI211_X1 U13418 ( .C1(n14148), .C2(n11527), .A(n11526), .B(n11525), .ZN(
        n11535) );
  OAI21_X1 U13419 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n11529), .A(n11528), .ZN(
        n15589) );
  INV_X1 U13420 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11530) );
  MUX2_X1 U13421 ( .A(n11530), .B(P2_REG1_REG_10__SCAN_IN), .S(n15597), .Z(
        n15590) );
  NOR2_X1 U13422 ( .A1(n15589), .A2(n15590), .ZN(n15587) );
  INV_X1 U13423 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11531) );
  MUX2_X1 U13424 ( .A(n11531), .B(P2_REG1_REG_11__SCAN_IN), .S(n12100), .Z(
        n11532) );
  AOI211_X1 U13425 ( .C1(n11533), .C2(n11532), .A(n15588), .B(n12099), .ZN(
        n11534) );
  AOI211_X1 U13426 ( .C1(n15583), .C2(n11536), .A(n11535), .B(n11534), .ZN(
        n11537) );
  INV_X1 U13427 ( .A(n11537), .ZN(P2_U3225) );
  MUX2_X1 U13428 ( .A(n12384), .B(n11538), .S(n13087), .Z(n12291) );
  XNOR2_X1 U13429 ( .A(n12291), .B(n12303), .ZN(n12293) );
  INV_X1 U13430 ( .A(n11539), .ZN(n11540) );
  MUX2_X1 U13431 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13087), .Z(n11544) );
  XNOR2_X1 U13432 ( .A(n11544), .B(n11553), .ZN(n15687) );
  XOR2_X1 U13433 ( .A(n12293), .B(n12294), .Z(n11563) );
  INV_X1 U13434 ( .A(n12303), .ZN(n12292) );
  INV_X1 U13435 ( .A(n11545), .ZN(n11547) );
  NAND2_X1 U13436 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11553), .ZN(n11548) );
  OAI21_X1 U13437 ( .B1(n11553), .B2(P3_REG1_REG_10__SCAN_IN), .A(n11548), 
        .ZN(n15695) );
  NOR2_X1 U13438 ( .A1(n15696), .A2(n15695), .ZN(n15694) );
  AOI21_X1 U13439 ( .B1(n11549), .B2(n11538), .A(n12281), .ZN(n11551) );
  INV_X1 U13440 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n13464) );
  NOR2_X1 U13441 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13464), .ZN(n12320) );
  AOI21_X1 U13442 ( .B1(n15702), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12320), 
        .ZN(n11550) );
  OAI21_X1 U13443 ( .B1(n11551), .B2(n15718), .A(n11550), .ZN(n11552) );
  AOI21_X1 U13444 ( .B1(n12292), .B2(n15704), .A(n11552), .ZN(n11562) );
  NAND2_X1 U13445 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11553), .ZN(n11558) );
  INV_X1 U13446 ( .A(n11553), .ZN(n15686) );
  AOI22_X1 U13447 ( .A1(n15686), .A2(n8392), .B1(P3_REG2_REG_10__SCAN_IN), 
        .B2(n11553), .ZN(n15691) );
  NAND2_X1 U13448 ( .A1(n11555), .A2(n11554), .ZN(n11557) );
  NAND2_X1 U13449 ( .A1(n11557), .A2(n11556), .ZN(n15690) );
  NAND2_X1 U13450 ( .A1(n15691), .A2(n15690), .ZN(n15689) );
  NAND2_X1 U13451 ( .A1(n11558), .A2(n15689), .ZN(n12304) );
  XNOR2_X1 U13452 ( .A(n12304), .B(n12292), .ZN(n11559) );
  NAND2_X1 U13453 ( .A1(P3_REG2_REG_11__SCAN_IN), .A2(n11559), .ZN(n12305) );
  OAI21_X1 U13454 ( .B1(n11559), .B2(P3_REG2_REG_11__SCAN_IN), .A(n12305), 
        .ZN(n11560) );
  NAND2_X1 U13455 ( .A1(n11560), .A2(n15711), .ZN(n11561) );
  OAI211_X1 U13456 ( .C1(n11563), .C2(n15681), .A(n11562), .B(n11561), .ZN(
        P3_U3193) );
  XOR2_X1 U13457 ( .A(n11578), .B(n14958), .Z(n15831) );
  XNOR2_X1 U13458 ( .A(n11616), .B(n14958), .ZN(n11570) );
  AOI21_X1 U13459 ( .B1(n11570), .B2(n15988), .A(n11569), .ZN(n15829) );
  MUX2_X1 U13460 ( .A(n11571), .B(n15829), .S(n15760), .Z(n11577) );
  INV_X1 U13461 ( .A(n11599), .ZN(n11660) );
  OAI211_X1 U13462 ( .C1(n15830), .C2(n11572), .A(n11660), .B(n15932), .ZN(
        n15828) );
  INV_X1 U13463 ( .A(n15828), .ZN(n11575) );
  OAI22_X1 U13464 ( .A1(n15317), .A2(n15830), .B1(n15755), .B2(n11573), .ZN(
        n11574) );
  AOI21_X1 U13465 ( .B1(n11575), .B2(n15951), .A(n11574), .ZN(n11576) );
  OAI211_X1 U13466 ( .C1(n15831), .C2(n15285), .A(n11577), .B(n11576), .ZN(
        P1_U3286) );
  NAND2_X1 U13467 ( .A1(n11578), .A2(n14958), .ZN(n11580) );
  INV_X1 U13468 ( .A(n11617), .ZN(n15048) );
  OR2_X1 U13469 ( .A1(n14796), .A2(n15048), .ZN(n11579) );
  XNOR2_X1 U13470 ( .A(n15848), .B(n15047), .ZN(n11654) );
  NAND2_X1 U13471 ( .A1(n15848), .A2(n15047), .ZN(n11581) );
  NAND2_X1 U13472 ( .A1(n11582), .A2(n14944), .ZN(n11585) );
  INV_X1 U13473 ( .A(n11583), .ZN(n15112) );
  AOI22_X1 U13474 ( .A1(n12597), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7182), 
        .B2(n15112), .ZN(n11584) );
  XNOR2_X1 U13475 ( .A(n15872), .B(n15046), .ZN(n14960) );
  OR2_X1 U13476 ( .A1(n15872), .A2(n15046), .ZN(n11586) );
  NAND2_X1 U13477 ( .A1(n11587), .A2(n14944), .ZN(n11590) );
  AOI22_X1 U13478 ( .A1(n12597), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n12596), 
        .B2(n11588), .ZN(n11589) );
  NAND2_X2 U13479 ( .A1(n11590), .A2(n11589), .ZN(n14815) );
  NAND2_X1 U13480 ( .A1(n12711), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11597) );
  INV_X1 U13481 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11591) );
  OR2_X1 U13482 ( .A1(n12686), .A2(n11591), .ZN(n11596) );
  NOR2_X1 U13483 ( .A1(n11592), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11593) );
  OR2_X1 U13484 ( .A1(n11603), .A2(n11593), .ZN(n11822) );
  OR2_X1 U13485 ( .A1(n7189), .A2(n11822), .ZN(n11595) );
  OR2_X1 U13486 ( .A1(n12705), .A2(n10404), .ZN(n11594) );
  OR2_X1 U13487 ( .A1(n14815), .A2(n11817), .ZN(n11741) );
  NAND2_X1 U13488 ( .A1(n14815), .A2(n11817), .ZN(n11598) );
  NAND2_X1 U13489 ( .A1(n11741), .A2(n11598), .ZN(n14959) );
  XNOR2_X1 U13490 ( .A(n11764), .B(n14959), .ZN(n15898) );
  INV_X1 U13491 ( .A(n15898), .ZN(n11628) );
  NAND2_X1 U13492 ( .A1(n11721), .A2(n14815), .ZN(n11600) );
  NAND2_X1 U13493 ( .A1(n11600), .A2(n15932), .ZN(n11601) );
  OR2_X1 U13494 ( .A1(n11760), .A2(n11601), .ZN(n11610) );
  NAND2_X1 U13495 ( .A1(n14924), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n11608) );
  OR2_X1 U13496 ( .A1(n14928), .A2(n11602), .ZN(n11607) );
  OR2_X1 U13497 ( .A1(n11603), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11604) );
  NAND2_X1 U13498 ( .A1(n11750), .A2(n11604), .ZN(n11914) );
  OR2_X1 U13499 ( .A1(n7189), .A2(n11914), .ZN(n11606) );
  OR2_X1 U13500 ( .A1(n12705), .A2(n10406), .ZN(n11605) );
  OR2_X1 U13501 ( .A1(n12269), .A2(n15195), .ZN(n11609) );
  AND2_X1 U13502 ( .A1(n11610), .A2(n11609), .ZN(n15892) );
  INV_X1 U13503 ( .A(n15892), .ZN(n11614) );
  INV_X1 U13504 ( .A(n14815), .ZN(n15893) );
  NAND2_X1 U13505 ( .A1(n15046), .A2(n15289), .ZN(n15891) );
  OAI22_X1 U13506 ( .A1(n15946), .A2(n15891), .B1(n11822), .B2(n15755), .ZN(
        n11611) );
  AOI21_X1 U13507 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n15946), .A(n11611), 
        .ZN(n11612) );
  OAI21_X1 U13508 ( .B1(n15893), .B2(n15317), .A(n11612), .ZN(n11613) );
  AOI21_X1 U13509 ( .B1(n11614), .B2(n15951), .A(n11613), .ZN(n11627) );
  NAND2_X1 U13510 ( .A1(n14796), .A2(n11617), .ZN(n11615) );
  NAND2_X1 U13511 ( .A1(n11616), .A2(n11615), .ZN(n11619) );
  OR2_X1 U13512 ( .A1(n14796), .A2(n11617), .ZN(n11618) );
  NAND2_X1 U13513 ( .A1(n11619), .A2(n11618), .ZN(n11653) );
  OR2_X1 U13514 ( .A1(n15848), .A2(n11620), .ZN(n11621) );
  NAND2_X1 U13515 ( .A1(n15872), .A2(n11821), .ZN(n11622) );
  NAND2_X1 U13516 ( .A1(n11625), .A2(n14959), .ZN(n15894) );
  NAND2_X1 U13517 ( .A1(n15760), .A2(n15988), .ZN(n15337) );
  INV_X1 U13518 ( .A(n15337), .ZN(n12224) );
  NAND3_X1 U13519 ( .A1(n15895), .A2(n15894), .A3(n12224), .ZN(n11626) );
  OAI211_X1 U13520 ( .C1(n11628), .C2(n15285), .A(n11627), .B(n11626), .ZN(
        P1_U3283) );
  AOI21_X1 U13521 ( .B1(n15841), .B2(n11879), .A(n11629), .ZN(n11630) );
  OAI211_X1 U13522 ( .C1(n11632), .C2(n14442), .A(n11631), .B(n11630), .ZN(
        n11634) );
  NAND2_X1 U13523 ( .A1(n11634), .A2(n14451), .ZN(n11633) );
  OAI21_X1 U13524 ( .B1(n14451), .B2(n11531), .A(n11633), .ZN(P2_U3510) );
  INV_X1 U13525 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11636) );
  NAND2_X1 U13526 ( .A1(n11634), .A2(n14469), .ZN(n11635) );
  OAI21_X1 U13527 ( .B1(n14469), .B2(n11636), .A(n11635), .ZN(P2_U3463) );
  INV_X1 U13528 ( .A(n15872), .ZN(n11651) );
  INV_X1 U13529 ( .A(n11637), .ZN(n11640) );
  INV_X1 U13530 ( .A(n11638), .ZN(n11639) );
  NAND2_X1 U13531 ( .A1(n15872), .A2(n14581), .ZN(n11642) );
  NAND2_X1 U13532 ( .A1(n15046), .A2(n14587), .ZN(n11641) );
  NAND2_X1 U13533 ( .A1(n11642), .A2(n11641), .ZN(n11643) );
  XNOR2_X1 U13534 ( .A(n11643), .B(n14628), .ZN(n11814) );
  AND2_X1 U13535 ( .A1(n15046), .A2(n14563), .ZN(n11644) );
  AOI21_X1 U13536 ( .B1(n15872), .B2(n14587), .A(n11644), .ZN(n11816) );
  XNOR2_X1 U13537 ( .A(n11814), .B(n11816), .ZN(n11645) );
  NAND2_X1 U13538 ( .A1(n11646), .A2(n11645), .ZN(n11815) );
  OAI211_X1 U13539 ( .C1(n11646), .C2(n11645), .A(n11815), .B(n14716), .ZN(
        n11650) );
  INV_X1 U13540 ( .A(n11723), .ZN(n11648) );
  INV_X1 U13541 ( .A(n14746), .ZN(n14667) );
  INV_X1 U13542 ( .A(n11817), .ZN(n15045) );
  AOI22_X1 U13543 ( .A1(n15045), .A2(n15342), .B1(n15289), .B2(n15047), .ZN(
        n11715) );
  NAND2_X1 U13544 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n15109) );
  OAI21_X1 U13545 ( .B1(n11715), .B2(n14665), .A(n15109), .ZN(n11647) );
  AOI21_X1 U13546 ( .B1(n11648), .B2(n14667), .A(n11647), .ZN(n11649) );
  OAI211_X1 U13547 ( .C1(n11651), .C2(n14725), .A(n11650), .B(n11649), .ZN(
        P1_U3231) );
  INV_X1 U13548 ( .A(n11654), .ZN(n14957) );
  XNOR2_X1 U13549 ( .A(n11652), .B(n14957), .ZN(n11658) );
  INV_X1 U13550 ( .A(n11658), .ZN(n15851) );
  XNOR2_X1 U13551 ( .A(n11653), .B(n11654), .ZN(n11656) );
  AOI22_X1 U13552 ( .A1(n15048), .A2(n15289), .B1(n15342), .B2(n15046), .ZN(
        n11655) );
  OAI21_X1 U13553 ( .B1(n11656), .B2(n15959), .A(n11655), .ZN(n11657) );
  AOI21_X1 U13554 ( .B1(n15880), .B2(n11658), .A(n11657), .ZN(n15850) );
  MUX2_X1 U13555 ( .A(n10383), .B(n15850), .S(n15760), .Z(n11665) );
  INV_X1 U13556 ( .A(n11720), .ZN(n11659) );
  AOI211_X1 U13557 ( .C1(n15848), .C2(n11660), .A(n15354), .B(n11659), .ZN(
        n15847) );
  OAI22_X1 U13558 ( .A1(n11662), .A2(n15317), .B1(n11661), .B2(n15755), .ZN(
        n11663) );
  AOI21_X1 U13559 ( .B1(n15847), .B2(n15951), .A(n11663), .ZN(n11664) );
  OAI211_X1 U13560 ( .C1(n15851), .C2(n15363), .A(n11665), .B(n11664), .ZN(
        P1_U3285) );
  OAI21_X1 U13561 ( .B1(n11667), .B2(n13054), .A(n11666), .ZN(n15799) );
  OAI211_X1 U13562 ( .C1(n11670), .C2(n11669), .A(n11668), .B(n13756), .ZN(
        n11672) );
  AOI22_X1 U13563 ( .A1(n13483), .A2(n13759), .B1(n13742), .B2(n13481), .ZN(
        n11671) );
  NAND2_X1 U13564 ( .A1(n11672), .A2(n11671), .ZN(n15798) );
  AOI21_X1 U13565 ( .B1(n15917), .B2(n15799), .A(n15798), .ZN(n11677) );
  OAI22_X1 U13566 ( .A1(n13960), .A2(n15805), .B1(n16000), .B2(n8358), .ZN(
        n11673) );
  INV_X1 U13567 ( .A(n11673), .ZN(n11674) );
  OAI21_X1 U13568 ( .B1(n11677), .B2(n16008), .A(n11674), .ZN(P3_U3408) );
  AOI22_X1 U13569 ( .A1(n16005), .A2(n11675), .B1(n16004), .B2(
        P3_REG1_REG_6__SCAN_IN), .ZN(n11676) );
  OAI21_X1 U13570 ( .B1(n11677), .B2(n16004), .A(n11676), .ZN(P3_U3465) );
  NOR2_X1 U13571 ( .A1(n15804), .A2(n10660), .ZN(n11679) );
  AOI211_X1 U13572 ( .C1(n11680), .C2(n12908), .A(n11679), .B(n11678), .ZN(
        n11684) );
  NAND2_X1 U13573 ( .A1(n15810), .A2(n11681), .ZN(n13702) );
  INV_X1 U13574 ( .A(n13702), .ZN(n11946) );
  AOI22_X1 U13575 ( .A1(n11682), .A2(n11946), .B1(n15802), .B2(
        P3_REG2_REG_2__SCAN_IN), .ZN(n11683) );
  OAI21_X1 U13576 ( .B1(n11684), .B2(n15802), .A(n11683), .ZN(P3_U3231) );
  OAI21_X1 U13577 ( .B1(n11686), .B2(n11696), .A(n11685), .ZN(n15795) );
  OAI211_X1 U13578 ( .C1(n11688), .C2(n15790), .A(n15932), .B(n11687), .ZN(
        n15789) );
  NOR2_X1 U13579 ( .A1(n15755), .A2(n11689), .ZN(n11690) );
  AOI21_X1 U13580 ( .B1(n15947), .B2(n14783), .A(n11690), .ZN(n11694) );
  INV_X1 U13581 ( .A(n11691), .ZN(n15788) );
  MUX2_X1 U13582 ( .A(n11692), .B(n15788), .S(n15760), .Z(n11693) );
  OAI211_X1 U13583 ( .C1(n15789), .C2(n15358), .A(n11694), .B(n11693), .ZN(
        n11698) );
  NAND2_X1 U13584 ( .A1(n11695), .A2(n11696), .ZN(n15791) );
  AND3_X1 U13585 ( .A1(n15792), .A2(n12224), .A3(n15791), .ZN(n11697) );
  AOI211_X1 U13586 ( .C1(n15952), .C2(n15795), .A(n11698), .B(n11697), .ZN(
        n11699) );
  INV_X1 U13587 ( .A(n11699), .ZN(P1_U3289) );
  INV_X1 U13588 ( .A(n12591), .ZN(n11774) );
  NAND2_X1 U13589 ( .A1(n11700), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11701) );
  XNOR2_X1 U13590 ( .A(n11701), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15129) );
  AOI22_X1 U13591 ( .A1(n15129), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n11702), .ZN(n11703) );
  OAI21_X1 U13592 ( .B1(n11774), .B2(n13160), .A(n11703), .ZN(P1_U3337) );
  INV_X1 U13593 ( .A(n12608), .ZN(n11867) );
  OAI222_X1 U13594 ( .A1(n15476), .A2(n12609), .B1(n13160), .B2(n11867), .C1(
        n7187), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U13595 ( .A(n11704), .ZN(n11713) );
  OAI22_X1 U13596 ( .A1(n15760), .A2(n11706), .B1(n11705), .B2(n15755), .ZN(
        n11707) );
  AOI21_X1 U13597 ( .B1(n15947), .B2(n14787), .A(n11707), .ZN(n11708) );
  OAI21_X1 U13598 ( .B1(n11709), .B2(n15358), .A(n11708), .ZN(n11710) );
  AOI21_X1 U13599 ( .B1(n11711), .B2(n15952), .A(n11710), .ZN(n11712) );
  OAI21_X1 U13600 ( .B1(n11713), .B2(n15946), .A(n11712), .ZN(P1_U3288) );
  XNOR2_X1 U13601 ( .A(n11714), .B(n14960), .ZN(n11716) );
  OAI21_X1 U13602 ( .B1(n11716), .B2(n15959), .A(n11715), .ZN(n15878) );
  INV_X1 U13603 ( .A(n15878), .ZN(n11728) );
  INV_X1 U13604 ( .A(n11717), .ZN(n11718) );
  AOI21_X1 U13605 ( .B1(n14960), .B2(n11719), .A(n11718), .ZN(n15876) );
  INV_X1 U13606 ( .A(n15876), .ZN(n15879) );
  AOI21_X1 U13607 ( .B1(n11720), .B2(n15872), .A(n15354), .ZN(n11722) );
  NAND2_X1 U13608 ( .A1(n11722), .A2(n11721), .ZN(n15874) );
  OAI22_X1 U13609 ( .A1(n15760), .A2(n10403), .B1(n11723), .B2(n15755), .ZN(
        n11724) );
  AOI21_X1 U13610 ( .B1(n15872), .B2(n15947), .A(n11724), .ZN(n11725) );
  OAI21_X1 U13611 ( .B1(n15874), .B2(n15358), .A(n11725), .ZN(n11726) );
  AOI21_X1 U13612 ( .B1(n15879), .B2(n15952), .A(n11726), .ZN(n11727) );
  OAI21_X1 U13613 ( .B1(n15946), .B2(n11728), .A(n11727), .ZN(P1_U3284) );
  INV_X1 U13614 ( .A(n11729), .ZN(n11730) );
  INV_X1 U13615 ( .A(n15755), .ZN(n15944) );
  AOI22_X1 U13616 ( .A1(n11731), .A2(n11730), .B1(n15944), .B2(n10352), .ZN(
        n11732) );
  AND2_X1 U13617 ( .A1(n11733), .A2(n11732), .ZN(n11735) );
  MUX2_X1 U13618 ( .A(n11735), .B(n11734), .S(n15946), .Z(n11738) );
  AOI22_X1 U13619 ( .A1(n11736), .A2(n15952), .B1(n15947), .B2(n14776), .ZN(
        n11737) );
  NAND2_X1 U13620 ( .A1(n11738), .A2(n11737), .ZN(P1_U3290) );
  NAND2_X1 U13621 ( .A1(n11739), .A2(n13973), .ZN(n11740) );
  OAI211_X1 U13622 ( .C1(n13390), .C2(n13969), .A(n11740), .B(n13091), .ZN(
        P3_U3272) );
  NAND2_X1 U13623 ( .A1(n11742), .A2(n14944), .ZN(n11745) );
  AOI22_X1 U13624 ( .A1(n12597), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7182), 
        .B2(n11743), .ZN(n11744) );
  NAND2_X1 U13625 ( .A1(n11745), .A2(n11744), .ZN(n15922) );
  OR2_X1 U13626 ( .A1(n15922), .A2(n12269), .ZN(n11997) );
  NAND2_X1 U13627 ( .A1(n15922), .A2(n12269), .ZN(n11746) );
  NAND2_X1 U13628 ( .A1(n11747), .A2(n14962), .ZN(n11998) );
  OAI211_X1 U13629 ( .C1(n11747), .C2(n14962), .A(n11998), .B(n15988), .ZN(
        n11759) );
  OR2_X1 U13630 ( .A1(n11817), .A2(n15345), .ZN(n11757) );
  NAND2_X1 U13631 ( .A1(n12711), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11755) );
  INV_X1 U13632 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11748) );
  OR2_X1 U13633 ( .A1(n12686), .A2(n11748), .ZN(n11754) );
  NAND2_X1 U13634 ( .A1(n11750), .A2(n11749), .ZN(n11751) );
  NAND2_X1 U13635 ( .A1(n11977), .A2(n11751), .ZN(n15943) );
  OR2_X1 U13636 ( .A1(n7189), .A2(n15943), .ZN(n11753) );
  OR2_X1 U13637 ( .A1(n12705), .A2(n10697), .ZN(n11752) );
  NAND4_X1 U13638 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n15043) );
  NAND2_X1 U13639 ( .A1(n15043), .A2(n15342), .ZN(n11756) );
  NAND2_X1 U13640 ( .A1(n11757), .A2(n11756), .ZN(n11917) );
  INV_X1 U13641 ( .A(n11917), .ZN(n11758) );
  NAND2_X1 U13642 ( .A1(n11759), .A2(n11758), .ZN(n15920) );
  INV_X1 U13643 ( .A(n15920), .ZN(n11772) );
  OAI21_X1 U13644 ( .B1(n11760), .B2(n11920), .A(n15932), .ZN(n11761) );
  NOR2_X1 U13645 ( .A1(n11761), .A2(n15933), .ZN(n15921) );
  NOR2_X1 U13646 ( .A1(n11920), .A2(n15317), .ZN(n11763) );
  OAI22_X1 U13647 ( .A1(n15760), .A2(n10406), .B1(n11914), .B2(n15755), .ZN(
        n11762) );
  AOI211_X1 U13648 ( .C1(n15921), .C2(n15951), .A(n11763), .B(n11762), .ZN(
        n11771) );
  NAND2_X1 U13649 ( .A1(n11764), .A2(n14959), .ZN(n11766) );
  OR2_X1 U13650 ( .A1(n14815), .A2(n15045), .ZN(n11765) );
  NAND2_X1 U13651 ( .A1(n11766), .A2(n11765), .ZN(n11769) );
  INV_X1 U13652 ( .A(n11769), .ZN(n11768) );
  NAND2_X1 U13653 ( .A1(n11768), .A2(n11767), .ZN(n11963) );
  NAND2_X1 U13654 ( .A1(n11769), .A2(n14962), .ZN(n15923) );
  NAND3_X1 U13655 ( .A1(n11963), .A2(n15923), .A3(n15952), .ZN(n11770) );
  OAI211_X1 U13656 ( .C1(n11772), .C2(n15946), .A(n11771), .B(n11770), .ZN(
        P1_U3282) );
  INV_X1 U13657 ( .A(n14122), .ZN(n14129) );
  OAI222_X1 U13658 ( .A1(P2_U3088), .A2(n14129), .B1(n14477), .B2(n11774), 
        .C1(n11773), .C2(n13150), .ZN(P2_U3309) );
  INV_X1 U13659 ( .A(n11775), .ZN(n12846) );
  NAND2_X1 U13660 ( .A1(n12846), .A2(n11776), .ZN(n11777) );
  NAND2_X1 U13661 ( .A1(n11778), .A2(n11777), .ZN(n11780) );
  XNOR2_X1 U13662 ( .A(n12854), .B(n12116), .ZN(n12788) );
  NAND2_X1 U13663 ( .A1(n14074), .A2(n12832), .ZN(n11781) );
  XNOR2_X1 U13664 ( .A(n12788), .B(n11781), .ZN(n12845) );
  NAND2_X1 U13665 ( .A1(n11780), .A2(n12845), .ZN(n12787) );
  INV_X1 U13666 ( .A(n12788), .ZN(n11782) );
  NAND2_X1 U13667 ( .A1(n11782), .A2(n11781), .ZN(n11783) );
  NAND2_X1 U13668 ( .A1(n12787), .A2(n11783), .ZN(n11784) );
  XNOR2_X1 U13669 ( .A(n12797), .B(n12116), .ZN(n11785) );
  NAND2_X1 U13670 ( .A1(n14073), .A2(n12832), .ZN(n11786) );
  XNOR2_X1 U13671 ( .A(n11785), .B(n11786), .ZN(n12786) );
  NAND2_X1 U13672 ( .A1(n11784), .A2(n12786), .ZN(n12803) );
  INV_X1 U13673 ( .A(n11785), .ZN(n11787) );
  NAND2_X1 U13674 ( .A1(n11787), .A2(n11786), .ZN(n11788) );
  NAND2_X1 U13675 ( .A1(n12803), .A2(n11788), .ZN(n11875) );
  AND2_X1 U13676 ( .A1(n14072), .A2(n12832), .ZN(n11789) );
  NAND2_X1 U13677 ( .A1(n13136), .A2(n11789), .ZN(n11795) );
  INV_X1 U13678 ( .A(n11789), .ZN(n11790) );
  NAND2_X1 U13679 ( .A1(n11791), .A2(n11790), .ZN(n11792) );
  NAND2_X1 U13680 ( .A1(n11795), .A2(n11792), .ZN(n11876) );
  INV_X1 U13681 ( .A(n11876), .ZN(n11793) );
  XNOR2_X1 U13682 ( .A(n11881), .B(n12116), .ZN(n11802) );
  NAND2_X1 U13683 ( .A1(n14071), .A2(n12832), .ZN(n11797) );
  XNOR2_X1 U13684 ( .A(n11802), .B(n11797), .ZN(n13139) );
  INV_X1 U13685 ( .A(n11802), .ZN(n11798) );
  XNOR2_X1 U13686 ( .A(n12134), .B(n12116), .ZN(n11896) );
  NAND2_X1 U13687 ( .A1(n13141), .A2(n12832), .ZN(n11890) );
  XNOR2_X1 U13688 ( .A(n11896), .B(n11890), .ZN(n11803) );
  INV_X1 U13689 ( .A(n12060), .ZN(n11800) );
  INV_X1 U13690 ( .A(n14031), .ZN(n14047) );
  AOI22_X1 U13691 ( .A1(n13142), .A2(n14070), .B1(n14047), .B2(n14071), .ZN(
        n11799) );
  NAND2_X1 U13692 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n12106)
         );
  OAI211_X1 U13693 ( .C1(n11800), .C2(n14030), .A(n11799), .B(n12106), .ZN(
        n11807) );
  INV_X1 U13694 ( .A(n11801), .ZN(n11805) );
  AOI22_X1 U13695 ( .A1(n11802), .A2(n14054), .B1(n13994), .B2(n14071), .ZN(
        n11804) );
  NOR3_X1 U13696 ( .A1(n11805), .A2(n11804), .A3(n11803), .ZN(n11806) );
  AOI211_X1 U13697 ( .C1(n12134), .C2(n14035), .A(n11807), .B(n11806), .ZN(
        n11808) );
  OAI21_X1 U13698 ( .B1(n11893), .B2(n10844), .A(n11808), .ZN(P2_U3206) );
  MUX2_X1 U13699 ( .A(n11810), .B(n11809), .S(n15997), .Z(n11813) );
  AOI22_X1 U13700 ( .A1(n11945), .A2(n12153), .B1(n11811), .B2(n16005), .ZN(
        n11812) );
  NAND2_X1 U13701 ( .A1(n11813), .A2(n11812), .ZN(P3_U3464) );
  NOR2_X1 U13702 ( .A1(n11817), .A2(n14626), .ZN(n11818) );
  AOI21_X1 U13703 ( .B1(n14815), .B2(n14587), .A(n11818), .ZN(n11904) );
  AOI22_X1 U13704 ( .A1(n14815), .A2(n14581), .B1(n14587), .B2(n15045), .ZN(
        n11819) );
  XNOR2_X1 U13705 ( .A(n11819), .B(n14628), .ZN(n11905) );
  XOR2_X1 U13706 ( .A(n11904), .B(n11905), .Z(n11908) );
  XNOR2_X1 U13707 ( .A(n11909), .B(n11908), .ZN(n11826) );
  OAI21_X1 U13708 ( .B1(n14743), .B2(n11821), .A(n11820), .ZN(n11824) );
  OAI22_X1 U13709 ( .A1(n12269), .A2(n14747), .B1(n14746), .B2(n11822), .ZN(
        n11823) );
  OAI21_X1 U13710 ( .B1(n11826), .B2(n14753), .A(n11825), .ZN(P1_U3217) );
  OAI21_X1 U13711 ( .B1(n11828), .B2(n12926), .A(n11827), .ZN(n12039) );
  OAI211_X1 U13712 ( .C1(n11829), .C2(n7766), .A(n11922), .B(n13756), .ZN(
        n11832) );
  OAI22_X1 U13713 ( .A1(n11935), .A2(n13833), .B1(n12892), .B2(n13835), .ZN(
        n11830) );
  INV_X1 U13714 ( .A(n11830), .ZN(n11831) );
  NAND2_X1 U13715 ( .A1(n11832), .A2(n11831), .ZN(n12036) );
  AOI21_X1 U13716 ( .B1(n15917), .B2(n12039), .A(n12036), .ZN(n11838) );
  INV_X1 U13717 ( .A(n11836), .ZN(n12928) );
  INV_X1 U13718 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n11833) );
  OAI22_X1 U13719 ( .A1(n13960), .A2(n12928), .B1(n16000), .B2(n11833), .ZN(
        n11834) );
  INV_X1 U13720 ( .A(n11834), .ZN(n11835) );
  OAI21_X1 U13721 ( .B1(n11838), .B2(n16008), .A(n11835), .ZN(P3_U3411) );
  AOI22_X1 U13722 ( .A1(n16005), .A2(n11836), .B1(n16004), .B2(
        P3_REG1_REG_7__SCAN_IN), .ZN(n11837) );
  OAI21_X1 U13723 ( .B1(n11838), .B2(n16004), .A(n11837), .ZN(P3_U3466) );
  INV_X1 U13724 ( .A(n12621), .ZN(n11861) );
  OAI222_X1 U13725 ( .A1(n15476), .A2(n12622), .B1(n13160), .B2(n11861), .C1(
        n14940), .C2(P1_U3086), .ZN(P1_U3334) );
  XNOR2_X1 U13726 ( .A(n11839), .B(n11841), .ZN(n11885) );
  AOI22_X1 U13727 ( .A1(n13141), .A2(n14355), .B1(n14072), .B2(n14353), .ZN(
        n11844) );
  OAI211_X1 U13728 ( .C1(n11842), .C2(n11841), .A(n11840), .B(n14358), .ZN(
        n11843) );
  OAI211_X1 U13729 ( .C1(n11885), .C2(n10019), .A(n11844), .B(n11843), .ZN(
        n11845) );
  INV_X1 U13730 ( .A(n11845), .ZN(n11884) );
  INV_X1 U13731 ( .A(n11846), .ZN(n11848) );
  INV_X1 U13732 ( .A(n12059), .ZN(n11847) );
  AOI21_X1 U13733 ( .B1(n11881), .B2(n11848), .A(n11847), .ZN(n11882) );
  AOI22_X1 U13734 ( .A1(n14359), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n13140), 
        .B2(n14345), .ZN(n11849) );
  OAI21_X1 U13735 ( .B1(n13145), .B2(n14349), .A(n11849), .ZN(n11851) );
  NOR2_X1 U13736 ( .A1(n11885), .A2(n14231), .ZN(n11850) );
  AOI211_X1 U13737 ( .C1(n11882), .C2(n14362), .A(n11851), .B(n11850), .ZN(
        n11852) );
  OAI21_X1 U13738 ( .B1(n14359), .B2(n11884), .A(n11852), .ZN(P2_U3253) );
  AOI211_X1 U13739 ( .C1(n11854), .C2(n11853), .A(n13222), .B(n7342), .ZN(
        n11855) );
  INV_X1 U13740 ( .A(n11855), .ZN(n11860) );
  OAI22_X1 U13741 ( .A1(n13255), .A2(n15805), .B1(n11856), .B2(n13247), .ZN(
        n11857) );
  AOI211_X1 U13742 ( .C1(n13245), .C2(n13481), .A(n11858), .B(n11857), .ZN(
        n11859) );
  OAI211_X1 U13743 ( .C1(n15803), .C2(n13200), .A(n11860), .B(n11859), .ZN(
        P3_U3179) );
  OAI222_X1 U13744 ( .A1(n13150), .A2(n11863), .B1(P2_U3088), .B2(n11862), 
        .C1(n14477), .C2(n11861), .ZN(P2_U3306) );
  INV_X1 U13745 ( .A(n12595), .ZN(n11865) );
  OAI222_X1 U13746 ( .A1(n13150), .A2(n11864), .B1(n14477), .B2(n11865), .C1(
        n9722), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13747 ( .A1(n15476), .A2(n11866), .B1(n13160), .B2(n11865), .C1(
        P1_U3086), .C2(n10342), .ZN(P1_U3336) );
  OAI222_X1 U13748 ( .A1(n13150), .A2(n11869), .B1(P2_U3088), .B2(n11868), 
        .C1(n14477), .C2(n11867), .ZN(P2_U3307) );
  INV_X1 U13749 ( .A(n11870), .ZN(n11873) );
  INV_X1 U13750 ( .A(n14002), .ZN(n14023) );
  AOI22_X1 U13751 ( .A1(n14023), .A2(n11871), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11872) );
  OAI21_X1 U13752 ( .B1(n11873), .B2(n14030), .A(n11872), .ZN(n11878) );
  INV_X1 U13753 ( .A(n13138), .ZN(n11874) );
  AOI211_X1 U13754 ( .C1(n11876), .C2(n11875), .A(n10844), .B(n11874), .ZN(
        n11877) );
  AOI211_X1 U13755 ( .C1(n11879), .C2(n14035), .A(n11878), .B(n11877), .ZN(
        n11880) );
  INV_X1 U13756 ( .A(n11880), .ZN(P2_U3208) );
  INV_X1 U13757 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U13758 ( .A1(n11882), .A2(n14445), .B1(n15841), .B2(n11881), .ZN(
        n11883) );
  OAI211_X1 U13759 ( .C1(n11885), .C2(n14449), .A(n11884), .B(n11883), .ZN(
        n11888) );
  NAND2_X1 U13760 ( .A1(n11888), .A2(n14469), .ZN(n11886) );
  OAI21_X1 U13761 ( .B1(n14469), .B2(n11887), .A(n11886), .ZN(P2_U3466) );
  INV_X1 U13762 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n12102) );
  NAND2_X1 U13763 ( .A1(n11888), .A2(n14451), .ZN(n11889) );
  OAI21_X1 U13764 ( .B1(n14451), .B2(n12102), .A(n11889), .ZN(P2_U3511) );
  INV_X1 U13765 ( .A(n11896), .ZN(n11891) );
  NAND2_X1 U13766 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  XNOR2_X1 U13767 ( .A(n12126), .B(n12116), .ZN(n12119) );
  NAND2_X1 U13768 ( .A1(n14070), .A2(n12832), .ZN(n12112) );
  XNOR2_X1 U13769 ( .A(n12119), .B(n12112), .ZN(n11897) );
  NAND2_X1 U13770 ( .A1(n11894), .A2(n11897), .ZN(n12115) );
  AOI22_X1 U13771 ( .A1(n14047), .A2(n13141), .B1(n13142), .B2(n14069), .ZN(
        n11895) );
  NAND2_X1 U13772 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n12371)
         );
  OAI211_X1 U13773 ( .C1(n11954), .C2(n14030), .A(n11895), .B(n12371), .ZN(
        n11901) );
  INV_X1 U13774 ( .A(n11893), .ZN(n11899) );
  AOI22_X1 U13775 ( .A1(n11896), .A2(n14054), .B1(n13994), .B2(n13141), .ZN(
        n11898) );
  NOR3_X1 U13776 ( .A1(n11899), .A2(n11898), .A3(n11897), .ZN(n11900) );
  AOI211_X1 U13777 ( .C1(n12126), .C2(n14035), .A(n11901), .B(n11900), .ZN(
        n11902) );
  OAI21_X1 U13778 ( .B1(n12115), .B2(n10844), .A(n11902), .ZN(P2_U3187) );
  OAI22_X1 U13779 ( .A1(n11920), .A2(n14572), .B1(n12269), .B2(n14626), .ZN(
        n12230) );
  OAI22_X1 U13780 ( .A1(n11920), .A2(n14627), .B1(n12269), .B2(n14572), .ZN(
        n11903) );
  XNOR2_X1 U13781 ( .A(n11903), .B(n14628), .ZN(n12229) );
  XOR2_X1 U13782 ( .A(n12230), .B(n12229), .Z(n11911) );
  INV_X1 U13783 ( .A(n11904), .ZN(n11907) );
  INV_X1 U13784 ( .A(n11905), .ZN(n11906) );
  OAI21_X1 U13785 ( .B1(n11911), .B2(n11910), .A(n12228), .ZN(n11912) );
  NAND2_X1 U13786 ( .A1(n11912), .A2(n14716), .ZN(n11919) );
  INV_X1 U13787 ( .A(n11913), .ZN(n11916) );
  NOR2_X1 U13788 ( .A1(n14746), .A2(n11914), .ZN(n11915) );
  AOI211_X1 U13789 ( .C1(n14694), .C2(n11917), .A(n11916), .B(n11915), .ZN(
        n11918) );
  OAI211_X1 U13790 ( .C1(n11920), .C2(n14725), .A(n11919), .B(n11918), .ZN(
        P1_U3236) );
  AND2_X1 U13791 ( .A1(n11922), .A2(n11921), .ZN(n11924) );
  OAI21_X1 U13792 ( .B1(n13059), .B2(n11924), .A(n11923), .ZN(n11925) );
  AOI222_X1 U13793 ( .A1(n13756), .A2(n11925), .B1(n13481), .B2(n13759), .C1(
        n7681), .C2(n13742), .ZN(n12147) );
  OAI21_X1 U13794 ( .B1(n11928), .B2(n11927), .A(n11926), .ZN(n12154) );
  NOR2_X1 U13795 ( .A1(n15810), .A2(n8244), .ZN(n11930) );
  OAI22_X1 U13796 ( .A1(n15806), .A2(n12891), .B1(n12090), .B2(n15804), .ZN(
        n11929) );
  AOI211_X1 U13797 ( .C1(n12154), .C2(n13820), .A(n11930), .B(n11929), .ZN(
        n11931) );
  OAI21_X1 U13798 ( .B1(n12147), .B2(n15802), .A(n11931), .ZN(P3_U3225) );
  XOR2_X1 U13799 ( .A(n11933), .B(n11932), .Z(n11934) );
  NAND2_X1 U13800 ( .A1(n11934), .A2(n13241), .ZN(n11939) );
  OAI22_X1 U13801 ( .A1(n13255), .A2(n12928), .B1(n11935), .B2(n13247), .ZN(
        n11936) );
  AOI211_X1 U13802 ( .C1(n13245), .C2(n13480), .A(n11937), .B(n11936), .ZN(
        n11938) );
  OAI211_X1 U13803 ( .C1(n13200), .C2(n12035), .A(n11939), .B(n11938), .ZN(
        P3_U3153) );
  OAI22_X1 U13804 ( .A1(n15806), .A2(n11941), .B1(n11940), .B2(n15804), .ZN(
        n11944) );
  MUX2_X1 U13805 ( .A(n11942), .B(P3_REG2_REG_5__SCAN_IN), .S(n15802), .Z(
        n11943) );
  AOI211_X1 U13806 ( .C1(n11946), .C2(n11945), .A(n11944), .B(n11943), .ZN(
        n11947) );
  INV_X1 U13807 ( .A(n11947), .ZN(P3_U3228) );
  XNOR2_X1 U13808 ( .A(n11948), .B(n11951), .ZN(n11949) );
  AOI222_X1 U13809 ( .A1(n14358), .A2(n11949), .B1(n14069), .B2(n14355), .C1(
        n13141), .C2(n14353), .ZN(n12129) );
  OAI21_X1 U13810 ( .B1(n11952), .B2(n11951), .A(n11950), .ZN(n12130) );
  NAND2_X1 U13811 ( .A1(n14347), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11953) );
  OAI21_X1 U13812 ( .B1(n14308), .B2(n11954), .A(n11953), .ZN(n11955) );
  AOI21_X1 U13813 ( .B1(n12126), .B2(n14271), .A(n11955), .ZN(n11959) );
  NAND2_X1 U13814 ( .A1(n12126), .A2(n12057), .ZN(n11957) );
  AND2_X1 U13815 ( .A1(n12401), .A2(n11957), .ZN(n12127) );
  NAND2_X1 U13816 ( .A1(n12127), .A2(n14362), .ZN(n11958) );
  OAI211_X1 U13817 ( .C1(n12130), .C2(n14364), .A(n11959), .B(n11958), .ZN(
        n11960) );
  INV_X1 U13818 ( .A(n11960), .ZN(n11961) );
  OAI21_X1 U13819 ( .B1(n14347), .B2(n12129), .A(n11961), .ZN(P2_U3251) );
  INV_X1 U13820 ( .A(n12269), .ZN(n15044) );
  NAND2_X1 U13821 ( .A1(n15922), .A2(n15044), .ZN(n11962) );
  NAND2_X1 U13822 ( .A1(n11963), .A2(n11962), .ZN(n11964) );
  NAND2_X1 U13823 ( .A1(n11965), .A2(n14944), .ZN(n11968) );
  AOI22_X1 U13824 ( .A1(n12597), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n12596), 
        .B2(n11966), .ZN(n11967) );
  NAND2_X2 U13825 ( .A1(n11968), .A2(n11967), .ZN(n15948) );
  XNOR2_X1 U13826 ( .A(n15948), .B(n15043), .ZN(n15928) );
  OR2_X1 U13827 ( .A1(n15948), .A2(n15043), .ZN(n11970) );
  NAND2_X1 U13828 ( .A1(n11971), .A2(n14944), .ZN(n11974) );
  AOI22_X1 U13829 ( .A1(n12597), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n12596), 
        .B2(n11972), .ZN(n11973) );
  NAND2_X1 U13830 ( .A1(n12711), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11983) );
  INV_X1 U13831 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11975) );
  OR2_X1 U13832 ( .A1(n12686), .A2(n11975), .ZN(n11982) );
  NAND2_X1 U13833 ( .A1(n11977), .A2(n11976), .ZN(n11978) );
  NAND2_X1 U13834 ( .A1(n11986), .A2(n11978), .ZN(n12238) );
  OR2_X1 U13835 ( .A1(n7189), .A2(n12238), .ZN(n11981) );
  OR2_X1 U13836 ( .A1(n12705), .A2(n11979), .ZN(n11980) );
  XNOR2_X1 U13837 ( .A(n14828), .B(n12268), .ZN(n14964) );
  XNOR2_X1 U13838 ( .A(n12026), .B(n14964), .ZN(n15964) );
  INV_X1 U13839 ( .A(n15948), .ZN(n15934) );
  AOI21_X1 U13840 ( .B1(n15931), .B2(n14828), .A(n15354), .ZN(n11984) );
  NAND2_X1 U13841 ( .A1(n11984), .A2(n12021), .ZN(n15958) );
  INV_X1 U13842 ( .A(n7189), .ZN(n12628) );
  AND2_X1 U13843 ( .A1(n11986), .A2(n11985), .ZN(n11987) );
  NOR2_X1 U13844 ( .A1(n12011), .A2(n11987), .ZN(n12429) );
  NAND2_X1 U13845 ( .A1(n12628), .A2(n12429), .ZN(n11993) );
  OR2_X1 U13846 ( .A1(n14928), .A2(n15978), .ZN(n11992) );
  INV_X1 U13847 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11988) );
  OR2_X1 U13848 ( .A1(n12686), .A2(n11988), .ZN(n11991) );
  OR2_X1 U13849 ( .A1(n12705), .A2(n11989), .ZN(n11990) );
  NAND4_X1 U13850 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n15041) );
  AOI22_X1 U13851 ( .A1(n15342), .A2(n15041), .B1(n15043), .B2(n15289), .ZN(
        n15957) );
  OAI22_X1 U13852 ( .A1(n15957), .A2(n15946), .B1(n12238), .B2(n15755), .ZN(
        n11995) );
  NOR2_X1 U13853 ( .A1(n7606), .A2(n15317), .ZN(n11994) );
  AOI211_X1 U13854 ( .C1(n15946), .C2(P1_REG2_REG_13__SCAN_IN), .A(n11995), 
        .B(n11994), .ZN(n11996) );
  OAI21_X1 U13855 ( .B1(n15358), .B2(n15958), .A(n11996), .ZN(n12003) );
  NAND2_X1 U13856 ( .A1(n11998), .A2(n11997), .ZN(n15935) );
  NAND2_X1 U13857 ( .A1(n15935), .A2(n15928), .ZN(n15938) );
  INV_X1 U13858 ( .A(n15043), .ZN(n12237) );
  OR2_X1 U13859 ( .A1(n15948), .A2(n12237), .ZN(n11999) );
  NAND2_X1 U13860 ( .A1(n15938), .A2(n11999), .ZN(n12001) );
  INV_X1 U13861 ( .A(n14964), .ZN(n12000) );
  NOR2_X1 U13862 ( .A1(n12001), .A2(n12000), .ZN(n15961) );
  NAND2_X1 U13863 ( .A1(n12001), .A2(n12000), .ZN(n12010) );
  INV_X1 U13864 ( .A(n12010), .ZN(n15960) );
  NOR3_X1 U13865 ( .A1(n15961), .A2(n15960), .A3(n15337), .ZN(n12002) );
  AOI211_X1 U13866 ( .C1(n15964), .C2(n15952), .A(n12003), .B(n12002), .ZN(
        n12004) );
  INV_X1 U13867 ( .A(n12004), .ZN(P1_U3280) );
  NAND2_X1 U13868 ( .A1(n12005), .A2(n14944), .ZN(n12008) );
  AOI22_X1 U13869 ( .A1(n12597), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n12006), 
        .B2(n7182), .ZN(n12007) );
  XNOR2_X1 U13870 ( .A(n15967), .B(n15041), .ZN(n14966) );
  OR2_X1 U13871 ( .A1(n14828), .A2(n12268), .ZN(n12009) );
  XOR2_X1 U13872 ( .A(n14966), .B(n12195), .Z(n15977) );
  INV_X1 U13873 ( .A(n15977), .ZN(n12034) );
  INV_X1 U13874 ( .A(n12268), .ZN(n15042) );
  OR2_X1 U13875 ( .A1(n12011), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12012) );
  AND2_X1 U13876 ( .A1(n12012), .A2(n12183), .ZN(n14744) );
  NAND2_X1 U13877 ( .A1(n12628), .A2(n14744), .ZN(n12018) );
  INV_X1 U13878 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n12013) );
  OR2_X1 U13879 ( .A1(n12686), .A2(n12013), .ZN(n12017) );
  INV_X1 U13880 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n12014) );
  OR2_X1 U13881 ( .A1(n14928), .A2(n12014), .ZN(n12016) );
  INV_X1 U13882 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12190) );
  OR2_X1 U13883 ( .A1(n12705), .A2(n12190), .ZN(n12015) );
  NAND4_X1 U13884 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n15040) );
  AOI22_X1 U13885 ( .A1(n15042), .A2(n15289), .B1(n15342), .B2(n15040), .ZN(
        n15968) );
  INV_X1 U13886 ( .A(n15968), .ZN(n12019) );
  AOI22_X1 U13887 ( .A1(n12019), .A2(n15760), .B1(n12429), .B2(n15944), .ZN(
        n12020) );
  OAI21_X1 U13888 ( .B1(n11989), .B2(n15760), .A(n12020), .ZN(n12025) );
  NAND2_X1 U13889 ( .A1(n15967), .A2(n12021), .ZN(n12022) );
  NAND2_X1 U13890 ( .A1(n12022), .A2(n15932), .ZN(n12023) );
  OR2_X1 U13891 ( .A1(n12191), .A2(n12023), .ZN(n15969) );
  NOR2_X1 U13892 ( .A1(n15969), .A2(n15358), .ZN(n12024) );
  AOI211_X1 U13893 ( .C1(n15947), .C2(n15967), .A(n12025), .B(n12024), .ZN(
        n12033) );
  OR2_X1 U13894 ( .A1(n14828), .A2(n15042), .ZN(n12027) );
  NAND2_X1 U13895 ( .A1(n12028), .A2(n12027), .ZN(n12031) );
  INV_X1 U13896 ( .A(n12031), .ZN(n12030) );
  NAND2_X1 U13897 ( .A1(n12031), .A2(n14966), .ZN(n15972) );
  NAND3_X1 U13898 ( .A1(n15974), .A2(n15972), .A3(n15952), .ZN(n12032) );
  OAI211_X1 U13899 ( .C1(n12034), .C2(n15337), .A(n12033), .B(n12032), .ZN(
        P1_U3279) );
  OAI22_X1 U13900 ( .A1(n15806), .A2(n12928), .B1(n12035), .B2(n15804), .ZN(
        n12038) );
  MUX2_X1 U13901 ( .A(n12036), .B(P3_REG2_REG_7__SCAN_IN), .S(n15802), .Z(
        n12037) );
  AOI211_X1 U13902 ( .C1(n13820), .C2(n12039), .A(n12038), .B(n12037), .ZN(
        n12040) );
  INV_X1 U13903 ( .A(n12040), .ZN(P3_U3226) );
  NAND2_X1 U13904 ( .A1(n12938), .A2(n12939), .ZN(n12941) );
  XNOR2_X1 U13905 ( .A(n12041), .B(n12941), .ZN(n12043) );
  OAI22_X1 U13906 ( .A1(n12379), .A2(n13835), .B1(n12892), .B2(n13833), .ZN(
        n12042) );
  AOI21_X1 U13907 ( .B1(n12043), .B2(n13756), .A(n12042), .ZN(n15869) );
  INV_X1 U13908 ( .A(n12941), .ZN(n13063) );
  XNOR2_X1 U13909 ( .A(n12044), .B(n13063), .ZN(n15864) );
  NOR2_X1 U13910 ( .A1(n15810), .A2(n12045), .ZN(n12047) );
  OAI22_X1 U13911 ( .A1(n15806), .A2(n12168), .B1(n12173), .B2(n15804), .ZN(
        n12046) );
  AOI211_X1 U13912 ( .C1(n15864), .C2(n13820), .A(n12047), .B(n12046), .ZN(
        n12048) );
  OAI21_X1 U13913 ( .B1(n15869), .B2(n15802), .A(n12048), .ZN(P3_U3224) );
  AOI21_X1 U13914 ( .B1(n12052), .B2(n12050), .A(n12049), .ZN(n12138) );
  AOI22_X1 U13915 ( .A1(n14070), .A2(n14355), .B1(n14353), .B2(n14071), .ZN(
        n12055) );
  OAI211_X1 U13916 ( .C1(n12053), .C2(n12052), .A(n12051), .B(n14358), .ZN(
        n12054) );
  OAI211_X1 U13917 ( .C1(n12138), .C2(n10019), .A(n12055), .B(n12054), .ZN(
        n12056) );
  INV_X1 U13918 ( .A(n12056), .ZN(n12137) );
  INV_X1 U13919 ( .A(n12057), .ZN(n12058) );
  AOI21_X1 U13920 ( .B1(n12134), .B2(n12059), .A(n12058), .ZN(n12135) );
  AOI22_X1 U13921 ( .A1(n14347), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n12060), 
        .B2(n14345), .ZN(n12061) );
  OAI21_X1 U13922 ( .B1(n12062), .B2(n14349), .A(n12061), .ZN(n12064) );
  NOR2_X1 U13923 ( .A1(n12138), .A2(n14231), .ZN(n12063) );
  AOI211_X1 U13924 ( .C1(n12135), .C2(n14362), .A(n12064), .B(n12063), .ZN(
        n12065) );
  OAI21_X1 U13925 ( .B1(n14359), .B2(n12137), .A(n12065), .ZN(P2_U3252) );
  OR2_X1 U13926 ( .A1(n12066), .A2(n12175), .ZN(n12071) );
  INV_X1 U13927 ( .A(n12071), .ZN(n12068) );
  INV_X1 U13928 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12748) );
  MUX2_X1 U13929 ( .A(n12748), .B(P1_REG2_REG_16__SCAN_IN), .S(n12205), .Z(
        n12067) );
  OAI21_X1 U13930 ( .B1(n12068), .B2(n12069), .A(n12067), .ZN(n12072) );
  AOI21_X1 U13931 ( .B1(n12755), .B2(n12748), .A(n12069), .ZN(n12070) );
  OAI211_X1 U13932 ( .C1(n12755), .C2(n12748), .A(n12071), .B(n12070), .ZN(
        n12747) );
  NAND3_X1 U13933 ( .A1(n12072), .A2(n15730), .A3(n12747), .ZN(n12081) );
  NAND2_X1 U13934 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14664)
         );
  XOR2_X1 U13935 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n12205), .Z(n12077) );
  AOI21_X1 U13936 ( .B1(n12075), .B2(n12074), .A(n12073), .ZN(n12076) );
  NAND2_X1 U13937 ( .A1(n12076), .A2(n12077), .ZN(n12753) );
  OAI211_X1 U13938 ( .C1(n12077), .C2(n12076), .A(n15739), .B(n12753), .ZN(
        n12078) );
  NAND2_X1 U13939 ( .A1(n14664), .A2(n12078), .ZN(n12079) );
  AOI21_X1 U13940 ( .B1(n15732), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n12079), 
        .ZN(n12080) );
  OAI211_X1 U13941 ( .C1(n12771), .C2(n12755), .A(n12081), .B(n12080), .ZN(
        P1_U3259) );
  XOR2_X1 U13942 ( .A(n12083), .B(n12082), .Z(n12084) );
  NAND2_X1 U13943 ( .A1(n12084), .A2(n13241), .ZN(n12089) );
  OAI22_X1 U13944 ( .A1(n13255), .A2(n12891), .B1(n12085), .B2(n13247), .ZN(
        n12086) );
  AOI211_X1 U13945 ( .C1(n13245), .C2(n7681), .A(n12087), .B(n12086), .ZN(
        n12088) );
  OAI211_X1 U13946 ( .C1(n12090), .C2(n13200), .A(n12089), .B(n12088), .ZN(
        P3_U3161) );
  INV_X1 U13947 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n12092) );
  NOR2_X1 U13948 ( .A1(n12367), .A2(n12092), .ZN(n12091) );
  AOI21_X1 U13949 ( .B1(n12367), .B2(n12092), .A(n12091), .ZN(n12097) );
  OAI21_X1 U13950 ( .B1(n12100), .B2(P2_REG2_REG_11__SCAN_IN), .A(n12093), 
        .ZN(n12094) );
  XNOR2_X1 U13951 ( .A(n12094), .B(n15574), .ZN(n15577) );
  INV_X1 U13952 ( .A(n12094), .ZN(n12095) );
  AOI211_X1 U13953 ( .C1(n12097), .C2(n12096), .A(n15592), .B(n12366), .ZN(
        n12111) );
  INV_X1 U13954 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n12140) );
  NOR2_X1 U13955 ( .A1(n12367), .A2(n12140), .ZN(n12098) );
  AOI21_X1 U13956 ( .B1(n12140), .B2(n12367), .A(n12098), .ZN(n12105) );
  NOR2_X1 U13957 ( .A1(n15574), .A2(n12102), .ZN(n12101) );
  AOI21_X1 U13958 ( .B1(n12102), .B2(n15574), .A(n12101), .ZN(n15580) );
  OAI21_X1 U13959 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n12103), .A(n15578), 
        .ZN(n12104) );
  NOR2_X1 U13960 ( .A1(n12104), .A2(n12105), .ZN(n12362) );
  AOI211_X1 U13961 ( .C1(n12105), .C2(n12104), .A(n15588), .B(n12362), .ZN(
        n12110) );
  NAND2_X1 U13962 ( .A1(n15522), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n12107) );
  OAI211_X1 U13963 ( .C1(n14148), .C2(n12108), .A(n12107), .B(n12106), .ZN(
        n12109) );
  OR3_X1 U13964 ( .A1(n12111), .A2(n12110), .A3(n12109), .ZN(P2_U3227) );
  INV_X1 U13965 ( .A(n12119), .ZN(n12113) );
  NAND2_X1 U13966 ( .A1(n12113), .A2(n12112), .ZN(n12114) );
  NAND2_X1 U13967 ( .A1(n12115), .A2(n12114), .ZN(n12117) );
  XNOR2_X1 U13968 ( .A(n14444), .B(n12116), .ZN(n13116) );
  NAND2_X1 U13969 ( .A1(n14069), .A2(n12832), .ZN(n12439) );
  XNOR2_X1 U13970 ( .A(n13116), .B(n12439), .ZN(n12120) );
  AOI22_X1 U13971 ( .A1(n13142), .A2(n14354), .B1(n14047), .B2(n14070), .ZN(
        n12118) );
  NAND2_X1 U13972 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14091)
         );
  OAI211_X1 U13973 ( .C1(n12402), .C2(n14030), .A(n12118), .B(n14091), .ZN(
        n12124) );
  INV_X1 U13974 ( .A(n12115), .ZN(n12122) );
  AOI22_X1 U13975 ( .A1(n12119), .A2(n14054), .B1(n13994), .B2(n14070), .ZN(
        n12121) );
  NOR3_X1 U13976 ( .A1(n12122), .A2(n12121), .A3(n12120), .ZN(n12123) );
  AOI211_X1 U13977 ( .C1(n14444), .C2(n14035), .A(n12124), .B(n12123), .ZN(
        n12125) );
  OAI21_X1 U13978 ( .B1(n12441), .B2(n10844), .A(n12125), .ZN(P2_U3213) );
  INV_X1 U13979 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U13980 ( .A1(n12127), .A2(n14445), .B1(n15841), .B2(n12126), .ZN(
        n12128) );
  OAI211_X1 U13981 ( .C1(n12130), .C2(n14442), .A(n12129), .B(n12128), .ZN(
        n12132) );
  NAND2_X1 U13982 ( .A1(n12132), .A2(n14451), .ZN(n12131) );
  OAI21_X1 U13983 ( .B1(n14451), .B2(n12361), .A(n12131), .ZN(P2_U3513) );
  NAND2_X1 U13984 ( .A1(n12132), .A2(n14469), .ZN(n12133) );
  OAI21_X1 U13985 ( .B1(n14469), .B2(n8960), .A(n12133), .ZN(P2_U3472) );
  AOI22_X1 U13986 ( .A1(n12135), .A2(n14445), .B1(n15841), .B2(n12134), .ZN(
        n12136) );
  OAI211_X1 U13987 ( .C1(n12138), .C2(n14449), .A(n12137), .B(n12136), .ZN(
        n12141) );
  NAND2_X1 U13988 ( .A1(n12141), .A2(n14451), .ZN(n12139) );
  OAI21_X1 U13989 ( .B1(n14451), .B2(n12140), .A(n12139), .ZN(P2_U3512) );
  INV_X1 U13990 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n12143) );
  NAND2_X1 U13991 ( .A1(n12141), .A2(n14469), .ZN(n12142) );
  OAI21_X1 U13992 ( .B1(n14469), .B2(n12143), .A(n12142), .ZN(P2_U3469) );
  OAI222_X1 U13993 ( .A1(n13150), .A2(n12146), .B1(P2_U3088), .B2(n12145), 
        .C1(n14477), .C2(n12144), .ZN(P2_U3305) );
  INV_X1 U13994 ( .A(n12147), .ZN(n12148) );
  AOI21_X1 U13995 ( .B1(n15769), .B2(n12154), .A(n12148), .ZN(n12156) );
  OAI22_X1 U13996 ( .A1(n13960), .A2(n12891), .B1(n16000), .B2(n8241), .ZN(
        n12149) );
  AOI21_X1 U13997 ( .B1(n12154), .B2(n15771), .A(n12149), .ZN(n12150) );
  OAI21_X1 U13998 ( .B1(n12156), .B2(n16008), .A(n12150), .ZN(P3_U3414) );
  INV_X1 U13999 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12151) );
  OAI22_X1 U14000 ( .A1(n13905), .A2(n12891), .B1(n15997), .B2(n12151), .ZN(
        n12152) );
  AOI21_X1 U14001 ( .B1(n12154), .B2(n12153), .A(n12152), .ZN(n12155) );
  OAI21_X1 U14002 ( .B1(n12156), .B2(n16004), .A(n12155), .ZN(P3_U3467) );
  INV_X1 U14003 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12655) );
  INV_X1 U14004 ( .A(n12654), .ZN(n12159) );
  OAI222_X1 U14005 ( .A1(n15476), .A2(n12655), .B1(n13160), .B2(n12159), .C1(
        n12157), .C2(P1_U3086), .ZN(P1_U3331) );
  OAI222_X1 U14006 ( .A1(n13150), .A2(n12160), .B1(n14477), .B2(n12159), .C1(
        n12158), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U14007 ( .A(n12669), .ZN(n12164) );
  OAI222_X1 U14008 ( .A1(n13150), .A2(n12162), .B1(n14477), .B2(n12164), .C1(
        n12161), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U14009 ( .A1(n15476), .A2(n12670), .B1(n13160), .B2(n12164), .C1(
        n12163), .C2(P1_U3086), .ZN(P1_U3330) );
  OAI21_X1 U14010 ( .B1(n12166), .B2(n12165), .A(n12244), .ZN(n12167) );
  NAND2_X1 U14011 ( .A1(n12167), .A2(n13241), .ZN(n12172) );
  OAI22_X1 U14012 ( .A1(n13255), .A2(n12168), .B1(n12892), .B2(n13247), .ZN(
        n12169) );
  AOI211_X1 U14013 ( .C1(n13245), .C2(n13479), .A(n12170), .B(n12169), .ZN(
        n12171) );
  OAI211_X1 U14014 ( .C1(n12173), .C2(n13200), .A(n12172), .B(n12171), .ZN(
        P3_U3171) );
  NAND2_X1 U14015 ( .A1(n12174), .A2(n14944), .ZN(n12177) );
  AOI22_X1 U14016 ( .A1(n12597), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n12596), 
        .B2(n12175), .ZN(n12176) );
  NAND2_X1 U14017 ( .A1(n15982), .A2(n15040), .ZN(n12178) );
  NAND2_X1 U14018 ( .A1(n12346), .A2(n12178), .ZN(n12209) );
  NAND2_X1 U14019 ( .A1(n15967), .A2(n15041), .ZN(n12179) );
  INV_X1 U14020 ( .A(n12354), .ZN(n12180) );
  AOI21_X1 U14021 ( .B1(n12209), .B2(n12181), .A(n12180), .ZN(n15986) );
  NAND2_X1 U14022 ( .A1(n12183), .A2(n12182), .ZN(n12184) );
  AND2_X1 U14023 ( .A1(n12215), .A2(n12184), .ZN(n14668) );
  NAND2_X1 U14024 ( .A1(n14668), .A2(n12628), .ZN(n12188) );
  NAND2_X1 U14025 ( .A1(n14924), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n12187) );
  NAND2_X1 U14026 ( .A1(n14923), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12186) );
  NAND2_X1 U14027 ( .A1(n12711), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n12185) );
  INV_X1 U14028 ( .A(n15041), .ZN(n14742) );
  OAI22_X1 U14029 ( .A1(n14748), .A2(n15195), .B1(n14742), .B2(n15345), .ZN(
        n15980) );
  AOI22_X1 U14030 ( .A1(n15980), .A2(n15760), .B1(n14744), .B2(n15944), .ZN(
        n12189) );
  OAI21_X1 U14031 ( .B1(n12190), .B2(n15760), .A(n12189), .ZN(n12193) );
  INV_X1 U14032 ( .A(n15982), .ZN(n14489) );
  NAND2_X1 U14033 ( .A1(n12191), .A2(n14489), .ZN(n12212) );
  OAI211_X1 U14034 ( .C1(n14489), .C2(n12191), .A(n15932), .B(n12212), .ZN(
        n15983) );
  NOR2_X1 U14035 ( .A1(n15983), .A2(n15358), .ZN(n12192) );
  AOI211_X1 U14036 ( .C1(n15947), .C2(n15982), .A(n12193), .B(n12192), .ZN(
        n12199) );
  NAND2_X1 U14037 ( .A1(n15967), .A2(n14742), .ZN(n12194) );
  NAND2_X1 U14038 ( .A1(n12195), .A2(n12194), .ZN(n12197) );
  OR2_X1 U14039 ( .A1(n15967), .A2(n14742), .ZN(n12196) );
  NAND2_X1 U14040 ( .A1(n12197), .A2(n12196), .ZN(n12210) );
  INV_X1 U14041 ( .A(n12209), .ZN(n14965) );
  XNOR2_X1 U14042 ( .A(n12210), .B(n14965), .ZN(n15989) );
  NAND2_X1 U14043 ( .A1(n15989), .A2(n12224), .ZN(n12198) );
  OAI211_X1 U14044 ( .C1(n15986), .C2(n15285), .A(n12199), .B(n12198), .ZN(
        P1_U3278) );
  NAND2_X1 U14045 ( .A1(n12650), .A2(n15481), .ZN(n12200) );
  OAI211_X1 U14046 ( .C1(n10568), .C2(n15476), .A(n12200), .B(n15013), .ZN(
        P1_U3332) );
  NAND2_X1 U14047 ( .A1(n12650), .A2(n12201), .ZN(n12203) );
  OAI211_X1 U14048 ( .C1(n10754), .C2(n13150), .A(n12203), .B(n12202), .ZN(
        P2_U3304) );
  NAND2_X1 U14049 ( .A1(n12354), .A2(n12346), .ZN(n12208) );
  NAND2_X1 U14050 ( .A1(n12204), .A2(n14944), .ZN(n12207) );
  AOI22_X1 U14051 ( .A1(n12597), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12596), 
        .B2(n12205), .ZN(n12206) );
  XNOR2_X1 U14052 ( .A(n14845), .B(n14748), .ZN(n12349) );
  INV_X1 U14053 ( .A(n12349), .ZN(n14967) );
  XNOR2_X1 U14054 ( .A(n12208), .B(n14967), .ZN(n15455) );
  INV_X1 U14055 ( .A(n15040), .ZN(n14488) );
  OR2_X1 U14056 ( .A1(n15982), .A2(n14488), .ZN(n12211) );
  XNOR2_X1 U14057 ( .A(n12327), .B(n12349), .ZN(n15453) );
  INV_X1 U14058 ( .A(n14845), .ZN(n15451) );
  INV_X1 U14059 ( .A(n12212), .ZN(n12213) );
  OAI211_X1 U14060 ( .C1(n15451), .C2(n12213), .A(n15932), .B(n12335), .ZN(
        n15450) );
  AND2_X1 U14061 ( .A1(n12215), .A2(n12214), .ZN(n12216) );
  OR2_X1 U14062 ( .A1(n12216), .A2(n12337), .ZN(n14675) );
  AOI22_X1 U14063 ( .A1(n12711), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n14924), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n12218) );
  INV_X1 U14064 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12344) );
  OR2_X1 U14065 ( .A1(n12705), .A2(n12344), .ZN(n12217) );
  OAI211_X1 U14066 ( .C1(n14675), .C2(n7189), .A(n12218), .B(n12217), .ZN(
        n15038) );
  AOI22_X1 U14067 ( .A1(n15038), .A2(n15342), .B1(n15289), .B2(n15040), .ZN(
        n15449) );
  INV_X1 U14068 ( .A(n14668), .ZN(n12219) );
  OAI22_X1 U14069 ( .A1(n15449), .A2(n15946), .B1(n12219), .B2(n15755), .ZN(
        n12221) );
  NOR2_X1 U14070 ( .A1(n15451), .A2(n15317), .ZN(n12220) );
  AOI211_X1 U14071 ( .C1(n15946), .C2(P1_REG2_REG_16__SCAN_IN), .A(n12221), 
        .B(n12220), .ZN(n12222) );
  OAI21_X1 U14072 ( .B1(n15358), .B2(n15450), .A(n12222), .ZN(n12223) );
  AOI21_X1 U14073 ( .B1(n15453), .B2(n12224), .A(n12223), .ZN(n12225) );
  OAI21_X1 U14074 ( .B1(n15455), .B2(n15285), .A(n12225), .ZN(P1_U3277) );
  AND2_X1 U14075 ( .A1(n15043), .A2(n14563), .ZN(n12226) );
  AOI21_X1 U14076 ( .B1(n15948), .B2(n14587), .A(n12226), .ZN(n12231) );
  INV_X1 U14077 ( .A(n12231), .ZN(n12233) );
  OAI22_X1 U14078 ( .A1(n15934), .A2(n14627), .B1(n12237), .B2(n14572), .ZN(
        n12227) );
  XNOR2_X1 U14079 ( .A(n12227), .B(n14628), .ZN(n12232) );
  XOR2_X1 U14080 ( .A(n12231), .B(n12232), .Z(n12276) );
  AOI22_X1 U14081 ( .A1(n14828), .A2(n14581), .B1(n14587), .B2(n15042), .ZN(
        n12234) );
  XNOR2_X1 U14082 ( .A(n12234), .B(n14628), .ZN(n12423) );
  NOR2_X1 U14083 ( .A1(n12268), .A2(n14626), .ZN(n12235) );
  AOI21_X1 U14084 ( .B1(n14828), .B2(n14587), .A(n12235), .ZN(n12424) );
  XNOR2_X1 U14085 ( .A(n12423), .B(n12424), .ZN(n12425) );
  XNOR2_X1 U14086 ( .A(n12426), .B(n12425), .ZN(n12242) );
  OAI21_X1 U14087 ( .B1(n14743), .B2(n12237), .A(n12236), .ZN(n12240) );
  OAI22_X1 U14088 ( .A1(n14742), .A2(n14747), .B1(n14746), .B2(n12238), .ZN(
        n12239) );
  AOI211_X1 U14089 ( .C1(n14828), .C2(n14751), .A(n12240), .B(n12239), .ZN(
        n12241) );
  OAI21_X1 U14090 ( .B1(n12242), .B2(n14753), .A(n12241), .ZN(P1_U3234) );
  AND2_X1 U14091 ( .A1(n12244), .A2(n12243), .ZN(n12247) );
  OAI211_X1 U14092 ( .C1(n12247), .C2(n12246), .A(n13241), .B(n12245), .ZN(
        n12253) );
  NAND2_X1 U14093 ( .A1(n13245), .A2(n13266), .ZN(n12251) );
  NAND2_X1 U14094 ( .A1(n13198), .A2(n7681), .ZN(n12250) );
  NAND2_X1 U14095 ( .A1(n13218), .A2(n12248), .ZN(n12249) );
  OR2_X1 U14096 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13448), .ZN(n15699) );
  AND4_X1 U14097 ( .A1(n12251), .A2(n12250), .A3(n12249), .A4(n15699), .ZN(
        n12252) );
  OAI211_X1 U14098 ( .C1(n12260), .C2(n13200), .A(n12253), .B(n12252), .ZN(
        P3_U3157) );
  XNOR2_X1 U14099 ( .A(n12254), .B(n13062), .ZN(n15884) );
  XNOR2_X1 U14100 ( .A(n12255), .B(n13062), .ZN(n12258) );
  OAI22_X1 U14101 ( .A1(n12256), .A2(n13833), .B1(n12552), .B2(n13835), .ZN(
        n12257) );
  AOI21_X1 U14102 ( .B1(n12258), .B2(n13756), .A(n12257), .ZN(n12259) );
  OAI21_X1 U14103 ( .B1(n13880), .B2(n15884), .A(n12259), .ZN(n15886) );
  NAND2_X1 U14104 ( .A1(n15886), .A2(n15810), .ZN(n12263) );
  OAI22_X1 U14105 ( .A1(n15806), .A2(n15885), .B1(n12260), .B2(n15804), .ZN(
        n12261) );
  AOI21_X1 U14106 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n15802), .A(n12261), 
        .ZN(n12262) );
  OAI211_X1 U14107 ( .C1(n15884), .C2(n13702), .A(n12263), .B(n12262), .ZN(
        P3_U3223) );
  INV_X1 U14108 ( .A(n12264), .ZN(n12265) );
  OAI222_X1 U14109 ( .A1(n12267), .A2(P3_U3151), .B1(n13969), .B2(n12266), 
        .C1(n13157), .C2(n12265), .ZN(P3_U3270) );
  OR2_X1 U14110 ( .A1(n12268), .A2(n15195), .ZN(n12271) );
  OR2_X1 U14111 ( .A1(n12269), .A2(n15345), .ZN(n12270) );
  NAND2_X1 U14112 ( .A1(n12271), .A2(n12270), .ZN(n15937) );
  NAND2_X1 U14113 ( .A1(n15937), .A2(n14694), .ZN(n12273) );
  OAI211_X1 U14114 ( .C1(n14746), .C2(n15943), .A(n12273), .B(n12272), .ZN(
        n12278) );
  AOI211_X1 U14115 ( .C1(n12276), .C2(n12275), .A(n14753), .B(n12274), .ZN(
        n12277) );
  AOI211_X1 U14116 ( .C1(n14751), .C2(n15948), .A(n12278), .B(n12277), .ZN(
        n12279) );
  INV_X1 U14117 ( .A(n12279), .ZN(P1_U3224) );
  INV_X1 U14118 ( .A(n12280), .ZN(n12282) );
  NAND2_X1 U14119 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12302), .ZN(n12283) );
  OAI21_X1 U14120 ( .B1(n12302), .B2(P3_REG1_REG_12__SCAN_IN), .A(n12283), 
        .ZN(n15715) );
  NAND2_X1 U14121 ( .A1(P3_REG1_REG_14__SCAN_IN), .A2(n13517), .ZN(n12287) );
  OAI21_X1 U14122 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n13517), .A(n12287), 
        .ZN(n12288) );
  AOI21_X1 U14123 ( .B1(n12289), .B2(n12288), .A(n13507), .ZN(n12316) );
  INV_X1 U14124 ( .A(n13517), .ZN(n12311) );
  INV_X1 U14125 ( .A(n15702), .ZN(n13577) );
  NAND2_X1 U14126 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n12484)
         );
  OAI21_X1 U14127 ( .B1(n13577), .B2(n9888), .A(n12484), .ZN(n12301) );
  MUX2_X1 U14128 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13087), .Z(n13518) );
  XNOR2_X1 U14129 ( .A(n13518), .B(n13517), .ZN(n12299) );
  MUX2_X1 U14130 ( .A(n12526), .B(n12290), .S(n13087), .Z(n12296) );
  INV_X1 U14131 ( .A(n12296), .ZN(n12297) );
  MUX2_X1 U14132 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13087), .Z(n12295) );
  INV_X1 U14133 ( .A(n12302), .ZN(n15703) );
  XNOR2_X1 U14134 ( .A(n12295), .B(n15703), .ZN(n15706) );
  AOI22_X1 U14135 ( .A1(n15705), .A2(n15706), .B1(n12295), .B2(n12302), .ZN(
        n13494) );
  XNOR2_X1 U14136 ( .A(n12296), .B(n13501), .ZN(n13493) );
  NAND2_X1 U14137 ( .A1(n13494), .A2(n13493), .ZN(n13492) );
  OAI21_X1 U14138 ( .B1(n12297), .B2(n13501), .A(n13492), .ZN(n12298) );
  NOR2_X1 U14139 ( .A1(n12298), .A2(n12299), .ZN(n13516) );
  AOI211_X1 U14140 ( .C1(n12299), .C2(n12298), .A(n15681), .B(n13516), .ZN(
        n12300) );
  AOI211_X1 U14141 ( .C1(n15704), .C2(n12311), .A(n12301), .B(n12300), .ZN(
        n12315) );
  NAND2_X1 U14142 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n12302), .ZN(n12307) );
  AOI22_X1 U14143 ( .A1(n15703), .A2(n12559), .B1(P3_REG2_REG_12__SCAN_IN), 
        .B2(n12302), .ZN(n15709) );
  NAND2_X1 U14144 ( .A1(n12304), .A2(n12303), .ZN(n12306) );
  NAND2_X1 U14145 ( .A1(n12306), .A2(n12305), .ZN(n15708) );
  NAND2_X1 U14146 ( .A1(n12308), .A2(n13501), .ZN(n12309) );
  NAND2_X1 U14147 ( .A1(n12311), .A2(n12310), .ZN(n13511) );
  OAI21_X1 U14148 ( .B1(n12311), .B2(n12310), .A(n13511), .ZN(n12313) );
  AOI21_X1 U14149 ( .B1(n13510), .B2(n12313), .A(n15677), .ZN(n12312) );
  OAI21_X1 U14150 ( .B1(n13510), .B2(n12313), .A(n12312), .ZN(n12314) );
  OAI211_X1 U14151 ( .C1(n12316), .C2(n15718), .A(n12315), .B(n12314), .ZN(
        P3_U3196) );
  XNOR2_X1 U14152 ( .A(n12318), .B(n12317), .ZN(n12326) );
  INV_X1 U14153 ( .A(n12383), .ZN(n12319) );
  NAND2_X1 U14154 ( .A1(n13250), .A2(n12319), .ZN(n12322) );
  AOI21_X1 U14155 ( .B1(n13245), .B2(n13264), .A(n12320), .ZN(n12321) );
  OAI211_X1 U14156 ( .C1(n12379), .C2(n13247), .A(n12322), .B(n12321), .ZN(
        n12323) );
  AOI21_X1 U14157 ( .B1(n12324), .B2(n13218), .A(n12323), .ZN(n12325) );
  OAI21_X1 U14158 ( .B1(n12326), .B2(n13222), .A(n12325), .ZN(P3_U3176) );
  NAND2_X1 U14159 ( .A1(n14845), .A2(n14748), .ZN(n12328) );
  NAND2_X1 U14160 ( .A1(n12329), .A2(n12328), .ZN(n12333) );
  NAND2_X1 U14161 ( .A1(n12330), .A2(n14944), .ZN(n12332) );
  AOI22_X1 U14162 ( .A1(n12597), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7182), 
        .B2(n12757), .ZN(n12331) );
  NAND2_X2 U14163 ( .A1(n12332), .A2(n12331), .ZN(n15445) );
  OAI21_X1 U14164 ( .B1(n12333), .B2(n14968), .A(n12590), .ZN(n12334) );
  INV_X1 U14165 ( .A(n12334), .ZN(n15448) );
  AOI21_X1 U14166 ( .B1(n15445), .B2(n12335), .A(n15354), .ZN(n12336) );
  AND2_X1 U14167 ( .A1(n12336), .A2(n15355), .ZN(n15443) );
  NAND2_X1 U14168 ( .A1(n15445), .A2(n15947), .ZN(n12343) );
  NOR2_X1 U14169 ( .A1(n12337), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n12338) );
  OR2_X1 U14170 ( .A1(n12600), .A2(n12338), .ZN(n15352) );
  AOI22_X1 U14171 ( .A1(n12711), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n14924), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n12340) );
  NAND2_X1 U14172 ( .A1(n14923), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n12339) );
  OAI211_X1 U14173 ( .C1(n15352), .C2(n7189), .A(n12340), .B(n12339), .ZN(
        n15037) );
  INV_X1 U14174 ( .A(n15037), .ZN(n14676) );
  OAI22_X1 U14175 ( .A1(n14676), .A2(n15195), .B1(n14748), .B2(n15345), .ZN(
        n15444) );
  INV_X1 U14176 ( .A(n14675), .ZN(n12341) );
  AOI22_X1 U14177 ( .A1(n15444), .A2(n15760), .B1(n12341), .B2(n15944), .ZN(
        n12342) );
  OAI211_X1 U14178 ( .C1(n15760), .C2(n12344), .A(n12343), .B(n12342), .ZN(
        n12345) );
  AOI21_X1 U14179 ( .B1(n15443), .B2(n15951), .A(n12345), .ZN(n12359) );
  INV_X1 U14180 ( .A(n14748), .ZN(n15039) );
  OR2_X1 U14181 ( .A1(n14845), .A2(n15039), .ZN(n12348) );
  AND2_X1 U14182 ( .A1(n12346), .A2(n12348), .ZN(n12353) );
  INV_X1 U14183 ( .A(n14968), .ZN(n12347) );
  AND2_X1 U14184 ( .A1(n12353), .A2(n12347), .ZN(n12352) );
  INV_X1 U14185 ( .A(n12348), .ZN(n12350) );
  OR2_X1 U14186 ( .A1(n12350), .A2(n12349), .ZN(n12355) );
  OR2_X1 U14187 ( .A1(n14968), .A2(n12355), .ZN(n12351) );
  NAND2_X1 U14188 ( .A1(n12354), .A2(n12353), .ZN(n12356) );
  AND2_X1 U14189 ( .A1(n12356), .A2(n12355), .ZN(n12357) );
  NAND2_X1 U14190 ( .A1(n12357), .A2(n14968), .ZN(n15442) );
  NAND3_X1 U14191 ( .A1(n12720), .A2(n15442), .A3(n15952), .ZN(n12358) );
  OAI211_X1 U14192 ( .C1(n15448), .C2(n15337), .A(n12359), .B(n12358), .ZN(
        P1_U3276) );
  NOR2_X1 U14193 ( .A1(n14084), .A2(n12361), .ZN(n12360) );
  AOI21_X1 U14194 ( .B1(n12361), .B2(n14084), .A(n12360), .ZN(n12364) );
  AOI211_X1 U14195 ( .C1(n12364), .C2(n12363), .A(n15588), .B(n14083), .ZN(
        n12365) );
  INV_X1 U14196 ( .A(n12365), .ZN(n12375) );
  NOR2_X1 U14197 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14084), .ZN(n14087) );
  INV_X1 U14198 ( .A(n14087), .ZN(n12368) );
  NAND2_X1 U14199 ( .A1(n14084), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14088) );
  NAND2_X1 U14200 ( .A1(n12368), .A2(n14088), .ZN(n12370) );
  OAI21_X1 U14201 ( .B1(n14089), .B2(n12370), .A(n15583), .ZN(n12369) );
  AOI21_X1 U14202 ( .B1(n14089), .B2(n12370), .A(n12369), .ZN(n12373) );
  INV_X1 U14203 ( .A(n12371), .ZN(n12372) );
  AOI211_X1 U14204 ( .C1(n15522), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n12373), 
        .B(n12372), .ZN(n12374) );
  OAI211_X1 U14205 ( .C1(n14148), .C2(n12376), .A(n12375), .B(n12374), .ZN(
        P2_U3228) );
  XNOR2_X1 U14206 ( .A(n12377), .B(n13061), .ZN(n12378) );
  OAI222_X1 U14207 ( .A1(n13835), .A2(n12380), .B1(n13833), .B2(n12379), .C1(
        n12378), .C2(n13831), .ZN(n15914) );
  INV_X1 U14208 ( .A(n15914), .ZN(n12388) );
  OAI21_X1 U14209 ( .B1(n12382), .B2(n13061), .A(n12381), .ZN(n15916) );
  NOR2_X1 U14210 ( .A1(n15806), .A2(n15913), .ZN(n12386) );
  OAI22_X1 U14211 ( .A1(n15810), .A2(n12384), .B1(n12383), .B2(n15804), .ZN(
        n12385) );
  AOI211_X1 U14212 ( .C1(n15916), .C2(n13820), .A(n12386), .B(n12385), .ZN(
        n12387) );
  OAI21_X1 U14213 ( .B1(n12388), .B2(n15802), .A(n12387), .ZN(P3_U3222) );
  INV_X1 U14214 ( .A(n12681), .ZN(n12390) );
  OAI222_X1 U14215 ( .A1(n10281), .A2(P1_U3086), .B1(n13160), .B2(n12390), 
        .C1(n12682), .C2(n15476), .ZN(P1_U3329) );
  OAI222_X1 U14216 ( .A1(n12391), .A2(P2_U3088), .B1(n14477), .B2(n12390), 
        .C1(n12389), .C2(n13150), .ZN(P2_U3301) );
  XOR2_X1 U14217 ( .A(n12392), .B(n12396), .Z(n12399) );
  OAI22_X1 U14218 ( .A1(n12394), .A2(n14322), .B1(n12393), .B2(n14320), .ZN(
        n12398) );
  AOI21_X1 U14219 ( .B1(n12396), .B2(n12395), .A(n7276), .ZN(n14450) );
  NOR2_X1 U14220 ( .A1(n14450), .A2(n10019), .ZN(n12397) );
  AOI211_X1 U14221 ( .C1(n12399), .C2(n14358), .A(n12398), .B(n12397), .ZN(
        n14448) );
  INV_X1 U14222 ( .A(n12470), .ZN(n12400) );
  AOI21_X1 U14223 ( .B1(n14444), .B2(n12401), .A(n12400), .ZN(n14446) );
  INV_X1 U14224 ( .A(n12402), .ZN(n12403) );
  AOI22_X1 U14225 ( .A1(n14347), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12403), 
        .B2(n14345), .ZN(n12404) );
  OAI21_X1 U14226 ( .B1(n9406), .B2(n14349), .A(n12404), .ZN(n12406) );
  NOR2_X1 U14227 ( .A1(n14450), .A2(n14231), .ZN(n12405) );
  AOI211_X1 U14228 ( .C1(n14446), .C2(n14362), .A(n12406), .B(n12405), .ZN(
        n12407) );
  OAI21_X1 U14229 ( .B1(n14448), .B2(n14359), .A(n12407), .ZN(P2_U3250) );
  NAND2_X1 U14230 ( .A1(n7993), .A2(n12409), .ZN(n12410) );
  XNOR2_X1 U14231 ( .A(n12411), .B(n12410), .ZN(n12416) );
  NAND2_X1 U14232 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n15720)
         );
  OAI21_X1 U14233 ( .B1(n13236), .B2(n12957), .A(n15720), .ZN(n12412) );
  AOI21_X1 U14234 ( .B1(n13198), .B2(n13266), .A(n12412), .ZN(n12413) );
  OAI21_X1 U14235 ( .B1(n13200), .B2(n12560), .A(n12413), .ZN(n12414) );
  AOI21_X1 U14236 ( .B1(n12566), .B2(n13218), .A(n12414), .ZN(n12415) );
  OAI21_X1 U14237 ( .B1(n12416), .B2(n13222), .A(n12415), .ZN(P3_U3164) );
  NAND2_X1 U14238 ( .A1(n15967), .A2(n14581), .ZN(n12418) );
  NAND2_X1 U14239 ( .A1(n15041), .A2(n14587), .ZN(n12417) );
  NAND2_X1 U14240 ( .A1(n12418), .A2(n12417), .ZN(n12419) );
  XNOR2_X1 U14241 ( .A(n12419), .B(n14584), .ZN(n12422) );
  AND2_X1 U14242 ( .A1(n15041), .A2(n14563), .ZN(n12420) );
  AOI21_X1 U14243 ( .B1(n15967), .B2(n14587), .A(n12420), .ZN(n12421) );
  NAND2_X1 U14244 ( .A1(n12422), .A2(n12421), .ZN(n14484) );
  OAI21_X1 U14245 ( .B1(n12422), .B2(n12421), .A(n14484), .ZN(n12428) );
  AOI21_X1 U14246 ( .B1(n12428), .B2(n12427), .A(n7339), .ZN(n12434) );
  NAND2_X1 U14247 ( .A1(n14667), .A2(n12429), .ZN(n12430) );
  OAI211_X1 U14248 ( .C1(n15968), .C2(n14665), .A(n12431), .B(n12430), .ZN(
        n12432) );
  AOI21_X1 U14249 ( .B1(n15967), .B2(n14751), .A(n12432), .ZN(n12433) );
  OAI21_X1 U14250 ( .B1(n12434), .B2(n14753), .A(n12433), .ZN(P1_U3215) );
  XNOR2_X1 U14251 ( .A(n14428), .B(n12804), .ZN(n12435) );
  AND2_X1 U14252 ( .A1(n14356), .A2(n12832), .ZN(n12436) );
  NAND2_X1 U14253 ( .A1(n12435), .A2(n12436), .ZN(n12499) );
  INV_X1 U14254 ( .A(n12435), .ZN(n12739) );
  INV_X1 U14255 ( .A(n12436), .ZN(n12437) );
  NAND2_X1 U14256 ( .A1(n12739), .A2(n12437), .ZN(n12438) );
  NAND2_X1 U14257 ( .A1(n12499), .A2(n12438), .ZN(n12450) );
  INV_X1 U14258 ( .A(n13116), .ZN(n12440) );
  XNOR2_X1 U14259 ( .A(n14438), .B(n12116), .ZN(n13106) );
  NAND2_X1 U14260 ( .A1(n14354), .A2(n12832), .ZN(n12442) );
  XNOR2_X1 U14261 ( .A(n13106), .B(n12442), .ZN(n13117) );
  INV_X1 U14262 ( .A(n13106), .ZN(n12443) );
  XNOR2_X1 U14263 ( .A(n14433), .B(n12116), .ZN(n12445) );
  NAND2_X1 U14264 ( .A1(n14068), .A2(n12832), .ZN(n12446) );
  XNOR2_X1 U14265 ( .A(n12445), .B(n12446), .ZN(n13107) );
  NAND2_X1 U14266 ( .A1(n12444), .A2(n13107), .ZN(n13113) );
  INV_X1 U14267 ( .A(n12445), .ZN(n12447) );
  NAND2_X1 U14268 ( .A1(n12447), .A2(n12446), .ZN(n12448) );
  NAND2_X1 U14269 ( .A1(n13113), .A2(n12448), .ZN(n12449) );
  AOI21_X1 U14270 ( .B1(n12450), .B2(n12449), .A(n10844), .ZN(n12453) );
  INV_X1 U14271 ( .A(n12449), .ZN(n12452) );
  NAND2_X1 U14272 ( .A1(n12453), .A2(n12737), .ZN(n12456) );
  AND2_X1 U14273 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14131) );
  OAI22_X1 U14274 ( .A1(n9224), .A2(n14050), .B1(n14031), .B2(n14321), .ZN(
        n12454) );
  AOI211_X1 U14275 ( .C1(n14046), .C2(n14330), .A(n14131), .B(n12454), .ZN(
        n12455) );
  OAI211_X1 U14276 ( .C1(n14333), .C2(n14044), .A(n12456), .B(n12455), .ZN(
        P2_U3210) );
  OAI211_X1 U14277 ( .C1(n12459), .C2(n12458), .A(n12457), .B(n13241), .ZN(
        n12465) );
  INV_X1 U14278 ( .A(n12958), .ZN(n12528) );
  INV_X1 U14279 ( .A(n12460), .ZN(n12527) );
  NAND2_X1 U14280 ( .A1(n13250), .A2(n12527), .ZN(n12462) );
  INV_X1 U14281 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n13468) );
  NOR2_X1 U14282 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13468), .ZN(n13499) );
  AOI21_X1 U14283 ( .B1(n13198), .B2(n13264), .A(n13499), .ZN(n12461) );
  OAI211_X1 U14284 ( .C1(n13248), .C2(n13236), .A(n12462), .B(n12461), .ZN(
        n12463) );
  AOI21_X1 U14285 ( .B1(n12528), .B2(n13218), .A(n12463), .ZN(n12464) );
  NAND2_X1 U14286 ( .A1(n12465), .A2(n12464), .ZN(P3_U3174) );
  INV_X1 U14287 ( .A(n12466), .ZN(n12467) );
  OAI222_X1 U14288 ( .A1(n13157), .A2(n12467), .B1(n13087), .B2(P3_U3151), 
        .C1(n13385), .C2(n13983), .ZN(P3_U3268) );
  XOR2_X1 U14289 ( .A(n12468), .B(n12475), .Z(n12469) );
  AOI222_X1 U14290 ( .A1(n14358), .A2(n12469), .B1(n14068), .B2(n14355), .C1(
        n14069), .C2(n14353), .ZN(n14441) );
  AOI21_X1 U14291 ( .B1(n14438), .B2(n12470), .A(n14340), .ZN(n14439) );
  INV_X1 U14292 ( .A(n13115), .ZN(n12471) );
  AOI22_X1 U14293 ( .A1(n14347), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12471), 
        .B2(n14345), .ZN(n12472) );
  OAI21_X1 U14294 ( .B1(n12473), .B2(n14349), .A(n12472), .ZN(n12478) );
  OAI21_X1 U14295 ( .B1(n12476), .B2(n12475), .A(n12474), .ZN(n14443) );
  NOR2_X1 U14296 ( .A1(n14443), .A2(n14364), .ZN(n12477) );
  AOI211_X1 U14297 ( .C1(n14439), .C2(n14362), .A(n12478), .B(n12477), .ZN(
        n12479) );
  OAI21_X1 U14298 ( .B1(n14347), .B2(n14441), .A(n12479), .ZN(P2_U3249) );
  OAI211_X1 U14299 ( .C1(n12482), .C2(n12481), .A(n12480), .B(n13241), .ZN(
        n12488) );
  INV_X1 U14300 ( .A(n12483), .ZN(n12494) );
  NAND2_X1 U14301 ( .A1(n13245), .A2(n13262), .ZN(n12485) );
  OAI211_X1 U14302 ( .C1(n12957), .C2(n13247), .A(n12485), .B(n12484), .ZN(
        n12486) );
  AOI21_X1 U14303 ( .B1(n12494), .B2(n13250), .A(n12486), .ZN(n12487) );
  OAI211_X1 U14304 ( .C1(n13255), .C2(n13913), .A(n12488), .B(n12487), .ZN(
        P3_U3155) );
  INV_X1 U14305 ( .A(n12586), .ZN(n12736) );
  OAI222_X1 U14306 ( .A1(n13150), .A2(n12490), .B1(n14477), .B2(n12736), .C1(
        P2_U3088), .C2(n12489), .ZN(P2_U3300) );
  XNOR2_X1 U14307 ( .A(n12491), .B(n7664), .ZN(n12492) );
  AOI222_X1 U14308 ( .A1(n13756), .A2(n12492), .B1(n9776), .B2(n13759), .C1(
        n13262), .C2(n13742), .ZN(n13912) );
  XNOR2_X1 U14309 ( .A(n12493), .B(n7664), .ZN(n13910) );
  AOI22_X1 U14310 ( .A1(n15802), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n13802), 
        .B2(n12494), .ZN(n12495) );
  OAI21_X1 U14311 ( .B1(n13913), .B2(n15806), .A(n12495), .ZN(n12496) );
  AOI21_X1 U14312 ( .B1(n13910), .B2(n13820), .A(n12496), .ZN(n12497) );
  OAI21_X1 U14313 ( .B1(n13912), .B2(n15802), .A(n12497), .ZN(P3_U3219) );
  AND2_X1 U14314 ( .A1(n14067), .A2(n12832), .ZN(n12498) );
  NAND2_X1 U14315 ( .A1(n12500), .A2(n12498), .ZN(n12502) );
  OAI21_X1 U14316 ( .B1(n12500), .B2(n12498), .A(n12502), .ZN(n12738) );
  NOR2_X1 U14317 ( .A1(n14038), .A2(n9224), .ZN(n12501) );
  AOI22_X1 U14318 ( .A1(n12746), .A2(n14054), .B1(n12501), .B2(n12500), .ZN(
        n12511) );
  NAND2_X1 U14319 ( .A1(n14066), .A2(n12832), .ZN(n12806) );
  XNOR2_X1 U14320 ( .A(n14418), .B(n12804), .ZN(n12805) );
  XOR2_X1 U14321 ( .A(n12806), .B(n12805), .Z(n12503) );
  INV_X1 U14322 ( .A(n12503), .ZN(n12510) );
  INV_X1 U14323 ( .A(n12502), .ZN(n12504) );
  OAI22_X1 U14324 ( .A1(n12505), .A2(n14322), .B1(n9224), .B2(n14320), .ZN(
        n14280) );
  AOI22_X1 U14325 ( .A1(n14280), .A2(n14023), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12507) );
  NAND2_X1 U14326 ( .A1(n14046), .A2(n14287), .ZN(n12506) );
  OAI211_X1 U14327 ( .C1(n14290), .C2(n14044), .A(n12507), .B(n12506), .ZN(
        n12508) );
  AOI21_X1 U14328 ( .B1(n12808), .B2(n14054), .A(n12508), .ZN(n12509) );
  OAI21_X1 U14329 ( .B1(n12511), .B2(n12510), .A(n12509), .ZN(P2_U3205) );
  INV_X1 U14330 ( .A(n12698), .ZN(n12579) );
  AOI21_X1 U14331 ( .B1(n14475), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n12512), 
        .ZN(n12513) );
  OAI21_X1 U14332 ( .B1(n12579), .B2(n14477), .A(n12513), .ZN(P2_U3299) );
  XNOR2_X1 U14333 ( .A(n12514), .B(n13065), .ZN(n12519) );
  INV_X1 U14334 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12520) );
  XNOR2_X1 U14335 ( .A(n12515), .B(n13065), .ZN(n12517) );
  AOI22_X1 U14336 ( .A1(n13264), .A2(n13759), .B1(n13263), .B2(n13742), .ZN(
        n12516) );
  OAI21_X1 U14337 ( .B1(n12517), .B2(n13831), .A(n12516), .ZN(n12518) );
  AOI21_X1 U14338 ( .B1(n12519), .B2(n15769), .A(n12518), .ZN(n12525) );
  MUX2_X1 U14339 ( .A(n12520), .B(n12525), .S(n16000), .Z(n12522) );
  INV_X1 U14340 ( .A(n13960), .ZN(n16009) );
  NAND2_X1 U14341 ( .A1(n16009), .A2(n12528), .ZN(n12521) );
  OAI211_X1 U14342 ( .C1(n12531), .C2(n13946), .A(n12522), .B(n12521), .ZN(
        P3_U3429) );
  MUX2_X1 U14343 ( .A(n12290), .B(n12525), .S(n15997), .Z(n12524) );
  NAND2_X1 U14344 ( .A1(n16005), .A2(n12528), .ZN(n12523) );
  OAI211_X1 U14345 ( .C1(n12531), .C2(n13885), .A(n12524), .B(n12523), .ZN(
        P3_U3472) );
  MUX2_X1 U14346 ( .A(n12526), .B(n12525), .S(n15810), .Z(n12530) );
  AOI22_X1 U14347 ( .A1(n13816), .A2(n12528), .B1(n13802), .B2(n12527), .ZN(
        n12529) );
  OAI211_X1 U14348 ( .C1(n12531), .C2(n13702), .A(n12530), .B(n12529), .ZN(
        P3_U3220) );
  XNOR2_X1 U14349 ( .A(n12532), .B(n13070), .ZN(n12533) );
  AOI222_X1 U14350 ( .A1(n13756), .A2(n12533), .B1(n13263), .B2(n13759), .C1(
        n13261), .C2(n13742), .ZN(n13909) );
  XNOR2_X1 U14351 ( .A(n12534), .B(n13070), .ZN(n13907) );
  INV_X1 U14352 ( .A(n12535), .ZN(n13251) );
  AOI22_X1 U14353 ( .A1(n15802), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n13802), 
        .B2(n13251), .ZN(n12536) );
  OAI21_X1 U14354 ( .B1(n13254), .B2(n15806), .A(n12536), .ZN(n12537) );
  AOI21_X1 U14355 ( .B1(n13907), .B2(n13820), .A(n12537), .ZN(n12538) );
  OAI21_X1 U14356 ( .B1(n13909), .B2(n15802), .A(n12538), .ZN(P3_U3218) );
  XNOR2_X1 U14357 ( .A(n12539), .B(n13260), .ZN(n12540) );
  XNOR2_X1 U14358 ( .A(n12541), .B(n12540), .ZN(n12546) );
  INV_X1 U14359 ( .A(n13900), .ZN(n13817) );
  NAND2_X1 U14360 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13555)
         );
  OAI21_X1 U14361 ( .B1(n13236), .B2(n13808), .A(n13555), .ZN(n12542) );
  AOI21_X1 U14362 ( .B1(n13198), .B2(n13261), .A(n12542), .ZN(n12543) );
  OAI21_X1 U14363 ( .B1(n13200), .B2(n13813), .A(n12543), .ZN(n12544) );
  AOI21_X1 U14364 ( .B1(n13817), .B2(n13218), .A(n12544), .ZN(n12545) );
  OAI21_X1 U14365 ( .B1(n12546), .B2(n13222), .A(n12545), .ZN(P3_U3168) );
  INV_X1 U14366 ( .A(n14945), .ZN(n13154) );
  OAI222_X1 U14367 ( .A1(n14477), .A2(n13154), .B1(P2_U3088), .B2(n12548), 
        .C1(n12547), .C2(n13150), .ZN(P2_U3298) );
  INV_X1 U14368 ( .A(n12549), .ZN(n13066) );
  XNOR2_X1 U14369 ( .A(n12550), .B(n13066), .ZN(n12569) );
  INV_X1 U14370 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12556) );
  XNOR2_X1 U14371 ( .A(n12551), .B(n13066), .ZN(n12555) );
  OAI22_X1 U14372 ( .A1(n12552), .A2(n13833), .B1(n12957), .B2(n13835), .ZN(
        n12554) );
  NOR2_X1 U14373 ( .A1(n12569), .A2(n13880), .ZN(n12553) );
  AOI211_X1 U14374 ( .C1(n13756), .C2(n12555), .A(n12554), .B(n12553), .ZN(
        n12564) );
  MUX2_X1 U14375 ( .A(n12556), .B(n12564), .S(n15997), .Z(n12558) );
  NAND2_X1 U14376 ( .A1(n16005), .A2(n12566), .ZN(n12557) );
  OAI211_X1 U14377 ( .C1(n12569), .C2(n13885), .A(n12558), .B(n12557), .ZN(
        P3_U3471) );
  MUX2_X1 U14378 ( .A(n12559), .B(n12564), .S(n15810), .Z(n12563) );
  INV_X1 U14379 ( .A(n12560), .ZN(n12561) );
  AOI22_X1 U14380 ( .A1(n13816), .A2(n12566), .B1(n13802), .B2(n12561), .ZN(
        n12562) );
  OAI211_X1 U14381 ( .C1(n12569), .C2(n13702), .A(n12563), .B(n12562), .ZN(
        P3_U3221) );
  MUX2_X1 U14382 ( .A(n12565), .B(n12564), .S(n16000), .Z(n12568) );
  NAND2_X1 U14383 ( .A1(n16009), .A2(n12566), .ZN(n12567) );
  OAI211_X1 U14384 ( .C1(n12569), .C2(n13946), .A(n12568), .B(n12567), .ZN(
        P3_U3426) );
  XNOR2_X1 U14385 ( .A(n12570), .B(n12571), .ZN(n12577) );
  NAND2_X1 U14386 ( .A1(n13198), .A2(n13260), .ZN(n12572) );
  NAND2_X1 U14387 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13575)
         );
  OAI211_X1 U14388 ( .C1(n13800), .C2(n13236), .A(n12572), .B(n13575), .ZN(
        n12575) );
  INV_X1 U14389 ( .A(n12573), .ZN(n13955) );
  NOR2_X1 U14390 ( .A1(n13955), .A2(n13255), .ZN(n12574) );
  AOI211_X1 U14391 ( .C1(n13801), .C2(n13250), .A(n12575), .B(n12574), .ZN(
        n12576) );
  OAI21_X1 U14392 ( .B1(n12577), .B2(n13222), .A(n12576), .ZN(P3_U3178) );
  AND2_X1 U14393 ( .A1(n12578), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U14394 ( .A1(n12578), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U14395 ( .A1(n12578), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U14396 ( .A1(n12578), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U14397 ( .A1(n12578), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U14398 ( .A1(n12578), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U14399 ( .A1(n12578), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U14400 ( .A1(n12578), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U14401 ( .A1(n12578), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U14402 ( .A1(n12578), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U14403 ( .A1(n12578), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U14404 ( .A1(n12578), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U14405 ( .A1(n12578), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U14406 ( .A1(n12578), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U14407 ( .A1(n12578), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U14408 ( .A1(n12578), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U14409 ( .A1(n12578), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U14410 ( .A1(n12578), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U14411 ( .A1(n12578), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U14412 ( .A1(n12578), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U14413 ( .A1(n12578), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U14414 ( .A1(n12578), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U14415 ( .A1(n12578), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U14416 ( .A1(n12578), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U14417 ( .A1(n12578), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U14418 ( .A1(n12578), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U14419 ( .A1(n12578), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U14420 ( .A1(n12578), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U14421 ( .A1(n12578), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U14422 ( .A1(n12578), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  OAI222_X1 U14423 ( .A1(n15476), .A2(n7845), .B1(n13160), .B2(n12579), .C1(
        n7409), .C2(P1_U3086), .ZN(P1_U3327) );
  NAND2_X1 U14424 ( .A1(n12711), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n12585) );
  INV_X1 U14425 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n12580) );
  OR2_X1 U14426 ( .A1(n12686), .A2(n12580), .ZN(n12584) );
  INV_X1 U14427 ( .A(n12660), .ZN(n12581) );
  NAND2_X1 U14428 ( .A1(n12687), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n12702) );
  OAI21_X1 U14429 ( .B1(n12687), .B2(P1_REG3_REG_27__SCAN_IN), .A(n12702), 
        .ZN(n15200) );
  OR2_X1 U14430 ( .A1(n7189), .A2(n15200), .ZN(n12583) );
  INV_X1 U14431 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n15201) );
  OR2_X1 U14432 ( .A1(n12705), .A2(n15201), .ZN(n12582) );
  NAND2_X1 U14433 ( .A1(n12586), .A2(n14944), .ZN(n12588) );
  OR2_X1 U14434 ( .A1(n14947), .A2(n7848), .ZN(n12587) );
  INV_X1 U14435 ( .A(n15038), .ZN(n15346) );
  NAND2_X1 U14436 ( .A1(n15445), .A2(n15346), .ZN(n12589) );
  NAND2_X1 U14437 ( .A1(n12591), .A2(n14944), .ZN(n12593) );
  AOI22_X1 U14438 ( .A1(n12597), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7182), 
        .B2(n15129), .ZN(n12592) );
  XNOR2_X1 U14439 ( .A(n15436), .B(n14676), .ZN(n15340) );
  NAND2_X1 U14440 ( .A1(n12595), .A2(n14944), .ZN(n12599) );
  AOI22_X1 U14441 ( .A1(n12597), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n12596), 
        .B2(n15140), .ZN(n12598) );
  NOR2_X1 U14442 ( .A1(n12600), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n12601) );
  OR2_X1 U14443 ( .A1(n12612), .A2(n12601), .ZN(n15329) );
  INV_X1 U14444 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15125) );
  NAND2_X1 U14445 ( .A1(n14924), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n12603) );
  NAND2_X1 U14446 ( .A1(n14923), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n12602) );
  OAI211_X1 U14447 ( .C1(n14928), .C2(n15125), .A(n12603), .B(n12602), .ZN(
        n12604) );
  INV_X1 U14448 ( .A(n12604), .ZN(n12605) );
  XNOR2_X1 U14449 ( .A(n15333), .B(n15343), .ZN(n15324) );
  NAND2_X1 U14450 ( .A1(n15333), .A2(n7974), .ZN(n12606) );
  NAND2_X1 U14451 ( .A1(n12608), .A2(n14944), .ZN(n12611) );
  OR2_X1 U14452 ( .A1(n14947), .A2(n12609), .ZN(n12610) );
  NOR2_X1 U14453 ( .A1(n12612), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n12613) );
  OR2_X1 U14454 ( .A1(n12625), .A2(n12613), .ZN(n15313) );
  INV_X1 U14455 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n12616) );
  NAND2_X1 U14456 ( .A1(n14923), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n12615) );
  NAND2_X1 U14457 ( .A1(n14924), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n12614) );
  OAI211_X1 U14458 ( .C1(n14928), .C2(n12616), .A(n12615), .B(n12614), .ZN(
        n12617) );
  INV_X1 U14459 ( .A(n12617), .ZN(n12618) );
  XNOR2_X1 U14460 ( .A(n15425), .B(n15290), .ZN(n12724) );
  INV_X1 U14461 ( .A(n15290), .ZN(n12619) );
  OR2_X1 U14462 ( .A1(n15425), .A2(n12619), .ZN(n12620) );
  NAND2_X1 U14463 ( .A1(n12621), .A2(n14944), .ZN(n12624) );
  OR2_X1 U14464 ( .A1(n14947), .A2(n12622), .ZN(n12623) );
  OR2_X1 U14465 ( .A1(n12625), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12627) );
  AND2_X1 U14466 ( .A1(n12627), .A2(n12626), .ZN(n15299) );
  NAND2_X1 U14467 ( .A1(n15299), .A2(n12628), .ZN(n12634) );
  INV_X1 U14468 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n12631) );
  NAND2_X1 U14469 ( .A1(n14923), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n12630) );
  NAND2_X1 U14470 ( .A1(n14924), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n12629) );
  OAI211_X1 U14471 ( .C1(n14928), .C2(n12631), .A(n12630), .B(n12629), .ZN(
        n12632) );
  INV_X1 U14472 ( .A(n12632), .ZN(n12633) );
  INV_X1 U14473 ( .A(n15295), .ZN(n12635) );
  NAND2_X1 U14474 ( .A1(n15288), .A2(n12635), .ZN(n12637) );
  OR2_X1 U14475 ( .A1(n15300), .A2(n14705), .ZN(n12636) );
  NAND2_X1 U14476 ( .A1(n12639), .A2(n12638), .ZN(n12640) );
  XNOR2_X1 U14477 ( .A(n12640), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15484) );
  NAND2_X1 U14478 ( .A1(n15484), .A2(n12641), .ZN(n14880) );
  NAND2_X1 U14479 ( .A1(n12711), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12648) );
  INV_X1 U14480 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n12642) );
  OR2_X1 U14481 ( .A1(n12686), .A2(n12642), .ZN(n12647) );
  OAI21_X1 U14482 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n12644), .A(n12643), 
        .ZN(n15278) );
  OR2_X1 U14483 ( .A1(n7189), .A2(n15278), .ZN(n12646) );
  INV_X1 U14484 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n15279) );
  OR2_X1 U14485 ( .A1(n12705), .A2(n15279), .ZN(n12645) );
  NAND4_X1 U14486 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n15291) );
  XNOR2_X1 U14487 ( .A(n14880), .B(n15291), .ZN(n15275) );
  OR2_X1 U14488 ( .A1(n14880), .A2(n15291), .ZN(n12649) );
  NAND2_X1 U14489 ( .A1(n12650), .A2(n14944), .ZN(n12652) );
  OR2_X1 U14490 ( .A1(n14947), .A2(n10568), .ZN(n12651) );
  NAND2_X2 U14491 ( .A1(n12652), .A2(n12651), .ZN(n15409) );
  XNOR2_X1 U14492 ( .A(n15409), .B(n15271), .ZN(n15262) );
  INV_X1 U14493 ( .A(n15271), .ZN(n14706) );
  NAND2_X1 U14494 ( .A1(n15409), .A2(n14706), .ZN(n12653) );
  NAND2_X1 U14495 ( .A1(n12654), .A2(n14944), .ZN(n12657) );
  OR2_X1 U14496 ( .A1(n14947), .A2(n12655), .ZN(n12656) );
  NAND2_X1 U14497 ( .A1(n14924), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n12666) );
  INV_X1 U14498 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n12658) );
  OR2_X1 U14499 ( .A1(n14928), .A2(n12658), .ZN(n12665) );
  INV_X1 U14500 ( .A(n12659), .ZN(n12675) );
  INV_X1 U14501 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n12661) );
  NAND2_X1 U14502 ( .A1(n12661), .A2(n12660), .ZN(n12662) );
  NAND2_X1 U14503 ( .A1(n12675), .A2(n12662), .ZN(n15247) );
  OR2_X1 U14504 ( .A1(n7189), .A2(n15247), .ZN(n12664) );
  INV_X1 U14505 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n15248) );
  OR2_X1 U14506 ( .A1(n12705), .A2(n15248), .ZN(n12663) );
  NAND4_X1 U14507 ( .A1(n12666), .A2(n12665), .A3(n12664), .A4(n12663), .ZN(
        n15036) );
  XNOR2_X1 U14508 ( .A(n15250), .B(n15036), .ZN(n15240) );
  INV_X1 U14509 ( .A(n15036), .ZN(n14599) );
  NAND2_X1 U14510 ( .A1(n12669), .A2(n14944), .ZN(n12672) );
  OR2_X1 U14511 ( .A1(n14947), .A2(n12670), .ZN(n12671) );
  NAND2_X1 U14512 ( .A1(n12711), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12680) );
  INV_X1 U14513 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n12673) );
  OR2_X1 U14514 ( .A1(n12686), .A2(n12673), .ZN(n12679) );
  INV_X1 U14515 ( .A(n12674), .ZN(n12688) );
  INV_X1 U14516 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14655) );
  NAND2_X1 U14517 ( .A1(n12675), .A2(n14655), .ZN(n12676) );
  NAND2_X1 U14518 ( .A1(n12688), .A2(n12676), .ZN(n15229) );
  INV_X1 U14519 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n15228) );
  OR2_X1 U14520 ( .A1(n12705), .A2(n15228), .ZN(n12677) );
  XNOR2_X1 U14521 ( .A(n15232), .B(n14733), .ZN(n15224) );
  NAND2_X1 U14522 ( .A1(n12681), .A2(n14944), .ZN(n12684) );
  OR2_X1 U14523 ( .A1(n14947), .A2(n12682), .ZN(n12683) );
  NAND2_X1 U14524 ( .A1(n12711), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12696) );
  INV_X1 U14525 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n12685) );
  OR2_X1 U14526 ( .A1(n12686), .A2(n12685), .ZN(n12695) );
  INV_X1 U14527 ( .A(n12687), .ZN(n12690) );
  INV_X1 U14528 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14732) );
  NAND2_X1 U14529 ( .A1(n12688), .A2(n14732), .ZN(n12689) );
  NAND2_X1 U14530 ( .A1(n12690), .A2(n12689), .ZN(n15210) );
  OR2_X1 U14531 ( .A1(n7189), .A2(n15210), .ZN(n12694) );
  INV_X1 U14532 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n12691) );
  OR2_X1 U14533 ( .A1(n12692), .A2(n12691), .ZN(n12693) );
  NAND2_X1 U14534 ( .A1(n15392), .A2(n15194), .ZN(n15190) );
  OR2_X1 U14535 ( .A1(n15392), .A2(n15194), .ZN(n12697) );
  NAND2_X1 U14536 ( .A1(n15190), .A2(n12697), .ZN(n15206) );
  INV_X1 U14537 ( .A(n15206), .ZN(n15216) );
  NAND2_X1 U14538 ( .A1(n15215), .A2(n15216), .ZN(n15214) );
  XNOR2_X1 U14539 ( .A(n15387), .B(n14734), .ZN(n15191) );
  AOI21_X1 U14540 ( .B1(n15214), .B2(n15190), .A(n15191), .ZN(n15189) );
  NAND2_X1 U14541 ( .A1(n12698), .A2(n14944), .ZN(n12700) );
  OR2_X1 U14542 ( .A1(n14947), .A2(n7845), .ZN(n12699) );
  NAND2_X1 U14543 ( .A1(n14924), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n12709) );
  INV_X1 U14544 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n12701) );
  OR2_X1 U14545 ( .A1(n14928), .A2(n12701), .ZN(n12708) );
  INV_X1 U14546 ( .A(n12702), .ZN(n12703) );
  NAND2_X1 U14547 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n12703), .ZN(n15166) );
  OAI21_X1 U14548 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n12703), .A(n15166), 
        .ZN(n14635) );
  OR2_X1 U14549 ( .A1(n7189), .A2(n14635), .ZN(n12707) );
  INV_X1 U14550 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n12731) );
  OR2_X1 U14551 ( .A1(n12705), .A2(n12731), .ZN(n12706) );
  NAND4_X1 U14552 ( .A1(n12709), .A2(n12708), .A3(n12707), .A4(n12706), .ZN(
        n15176) );
  XNOR2_X1 U14553 ( .A(n15378), .B(n15176), .ZN(n14975) );
  XNOR2_X1 U14554 ( .A(n15179), .B(n12710), .ZN(n12718) );
  NAND2_X1 U14555 ( .A1(n12711), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12715) );
  NAND2_X1 U14556 ( .A1(n14924), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12714) );
  OR2_X1 U14557 ( .A1(n7189), .A2(n15166), .ZN(n12713) );
  INV_X1 U14558 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n15170) );
  OR2_X1 U14559 ( .A1(n12705), .A2(n15170), .ZN(n12712) );
  NAND4_X1 U14560 ( .A1(n12715), .A2(n12714), .A3(n12713), .A4(n12712), .ZN(
        n15034) );
  NAND2_X1 U14561 ( .A1(n15034), .A2(n15342), .ZN(n12716) );
  NAND2_X1 U14562 ( .A1(n15445), .A2(n15038), .ZN(n12719) );
  OR2_X1 U14563 ( .A1(n15436), .A2(n15037), .ZN(n12721) );
  NAND2_X1 U14564 ( .A1(n15338), .A2(n12721), .ZN(n12723) );
  NAND2_X1 U14565 ( .A1(n15436), .A2(n15037), .ZN(n12722) );
  NAND2_X1 U14566 ( .A1(n15425), .A2(n15290), .ZN(n15293) );
  AND2_X1 U14567 ( .A1(n15295), .A2(n15293), .ZN(n12725) );
  OR2_X1 U14568 ( .A1(n15300), .A2(n15272), .ZN(n12726) );
  NAND2_X1 U14569 ( .A1(n15294), .A2(n12726), .ZN(n15276) );
  INV_X1 U14570 ( .A(n15291), .ZN(n14881) );
  NAND2_X1 U14571 ( .A1(n14880), .A2(n14881), .ZN(n12727) );
  NAND2_X1 U14572 ( .A1(n15409), .A2(n15271), .ZN(n12729) );
  OAI21_X1 U14573 ( .B1(n15398), .B2(n14733), .A(n15223), .ZN(n15207) );
  INV_X1 U14574 ( .A(n15194), .ZN(n15035) );
  NAND2_X1 U14575 ( .A1(n15188), .A2(n15191), .ZN(n15187) );
  OAI21_X1 U14576 ( .B1(n15217), .B2(n15387), .A(n15187), .ZN(n12730) );
  NOR2_X1 U14577 ( .A1(n12730), .A2(n14975), .ZN(n15161) );
  AOI21_X1 U14578 ( .B1(n14975), .B2(n12730), .A(n15161), .ZN(n15377) );
  INV_X1 U14579 ( .A(n15300), .ZN(n15298) );
  NAND2_X1 U14580 ( .A1(n15311), .A2(n15298), .ZN(n15297) );
  OAI211_X1 U14581 ( .C1(n7224), .C2(n15177), .A(n15932), .B(n15171), .ZN(
        n15380) );
  OAI22_X1 U14582 ( .A1(n15760), .A2(n12731), .B1(n14635), .B2(n15755), .ZN(
        n12732) );
  AOI21_X1 U14583 ( .B1(n15378), .B2(n15947), .A(n12732), .ZN(n12733) );
  OAI21_X1 U14584 ( .B1(n15380), .B2(n15358), .A(n12733), .ZN(n12734) );
  AOI21_X1 U14585 ( .B1(n15377), .B2(n15952), .A(n12734), .ZN(n12735) );
  OAI21_X1 U14586 ( .B1(n15384), .B2(n15946), .A(n12735), .ZN(P1_U3265) );
  OAI222_X1 U14587 ( .A1(n15476), .A2(n7848), .B1(n13160), .B2(n12736), .C1(
        P1_U3086), .C2(n7200), .ZN(P1_U3328) );
  AOI21_X1 U14588 ( .B1(n12738), .B2(n12737), .A(n10844), .ZN(n12741) );
  INV_X1 U14589 ( .A(n14356), .ZN(n14301) );
  NOR3_X1 U14590 ( .A1(n12739), .A2(n14301), .A3(n14038), .ZN(n12740) );
  NOR2_X1 U14591 ( .A1(n12741), .A2(n12740), .ZN(n12745) );
  AOI22_X1 U14592 ( .A1(n14047), .A2(n14356), .B1(n13142), .B2(n14066), .ZN(
        n12742) );
  NAND2_X1 U14593 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n14146)
         );
  OAI211_X1 U14594 ( .C1(n14030), .C2(n14309), .A(n12742), .B(n14146), .ZN(
        n12743) );
  AOI21_X1 U14595 ( .B1(n14424), .B2(n14035), .A(n12743), .ZN(n12744) );
  OAI21_X1 U14596 ( .B1(n12746), .B2(n12745), .A(n12744), .ZN(P2_U3191) );
  NAND2_X1 U14597 ( .A1(n12757), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n12752) );
  OAI21_X1 U14598 ( .B1(n12748), .B2(n12755), .A(n12747), .ZN(n12764) );
  OR2_X1 U14599 ( .A1(n12757), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U14600 ( .A1(n12749), .A2(n12752), .ZN(n12765) );
  INV_X1 U14601 ( .A(n12765), .ZN(n12750) );
  NAND2_X1 U14602 ( .A1(n12764), .A2(n12750), .ZN(n12751) );
  NAND2_X1 U14603 ( .A1(n12752), .A2(n12751), .ZN(n15130) );
  XNOR2_X1 U14604 ( .A(n15130), .B(n15129), .ZN(n15127) );
  INV_X1 U14605 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15353) );
  XNOR2_X1 U14606 ( .A(n15127), .B(n15353), .ZN(n12763) );
  NAND2_X1 U14607 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14719)
         );
  INV_X1 U14608 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n12754) );
  OAI21_X1 U14609 ( .B1(n12755), .B2(n12754), .A(n12753), .ZN(n12766) );
  INV_X1 U14610 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n12756) );
  XNOR2_X1 U14611 ( .A(n12757), .B(n12756), .ZN(n12767) );
  AOI22_X1 U14612 ( .A1(n12766), .A2(n12767), .B1(n12757), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n15121) );
  XNOR2_X1 U14613 ( .A(n15121), .B(n15129), .ZN(n12758) );
  NAND2_X1 U14614 ( .A1(n12758), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n15124) );
  OAI211_X1 U14615 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n12758), .A(n15739), 
        .B(n15124), .ZN(n12759) );
  NAND2_X1 U14616 ( .A1(n14719), .A2(n12759), .ZN(n12760) );
  AOI21_X1 U14617 ( .B1(n15732), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n12760), 
        .ZN(n12762) );
  NAND2_X1 U14618 ( .A1(n15741), .A2(n15129), .ZN(n12761) );
  OAI211_X1 U14619 ( .C1(n12763), .C2(n15087), .A(n12762), .B(n12761), .ZN(
        P1_U3261) );
  XOR2_X1 U14620 ( .A(n12765), .B(n12764), .Z(n12775) );
  NAND2_X1 U14621 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14674)
         );
  XOR2_X1 U14622 ( .A(n12767), .B(n12766), .Z(n12768) );
  NAND2_X1 U14623 ( .A1(n15739), .A2(n12768), .ZN(n12769) );
  NAND2_X1 U14624 ( .A1(n14674), .A2(n12769), .ZN(n12773) );
  NOR2_X1 U14625 ( .A1(n12771), .A2(n12770), .ZN(n12772) );
  AOI211_X1 U14626 ( .C1(n15732), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n12773), 
        .B(n12772), .ZN(n12774) );
  OAI21_X1 U14627 ( .B1(n12775), .B2(n15087), .A(n12774), .ZN(P1_U3260) );
  OAI21_X1 U14628 ( .B1(n12778), .B2(n12777), .A(n12776), .ZN(n12779) );
  NAND2_X1 U14629 ( .A1(n12779), .A2(n14716), .ZN(n12785) );
  INV_X1 U14630 ( .A(n15052), .ZN(n12781) );
  OAI22_X1 U14631 ( .A1(n12781), .A2(n14747), .B1(n14743), .B2(n12780), .ZN(
        n12782) );
  AOI21_X1 U14632 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n12783), .A(n12782), .ZN(
        n12784) );
  OAI211_X1 U14633 ( .C1(n15775), .C2(n14725), .A(n12785), .B(n12784), .ZN(
        P1_U3237) );
  INV_X1 U14634 ( .A(n12786), .ZN(n12791) );
  NAND2_X1 U14635 ( .A1(n12788), .A2(n14054), .ZN(n12789) );
  OAI21_X1 U14636 ( .B1(n12795), .B2(n14038), .A(n12789), .ZN(n12790) );
  NAND3_X1 U14637 ( .A1(n12791), .A2(n12787), .A3(n12790), .ZN(n12801) );
  NAND2_X1 U14638 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n15599)
         );
  INV_X1 U14639 ( .A(n15599), .ZN(n12792) );
  AOI21_X1 U14640 ( .B1(n14046), .B2(n12793), .A(n12792), .ZN(n12800) );
  OAI22_X1 U14641 ( .A1(n12795), .A2(n14031), .B1(n14050), .B2(n12794), .ZN(
        n12796) );
  INV_X1 U14642 ( .A(n12796), .ZN(n12799) );
  NAND2_X1 U14643 ( .A1(n12797), .A2(n14035), .ZN(n12798) );
  AND4_X1 U14644 ( .A1(n12801), .A2(n12800), .A3(n12799), .A4(n12798), .ZN(
        n12802) );
  OAI21_X1 U14645 ( .B1(n12803), .B2(n10844), .A(n12802), .ZN(P2_U3189) );
  XNOR2_X1 U14646 ( .A(n14413), .B(n12804), .ZN(n12809) );
  NAND2_X1 U14647 ( .A1(n14251), .A2(n12832), .ZN(n12810) );
  INV_X1 U14648 ( .A(n12805), .ZN(n12807) );
  XNOR2_X1 U14649 ( .A(n12809), .B(n12810), .ZN(n14007) );
  XNOR2_X1 U14650 ( .A(n14407), .B(n12116), .ZN(n12812) );
  XNOR2_X1 U14651 ( .A(n12813), .B(n12812), .ZN(n13095) );
  XNOR2_X1 U14652 ( .A(n14403), .B(n12116), .ZN(n12814) );
  NAND2_X1 U14653 ( .A1(n14252), .A2(n12832), .ZN(n13995) );
  INV_X1 U14654 ( .A(n12814), .ZN(n12815) );
  AND2_X1 U14655 ( .A1(n12816), .A2(n12815), .ZN(n12817) );
  XNOR2_X1 U14656 ( .A(n14396), .B(n7540), .ZN(n14014) );
  NAND2_X1 U14657 ( .A1(n14064), .A2(n12832), .ZN(n12819) );
  NOR2_X1 U14658 ( .A1(n14014), .A2(n12819), .ZN(n12820) );
  AOI21_X1 U14659 ( .B1(n14014), .B2(n12819), .A(n12820), .ZN(n14027) );
  INV_X1 U14660 ( .A(n12820), .ZN(n12821) );
  NAND2_X1 U14661 ( .A1(n14026), .A2(n12821), .ZN(n12827) );
  XNOR2_X1 U14662 ( .A(n14392), .B(n12116), .ZN(n12822) );
  AND2_X1 U14663 ( .A1(n14221), .A2(n12832), .ZN(n12823) );
  NAND2_X1 U14664 ( .A1(n12822), .A2(n12823), .ZN(n12828) );
  INV_X1 U14665 ( .A(n12822), .ZN(n14040) );
  INV_X1 U14666 ( .A(n12823), .ZN(n12824) );
  NAND2_X1 U14667 ( .A1(n14040), .A2(n12824), .ZN(n12825) );
  NAND2_X1 U14668 ( .A1(n12828), .A2(n12825), .ZN(n14015) );
  XNOR2_X1 U14669 ( .A(n14386), .B(n7540), .ZN(n12831) );
  NAND2_X1 U14670 ( .A1(n14063), .A2(n12832), .ZN(n12830) );
  XNOR2_X1 U14671 ( .A(n12831), .B(n12830), .ZN(n14043) );
  INV_X1 U14672 ( .A(n12828), .ZN(n12829) );
  XNOR2_X1 U14673 ( .A(n14377), .B(n7540), .ZN(n12834) );
  NAND2_X1 U14674 ( .A1(n14190), .A2(n12832), .ZN(n12833) );
  NOR2_X1 U14675 ( .A1(n12834), .A2(n12833), .ZN(n12835) );
  AOI21_X1 U14676 ( .B1(n12834), .B2(n12833), .A(n12835), .ZN(n13986) );
  MUX2_X1 U14677 ( .A(n14373), .B(n12836), .S(n12832), .Z(n12837) );
  XNOR2_X1 U14678 ( .A(n12837), .B(n12116), .ZN(n12838) );
  XNOR2_X1 U14679 ( .A(n12839), .B(n12838), .ZN(n12844) );
  AOI22_X1 U14680 ( .A1(n14190), .A2(n14353), .B1(n14061), .B2(n14355), .ZN(
        n14168) );
  INV_X1 U14681 ( .A(n14173), .ZN(n12840) );
  AOI22_X1 U14682 ( .A1(n12840), .A2(n14046), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12841) );
  OAI21_X1 U14683 ( .B1(n14168), .B2(n14002), .A(n12841), .ZN(n12842) );
  AOI21_X1 U14684 ( .B1(n14373), .B2(n14035), .A(n12842), .ZN(n12843) );
  OAI21_X1 U14685 ( .B1(n12844), .B2(n10844), .A(n12843), .ZN(P2_U3192) );
  INV_X1 U14686 ( .A(n12845), .ZN(n12848) );
  OAI22_X1 U14687 ( .A1(n14038), .A2(n12852), .B1(n12846), .B2(n10844), .ZN(
        n12847) );
  NAND3_X1 U14688 ( .A1(n12848), .A2(n11778), .A3(n12847), .ZN(n12858) );
  AOI21_X1 U14689 ( .B1(n14046), .B2(n12850), .A(n12849), .ZN(n12857) );
  OAI22_X1 U14690 ( .A1(n12852), .A2(n14031), .B1(n14050), .B2(n12851), .ZN(
        n12853) );
  INV_X1 U14691 ( .A(n12853), .ZN(n12856) );
  NAND2_X1 U14692 ( .A1(n14035), .A2(n12854), .ZN(n12855) );
  AND4_X1 U14693 ( .A1(n12858), .A2(n12857), .A3(n12856), .A4(n12855), .ZN(
        n12859) );
  OAI21_X1 U14694 ( .B1(n12787), .B2(n10844), .A(n12859), .ZN(P2_U3203) );
  INV_X1 U14695 ( .A(n12860), .ZN(n12865) );
  NAND2_X1 U14696 ( .A1(n12861), .A2(n14362), .ZN(n12864) );
  AOI22_X1 U14697 ( .A1(n12862), .A2(n14345), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14359), .ZN(n12863) );
  OAI211_X1 U14698 ( .C1(n12865), .C2(n14349), .A(n12864), .B(n12863), .ZN(
        n12866) );
  AOI21_X1 U14699 ( .B1(n12867), .B2(n14292), .A(n12866), .ZN(n12868) );
  OAI21_X1 U14700 ( .B1(n12869), .B2(n14359), .A(n12868), .ZN(P2_U3236) );
  INV_X1 U14701 ( .A(n12870), .ZN(n12871) );
  OAI222_X1 U14702 ( .A1(n12873), .A2(P3_U3151), .B1(n13983), .B2(n12872), 
        .C1(n13157), .C2(n12871), .ZN(P3_U3269) );
  AND2_X2 U14703 ( .A1(n12886), .A2(n12874), .ZN(n13693) );
  OAI21_X1 U14704 ( .B1(n13925), .B2(n13691), .A(n12876), .ZN(n12878) );
  NAND2_X1 U14705 ( .A1(n12878), .A2(n12877), .ZN(n12881) );
  INV_X1 U14706 ( .A(n12879), .ZN(n12880) );
  AOI21_X1 U14707 ( .B1(n12882), .B2(n12881), .A(n12880), .ZN(n12885) );
  AOI21_X1 U14708 ( .B1(n12887), .B2(n12883), .A(n13012), .ZN(n12888) );
  NOR3_X1 U14709 ( .A1(n12884), .A2(n12885), .A3(n12889), .ZN(n13007) );
  AOI21_X1 U14710 ( .B1(n12887), .B2(n12886), .A(n12885), .ZN(n12890) );
  MUX2_X1 U14711 ( .A(n12892), .B(n12891), .S(n13012), .Z(n12932) );
  INV_X1 U14712 ( .A(n12932), .ZN(n12937) );
  OAI21_X1 U14713 ( .B1(n12896), .B2(n12895), .A(n12894), .ZN(n12903) );
  NOR2_X1 U14714 ( .A1(n12901), .A2(n12900), .ZN(n12907) );
  AOI21_X1 U14715 ( .B1(n12903), .B2(n12902), .A(n13012), .ZN(n12906) );
  OAI21_X1 U14716 ( .B1(n12914), .B2(n12904), .A(n13012), .ZN(n12905) );
  OAI21_X1 U14717 ( .B1(n12909), .B2(n12908), .A(n12911), .ZN(n12910) );
  AOI22_X1 U14718 ( .A1(n12912), .A2(n12911), .B1(n13002), .B2(n12910), .ZN(
        n12913) );
  MUX2_X1 U14719 ( .A(n12916), .B(n12915), .S(n13012), .Z(n12917) );
  OAI211_X1 U14720 ( .C1(n12918), .C2(n13053), .A(n13055), .B(n12917), .ZN(
        n12922) );
  MUX2_X1 U14721 ( .A(n12920), .B(n12919), .S(n13012), .Z(n12921) );
  NAND3_X1 U14722 ( .A1(n12922), .A2(n13054), .A3(n12921), .ZN(n12927) );
  MUX2_X1 U14723 ( .A(n12924), .B(n12923), .S(n13012), .Z(n12925) );
  NAND3_X1 U14724 ( .A1(n12927), .A2(n12926), .A3(n12925), .ZN(n12934) );
  NAND2_X1 U14725 ( .A1(n13481), .A2(n12928), .ZN(n12930) );
  MUX2_X1 U14726 ( .A(n12930), .B(n12929), .S(n13012), .Z(n12933) );
  AOI22_X1 U14727 ( .A1(n12934), .A2(n12933), .B1(n12932), .B2(n12931), .ZN(
        n12935) );
  MUX2_X1 U14728 ( .A(n12939), .B(n12938), .S(n13012), .Z(n12940) );
  OAI211_X1 U14729 ( .C1(n12942), .C2(n12941), .A(n13062), .B(n12940), .ZN(
        n12946) );
  MUX2_X1 U14730 ( .A(n12944), .B(n12943), .S(n13002), .Z(n12945) );
  NAND3_X1 U14731 ( .A1(n12946), .A2(n13061), .A3(n12945), .ZN(n12951) );
  NAND3_X1 U14732 ( .A1(n12951), .A2(n12953), .A3(n12947), .ZN(n12949) );
  NAND2_X1 U14733 ( .A1(n12949), .A2(n12948), .ZN(n12956) );
  NAND2_X1 U14734 ( .A1(n12951), .A2(n12950), .ZN(n12954) );
  AOI21_X1 U14735 ( .B1(n12954), .B2(n12953), .A(n12952), .ZN(n12955) );
  NOR2_X1 U14736 ( .A1(n12957), .A2(n13002), .ZN(n12959) );
  OAI21_X1 U14737 ( .B1(n12962), .B2(n12961), .A(n12963), .ZN(n12964) );
  MUX2_X1 U14738 ( .A(n12964), .B(n12963), .S(n13012), .Z(n12965) );
  OAI211_X1 U14739 ( .C1(n12966), .C2(n13067), .A(n13070), .B(n12965), .ZN(
        n12975) );
  MUX2_X1 U14740 ( .A(n13261), .B(n13836), .S(n13012), .Z(n12971) );
  INV_X1 U14741 ( .A(n13254), .ZN(n13906) );
  NOR2_X1 U14742 ( .A1(n13906), .A2(n13832), .ZN(n12968) );
  MUX2_X1 U14743 ( .A(n12968), .B(n12967), .S(n13012), .Z(n12969) );
  AOI21_X1 U14744 ( .B1(n12970), .B2(n12971), .A(n12969), .ZN(n12974) );
  OAI21_X1 U14745 ( .B1(n12972), .B2(n12971), .A(n13818), .ZN(n12973) );
  INV_X1 U14746 ( .A(n12979), .ZN(n12978) );
  OAI211_X1 U14747 ( .C1(n12978), .C2(n12977), .A(n12983), .B(n12976), .ZN(
        n12982) );
  OAI211_X1 U14748 ( .C1(n12980), .C2(n13790), .A(n12984), .B(n12979), .ZN(
        n12981) );
  MUX2_X1 U14749 ( .A(n12982), .B(n12981), .S(n13012), .Z(n12986) );
  MUX2_X1 U14750 ( .A(n12984), .B(n12983), .S(n13012), .Z(n12985) );
  OAI211_X1 U14751 ( .C1(n12987), .C2(n12986), .A(n13765), .B(n12985), .ZN(
        n12991) );
  MUX2_X1 U14752 ( .A(n12989), .B(n12988), .S(n13012), .Z(n12990) );
  AND3_X1 U14753 ( .A1(n12991), .A2(n13073), .A3(n12990), .ZN(n12996) );
  INV_X1 U14754 ( .A(n13717), .ZN(n12994) );
  INV_X1 U14755 ( .A(n12992), .ZN(n12993) );
  MUX2_X1 U14756 ( .A(n12994), .B(n12993), .S(n13012), .Z(n12995) );
  AND2_X1 U14757 ( .A1(n13870), .A2(n13710), .ZN(n12998) );
  MUX2_X1 U14758 ( .A(n12998), .B(n12997), .S(n13002), .Z(n13000) );
  OAI33_X1 U14759 ( .A1(n13933), .A2(n13727), .A3(n13002), .B1(n13001), .B2(
        n13000), .B3(n12999), .ZN(n13003) );
  OAI211_X1 U14760 ( .C1(n13009), .C2(n13012), .A(n13008), .B(n13051), .ZN(
        n13015) );
  INV_X1 U14761 ( .A(n13015), .ZN(n13011) );
  INV_X1 U14762 ( .A(n13043), .ZN(n13013) );
  NAND2_X1 U14763 ( .A1(n13015), .A2(n13040), .ZN(n13016) );
  OAI22_X1 U14764 ( .A1(n7868), .A2(n13151), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13024) );
  INV_X1 U14765 ( .A(n13156), .ZN(n13022) );
  INV_X1 U14766 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15477) );
  AOI22_X1 U14767 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n9630), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n15477), .ZN(n13025) );
  INV_X1 U14768 ( .A(SI_31_), .ZN(n13970) );
  NOR2_X1 U14769 ( .A1(n13026), .A2(n13970), .ZN(n13027) );
  INV_X1 U14770 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13034) );
  NAND2_X1 U14771 ( .A1(n13029), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13032) );
  NAND2_X1 U14772 ( .A1(n13030), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13031) );
  OAI211_X1 U14773 ( .C1(n13034), .C2(n13033), .A(n13032), .B(n13031), .ZN(
        n13035) );
  INV_X1 U14774 ( .A(n13035), .ZN(n13036) );
  NAND2_X1 U14775 ( .A1(n13037), .A2(n13036), .ZN(n13618) );
  NAND2_X1 U14776 ( .A1(n15995), .A2(n13256), .ZN(n13045) );
  OAI21_X1 U14777 ( .B1(n16003), .B2(n13618), .A(n13045), .ZN(n13050) );
  NAND2_X1 U14778 ( .A1(n16003), .A2(n13618), .ZN(n13041) );
  OAI21_X1 U14779 ( .B1(n13038), .B2(n13050), .A(n13041), .ZN(n13085) );
  OAI21_X1 U14780 ( .B1(n15995), .B2(n13618), .A(n13040), .ZN(n13042) );
  NAND2_X1 U14781 ( .A1(n13041), .A2(n7242), .ZN(n13049) );
  AOI21_X1 U14782 ( .B1(n13045), .B2(n13618), .A(n16003), .ZN(n13046) );
  INV_X1 U14783 ( .A(n13049), .ZN(n13080) );
  INV_X1 U14784 ( .A(n13050), .ZN(n13079) );
  INV_X1 U14785 ( .A(n13051), .ZN(n13077) );
  INV_X1 U14786 ( .A(n13765), .ZN(n13757) );
  NOR3_X1 U14787 ( .A1(n13053), .A2(n8680), .A3(n8678), .ZN(n13056) );
  NAND4_X1 U14788 ( .A1(n13057), .A2(n13056), .A3(n13055), .A4(n13054), .ZN(
        n13060) );
  NOR4_X1 U14789 ( .A1(n13060), .A2(n13059), .A3(n13058), .A4(n7766), .ZN(
        n13064) );
  NAND4_X1 U14790 ( .A1(n13064), .A2(n13063), .A3(n13062), .A4(n13061), .ZN(
        n13068) );
  NOR4_X1 U14791 ( .A1(n13068), .A2(n13067), .A3(n7665), .A4(n13066), .ZN(
        n13069) );
  NAND4_X1 U14792 ( .A1(n13818), .A2(n13070), .A3(n13069), .A4(n13829), .ZN(
        n13071) );
  NOR4_X1 U14793 ( .A1(n13757), .A2(n13795), .A3(n13781), .A4(n13071), .ZN(
        n13072) );
  INV_X1 U14794 ( .A(n13728), .ZN(n13724) );
  NAND4_X1 U14795 ( .A1(n13719), .A2(n13073), .A3(n13072), .A4(n13724), .ZN(
        n13074) );
  NOR4_X1 U14796 ( .A1(n13077), .A2(n13076), .A3(n13075), .A4(n13074), .ZN(
        n13078) );
  NAND3_X1 U14797 ( .A1(n13080), .A2(n13079), .A3(n13078), .ZN(n13081) );
  XOR2_X1 U14798 ( .A(n13610), .B(n13081), .Z(n13082) );
  INV_X1 U14799 ( .A(n7186), .ZN(n13088) );
  NAND3_X1 U14800 ( .A1(n13089), .A2(n13088), .A3(n13087), .ZN(n13090) );
  OAI211_X1 U14801 ( .C1(n13092), .C2(n13091), .A(n13090), .B(P3_B_REG_SCAN_IN), .ZN(n13093) );
  NAND2_X1 U14802 ( .A1(n13094), .A2(n13093), .ZN(P3_U3296) );
  INV_X1 U14803 ( .A(n13095), .ZN(n13096) );
  AOI22_X1 U14804 ( .A1(n13096), .A2(n14054), .B1(n13994), .B2(n14065), .ZN(
        n13102) );
  NAND2_X1 U14805 ( .A1(n14047), .A2(n14251), .ZN(n13099) );
  INV_X1 U14806 ( .A(n13097), .ZN(n14255) );
  AOI22_X1 U14807 ( .A1(n14046), .A2(n14255), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13098) );
  OAI211_X1 U14808 ( .C1(n14032), .C2(n14050), .A(n13099), .B(n13098), .ZN(
        n13100) );
  AOI21_X1 U14809 ( .B1(n14407), .B2(n14035), .A(n13100), .ZN(n13101) );
  OAI21_X1 U14810 ( .B1(n13103), .B2(n13102), .A(n13101), .ZN(P2_U3207) );
  AOI22_X1 U14811 ( .A1(n14047), .A2(n14354), .B1(n13142), .B2(n14356), .ZN(
        n13104) );
  NAND2_X1 U14812 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n15561)
         );
  OAI211_X1 U14813 ( .C1(n14344), .C2(n14030), .A(n13104), .B(n15561), .ZN(
        n13111) );
  INV_X1 U14814 ( .A(n13105), .ZN(n13109) );
  AOI22_X1 U14815 ( .A1(n13106), .A2(n14054), .B1(n13994), .B2(n14354), .ZN(
        n13108) );
  NOR3_X1 U14816 ( .A1(n13109), .A2(n13108), .A3(n13107), .ZN(n13110) );
  AOI211_X1 U14817 ( .C1(n14433), .C2(n14035), .A(n13111), .B(n13110), .ZN(
        n13112) );
  OAI21_X1 U14818 ( .B1(n13113), .B2(n10844), .A(n13112), .ZN(P2_U3200) );
  AOI22_X1 U14819 ( .A1(n14047), .A2(n14069), .B1(n13142), .B2(n14068), .ZN(
        n13114) );
  NAND2_X1 U14820 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14110)
         );
  OAI211_X1 U14821 ( .C1(n13115), .C2(n14030), .A(n13114), .B(n14110), .ZN(
        n13121) );
  INV_X1 U14822 ( .A(n12441), .ZN(n13119) );
  AOI22_X1 U14823 ( .A1(n13116), .A2(n14054), .B1(n13994), .B2(n14069), .ZN(
        n13118) );
  NOR3_X1 U14824 ( .A1(n13119), .A2(n13118), .A3(n13117), .ZN(n13120) );
  AOI211_X1 U14825 ( .C1(n14438), .C2(n14035), .A(n13121), .B(n13120), .ZN(
        n13122) );
  OAI21_X1 U14826 ( .B1(n13105), .B2(n10844), .A(n13122), .ZN(P2_U3198) );
  INV_X1 U14827 ( .A(n13123), .ZN(n13133) );
  OAI22_X1 U14828 ( .A1(n14038), .A2(n13125), .B1(n13124), .B2(n10844), .ZN(
        n13132) );
  OAI22_X1 U14829 ( .A1(n14044), .A2(n13127), .B1(n13126), .B2(n11210), .ZN(
        n13131) );
  OAI22_X1 U14830 ( .A1(n13129), .A2(n14031), .B1(n14050), .B2(n13128), .ZN(
        n13130) );
  AOI211_X1 U14831 ( .C1(n13133), .C2(n13132), .A(n13131), .B(n13130), .ZN(
        n13134) );
  OAI21_X1 U14832 ( .B1(n13135), .B2(n10844), .A(n13134), .ZN(P2_U3194) );
  NAND3_X1 U14833 ( .A1(n13136), .A2(n13994), .A3(n14072), .ZN(n13137) );
  OAI21_X1 U14834 ( .B1(n13138), .B2(n10844), .A(n13137), .ZN(n13148) );
  INV_X1 U14835 ( .A(n13139), .ZN(n13147) );
  AOI22_X1 U14836 ( .A1(n14046), .A2(n13140), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13144) );
  AOI22_X1 U14837 ( .A1(n13142), .A2(n13141), .B1(n14047), .B2(n14072), .ZN(
        n13143) );
  OAI211_X1 U14838 ( .C1(n13145), .C2(n14044), .A(n13144), .B(n13143), .ZN(
        n13146) );
  AOI21_X1 U14839 ( .B1(n13148), .B2(n13147), .A(n13146), .ZN(n13149) );
  OAI21_X1 U14840 ( .B1(n11801), .B2(n10844), .A(n13149), .ZN(P2_U3196) );
  OAI222_X1 U14841 ( .A1(n15476), .A2(n14946), .B1(n13160), .B2(n13154), .C1(
        n13153), .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U14842 ( .A(SI_30_), .ZN(n13155) );
  OAI222_X1 U14843 ( .A1(n13158), .A2(P3_U3151), .B1(n13157), .B2(n13156), 
        .C1(n13155), .C2(n13983), .ZN(P3_U3265) );
  OAI222_X1 U14844 ( .A1(n15476), .A2(n7868), .B1(n13160), .B2(n14930), .C1(
        n13159), .C2(P1_U3086), .ZN(P1_U3325) );
  INV_X1 U14845 ( .A(n13206), .ZN(n13161) );
  AOI21_X1 U14846 ( .B1(n13690), .B2(n13162), .A(n13161), .ZN(n13167) );
  OAI22_X1 U14847 ( .A1(n13710), .A2(n13247), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13378), .ZN(n13164) );
  NOR2_X1 U14848 ( .A1(n13674), .A2(n13236), .ZN(n13163) );
  AOI211_X1 U14849 ( .C1(n13713), .C2(n13250), .A(n13164), .B(n13163), .ZN(
        n13166) );
  NAND2_X1 U14850 ( .A1(n13933), .A2(n13218), .ZN(n13165) );
  OAI211_X1 U14851 ( .C1(n13167), .C2(n13222), .A(n13166), .B(n13165), .ZN(
        P3_U3156) );
  XNOR2_X1 U14852 ( .A(n13169), .B(n13168), .ZN(n13174) );
  NAND2_X1 U14853 ( .A1(n13250), .A2(n13785), .ZN(n13171) );
  NOR2_X1 U14854 ( .A1(n13446), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13608) );
  AOI21_X1 U14855 ( .B1(n13245), .B2(n13741), .A(n13608), .ZN(n13170) );
  OAI211_X1 U14856 ( .C1(n13808), .C2(n13247), .A(n13171), .B(n13170), .ZN(
        n13172) );
  AOI21_X1 U14857 ( .B1(n13784), .B2(n13218), .A(n13172), .ZN(n13173) );
  OAI21_X1 U14858 ( .B1(n13174), .B2(n13222), .A(n13173), .ZN(P3_U3159) );
  XOR2_X1 U14859 ( .A(n13175), .B(n13176), .Z(n13181) );
  NAND2_X1 U14860 ( .A1(n13250), .A2(n13749), .ZN(n13178) );
  AOI22_X1 U14861 ( .A1(n13198), .A2(n13741), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13177) );
  OAI211_X1 U14862 ( .C1(n13710), .C2(n13236), .A(n13178), .B(n13177), .ZN(
        n13179) );
  AOI21_X1 U14863 ( .B1(n13873), .B2(n13218), .A(n13179), .ZN(n13180) );
  OAI21_X1 U14864 ( .B1(n13181), .B2(n13222), .A(n13180), .ZN(P3_U3163) );
  INV_X1 U14865 ( .A(n13182), .ZN(n13208) );
  INV_X1 U14866 ( .A(n13183), .ZN(n13185) );
  NOR3_X1 U14867 ( .A1(n13208), .A2(n13185), .A3(n13184), .ZN(n13188) );
  INV_X1 U14868 ( .A(n13186), .ZN(n13187) );
  OAI21_X1 U14869 ( .B1(n13188), .B2(n13187), .A(n13241), .ZN(n13192) );
  INV_X1 U14870 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n13369) );
  OAI22_X1 U14871 ( .A1(n13674), .A2(n13247), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13369), .ZN(n13190) );
  NOR2_X1 U14872 ( .A1(n13675), .A2(n13236), .ZN(n13189) );
  AOI211_X1 U14873 ( .C1(n13679), .C2(n13250), .A(n13190), .B(n13189), .ZN(
        n13191) );
  OAI211_X1 U14874 ( .C1(n13925), .C2(n13255), .A(n13192), .B(n13191), .ZN(
        P3_U3165) );
  XNOR2_X1 U14875 ( .A(n13193), .B(n13262), .ZN(n13244) );
  NAND2_X1 U14876 ( .A1(n13244), .A2(n13243), .ZN(n13242) );
  OAI21_X1 U14877 ( .B1(n13832), .B2(n13193), .A(n13242), .ZN(n13196) );
  XNOR2_X1 U14878 ( .A(n13194), .B(n13809), .ZN(n13195) );
  XNOR2_X1 U14879 ( .A(n13196), .B(n13195), .ZN(n13203) );
  NAND2_X1 U14880 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13546)
         );
  OAI21_X1 U14881 ( .B1(n13236), .B2(n13834), .A(n13546), .ZN(n13197) );
  AOI21_X1 U14882 ( .B1(n13198), .B2(n13262), .A(n13197), .ZN(n13199) );
  OAI21_X1 U14883 ( .B1(n13200), .B2(n13837), .A(n13199), .ZN(n13201) );
  AOI21_X1 U14884 ( .B1(n13836), .B2(n13218), .A(n13201), .ZN(n13202) );
  OAI21_X1 U14885 ( .B1(n13203), .B2(n13222), .A(n13202), .ZN(P3_U3166) );
  AND3_X1 U14886 ( .A1(n13206), .A2(n13205), .A3(n13204), .ZN(n13207) );
  OAI21_X1 U14887 ( .B1(n13208), .B2(n13207), .A(n13241), .ZN(n13212) );
  AOI22_X1 U14888 ( .A1(n13691), .A2(n13245), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13209) );
  OAI21_X1 U14889 ( .B1(n13727), .B2(n13247), .A(n13209), .ZN(n13210) );
  AOI21_X1 U14890 ( .B1(n13698), .B2(n13250), .A(n13210), .ZN(n13211) );
  OAI211_X1 U14891 ( .C1(n13255), .C2(n13927), .A(n13212), .B(n13211), .ZN(
        P3_U3169) );
  XNOR2_X1 U14892 ( .A(n13213), .B(n13214), .ZN(n13223) );
  NOR2_X1 U14893 ( .A1(n13247), .A2(n13800), .ZN(n13217) );
  INV_X1 U14894 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n13215) );
  OAI22_X1 U14895 ( .A1(n13236), .A2(n13763), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13215), .ZN(n13216) );
  AOI211_X1 U14896 ( .C1(n13768), .C2(n13250), .A(n13217), .B(n13216), .ZN(
        n13221) );
  NAND2_X1 U14897 ( .A1(n13219), .A2(n13218), .ZN(n13220) );
  OAI211_X1 U14898 ( .C1(n13223), .C2(n13222), .A(n13221), .B(n13220), .ZN(
        P3_U3173) );
  INV_X1 U14899 ( .A(n13870), .ZN(n13734) );
  OAI21_X1 U14900 ( .B1(n9798), .B2(n13710), .A(n13225), .ZN(n13226) );
  NAND2_X1 U14901 ( .A1(n13226), .A2(n13241), .ZN(n13231) );
  OAI22_X1 U14902 ( .A1(n13247), .A2(n13763), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13227), .ZN(n13229) );
  NOR2_X1 U14903 ( .A1(n13727), .A2(n13236), .ZN(n13228) );
  AOI211_X1 U14904 ( .C1(n13732), .C2(n13250), .A(n13229), .B(n13228), .ZN(
        n13230) );
  OAI211_X1 U14905 ( .C1(n13734), .C2(n13255), .A(n13231), .B(n13230), .ZN(
        P3_U3175) );
  OAI21_X1 U14906 ( .B1(n13234), .B2(n13233), .A(n13232), .ZN(n13235) );
  NAND2_X1 U14907 ( .A1(n13235), .A2(n13241), .ZN(n13240) );
  INV_X1 U14908 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n13269) );
  OAI22_X1 U14909 ( .A1(n13662), .A2(n13247), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13269), .ZN(n13238) );
  NOR2_X1 U14910 ( .A1(n13663), .A2(n13236), .ZN(n13237) );
  AOI211_X1 U14911 ( .C1(n13666), .C2(n13250), .A(n13238), .B(n13237), .ZN(
        n13239) );
  OAI211_X1 U14912 ( .C1(n13921), .C2(n13255), .A(n13240), .B(n13239), .ZN(
        P3_U3180) );
  OAI211_X1 U14913 ( .C1(n13244), .C2(n13243), .A(n13242), .B(n13241), .ZN(
        n13253) );
  INV_X1 U14914 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13268) );
  NOR2_X1 U14915 ( .A1(n13268), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13513) );
  AOI21_X1 U14916 ( .B1(n13245), .B2(n13261), .A(n13513), .ZN(n13246) );
  OAI21_X1 U14917 ( .B1(n13248), .B2(n13247), .A(n13246), .ZN(n13249) );
  AOI21_X1 U14918 ( .B1(n13251), .B2(n13250), .A(n13249), .ZN(n13252) );
  OAI211_X1 U14919 ( .C1(n13255), .C2(n13254), .A(n13253), .B(n13252), .ZN(
        P3_U3181) );
  MUX2_X1 U14920 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13618), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14921 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n13256), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14922 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13652), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14923 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13257), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14924 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13651), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14925 ( .A(n13691), .B(P3_DATAO_REG_25__SCAN_IN), .S(n13265), .Z(
        P3_U3516) );
  MUX2_X1 U14926 ( .A(n13708), .B(P3_DATAO_REG_24__SCAN_IN), .S(n13265), .Z(
        P3_U3515) );
  MUX2_X1 U14927 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13690), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14928 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13743), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14929 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13258), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14930 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13741), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14931 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13760), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14932 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13259), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14933 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13260), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14934 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13261), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14935 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13262), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14936 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13263), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14937 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n9776), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14938 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13264), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14939 ( .A(n13266), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13265), .Z(
        n13478) );
  OAI22_X1 U14940 ( .A1(n13269), .A2(keyinput_62), .B1(n13268), .B2(
        keyinput_63), .ZN(n13267) );
  AOI221_X1 U14941 ( .B1(n13269), .B2(keyinput_62), .C1(keyinput_63), .C2(
        n13268), .A(n13267), .ZN(n13476) );
  OAI22_X1 U14942 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_57), .B1(
        P3_REG3_REG_13__SCAN_IN), .B2(keyinput_56), .ZN(n13270) );
  AOI221_X1 U14943 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .C1(
        keyinput_56), .C2(P3_REG3_REG_13__SCAN_IN), .A(n13270), .ZN(n13357) );
  INV_X1 U14944 ( .A(keyinput_44), .ZN(n13340) );
  INV_X1 U14945 ( .A(keyinput_43), .ZN(n13338) );
  AOI22_X1 U14946 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_39), .B1(
        P3_REG3_REG_19__SCAN_IN), .B2(keyinput_41), .ZN(n13271) );
  OAI221_X1 U14947 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_41), .A(n13271), .ZN(n13335) );
  XOR2_X1 U14948 ( .A(n13272), .B(keyinput_18), .Z(n13302) );
  INV_X1 U14949 ( .A(keyinput_17), .ZN(n13297) );
  INV_X1 U14950 ( .A(keyinput_16), .ZN(n13295) );
  INV_X1 U14951 ( .A(keyinput_15), .ZN(n13293) );
  OAI22_X1 U14952 ( .A1(n13403), .A2(keyinput_13), .B1(SI_20_), .B2(
        keyinput_12), .ZN(n13273) );
  AOI221_X1 U14953 ( .B1(n13403), .B2(keyinput_13), .C1(keyinput_12), .C2(
        SI_20_), .A(n13273), .ZN(n13289) );
  INV_X1 U14954 ( .A(keyinput_11), .ZN(n13287) );
  OAI22_X1 U14955 ( .A1(SI_29_), .A2(keyinput_3), .B1(SI_30_), .B2(keyinput_2), 
        .ZN(n13274) );
  AOI221_X1 U14956 ( .B1(SI_29_), .B2(keyinput_3), .C1(keyinput_2), .C2(SI_30_), .A(n13274), .ZN(n13279) );
  AOI22_X1 U14957 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n13275) );
  OAI221_X1 U14958 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n13275), .ZN(n13278) );
  AOI22_X1 U14959 ( .A1(SI_27_), .A2(keyinput_5), .B1(SI_28_), .B2(keyinput_4), 
        .ZN(n13276) );
  OAI221_X1 U14960 ( .B1(SI_27_), .B2(keyinput_5), .C1(SI_28_), .C2(keyinput_4), .A(n13276), .ZN(n13277) );
  AOI21_X1 U14961 ( .B1(n13279), .B2(n13278), .A(n13277), .ZN(n13285) );
  XNOR2_X1 U14962 ( .A(SI_26_), .B(keyinput_6), .ZN(n13284) );
  OAI22_X1 U14963 ( .A1(SI_25_), .A2(keyinput_7), .B1(SI_22_), .B2(keyinput_10), .ZN(n13280) );
  AOI221_X1 U14964 ( .B1(SI_25_), .B2(keyinput_7), .C1(keyinput_10), .C2(
        SI_22_), .A(n13280), .ZN(n13283) );
  OAI22_X1 U14965 ( .A1(SI_24_), .A2(keyinput_8), .B1(SI_23_), .B2(keyinput_9), 
        .ZN(n13281) );
  AOI221_X1 U14966 ( .B1(SI_24_), .B2(keyinput_8), .C1(keyinput_9), .C2(SI_23_), .A(n13281), .ZN(n13282) );
  OAI211_X1 U14967 ( .C1(n13285), .C2(n13284), .A(n13283), .B(n13282), .ZN(
        n13286) );
  OAI221_X1 U14968 ( .B1(SI_21_), .B2(keyinput_11), .C1(n13398), .C2(n13287), 
        .A(n13286), .ZN(n13288) );
  OAI211_X1 U14969 ( .C1(n13291), .C2(keyinput_14), .A(n13289), .B(n13288), 
        .ZN(n13290) );
  AOI21_X1 U14970 ( .B1(n13291), .B2(keyinput_14), .A(n13290), .ZN(n13292) );
  AOI221_X1 U14971 ( .B1(SI_17_), .B2(keyinput_15), .C1(n13405), .C2(n13293), 
        .A(n13292), .ZN(n13294) );
  AOI221_X1 U14972 ( .B1(SI_16_), .B2(n13295), .C1(n13409), .C2(keyinput_16), 
        .A(n13294), .ZN(n13296) );
  AOI221_X1 U14973 ( .B1(SI_15_), .B2(keyinput_17), .C1(n13412), .C2(n13297), 
        .A(n13296), .ZN(n13301) );
  OAI22_X1 U14974 ( .A1(n13299), .A2(keyinput_19), .B1(keyinput_20), .B2(
        SI_12_), .ZN(n13298) );
  AOI221_X1 U14975 ( .B1(n13299), .B2(keyinput_19), .C1(SI_12_), .C2(
        keyinput_20), .A(n13298), .ZN(n13300) );
  OAI21_X1 U14976 ( .B1(n13302), .B2(n13301), .A(n13300), .ZN(n13311) );
  OAI22_X1 U14977 ( .A1(n13304), .A2(keyinput_22), .B1(keyinput_21), .B2(
        SI_11_), .ZN(n13303) );
  AOI221_X1 U14978 ( .B1(n13304), .B2(keyinput_22), .C1(SI_11_), .C2(
        keyinput_21), .A(n13303), .ZN(n13310) );
  AOI22_X1 U14979 ( .A1(SI_6_), .A2(keyinput_26), .B1(SI_7_), .B2(keyinput_25), 
        .ZN(n13305) );
  OAI221_X1 U14980 ( .B1(SI_6_), .B2(keyinput_26), .C1(SI_7_), .C2(keyinput_25), .A(n13305), .ZN(n13309) );
  XNOR2_X1 U14981 ( .A(SI_9_), .B(keyinput_23), .ZN(n13307) );
  XNOR2_X1 U14982 ( .A(SI_8_), .B(keyinput_24), .ZN(n13306) );
  NAND2_X1 U14983 ( .A1(n13307), .A2(n13306), .ZN(n13308) );
  AOI211_X1 U14984 ( .C1(n13311), .C2(n13310), .A(n13309), .B(n13308), .ZN(
        n13316) );
  INV_X1 U14985 ( .A(keyinput_27), .ZN(n13312) );
  MUX2_X1 U14986 ( .A(keyinput_27), .B(n13312), .S(SI_5_), .Z(n13315) );
  XOR2_X1 U14987 ( .A(SI_4_), .B(keyinput_28), .Z(n13314) );
  XNOR2_X1 U14988 ( .A(SI_3_), .B(keyinput_29), .ZN(n13313) );
  OAI211_X1 U14989 ( .C1(n13316), .C2(n13315), .A(n13314), .B(n13313), .ZN(
        n13318) );
  NAND2_X1 U14990 ( .A1(SI_2_), .A2(keyinput_30), .ZN(n13317) );
  OAI211_X1 U14991 ( .C1(SI_2_), .C2(keyinput_30), .A(n13318), .B(n13317), 
        .ZN(n13321) );
  INV_X1 U14992 ( .A(keyinput_31), .ZN(n13319) );
  MUX2_X1 U14993 ( .A(keyinput_31), .B(n13319), .S(SI_1_), .Z(n13320) );
  NAND2_X1 U14994 ( .A1(n13321), .A2(n13320), .ZN(n13324) );
  INV_X1 U14995 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15723) );
  OAI22_X1 U14996 ( .A1(n15723), .A2(keyinput_33), .B1(SI_0_), .B2(keyinput_32), .ZN(n13322) );
  AOI221_X1 U14997 ( .B1(n15723), .B2(keyinput_33), .C1(keyinput_32), .C2(
        SI_0_), .A(n13322), .ZN(n13323) );
  AOI22_X1 U14998 ( .A1(n13324), .A2(n13323), .B1(P3_STATE_REG_SCAN_IN), .B2(
        keyinput_34), .ZN(n13327) );
  AOI22_X1 U14999 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_36), .B1(n13378), .B2(keyinput_38), .ZN(n13325) );
  OAI221_X1 U15000 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_36), .C1(
        n13378), .C2(keyinput_38), .A(n13325), .ZN(n13326) );
  AOI221_X1 U15001 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n13327), .C1(keyinput_34), 
        .C2(n13327), .A(n13326), .ZN(n13331) );
  OAI22_X1 U15002 ( .A1(n13379), .A2(keyinput_37), .B1(n13329), .B2(
        keyinput_35), .ZN(n13328) );
  AOI221_X1 U15003 ( .B1(n13379), .B2(keyinput_37), .C1(keyinput_35), .C2(
        n13329), .A(n13328), .ZN(n13330) );
  AOI22_X1 U15004 ( .A1(n13331), .A2(n13330), .B1(keyinput_40), .B2(n13333), 
        .ZN(n13332) );
  OAI21_X1 U15005 ( .B1(keyinput_40), .B2(n13333), .A(n13332), .ZN(n13334) );
  OAI22_X1 U15006 ( .A1(n13335), .A2(n13334), .B1(keyinput_42), .B2(
        P3_REG3_REG_28__SCAN_IN), .ZN(n13336) );
  AOI21_X1 U15007 ( .B1(keyinput_42), .B2(P3_REG3_REG_28__SCAN_IN), .A(n13336), 
        .ZN(n13337) );
  AOI221_X1 U15008 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .C1(n13454), .C2(n13338), .A(n13337), .ZN(n13339) );
  AOI221_X1 U15009 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .C1(n10513), .C2(n13340), .A(n13339), .ZN(n13355) );
  OAI22_X1 U15010 ( .A1(n13369), .A2(keyinput_47), .B1(keyinput_49), .B2(
        P3_REG3_REG_5__SCAN_IN), .ZN(n13341) );
  AOI221_X1 U15011 ( .B1(n13369), .B2(keyinput_47), .C1(P3_REG3_REG_5__SCAN_IN), .C2(keyinput_49), .A(n13341), .ZN(n13350) );
  INV_X1 U15012 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13343) );
  OAI22_X1 U15013 ( .A1(n13344), .A2(keyinput_50), .B1(n13343), .B2(
        keyinput_46), .ZN(n13342) );
  AOI221_X1 U15014 ( .B1(n13344), .B2(keyinput_50), .C1(keyinput_46), .C2(
        n13343), .A(n13342), .ZN(n13349) );
  OAI22_X1 U15015 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_51), .B1(
        keyinput_48), .B2(P3_REG3_REG_16__SCAN_IN), .ZN(n13345) );
  AOI221_X1 U15016 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput_48), .A(n13345), .ZN(n13348) );
  OAI22_X1 U15017 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_45), .B1(
        P3_REG3_REG_4__SCAN_IN), .B2(keyinput_52), .ZN(n13346) );
  AOI221_X1 U15018 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(
        keyinput_52), .C2(P3_REG3_REG_4__SCAN_IN), .A(n13346), .ZN(n13347) );
  NAND4_X1 U15019 ( .A1(n13350), .A2(n13349), .A3(n13348), .A4(n13347), .ZN(
        n13354) );
  OAI22_X1 U15020 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_53), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .ZN(n13351) );
  AOI221_X1 U15021 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_53), .C1(
        keyinput_54), .C2(P3_REG3_REG_0__SCAN_IN), .A(n13351), .ZN(n13353) );
  XNOR2_X1 U15022 ( .A(P3_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n13352)
         );
  OAI211_X1 U15023 ( .C1(n13355), .C2(n13354), .A(n13353), .B(n13352), .ZN(
        n13356) );
  OAI211_X1 U15024 ( .C1(P3_REG3_REG_11__SCAN_IN), .C2(keyinput_58), .A(n13357), .B(n13356), .ZN(n13358) );
  AOI21_X1 U15025 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .A(n13358), 
        .ZN(n13362) );
  AOI22_X1 U15026 ( .A1(n10660), .A2(keyinput_59), .B1(n13360), .B2(
        keyinput_60), .ZN(n13359) );
  OAI221_X1 U15027 ( .B1(n10660), .B2(keyinput_59), .C1(n13360), .C2(
        keyinput_60), .A(n13359), .ZN(n13361) );
  AOI211_X1 U15028 ( .C1(n13364), .C2(keyinput_61), .A(n13362), .B(n13361), 
        .ZN(n13363) );
  OAI21_X1 U15029 ( .B1(n13364), .B2(keyinput_61), .A(n13363), .ZN(n13475) );
  OAI22_X1 U15030 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_124), .B1(
        keyinput_123), .B2(P3_REG3_REG_2__SCAN_IN), .ZN(n13365) );
  AOI221_X1 U15031 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_124), .C1(
        P3_REG3_REG_2__SCAN_IN), .C2(keyinput_123), .A(n13365), .ZN(n13470) );
  AOI22_X1 U15032 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_110), .B1(
        n13367), .B2(keyinput_116), .ZN(n13366) );
  OAI221_X1 U15033 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .C1(
        n13367), .C2(keyinput_116), .A(n13366), .ZN(n13376) );
  AOI22_X1 U15034 ( .A1(n13370), .A2(keyinput_112), .B1(n13369), .B2(
        keyinput_111), .ZN(n13368) );
  OAI221_X1 U15035 ( .B1(n13370), .B2(keyinput_112), .C1(n13369), .C2(
        keyinput_111), .A(n13368), .ZN(n13375) );
  AOI22_X1 U15036 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput_113), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_114), .ZN(n13371) );
  OAI221_X1 U15037 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_114), .A(n13371), .ZN(n13374)
         );
  AOI22_X1 U15038 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(keyinput_109), .B1(
        P3_REG3_REG_24__SCAN_IN), .B2(keyinput_115), .ZN(n13372) );
  OAI221_X1 U15039 ( .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_109), .C1(
        P3_REG3_REG_24__SCAN_IN), .C2(keyinput_115), .A(n13372), .ZN(n13373)
         );
  NOR4_X1 U15040 ( .A1(n13376), .A2(n13375), .A3(n13374), .A4(n13373), .ZN(
        n13462) );
  INV_X1 U15041 ( .A(keyinput_108), .ZN(n13456) );
  INV_X1 U15042 ( .A(keyinput_107), .ZN(n13453) );
  AOI22_X1 U15043 ( .A1(n13379), .A2(keyinput_101), .B1(n13378), .B2(
        keyinput_102), .ZN(n13377) );
  OAI221_X1 U15044 ( .B1(n13379), .B2(keyinput_101), .C1(n13378), .C2(
        keyinput_102), .A(n13377), .ZN(n13444) );
  XOR2_X1 U15045 ( .A(SI_14_), .B(keyinput_82), .Z(n13417) );
  INV_X1 U15046 ( .A(keyinput_81), .ZN(n13411) );
  INV_X1 U15047 ( .A(keyinput_80), .ZN(n13408) );
  INV_X1 U15048 ( .A(keyinput_79), .ZN(n13406) );
  OAI22_X1 U15049 ( .A1(n13381), .A2(keyinput_76), .B1(SI_18_), .B2(
        keyinput_78), .ZN(n13380) );
  AOI221_X1 U15050 ( .B1(n13381), .B2(keyinput_76), .C1(keyinput_78), .C2(
        SI_18_), .A(n13380), .ZN(n13401) );
  INV_X1 U15051 ( .A(keyinput_75), .ZN(n13399) );
  OAI22_X1 U15052 ( .A1(SI_29_), .A2(keyinput_67), .B1(keyinput_66), .B2(
        SI_30_), .ZN(n13382) );
  AOI221_X1 U15053 ( .B1(SI_29_), .B2(keyinput_67), .C1(SI_30_), .C2(
        keyinput_66), .A(n13382), .ZN(n13388) );
  AOI22_X1 U15054 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_64), .B1(SI_31_), 
        .B2(keyinput_65), .ZN(n13383) );
  OAI221_X1 U15055 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_64), .C1(SI_31_), 
        .C2(keyinput_65), .A(n13383), .ZN(n13387) );
  AOI22_X1 U15056 ( .A1(SI_28_), .A2(keyinput_68), .B1(n13385), .B2(
        keyinput_69), .ZN(n13384) );
  OAI221_X1 U15057 ( .B1(SI_28_), .B2(keyinput_68), .C1(n13385), .C2(
        keyinput_69), .A(n13384), .ZN(n13386) );
  AOI21_X1 U15058 ( .B1(n13388), .B2(n13387), .A(n13386), .ZN(n13396) );
  XNOR2_X1 U15059 ( .A(SI_26_), .B(keyinput_70), .ZN(n13395) );
  OAI22_X1 U15060 ( .A1(n13391), .A2(keyinput_72), .B1(n13390), .B2(
        keyinput_73), .ZN(n13389) );
  AOI221_X1 U15061 ( .B1(n13391), .B2(keyinput_72), .C1(keyinput_73), .C2(
        n13390), .A(n13389), .ZN(n13394) );
  OAI22_X1 U15062 ( .A1(SI_25_), .A2(keyinput_71), .B1(keyinput_74), .B2(
        SI_22_), .ZN(n13392) );
  AOI221_X1 U15063 ( .B1(SI_25_), .B2(keyinput_71), .C1(SI_22_), .C2(
        keyinput_74), .A(n13392), .ZN(n13393) );
  OAI211_X1 U15064 ( .C1(n13396), .C2(n13395), .A(n13394), .B(n13393), .ZN(
        n13397) );
  OAI221_X1 U15065 ( .B1(SI_21_), .B2(n13399), .C1(n13398), .C2(keyinput_75), 
        .A(n13397), .ZN(n13400) );
  OAI211_X1 U15066 ( .C1(n13403), .C2(keyinput_77), .A(n13401), .B(n13400), 
        .ZN(n13402) );
  AOI21_X1 U15067 ( .B1(n13403), .B2(keyinput_77), .A(n13402), .ZN(n13404) );
  AOI221_X1 U15068 ( .B1(SI_17_), .B2(n13406), .C1(n13405), .C2(keyinput_79), 
        .A(n13404), .ZN(n13407) );
  AOI221_X1 U15069 ( .B1(SI_16_), .B2(keyinput_80), .C1(n13409), .C2(n13408), 
        .A(n13407), .ZN(n13410) );
  AOI221_X1 U15070 ( .B1(SI_15_), .B2(keyinput_81), .C1(n13412), .C2(n13411), 
        .A(n13410), .ZN(n13416) );
  OAI22_X1 U15071 ( .A1(n13414), .A2(keyinput_84), .B1(SI_13_), .B2(
        keyinput_83), .ZN(n13413) );
  AOI221_X1 U15072 ( .B1(n13414), .B2(keyinput_84), .C1(keyinput_83), .C2(
        SI_13_), .A(n13413), .ZN(n13415) );
  OAI21_X1 U15073 ( .B1(n13417), .B2(n13416), .A(n13415), .ZN(n13426) );
  OAI22_X1 U15074 ( .A1(n13419), .A2(keyinput_85), .B1(keyinput_86), .B2(
        SI_10_), .ZN(n13418) );
  AOI221_X1 U15075 ( .B1(n13419), .B2(keyinput_85), .C1(SI_10_), .C2(
        keyinput_86), .A(n13418), .ZN(n13425) );
  AOI22_X1 U15076 ( .A1(SI_8_), .A2(keyinput_88), .B1(SI_9_), .B2(keyinput_87), 
        .ZN(n13420) );
  OAI221_X1 U15077 ( .B1(SI_8_), .B2(keyinput_88), .C1(SI_9_), .C2(keyinput_87), .A(n13420), .ZN(n13424) );
  XNOR2_X1 U15078 ( .A(SI_7_), .B(keyinput_89), .ZN(n13422) );
  XNOR2_X1 U15079 ( .A(SI_6_), .B(keyinput_90), .ZN(n13421) );
  NAND2_X1 U15080 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  AOI211_X1 U15081 ( .C1(n13426), .C2(n13425), .A(n13424), .B(n13423), .ZN(
        n13431) );
  INV_X1 U15082 ( .A(keyinput_91), .ZN(n13427) );
  MUX2_X1 U15083 ( .A(keyinput_91), .B(n13427), .S(SI_5_), .Z(n13430) );
  XOR2_X1 U15084 ( .A(SI_4_), .B(keyinput_92), .Z(n13429) );
  XNOR2_X1 U15085 ( .A(SI_3_), .B(keyinput_93), .ZN(n13428) );
  OAI211_X1 U15086 ( .C1(n13431), .C2(n13430), .A(n13429), .B(n13428), .ZN(
        n13435) );
  XNOR2_X1 U15087 ( .A(SI_2_), .B(keyinput_94), .ZN(n13434) );
  INV_X1 U15088 ( .A(keyinput_95), .ZN(n13432) );
  MUX2_X1 U15089 ( .A(keyinput_95), .B(n13432), .S(SI_1_), .Z(n13433) );
  AOI21_X1 U15090 ( .B1(n13435), .B2(n13434), .A(n13433), .ZN(n13439) );
  XOR2_X1 U15091 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_97), .Z(n13437) );
  XNOR2_X1 U15092 ( .A(SI_0_), .B(keyinput_96), .ZN(n13436) );
  NAND2_X1 U15093 ( .A1(n13437), .A2(n13436), .ZN(n13438) );
  OAI22_X1 U15094 ( .A1(n13439), .A2(n13438), .B1(P3_STATE_REG_SCAN_IN), .B2(
        keyinput_98), .ZN(n13442) );
  OAI22_X1 U15095 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_100), .B1(
        keyinput_99), .B2(P3_REG3_REG_7__SCAN_IN), .ZN(n13440) );
  AOI221_X1 U15096 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_100), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput_99), .A(n13440), .ZN(n13441) );
  OAI221_X1 U15097 ( .B1(n13442), .B2(keyinput_98), .C1(n13442), .C2(
        P3_STATE_REG_SCAN_IN), .A(n13441), .ZN(n13443) );
  OAI22_X1 U15098 ( .A1(n13444), .A2(n13443), .B1(n13446), .B2(keyinput_105), 
        .ZN(n13445) );
  AOI21_X1 U15099 ( .B1(n13446), .B2(keyinput_105), .A(n13445), .ZN(n13450) );
  OAI22_X1 U15100 ( .A1(n13448), .A2(keyinput_103), .B1(keyinput_104), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n13447) );
  AOI221_X1 U15101 ( .B1(n13448), .B2(keyinput_103), .C1(
        P3_REG3_REG_3__SCAN_IN), .C2(keyinput_104), .A(n13447), .ZN(n13449) );
  AOI22_X1 U15102 ( .A1(n13450), .A2(n13449), .B1(keyinput_106), .B2(
        P3_REG3_REG_28__SCAN_IN), .ZN(n13451) );
  OAI21_X1 U15103 ( .B1(keyinput_106), .B2(P3_REG3_REG_28__SCAN_IN), .A(n13451), .ZN(n13452) );
  OAI221_X1 U15104 ( .B1(P3_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        n13454), .C2(n13453), .A(n13452), .ZN(n13455) );
  OAI221_X1 U15105 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n13456), .C1(n10513), 
        .C2(keyinput_108), .A(n13455), .ZN(n13461) );
  XNOR2_X1 U15106 ( .A(keyinput_118), .B(n13457), .ZN(n13460) );
  AOI22_X1 U15107 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(keyinput_119), .B1(n8154), .B2(keyinput_117), .ZN(n13458) );
  OAI221_X1 U15108 ( .B1(P3_REG3_REG_20__SCAN_IN), .B2(keyinput_119), .C1(
        n8154), .C2(keyinput_117), .A(n13458), .ZN(n13459) );
  AOI211_X1 U15109 ( .C1(n13462), .C2(n13461), .A(n13460), .B(n13459), .ZN(
        n13466) );
  AOI22_X1 U15110 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput_121), .B1(
        n13464), .B2(keyinput_122), .ZN(n13463) );
  OAI221_X1 U15111 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .C1(
        n13464), .C2(keyinput_122), .A(n13463), .ZN(n13465) );
  AOI211_X1 U15112 ( .C1(n13468), .C2(keyinput_120), .A(n13466), .B(n13465), 
        .ZN(n13467) );
  OAI21_X1 U15113 ( .B1(n13468), .B2(keyinput_120), .A(n13467), .ZN(n13469) );
  OAI211_X1 U15114 ( .C1(P3_REG3_REG_6__SCAN_IN), .C2(keyinput_125), .A(n13470), .B(n13469), .ZN(n13471) );
  AOI21_X1 U15115 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_125), .A(n13471), 
        .ZN(n13474) );
  AOI22_X1 U15116 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_127), .B1(
        P3_REG3_REG_26__SCAN_IN), .B2(keyinput_126), .ZN(n13472) );
  OAI221_X1 U15117 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_127), .C1(
        P3_REG3_REG_26__SCAN_IN), .C2(keyinput_126), .A(n13472), .ZN(n13473)
         );
  AOI211_X1 U15118 ( .C1(n13476), .C2(n13475), .A(n13474), .B(n13473), .ZN(
        n13477) );
  XOR2_X1 U15119 ( .A(n13478), .B(n13477), .Z(P3_U3502) );
  MUX2_X1 U15120 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13479), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15121 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n7681), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15122 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13480), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15123 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13481), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15124 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13482), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15125 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13483), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15126 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13484), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15127 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13485), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15128 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13486), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15129 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13487), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15130 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n13488), .S(P3_U3897), .Z(
        P3_U3491) );
  OAI21_X1 U15131 ( .B1(n13490), .B2(P3_REG2_REG_13__SCAN_IN), .A(n13489), 
        .ZN(n13491) );
  INV_X1 U15132 ( .A(n13491), .ZN(n13505) );
  OAI21_X1 U15133 ( .B1(n13494), .B2(n13493), .A(n13492), .ZN(n13503) );
  AOI21_X1 U15134 ( .B1(n13496), .B2(n12290), .A(n13495), .ZN(n13497) );
  NOR2_X1 U15135 ( .A1(n15718), .A2(n13497), .ZN(n13498) );
  AOI211_X1 U15136 ( .C1(n15702), .C2(P3_ADDR_REG_13__SCAN_IN), .A(n13499), 
        .B(n13498), .ZN(n13500) );
  OAI21_X1 U15137 ( .B1(n13501), .B2(n13611), .A(n13500), .ZN(n13502) );
  AOI21_X1 U15138 ( .B1(n13503), .B2(n15712), .A(n13502), .ZN(n13504) );
  OAI21_X1 U15139 ( .B1(n13505), .B2(n15677), .A(n13504), .ZN(P3_U3195) );
  AND2_X1 U15140 ( .A1(n13517), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13506) );
  OAI21_X1 U15141 ( .B1(n13508), .B2(n13536), .A(n13528), .ZN(n13509) );
  AOI21_X1 U15142 ( .B1(n13509), .B2(n13519), .A(n13529), .ZN(n13527) );
  INV_X1 U15143 ( .A(n13536), .ZN(n13525) );
  AOI22_X1 U15144 ( .A1(n13517), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n13511), 
        .B2(n13510), .ZN(n13512) );
  NOR2_X1 U15145 ( .A1(n13512), .A2(n13525), .ZN(n13540) );
  AOI21_X1 U15146 ( .B1(n7221), .B2(n13520), .A(n13539), .ZN(n13515) );
  AOI21_X1 U15147 ( .B1(n15702), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13513), 
        .ZN(n13514) );
  OAI21_X1 U15148 ( .B1(n13515), .B2(n15677), .A(n13514), .ZN(n13524) );
  MUX2_X1 U15149 ( .A(n13520), .B(n13519), .S(n13087), .Z(n13521) );
  NOR2_X1 U15150 ( .A1(n13522), .A2(n13521), .ZN(n13534) );
  AOI211_X1 U15151 ( .C1(n13522), .C2(n13521), .A(n15681), .B(n13534), .ZN(
        n13523) );
  AOI211_X1 U15152 ( .C1(n15704), .C2(n13525), .A(n13524), .B(n13523), .ZN(
        n13526) );
  OAI21_X1 U15153 ( .B1(n13527), .B2(n15718), .A(n13526), .ZN(P3_U3197) );
  INV_X1 U15154 ( .A(n13528), .ZN(n13530) );
  AOI22_X1 U15155 ( .A1(n13541), .A2(P3_REG1_REG_16__SCAN_IN), .B1(n13903), 
        .B2(n13564), .ZN(n13531) );
  AOI21_X1 U15156 ( .B1(n13532), .B2(n13531), .A(n13552), .ZN(n13551) );
  INV_X1 U15157 ( .A(n13533), .ZN(n13535) );
  MUX2_X1 U15158 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13087), .Z(n13558) );
  XNOR2_X1 U15159 ( .A(n13558), .B(n13541), .ZN(n13537) );
  NAND2_X1 U15160 ( .A1(n13538), .A2(n13537), .ZN(n13557) );
  OAI21_X1 U15161 ( .B1(n13538), .B2(n13537), .A(n13557), .ZN(n13549) );
  AOI22_X1 U15162 ( .A1(n13541), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n13838), 
        .B2(n13564), .ZN(n13542) );
  AOI21_X1 U15163 ( .B1(n13543), .B2(n13542), .A(n13563), .ZN(n13544) );
  NOR2_X1 U15164 ( .A1(n13544), .A2(n15677), .ZN(n13548) );
  NAND2_X1 U15165 ( .A1(n15702), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n13545) );
  OAI211_X1 U15166 ( .C1(n13611), .C2(n13564), .A(n13546), .B(n13545), .ZN(
        n13547) );
  AOI211_X1 U15167 ( .C1(n13549), .C2(n15712), .A(n13548), .B(n13547), .ZN(
        n13550) );
  OAI21_X1 U15168 ( .B1(n13551), .B2(n15718), .A(n13550), .ZN(P3_U3198) );
  NOR2_X1 U15169 ( .A1(n13554), .A2(n13553), .ZN(n13571) );
  AOI21_X1 U15170 ( .B1(n13554), .B2(n13553), .A(n13571), .ZN(n13569) );
  OAI21_X1 U15171 ( .B1(n13577), .B2(n13556), .A(n13555), .ZN(n13562) );
  MUX2_X1 U15172 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13087), .Z(n13580) );
  XNOR2_X1 U15173 ( .A(n13580), .B(n13579), .ZN(n13560) );
  OAI21_X1 U15174 ( .B1(n13558), .B2(n13564), .A(n13557), .ZN(n13559) );
  NOR2_X1 U15175 ( .A1(n13559), .A2(n13560), .ZN(n13578) );
  AOI211_X1 U15176 ( .C1(n13560), .C2(n13559), .A(n15681), .B(n13578), .ZN(
        n13561) );
  AOI211_X1 U15177 ( .C1(n15704), .C2(n7561), .A(n13562), .B(n13561), .ZN(
        n13568) );
  AOI21_X1 U15178 ( .B1(n13565), .B2(n13814), .A(n13586), .ZN(n13566) );
  OR2_X1 U15179 ( .A1(n13566), .A2(n15677), .ZN(n13567) );
  OAI211_X1 U15180 ( .C1(n13569), .C2(n15718), .A(n13568), .B(n13567), .ZN(
        P3_U3199) );
  NOR2_X1 U15181 ( .A1(n7561), .A2(n13570), .ZN(n13572) );
  NAND2_X1 U15182 ( .A1(n13588), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13595) );
  OAI21_X1 U15183 ( .B1(n13588), .B2(P3_REG1_REG_18__SCAN_IN), .A(n13595), 
        .ZN(n13573) );
  AOI21_X1 U15184 ( .B1(n13574), .B2(n13573), .A(n13596), .ZN(n13594) );
  OAI21_X1 U15185 ( .B1(n13577), .B2(n13576), .A(n13575), .ZN(n13584) );
  MUX2_X1 U15186 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13087), .Z(n13582) );
  XNOR2_X1 U15187 ( .A(n13600), .B(n13599), .ZN(n13581) );
  NOR2_X1 U15188 ( .A1(n13581), .A2(n13582), .ZN(n13598) );
  AOI211_X1 U15189 ( .C1(n15704), .C2(n13599), .A(n13584), .B(n13583), .ZN(
        n13593) );
  NOR2_X1 U15190 ( .A1(n7561), .A2(n13585), .ZN(n13587) );
  NOR2_X1 U15191 ( .A1(n13587), .A2(n13586), .ZN(n13590) );
  NAND2_X1 U15192 ( .A1(n13588), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n13604) );
  OAI21_X1 U15193 ( .B1(n13588), .B2(P3_REG2_REG_18__SCAN_IN), .A(n13604), 
        .ZN(n13589) );
  NOR2_X1 U15194 ( .A1(n13590), .A2(n13589), .ZN(n13606) );
  AOI21_X1 U15195 ( .B1(n13590), .B2(n13589), .A(n13606), .ZN(n13591) );
  OR2_X1 U15196 ( .A1(n13591), .A2(n15677), .ZN(n13592) );
  OAI211_X1 U15197 ( .C1(n13594), .C2(n15718), .A(n13593), .B(n13592), .ZN(
        P3_U3200) );
  XNOR2_X1 U15198 ( .A(n13610), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13601) );
  INV_X1 U15199 ( .A(n13601), .ZN(n13597) );
  AOI21_X1 U15200 ( .B1(n13600), .B2(n13599), .A(n13598), .ZN(n13603) );
  XNOR2_X1 U15201 ( .A(n13610), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13607) );
  MUX2_X1 U15202 ( .A(n13607), .B(n13601), .S(n13087), .Z(n13602) );
  XNOR2_X1 U15203 ( .A(n13603), .B(n13602), .ZN(n13613) );
  INV_X1 U15204 ( .A(n13604), .ZN(n13605) );
  AOI21_X1 U15205 ( .B1(n15702), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n13608), 
        .ZN(n13609) );
  OAI21_X1 U15206 ( .B1(n13611), .B2(n13610), .A(n13609), .ZN(n13612) );
  NAND2_X1 U15207 ( .A1(n13615), .A2(n13802), .ZN(n13624) );
  INV_X1 U15208 ( .A(n13616), .ZN(n13617) );
  NAND2_X1 U15209 ( .A1(n13618), .A2(n13617), .ZN(n15996) );
  NAND3_X1 U15210 ( .A1(n13624), .A2(n15810), .A3(n15996), .ZN(n13620) );
  OAI21_X1 U15211 ( .B1(n15810), .B2(P3_REG2_REG_31__SCAN_IN), .A(n13620), 
        .ZN(n13619) );
  OAI21_X1 U15212 ( .B1(n16003), .B2(n15806), .A(n13619), .ZN(P3_U3202) );
  OAI21_X1 U15213 ( .B1(n15810), .B2(P3_REG2_REG_30__SCAN_IN), .A(n13620), 
        .ZN(n13621) );
  OAI21_X1 U15214 ( .B1(n15995), .B2(n15806), .A(n13621), .ZN(P3_U3203) );
  INV_X1 U15215 ( .A(n13622), .ZN(n13629) );
  NAND2_X1 U15216 ( .A1(n15802), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n13623) );
  OAI211_X1 U15217 ( .C1(n13625), .C2(n15806), .A(n13624), .B(n13623), .ZN(
        n13626) );
  AOI21_X1 U15218 ( .B1(n13627), .B2(n13820), .A(n13626), .ZN(n13628) );
  OAI21_X1 U15219 ( .B1(n13629), .B2(n15802), .A(n13628), .ZN(P3_U3204) );
  OAI22_X1 U15220 ( .A1(n13634), .A2(n13835), .B1(n13663), .B2(n13833), .ZN(
        n13635) );
  NOR2_X1 U15221 ( .A1(n13639), .A2(n7752), .ZN(n13641) );
  NAND2_X1 U15222 ( .A1(n13845), .A2(n13820), .ZN(n13644) );
  AOI22_X1 U15223 ( .A1(n13642), .A2(n13802), .B1(n15802), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13643) );
  OAI211_X1 U15224 ( .C1(n13916), .C2(n15806), .A(n13644), .B(n13643), .ZN(
        n13645) );
  AOI21_X1 U15225 ( .B1(n13844), .B2(n15810), .A(n13645), .ZN(n13646) );
  INV_X1 U15226 ( .A(n13646), .ZN(P3_U3205) );
  XNOR2_X1 U15227 ( .A(n13647), .B(n13649), .ZN(n13850) );
  INV_X1 U15228 ( .A(n13820), .ZN(n13842) );
  OAI21_X1 U15229 ( .B1(n13650), .B2(n13649), .A(n13648), .ZN(n13653) );
  AOI222_X1 U15230 ( .A1(n13756), .A2(n13653), .B1(n13652), .B2(n13742), .C1(
        n13651), .C2(n13759), .ZN(n13849) );
  INV_X1 U15231 ( .A(n13849), .ZN(n13658) );
  AOI22_X1 U15232 ( .A1(n13654), .A2(n13802), .B1(n15802), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13655) );
  OAI21_X1 U15233 ( .B1(n13656), .B2(n15806), .A(n13655), .ZN(n13657) );
  AOI21_X1 U15234 ( .B1(n13658), .B2(n15810), .A(n13657), .ZN(n13659) );
  OAI21_X1 U15235 ( .B1(n13850), .B2(n13842), .A(n13659), .ZN(P3_U3206) );
  XOR2_X1 U15236 ( .A(n13665), .B(n13660), .Z(n13661) );
  OAI222_X1 U15237 ( .A1(n13835), .A2(n13663), .B1(n13833), .B2(n13662), .C1(
        n13661), .C2(n13831), .ZN(n13851) );
  INV_X1 U15238 ( .A(n13851), .ZN(n13670) );
  XOR2_X1 U15239 ( .A(n13664), .B(n13665), .Z(n13852) );
  AOI22_X1 U15240 ( .A1(n13666), .A2(n13802), .B1(n15802), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13667) );
  OAI21_X1 U15241 ( .B1(n13921), .B2(n15806), .A(n13667), .ZN(n13668) );
  AOI21_X1 U15242 ( .B1(n13852), .B2(n13820), .A(n13668), .ZN(n13669) );
  OAI21_X1 U15243 ( .B1(n13670), .B2(n15802), .A(n13669), .ZN(P3_U3207) );
  NAND2_X1 U15244 ( .A1(n13671), .A2(n13684), .ZN(n13672) );
  NAND3_X1 U15245 ( .A1(n13673), .A2(n13756), .A3(n13672), .ZN(n13678) );
  OAI22_X1 U15246 ( .A1(n13675), .A2(n13835), .B1(n13674), .B2(n13833), .ZN(
        n13676) );
  INV_X1 U15247 ( .A(n13676), .ZN(n13677) );
  AND2_X1 U15248 ( .A1(n13678), .A2(n13677), .ZN(n13857) );
  INV_X1 U15249 ( .A(n13679), .ZN(n13681) );
  INV_X1 U15250 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n13680) );
  OAI22_X1 U15251 ( .A1(n13681), .A2(n15804), .B1(n15810), .B2(n13680), .ZN(
        n13682) );
  AOI21_X1 U15252 ( .B1(n13683), .B2(n13816), .A(n13682), .ZN(n13688) );
  INV_X1 U15253 ( .A(n13684), .ZN(n13685) );
  XNOR2_X1 U15254 ( .A(n13686), .B(n13685), .ZN(n13855) );
  NAND2_X1 U15255 ( .A1(n13855), .A2(n13820), .ZN(n13687) );
  OAI211_X1 U15256 ( .C1(n13857), .C2(n15802), .A(n13688), .B(n13687), .ZN(
        P3_U3208) );
  XNOR2_X1 U15257 ( .A(n13689), .B(n13693), .ZN(n13928) );
  AOI22_X1 U15258 ( .A1(n13691), .A2(n13742), .B1(n13690), .B2(n13759), .ZN(
        n13696) );
  XNOR2_X1 U15259 ( .A(n13692), .B(n13693), .ZN(n13694) );
  NAND2_X1 U15260 ( .A1(n13694), .A2(n13756), .ZN(n13695) );
  OAI211_X1 U15261 ( .C1(n13928), .C2(n13880), .A(n13696), .B(n13695), .ZN(
        n13926) );
  MUX2_X1 U15262 ( .A(n13926), .B(P3_REG2_REG_24__SCAN_IN), .S(n15802), .Z(
        n13697) );
  INV_X1 U15263 ( .A(n13697), .ZN(n13701) );
  AOI22_X1 U15264 ( .A1(n13699), .A2(n13816), .B1(n13802), .B2(n13698), .ZN(
        n13700) );
  OAI211_X1 U15265 ( .C1(n13928), .C2(n13702), .A(n13701), .B(n13700), .ZN(
        P3_U3209) );
  NAND2_X1 U15266 ( .A1(n13740), .A2(n13704), .ZN(n13706) );
  AND2_X1 U15267 ( .A1(n13706), .A2(n13705), .ZN(n13707) );
  XNOR2_X1 U15268 ( .A(n13707), .B(n13719), .ZN(n13712) );
  NAND2_X1 U15269 ( .A1(n13708), .A2(n13742), .ZN(n13709) );
  OAI21_X1 U15270 ( .B1(n13710), .B2(n13833), .A(n13709), .ZN(n13711) );
  AOI21_X1 U15271 ( .B1(n13712), .B2(n13756), .A(n13711), .ZN(n13865) );
  INV_X1 U15272 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13715) );
  INV_X1 U15273 ( .A(n13713), .ZN(n13714) );
  OAI22_X1 U15274 ( .A1(n15810), .A2(n13715), .B1(n13714), .B2(n15804), .ZN(
        n13716) );
  AOI21_X1 U15275 ( .B1(n13933), .B2(n13816), .A(n13716), .ZN(n13722) );
  NAND2_X1 U15276 ( .A1(n13748), .A2(n13717), .ZN(n13729) );
  NAND2_X1 U15277 ( .A1(n13731), .A2(n13718), .ZN(n13720) );
  OR2_X1 U15278 ( .A1(n13720), .A2(n13719), .ZN(n13863) );
  NAND3_X1 U15279 ( .A1(n13863), .A2(n13862), .A3(n13820), .ZN(n13721) );
  OAI211_X1 U15280 ( .C1(n13865), .C2(n15802), .A(n13722), .B(n13721), .ZN(
        P3_U3210) );
  NAND2_X1 U15281 ( .A1(n13740), .A2(n13745), .ZN(n13739) );
  NAND2_X1 U15282 ( .A1(n13739), .A2(n13723), .ZN(n13725) );
  XNOR2_X1 U15283 ( .A(n13725), .B(n13724), .ZN(n13726) );
  OAI222_X1 U15284 ( .A1(n13835), .A2(n13727), .B1(n13833), .B2(n13763), .C1(
        n13726), .C2(n13831), .ZN(n13868) );
  INV_X1 U15285 ( .A(n13868), .ZN(n13738) );
  NAND2_X1 U15286 ( .A1(n13729), .A2(n13728), .ZN(n13730) );
  NAND2_X1 U15287 ( .A1(n13731), .A2(n13730), .ZN(n13938) );
  INV_X1 U15288 ( .A(n13938), .ZN(n13736) );
  AOI22_X1 U15289 ( .A1(n15802), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n13802), 
        .B2(n13732), .ZN(n13733) );
  OAI21_X1 U15290 ( .B1(n13734), .B2(n15806), .A(n13733), .ZN(n13735) );
  AOI21_X1 U15291 ( .B1(n13736), .B2(n13820), .A(n13735), .ZN(n13737) );
  OAI21_X1 U15292 ( .B1(n13738), .B2(n15802), .A(n13737), .ZN(P3_U3211) );
  OAI21_X1 U15293 ( .B1(n13740), .B2(n13745), .A(n13739), .ZN(n13744) );
  AOI222_X1 U15294 ( .A1(n13756), .A2(n13744), .B1(n13743), .B2(n13742), .C1(
        n13741), .C2(n13759), .ZN(n13876) );
  NAND2_X1 U15295 ( .A1(n13746), .A2(n13745), .ZN(n13747) );
  NAND2_X1 U15296 ( .A1(n13748), .A2(n13747), .ZN(n13874) );
  INV_X1 U15297 ( .A(n13873), .ZN(n13751) );
  AOI22_X1 U15298 ( .A1(n15802), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13802), 
        .B2(n13749), .ZN(n13750) );
  OAI21_X1 U15299 ( .B1(n13751), .B2(n15806), .A(n13750), .ZN(n13752) );
  AOI21_X1 U15300 ( .B1(n13874), .B2(n13820), .A(n13752), .ZN(n13753) );
  OAI21_X1 U15301 ( .B1(n13876), .B2(n15802), .A(n13753), .ZN(P3_U3212) );
  INV_X1 U15302 ( .A(n13754), .ZN(n13758) );
  OAI211_X1 U15303 ( .C1(n13758), .C2(n13757), .A(n13756), .B(n13755), .ZN(
        n13762) );
  NAND2_X1 U15304 ( .A1(n13760), .A2(n13759), .ZN(n13761) );
  OAI211_X1 U15305 ( .C1(n13763), .C2(n13835), .A(n13762), .B(n13761), .ZN(
        n13882) );
  INV_X1 U15306 ( .A(n13882), .ZN(n13773) );
  NAND2_X1 U15307 ( .A1(n13764), .A2(n13767), .ZN(n13947) );
  INV_X1 U15308 ( .A(n13947), .ZN(n13771) );
  AOI22_X1 U15309 ( .A1(n15802), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n13802), 
        .B2(n13768), .ZN(n13769) );
  OAI21_X1 U15310 ( .B1(n13879), .B2(n15806), .A(n13769), .ZN(n13770) );
  AOI21_X1 U15311 ( .B1(n13771), .B2(n13820), .A(n13770), .ZN(n13772) );
  OAI21_X1 U15312 ( .B1(n13773), .B2(n15802), .A(n13772), .ZN(P3_U3213) );
  XOR2_X1 U15313 ( .A(n13781), .B(n13774), .Z(n13775) );
  OAI222_X1 U15314 ( .A1(n13835), .A2(n13776), .B1(n13833), .B2(n13808), .C1(
        n13831), .C2(n13775), .ZN(n13888) );
  NAND2_X1 U15315 ( .A1(n13819), .A2(n13777), .ZN(n13780) );
  NAND2_X1 U15316 ( .A1(n13780), .A2(n13778), .ZN(n13889) );
  INV_X1 U15317 ( .A(n13889), .ZN(n13783) );
  NAND2_X1 U15318 ( .A1(n13780), .A2(n13779), .ZN(n13782) );
  AND2_X1 U15319 ( .A1(n13782), .A2(n13781), .ZN(n13887) );
  NOR3_X1 U15320 ( .A1(n13783), .A2(n13887), .A3(n13842), .ZN(n13788) );
  INV_X1 U15321 ( .A(n13784), .ZN(n13951) );
  AOI22_X1 U15322 ( .A1(n15802), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13802), 
        .B2(n13785), .ZN(n13786) );
  OAI21_X1 U15323 ( .B1(n13951), .B2(n15806), .A(n13786), .ZN(n13787) );
  AOI211_X1 U15324 ( .C1(n13888), .C2(n15810), .A(n13788), .B(n13787), .ZN(
        n13789) );
  INV_X1 U15325 ( .A(n13789), .ZN(P3_U3214) );
  NAND2_X1 U15326 ( .A1(n13819), .A2(n13818), .ZN(n13791) );
  NAND2_X1 U15327 ( .A1(n13791), .A2(n13790), .ZN(n13793) );
  INV_X1 U15328 ( .A(n13795), .ZN(n13792) );
  XNOR2_X1 U15329 ( .A(n13793), .B(n13792), .ZN(n13894) );
  INV_X1 U15330 ( .A(n13894), .ZN(n13806) );
  INV_X1 U15331 ( .A(n13794), .ZN(n13798) );
  AOI21_X1 U15332 ( .B1(n13811), .B2(n13796), .A(n13795), .ZN(n13797) );
  NOR2_X1 U15333 ( .A1(n13798), .A2(n13797), .ZN(n13799) );
  OAI222_X1 U15334 ( .A1(n13835), .A2(n13800), .B1(n13833), .B2(n13834), .C1(
        n13831), .C2(n13799), .ZN(n13893) );
  AOI22_X1 U15335 ( .A1(n15802), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n13802), 
        .B2(n13801), .ZN(n13803) );
  OAI21_X1 U15336 ( .B1(n13955), .B2(n15806), .A(n13803), .ZN(n13804) );
  AOI21_X1 U15337 ( .B1(n13893), .B2(n15810), .A(n13804), .ZN(n13805) );
  OAI21_X1 U15338 ( .B1(n13842), .B2(n13806), .A(n13805), .ZN(P3_U3215) );
  AOI21_X1 U15339 ( .B1(n13807), .B2(n13818), .A(n13831), .ZN(n13812) );
  OAI22_X1 U15340 ( .A1(n13809), .A2(n13833), .B1(n13808), .B2(n13835), .ZN(
        n13810) );
  AOI21_X1 U15341 ( .B1(n13812), .B2(n13811), .A(n13810), .ZN(n13899) );
  OAI22_X1 U15342 ( .A1(n15810), .A2(n13814), .B1(n13813), .B2(n15804), .ZN(
        n13815) );
  AOI21_X1 U15343 ( .B1(n13817), .B2(n13816), .A(n13815), .ZN(n13822) );
  XNOR2_X1 U15344 ( .A(n13819), .B(n13818), .ZN(n13897) );
  NAND2_X1 U15345 ( .A1(n13897), .A2(n13820), .ZN(n13821) );
  OAI211_X1 U15346 ( .C1(n13899), .C2(n15802), .A(n13822), .B(n13821), .ZN(
        P3_U3216) );
  NAND2_X1 U15347 ( .A1(n13824), .A2(n13823), .ZN(n13825) );
  XNOR2_X1 U15348 ( .A(n13825), .B(n13829), .ZN(n13902) );
  INV_X1 U15349 ( .A(n13902), .ZN(n13843) );
  INV_X1 U15350 ( .A(n13826), .ZN(n13827) );
  AOI21_X1 U15351 ( .B1(n13829), .B2(n13828), .A(n13827), .ZN(n13830) );
  OAI222_X1 U15352 ( .A1(n13835), .A2(n13834), .B1(n13833), .B2(n13832), .C1(
        n13831), .C2(n13830), .ZN(n13901) );
  INV_X1 U15353 ( .A(n13836), .ZN(n13961) );
  NOR2_X1 U15354 ( .A1(n13961), .A2(n15806), .ZN(n13840) );
  OAI22_X1 U15355 ( .A1(n15810), .A2(n13838), .B1(n13837), .B2(n15804), .ZN(
        n13839) );
  AOI211_X1 U15356 ( .C1(n13901), .C2(n15810), .A(n13840), .B(n13839), .ZN(
        n13841) );
  OAI21_X1 U15357 ( .B1(n13843), .B2(n13842), .A(n13841), .ZN(P3_U3217) );
  INV_X1 U15358 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13846) );
  OAI21_X1 U15359 ( .B1(n13916), .B2(n13905), .A(n13847), .ZN(P3_U3487) );
  INV_X1 U15360 ( .A(n15917), .ZN(n13886) );
  NAND2_X1 U15361 ( .A1(n8647), .A2(n15865), .ZN(n13848) );
  OAI211_X1 U15362 ( .C1(n13886), .C2(n13850), .A(n13849), .B(n13848), .ZN(
        n13917) );
  MUX2_X1 U15363 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13917), .S(n15997), .Z(
        P3_U3486) );
  INV_X1 U15364 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13853) );
  AOI21_X1 U15365 ( .B1(n15917), .B2(n13852), .A(n13851), .ZN(n13918) );
  MUX2_X1 U15366 ( .A(n13853), .B(n13918), .S(n15997), .Z(n13854) );
  OAI21_X1 U15367 ( .B1(n13921), .B2(n13905), .A(n13854), .ZN(P3_U3485) );
  NAND2_X1 U15368 ( .A1(n13855), .A2(n15917), .ZN(n13856) );
  AND2_X1 U15369 ( .A1(n13857), .A2(n13856), .ZN(n13923) );
  INV_X1 U15370 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13858) );
  MUX2_X1 U15371 ( .A(n13923), .B(n13858), .S(n16004), .Z(n13859) );
  OAI21_X1 U15372 ( .B1(n13925), .B2(n13905), .A(n13859), .ZN(P3_U3484) );
  MUX2_X1 U15373 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13926), .S(n15997), .Z(
        n13861) );
  OAI22_X1 U15374 ( .A1(n13928), .A2(n13885), .B1(n13927), .B2(n13905), .ZN(
        n13860) );
  NAND3_X1 U15375 ( .A1(n13863), .A2(n13862), .A3(n15917), .ZN(n13864) );
  NAND2_X1 U15376 ( .A1(n13865), .A2(n13864), .ZN(n13931) );
  MUX2_X1 U15377 ( .A(n13931), .B(P3_REG1_REG_23__SCAN_IN), .S(n16004), .Z(
        n13866) );
  AOI21_X1 U15378 ( .B1(n16005), .B2(n13933), .A(n13866), .ZN(n13867) );
  INV_X1 U15379 ( .A(n13867), .ZN(P3_U3482) );
  INV_X1 U15380 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13871) );
  NOR2_X1 U15381 ( .A1(n13938), .A2(n13880), .ZN(n13869) );
  AOI211_X1 U15382 ( .C1(n15865), .C2(n13870), .A(n13869), .B(n13868), .ZN(
        n13935) );
  MUX2_X1 U15383 ( .A(n13871), .B(n13935), .S(n15997), .Z(n13872) );
  OAI21_X1 U15384 ( .B1(n13938), .B2(n13885), .A(n13872), .ZN(P3_U3481) );
  INV_X1 U15385 ( .A(n13874), .ZN(n13942) );
  INV_X1 U15386 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13877) );
  AOI22_X1 U15387 ( .A1(n13874), .A2(n15769), .B1(n15865), .B2(n13873), .ZN(
        n13875) );
  AND2_X1 U15388 ( .A1(n13876), .A2(n13875), .ZN(n13939) );
  MUX2_X1 U15389 ( .A(n13877), .B(n13939), .S(n15997), .Z(n13878) );
  OAI21_X1 U15390 ( .B1(n13942), .B2(n13885), .A(n13878), .ZN(P3_U3480) );
  OAI22_X1 U15391 ( .A1(n13947), .A2(n13880), .B1(n13879), .B2(n15912), .ZN(
        n13881) );
  NOR2_X1 U15392 ( .A1(n13882), .A2(n13881), .ZN(n13944) );
  INV_X1 U15393 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13883) );
  MUX2_X1 U15394 ( .A(n13944), .B(n13883), .S(n16004), .Z(n13884) );
  OAI21_X1 U15395 ( .B1(n13947), .B2(n13885), .A(n13884), .ZN(P3_U3479) );
  NOR2_X1 U15396 ( .A1(n13887), .A2(n13886), .ZN(n13890) );
  AOI21_X1 U15397 ( .B1(n13890), .B2(n13889), .A(n13888), .ZN(n13948) );
  MUX2_X1 U15398 ( .A(n13891), .B(n13948), .S(n15997), .Z(n13892) );
  OAI21_X1 U15399 ( .B1(n13951), .B2(n13905), .A(n13892), .ZN(P3_U3478) );
  AOI21_X1 U15400 ( .B1(n13894), .B2(n15917), .A(n13893), .ZN(n13952) );
  MUX2_X1 U15401 ( .A(n13895), .B(n13952), .S(n15997), .Z(n13896) );
  OAI21_X1 U15402 ( .B1(n13955), .B2(n13905), .A(n13896), .ZN(P3_U3477) );
  NAND2_X1 U15403 ( .A1(n13897), .A2(n15917), .ZN(n13898) );
  OAI211_X1 U15404 ( .C1(n15912), .C2(n13900), .A(n13899), .B(n13898), .ZN(
        n13956) );
  MUX2_X1 U15405 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13956), .S(n15997), .Z(
        P3_U3476) );
  AOI21_X1 U15406 ( .B1(n15917), .B2(n13902), .A(n13901), .ZN(n13957) );
  MUX2_X1 U15407 ( .A(n13903), .B(n13957), .S(n15997), .Z(n13904) );
  OAI21_X1 U15408 ( .B1(n13961), .B2(n13905), .A(n13904), .ZN(P3_U3475) );
  AOI22_X1 U15409 ( .A1(n13907), .A2(n15917), .B1(n13906), .B2(n15865), .ZN(
        n13908) );
  NAND2_X1 U15410 ( .A1(n13909), .A2(n13908), .ZN(n13962) );
  MUX2_X1 U15411 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13962), .S(n15997), .Z(
        P3_U3474) );
  NAND2_X1 U15412 ( .A1(n13910), .A2(n15917), .ZN(n13911) );
  OAI211_X1 U15413 ( .C1(n15912), .C2(n13913), .A(n13912), .B(n13911), .ZN(
        n13963) );
  MUX2_X1 U15414 ( .A(P3_REG1_REG_14__SCAN_IN), .B(n13963), .S(n15997), .Z(
        P3_U3473) );
  MUX2_X1 U15415 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13917), .S(n16000), .Z(
        P3_U3454) );
  MUX2_X1 U15416 ( .A(n13919), .B(n13918), .S(n16000), .Z(n13920) );
  OAI21_X1 U15417 ( .B1(n13921), .B2(n13960), .A(n13920), .ZN(P3_U3453) );
  MUX2_X1 U15418 ( .A(n13923), .B(n13922), .S(n16008), .Z(n13924) );
  OAI21_X1 U15419 ( .B1(n13925), .B2(n13960), .A(n13924), .ZN(P3_U3452) );
  MUX2_X1 U15420 ( .A(n13926), .B(P3_REG0_REG_24__SCAN_IN), .S(n16008), .Z(
        n13930) );
  OAI22_X1 U15421 ( .A1(n13928), .A2(n13946), .B1(n13927), .B2(n13960), .ZN(
        n13929) );
  MUX2_X1 U15422 ( .A(n13931), .B(P3_REG0_REG_23__SCAN_IN), .S(n16008), .Z(
        n13932) );
  AOI21_X1 U15423 ( .B1(n16009), .B2(n13933), .A(n13932), .ZN(n13934) );
  INV_X1 U15424 ( .A(n13934), .ZN(P3_U3450) );
  MUX2_X1 U15425 ( .A(n13936), .B(n13935), .S(n16000), .Z(n13937) );
  OAI21_X1 U15426 ( .B1(n13938), .B2(n13946), .A(n13937), .ZN(P3_U3449) );
  INV_X1 U15427 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13940) );
  MUX2_X1 U15428 ( .A(n13940), .B(n13939), .S(n16000), .Z(n13941) );
  OAI21_X1 U15429 ( .B1(n13942), .B2(n13946), .A(n13941), .ZN(P3_U3448) );
  MUX2_X1 U15430 ( .A(n13944), .B(n13943), .S(n16008), .Z(n13945) );
  OAI21_X1 U15431 ( .B1(n13947), .B2(n13946), .A(n13945), .ZN(P3_U3447) );
  MUX2_X1 U15432 ( .A(n13949), .B(n13948), .S(n16000), .Z(n13950) );
  OAI21_X1 U15433 ( .B1(n13951), .B2(n13960), .A(n13950), .ZN(P3_U3446) );
  MUX2_X1 U15434 ( .A(n13953), .B(n13952), .S(n16000), .Z(n13954) );
  OAI21_X1 U15435 ( .B1(n13955), .B2(n13960), .A(n13954), .ZN(P3_U3444) );
  MUX2_X1 U15436 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13956), .S(n16000), .Z(
        P3_U3441) );
  INV_X1 U15437 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13958) );
  MUX2_X1 U15438 ( .A(n13958), .B(n13957), .S(n16000), .Z(n13959) );
  OAI21_X1 U15439 ( .B1(n13961), .B2(n13960), .A(n13959), .ZN(P3_U3438) );
  MUX2_X1 U15440 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13962), .S(n16000), .Z(
        P3_U3435) );
  MUX2_X1 U15441 ( .A(P3_REG0_REG_14__SCAN_IN), .B(n13963), .S(n16000), .Z(
        P3_U3432) );
  MUX2_X1 U15442 ( .A(n13965), .B(P3_D_REG_1__SCAN_IN), .S(n13964), .Z(
        P3_U3377) );
  MUX2_X1 U15443 ( .A(P3_D_REG_0__SCAN_IN), .B(n9744), .S(n13966), .Z(P3_U3376) );
  INV_X1 U15444 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13968) );
  NAND3_X1 U15445 ( .A1(n13968), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13971) );
  OAI22_X1 U15446 ( .A1(n13967), .A2(n13971), .B1(n13970), .B2(n13969), .ZN(
        n13972) );
  AOI21_X1 U15447 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n13975) );
  INV_X1 U15448 ( .A(n13975), .ZN(P3_U3264) );
  INV_X1 U15449 ( .A(n13976), .ZN(n13979) );
  OAI222_X1 U15450 ( .A1(n13157), .A2(n13979), .B1(n13978), .B2(P3_U3151), 
        .C1(n13977), .C2(n13983), .ZN(P3_U3266) );
  INV_X1 U15451 ( .A(n13980), .ZN(n13981) );
  OAI222_X1 U15452 ( .A1(P3_U3151), .A2(n7186), .B1(n13983), .B2(n13982), .C1(
        n13157), .C2(n13981), .ZN(P3_U3267) );
  MUX2_X1 U15453 ( .A(n13984), .B(n8719), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3271) );
  OAI211_X1 U15454 ( .C1(n13987), .C2(n13986), .A(n13985), .B(n14054), .ZN(
        n13993) );
  OAI22_X1 U15455 ( .A1(n13988), .A2(n14322), .B1(n14019), .B2(n14320), .ZN(
        n14179) );
  INV_X1 U15456 ( .A(n14181), .ZN(n13990) );
  OAI22_X1 U15457 ( .A1(n13990), .A2(n14030), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13989), .ZN(n13991) );
  AOI21_X1 U15458 ( .B1(n14179), .B2(n14023), .A(n13991), .ZN(n13992) );
  OAI211_X1 U15459 ( .C1(n14183), .C2(n14044), .A(n13993), .B(n13992), .ZN(
        P2_U3186) );
  NAND2_X1 U15460 ( .A1(n13994), .A2(n14252), .ZN(n13998) );
  NAND2_X1 U15461 ( .A1(n13995), .A2(n14054), .ZN(n13997) );
  MUX2_X1 U15462 ( .A(n13998), .B(n13997), .S(n13996), .Z(n14005) );
  INV_X1 U15463 ( .A(n13999), .ZN(n14245) );
  AND2_X1 U15464 ( .A1(n14065), .A2(n14353), .ZN(n14000) );
  AOI21_X1 U15465 ( .B1(n14064), .B2(n14355), .A(n14000), .ZN(n14238) );
  OAI22_X1 U15466 ( .A1(n14238), .A2(n14002), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14001), .ZN(n14003) );
  AOI21_X1 U15467 ( .B1(n14245), .B2(n14046), .A(n14003), .ZN(n14004) );
  OAI211_X1 U15468 ( .C1(n9407), .C2(n14044), .A(n14005), .B(n14004), .ZN(
        P2_U3188) );
  OAI211_X1 U15469 ( .C1(n14008), .C2(n14007), .A(n14006), .B(n14054), .ZN(
        n14013) );
  OAI22_X1 U15470 ( .A1(n14009), .A2(n14322), .B1(n14302), .B2(n14320), .ZN(
        n14264) );
  AOI22_X1 U15471 ( .A1(n14264), .A2(n14023), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14010) );
  OAI21_X1 U15472 ( .B1(n14269), .B2(n14030), .A(n14010), .ZN(n14011) );
  AOI21_X1 U15473 ( .B1(n14413), .B2(n14035), .A(n14011), .ZN(n14012) );
  NAND2_X1 U15474 ( .A1(n14013), .A2(n14012), .ZN(P2_U3195) );
  NOR3_X1 U15475 ( .A1(n14014), .A2(n14018), .A3(n14038), .ZN(n14017) );
  AOI21_X1 U15476 ( .B1(n14026), .B2(n14015), .A(n10844), .ZN(n14016) );
  OAI21_X1 U15477 ( .B1(n14017), .B2(n14016), .A(n7531), .ZN(n14025) );
  OAI22_X1 U15478 ( .A1(n14019), .A2(n14322), .B1(n14018), .B2(n14320), .ZN(
        n14202) );
  INV_X1 U15479 ( .A(n14210), .ZN(n14021) );
  OAI22_X1 U15480 ( .A1(n14021), .A2(n14030), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14020), .ZN(n14022) );
  AOI21_X1 U15481 ( .B1(n14202), .B2(n14023), .A(n14022), .ZN(n14024) );
  OAI211_X1 U15482 ( .C1(n14213), .C2(n14044), .A(n14025), .B(n14024), .ZN(
        P2_U3197) );
  OAI211_X1 U15483 ( .C1(n14028), .C2(n14027), .A(n14026), .B(n14054), .ZN(
        n14037) );
  OAI22_X1 U15484 ( .A1(n14030), .A2(n14226), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14029), .ZN(n14034) );
  INV_X1 U15485 ( .A(n14221), .ZN(n14039) );
  OAI22_X1 U15486 ( .A1(n14039), .A2(n14050), .B1(n14032), .B2(n14031), .ZN(
        n14033) );
  AOI211_X1 U15487 ( .C1(n14396), .C2(n14035), .A(n14034), .B(n14033), .ZN(
        n14036) );
  NAND2_X1 U15488 ( .A1(n14037), .A2(n14036), .ZN(P2_U3201) );
  NOR3_X1 U15489 ( .A1(n14040), .A2(n14039), .A3(n14038), .ZN(n14041) );
  AOI21_X1 U15490 ( .B1(n14042), .B2(n14054), .A(n14041), .ZN(n14058) );
  INV_X1 U15491 ( .A(n14043), .ZN(n14057) );
  NOR2_X1 U15492 ( .A1(n14194), .A2(n14044), .ZN(n14053) );
  INV_X1 U15493 ( .A(n14045), .ZN(n14192) );
  AOI22_X1 U15494 ( .A1(n14192), .A2(n14046), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14049) );
  NAND2_X1 U15495 ( .A1(n14221), .A2(n14047), .ZN(n14048) );
  OAI211_X1 U15496 ( .C1(n14051), .C2(n14050), .A(n14049), .B(n14048), .ZN(
        n14052) );
  AOI211_X1 U15497 ( .C1(n14055), .C2(n14054), .A(n14053), .B(n14052), .ZN(
        n14056) );
  OAI21_X1 U15498 ( .B1(n14058), .B2(n14057), .A(n14056), .ZN(P2_U3212) );
  INV_X2 U15499 ( .A(P2_U3947), .ZN(n14082) );
  MUX2_X1 U15500 ( .A(n14059), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14082), .Z(
        P2_U3562) );
  MUX2_X1 U15501 ( .A(n14060), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14082), .Z(
        P2_U3561) );
  MUX2_X1 U15502 ( .A(n14061), .B(P2_DATAO_REG_29__SCAN_IN), .S(n14082), .Z(
        P2_U3560) );
  MUX2_X1 U15503 ( .A(n14062), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14082), .Z(
        P2_U3559) );
  MUX2_X1 U15504 ( .A(n14190), .B(P2_DATAO_REG_27__SCAN_IN), .S(n14082), .Z(
        P2_U3558) );
  MUX2_X1 U15505 ( .A(n14063), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14082), .Z(
        P2_U3557) );
  MUX2_X1 U15506 ( .A(n14221), .B(P2_DATAO_REG_25__SCAN_IN), .S(n14082), .Z(
        P2_U3556) );
  MUX2_X1 U15507 ( .A(n14064), .B(P2_DATAO_REG_24__SCAN_IN), .S(n14082), .Z(
        P2_U3555) );
  MUX2_X1 U15508 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14065), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15509 ( .A(n14251), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14082), .Z(
        P2_U3552) );
  MUX2_X1 U15510 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n14066), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15511 ( .A(n14067), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14082), .Z(
        P2_U3550) );
  MUX2_X1 U15512 ( .A(n14356), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14082), .Z(
        P2_U3549) );
  MUX2_X1 U15513 ( .A(n14068), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14082), .Z(
        P2_U3548) );
  MUX2_X1 U15514 ( .A(n14354), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14082), .Z(
        P2_U3547) );
  MUX2_X1 U15515 ( .A(n14069), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14082), .Z(
        P2_U3546) );
  MUX2_X1 U15516 ( .A(n14070), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14082), .Z(
        P2_U3545) );
  MUX2_X1 U15517 ( .A(n14071), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14082), .Z(
        P2_U3543) );
  MUX2_X1 U15518 ( .A(n14072), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14082), .Z(
        P2_U3542) );
  MUX2_X1 U15519 ( .A(n14073), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14082), .Z(
        P2_U3541) );
  MUX2_X1 U15520 ( .A(n14074), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14082), .Z(
        P2_U3540) );
  MUX2_X1 U15521 ( .A(n14075), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14082), .Z(
        P2_U3539) );
  MUX2_X1 U15522 ( .A(n14076), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14082), .Z(
        P2_U3538) );
  MUX2_X1 U15523 ( .A(n14077), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14082), .Z(
        P2_U3537) );
  MUX2_X1 U15524 ( .A(n14078), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14082), .Z(
        P2_U3536) );
  MUX2_X1 U15525 ( .A(n14079), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14082), .Z(
        P2_U3535) );
  MUX2_X1 U15526 ( .A(n14080), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14082), .Z(
        P2_U3534) );
  MUX2_X1 U15527 ( .A(n14081), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14082), .Z(
        P2_U3533) );
  MUX2_X1 U15528 ( .A(n9000), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14082), .Z(
        P2_U3532) );
  MUX2_X1 U15529 ( .A(n9450), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14082), .Z(
        P2_U3531) );
  INV_X1 U15530 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14085) );
  NOR2_X1 U15531 ( .A1(n14085), .A2(n14086), .ZN(n14099) );
  AOI211_X1 U15532 ( .C1(n14086), .C2(n14085), .A(n14099), .B(n15588), .ZN(
        n14096) );
  OAI211_X1 U15533 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14090), .A(n15583), 
        .B(n14105), .ZN(n14094) );
  INV_X1 U15534 ( .A(n14091), .ZN(n14092) );
  AOI21_X1 U15535 ( .B1(n15522), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n14092), 
        .ZN(n14093) );
  OAI211_X1 U15536 ( .C1(n14148), .C2(n14097), .A(n14094), .B(n14093), .ZN(
        n14095) );
  OR2_X1 U15537 ( .A1(n14096), .A2(n14095), .ZN(P2_U3229) );
  NOR2_X1 U15538 ( .A1(n14098), .A2(n14097), .ZN(n14100) );
  NOR2_X1 U15539 ( .A1(n14100), .A2(n14099), .ZN(n14102) );
  XNOR2_X1 U15540 ( .A(n14127), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14101) );
  NOR2_X1 U15541 ( .A1(n14102), .A2(n14101), .ZN(n14126) );
  AOI211_X1 U15542 ( .C1(n14102), .C2(n14101), .A(n15588), .B(n14126), .ZN(
        n14115) );
  NAND2_X1 U15543 ( .A1(n14104), .A2(n14103), .ZN(n14106) );
  NAND2_X1 U15544 ( .A1(n14117), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14107) );
  OAI21_X1 U15545 ( .B1(n14117), .B2(P2_REG2_REG_16__SCAN_IN), .A(n14107), 
        .ZN(n14108) );
  OAI211_X1 U15546 ( .C1(n14109), .C2(n14108), .A(n14116), .B(n15583), .ZN(
        n14113) );
  INV_X1 U15547 ( .A(n14110), .ZN(n14111) );
  AOI21_X1 U15548 ( .B1(n15522), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n14111), 
        .ZN(n14112) );
  OAI211_X1 U15549 ( .C1(n14148), .C2(n14117), .A(n14113), .B(n14112), .ZN(
        n14114) );
  OR2_X1 U15550 ( .A1(n14115), .A2(n14114), .ZN(P2_U3230) );
  NAND2_X1 U15551 ( .A1(n15567), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14121) );
  INV_X1 U15552 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14118) );
  INV_X1 U15553 ( .A(n14121), .ZN(n14119) );
  AOI21_X1 U15554 ( .B1(n9178), .B2(n14120), .A(n14119), .ZN(n15569) );
  NAND2_X1 U15555 ( .A1(n15570), .A2(n15569), .ZN(n15568) );
  NAND2_X1 U15556 ( .A1(n14121), .A2(n15568), .ZN(n14123) );
  INV_X1 U15557 ( .A(n14123), .ZN(n14124) );
  OAI21_X1 U15558 ( .B1(n14124), .B2(n14129), .A(n14141), .ZN(n14125) );
  AOI21_X1 U15559 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14125), .A(n14143), 
        .ZN(n14134) );
  AOI21_X1 U15560 ( .B1(n14127), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14126), 
        .ZN(n15564) );
  XNOR2_X1 U15561 ( .A(n15567), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15563) );
  NAND2_X1 U15562 ( .A1(n14128), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n14137) );
  OAI211_X1 U15563 ( .C1(n14128), .C2(P2_REG1_REG_18__SCAN_IN), .A(n14137), 
        .B(n15581), .ZN(n14133) );
  NOR2_X1 U15564 ( .A1(n14148), .A2(n14129), .ZN(n14130) );
  AOI211_X1 U15565 ( .C1(n15522), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n14131), 
        .B(n14130), .ZN(n14132) );
  OAI211_X1 U15566 ( .C1(n14134), .C2(n15592), .A(n14133), .B(n14132), .ZN(
        P2_U3232) );
  INV_X1 U15567 ( .A(n14135), .ZN(n14136) );
  NAND2_X1 U15568 ( .A1(n14137), .A2(n14136), .ZN(n14139) );
  XNOR2_X1 U15569 ( .A(n9722), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14138) );
  XNOR2_X1 U15570 ( .A(n14139), .B(n14138), .ZN(n14151) );
  MUX2_X1 U15571 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n14310), .S(n14140), .Z(
        n14145) );
  INV_X1 U15572 ( .A(n14141), .ZN(n14142) );
  NOR2_X1 U15573 ( .A1(n14143), .A2(n14142), .ZN(n14144) );
  NAND2_X1 U15574 ( .A1(n15522), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n14147) );
  OAI211_X1 U15575 ( .C1(n14148), .C2(n9722), .A(n14147), .B(n14146), .ZN(
        n14149) );
  OAI21_X1 U15576 ( .B1(n14151), .B2(n15588), .A(n14150), .ZN(P2_U3233) );
  XNOR2_X1 U15577 ( .A(n14157), .B(n14365), .ZN(n14367) );
  NOR2_X1 U15578 ( .A1(n14153), .A2(n14152), .ZN(n14368) );
  INV_X1 U15579 ( .A(n14368), .ZN(n14154) );
  NOR2_X1 U15580 ( .A1(n14359), .A2(n14154), .ZN(n14161) );
  AOI21_X1 U15581 ( .B1(n14359), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14161), 
        .ZN(n14156) );
  NAND2_X1 U15582 ( .A1(n14365), .A2(n14271), .ZN(n14155) );
  OAI211_X1 U15583 ( .C1(n14367), .C2(n14163), .A(n14156), .B(n14155), .ZN(
        P2_U3234) );
  OAI21_X1 U15584 ( .B1(n14159), .B2(n14158), .A(n14157), .ZN(n14371) );
  NOR2_X1 U15585 ( .A1(n14159), .A2(n14349), .ZN(n14160) );
  AOI211_X1 U15586 ( .C1(n14359), .C2(P2_REG2_REG_30__SCAN_IN), .A(n14161), 
        .B(n14160), .ZN(n14162) );
  OAI21_X1 U15587 ( .B1(n14163), .B2(n14371), .A(n14162), .ZN(P2_U3235) );
  AOI21_X1 U15588 ( .B1(n14167), .B2(n14165), .A(n14164), .ZN(n14376) );
  INV_X1 U15589 ( .A(n14170), .ZN(n14171) );
  AOI211_X1 U15590 ( .C1(n14373), .C2(n7245), .A(n15821), .B(n14171), .ZN(
        n14372) );
  NAND2_X1 U15591 ( .A1(n14372), .A2(n9722), .ZN(n14172) );
  OAI211_X1 U15592 ( .C1(n14308), .C2(n14173), .A(n14375), .B(n14172), .ZN(
        n14174) );
  NAND2_X1 U15593 ( .A1(n14174), .A2(n14311), .ZN(n14176) );
  AOI22_X1 U15594 ( .A1(n14373), .A2(n14271), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14359), .ZN(n14175) );
  OAI211_X1 U15595 ( .C1(n14364), .C2(n14376), .A(n14176), .B(n14175), .ZN(
        P2_U3237) );
  XNOR2_X1 U15596 ( .A(n14178), .B(n14177), .ZN(n14180) );
  AOI21_X1 U15597 ( .B1(n14180), .B2(n14358), .A(n14179), .ZN(n14383) );
  XNOR2_X1 U15598 ( .A(n14183), .B(n14191), .ZN(n14378) );
  AOI22_X1 U15599 ( .A1(n14181), .A2(n14345), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14359), .ZN(n14182) );
  OAI21_X1 U15600 ( .B1(n14183), .B2(n14349), .A(n14182), .ZN(n14184) );
  AOI21_X1 U15601 ( .B1(n14378), .B2(n14362), .A(n14184), .ZN(n14188) );
  OR2_X1 U15602 ( .A1(n14186), .A2(n14185), .ZN(n14380) );
  NAND3_X1 U15603 ( .A1(n14380), .A2(n14379), .A3(n14292), .ZN(n14187) );
  OAI211_X1 U15604 ( .C1(n14383), .C2(n14359), .A(n14188), .B(n14187), .ZN(
        P2_U3238) );
  OAI21_X1 U15605 ( .B1(n14209), .B2(n14194), .A(n14191), .ZN(n14384) );
  INV_X1 U15606 ( .A(n14384), .ZN(n14199) );
  AOI22_X1 U15607 ( .A1(n14192), .A2(n14345), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14347), .ZN(n14193) );
  OAI21_X1 U15608 ( .B1(n14194), .B2(n14349), .A(n14193), .ZN(n14198) );
  XNOR2_X1 U15609 ( .A(n14196), .B(n14195), .ZN(n14389) );
  NOR2_X1 U15610 ( .A1(n14389), .A2(n14364), .ZN(n14197) );
  AOI211_X1 U15611 ( .C1(n14199), .C2(n14362), .A(n14198), .B(n14197), .ZN(
        n14200) );
  OAI21_X1 U15612 ( .B1(n14388), .B2(n14347), .A(n14200), .ZN(P2_U3239) );
  XNOR2_X1 U15613 ( .A(n14201), .B(n14205), .ZN(n14203) );
  AOI21_X1 U15614 ( .B1(n14203), .B2(n14358), .A(n14202), .ZN(n14394) );
  OAI21_X1 U15615 ( .B1(n14206), .B2(n14205), .A(n14204), .ZN(n14390) );
  NAND2_X1 U15616 ( .A1(n14225), .A2(n14392), .ZN(n14207) );
  NAND2_X1 U15617 ( .A1(n14207), .A2(n14445), .ZN(n14208) );
  NOR2_X1 U15618 ( .A1(n14209), .A2(n14208), .ZN(n14391) );
  NAND2_X1 U15619 ( .A1(n14391), .A2(n14314), .ZN(n14212) );
  AOI22_X1 U15620 ( .A1(n14210), .A2(n14345), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14347), .ZN(n14211) );
  OAI211_X1 U15621 ( .C1(n14213), .C2(n14349), .A(n14212), .B(n14211), .ZN(
        n14214) );
  AOI21_X1 U15622 ( .B1(n14390), .B2(n14292), .A(n14214), .ZN(n14215) );
  OAI21_X1 U15623 ( .B1(n14394), .B2(n14359), .A(n14215), .ZN(P2_U3240) );
  OAI21_X1 U15624 ( .B1(n14217), .B2(n14220), .A(n14216), .ZN(n14230) );
  AOI21_X1 U15625 ( .B1(n14220), .B2(n14219), .A(n14218), .ZN(n14223) );
  AOI22_X1 U15626 ( .A1(n14221), .A2(n14355), .B1(n14353), .B2(n14252), .ZN(
        n14222) );
  OAI21_X1 U15627 ( .B1(n14223), .B2(n14298), .A(n14222), .ZN(n14224) );
  AOI21_X1 U15628 ( .B1(n14305), .B2(n14230), .A(n14224), .ZN(n14399) );
  AOI21_X1 U15629 ( .B1(n14396), .B2(n7215), .A(n7577), .ZN(n14397) );
  INV_X1 U15630 ( .A(n14396), .ZN(n14229) );
  INV_X1 U15631 ( .A(n14226), .ZN(n14227) );
  AOI22_X1 U15632 ( .A1(n14227), .A2(n14345), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14347), .ZN(n14228) );
  OAI21_X1 U15633 ( .B1(n14229), .B2(n14349), .A(n14228), .ZN(n14233) );
  INV_X1 U15634 ( .A(n14230), .ZN(n14400) );
  NOR2_X1 U15635 ( .A1(n14400), .A2(n14231), .ZN(n14232) );
  AOI211_X1 U15636 ( .C1(n14397), .C2(n14362), .A(n14233), .B(n14232), .ZN(
        n14234) );
  OAI21_X1 U15637 ( .B1(n14399), .B2(n14347), .A(n14234), .ZN(P2_U3241) );
  OAI211_X1 U15638 ( .C1(n14237), .C2(n14236), .A(n14235), .B(n14358), .ZN(
        n14239) );
  OAI21_X1 U15639 ( .B1(n14242), .B2(n14241), .A(n14240), .ZN(n14401) );
  AOI21_X1 U15640 ( .B1(n14403), .B2(n14254), .A(n15821), .ZN(n14244) );
  AND2_X1 U15641 ( .A1(n14244), .A2(n7215), .ZN(n14402) );
  NAND2_X1 U15642 ( .A1(n14402), .A2(n14314), .ZN(n14247) );
  AOI22_X1 U15643 ( .A1(n14245), .A2(n14345), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14359), .ZN(n14246) );
  OAI211_X1 U15644 ( .C1(n9407), .C2(n14349), .A(n14247), .B(n14246), .ZN(
        n14248) );
  AOI21_X1 U15645 ( .B1(n14401), .B2(n14292), .A(n14248), .ZN(n14249) );
  OAI21_X1 U15646 ( .B1(n14405), .B2(n14359), .A(n14249), .ZN(P2_U3242) );
  XNOR2_X1 U15647 ( .A(n14250), .B(n14258), .ZN(n14253) );
  AOI222_X1 U15648 ( .A1(n14358), .A2(n14253), .B1(n14252), .B2(n14355), .C1(
        n14251), .C2(n14353), .ZN(n14410) );
  AOI21_X1 U15649 ( .B1(n14407), .B2(n14274), .A(n14243), .ZN(n14408) );
  AOI22_X1 U15650 ( .A1(n14255), .A2(n14345), .B1(n14347), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n14256) );
  OAI21_X1 U15651 ( .B1(n14257), .B2(n14349), .A(n14256), .ZN(n14261) );
  XNOR2_X1 U15652 ( .A(n14259), .B(n14258), .ZN(n14411) );
  NOR2_X1 U15653 ( .A1(n14411), .A2(n14364), .ZN(n14260) );
  AOI211_X1 U15654 ( .C1(n14408), .C2(n14362), .A(n14261), .B(n14260), .ZN(
        n14262) );
  OAI21_X1 U15655 ( .B1(n14359), .B2(n14410), .A(n14262), .ZN(P2_U3243) );
  XOR2_X1 U15656 ( .A(n14266), .B(n14263), .Z(n14265) );
  AOI21_X1 U15657 ( .B1(n14265), .B2(n14358), .A(n14264), .ZN(n14415) );
  XOR2_X1 U15658 ( .A(n14267), .B(n14266), .Z(n14416) );
  NAND2_X1 U15659 ( .A1(n14347), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n14268) );
  OAI21_X1 U15660 ( .B1(n14308), .B2(n14269), .A(n14268), .ZN(n14270) );
  AOI21_X1 U15661 ( .B1(n14413), .B2(n14271), .A(n14270), .ZN(n14276) );
  OR2_X1 U15662 ( .A1(n14286), .A2(n14272), .ZN(n14273) );
  AND3_X1 U15663 ( .A1(n14274), .A2(n14445), .A3(n14273), .ZN(n14412) );
  NAND2_X1 U15664 ( .A1(n14412), .A2(n14314), .ZN(n14275) );
  OAI211_X1 U15665 ( .C1(n14416), .C2(n14364), .A(n14276), .B(n14275), .ZN(
        n14277) );
  INV_X1 U15666 ( .A(n14277), .ZN(n14278) );
  OAI21_X1 U15667 ( .B1(n14347), .B2(n14415), .A(n14278), .ZN(P2_U3244) );
  XNOR2_X1 U15668 ( .A(n14279), .B(n14282), .ZN(n14281) );
  AOI21_X1 U15669 ( .B1(n14281), .B2(n14358), .A(n14280), .ZN(n14420) );
  XNOR2_X1 U15670 ( .A(n14283), .B(n14282), .ZN(n14421) );
  INV_X1 U15671 ( .A(n14421), .ZN(n14293) );
  NAND2_X1 U15672 ( .A1(n14306), .A2(n14418), .ZN(n14284) );
  NAND2_X1 U15673 ( .A1(n14284), .A2(n14445), .ZN(n14285) );
  NOR2_X1 U15674 ( .A1(n14286), .A2(n14285), .ZN(n14417) );
  NAND2_X1 U15675 ( .A1(n14417), .A2(n14314), .ZN(n14289) );
  AOI22_X1 U15676 ( .A1(n14347), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14287), 
        .B2(n14345), .ZN(n14288) );
  OAI211_X1 U15677 ( .C1(n14290), .C2(n14349), .A(n14289), .B(n14288), .ZN(
        n14291) );
  AOI21_X1 U15678 ( .B1(n14293), .B2(n14292), .A(n14291), .ZN(n14294) );
  OAI21_X1 U15679 ( .B1(n14359), .B2(n14420), .A(n14294), .ZN(P2_U3245) );
  OAI21_X1 U15680 ( .B1(n14296), .B2(n14300), .A(n14295), .ZN(n14422) );
  AOI211_X1 U15681 ( .C1(n14300), .C2(n14299), .A(n14298), .B(n14297), .ZN(
        n14304) );
  OAI22_X1 U15682 ( .A1(n14302), .A2(n14322), .B1(n14301), .B2(n14320), .ZN(
        n14303) );
  AOI211_X1 U15683 ( .C1(n14422), .C2(n14305), .A(n14304), .B(n14303), .ZN(
        n14426) );
  INV_X1 U15684 ( .A(n14306), .ZN(n14307) );
  AOI211_X1 U15685 ( .C1(n14424), .C2(n14329), .A(n15821), .B(n14307), .ZN(
        n14423) );
  NOR2_X1 U15686 ( .A1(n7585), .A2(n14349), .ZN(n14313) );
  OAI22_X1 U15687 ( .A1(n14311), .A2(n14310), .B1(n14309), .B2(n14308), .ZN(
        n14312) );
  AOI211_X1 U15688 ( .C1(n14423), .C2(n14314), .A(n14313), .B(n14312), .ZN(
        n14316) );
  NAND2_X1 U15689 ( .A1(n14422), .A2(n14335), .ZN(n14315) );
  OAI211_X1 U15690 ( .C1(n14426), .C2(n14359), .A(n14316), .B(n14315), .ZN(
        P2_U3246) );
  OAI21_X1 U15691 ( .B1(n14319), .B2(n14318), .A(n14317), .ZN(n14328) );
  OAI22_X1 U15692 ( .A1(n9224), .A2(n14322), .B1(n14321), .B2(n14320), .ZN(
        n14327) );
  OAI21_X1 U15693 ( .B1(n14325), .B2(n14324), .A(n14323), .ZN(n14336) );
  INV_X1 U15694 ( .A(n14336), .ZN(n14432) );
  NOR2_X1 U15695 ( .A1(n14432), .A2(n10019), .ZN(n14326) );
  AOI211_X1 U15696 ( .C1(n14358), .C2(n14328), .A(n14327), .B(n14326), .ZN(
        n14431) );
  AOI21_X1 U15697 ( .B1(n14428), .B2(n14341), .A(n7586), .ZN(n14429) );
  NAND2_X1 U15698 ( .A1(n14429), .A2(n14362), .ZN(n14332) );
  AOI22_X1 U15699 ( .A1(n14347), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14330), 
        .B2(n14345), .ZN(n14331) );
  OAI211_X1 U15700 ( .C1(n14333), .C2(n14349), .A(n14332), .B(n14331), .ZN(
        n14334) );
  AOI21_X1 U15701 ( .B1(n14336), .B2(n14335), .A(n14334), .ZN(n14337) );
  OAI21_X1 U15702 ( .B1(n14431), .B2(n14359), .A(n14337), .ZN(P2_U3247) );
  XNOR2_X1 U15703 ( .A(n14339), .B(n14338), .ZN(n14437) );
  INV_X1 U15704 ( .A(n14340), .ZN(n14343) );
  INV_X1 U15705 ( .A(n14341), .ZN(n14342) );
  AOI21_X1 U15706 ( .B1(n14433), .B2(n14343), .A(n14342), .ZN(n14434) );
  INV_X1 U15707 ( .A(n14344), .ZN(n14346) );
  AOI22_X1 U15708 ( .A1(n14347), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14346), 
        .B2(n14345), .ZN(n14348) );
  OAI21_X1 U15709 ( .B1(n14350), .B2(n14349), .A(n14348), .ZN(n14361) );
  XNOR2_X1 U15710 ( .A(n14352), .B(n14351), .ZN(n14357) );
  AOI222_X1 U15711 ( .A1(n14358), .A2(n14357), .B1(n14356), .B2(n14355), .C1(
        n14354), .C2(n14353), .ZN(n14436) );
  NOR2_X1 U15712 ( .A1(n14436), .A2(n14359), .ZN(n14360) );
  AOI211_X1 U15713 ( .C1(n14434), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14363) );
  OAI21_X1 U15714 ( .B1(n14364), .B2(n14437), .A(n14363), .ZN(P2_U3248) );
  AOI21_X1 U15715 ( .B1(n14365), .B2(n15841), .A(n14368), .ZN(n14366) );
  OAI21_X1 U15716 ( .B1(n14367), .B2(n15821), .A(n14366), .ZN(n14454) );
  MUX2_X1 U15717 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14454), .S(n14451), .Z(
        P2_U3530) );
  AOI21_X1 U15718 ( .B1(n14369), .B2(n15841), .A(n14368), .ZN(n14370) );
  OAI21_X1 U15719 ( .B1(n14371), .B2(n15821), .A(n14370), .ZN(n14455) );
  MUX2_X1 U15720 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14455), .S(n14451), .Z(
        P2_U3529) );
  AOI21_X1 U15721 ( .B1(n15841), .B2(n14373), .A(n14372), .ZN(n14374) );
  MUX2_X1 U15722 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14456), .S(n14451), .Z(
        P2_U3527) );
  AOI22_X1 U15723 ( .A1(n14378), .A2(n14445), .B1(n15841), .B2(n14377), .ZN(
        n14382) );
  NAND3_X1 U15724 ( .A1(n14380), .A2(n14379), .A3(n15860), .ZN(n14381) );
  NAND3_X1 U15725 ( .A1(n14383), .A2(n14382), .A3(n14381), .ZN(n14457) );
  MUX2_X1 U15726 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14457), .S(n14451), .Z(
        P2_U3526) );
  NOR2_X1 U15727 ( .A1(n14384), .A2(n15821), .ZN(n14385) );
  AOI21_X1 U15728 ( .B1(n15841), .B2(n14386), .A(n14385), .ZN(n14387) );
  OAI211_X1 U15729 ( .C1(n14442), .C2(n14389), .A(n14388), .B(n14387), .ZN(
        n14458) );
  MUX2_X1 U15730 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14458), .S(n14451), .Z(
        P2_U3525) );
  INV_X1 U15731 ( .A(n14390), .ZN(n14395) );
  AOI21_X1 U15732 ( .B1(n15841), .B2(n14392), .A(n14391), .ZN(n14393) );
  OAI211_X1 U15733 ( .C1(n14442), .C2(n14395), .A(n14394), .B(n14393), .ZN(
        n14459) );
  MUX2_X1 U15734 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14459), .S(n14451), .Z(
        P2_U3524) );
  AOI22_X1 U15735 ( .A1(n14397), .A2(n14445), .B1(n15841), .B2(n14396), .ZN(
        n14398) );
  OAI211_X1 U15736 ( .C1(n14400), .C2(n14449), .A(n14399), .B(n14398), .ZN(
        n14460) );
  MUX2_X1 U15737 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14460), .S(n14451), .Z(
        P2_U3523) );
  INV_X1 U15738 ( .A(n14401), .ZN(n14406) );
  AOI21_X1 U15739 ( .B1(n15841), .B2(n14403), .A(n14402), .ZN(n14404) );
  OAI211_X1 U15740 ( .C1(n14406), .C2(n14442), .A(n14405), .B(n14404), .ZN(
        n14461) );
  MUX2_X1 U15741 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14461), .S(n14451), .Z(
        P2_U3522) );
  AOI22_X1 U15742 ( .A1(n14408), .A2(n14445), .B1(n15841), .B2(n14407), .ZN(
        n14409) );
  OAI211_X1 U15743 ( .C1(n14411), .C2(n14442), .A(n14410), .B(n14409), .ZN(
        n14462) );
  MUX2_X1 U15744 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14462), .S(n14451), .Z(
        P2_U3521) );
  AOI21_X1 U15745 ( .B1(n15841), .B2(n14413), .A(n14412), .ZN(n14414) );
  OAI211_X1 U15746 ( .C1(n14416), .C2(n14442), .A(n14415), .B(n14414), .ZN(
        n14463) );
  MUX2_X1 U15747 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14463), .S(n14451), .Z(
        P2_U3520) );
  AOI21_X1 U15748 ( .B1(n15841), .B2(n14418), .A(n14417), .ZN(n14419) );
  OAI211_X1 U15749 ( .C1(n14421), .C2(n14442), .A(n14420), .B(n14419), .ZN(
        n14464) );
  MUX2_X1 U15750 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14464), .S(n14451), .Z(
        P2_U3519) );
  INV_X1 U15751 ( .A(n14422), .ZN(n14427) );
  AOI21_X1 U15752 ( .B1(n15841), .B2(n14424), .A(n14423), .ZN(n14425) );
  OAI211_X1 U15753 ( .C1(n14427), .C2(n14449), .A(n14426), .B(n14425), .ZN(
        n14465) );
  MUX2_X1 U15754 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14465), .S(n14451), .Z(
        P2_U3518) );
  AOI22_X1 U15755 ( .A1(n14429), .A2(n14445), .B1(n15841), .B2(n14428), .ZN(
        n14430) );
  OAI211_X1 U15756 ( .C1(n14432), .C2(n14449), .A(n14431), .B(n14430), .ZN(
        n14466) );
  MUX2_X1 U15757 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14466), .S(n14451), .Z(
        P2_U3517) );
  AOI22_X1 U15758 ( .A1(n14434), .A2(n14445), .B1(n15841), .B2(n14433), .ZN(
        n14435) );
  OAI211_X1 U15759 ( .C1(n14437), .C2(n14442), .A(n14436), .B(n14435), .ZN(
        n14467) );
  MUX2_X1 U15760 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14467), .S(n14451), .Z(
        P2_U3516) );
  AOI22_X1 U15761 ( .A1(n14439), .A2(n14445), .B1(n15841), .B2(n14438), .ZN(
        n14440) );
  OAI211_X1 U15762 ( .C1(n14443), .C2(n14442), .A(n14441), .B(n14440), .ZN(
        n14468) );
  MUX2_X1 U15763 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14468), .S(n14451), .Z(
        P2_U3515) );
  AOI22_X1 U15764 ( .A1(n14446), .A2(n14445), .B1(n15841), .B2(n14444), .ZN(
        n14447) );
  OAI211_X1 U15765 ( .C1(n14450), .C2(n14449), .A(n14448), .B(n14447), .ZN(
        n14470) );
  MUX2_X1 U15766 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14470), .S(n14451), .Z(
        P2_U3514) );
  MUX2_X1 U15767 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n14452), .S(n14451), .Z(
        P2_U3502) );
  MUX2_X1 U15768 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n14453), .S(n14451), .Z(
        P2_U3501) );
  MUX2_X1 U15769 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14454), .S(n14469), .Z(
        P2_U3498) );
  MUX2_X1 U15770 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14455), .S(n14469), .Z(
        P2_U3497) );
  MUX2_X1 U15771 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14456), .S(n14469), .Z(
        P2_U3495) );
  MUX2_X1 U15772 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14457), .S(n14469), .Z(
        P2_U3494) );
  MUX2_X1 U15773 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14458), .S(n14469), .Z(
        P2_U3493) );
  MUX2_X1 U15774 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14459), .S(n14469), .Z(
        P2_U3492) );
  MUX2_X1 U15775 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14460), .S(n14469), .Z(
        P2_U3491) );
  MUX2_X1 U15776 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14461), .S(n14469), .Z(
        P2_U3490) );
  MUX2_X1 U15777 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14462), .S(n14469), .Z(
        P2_U3489) );
  MUX2_X1 U15778 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14463), .S(n14469), .Z(
        P2_U3488) );
  MUX2_X1 U15779 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14464), .S(n14469), .Z(
        P2_U3487) );
  MUX2_X1 U15780 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14465), .S(n14469), .Z(
        P2_U3486) );
  MUX2_X1 U15781 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14466), .S(n14469), .Z(
        P2_U3484) );
  MUX2_X1 U15782 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14467), .S(n14469), .Z(
        P2_U3481) );
  MUX2_X1 U15783 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14468), .S(n14469), .Z(
        P2_U3478) );
  MUX2_X1 U15784 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14470), .S(n14469), .Z(
        P2_U3475) );
  INV_X1 U15785 ( .A(n15482), .ZN(n14478) );
  INV_X1 U15786 ( .A(n14471), .ZN(n14473) );
  NOR4_X1 U15787 ( .A1(n14473), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8875), .A4(
        P2_U3088), .ZN(n14474) );
  AOI21_X1 U15788 ( .B1(n14475), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14474), 
        .ZN(n14476) );
  OAI21_X1 U15789 ( .B1(n14478), .B2(n14477), .A(n14476), .ZN(P2_U3296) );
  MUX2_X1 U15790 ( .A(n14480), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15791 ( .A(n15387), .ZN(n15199) );
  OAI22_X1 U15792 ( .A1(n15199), .A2(n14572), .B1(n14734), .B2(n14626), .ZN(
        n14621) );
  NAND2_X1 U15793 ( .A1(n15387), .A2(n14581), .ZN(n14482) );
  OR2_X1 U15794 ( .A1(n14734), .A2(n14572), .ZN(n14481) );
  NAND2_X1 U15795 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  XNOR2_X1 U15796 ( .A(n14483), .B(n14628), .ZN(n14620) );
  XOR2_X1 U15797 ( .A(n14621), .B(n14620), .Z(n14624) );
  NAND2_X1 U15798 ( .A1(n15982), .A2(n14581), .ZN(n14486) );
  NAND2_X1 U15799 ( .A1(n15040), .A2(n14587), .ZN(n14485) );
  NAND2_X1 U15800 ( .A1(n14486), .A2(n14485), .ZN(n14487) );
  XNOR2_X1 U15801 ( .A(n14487), .B(n14584), .ZN(n14490) );
  XNOR2_X1 U15802 ( .A(n14492), .B(n14490), .ZN(n14739) );
  OAI22_X1 U15803 ( .A1(n14489), .A2(n14572), .B1(n14488), .B2(n14626), .ZN(
        n14740) );
  INV_X1 U15804 ( .A(n14490), .ZN(n14491) );
  NAND2_X1 U15805 ( .A1(n14845), .A2(n14581), .ZN(n14494) );
  OR2_X1 U15806 ( .A1(n14748), .A2(n14572), .ZN(n14493) );
  NAND2_X1 U15807 ( .A1(n14494), .A2(n14493), .ZN(n14495) );
  XNOR2_X1 U15808 ( .A(n14495), .B(n14584), .ZN(n14498) );
  INV_X1 U15809 ( .A(n14498), .ZN(n14500) );
  NOR2_X1 U15810 ( .A1(n14748), .A2(n14626), .ZN(n14496) );
  AOI21_X1 U15811 ( .B1(n14845), .B2(n14587), .A(n14496), .ZN(n14497) );
  INV_X1 U15812 ( .A(n14497), .ZN(n14499) );
  AND2_X1 U15813 ( .A1(n14498), .A2(n14497), .ZN(n14501) );
  AOI21_X1 U15814 ( .B1(n14500), .B2(n14499), .A(n14501), .ZN(n14662) );
  NAND2_X1 U15815 ( .A1(n14661), .A2(n14662), .ZN(n14660) );
  INV_X1 U15816 ( .A(n14501), .ZN(n14672) );
  NAND2_X1 U15817 ( .A1(n15445), .A2(n14581), .ZN(n14503) );
  NAND2_X1 U15818 ( .A1(n15038), .A2(n14587), .ZN(n14502) );
  NAND2_X1 U15819 ( .A1(n14503), .A2(n14502), .ZN(n14504) );
  XNOR2_X1 U15820 ( .A(n14504), .B(n14584), .ZN(n14506) );
  AND2_X1 U15821 ( .A1(n15038), .A2(n14563), .ZN(n14505) );
  AOI21_X1 U15822 ( .B1(n15445), .B2(n14587), .A(n14505), .ZN(n14507) );
  NAND2_X1 U15823 ( .A1(n14506), .A2(n14507), .ZN(n14511) );
  INV_X1 U15824 ( .A(n14506), .ZN(n14509) );
  INV_X1 U15825 ( .A(n14507), .ZN(n14508) );
  NAND2_X1 U15826 ( .A1(n14509), .A2(n14508), .ZN(n14510) );
  NAND2_X1 U15827 ( .A1(n14511), .A2(n14510), .ZN(n14671) );
  INV_X1 U15828 ( .A(n14511), .ZN(n14714) );
  NAND2_X1 U15829 ( .A1(n15436), .A2(n14581), .ZN(n14513) );
  NAND2_X1 U15830 ( .A1(n15037), .A2(n14587), .ZN(n14512) );
  NAND2_X1 U15831 ( .A1(n14513), .A2(n14512), .ZN(n14514) );
  XNOR2_X1 U15832 ( .A(n14514), .B(n14584), .ZN(n14516) );
  AND2_X1 U15833 ( .A1(n15037), .A2(n14563), .ZN(n14515) );
  AOI21_X1 U15834 ( .B1(n15436), .B2(n14587), .A(n14515), .ZN(n14517) );
  NAND2_X1 U15835 ( .A1(n14516), .A2(n14517), .ZN(n14521) );
  INV_X1 U15836 ( .A(n14516), .ZN(n14519) );
  INV_X1 U15837 ( .A(n14517), .ZN(n14518) );
  NAND2_X1 U15838 ( .A1(n14519), .A2(n14518), .ZN(n14520) );
  AND2_X1 U15839 ( .A1(n14521), .A2(n14520), .ZN(n14713) );
  NAND2_X1 U15840 ( .A1(n15333), .A2(n14581), .ZN(n14523) );
  NAND2_X1 U15841 ( .A1(n15343), .A2(n14587), .ZN(n14522) );
  NAND2_X1 U15842 ( .A1(n14523), .A2(n14522), .ZN(n14524) );
  XNOR2_X1 U15843 ( .A(n14524), .B(n14628), .ZN(n14525) );
  AOI22_X1 U15844 ( .A1(n15333), .A2(n14587), .B1(n14563), .B2(n15343), .ZN(
        n14526) );
  XNOR2_X1 U15845 ( .A(n14525), .B(n14526), .ZN(n14613) );
  NAND2_X2 U15846 ( .A1(n14612), .A2(n14613), .ZN(n14693) );
  INV_X1 U15847 ( .A(n14525), .ZN(n14527) );
  NAND2_X1 U15848 ( .A1(n14527), .A2(n14526), .ZN(n14692) );
  NAND2_X1 U15849 ( .A1(n15425), .A2(n14581), .ZN(n14529) );
  NAND2_X1 U15850 ( .A1(n15290), .A2(n14587), .ZN(n14528) );
  NAND2_X1 U15851 ( .A1(n14529), .A2(n14528), .ZN(n14530) );
  XNOR2_X1 U15852 ( .A(n14530), .B(n14628), .ZN(n14539) );
  AND2_X1 U15853 ( .A1(n15290), .A2(n14563), .ZN(n14531) );
  AOI21_X1 U15854 ( .B1(n15425), .B2(n14587), .A(n14531), .ZN(n14537) );
  XNOR2_X1 U15855 ( .A(n14539), .B(n14537), .ZN(n14691) );
  NAND2_X1 U15856 ( .A1(n15300), .A2(n14581), .ZN(n14534) );
  NAND2_X1 U15857 ( .A1(n15272), .A2(n14587), .ZN(n14533) );
  NAND2_X1 U15858 ( .A1(n14534), .A2(n14533), .ZN(n14535) );
  XNOR2_X1 U15859 ( .A(n14535), .B(n14628), .ZN(n14544) );
  NOR2_X1 U15860 ( .A1(n14705), .A2(n14626), .ZN(n14536) );
  AOI21_X1 U15861 ( .B1(n15300), .B2(n14587), .A(n14536), .ZN(n14545) );
  XNOR2_X1 U15862 ( .A(n14544), .B(n14545), .ZN(n14640) );
  INV_X1 U15863 ( .A(n14537), .ZN(n14538) );
  NAND2_X1 U15864 ( .A1(n14539), .A2(n14538), .ZN(n14641) );
  OAI22_X1 U15865 ( .A1(n14880), .A2(n14627), .B1(n14881), .B2(n14572), .ZN(
        n14541) );
  XNOR2_X1 U15866 ( .A(n14541), .B(n14584), .ZN(n14555) );
  OR2_X1 U15867 ( .A1(n14880), .A2(n14572), .ZN(n14543) );
  NAND2_X1 U15868 ( .A1(n15291), .A2(n14563), .ZN(n14542) );
  NAND2_X1 U15869 ( .A1(n14543), .A2(n14542), .ZN(n14556) );
  XNOR2_X1 U15870 ( .A(n14555), .B(n14556), .ZN(n14701) );
  INV_X1 U15871 ( .A(n14544), .ZN(n14546) );
  NAND2_X1 U15872 ( .A1(n14546), .A2(n14545), .ZN(n14702) );
  NAND2_X1 U15873 ( .A1(n15409), .A2(n14581), .ZN(n14549) );
  NAND2_X1 U15874 ( .A1(n15271), .A2(n14587), .ZN(n14548) );
  NAND2_X1 U15875 ( .A1(n14549), .A2(n14548), .ZN(n14550) );
  XNOR2_X1 U15876 ( .A(n14550), .B(n14628), .ZN(n14554) );
  NAND2_X1 U15877 ( .A1(n15409), .A2(n14587), .ZN(n14552) );
  NAND2_X1 U15878 ( .A1(n15271), .A2(n14563), .ZN(n14551) );
  NAND2_X1 U15879 ( .A1(n14552), .A2(n14551), .ZN(n14553) );
  NOR2_X1 U15880 ( .A1(n14554), .A2(n14553), .ZN(n14682) );
  AOI21_X1 U15881 ( .B1(n14554), .B2(n14553), .A(n14682), .ZN(n14596) );
  INV_X1 U15882 ( .A(n14555), .ZN(n14557) );
  NAND2_X1 U15883 ( .A1(n14557), .A2(n14556), .ZN(n14597) );
  INV_X1 U15884 ( .A(n14682), .ZN(n14559) );
  NAND2_X1 U15885 ( .A1(n14595), .A2(n14559), .ZN(n14570) );
  NAND2_X1 U15886 ( .A1(n15250), .A2(n14581), .ZN(n14561) );
  NAND2_X1 U15887 ( .A1(n15036), .A2(n11286), .ZN(n14560) );
  NAND2_X1 U15888 ( .A1(n14561), .A2(n14560), .ZN(n14562) );
  XNOR2_X1 U15889 ( .A(n14562), .B(n14584), .ZN(n14565) );
  AND2_X1 U15890 ( .A1(n15036), .A2(n14563), .ZN(n14564) );
  AOI21_X1 U15891 ( .B1(n15250), .B2(n11286), .A(n14564), .ZN(n14566) );
  NAND2_X1 U15892 ( .A1(n14565), .A2(n14566), .ZN(n14571) );
  INV_X1 U15893 ( .A(n14565), .ZN(n14568) );
  INV_X1 U15894 ( .A(n14566), .ZN(n14567) );
  NAND2_X1 U15895 ( .A1(n14568), .A2(n14567), .ZN(n14569) );
  AND2_X1 U15896 ( .A1(n14571), .A2(n14569), .ZN(n14681) );
  NAND2_X1 U15897 ( .A1(n14683), .A2(n14571), .ZN(n14652) );
  OAI22_X1 U15898 ( .A1(n15398), .A2(n14572), .B1(n14733), .B2(n14626), .ZN(
        n14577) );
  NAND2_X1 U15899 ( .A1(n15232), .A2(n14581), .ZN(n14574) );
  OR2_X1 U15900 ( .A1(n14733), .A2(n14572), .ZN(n14573) );
  NAND2_X1 U15901 ( .A1(n14574), .A2(n14573), .ZN(n14575) );
  XNOR2_X1 U15902 ( .A(n14575), .B(n14628), .ZN(n14576) );
  XOR2_X1 U15903 ( .A(n14577), .B(n14576), .Z(n14653) );
  INV_X1 U15904 ( .A(n14576), .ZN(n14579) );
  INV_X1 U15905 ( .A(n14577), .ZN(n14578) );
  NAND2_X1 U15906 ( .A1(n14579), .A2(n14578), .ZN(n14580) );
  NAND2_X1 U15907 ( .A1(n15392), .A2(n14581), .ZN(n14583) );
  OR2_X1 U15908 ( .A1(n15194), .A2(n14572), .ZN(n14582) );
  NAND2_X1 U15909 ( .A1(n14583), .A2(n14582), .ZN(n14585) );
  XNOR2_X1 U15910 ( .A(n14585), .B(n14584), .ZN(n14589) );
  NOR2_X1 U15911 ( .A1(n15194), .A2(n14626), .ZN(n14586) );
  AOI21_X1 U15912 ( .B1(n15392), .B2(n14587), .A(n14586), .ZN(n14588) );
  OR2_X1 U15913 ( .A1(n14589), .A2(n14588), .ZN(n14728) );
  NAND2_X1 U15914 ( .A1(n14589), .A2(n14588), .ZN(n14730) );
  XOR2_X1 U15915 ( .A(n14624), .B(n14625), .Z(n14594) );
  INV_X1 U15916 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14590) );
  OAI22_X1 U15917 ( .A1(n14743), .A2(n15194), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14590), .ZN(n14592) );
  OAI22_X1 U15918 ( .A1(n15196), .A2(n14747), .B1(n14746), .B2(n15200), .ZN(
        n14591) );
  AOI211_X1 U15919 ( .C1(n15387), .C2(n14751), .A(n14592), .B(n14591), .ZN(
        n14593) );
  OAI21_X1 U15920 ( .B1(n14594), .B2(n14753), .A(n14593), .ZN(P1_U3214) );
  AOI21_X1 U15921 ( .B1(n14700), .B2(n14597), .A(n14596), .ZN(n14598) );
  OAI21_X1 U15922 ( .B1(n7807), .B2(n14598), .A(n14716), .ZN(n14603) );
  OAI22_X1 U15923 ( .A1(n14599), .A2(n15195), .B1(n14881), .B2(n15345), .ZN(
        n15264) );
  AOI22_X1 U15924 ( .A1(n15264), .A2(n14694), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14600) );
  OAI21_X1 U15925 ( .B1(n15266), .B2(n14746), .A(n14600), .ZN(n14601) );
  AOI21_X1 U15926 ( .B1(n15409), .B2(n14751), .A(n14601), .ZN(n14602) );
  NAND2_X1 U15927 ( .A1(n14603), .A2(n14602), .ZN(P1_U3216) );
  OAI211_X1 U15928 ( .C1(n14606), .C2(n14605), .A(n14604), .B(n14716), .ZN(
        n14611) );
  AOI22_X1 U15929 ( .A1(n14644), .A2(n15051), .B1(n14667), .B2(n10352), .ZN(
        n14610) );
  NAND2_X1 U15930 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n15091) );
  OAI21_X1 U15931 ( .B1(n14743), .B2(n14607), .A(n15091), .ZN(n14608) );
  AOI21_X1 U15932 ( .B1(n14751), .B2(n14776), .A(n14608), .ZN(n14609) );
  NAND3_X1 U15933 ( .A1(n14611), .A2(n14610), .A3(n14609), .ZN(P1_U3218) );
  OAI21_X1 U15934 ( .B1(n14613), .B2(n14612), .A(n14693), .ZN(n14614) );
  NAND2_X1 U15935 ( .A1(n14614), .A2(n14716), .ZN(n14619) );
  INV_X1 U15936 ( .A(n15329), .ZN(n14617) );
  AND2_X1 U15937 ( .A1(n15037), .A2(n15289), .ZN(n14615) );
  AOI21_X1 U15938 ( .B1(n15290), .B2(n15342), .A(n14615), .ZN(n15430) );
  NAND2_X1 U15939 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15143)
         );
  OAI21_X1 U15940 ( .B1(n15430), .B2(n14665), .A(n15143), .ZN(n14616) );
  AOI21_X1 U15941 ( .B1(n14617), .B2(n14667), .A(n14616), .ZN(n14618) );
  OAI211_X1 U15942 ( .C1(n7975), .C2(n14725), .A(n14619), .B(n14618), .ZN(
        P1_U3219) );
  INV_X1 U15943 ( .A(n14620), .ZN(n14623) );
  INV_X1 U15944 ( .A(n14621), .ZN(n14622) );
  OAI22_X1 U15945 ( .A1(n15177), .A2(n14572), .B1(n15196), .B2(n14626), .ZN(
        n14631) );
  OAI22_X1 U15946 ( .A1(n15177), .A2(n14627), .B1(n15196), .B2(n14572), .ZN(
        n14629) );
  XNOR2_X1 U15947 ( .A(n14629), .B(n14628), .ZN(n14630) );
  XOR2_X1 U15948 ( .A(n14631), .B(n14630), .Z(n14632) );
  INV_X1 U15949 ( .A(n15034), .ZN(n14634) );
  INV_X1 U15950 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n14633) );
  OAI22_X1 U15951 ( .A1(n14747), .A2(n14634), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14633), .ZN(n14637) );
  OAI22_X1 U15952 ( .A1(n14734), .A2(n14743), .B1(n14746), .B2(n14635), .ZN(
        n14636) );
  AOI211_X1 U15953 ( .C1(n15378), .C2(n14751), .A(n14637), .B(n14636), .ZN(
        n14638) );
  OAI21_X1 U15954 ( .B1(n14639), .B2(n14753), .A(n14638), .ZN(P1_U3220) );
  INV_X1 U15955 ( .A(n14703), .ZN(n14643) );
  AOI21_X1 U15956 ( .B1(n14690), .B2(n14641), .A(n14640), .ZN(n14642) );
  OAI21_X1 U15957 ( .B1(n14643), .B2(n14642), .A(n14716), .ZN(n14650) );
  INV_X1 U15958 ( .A(n14743), .ZN(n14722) );
  AOI22_X1 U15959 ( .A1(n15290), .A2(n14722), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14649) );
  AOI22_X1 U15960 ( .A1(n15299), .A2(n14667), .B1(n14644), .B2(n15291), .ZN(
        n14648) );
  NAND2_X1 U15961 ( .A1(n15300), .A2(n15981), .ZN(n15421) );
  INV_X1 U15962 ( .A(n15421), .ZN(n14646) );
  NAND2_X1 U15963 ( .A1(n14646), .A2(n14645), .ZN(n14647) );
  NAND4_X1 U15964 ( .A1(n14650), .A2(n14649), .A3(n14648), .A4(n14647), .ZN(
        P1_U3223) );
  OAI21_X1 U15965 ( .B1(n14653), .B2(n14652), .A(n14651), .ZN(n14654) );
  NAND2_X1 U15966 ( .A1(n14654), .A2(n14716), .ZN(n14659) );
  INV_X1 U15967 ( .A(n15229), .ZN(n14657) );
  AOI22_X1 U15968 ( .A1(n15035), .A2(n15342), .B1(n15289), .B2(n15036), .ZN(
        n15396) );
  OAI22_X1 U15969 ( .A1(n15396), .A2(n14665), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14655), .ZN(n14656) );
  AOI21_X1 U15970 ( .B1(n14657), .B2(n14667), .A(n14656), .ZN(n14658) );
  OAI211_X1 U15971 ( .C1(n15398), .C2(n14725), .A(n14659), .B(n14658), .ZN(
        P1_U3225) );
  OAI21_X1 U15972 ( .B1(n14662), .B2(n14661), .A(n14660), .ZN(n14663) );
  NAND2_X1 U15973 ( .A1(n14663), .A2(n14716), .ZN(n14670) );
  OAI21_X1 U15974 ( .B1(n15449), .B2(n14665), .A(n14664), .ZN(n14666) );
  AOI21_X1 U15975 ( .B1(n14668), .B2(n14667), .A(n14666), .ZN(n14669) );
  OAI211_X1 U15976 ( .C1(n15451), .C2(n14725), .A(n14670), .B(n14669), .ZN(
        P1_U3226) );
  AND3_X1 U15977 ( .A1(n14660), .A2(n14672), .A3(n14671), .ZN(n14673) );
  OAI21_X1 U15978 ( .B1(n14715), .B2(n14673), .A(n14716), .ZN(n14680) );
  INV_X1 U15979 ( .A(n14674), .ZN(n14678) );
  OAI22_X1 U15980 ( .A1(n14676), .A2(n14747), .B1(n14675), .B2(n14746), .ZN(
        n14677) );
  AOI211_X1 U15981 ( .C1(n14722), .C2(n15039), .A(n14678), .B(n14677), .ZN(
        n14679) );
  OAI211_X1 U15982 ( .C1(n7617), .C2(n14725), .A(n14680), .B(n14679), .ZN(
        P1_U3228) );
  NOR3_X1 U15983 ( .A1(n7807), .A2(n14682), .A3(n14681), .ZN(n14685) );
  INV_X1 U15984 ( .A(n14683), .ZN(n14684) );
  OAI21_X1 U15985 ( .B1(n14685), .B2(n14684), .A(n14716), .ZN(n14689) );
  NOR2_X1 U15986 ( .A1(n14743), .A2(n14706), .ZN(n14687) );
  OAI22_X1 U15987 ( .A1(n14733), .A2(n14747), .B1(n14746), .B2(n15247), .ZN(
        n14686) );
  AOI211_X1 U15988 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n14687), 
        .B(n14686), .ZN(n14688) );
  OAI211_X1 U15989 ( .C1(n12667), .C2(n14725), .A(n14689), .B(n14688), .ZN(
        P1_U3229) );
  NAND2_X1 U15990 ( .A1(n14690), .A2(n14716), .ZN(n14699) );
  AOI21_X1 U15991 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(n14698) );
  OAI22_X1 U15992 ( .A1(n14705), .A2(n15195), .B1(n7974), .B2(n15345), .ZN(
        n15424) );
  AOI22_X1 U15993 ( .A1(n15424), .A2(n14694), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14695) );
  OAI21_X1 U15994 ( .B1(n15313), .B2(n14746), .A(n14695), .ZN(n14696) );
  AOI21_X1 U15995 ( .B1(n15425), .B2(n14751), .A(n14696), .ZN(n14697) );
  OAI21_X1 U15996 ( .B1(n14699), .B2(n14698), .A(n14697), .ZN(P1_U3233) );
  NAND2_X1 U15997 ( .A1(n14700), .A2(n14716), .ZN(n14711) );
  AOI21_X1 U15998 ( .B1(n14703), .B2(n14702), .A(n14701), .ZN(n14710) );
  INV_X1 U15999 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14704) );
  OAI22_X1 U16000 ( .A1(n14705), .A2(n14743), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14704), .ZN(n14708) );
  OAI22_X1 U16001 ( .A1(n14706), .A2(n14747), .B1(n14746), .B2(n15278), .ZN(
        n14707) );
  AOI211_X1 U16002 ( .C1(n15414), .C2(n14751), .A(n14708), .B(n14707), .ZN(
        n14709) );
  OAI21_X1 U16003 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(P1_U3235) );
  INV_X1 U16004 ( .A(n14712), .ZN(n14718) );
  NOR3_X1 U16005 ( .A1(n14715), .A2(n14714), .A3(n14713), .ZN(n14717) );
  OAI21_X1 U16006 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(n14724) );
  INV_X1 U16007 ( .A(n14719), .ZN(n14721) );
  OAI22_X1 U16008 ( .A1(n7974), .A2(n14747), .B1(n15352), .B2(n14746), .ZN(
        n14720) );
  AOI211_X1 U16009 ( .C1(n14722), .C2(n15038), .A(n14721), .B(n14720), .ZN(
        n14723) );
  OAI211_X1 U16010 ( .C1(n7615), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        P1_U3238) );
  INV_X1 U16011 ( .A(n14726), .ZN(n14731) );
  AOI21_X1 U16012 ( .B1(n14730), .B2(n14728), .A(n14727), .ZN(n14729) );
  AOI21_X1 U16013 ( .B1(n14731), .B2(n14730), .A(n14729), .ZN(n14738) );
  OAI22_X1 U16014 ( .A1(n14743), .A2(n14733), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14732), .ZN(n14736) );
  OAI22_X1 U16015 ( .A1(n14734), .A2(n14747), .B1(n14746), .B2(n15210), .ZN(
        n14735) );
  AOI211_X1 U16016 ( .C1(n15392), .C2(n14751), .A(n14736), .B(n14735), .ZN(
        n14737) );
  OAI21_X1 U16017 ( .B1(n14738), .B2(n14753), .A(n14737), .ZN(P1_U3240) );
  XNOR2_X1 U16018 ( .A(n14739), .B(n14740), .ZN(n14754) );
  OAI22_X1 U16019 ( .A1(n14743), .A2(n14742), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14741), .ZN(n14750) );
  INV_X1 U16020 ( .A(n14744), .ZN(n14745) );
  OAI22_X1 U16021 ( .A1(n14748), .A2(n14747), .B1(n14746), .B2(n14745), .ZN(
        n14749) );
  AOI211_X1 U16022 ( .C1(n15982), .C2(n14751), .A(n14750), .B(n14749), .ZN(
        n14752) );
  OAI21_X1 U16023 ( .B1(n14754), .B2(n14753), .A(n14752), .ZN(P1_U3241) );
  MUX2_X1 U16024 ( .A(n15035), .B(n15392), .S(n7414), .Z(n14909) );
  INV_X1 U16025 ( .A(n14909), .ZN(n14913) );
  NAND2_X1 U16026 ( .A1(n14759), .A2(n14758), .ZN(n14761) );
  NAND4_X1 U16027 ( .A1(n14768), .A2(n14761), .A3(n14762), .A4(n14760), .ZN(
        n14775) );
  NAND2_X1 U16028 ( .A1(n14763), .A2(n14762), .ZN(n14766) );
  NAND4_X1 U16029 ( .A1(n14766), .A2(n14941), .A3(n14765), .A4(n14764), .ZN(
        n14774) );
  NAND2_X1 U16030 ( .A1(n14768), .A2(n14767), .ZN(n14773) );
  OAI21_X1 U16031 ( .B1(n15053), .B2(n14941), .A(n14769), .ZN(n14771) );
  CLKBUF_X1 U16032 ( .A(n14814), .Z(n14907) );
  MUX2_X1 U16033 ( .A(n14776), .B(n15052), .S(n14907), .Z(n14777) );
  INV_X1 U16034 ( .A(n14780), .ZN(n14781) );
  NAND2_X1 U16035 ( .A1(n7183), .A2(n14781), .ZN(n14782) );
  AOI21_X1 U16036 ( .B1(n15051), .B2(n14941), .A(n14783), .ZN(n14786) );
  AOI21_X1 U16037 ( .B1(n14784), .B2(n14991), .A(n15790), .ZN(n14785) );
  MUX2_X1 U16038 ( .A(n15050), .B(n14787), .S(n14991), .Z(n14791) );
  MUX2_X1 U16039 ( .A(n15050), .B(n14787), .S(n14941), .Z(n14788) );
  INV_X1 U16040 ( .A(n14790), .ZN(n14793) );
  INV_X1 U16041 ( .A(n14791), .ZN(n14792) );
  MUX2_X1 U16042 ( .A(n15049), .B(n15813), .S(n14941), .Z(n14795) );
  MUX2_X1 U16043 ( .A(n15813), .B(n15049), .S(n14941), .Z(n14794) );
  MUX2_X1 U16044 ( .A(n15048), .B(n14796), .S(n14991), .Z(n14800) );
  MUX2_X1 U16045 ( .A(n15048), .B(n14796), .S(n7414), .Z(n14797) );
  NAND2_X1 U16046 ( .A1(n14798), .A2(n14797), .ZN(n14804) );
  INV_X1 U16047 ( .A(n14799), .ZN(n14802) );
  INV_X1 U16048 ( .A(n14800), .ZN(n14801) );
  NAND2_X1 U16049 ( .A1(n14802), .A2(n14801), .ZN(n14803) );
  MUX2_X1 U16050 ( .A(n15047), .B(n15848), .S(n14941), .Z(n14806) );
  MUX2_X1 U16051 ( .A(n15047), .B(n15848), .S(n14991), .Z(n14805) );
  MUX2_X1 U16052 ( .A(n15046), .B(n15872), .S(n14991), .Z(n14811) );
  NAND2_X1 U16053 ( .A1(n14810), .A2(n14811), .ZN(n14809) );
  MUX2_X1 U16054 ( .A(n15046), .B(n15872), .S(n7414), .Z(n14808) );
  INV_X1 U16055 ( .A(n14810), .ZN(n14813) );
  INV_X1 U16056 ( .A(n14811), .ZN(n14812) );
  MUX2_X1 U16057 ( .A(n15045), .B(n14815), .S(n7414), .Z(n14817) );
  MUX2_X1 U16058 ( .A(n15045), .B(n14815), .S(n14991), .Z(n14816) );
  MUX2_X1 U16059 ( .A(n15044), .B(n15922), .S(n14991), .Z(n14821) );
  MUX2_X1 U16060 ( .A(n15044), .B(n15922), .S(n7414), .Z(n14818) );
  NAND2_X1 U16061 ( .A1(n14819), .A2(n14818), .ZN(n14825) );
  INV_X1 U16062 ( .A(n14820), .ZN(n14823) );
  INV_X1 U16063 ( .A(n14821), .ZN(n14822) );
  NAND2_X1 U16064 ( .A1(n14823), .A2(n14822), .ZN(n14824) );
  MUX2_X1 U16065 ( .A(n15043), .B(n15948), .S(n7414), .Z(n14827) );
  MUX2_X1 U16066 ( .A(n15043), .B(n15948), .S(n14991), .Z(n14826) );
  MUX2_X1 U16067 ( .A(n15042), .B(n14828), .S(n14991), .Z(n14832) );
  NAND2_X1 U16068 ( .A1(n14831), .A2(n14832), .ZN(n14830) );
  MUX2_X1 U16069 ( .A(n15042), .B(n14828), .S(n7414), .Z(n14829) );
  NAND2_X1 U16070 ( .A1(n14830), .A2(n14829), .ZN(n14836) );
  INV_X1 U16071 ( .A(n14831), .ZN(n14834) );
  INV_X1 U16072 ( .A(n14832), .ZN(n14833) );
  NAND2_X1 U16073 ( .A1(n14834), .A2(n14833), .ZN(n14835) );
  NAND2_X1 U16074 ( .A1(n14836), .A2(n14835), .ZN(n14839) );
  MUX2_X1 U16075 ( .A(n15041), .B(n15967), .S(n7414), .Z(n14840) );
  NAND2_X1 U16076 ( .A1(n14839), .A2(n14840), .ZN(n14838) );
  MUX2_X1 U16077 ( .A(n15041), .B(n15967), .S(n14991), .Z(n14837) );
  INV_X1 U16078 ( .A(n14839), .ZN(n14842) );
  INV_X1 U16079 ( .A(n14840), .ZN(n14841) );
  MUX2_X1 U16080 ( .A(n15040), .B(n15982), .S(n14991), .Z(n14844) );
  MUX2_X1 U16081 ( .A(n15040), .B(n15982), .S(n7414), .Z(n14843) );
  MUX2_X1 U16082 ( .A(n15039), .B(n14845), .S(n7414), .Z(n14849) );
  NAND2_X1 U16083 ( .A1(n14848), .A2(n14849), .ZN(n14847) );
  MUX2_X1 U16084 ( .A(n15039), .B(n14845), .S(n14991), .Z(n14846) );
  NAND2_X1 U16085 ( .A1(n14847), .A2(n14846), .ZN(n14853) );
  INV_X1 U16086 ( .A(n14848), .ZN(n14851) );
  INV_X1 U16087 ( .A(n14849), .ZN(n14850) );
  NAND2_X1 U16088 ( .A1(n14851), .A2(n14850), .ZN(n14852) );
  MUX2_X1 U16089 ( .A(n15038), .B(n15445), .S(n14991), .Z(n14857) );
  NAND2_X1 U16090 ( .A1(n14856), .A2(n14857), .ZN(n14855) );
  MUX2_X1 U16091 ( .A(n15038), .B(n15445), .S(n7414), .Z(n14854) );
  NAND2_X1 U16092 ( .A1(n14855), .A2(n14854), .ZN(n14861) );
  INV_X1 U16093 ( .A(n14856), .ZN(n14859) );
  INV_X1 U16094 ( .A(n14857), .ZN(n14858) );
  NAND2_X1 U16095 ( .A1(n14859), .A2(n14858), .ZN(n14860) );
  MUX2_X1 U16096 ( .A(n15037), .B(n15436), .S(n7414), .Z(n14863) );
  MUX2_X1 U16097 ( .A(n15037), .B(n15436), .S(n14991), .Z(n14862) );
  MUX2_X1 U16098 ( .A(n15343), .B(n15333), .S(n14991), .Z(n14867) );
  MUX2_X1 U16099 ( .A(n15343), .B(n15333), .S(n7414), .Z(n14864) );
  NAND2_X1 U16100 ( .A1(n14865), .A2(n14864), .ZN(n14871) );
  INV_X1 U16101 ( .A(n14866), .ZN(n14869) );
  INV_X1 U16102 ( .A(n14867), .ZN(n14868) );
  NAND2_X1 U16103 ( .A1(n14869), .A2(n14868), .ZN(n14870) );
  NAND2_X1 U16104 ( .A1(n14871), .A2(n14870), .ZN(n14874) );
  MUX2_X1 U16105 ( .A(n15290), .B(n15425), .S(n7414), .Z(n14875) );
  NAND2_X1 U16106 ( .A1(n14874), .A2(n14875), .ZN(n14873) );
  MUX2_X1 U16107 ( .A(n15290), .B(n15425), .S(n14991), .Z(n14872) );
  INV_X1 U16108 ( .A(n14874), .ZN(n14877) );
  INV_X1 U16109 ( .A(n14875), .ZN(n14876) );
  MUX2_X1 U16110 ( .A(n15272), .B(n15300), .S(n14907), .Z(n14879) );
  MUX2_X1 U16111 ( .A(n15272), .B(n15300), .S(n7414), .Z(n14878) );
  MUX2_X1 U16112 ( .A(n15291), .B(n15414), .S(n7414), .Z(n14886) );
  NAND2_X1 U16113 ( .A1(n14885), .A2(n14886), .ZN(n14884) );
  MUX2_X1 U16114 ( .A(n14881), .B(n14880), .S(n14991), .Z(n14882) );
  INV_X1 U16115 ( .A(n14882), .ZN(n14883) );
  NAND2_X1 U16116 ( .A1(n14884), .A2(n14883), .ZN(n14890) );
  INV_X1 U16117 ( .A(n14885), .ZN(n14888) );
  INV_X1 U16118 ( .A(n14886), .ZN(n14887) );
  NAND2_X1 U16119 ( .A1(n14888), .A2(n14887), .ZN(n14889) );
  NAND2_X1 U16120 ( .A1(n14890), .A2(n14889), .ZN(n14893) );
  MUX2_X1 U16121 ( .A(n15271), .B(n15409), .S(n14907), .Z(n14894) );
  NAND2_X1 U16122 ( .A1(n14893), .A2(n14894), .ZN(n14892) );
  MUX2_X1 U16123 ( .A(n15271), .B(n15409), .S(n7414), .Z(n14891) );
  NAND2_X1 U16124 ( .A1(n14892), .A2(n14891), .ZN(n14898) );
  INV_X1 U16125 ( .A(n14893), .ZN(n14896) );
  INV_X1 U16126 ( .A(n14894), .ZN(n14895) );
  NAND2_X1 U16127 ( .A1(n14896), .A2(n14895), .ZN(n14897) );
  MUX2_X1 U16128 ( .A(n15036), .B(n15250), .S(n7414), .Z(n14900) );
  MUX2_X1 U16129 ( .A(n15036), .B(n15250), .S(n14991), .Z(n14899) );
  INV_X1 U16130 ( .A(n14900), .ZN(n14901) );
  MUX2_X1 U16131 ( .A(n15241), .B(n15232), .S(n14991), .Z(n14903) );
  MUX2_X1 U16132 ( .A(n15241), .B(n15232), .S(n7414), .Z(n14902) );
  INV_X1 U16133 ( .A(n14903), .ZN(n14904) );
  NAND2_X1 U16134 ( .A1(n7185), .A2(n14904), .ZN(n14905) );
  NAND2_X1 U16135 ( .A1(n14906), .A2(n14905), .ZN(n14910) );
  INV_X1 U16136 ( .A(n14910), .ZN(n14912) );
  INV_X1 U16137 ( .A(n15392), .ZN(n15213) );
  MUX2_X1 U16138 ( .A(n15194), .B(n15213), .S(n14907), .Z(n14908) );
  MUX2_X1 U16140 ( .A(n15217), .B(n15387), .S(n14991), .Z(n14915) );
  INV_X1 U16141 ( .A(n14915), .ZN(n14919) );
  INV_X1 U16142 ( .A(n14914), .ZN(n14916) );
  NAND2_X1 U16143 ( .A1(n14916), .A2(n14915), .ZN(n14918) );
  MUX2_X1 U16144 ( .A(n15217), .B(n15387), .S(n7414), .Z(n14917) );
  MUX2_X1 U16145 ( .A(n15196), .B(n15177), .S(n7414), .Z(n14922) );
  MUX2_X1 U16146 ( .A(n15176), .B(n15378), .S(n14907), .Z(n14921) );
  AND2_X1 U16147 ( .A1(n14922), .A2(n14921), .ZN(n15005) );
  OAI21_X1 U16148 ( .B1(n15031), .B2(n15005), .A(n8150), .ZN(n14995) );
  INV_X1 U16149 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14927) );
  NAND2_X1 U16150 ( .A1(n14923), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14926) );
  NAND2_X1 U16151 ( .A1(n14924), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n14925) );
  OAI211_X1 U16152 ( .C1(n14928), .C2(n14927), .A(n14926), .B(n14925), .ZN(
        n15164) );
  OAI21_X1 U16153 ( .B1(n15151), .B2(n7187), .A(n15164), .ZN(n14933) );
  OR2_X1 U16154 ( .A1(n14947), .A2(n7868), .ZN(n14931) );
  MUX2_X1 U16155 ( .A(n14933), .B(n15368), .S(n7414), .Z(n15008) );
  NOR2_X1 U16156 ( .A1(n15008), .A2(n15013), .ZN(n15015) );
  OR2_X1 U16157 ( .A1(n14947), .A2(n15477), .ZN(n14934) );
  INV_X1 U16158 ( .A(n15153), .ZN(n15365) );
  NOR2_X1 U16159 ( .A1(n15365), .A2(n14991), .ZN(n14978) );
  NAND2_X1 U16160 ( .A1(n14755), .A2(n7187), .ZN(n14936) );
  NAND2_X1 U16161 ( .A1(n14937), .A2(n14936), .ZN(n14939) );
  NAND2_X1 U16162 ( .A1(n14939), .A2(n14938), .ZN(n15002) );
  NAND2_X1 U16163 ( .A1(n14940), .A2(n8111), .ZN(n14986) );
  NAND2_X1 U16164 ( .A1(n15002), .A2(n14986), .ZN(n14999) );
  NOR2_X1 U16165 ( .A1(n15153), .A2(n7414), .ZN(n14980) );
  NAND2_X1 U16166 ( .A1(n14980), .A2(n15151), .ZN(n14983) );
  INV_X1 U16167 ( .A(n14983), .ZN(n14942) );
  AOI211_X1 U16168 ( .C1(n14943), .C2(n14978), .A(n14999), .B(n14942), .ZN(
        n15016) );
  XNOR2_X1 U16169 ( .A(n15153), .B(n14943), .ZN(n15003) );
  NAND2_X1 U16170 ( .A1(n14945), .A2(n14944), .ZN(n14949) );
  OR2_X1 U16171 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  XNOR2_X1 U16172 ( .A(n15372), .B(n15034), .ZN(n15180) );
  INV_X1 U16173 ( .A(n15180), .ZN(n14977) );
  NOR4_X1 U16174 ( .A1(n14951), .A2(n14950), .A3(n10525), .A4(n15758), .ZN(
        n14955) );
  NAND4_X1 U16175 ( .A1(n14955), .A2(n14954), .A3(n14953), .A4(n14952), .ZN(
        n14956) );
  NOR4_X1 U16176 ( .A1(n14959), .A2(n14958), .A3(n14957), .A4(n14956), .ZN(
        n14961) );
  NAND4_X1 U16177 ( .A1(n15928), .A2(n14962), .A3(n14961), .A4(n14960), .ZN(
        n14963) );
  NOR3_X1 U16178 ( .A1(n14965), .A2(n14964), .A3(n14963), .ZN(n14969) );
  NAND4_X1 U16179 ( .A1(n14969), .A2(n14968), .A3(n14967), .A4(n14966), .ZN(
        n14970) );
  NOR4_X1 U16180 ( .A1(n15295), .A2(n15340), .A3(n7972), .A4(n14970), .ZN(
        n14971) );
  NAND4_X1 U16181 ( .A1(n15216), .A2(n14971), .A3(n15324), .A4(n15240), .ZN(
        n14972) );
  NOR3_X1 U16182 ( .A1(n14972), .A2(n15224), .A3(n15275), .ZN(n14974) );
  INV_X1 U16183 ( .A(n15191), .ZN(n14973) );
  NAND4_X1 U16184 ( .A1(n14975), .A2(n14974), .A3(n14973), .A4(n15262), .ZN(
        n14976) );
  XNOR2_X1 U16185 ( .A(n14978), .B(n15002), .ZN(n14979) );
  NOR2_X1 U16186 ( .A1(n14979), .A2(n15151), .ZN(n14985) );
  INV_X1 U16187 ( .A(n14980), .ZN(n14981) );
  NAND3_X1 U16188 ( .A1(n14981), .A2(n15151), .A3(n15002), .ZN(n14982) );
  OAI211_X1 U16189 ( .C1(n14983), .C2(n15002), .A(n14986), .B(n14982), .ZN(
        n14984) );
  OAI22_X1 U16190 ( .A1(n14987), .A2(n14986), .B1(n14985), .B2(n14984), .ZN(
        n15000) );
  OAI21_X1 U16191 ( .B1(n15151), .B2(n14988), .A(n15164), .ZN(n14989) );
  INV_X1 U16192 ( .A(n14989), .ZN(n14990) );
  MUX2_X1 U16193 ( .A(n14990), .B(n15146), .S(n14991), .Z(n15009) );
  MUX2_X1 U16194 ( .A(n15034), .B(n15372), .S(n14991), .Z(n14997) );
  INV_X1 U16195 ( .A(n14997), .ZN(n14993) );
  MUX2_X1 U16196 ( .A(n15034), .B(n15372), .S(n7414), .Z(n14996) );
  NOR2_X1 U16197 ( .A1(n14993), .A2(n14996), .ZN(n15023) );
  NAND2_X1 U16198 ( .A1(n14995), .A2(n14994), .ZN(n15033) );
  INV_X1 U16199 ( .A(n14996), .ZN(n14998) );
  NOR2_X1 U16200 ( .A1(n14998), .A2(n14997), .ZN(n15029) );
  INV_X1 U16201 ( .A(n14999), .ZN(n15001) );
  AOI211_X1 U16202 ( .C1(n15001), .C2(n7631), .A(n15013), .B(n15000), .ZN(
        n15028) );
  NOR2_X1 U16203 ( .A1(n15003), .A2(n15002), .ZN(n15007) );
  INV_X1 U16204 ( .A(n15013), .ZN(n15004) );
  OAI211_X1 U16205 ( .C1(n15008), .C2(n15009), .A(n15007), .B(n15004), .ZN(
        n15006) );
  NOR2_X1 U16206 ( .A1(n15006), .A2(n15029), .ZN(n15030) );
  INV_X1 U16207 ( .A(n15030), .ZN(n15026) );
  INV_X1 U16208 ( .A(n15005), .ZN(n15025) );
  INV_X1 U16209 ( .A(n15006), .ZN(n15022) );
  INV_X1 U16210 ( .A(n15007), .ZN(n15011) );
  INV_X1 U16211 ( .A(n15008), .ZN(n15010) );
  INV_X1 U16212 ( .A(n15009), .ZN(n15014) );
  NOR4_X1 U16213 ( .A1(n15011), .A2(n15010), .A3(n15014), .A4(n15013), .ZN(
        n15021) );
  NOR3_X1 U16214 ( .A1(n15012), .A2(n7200), .A3(n15345), .ZN(n15019) );
  OAI21_X1 U16215 ( .B1(n15013), .B2(n10343), .A(P1_B_REG_SCAN_IN), .ZN(n15018) );
  NAND3_X1 U16216 ( .A1(n15016), .A2(n15015), .A3(n15014), .ZN(n15017) );
  OAI21_X1 U16217 ( .B1(n15019), .B2(n15018), .A(n15017), .ZN(n15020) );
  AOI211_X1 U16218 ( .C1(n15023), .C2(n15022), .A(n15021), .B(n15020), .ZN(
        n15024) );
  OAI21_X1 U16219 ( .B1(n15026), .B2(n15025), .A(n15024), .ZN(n15027) );
  NAND3_X1 U16220 ( .A1(n7181), .A2(n15030), .A3(n8150), .ZN(n15032) );
  MUX2_X1 U16221 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15164), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16222 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n15034), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16223 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15176), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16224 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15217), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16225 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15035), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16226 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15241), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16227 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15036), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16228 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n15291), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16229 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15272), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16230 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15290), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16231 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15343), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16232 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15037), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16233 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15038), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16234 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15039), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16235 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15040), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16236 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15041), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16237 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15042), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16238 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n15043), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16239 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n15044), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16240 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n15045), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16241 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n15046), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16242 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n15047), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16243 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n15048), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16244 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n15049), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16245 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n15050), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16246 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n15051), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16247 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n15052), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16248 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n7377), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16249 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n15054), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16250 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n7381), .S(P1_U4016), .Z(
        P1_U3560) );
  INV_X1 U16251 ( .A(n15056), .ZN(n15071) );
  MUX2_X1 U16252 ( .A(n10181), .B(P1_REG2_REG_1__SCAN_IN), .S(n15057), .Z(
        n15059) );
  OAI211_X1 U16253 ( .C1(n15071), .C2(n15059), .A(n15730), .B(n15058), .ZN(
        n15068) );
  AOI22_X1 U16254 ( .A1(n15732), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n15067) );
  OAI211_X1 U16255 ( .C1(n15063), .C2(n15062), .A(n15739), .B(n15061), .ZN(
        n15066) );
  NAND2_X1 U16256 ( .A1(n15741), .A2(n15064), .ZN(n15065) );
  NAND4_X1 U16257 ( .A1(n15068), .A2(n15067), .A3(n15066), .A4(n15065), .ZN(
        P1_U3244) );
  MUX2_X1 U16258 ( .A(n15071), .B(n15070), .S(n7200), .Z(n15073) );
  NAND2_X1 U16259 ( .A1(n15073), .A2(n15072), .ZN(n15075) );
  OAI211_X1 U16260 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n15076), .A(n15075), .B(
        P1_U4016), .ZN(n15746) );
  AOI22_X1 U16261 ( .A1(n15732), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n15090) );
  XNOR2_X1 U16262 ( .A(n15078), .B(n15077), .ZN(n15086) );
  INV_X1 U16263 ( .A(n15079), .ZN(n15080) );
  NAND2_X1 U16264 ( .A1(n15741), .A2(n15080), .ZN(n15085) );
  OAI21_X1 U16265 ( .B1(n15082), .B2(n15081), .A(n15099), .ZN(n15083) );
  OR2_X1 U16266 ( .A1(n15135), .A2(n15083), .ZN(n15084) );
  OAI211_X1 U16267 ( .C1(n15087), .C2(n15086), .A(n15085), .B(n15084), .ZN(
        n15088) );
  INV_X1 U16268 ( .A(n15088), .ZN(n15089) );
  NAND3_X1 U16269 ( .A1(n15746), .A2(n15090), .A3(n15089), .ZN(P1_U3245) );
  INV_X1 U16270 ( .A(n15096), .ZN(n15093) );
  OAI21_X1 U16271 ( .B1(n15145), .B2(n7694), .A(n15091), .ZN(n15092) );
  AOI21_X1 U16272 ( .B1(n15093), .B2(n15741), .A(n15092), .ZN(n15103) );
  OAI211_X1 U16273 ( .C1(n15095), .C2(n15094), .A(n15730), .B(n15726), .ZN(
        n15102) );
  MUX2_X1 U16274 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10330), .S(n15096), .Z(
        n15097) );
  NAND3_X1 U16275 ( .A1(n15099), .A2(n15098), .A3(n15097), .ZN(n15100) );
  NAND3_X1 U16276 ( .A1(n15739), .A2(n15736), .A3(n15100), .ZN(n15101) );
  NAND3_X1 U16277 ( .A1(n15103), .A2(n15102), .A3(n15101), .ZN(P1_U3246) );
  AND3_X1 U16278 ( .A1(n15106), .A2(n15105), .A3(n15104), .ZN(n15107) );
  OAI21_X1 U16279 ( .B1(n15108), .B2(n15107), .A(n15739), .ZN(n15120) );
  OAI21_X1 U16280 ( .B1(n15145), .B2(n15110), .A(n15109), .ZN(n15111) );
  AOI21_X1 U16281 ( .B1(n15112), .B2(n15741), .A(n15111), .ZN(n15119) );
  OR3_X1 U16282 ( .A1(n15115), .A2(n15114), .A3(n15113), .ZN(n15116) );
  NAND3_X1 U16283 ( .A1(n15117), .A2(n15730), .A3(n15116), .ZN(n15118) );
  NAND3_X1 U16284 ( .A1(n15120), .A2(n15119), .A3(n15118), .ZN(P1_U3252) );
  INV_X1 U16285 ( .A(n15121), .ZN(n15122) );
  NAND2_X1 U16286 ( .A1(n15122), .A2(n15129), .ZN(n15123) );
  NAND2_X1 U16287 ( .A1(n15124), .A2(n15123), .ZN(n15126) );
  XNOR2_X1 U16288 ( .A(n15126), .B(n15125), .ZN(n15136) );
  INV_X1 U16289 ( .A(n15127), .ZN(n15128) );
  NAND2_X1 U16290 ( .A1(n15128), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n15132) );
  NAND2_X1 U16291 ( .A1(n15130), .A2(n15129), .ZN(n15131) );
  NAND2_X1 U16292 ( .A1(n15132), .A2(n15131), .ZN(n15133) );
  XOR2_X1 U16293 ( .A(n15133), .B(P1_REG2_REG_19__SCAN_IN), .Z(n15134) );
  AOI22_X1 U16294 ( .A1(n15136), .A2(n15739), .B1(n15730), .B2(n15134), .ZN(
        n15142) );
  INV_X1 U16295 ( .A(n15134), .ZN(n15138) );
  NOR2_X1 U16296 ( .A1(n15136), .A2(n15135), .ZN(n15137) );
  AOI211_X1 U16297 ( .C1(n15139), .C2(n15138), .A(n15741), .B(n15137), .ZN(
        n15141) );
  MUX2_X1 U16298 ( .A(n15142), .B(n15141), .S(n15140), .Z(n15144) );
  OAI211_X1 U16299 ( .C1(n8223), .C2(n15145), .A(n15144), .B(n15143), .ZN(
        P1_U3262) );
  OR2_X2 U16300 ( .A1(n15171), .A2(n15372), .ZN(n15172) );
  XNOR2_X1 U16301 ( .A(n15155), .B(n15153), .ZN(n15147) );
  NAND2_X1 U16302 ( .A1(n15147), .A2(n15932), .ZN(n15364) );
  NOR2_X1 U16303 ( .A1(n15760), .A2(n15148), .ZN(n15152) );
  AND2_X1 U16304 ( .A1(n15149), .A2(P1_B_REG_SCAN_IN), .ZN(n15150) );
  NOR2_X1 U16305 ( .A1(n15195), .A2(n15150), .ZN(n15163) );
  NAND2_X1 U16306 ( .A1(n15151), .A2(n15163), .ZN(n15366) );
  NOR2_X1 U16307 ( .A1(n15366), .A2(n15946), .ZN(n15159) );
  AOI211_X1 U16308 ( .C1(n15153), .C2(n15947), .A(n15152), .B(n15159), .ZN(
        n15154) );
  OAI21_X1 U16309 ( .B1(n15364), .B2(n15358), .A(n15154), .ZN(P1_U3263) );
  INV_X1 U16310 ( .A(n15172), .ZN(n15157) );
  INV_X1 U16311 ( .A(n15155), .ZN(n15156) );
  OAI211_X1 U16312 ( .C1(n15368), .C2(n15157), .A(n15156), .B(n15932), .ZN(
        n15367) );
  NOR2_X1 U16313 ( .A1(n15368), .A2(n15317), .ZN(n15158) );
  AOI211_X1 U16314 ( .C1(n15946), .C2(P1_REG2_REG_30__SCAN_IN), .A(n15159), 
        .B(n15158), .ZN(n15160) );
  OAI21_X1 U16315 ( .B1(n15358), .B2(n15367), .A(n15160), .ZN(P1_U3264) );
  XNOR2_X1 U16316 ( .A(n15162), .B(n14977), .ZN(n15369) );
  INV_X1 U16317 ( .A(n15369), .ZN(n15186) );
  AND2_X1 U16318 ( .A1(n15164), .A2(n15163), .ZN(n15371) );
  INV_X1 U16319 ( .A(n15165), .ZN(n15168) );
  NOR2_X1 U16320 ( .A1(n15755), .A2(n15166), .ZN(n15167) );
  AOI21_X1 U16321 ( .B1(n15371), .B2(n15168), .A(n15167), .ZN(n15169) );
  OAI21_X1 U16322 ( .B1(n15170), .B2(n15760), .A(n15169), .ZN(n15175) );
  AOI21_X1 U16323 ( .B1(n15171), .B2(n15372), .A(n15354), .ZN(n15173) );
  NAND2_X1 U16324 ( .A1(n15173), .A2(n15172), .ZN(n15374) );
  NOR2_X1 U16325 ( .A1(n15374), .A2(n15358), .ZN(n15174) );
  AOI211_X1 U16326 ( .C1(n15947), .C2(n15372), .A(n15175), .B(n15174), .ZN(
        n15185) );
  NOR2_X1 U16327 ( .A1(n15378), .A2(n15196), .ZN(n15178) );
  OAI22_X1 U16328 ( .A1(n15179), .A2(n15178), .B1(n15177), .B2(n15176), .ZN(
        n15181) );
  XNOR2_X1 U16329 ( .A(n15181), .B(n15180), .ZN(n15182) );
  INV_X1 U16330 ( .A(n15376), .ZN(n15183) );
  NOR2_X1 U16331 ( .A1(n15196), .A2(n15345), .ZN(n15370) );
  OAI21_X1 U16332 ( .B1(n15183), .B2(n15370), .A(n15760), .ZN(n15184) );
  OAI211_X1 U16333 ( .C1(n15186), .C2(n15285), .A(n15185), .B(n15184), .ZN(
        P1_U3356) );
  OAI21_X1 U16334 ( .B1(n15188), .B2(n15191), .A(n15187), .ZN(n15385) );
  INV_X1 U16335 ( .A(n15189), .ZN(n15193) );
  NAND3_X1 U16336 ( .A1(n15214), .A2(n15191), .A3(n15190), .ZN(n15192) );
  AOI21_X1 U16337 ( .B1(n15193), .B2(n15192), .A(n15959), .ZN(n15198) );
  OAI22_X1 U16338 ( .A1(n15196), .A2(n15195), .B1(n15194), .B2(n15345), .ZN(
        n15197) );
  AOI211_X1 U16339 ( .C1(n15387), .C2(n15208), .A(n15354), .B(n7224), .ZN(
        n15386) );
  NOR2_X1 U16340 ( .A1(n15199), .A2(n15317), .ZN(n15203) );
  OAI22_X1 U16341 ( .A1(n15760), .A2(n15201), .B1(n15200), .B2(n15755), .ZN(
        n15202) );
  AOI211_X1 U16342 ( .C1(n15386), .C2(n15951), .A(n15203), .B(n15202), .ZN(
        n15205) );
  INV_X1 U16343 ( .A(n15363), .ZN(n15815) );
  NAND2_X1 U16344 ( .A1(n15385), .A2(n15815), .ZN(n15204) );
  OAI211_X1 U16345 ( .C1(n15389), .C2(n15946), .A(n15205), .B(n15204), .ZN(
        P1_U3266) );
  XNOR2_X1 U16346 ( .A(n15207), .B(n15206), .ZN(n15395) );
  INV_X1 U16347 ( .A(n15208), .ZN(n15209) );
  AOI211_X1 U16348 ( .C1(n15392), .C2(n15227), .A(n15354), .B(n15209), .ZN(
        n15391) );
  INV_X1 U16349 ( .A(n15210), .ZN(n15211) );
  AOI22_X1 U16350 ( .A1(n15946), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n15211), 
        .B2(n15944), .ZN(n15212) );
  OAI21_X1 U16351 ( .B1(n15213), .B2(n15317), .A(n15212), .ZN(n15220) );
  OAI21_X1 U16352 ( .B1(n15216), .B2(n15215), .A(n15214), .ZN(n15218) );
  AOI222_X1 U16353 ( .A1(n15988), .A2(n15218), .B1(n15241), .B2(n15289), .C1(
        n15217), .C2(n15342), .ZN(n15394) );
  NOR2_X1 U16354 ( .A1(n15394), .A2(n15946), .ZN(n15219) );
  AOI211_X1 U16355 ( .C1(n15391), .C2(n15951), .A(n15220), .B(n15219), .ZN(
        n15221) );
  OAI21_X1 U16356 ( .B1(n15285), .B2(n15395), .A(n15221), .ZN(P1_U3267) );
  XOR2_X1 U16357 ( .A(n15224), .B(n15222), .Z(n15402) );
  OAI21_X1 U16358 ( .B1(n15225), .B2(n15224), .A(n15223), .ZN(n15226) );
  INV_X1 U16359 ( .A(n15226), .ZN(n15400) );
  OAI211_X1 U16360 ( .C1(n15246), .C2(n15398), .A(n15932), .B(n15227), .ZN(
        n15397) );
  NOR2_X1 U16361 ( .A1(n15760), .A2(n15228), .ZN(n15231) );
  OAI22_X1 U16362 ( .A1(n15396), .A2(n15946), .B1(n15229), .B2(n15755), .ZN(
        n15230) );
  AOI211_X1 U16363 ( .C1(n15232), .C2(n15947), .A(n15231), .B(n15230), .ZN(
        n15233) );
  OAI21_X1 U16364 ( .B1(n15397), .B2(n15358), .A(n15233), .ZN(n15234) );
  AOI21_X1 U16365 ( .B1(n15400), .B2(n15952), .A(n15234), .ZN(n15235) );
  OAI21_X1 U16366 ( .B1(n15402), .B2(n15337), .A(n15235), .ZN(P1_U3268) );
  AND2_X1 U16367 ( .A1(n15236), .A2(n15240), .ZN(n15238) );
  OR2_X1 U16368 ( .A1(n15238), .A2(n15237), .ZN(n15405) );
  OAI211_X1 U16369 ( .C1(n7313), .C2(n15240), .A(n15239), .B(n15988), .ZN(
        n15243) );
  AOI22_X1 U16370 ( .A1(n15241), .A2(n15342), .B1(n15289), .B2(n15271), .ZN(
        n15242) );
  NAND2_X1 U16371 ( .A1(n15243), .A2(n15242), .ZN(n15244) );
  AOI21_X1 U16372 ( .B1(n15405), .B2(n15880), .A(n15244), .ZN(n15407) );
  NOR2_X1 U16373 ( .A1(n15257), .A2(n12667), .ZN(n15245) );
  OR3_X1 U16374 ( .A1(n15246), .A2(n15245), .A3(n15354), .ZN(n15403) );
  OAI22_X1 U16375 ( .A1(n15760), .A2(n15248), .B1(n15247), .B2(n15755), .ZN(
        n15249) );
  AOI21_X1 U16376 ( .B1(n15250), .B2(n15947), .A(n15249), .ZN(n15251) );
  OAI21_X1 U16377 ( .B1(n15403), .B2(n15358), .A(n15251), .ZN(n15252) );
  AOI21_X1 U16378 ( .B1(n15405), .B2(n15815), .A(n15252), .ZN(n15253) );
  OAI21_X1 U16379 ( .B1(n15407), .B2(n15946), .A(n15253), .ZN(P1_U3269) );
  OAI21_X1 U16380 ( .B1(n8149), .B2(n12728), .A(n7412), .ZN(n15412) );
  NAND2_X1 U16381 ( .A1(n15409), .A2(n15282), .ZN(n15255) );
  NAND2_X1 U16382 ( .A1(n15255), .A2(n15932), .ZN(n15256) );
  NOR2_X1 U16383 ( .A1(n15257), .A2(n15256), .ZN(n15408) );
  NAND2_X1 U16384 ( .A1(n15409), .A2(n15947), .ZN(n15258) );
  OAI21_X1 U16385 ( .B1(n15760), .B2(n15259), .A(n15258), .ZN(n15260) );
  AOI21_X1 U16386 ( .B1(n15408), .B2(n15951), .A(n15260), .ZN(n15269) );
  OAI21_X1 U16387 ( .B1(n15263), .B2(n15262), .A(n15261), .ZN(n15265) );
  AOI21_X1 U16388 ( .B1(n15265), .B2(n15988), .A(n15264), .ZN(n15411) );
  OAI21_X1 U16389 ( .B1(n15266), .B2(n15755), .A(n15411), .ZN(n15267) );
  NAND2_X1 U16390 ( .A1(n15267), .A2(n15760), .ZN(n15268) );
  OAI211_X1 U16391 ( .C1(n15412), .C2(n15285), .A(n15269), .B(n15268), .ZN(
        P1_U3270) );
  XNOR2_X1 U16392 ( .A(n15270), .B(n15275), .ZN(n15273) );
  AOI222_X1 U16393 ( .A1(n15988), .A2(n15273), .B1(n15272), .B2(n15289), .C1(
        n15271), .C2(n15342), .ZN(n15416) );
  OAI21_X1 U16394 ( .B1(n15276), .B2(n15275), .A(n15274), .ZN(n15277) );
  INV_X1 U16395 ( .A(n15277), .ZN(n15417) );
  OAI22_X1 U16396 ( .A1(n15760), .A2(n15279), .B1(n15278), .B2(n15755), .ZN(
        n15280) );
  AOI21_X1 U16397 ( .B1(n15414), .B2(n15947), .A(n15280), .ZN(n15284) );
  NAND2_X1 U16398 ( .A1(n15414), .A2(n15297), .ZN(n15281) );
  AND3_X1 U16399 ( .A1(n15282), .A2(n15281), .A3(n15932), .ZN(n15413) );
  NAND2_X1 U16400 ( .A1(n15413), .A2(n15951), .ZN(n15283) );
  OAI211_X1 U16401 ( .C1(n15417), .C2(n15285), .A(n15284), .B(n15283), .ZN(
        n15286) );
  INV_X1 U16402 ( .A(n15286), .ZN(n15287) );
  OAI21_X1 U16403 ( .B1(n15946), .B2(n15416), .A(n15287), .ZN(P1_U3271) );
  XNOR2_X1 U16404 ( .A(n15288), .B(n15295), .ZN(n15292) );
  AOI222_X1 U16405 ( .A1(n15988), .A2(n15292), .B1(n15291), .B2(n15342), .C1(
        n15290), .C2(n15289), .ZN(n15422) );
  AND2_X1 U16406 ( .A1(n15308), .A2(n15293), .ZN(n15296) );
  OAI21_X1 U16407 ( .B1(n15296), .B2(n15295), .A(n15294), .ZN(n15418) );
  OAI211_X1 U16408 ( .C1(n15311), .C2(n15298), .A(n15932), .B(n15297), .ZN(
        n15419) );
  AOI22_X1 U16409 ( .A1(n15299), .A2(n15944), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n15946), .ZN(n15302) );
  NAND2_X1 U16410 ( .A1(n15300), .A2(n15947), .ZN(n15301) );
  OAI211_X1 U16411 ( .C1(n15419), .C2(n15358), .A(n15302), .B(n15301), .ZN(
        n15303) );
  AOI21_X1 U16412 ( .B1(n15418), .B2(n15952), .A(n15303), .ZN(n15304) );
  OAI21_X1 U16413 ( .B1(n15422), .B2(n15946), .A(n15304), .ZN(P1_U3272) );
  INV_X1 U16414 ( .A(n15305), .ZN(n15306) );
  AOI21_X1 U16415 ( .B1(n7972), .B2(n15307), .A(n15306), .ZN(n15426) );
  INV_X1 U16416 ( .A(n15426), .ZN(n15322) );
  OAI21_X1 U16417 ( .B1(n7336), .B2(n7972), .A(n15308), .ZN(n15429) );
  INV_X1 U16418 ( .A(n15429), .ZN(n15320) );
  INV_X1 U16419 ( .A(n15425), .ZN(n15318) );
  NAND2_X1 U16420 ( .A1(n15327), .A2(n15425), .ZN(n15309) );
  NAND2_X1 U16421 ( .A1(n15309), .A2(n15932), .ZN(n15310) );
  NOR2_X1 U16422 ( .A1(n15311), .A2(n15310), .ZN(n15423) );
  NAND2_X1 U16423 ( .A1(n15423), .A2(n15951), .ZN(n15316) );
  INV_X1 U16424 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n15312) );
  OAI22_X1 U16425 ( .A1(n15313), .A2(n15755), .B1(n15312), .B2(n15760), .ZN(
        n15314) );
  AOI21_X1 U16426 ( .B1(n15424), .B2(n15760), .A(n15314), .ZN(n15315) );
  OAI211_X1 U16427 ( .C1(n15318), .C2(n15317), .A(n15316), .B(n15315), .ZN(
        n15319) );
  AOI21_X1 U16428 ( .B1(n15320), .B2(n15952), .A(n15319), .ZN(n15321) );
  OAI21_X1 U16429 ( .B1(n15337), .B2(n15322), .A(n15321), .ZN(P1_U3273) );
  XNOR2_X1 U16430 ( .A(n15323), .B(n15324), .ZN(n15435) );
  XNOR2_X1 U16431 ( .A(n15325), .B(n15324), .ZN(n15433) );
  NAND2_X1 U16432 ( .A1(n15333), .A2(n15356), .ZN(n15326) );
  NAND3_X1 U16433 ( .A1(n15327), .A2(n15932), .A3(n15326), .ZN(n15431) );
  INV_X1 U16434 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15328) );
  OAI22_X1 U16435 ( .A1(n15329), .A2(n15755), .B1(n15328), .B2(n15760), .ZN(
        n15330) );
  INV_X1 U16436 ( .A(n15330), .ZN(n15331) );
  OAI21_X1 U16437 ( .B1(n15430), .B2(n15946), .A(n15331), .ZN(n15332) );
  AOI21_X1 U16438 ( .B1(n15333), .B2(n15947), .A(n15332), .ZN(n15334) );
  OAI21_X1 U16439 ( .B1(n15431), .B2(n15358), .A(n15334), .ZN(n15335) );
  AOI21_X1 U16440 ( .B1(n15433), .B2(n15952), .A(n15335), .ZN(n15336) );
  OAI21_X1 U16441 ( .B1(n15337), .B2(n15435), .A(n15336), .ZN(P1_U3274) );
  XNOR2_X1 U16442 ( .A(n15338), .B(n15340), .ZN(n15439) );
  INV_X1 U16443 ( .A(n15439), .ZN(n15339) );
  NAND2_X1 U16444 ( .A1(n15339), .A2(n15880), .ZN(n15351) );
  AOI21_X1 U16445 ( .B1(n15341), .B2(n15340), .A(n15959), .ZN(n15349) );
  NAND2_X1 U16446 ( .A1(n15343), .A2(n15342), .ZN(n15344) );
  OAI21_X1 U16447 ( .B1(n15346), .B2(n15345), .A(n15344), .ZN(n15347) );
  AOI21_X1 U16448 ( .B1(n15349), .B2(n15348), .A(n15347), .ZN(n15350) );
  NAND2_X1 U16449 ( .A1(n15351), .A2(n15350), .ZN(n15441) );
  NAND2_X1 U16450 ( .A1(n15441), .A2(n15760), .ZN(n15362) );
  OAI22_X1 U16451 ( .A1(n15353), .A2(n15760), .B1(n15352), .B2(n15755), .ZN(
        n15360) );
  AOI21_X1 U16452 ( .B1(n15436), .B2(n15355), .A(n15354), .ZN(n15357) );
  NAND2_X1 U16453 ( .A1(n15357), .A2(n15356), .ZN(n15437) );
  NOR2_X1 U16454 ( .A1(n15437), .A2(n15358), .ZN(n15359) );
  AOI211_X1 U16455 ( .C1(n15947), .C2(n15436), .A(n15360), .B(n15359), .ZN(
        n15361) );
  OAI211_X1 U16456 ( .C1(n15439), .C2(n15363), .A(n15362), .B(n15361), .ZN(
        P1_U3275) );
  OAI211_X1 U16457 ( .C1(n15365), .C2(n15970), .A(n15364), .B(n15366), .ZN(
        n15456) );
  MUX2_X1 U16458 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15456), .S(n15991), .Z(
        P1_U3559) );
  MUX2_X1 U16459 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15457), .S(n15991), .Z(
        P1_U3557) );
  NAND2_X1 U16460 ( .A1(n15377), .A2(n15973), .ZN(n15382) );
  NAND2_X1 U16461 ( .A1(n15378), .A2(n15981), .ZN(n15379) );
  MUX2_X1 U16462 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15458), .S(n15991), .Z(
        P1_U3556) );
  INV_X1 U16463 ( .A(n15385), .ZN(n15390) );
  AOI21_X1 U16464 ( .B1(n15981), .B2(n15387), .A(n15386), .ZN(n15388) );
  OAI211_X1 U16465 ( .C1(n15390), .C2(n15875), .A(n15389), .B(n15388), .ZN(
        n15459) );
  MUX2_X1 U16466 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15459), .S(n15991), .Z(
        P1_U3555) );
  AOI21_X1 U16467 ( .B1(n15981), .B2(n15392), .A(n15391), .ZN(n15393) );
  OAI211_X1 U16468 ( .C1(n15395), .C2(n15985), .A(n15394), .B(n15393), .ZN(
        n15460) );
  MUX2_X1 U16469 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15460), .S(n15991), .Z(
        P1_U3554) );
  OAI211_X1 U16470 ( .C1(n15398), .C2(n15970), .A(n15397), .B(n15396), .ZN(
        n15399) );
  AOI21_X1 U16471 ( .B1(n15400), .B2(n15973), .A(n15399), .ZN(n15401) );
  OAI21_X1 U16472 ( .B1(n15959), .B2(n15402), .A(n15401), .ZN(n15461) );
  MUX2_X1 U16473 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15461), .S(n15991), .Z(
        P1_U3553) );
  OAI21_X1 U16474 ( .B1(n12667), .B2(n15970), .A(n15403), .ZN(n15404) );
  AOI21_X1 U16475 ( .B1(n15405), .B2(n15779), .A(n15404), .ZN(n15406) );
  NAND2_X1 U16476 ( .A1(n15407), .A2(n15406), .ZN(n15462) );
  MUX2_X1 U16477 ( .A(n15462), .B(P1_REG1_REG_24__SCAN_IN), .S(n15990), .Z(
        P1_U3552) );
  AOI21_X1 U16478 ( .B1(n15981), .B2(n15409), .A(n15408), .ZN(n15410) );
  OAI211_X1 U16479 ( .C1(n15412), .C2(n15985), .A(n15411), .B(n15410), .ZN(
        n15463) );
  MUX2_X1 U16480 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15463), .S(n15991), .Z(
        P1_U3551) );
  AOI21_X1 U16481 ( .B1(n15981), .B2(n15414), .A(n15413), .ZN(n15415) );
  OAI211_X1 U16482 ( .C1(n15985), .C2(n15417), .A(n15416), .B(n15415), .ZN(
        n15464) );
  MUX2_X1 U16483 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15464), .S(n15991), .Z(
        P1_U3550) );
  NAND2_X1 U16484 ( .A1(n15418), .A2(n15973), .ZN(n15420) );
  NAND4_X1 U16485 ( .A1(n15422), .A2(n15421), .A3(n15420), .A4(n15419), .ZN(
        n15465) );
  MUX2_X1 U16486 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15465), .S(n15991), .Z(
        P1_U3549) );
  AOI211_X1 U16487 ( .C1(n15981), .C2(n15425), .A(n15424), .B(n15423), .ZN(
        n15428) );
  NAND2_X1 U16488 ( .A1(n15426), .A2(n15988), .ZN(n15427) );
  OAI211_X1 U16489 ( .C1(n15429), .C2(n15985), .A(n15428), .B(n15427), .ZN(
        n15466) );
  MUX2_X1 U16490 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15466), .S(n15991), .Z(
        P1_U3548) );
  OAI211_X1 U16491 ( .C1(n7975), .C2(n15970), .A(n15431), .B(n15430), .ZN(
        n15432) );
  AOI21_X1 U16492 ( .B1(n15433), .B2(n15973), .A(n15432), .ZN(n15434) );
  OAI21_X1 U16493 ( .B1(n15959), .B2(n15435), .A(n15434), .ZN(n15467) );
  MUX2_X1 U16494 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15467), .S(n15991), .Z(
        P1_U3547) );
  NAND2_X1 U16495 ( .A1(n15436), .A2(n15981), .ZN(n15438) );
  OAI211_X1 U16496 ( .C1(n15439), .C2(n15875), .A(n15438), .B(n15437), .ZN(
        n15440) );
  MUX2_X1 U16497 ( .A(n15468), .B(P1_REG1_REG_18__SCAN_IN), .S(n15990), .Z(
        P1_U3546) );
  NAND3_X1 U16498 ( .A1(n12720), .A2(n15973), .A3(n15442), .ZN(n15447) );
  AOI211_X1 U16499 ( .C1(n15981), .C2(n15445), .A(n15444), .B(n15443), .ZN(
        n15446) );
  OAI211_X1 U16500 ( .C1(n15959), .C2(n15448), .A(n15447), .B(n15446), .ZN(
        n15469) );
  MUX2_X1 U16501 ( .A(n15469), .B(P1_REG1_REG_17__SCAN_IN), .S(n15990), .Z(
        P1_U3545) );
  OAI211_X1 U16502 ( .C1(n15451), .C2(n15970), .A(n15450), .B(n15449), .ZN(
        n15452) );
  AOI21_X1 U16503 ( .B1(n15453), .B2(n15988), .A(n15452), .ZN(n15454) );
  OAI21_X1 U16504 ( .B1(n15455), .B2(n15985), .A(n15454), .ZN(n15470) );
  MUX2_X1 U16505 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15470), .S(n15991), .Z(
        P1_U3544) );
  MUX2_X1 U16506 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15456), .S(n15994), .Z(
        P1_U3527) );
  MUX2_X1 U16507 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15457), .S(n15994), .Z(
        P1_U3525) );
  MUX2_X1 U16508 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15458), .S(n15994), .Z(
        P1_U3524) );
  MUX2_X1 U16509 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15459), .S(n15994), .Z(
        P1_U3523) );
  MUX2_X1 U16510 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15460), .S(n15994), .Z(
        P1_U3522) );
  MUX2_X1 U16511 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15461), .S(n15994), .Z(
        P1_U3521) );
  MUX2_X1 U16512 ( .A(n15462), .B(P1_REG0_REG_24__SCAN_IN), .S(n15992), .Z(
        P1_U3520) );
  MUX2_X1 U16513 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15463), .S(n15994), .Z(
        P1_U3519) );
  MUX2_X1 U16514 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15464), .S(n15994), .Z(
        P1_U3518) );
  MUX2_X1 U16515 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15465), .S(n15994), .Z(
        P1_U3517) );
  MUX2_X1 U16516 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15466), .S(n15994), .Z(
        P1_U3516) );
  MUX2_X1 U16517 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15467), .S(n15994), .Z(
        P1_U3515) );
  MUX2_X1 U16518 ( .A(n15468), .B(P1_REG0_REG_18__SCAN_IN), .S(n15992), .Z(
        P1_U3513) );
  MUX2_X1 U16519 ( .A(n15469), .B(P1_REG0_REG_17__SCAN_IN), .S(n15992), .Z(
        P1_U3510) );
  MUX2_X1 U16520 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15470), .S(n15994), .Z(
        P1_U3507) );
  MUX2_X1 U16521 ( .A(P1_D_REG_1__SCAN_IN), .B(n15473), .S(n15517), .Z(
        P1_U3446) );
  MUX2_X1 U16522 ( .A(P1_D_REG_0__SCAN_IN), .B(n15474), .S(n15517), .Z(
        P1_U3445) );
  NAND3_X1 U16523 ( .A1(n15475), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n15478) );
  OAI22_X1 U16524 ( .A1(n15479), .A2(n15478), .B1(n15477), .B2(n15476), .ZN(
        n15480) );
  AOI21_X1 U16525 ( .B1(n15482), .B2(n15481), .A(n15480), .ZN(n15483) );
  INV_X1 U16526 ( .A(n15483), .ZN(P1_U3324) );
  MUX2_X1 U16527 ( .A(n10343), .B(n15484), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16528 ( .A(n15485), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16529 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15486) );
  NOR2_X1 U16530 ( .A1(n15517), .A2(n15486), .ZN(P1_U3323) );
  INV_X1 U16531 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15487) );
  NOR2_X1 U16532 ( .A1(n15517), .A2(n15487), .ZN(P1_U3322) );
  INV_X1 U16533 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15488) );
  NOR2_X1 U16534 ( .A1(n15517), .A2(n15488), .ZN(P1_U3321) );
  INV_X1 U16535 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15489) );
  NOR2_X1 U16536 ( .A1(n15517), .A2(n15489), .ZN(P1_U3320) );
  INV_X1 U16537 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n15490) );
  NOR2_X1 U16538 ( .A1(n15517), .A2(n15490), .ZN(P1_U3319) );
  INV_X1 U16539 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15491) );
  NOR2_X1 U16540 ( .A1(n15517), .A2(n15491), .ZN(P1_U3318) );
  INV_X1 U16541 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15492) );
  NOR2_X1 U16542 ( .A1(n15502), .A2(n15492), .ZN(P1_U3317) );
  INV_X1 U16543 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15493) );
  NOR2_X1 U16544 ( .A1(n15502), .A2(n15493), .ZN(P1_U3316) );
  INV_X1 U16545 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n15494) );
  NOR2_X1 U16546 ( .A1(n15502), .A2(n15494), .ZN(P1_U3315) );
  INV_X1 U16547 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15495) );
  NOR2_X1 U16548 ( .A1(n15502), .A2(n15495), .ZN(P1_U3314) );
  INV_X1 U16549 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15496) );
  NOR2_X1 U16550 ( .A1(n15502), .A2(n15496), .ZN(P1_U3313) );
  INV_X1 U16551 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n15497) );
  NOR2_X1 U16552 ( .A1(n15502), .A2(n15497), .ZN(P1_U3312) );
  INV_X1 U16553 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15498) );
  NOR2_X1 U16554 ( .A1(n15502), .A2(n15498), .ZN(P1_U3311) );
  INV_X1 U16555 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15499) );
  NOR2_X1 U16556 ( .A1(n15502), .A2(n15499), .ZN(P1_U3310) );
  INV_X1 U16557 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15500) );
  NOR2_X1 U16558 ( .A1(n15502), .A2(n15500), .ZN(P1_U3309) );
  INV_X1 U16559 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n15501) );
  NOR2_X1 U16560 ( .A1(n15502), .A2(n15501), .ZN(P1_U3308) );
  INV_X1 U16561 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15503) );
  NOR2_X1 U16562 ( .A1(n15517), .A2(n15503), .ZN(P1_U3307) );
  INV_X1 U16563 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n15504) );
  NOR2_X1 U16564 ( .A1(n15517), .A2(n15504), .ZN(P1_U3306) );
  INV_X1 U16565 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15505) );
  NOR2_X1 U16566 ( .A1(n15517), .A2(n15505), .ZN(P1_U3305) );
  INV_X1 U16567 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15506) );
  NOR2_X1 U16568 ( .A1(n15517), .A2(n15506), .ZN(P1_U3304) );
  INV_X1 U16569 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n15507) );
  NOR2_X1 U16570 ( .A1(n15517), .A2(n15507), .ZN(P1_U3303) );
  INV_X1 U16571 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15508) );
  NOR2_X1 U16572 ( .A1(n15517), .A2(n15508), .ZN(P1_U3302) );
  INV_X1 U16573 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15509) );
  NOR2_X1 U16574 ( .A1(n15517), .A2(n15509), .ZN(P1_U3301) );
  INV_X1 U16575 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15510) );
  NOR2_X1 U16576 ( .A1(n15517), .A2(n15510), .ZN(P1_U3300) );
  INV_X1 U16577 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n15511) );
  NOR2_X1 U16578 ( .A1(n15517), .A2(n15511), .ZN(P1_U3299) );
  INV_X1 U16579 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15512) );
  NOR2_X1 U16580 ( .A1(n15517), .A2(n15512), .ZN(P1_U3298) );
  INV_X1 U16581 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15513) );
  NOR2_X1 U16582 ( .A1(n15517), .A2(n15513), .ZN(P1_U3297) );
  INV_X1 U16583 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15514) );
  NOR2_X1 U16584 ( .A1(n15517), .A2(n15514), .ZN(P1_U3296) );
  INV_X1 U16585 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15515) );
  NOR2_X1 U16586 ( .A1(n15517), .A2(n15515), .ZN(P1_U3295) );
  INV_X1 U16587 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15516) );
  NOR2_X1 U16588 ( .A1(n15517), .A2(n15516), .ZN(P1_U3294) );
  INV_X1 U16589 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U16590 ( .A1(n15526), .A2(n15519), .B1(n15518), .B2(n15523), .ZN(
        P2_U3417) );
  AND2_X1 U16591 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15521), .ZN(P2_U3295) );
  AND2_X1 U16592 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15521), .ZN(P2_U3294) );
  AND2_X1 U16593 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15521), .ZN(P2_U3293) );
  AND2_X1 U16594 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15521), .ZN(P2_U3292) );
  AND2_X1 U16595 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15521), .ZN(P2_U3291) );
  AND2_X1 U16596 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15521), .ZN(P2_U3290) );
  AND2_X1 U16597 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15521), .ZN(P2_U3289) );
  AND2_X1 U16598 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15521), .ZN(P2_U3288) );
  AND2_X1 U16599 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15521), .ZN(P2_U3287) );
  AND2_X1 U16600 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15521), .ZN(P2_U3286) );
  AND2_X1 U16601 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15521), .ZN(P2_U3285) );
  AND2_X1 U16602 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15521), .ZN(P2_U3284) );
  AND2_X1 U16603 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15521), .ZN(P2_U3283) );
  AND2_X1 U16604 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15521), .ZN(P2_U3282) );
  AND2_X1 U16605 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15521), .ZN(P2_U3281) );
  AND2_X1 U16606 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15521), .ZN(P2_U3280) );
  AND2_X1 U16607 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15521), .ZN(P2_U3279) );
  AND2_X1 U16608 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15521), .ZN(P2_U3278) );
  AND2_X1 U16609 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15521), .ZN(P2_U3277) );
  AND2_X1 U16610 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15521), .ZN(P2_U3276) );
  AND2_X1 U16611 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15521), .ZN(P2_U3275) );
  AND2_X1 U16612 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15521), .ZN(P2_U3274) );
  AND2_X1 U16613 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15521), .ZN(P2_U3273) );
  AND2_X1 U16614 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15521), .ZN(P2_U3272) );
  AND2_X1 U16615 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15521), .ZN(P2_U3271) );
  AND2_X1 U16616 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15521), .ZN(P2_U3270) );
  AND2_X1 U16617 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15521), .ZN(P2_U3269) );
  AND2_X1 U16618 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15521), .ZN(P2_U3268) );
  AND2_X1 U16619 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15521), .ZN(P2_U3267) );
  AND2_X1 U16620 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15521), .ZN(P2_U3266) );
  NOR2_X1 U16621 ( .A1(n15522), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U16622 ( .A1(P3_U3897), .A2(n15702), .ZN(P3_U3150) );
  INV_X1 U16623 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15524) );
  AOI22_X1 U16624 ( .A1(n15526), .A2(n15525), .B1(n15524), .B2(n15523), .ZN(
        P2_U3416) );
  AOI211_X1 U16625 ( .C1(n15529), .C2(n15528), .A(n15588), .B(n15527), .ZN(
        n15534) );
  AOI211_X1 U16626 ( .C1(n15532), .C2(n15531), .A(n15592), .B(n15530), .ZN(
        n15533) );
  AOI211_X1 U16627 ( .C1(n15598), .C2(n15535), .A(n15534), .B(n15533), .ZN(
        n15537) );
  OAI211_X1 U16628 ( .C1(n15601), .C2(n15615), .A(n15537), .B(n15536), .ZN(
        P2_U3219) );
  INV_X1 U16629 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n15669) );
  AOI211_X1 U16630 ( .C1(n15540), .C2(n15539), .A(n15588), .B(n15538), .ZN(
        n15545) );
  AOI211_X1 U16631 ( .C1(n15543), .C2(n15542), .A(n15592), .B(n15541), .ZN(
        n15544) );
  AOI211_X1 U16632 ( .C1(n15598), .C2(n15546), .A(n15545), .B(n15544), .ZN(
        n15548) );
  OAI211_X1 U16633 ( .C1(n15601), .C2(n15669), .A(n15548), .B(n15547), .ZN(
        P2_U3220) );
  AOI211_X1 U16634 ( .C1(n15551), .C2(n15550), .A(n15588), .B(n15549), .ZN(
        n15556) );
  AOI211_X1 U16635 ( .C1(n15554), .C2(n15553), .A(n15592), .B(n15552), .ZN(
        n15555) );
  AOI211_X1 U16636 ( .C1(n15598), .C2(n15557), .A(n15556), .B(n15555), .ZN(
        n15559) );
  OAI211_X1 U16637 ( .C1(n15601), .C2(n15560), .A(n15559), .B(n15558), .ZN(
        P2_U3221) );
  INV_X1 U16638 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15573) );
  INV_X1 U16639 ( .A(n15561), .ZN(n15566) );
  AOI211_X1 U16640 ( .C1(n15564), .C2(n15563), .A(n15588), .B(n15562), .ZN(
        n15565) );
  AOI211_X1 U16641 ( .C1(n15598), .C2(n15567), .A(n15566), .B(n15565), .ZN(
        n15572) );
  OAI211_X1 U16642 ( .C1(n15570), .C2(n15569), .A(n15568), .B(n15583), .ZN(
        n15571) );
  OAI211_X1 U16643 ( .C1(n15601), .C2(n15573), .A(n15572), .B(n15571), .ZN(
        P2_U3231) );
  OAI21_X1 U16644 ( .B1(n15575), .B2(n15574), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15576) );
  OAI21_X1 U16645 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15576), .ZN(n15586) );
  XNOR2_X1 U16646 ( .A(n15577), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n15584) );
  OAI21_X1 U16647 ( .B1(n15580), .B2(n15579), .A(n15578), .ZN(n15582) );
  AOI22_X1 U16648 ( .A1(n15584), .A2(n15583), .B1(n15582), .B2(n15581), .ZN(
        n15585) );
  OAI211_X1 U16649 ( .C1(n15639), .C2(n15601), .A(n15586), .B(n15585), .ZN(
        P2_U3226) );
  INV_X1 U16650 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15602) );
  AOI211_X1 U16651 ( .C1(n15590), .C2(n15589), .A(n15588), .B(n15587), .ZN(
        n15596) );
  AOI211_X1 U16652 ( .C1(n15594), .C2(n15593), .A(n15592), .B(n15591), .ZN(
        n15595) );
  AOI211_X1 U16653 ( .C1(n15598), .C2(n15597), .A(n15596), .B(n15595), .ZN(
        n15600) );
  OAI211_X1 U16654 ( .C1(n15602), .C2(n15601), .A(n15600), .B(n15599), .ZN(
        P2_U3224) );
  XOR2_X1 U16655 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15603), .Z(SUB_1596_U53) );
  OAI21_X1 U16656 ( .B1(n15606), .B2(n15605), .A(n15604), .ZN(n15607) );
  XNOR2_X1 U16657 ( .A(n15607), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  OAI21_X1 U16658 ( .B1(n15610), .B2(n15609), .A(n15608), .ZN(SUB_1596_U60) );
  AOI21_X1 U16659 ( .B1(n15613), .B2(n15612), .A(n15611), .ZN(SUB_1596_U59) );
  AOI21_X1 U16660 ( .B1(n15616), .B2(n15615), .A(n15614), .ZN(SUB_1596_U58) );
  OAI21_X1 U16661 ( .B1(n15619), .B2(n15618), .A(n15617), .ZN(SUB_1596_U56) );
  OAI222_X1 U16662 ( .A1(n15624), .A2(n15623), .B1(n15624), .B2(n15622), .C1(
        n15621), .C2(n15620), .ZN(SUB_1596_U55) );
  OAI222_X1 U16663 ( .A1(n15629), .A2(n15628), .B1(n15629), .B2(n15627), .C1(
        n15626), .C2(n15625), .ZN(SUB_1596_U54) );
  AOI21_X1 U16664 ( .B1(n15632), .B2(n15631), .A(n15630), .ZN(n15633) );
  XOR2_X1 U16665 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n15633), .Z(SUB_1596_U70)
         );
  AOI21_X1 U16666 ( .B1(n15636), .B2(n15635), .A(n15634), .ZN(n15637) );
  XOR2_X1 U16667 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n15637), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16668 ( .B1(n15640), .B2(n15639), .A(n15638), .ZN(SUB_1596_U68) );
  OAI21_X1 U16669 ( .B1(n15643), .B2(n15642), .A(n15641), .ZN(n15644) );
  XNOR2_X1 U16670 ( .A(n15644), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI222_X1 U16671 ( .A1(n15649), .A2(n15648), .B1(n15649), .B2(n15647), .C1(
        n15646), .C2(n15645), .ZN(SUB_1596_U66) );
  AOI21_X1 U16672 ( .B1(n15652), .B2(n15651), .A(n15650), .ZN(n15653) );
  XOR2_X1 U16673 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15653), .Z(SUB_1596_U65)
         );
  OAI222_X1 U16674 ( .A1(n15658), .A2(n15657), .B1(n15658), .B2(n15656), .C1(
        n15655), .C2(n15654), .ZN(SUB_1596_U64) );
  AOI21_X1 U16675 ( .B1(n15661), .B2(n15660), .A(n15659), .ZN(SUB_1596_U63) );
  XOR2_X1 U16676 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n15665), .Z(SUB_1596_U62)
         );
  AOI21_X1 U16677 ( .B1(n15668), .B2(n15667), .A(n15666), .ZN(n15670) );
  XNOR2_X1 U16678 ( .A(n15670), .B(n15669), .ZN(SUB_1596_U57) );
  AOI21_X1 U16679 ( .B1(n15673), .B2(n15672), .A(n15671), .ZN(SUB_1596_U5) );
  AOI22_X1 U16680 ( .A1(n15711), .A2(n15676), .B1(n15675), .B2(n15674), .ZN(
        n15685) );
  AOI22_X1 U16681 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n15702), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n15684) );
  NAND3_X1 U16682 ( .A1(n15677), .A2(n15718), .A3(n15681), .ZN(n15678) );
  AOI22_X1 U16683 ( .A1(n15704), .A2(P3_IR_REG_0__SCAN_IN), .B1(n15679), .B2(
        n15678), .ZN(n15683) );
  OR3_X1 U16684 ( .A1(n15681), .A2(P3_IR_REG_0__SCAN_IN), .A3(n15680), .ZN(
        n15682) );
  NAND4_X1 U16685 ( .A1(n15685), .A2(n15684), .A3(n15683), .A4(n15682), .ZN(
        P3_U3182) );
  AOI22_X1 U16686 ( .A1(n15704), .A2(n15686), .B1(n15702), .B2(
        P3_ADDR_REG_10__SCAN_IN), .ZN(n15701) );
  XNOR2_X1 U16687 ( .A(n15688), .B(n15687), .ZN(n15693) );
  OAI21_X1 U16688 ( .B1(n15691), .B2(n15690), .A(n15689), .ZN(n15692) );
  AOI22_X1 U16689 ( .A1(n15693), .A2(n15712), .B1(n15711), .B2(n15692), .ZN(
        n15700) );
  AOI21_X1 U16690 ( .B1(n15696), .B2(n15695), .A(n15694), .ZN(n15697) );
  OR2_X1 U16691 ( .A1(n15697), .A2(n15718), .ZN(n15698) );
  NAND4_X1 U16692 ( .A1(n15701), .A2(n15700), .A3(n15699), .A4(n15698), .ZN(
        P3_U3192) );
  AOI22_X1 U16693 ( .A1(n15704), .A2(n15703), .B1(n15702), .B2(
        P3_ADDR_REG_12__SCAN_IN), .ZN(n15722) );
  XOR2_X1 U16694 ( .A(n15706), .B(n15705), .Z(n15713) );
  OAI21_X1 U16695 ( .B1(n15709), .B2(n15708), .A(n15707), .ZN(n15710) );
  AOI22_X1 U16696 ( .A1(n15713), .A2(n15712), .B1(n15711), .B2(n15710), .ZN(
        n15721) );
  AOI21_X1 U16697 ( .B1(n15716), .B2(n15715), .A(n15714), .ZN(n15717) );
  OR2_X1 U16698 ( .A1(n15718), .A2(n15717), .ZN(n15719) );
  NAND4_X1 U16699 ( .A1(n15722), .A2(n15721), .A3(n15720), .A4(n15719), .ZN(
        P3_U3194) );
  OAI221_X1 U16700 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n8224), .C2(n8222), .A(n15723), .ZN(U29) );
  MUX2_X1 U16701 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11692), .S(n15724), .Z(
        n15727) );
  NAND3_X1 U16702 ( .A1(n15727), .A2(n15726), .A3(n15725), .ZN(n15728) );
  NAND3_X1 U16703 ( .A1(n15730), .A2(n15729), .A3(n15728), .ZN(n15745) );
  AND2_X1 U16704 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n15731) );
  AOI21_X1 U16705 ( .B1(n15732), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n15731), .ZN(
        n15744) );
  INV_X1 U16706 ( .A(n15733), .ZN(n15738) );
  NAND3_X1 U16707 ( .A1(n15736), .A2(n15735), .A3(n15734), .ZN(n15737) );
  NAND3_X1 U16708 ( .A1(n15739), .A2(n15738), .A3(n15737), .ZN(n15743) );
  NAND2_X1 U16709 ( .A1(n15741), .A2(n15740), .ZN(n15742) );
  AND4_X1 U16710 ( .A1(n15745), .A2(n15744), .A3(n15743), .A4(n15742), .ZN(
        n15747) );
  NAND2_X1 U16711 ( .A1(n15747), .A2(n15746), .ZN(P1_U3247) );
  INV_X1 U16712 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15748) );
  AOI22_X1 U16713 ( .A1(n15994), .A2(n15749), .B1(n15748), .B2(n15992), .ZN(
        P1_U3459) );
  INV_X1 U16714 ( .A(n15750), .ZN(n15751) );
  NAND2_X1 U16715 ( .A1(n15752), .A2(n15751), .ZN(n15753) );
  OAI21_X1 U16716 ( .B1(n15755), .B2(n15754), .A(n15753), .ZN(n15757) );
  AOI211_X1 U16717 ( .C1(n15759), .C2(n15758), .A(n15757), .B(n15756), .ZN(
        n15761) );
  AOI22_X1 U16718 ( .A1(n15946), .A2(n15762), .B1(n15761), .B2(n15760), .ZN(
        P1_U3293) );
  INV_X1 U16719 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15763) );
  AOI22_X1 U16720 ( .A1(n14469), .A2(n15764), .B1(n15763), .B2(n15909), .ZN(
        P2_U3430) );
  OR2_X1 U16721 ( .A1(n15766), .A2(n15765), .ZN(n15768) );
  AOI21_X1 U16722 ( .B1(n15917), .B2(n15770), .A(n15768), .ZN(n15767) );
  AOI22_X1 U16723 ( .A1(n15997), .A2(n15767), .B1(n8269), .B2(n16004), .ZN(
        P3_U3460) );
  AOI21_X1 U16724 ( .B1(n15769), .B2(n15770), .A(n15768), .ZN(n15773) );
  AOI22_X1 U16725 ( .A1(n15771), .A2(n15770), .B1(P3_REG0_REG_1__SCAN_IN), 
        .B2(n16008), .ZN(n15772) );
  OAI21_X1 U16726 ( .B1(n15773), .B2(n16008), .A(n15772), .ZN(P3_U3393) );
  OAI21_X1 U16727 ( .B1(n15775), .B2(n15970), .A(n15774), .ZN(n15777) );
  AOI211_X1 U16728 ( .C1(n15779), .C2(n15778), .A(n15777), .B(n15776), .ZN(
        n15781) );
  AOI22_X1 U16729 ( .A1(n15991), .A2(n15781), .B1(n10320), .B2(n15990), .ZN(
        P1_U3530) );
  INV_X1 U16730 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15780) );
  AOI22_X1 U16731 ( .A1(n15994), .A2(n15781), .B1(n15780), .B2(n15992), .ZN(
        P1_U3465) );
  NOR2_X1 U16732 ( .A1(n15782), .A2(n15912), .ZN(n15784) );
  AOI211_X1 U16733 ( .C1(n15917), .C2(n15785), .A(n15784), .B(n15783), .ZN(
        n15787) );
  AOI22_X1 U16734 ( .A1(n15997), .A2(n15787), .B1(n8306), .B2(n16004), .ZN(
        P3_U3462) );
  INV_X1 U16735 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15786) );
  AOI22_X1 U16736 ( .A1(n16000), .A2(n15787), .B1(n15786), .B2(n16008), .ZN(
        P3_U3399) );
  OAI211_X1 U16737 ( .C1(n15790), .C2(n15970), .A(n15789), .B(n15788), .ZN(
        n15794) );
  AND3_X1 U16738 ( .A1(n15792), .A2(n15791), .A3(n15988), .ZN(n15793) );
  AOI211_X1 U16739 ( .C1(n15973), .C2(n15795), .A(n15794), .B(n15793), .ZN(
        n15797) );
  AOI22_X1 U16740 ( .A1(n15991), .A2(n15797), .B1(n10355), .B2(n15990), .ZN(
        P1_U3532) );
  INV_X1 U16741 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15796) );
  AOI22_X1 U16742 ( .A1(n15994), .A2(n15797), .B1(n15796), .B2(n15992), .ZN(
        P1_U3471) );
  AOI21_X1 U16743 ( .B1(n15800), .B2(n15799), .A(n15798), .ZN(n15801) );
  OAI222_X1 U16744 ( .A1(n15806), .A2(n15805), .B1(n15804), .B2(n15803), .C1(
        n15802), .C2(n15801), .ZN(n15807) );
  INV_X1 U16745 ( .A(n15807), .ZN(n15808) );
  OAI21_X1 U16746 ( .B1(n15810), .B2(n15809), .A(n15808), .ZN(P3_U3227) );
  INV_X1 U16747 ( .A(n15811), .ZN(n15812) );
  AOI222_X1 U16748 ( .A1(n15813), .A2(n15947), .B1(n15812), .B2(n15944), .C1(
        P1_REG2_REG_6__SCAN_IN), .C2(n15946), .ZN(n15818) );
  AOI22_X1 U16749 ( .A1(n15816), .A2(n15815), .B1(n15951), .B2(n15814), .ZN(
        n15817) );
  OAI211_X1 U16750 ( .C1(n15946), .C2(n15819), .A(n15818), .B(n15817), .ZN(
        P1_U3287) );
  OAI22_X1 U16751 ( .A1(n15822), .A2(n15821), .B1(n15820), .B2(n15903), .ZN(
        n15824) );
  AOI211_X1 U16752 ( .C1(n15825), .C2(n15860), .A(n15824), .B(n15823), .ZN(
        n15827) );
  AOI22_X1 U16753 ( .A1(n14451), .A2(n15827), .B1(n10869), .B2(n15908), .ZN(
        P2_U3505) );
  INV_X1 U16754 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15826) );
  AOI22_X1 U16755 ( .A1(n14469), .A2(n15827), .B1(n15826), .B2(n15909), .ZN(
        P2_U3448) );
  INV_X1 U16756 ( .A(n15831), .ZN(n15834) );
  OAI211_X1 U16757 ( .C1(n15830), .C2(n15970), .A(n15829), .B(n15828), .ZN(
        n15833) );
  NOR2_X1 U16758 ( .A1(n15831), .A2(n15875), .ZN(n15832) );
  AOI211_X1 U16759 ( .C1(n15834), .C2(n15880), .A(n15833), .B(n15832), .ZN(
        n15836) );
  AOI22_X1 U16760 ( .A1(n15991), .A2(n15836), .B1(n15835), .B2(n15990), .ZN(
        P1_U3535) );
  AOI22_X1 U16761 ( .A1(n15994), .A2(n15836), .B1(n11036), .B2(n15992), .ZN(
        P1_U3480) );
  NAND3_X1 U16762 ( .A1(n15838), .A2(n15837), .A3(n15860), .ZN(n15844) );
  AOI21_X1 U16763 ( .B1(n15841), .B2(n15840), .A(n15839), .ZN(n15842) );
  AND3_X1 U16764 ( .A1(n15844), .A2(n15843), .A3(n15842), .ZN(n15846) );
  AOI22_X1 U16765 ( .A1(n14451), .A2(n15846), .B1(n10870), .B2(n15908), .ZN(
        P2_U3506) );
  INV_X1 U16766 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15845) );
  AOI22_X1 U16767 ( .A1(n14469), .A2(n15846), .B1(n15845), .B2(n15909), .ZN(
        P2_U3451) );
  AOI21_X1 U16768 ( .B1(n15981), .B2(n15848), .A(n15847), .ZN(n15849) );
  OAI211_X1 U16769 ( .C1(n15875), .C2(n15851), .A(n15850), .B(n15849), .ZN(
        n15852) );
  INV_X1 U16770 ( .A(n15852), .ZN(n15855) );
  AOI22_X1 U16771 ( .A1(n15991), .A2(n15855), .B1(n15853), .B2(n15990), .ZN(
        P1_U3536) );
  INV_X1 U16772 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15854) );
  AOI22_X1 U16773 ( .A1(n15994), .A2(n15855), .B1(n15854), .B2(n15992), .ZN(
        P1_U3483) );
  OAI21_X1 U16774 ( .B1(n15857), .B2(n15903), .A(n15856), .ZN(n15859) );
  AOI211_X1 U16775 ( .C1(n15861), .C2(n15860), .A(n15859), .B(n15858), .ZN(
        n15863) );
  AOI22_X1 U16776 ( .A1(n14451), .A2(n15863), .B1(n10871), .B2(n15908), .ZN(
        P2_U3507) );
  INV_X1 U16777 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15862) );
  AOI22_X1 U16778 ( .A1(n14469), .A2(n15863), .B1(n15862), .B2(n15909), .ZN(
        P2_U3454) );
  NAND2_X1 U16779 ( .A1(n15864), .A2(n15917), .ZN(n15868) );
  NAND2_X1 U16780 ( .A1(n15866), .A2(n15865), .ZN(n15867) );
  AOI22_X1 U16781 ( .A1(n15997), .A2(n15871), .B1(n8372), .B2(n16004), .ZN(
        P3_U3468) );
  INV_X1 U16782 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15870) );
  AOI22_X1 U16783 ( .A1(n16000), .A2(n15871), .B1(n15870), .B2(n16008), .ZN(
        P3_U3417) );
  NAND2_X1 U16784 ( .A1(n15872), .A2(n15981), .ZN(n15873) );
  OAI211_X1 U16785 ( .C1(n15876), .C2(n15875), .A(n15874), .B(n15873), .ZN(
        n15877) );
  AOI211_X1 U16786 ( .C1(n15880), .C2(n15879), .A(n15878), .B(n15877), .ZN(
        n15883) );
  AOI22_X1 U16787 ( .A1(n15991), .A2(n15883), .B1(n15881), .B2(n15990), .ZN(
        P1_U3537) );
  INV_X1 U16788 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15882) );
  AOI22_X1 U16789 ( .A1(n15994), .A2(n15883), .B1(n15882), .B2(n15992), .ZN(
        P1_U3486) );
  INV_X1 U16790 ( .A(n15884), .ZN(n15888) );
  NOR2_X1 U16791 ( .A1(n15885), .A2(n15912), .ZN(n15887) );
  AOI211_X1 U16792 ( .C1(n15889), .C2(n15888), .A(n15887), .B(n15886), .ZN(
        n15890) );
  AOI22_X1 U16793 ( .A1(n15997), .A2(n15890), .B1(n7733), .B2(n16004), .ZN(
        P3_U3469) );
  AOI22_X1 U16794 ( .A1(n16000), .A2(n15890), .B1(n8395), .B2(n16008), .ZN(
        P3_U3420) );
  OAI211_X1 U16795 ( .C1(n15893), .C2(n15970), .A(n15892), .B(n15891), .ZN(
        n15897) );
  AND3_X1 U16796 ( .A1(n15895), .A2(n15988), .A3(n15894), .ZN(n15896) );
  AOI211_X1 U16797 ( .C1(n15973), .C2(n15898), .A(n15897), .B(n15896), .ZN(
        n15900) );
  AOI22_X1 U16798 ( .A1(n15991), .A2(n15900), .B1(n15899), .B2(n15990), .ZN(
        P1_U3538) );
  AOI22_X1 U16799 ( .A1(n15994), .A2(n15900), .B1(n11591), .B2(n15992), .ZN(
        P1_U3489) );
  INV_X1 U16800 ( .A(n15901), .ZN(n15907) );
  OAI21_X1 U16801 ( .B1(n15904), .B2(n15903), .A(n15902), .ZN(n15906) );
  AOI211_X1 U16802 ( .C1(n9444), .C2(n15907), .A(n15906), .B(n15905), .ZN(
        n15911) );
  AOI22_X1 U16803 ( .A1(n14451), .A2(n15911), .B1(n11530), .B2(n15908), .ZN(
        P2_U3509) );
  INV_X1 U16804 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15910) );
  AOI22_X1 U16805 ( .A1(n14469), .A2(n15911), .B1(n15910), .B2(n15909), .ZN(
        P2_U3460) );
  NOR2_X1 U16806 ( .A1(n15913), .A2(n15912), .ZN(n15915) );
  AOI211_X1 U16807 ( .C1(n15917), .C2(n15916), .A(n15915), .B(n15914), .ZN(
        n15919) );
  AOI22_X1 U16808 ( .A1(n15997), .A2(n15919), .B1(n11538), .B2(n16004), .ZN(
        P3_U3470) );
  INV_X1 U16809 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15918) );
  AOI22_X1 U16810 ( .A1(n16000), .A2(n15919), .B1(n15918), .B2(n16008), .ZN(
        P3_U3423) );
  AOI211_X1 U16811 ( .C1(n15981), .C2(n15922), .A(n15921), .B(n15920), .ZN(
        n15925) );
  NAND3_X1 U16812 ( .A1(n11963), .A2(n15923), .A3(n15973), .ZN(n15924) );
  AOI22_X1 U16813 ( .A1(n15991), .A2(n15927), .B1(n11602), .B2(n15990), .ZN(
        P1_U3539) );
  INV_X1 U16814 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n15926) );
  AOI22_X1 U16815 ( .A1(n15994), .A2(n15927), .B1(n15926), .B2(n15992), .ZN(
        P1_U3492) );
  OAI21_X1 U16816 ( .B1(n15930), .B2(n11969), .A(n15929), .ZN(n15953) );
  OAI211_X1 U16817 ( .C1(n15933), .C2(n15934), .A(n15932), .B(n15931), .ZN(
        n15949) );
  OAI21_X1 U16818 ( .B1(n15934), .B2(n15970), .A(n15949), .ZN(n15941) );
  INV_X1 U16819 ( .A(n15935), .ZN(n15936) );
  AOI21_X1 U16820 ( .B1(n15936), .B2(n11969), .A(n15959), .ZN(n15939) );
  AOI21_X1 U16821 ( .B1(n15939), .B2(n15938), .A(n15937), .ZN(n15956) );
  INV_X1 U16822 ( .A(n15956), .ZN(n15940) );
  AOI211_X1 U16823 ( .C1(n15973), .C2(n15953), .A(n15941), .B(n15940), .ZN(
        n15942) );
  AOI22_X1 U16824 ( .A1(n15991), .A2(n15942), .B1(n10693), .B2(n15990), .ZN(
        P1_U3540) );
  AOI22_X1 U16825 ( .A1(n15994), .A2(n15942), .B1(n11748), .B2(n15992), .ZN(
        P1_U3495) );
  INV_X1 U16826 ( .A(n15943), .ZN(n15945) );
  AOI222_X1 U16827 ( .A1(n15948), .A2(n15947), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n15946), .C1(n15945), .C2(n15944), .ZN(n15955) );
  INV_X1 U16828 ( .A(n15949), .ZN(n15950) );
  AOI22_X1 U16829 ( .A1(n15953), .A2(n15952), .B1(n15951), .B2(n15950), .ZN(
        n15954) );
  OAI211_X1 U16830 ( .C1(n15946), .C2(n15956), .A(n15955), .B(n15954), .ZN(
        P1_U3281) );
  OAI211_X1 U16831 ( .C1(n7606), .C2(n15970), .A(n15958), .B(n15957), .ZN(
        n15963) );
  NOR3_X1 U16832 ( .A1(n15961), .A2(n15960), .A3(n15959), .ZN(n15962) );
  AOI211_X1 U16833 ( .C1(n15964), .C2(n15973), .A(n15963), .B(n15962), .ZN(
        n15966) );
  AOI22_X1 U16834 ( .A1(n15991), .A2(n15966), .B1(n15965), .B2(n15990), .ZN(
        P1_U3541) );
  AOI22_X1 U16835 ( .A1(n15994), .A2(n15966), .B1(n11975), .B2(n15992), .ZN(
        P1_U3498) );
  INV_X1 U16836 ( .A(n15967), .ZN(n15971) );
  OAI211_X1 U16837 ( .C1(n15971), .C2(n15970), .A(n15969), .B(n15968), .ZN(
        n15976) );
  AND3_X1 U16838 ( .A1(n15974), .A2(n15973), .A3(n15972), .ZN(n15975) );
  AOI211_X1 U16839 ( .C1(n15977), .C2(n15988), .A(n15976), .B(n15975), .ZN(
        n15979) );
  AOI22_X1 U16840 ( .A1(n15991), .A2(n15979), .B1(n15978), .B2(n15990), .ZN(
        P1_U3542) );
  AOI22_X1 U16841 ( .A1(n15994), .A2(n15979), .B1(n11988), .B2(n15992), .ZN(
        P1_U3501) );
  AOI21_X1 U16842 ( .B1(n15982), .B2(n15981), .A(n15980), .ZN(n15984) );
  OAI211_X1 U16843 ( .C1(n15986), .C2(n15985), .A(n15984), .B(n15983), .ZN(
        n15987) );
  AOI21_X1 U16844 ( .B1(n15989), .B2(n15988), .A(n15987), .ZN(n15993) );
  AOI22_X1 U16845 ( .A1(n15991), .A2(n15993), .B1(n12014), .B2(n15990), .ZN(
        P1_U3543) );
  AOI22_X1 U16846 ( .A1(n15994), .A2(n15993), .B1(n12013), .B2(n15992), .ZN(
        P1_U3504) );
  INV_X1 U16847 ( .A(n15995), .ZN(n15999) );
  AOI22_X1 U16848 ( .A1(n15999), .A2(n16005), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n16004), .ZN(n15998) );
  INV_X1 U16849 ( .A(n15996), .ZN(n16001) );
  NAND2_X1 U16850 ( .A1(n16001), .A2(n15997), .ZN(n16006) );
  NAND2_X1 U16851 ( .A1(n15998), .A2(n16006), .ZN(P3_U3489) );
  AOI22_X1 U16852 ( .A1(n15999), .A2(n16009), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n16008), .ZN(n16002) );
  NAND2_X1 U16853 ( .A1(n16001), .A2(n16000), .ZN(n16011) );
  NAND2_X1 U16854 ( .A1(n16002), .A2(n16011), .ZN(P3_U3457) );
  INV_X1 U16855 ( .A(n16003), .ZN(n16010) );
  AOI22_X1 U16856 ( .A1(n16010), .A2(n16005), .B1(P3_REG1_REG_31__SCAN_IN), 
        .B2(n16004), .ZN(n16007) );
  NAND2_X1 U16857 ( .A1(n16007), .A2(n16006), .ZN(P3_U3490) );
  AOI22_X1 U16858 ( .A1(n16010), .A2(n16009), .B1(P3_REG0_REG_31__SCAN_IN), 
        .B2(n16008), .ZN(n16012) );
  NAND2_X1 U16859 ( .A1(n16012), .A2(n16011), .ZN(P3_U3458) );
  AOI21_X1 U16860 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16013) );
  OAI21_X1 U16861 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16013), 
        .ZN(U28) );
  INV_X1 U9516 ( .A(n8270), .ZN(n13029) );
  CLKBUF_X1 U7299 ( .A(n9475), .Z(n9604) );
  CLKBUF_X1 U7379 ( .A(n14914), .Z(n14920) );
  MUX2_X1 U8808 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15485), .S(n7201), .Z(n10484)
         );
  INV_X1 U11363 ( .A(n8172), .ZN(n13158) );
  CLKBUF_X1 U12204 ( .A(n14935), .Z(n7187) );
endmodule

