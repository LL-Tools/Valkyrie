

module b15_C_SARLock_k_64_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2970, n2974, n2975, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796;

  CLKBUF_X1 U3419 ( .A(n3576), .Z(n2985) );
  OAI21_X1 U3420 ( .B1(n4703), .B2(n3363), .A(n3362), .ZN(n6269) );
  INV_X1 U3421 ( .A(n4304), .ZN(n4315) );
  INV_X1 U3422 ( .A(n4323), .ZN(n3523) );
  CLKBUF_X1 U3424 ( .A(n2978), .Z(n2979) );
  BUF_X1 U3426 ( .A(n3194), .Z(n2989) );
  AND2_X2 U3427 ( .A1(n3116), .A2(n4500), .ZN(n2997) );
  AND2_X1 U3428 ( .A1(n3116), .A2(n4490), .ZN(n3266) );
  AND2_X1 U3429 ( .A1(n4506), .A2(n3114), .ZN(n3193) );
  AND2_X4 U3430 ( .A1(n4490), .A2(n3035), .ZN(n2984) );
  CLKBUF_X2 U3431 ( .A(n3158), .Z(n2975) );
  INV_X2 U3432 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3109) );
  AND2_X1 U3434 ( .A1(n3353), .A2(n3325), .ZN(n3331) );
  NAND2_X1 U3435 ( .A1(n3331), .A2(n3330), .ZN(n3342) );
  AND4_X1 U3436 ( .A1(n3126), .A2(n3125), .A3(n3124), .A4(n3123), .ZN(n3132)
         );
  OR2_X1 U3439 ( .A1(n3459), .A2(n3458), .ZN(n3461) );
  NAND2_X1 U3440 ( .A1(n3155), .A2(n4304), .ZN(n3241) );
  AND2_X2 U3441 ( .A1(n3132), .A2(n3131), .ZN(n4304) );
  INV_X1 U3442 ( .A(n4874), .ZN(n3339) );
  INV_X1 U3444 ( .A(n3155), .ZN(n3214) );
  AND2_X1 U34450 ( .A1(n3508), .A2(n5582), .ZN(n3022) );
  INV_X1 U34460 ( .A(n3493), .ZN(n5917) );
  OR2_X1 U34470 ( .A1(n3345), .A2(n3344), .ZN(n3347) );
  NAND3_X1 U34480 ( .A1(n3029), .A2(n3038), .A3(n3028), .ZN(n4330) );
  NAND2_X2 U3449 ( .A1(n3347), .A2(n3346), .ZN(n4259) );
  OR2_X2 U3450 ( .A1(n3143), .A2(n3142), .ZN(n4645) );
  AND2_X1 U34510 ( .A1(n5604), .A2(n3097), .ZN(n5588) );
  OR2_X2 U34520 ( .A1(n3200), .A2(n3199), .ZN(n4874) );
  XNOR2_X1 U34530 ( .A(n3468), .B(n6311), .ZN(n4914) );
  OR2_X1 U3454 ( .A1(n3357), .A2(n3356), .ZN(n4703) );
  INV_X1 U34560 ( .A(n6072), .ZN(n6103) );
  INV_X2 U3457 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3108) );
  AND2_X1 U3458 ( .A1(n3295), .A2(n3235), .ZN(n3279) );
  XNOR2_X1 U34590 ( .A(n3295), .B(n3294), .ZN(n3576) );
  AND2_X1 U34600 ( .A1(n4500), .A2(n3035), .ZN(n2970) );
  AND2_X2 U34610 ( .A1(n4833), .A2(n3012), .ZN(n5184) );
  AND2_X1 U34620 ( .A1(n4803), .A2(n4801), .ZN(n4833) );
  NAND2_X1 U34630 ( .A1(n4649), .A2(n3088), .ZN(n4781) );
  INV_X2 U34640 ( .A(n3079), .ZN(n4655) );
  CLKBUF_X2 U34650 ( .A(n6166), .Z(n6228) );
  AND2_X1 U3466 ( .A1(n5131), .A2(n4116), .ZN(n5189) );
  AND3_X1 U3467 ( .A1(n3234), .A2(n4192), .A3(n3233), .ZN(n3294) );
  CLKBUF_X2 U34680 ( .A(n3259), .Z(n5282) );
  CLKBUF_X2 U34690 ( .A(n5283), .Z(n4014) );
  CLKBUF_X2 U34700 ( .A(n3157), .Z(n3873) );
  AND2_X1 U34710 ( .A1(n3109), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4507) );
  AND2_X1 U34720 ( .A1(n4512), .A2(n3115), .ZN(n3194) );
  AND2_X2 U34730 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3035) );
  NAND2_X1 U34740 ( .A1(n3070), .A2(n3069), .ZN(n5615) );
  OAI21_X1 U3475 ( .B1(n5522), .B2(n5872), .A(n3052), .ZN(n3051) );
  INV_X1 U3476 ( .A(n5552), .ZN(n5522) );
  OAI21_X1 U3477 ( .B1(n4029), .B2(n4030), .A(n5353), .ZN(n5380) );
  NAND2_X1 U3478 ( .A1(n3091), .A2(n3094), .ZN(n5353) );
  AND2_X1 U3479 ( .A1(n5391), .A2(n5570), .ZN(n5891) );
  XOR2_X1 U3480 ( .A(n5355), .B(n5354), .Z(n5374) );
  NOR2_X1 U3481 ( .A1(n5391), .A2(n5392), .ZN(n4029) );
  AND2_X1 U3482 ( .A1(n5569), .A2(n3090), .ZN(n5354) );
  AOI21_X1 U3483 ( .B1(n5537), .B2(n5536), .A(n5535), .ZN(n6105) );
  AND2_X1 U3484 ( .A1(n5509), .A2(n5508), .ZN(n6124) );
  AND2_X1 U3485 ( .A1(n5534), .A2(n5456), .ZN(n5461) );
  OR2_X1 U3486 ( .A1(n5428), .A2(n5414), .ZN(n5633) );
  OR2_X1 U3487 ( .A1(n5536), .A2(n5537), .ZN(n5534) );
  AND2_X1 U3488 ( .A1(n5460), .A2(n5459), .ZN(n5507) );
  NAND2_X1 U3489 ( .A1(n3057), .A2(n3055), .ZN(n5256) );
  XNOR2_X1 U3490 ( .A(n4182), .B(n4181), .ZN(n5477) );
  NAND2_X1 U3491 ( .A1(n5320), .A2(n5319), .ZN(n5671) );
  AOI21_X1 U3492 ( .B1(n3060), .B2(n3496), .A(n3006), .ZN(n3059) );
  NAND2_X1 U3493 ( .A1(n5700), .A2(n5393), .ZN(n5395) );
  NOR2_X1 U3494 ( .A1(n3063), .A2(n5231), .ZN(n3060) );
  NAND2_X1 U3495 ( .A1(n3496), .A2(n3062), .ZN(n3061) );
  AND2_X1 U3496 ( .A1(n5207), .A2(n3495), .ZN(n3496) );
  NAND2_X1 U3497 ( .A1(n3589), .A2(n3588), .ZN(n4649) );
  NAND2_X1 U3498 ( .A1(n3617), .A2(n3616), .ZN(n4780) );
  NOR2_X1 U3499 ( .A1(n3092), .A2(n3987), .ZN(n3090) );
  AND2_X1 U3500 ( .A1(n4650), .A2(n3089), .ZN(n3088) );
  OR2_X1 U3501 ( .A1(n3587), .A2(n4378), .ZN(n4436) );
  NAND2_X1 U3502 ( .A1(n3096), .A2(n3926), .ZN(n3587) );
  AND2_X1 U3503 ( .A1(n4376), .A2(n4375), .ZN(n4378) );
  NAND2_X1 U3504 ( .A1(n3398), .A2(n3397), .ZN(n3399) );
  INV_X1 U3505 ( .A(n3423), .ZN(n3033) );
  AOI21_X1 U3506 ( .B1(n4277), .B2(n4276), .A(n3368), .ZN(n6255) );
  NAND2_X1 U3507 ( .A1(n5786), .A2(n4135), .ZN(n5511) );
  NAND2_X1 U3508 ( .A1(n3392), .A2(n3391), .ZN(n4284) );
  CLKBUF_X1 U3509 ( .A(n4286), .Z(n2990) );
  NOR2_X1 U3511 ( .A1(n4651), .A2(n4742), .ZN(n6446) );
  NAND2_X1 U3512 ( .A1(n3037), .A2(n3036), .ZN(n6052) );
  INV_X1 U3513 ( .A(n4608), .ZN(n3037) );
  NAND2_X1 U3514 ( .A1(n3257), .A2(n3256), .ZN(n3258) );
  NAND2_X1 U3515 ( .A1(n3221), .A2(n3220), .ZN(n3295) );
  NAND2_X1 U3516 ( .A1(n4562), .A2(n4561), .ZN(n4608) );
  AND2_X1 U3517 ( .A1(n4698), .A2(n4311), .ZN(n4562) );
  NOR2_X1 U3518 ( .A1(n4433), .A2(n3048), .ZN(n4698) );
  NAND2_X1 U3519 ( .A1(n3242), .A2(n3101), .ZN(n5976) );
  INV_X1 U3520 ( .A(n4607), .ZN(n3036) );
  AND2_X1 U3521 ( .A1(n3205), .A2(n4195), .ZN(n3231) );
  NOR2_X1 U3522 ( .A1(n3543), .A2(n4050), .ZN(n3216) );
  NAND2_X1 U3523 ( .A1(n4083), .A2(n5444), .ZN(n4344) );
  CLKBUF_X1 U3524 ( .A(n3224), .Z(n6152) );
  AND2_X1 U3525 ( .A1(n5444), .A2(n4307), .ZN(n4158) );
  INV_X1 U3526 ( .A(n3223), .ZN(n3575) );
  INV_X1 U3527 ( .A(n4642), .ZN(n4050) );
  INV_X1 U3528 ( .A(n4077), .ZN(n3204) );
  NAND2_X1 U3529 ( .A1(n4323), .A2(n4330), .ZN(n4077) );
  AND2_X2 U3530 ( .A1(n4874), .A2(n4323), .ZN(n4307) );
  OR2_X1 U3531 ( .A1(n3306), .A2(n3305), .ZN(n3484) );
  AND4_X1 U3532 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3167)
         );
  AND4_X1 U3533 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .ZN(n3131)
         );
  AND2_X1 U3534 ( .A1(n3175), .A2(n3172), .ZN(n3028) );
  AOI21_X1 U3535 ( .B1(n3193), .B2(INSTQUEUE_REG_10__7__SCAN_IN), .A(n3137), 
        .ZN(n3141) );
  INV_X2 U3536 ( .A(n2993), .ZN(n2994) );
  AND2_X1 U3537 ( .A1(n3171), .A2(n3170), .ZN(n3038) );
  INV_X2 U3538 ( .A(n6271), .ZN(n6258) );
  BUF_X2 U3540 ( .A(n3307), .Z(n5285) );
  BUF_X2 U3542 ( .A(n3266), .Z(n3992) );
  INV_X2 U3543 ( .A(n6622), .ZN(n6608) );
  BUF_X4 U3544 ( .A(n2978), .Z(n2974) );
  AND2_X2 U3545 ( .A1(n5340), .A2(n3035), .ZN(n3259) );
  AND2_X2 U3546 ( .A1(n3108), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5340)
         );
  AND2_X1 U3547 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4512) );
  NOR2_X1 U3548 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4864) );
  NAND2_X4 U3549 ( .A1(n3122), .A2(n3121), .ZN(n3155) );
  AOI21_X1 U3550 ( .B1(n3609), .B2(n3732), .A(n3608), .ZN(n4300) );
  XNOR2_X1 U3551 ( .A(n3459), .B(n3457), .ZN(n3610) );
  INV_X1 U3552 ( .A(n3193), .ZN(n2993) );
  NAND2_X2 U3553 ( .A1(n3022), .A2(n3509), .ZN(n3021) );
  NAND2_X2 U3554 ( .A1(n3214), .A2(n4319), .ZN(n3209) );
  NAND2_X2 U3555 ( .A1(n5605), .A2(n3505), .ZN(n5592) );
  XNOR2_X1 U3556 ( .A(n3423), .B(n3424), .ZN(n3609) );
  NOR2_X2 U3557 ( .A1(n3236), .A2(n4049), .ZN(n4494) );
  AND2_X1 U3558 ( .A1(n3114), .A2(n3116), .ZN(n2978) );
  AND2_X1 U3559 ( .A1(n3114), .A2(n3116), .ZN(n3158) );
  AND2_X1 U3560 ( .A1(n4506), .A2(n4490), .ZN(n2992) );
  AND2_X2 U3561 ( .A1(n4506), .A2(n4490), .ZN(n3265) );
  AND2_X2 U3562 ( .A1(n4914), .A2(n3446), .ZN(n3076) );
  NAND2_X2 U3563 ( .A1(n3467), .A2(n3466), .ZN(n3468) );
  NAND2_X2 U3564 ( .A1(n3018), .A2(n5108), .ZN(n5116) );
  XNOR2_X2 U3565 ( .A(n3279), .B(n3281), .ZN(n4262) );
  AND2_X1 U3566 ( .A1(n4507), .A2(n4500), .ZN(n2982) );
  AND2_X1 U3567 ( .A1(n4507), .A2(n4500), .ZN(n2986) );
  AND2_X4 U3568 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4500) );
  AND2_X1 U3569 ( .A1(n4490), .A2(n3035), .ZN(n2983) );
  AND2_X1 U3570 ( .A1(n4490), .A2(n3035), .ZN(n5284) );
  AOI21_X2 U3571 ( .B1(n3576), .B2(n6669), .A(n3323), .ZN(n3353) );
  AND2_X2 U3572 ( .A1(n4507), .A2(n4500), .ZN(n3403) );
  BUF_X4 U3573 ( .A(n3194), .Z(n2987) );
  AND2_X2 U3574 ( .A1(n4506), .A2(n4490), .ZN(n2991) );
  AND2_X4 U3575 ( .A1(n4506), .A2(n4500), .ZN(n2995) );
  AND2_X1 U3576 ( .A1(n3116), .A2(n4500), .ZN(n2996) );
  AND2_X1 U3578 ( .A1(n3116), .A2(n4500), .ZN(n3260) );
  AND2_X4 U3579 ( .A1(n5340), .A2(n3116), .ZN(n3000) );
  AND2_X4 U3580 ( .A1(n5340), .A2(n3116), .ZN(n3380) );
  NOR2_X4 U3581 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4490) );
  AND2_X1 U3582 ( .A1(n6084), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5359) );
  AND2_X1 U3583 ( .A1(n4480), .A2(n6490), .ZN(n6149) );
  NAND2_X1 U3584 ( .A1(n3402), .A2(n4284), .ZN(n3423) );
  NOR2_X1 U3585 ( .A1(n3258), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3065) );
  NAND2_X1 U3586 ( .A1(n4494), .A2(n3023), .ZN(n3026) );
  INV_X1 U3587 ( .A(n3379), .ZN(n3276) );
  NAND2_X1 U3588 ( .A1(n3379), .A2(n3378), .ZN(n3559) );
  INV_X1 U3589 ( .A(n4319), .ZN(n3570) );
  INV_X1 U3590 ( .A(n5404), .ZN(n3931) );
  OAI21_X1 U3591 ( .B1(n5228), .B2(n3016), .A(n3081), .ZN(n5263) );
  INV_X1 U3592 ( .A(n5218), .ZN(n3086) );
  AND2_X1 U3593 ( .A1(n3155), .A2(n4323), .ZN(n3519) );
  NAND2_X1 U3594 ( .A1(n4304), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3378) );
  NAND2_X1 U3595 ( .A1(n3570), .A2(n4645), .ZN(n3223) );
  OR3_X1 U3596 ( .A1(n6614), .A2(n6495), .A3(n4866), .ZN(n6084) );
  NAND2_X1 U3597 ( .A1(n3155), .A2(n3570), .ZN(n4642) );
  NAND2_X1 U3598 ( .A1(n4913), .A2(n3479), .ZN(n4900) );
  NAND2_X1 U3599 ( .A1(n4071), .A2(n4070), .ZN(n4204) );
  INV_X1 U3600 ( .A(n3274), .ZN(n3543) );
  AOI21_X1 U3601 ( .B1(n4923), .B2(n3241), .A(n3222), .ZN(n4191) );
  INV_X1 U3602 ( .A(n4864), .ZN(n5279) );
  INV_X1 U3603 ( .A(n5279), .ZN(n4028) );
  NAND2_X1 U3604 ( .A1(n5408), .A2(n5716), .ZN(n3045) );
  NAND2_X1 U3605 ( .A1(n3493), .A2(n6659), .ZN(n3075) );
  INV_X1 U3606 ( .A(n5621), .ZN(n3073) );
  NOR2_X1 U3607 ( .A1(n3078), .A2(n3010), .ZN(n3027) );
  OR2_X1 U3608 ( .A1(n3318), .A2(n3317), .ZN(n3360) );
  XNOR2_X1 U3609 ( .A(n3278), .B(n3277), .ZN(n3337) );
  OAI211_X1 U3610 ( .C1(n3068), .C2(n3067), .A(n3066), .B(n3007), .ZN(n3278)
         );
  NAND2_X1 U3611 ( .A1(n3377), .A2(n3376), .ZN(n4263) );
  AND2_X1 U3612 ( .A1(n6592), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3566) );
  OR2_X1 U3613 ( .A1(n4187), .A2(n3155), .ZN(n3236) );
  AND2_X1 U3614 ( .A1(n4143), .A2(n4142), .ZN(n5445) );
  INV_X1 U3615 ( .A(n3594), .ZN(n5351) );
  NAND2_X1 U3616 ( .A1(n3094), .A2(n3093), .ZN(n3092) );
  INV_X1 U3617 ( .A(n5352), .ZN(n3093) );
  INV_X1 U3618 ( .A(n5391), .ZN(n3091) );
  AND2_X1 U3619 ( .A1(n5278), .A2(n4009), .ZN(n5382) );
  NOR2_X1 U3620 ( .A1(n5585), .A2(n3099), .ZN(n3097) );
  NAND2_X1 U3621 ( .A1(n5604), .A2(n3098), .ZN(n5586) );
  INV_X1 U3622 ( .A(n5231), .ZN(n3062) );
  NAND2_X1 U3623 ( .A1(n3712), .A2(n3711), .ZN(n5228) );
  NOR2_X1 U3624 ( .A1(n6233), .A2(n3482), .ZN(n3489) );
  NOR2_X1 U3625 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  NAND2_X1 U3626 ( .A1(n3629), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3647)
         );
  INV_X1 U3627 ( .A(n4300), .ZN(n3089) );
  NAND2_X1 U3628 ( .A1(n3021), .A2(n3009), .ZN(n5566) );
  NAND2_X1 U3629 ( .A1(n5418), .A2(n5417), .ZN(n5497) );
  NAND2_X1 U3630 ( .A1(n5917), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U3631 ( .A1(n5910), .A2(n5593), .ZN(n5628) );
  OR2_X1 U3632 ( .A1(n3493), .A2(n5932), .ZN(n5593) );
  OR2_X1 U3633 ( .A1(n6597), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4034) );
  NOR2_X1 U3634 ( .A1(n3497), .A2(n3064), .ZN(n3063) );
  INV_X1 U3635 ( .A(n5115), .ZN(n3064) );
  NAND2_X1 U3636 ( .A1(n5106), .A2(n5107), .ZN(n3018) );
  AND2_X1 U3637 ( .A1(n6362), .A2(n5950), .ZN(n5118) );
  AND2_X1 U3638 ( .A1(n4092), .A2(n4091), .ZN(n4696) );
  OR2_X1 U3639 ( .A1(n5118), .A2(n4278), .ZN(n4554) );
  OR2_X1 U3640 ( .A1(n3241), .A2(n4874), .ZN(n4047) );
  NAND3_X1 U3641 ( .A1(n3215), .A2(n3225), .A3(n4645), .ZN(n4048) );
  NAND2_X1 U3642 ( .A1(n3211), .A2(n3176), .ZN(n3212) );
  NOR2_X1 U3643 ( .A1(n3041), .A2(n3040), .ZN(n3039) );
  NAND2_X1 U3644 ( .A1(n3565), .A2(n3564), .ZN(n4480) );
  NAND2_X1 U3645 ( .A1(n3561), .A2(n3560), .ZN(n3565) );
  AND2_X1 U3646 ( .A1(n3566), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6490) );
  AND2_X1 U3647 ( .A1(n5364), .A2(REIP_REG_30__SCAN_IN), .ZN(n3054) );
  INV_X1 U3648 ( .A(n5323), .ZN(n3053) );
  AND2_X1 U3649 ( .A1(n5359), .A2(n4881), .ZN(n6090) );
  INV_X1 U3650 ( .A(n6090), .ZN(n6079) );
  AND2_X1 U3651 ( .A1(n5544), .A2(n4644), .ZN(n6122) );
  AND2_X1 U3652 ( .A1(n5544), .A2(n4646), .ZN(n6126) );
  NOR2_X1 U3653 ( .A1(n5278), .A2(n5321), .ZN(n4863) );
  INV_X1 U3654 ( .A(n6264), .ZN(n5649) );
  AND2_X1 U3655 ( .A1(n6149), .A2(n4229), .ZN(n6257) );
  AND2_X1 U3656 ( .A1(n3240), .A2(n4874), .ZN(n3023) );
  NOR2_X1 U3657 ( .A1(n3237), .A2(n3528), .ZN(n3547) );
  AND2_X1 U3658 ( .A1(n3733), .A2(n5250), .ZN(n3082) );
  OR2_X1 U3659 ( .A1(n3733), .A2(n3084), .ZN(n3083) );
  INV_X1 U3660 ( .A(n5250), .ZN(n3084) );
  NAND2_X1 U3661 ( .A1(n3033), .A2(n3424), .ZN(n3459) );
  OR2_X1 U3662 ( .A1(n3456), .A2(n3455), .ZN(n3474) );
  OR2_X1 U3663 ( .A1(n3413), .A2(n3412), .ZN(n3437) );
  OR2_X1 U3664 ( .A1(n3291), .A2(n3290), .ZN(n3348) );
  NAND2_X1 U3665 ( .A1(n3258), .A2(n6669), .ZN(n3067) );
  OR2_X1 U3666 ( .A1(n3273), .A2(n3272), .ZN(n3275) );
  AND2_X1 U3667 ( .A1(n4030), .A2(n3095), .ZN(n3094) );
  INV_X1 U3668 ( .A(n5392), .ZN(n3095) );
  NOR2_X1 U3669 ( .A1(n3818), .A2(n3734), .ZN(n3803) );
  AND2_X1 U3670 ( .A1(n3662), .A2(n4832), .ZN(n3087) );
  INV_X1 U3671 ( .A(n4931), .ZN(n3662) );
  NAND2_X1 U3672 ( .A1(n4655), .A2(n3732), .ZN(n3096) );
  INV_X1 U3673 ( .A(n3275), .ZN(n3393) );
  NAND2_X1 U3674 ( .A1(n6254), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3369)
         );
  INV_X1 U3675 ( .A(n3348), .ZN(n3326) );
  INV_X1 U3676 ( .A(n3342), .ZN(n3332) );
  OR2_X1 U3677 ( .A1(n3247), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3248)
         );
  INV_X1 U3678 ( .A(n3566), .ZN(n3255) );
  AOI21_X1 U3679 ( .B1(n4048), .B2(n3276), .A(n3216), .ZN(n3217) );
  AND4_X1 U3680 ( .A1(n4191), .A2(n3227), .A3(n4515), .A4(n3226), .ZN(n3234)
         );
  NOR2_X1 U3681 ( .A1(n3210), .A2(n4330), .ZN(n4305) );
  AOI22_X1 U3682 ( .A1(n2982), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3195) );
  NAND2_X1 U3683 ( .A1(n2989), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U3684 ( .A1(n3193), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U3685 ( .A1(n3185), .A2(n3187), .ZN(n3041) );
  NAND3_X1 U3686 ( .A1(n3168), .A2(n3174), .A3(n3173), .ZN(n3030) );
  AOI22_X1 U3687 ( .A1(n2982), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U3688 ( .A1(n4286), .A2(n6669), .ZN(n3392) );
  AND2_X1 U3689 ( .A1(n3558), .A2(n3557), .ZN(n4060) );
  OR2_X1 U3690 ( .A1(n3556), .A2(n3555), .ZN(n3558) );
  AOI21_X1 U3691 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6669), .A(n3554), 
        .ZN(n3561) );
  OAI21_X1 U3692 ( .B1(n4061), .B2(n3563), .A(n3553), .ZN(n3554) );
  INV_X1 U3693 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6478) );
  INV_X1 U3694 ( .A(n5448), .ZN(n6095) );
  NOR2_X1 U3695 ( .A1(n5252), .A2(n5251), .ZN(n5266) );
  AND2_X1 U3696 ( .A1(n6149), .A2(n4248), .ZN(n6129) );
  NAND2_X1 U3697 ( .A1(n6149), .A2(n4227), .ZN(n6150) );
  OR2_X1 U3698 ( .A1(n5550), .A2(n5279), .ZN(n5304) );
  OR2_X1 U3699 ( .A1(n4008), .A2(n4035), .ZN(n5278) );
  NAND2_X1 U3700 ( .A1(n3988), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4008)
         );
  NOR2_X1 U3701 ( .A1(n3933), .A2(n5827), .ZN(n3969) );
  AND2_X1 U3702 ( .A1(n3913), .A2(n3912), .ZN(n5603) );
  OR2_X1 U3703 ( .A1(n5841), .A2(n5279), .ZN(n3913) );
  NAND2_X1 U3704 ( .A1(n5604), .A2(n5603), .ZN(n5602) );
  OR2_X1 U3705 ( .A1(n3886), .A2(n3908), .ZN(n3932) );
  NAND2_X1 U3706 ( .A1(n3751), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3853)
         );
  AND2_X1 U3707 ( .A1(n3851), .A2(n5426), .ZN(n3852) );
  NOR2_X1 U3708 ( .A1(n3799), .A2(n5451), .ZN(n3752) );
  AND2_X1 U3709 ( .A1(n3752), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3751)
         );
  AND2_X1 U3710 ( .A1(n3803), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3800)
         );
  NAND2_X1 U3711 ( .A1(n3800), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3799)
         );
  NOR2_X1 U3712 ( .A1(n3717), .A2(n3714), .ZN(n3843) );
  AOI21_X1 U3713 ( .B1(n3059), .B2(n3061), .A(n3056), .ZN(n3055) );
  NAND2_X1 U3714 ( .A1(n5116), .A2(n3059), .ZN(n3057) );
  INV_X1 U3715 ( .A(n5257), .ZN(n3056) );
  NOR2_X1 U3716 ( .A1(n3694), .A2(n5195), .ZN(n3713) );
  NAND2_X1 U3717 ( .A1(n3690), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3694)
         );
  NOR2_X1 U3718 ( .A1(n3664), .A2(n3663), .ZN(n3690) );
  OR2_X1 U3719 ( .A1(n3647), .A2(n4896), .ZN(n3664) );
  NAND2_X1 U3720 ( .A1(n4833), .A2(n3087), .ZN(n5219) );
  NAND2_X1 U3721 ( .A1(n4833), .A2(n4832), .ZN(n4932) );
  NAND2_X1 U3722 ( .A1(n3633), .A2(n3632), .ZN(n4801) );
  NAND2_X1 U3723 ( .A1(n4780), .A2(n4605), .ZN(n3625) );
  NAND2_X1 U3724 ( .A1(n3611), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3628)
         );
  NOR2_X1 U3725 ( .A1(n3605), .A2(n3604), .ZN(n3611) );
  NAND2_X1 U3726 ( .A1(n3592), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3605)
         );
  NAND2_X1 U3727 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3591) );
  OR2_X1 U3728 ( .A1(n5715), .A2(n4219), .ZN(n5686) );
  OR3_X1 U3729 ( .A1(n3045), .A2(n5737), .A3(n5486), .ZN(n3044) );
  NOR2_X2 U3730 ( .A1(n3002), .A2(n5698), .ZN(n5700) );
  NOR3_X1 U3731 ( .A1(n5736), .A2(n5737), .A3(n3046), .ZN(n5717) );
  NOR2_X1 U3732 ( .A1(n5736), .A2(n5737), .ZN(n5735) );
  NAND2_X1 U3733 ( .A1(n3072), .A2(n3001), .ZN(n3069) );
  NOR2_X1 U3734 ( .A1(n4146), .A2(n5870), .ZN(n5418) );
  NAND2_X1 U3735 ( .A1(n5592), .A2(n5911), .ZN(n5910) );
  NAND2_X1 U3736 ( .A1(n3043), .A2(n3042), .ZN(n5870) );
  INV_X1 U3737 ( .A(n5867), .ZN(n3042) );
  INV_X1 U3738 ( .A(n3043), .ZN(n5513) );
  OR2_X1 U3739 ( .A1(n5235), .A2(n5234), .ZN(n5252) );
  NAND2_X1 U3740 ( .A1(n5189), .A2(n5188), .ZN(n5235) );
  NAND2_X1 U3741 ( .A1(n4826), .A2(n3422), .ZN(n4559) );
  XNOR2_X1 U3742 ( .A(n3445), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4558)
         );
  INV_X1 U3743 ( .A(n4696), .ZN(n3049) );
  NAND2_X1 U3744 ( .A1(n3047), .A2(n4088), .ZN(n4697) );
  INV_X1 U3745 ( .A(n4433), .ZN(n3047) );
  AND2_X1 U3746 ( .A1(n3355), .A2(n3354), .ZN(n3323) );
  NAND2_X1 U3747 ( .A1(n3337), .A2(n3336), .ZN(n3401) );
  NAND2_X1 U3748 ( .A1(n3068), .A2(n3258), .ZN(n4487) );
  INV_X1 U3749 ( .A(n4259), .ZN(n4702) );
  AND2_X1 U3750 ( .A1(n4806), .A2(n4702), .ZN(n4710) );
  NAND2_X1 U3751 ( .A1(n6669), .A2(n4271), .ZN(n4742) );
  INV_X1 U3752 ( .A(n4742), .ZN(n4442) );
  AOI22_X1 U3753 ( .A1(n2982), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5283), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3144) );
  AND2_X1 U3754 ( .A1(n5329), .A2(n4271), .ZN(n4337) );
  INV_X1 U3755 ( .A(n4812), .ZN(n5016) );
  INV_X1 U3756 ( .A(n3035), .ZN(n4524) );
  NAND2_X1 U3757 ( .A1(n6150), .A2(n5804), .ZN(n6614) );
  AND2_X1 U3758 ( .A1(n6095), .A2(n4871), .ZN(n6066) );
  AND2_X1 U3759 ( .A1(n5359), .A2(n4877), .ZN(n6091) );
  AND2_X1 U3760 ( .A1(n5369), .A2(n4868), .ZN(n6072) );
  INV_X1 U3761 ( .A(n5886), .ZN(n6116) );
  NAND2_X1 U3762 ( .A1(n4303), .A2(n6118), .ZN(n5885) );
  AND2_X2 U3763 ( .A1(n4310), .A2(n6490), .ZN(n6118) );
  OR2_X1 U3764 ( .A1(n6122), .A2(n6126), .ZN(n5538) );
  NAND2_X1 U3765 ( .A1(n4641), .A2(n6226), .ZN(n5544) );
  OAI21_X1 U3766 ( .B1(n4638), .B2(n4637), .A(n6490), .ZN(n4641) );
  INV_X1 U3767 ( .A(n5538), .ZN(n5543) );
  BUF_X1 U3768 ( .A(n4600), .Z(n6609) );
  XNOR2_X1 U3769 ( .A(n5228), .B(n3733), .ZN(n5249) );
  AND2_X1 U3770 ( .A1(n4900), .A2(n3019), .ZN(n4903) );
  INV_X1 U3771 ( .A(n3489), .ZN(n3019) );
  AND2_X1 U3772 ( .A1(n4557), .A2(n3446), .ZN(n4915) );
  OR2_X1 U3773 ( .A1(n6257), .A2(n4031), .ZN(n5646) );
  NAND2_X1 U3774 ( .A1(n4649), .A2(n4650), .ZN(n4301) );
  NAND2_X1 U3775 ( .A1(n5646), .A2(n6275), .ZN(n6264) );
  INV_X1 U3776 ( .A(n5646), .ZN(n6276) );
  OR2_X1 U3777 ( .A1(n3021), .A2(n4043), .ZN(n3102) );
  AND2_X1 U3778 ( .A1(n5745), .A2(n4218), .ZN(n5726) );
  OAI21_X1 U3779 ( .B1(n5609), .B2(n5608), .A(n5607), .ZN(n5610) );
  NAND2_X1 U3780 ( .A1(n5917), .A2(n6692), .ZN(n5608) );
  NAND2_X1 U3781 ( .A1(n3074), .A2(n5594), .ZN(n5620) );
  AND2_X1 U3782 ( .A1(n5935), .A2(n4210), .ZN(n5926) );
  NAND2_X1 U3783 ( .A1(n5635), .A2(n3503), .ZN(n5643) );
  NAND2_X1 U3784 ( .A1(n5116), .A2(n3063), .ZN(n3058) );
  NAND2_X1 U3785 ( .A1(n5116), .A2(n5115), .ZN(n5208) );
  AND2_X1 U3786 ( .A1(n4204), .A2(n4185), .ZN(n6340) );
  INV_X1 U3787 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5005) );
  INV_X1 U3788 ( .A(n4817), .ZN(n4657) );
  INV_X1 U3789 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6365) );
  INV_X1 U3790 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6592) );
  INV_X1 U3791 ( .A(n4048), .ZN(n3242) );
  INV_X1 U3792 ( .A(n5182), .ZN(n5137) );
  NAND2_X1 U3793 ( .A1(n4710), .A2(n5008), .ZN(n4966) );
  NOR2_X1 U3794 ( .A1(n4647), .A2(n4742), .ZN(n6784) );
  NOR2_X1 U3795 ( .A1(n4653), .A2(n4742), .ZN(n6436) );
  NOR2_X1 U3796 ( .A1(n4782), .A2(n4742), .ZN(n6452) );
  NOR2_X1 U3797 ( .A1(n4654), .A2(n4742), .ZN(n6382) );
  INV_X1 U3798 ( .A(n6430), .ZN(n5097) );
  INV_X1 U3799 ( .A(n6422), .ZN(n5089) );
  INV_X1 U3800 ( .A(n6382), .ZN(n5084) );
  INV_X1 U3801 ( .A(n4468), .ZN(n4542) );
  NAND2_X1 U3802 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4480), .ZN(n6497) );
  OAI21_X1 U3803 ( .B1(n5671), .B2(n6079), .A(n3050), .ZN(U2797) );
  INV_X1 U3804 ( .A(n3051), .ZN(n3050) );
  NOR3_X1 U3805 ( .A1(n3054), .A2(n3053), .A3(n5365), .ZN(n3052) );
  NOR2_X1 U3806 ( .A1(n4040), .A2(n4039), .ZN(n4041) );
  NAND2_X1 U3807 ( .A1(n4038), .A2(n4037), .ZN(n4039) );
  AND2_X2 U3808 ( .A1(n4507), .A2(n4490), .ZN(n3307) );
  AND2_X2 U3809 ( .A1(n5340), .A2(n4507), .ZN(n3296) );
  OAI21_X1 U3810 ( .B1(n3068), .B2(n3258), .A(n4487), .ZN(n4261) );
  NOR2_X1 U3811 ( .A1(n4874), .A2(n4323), .ZN(n3237) );
  NAND2_X1 U3812 ( .A1(n3493), .A2(n5746), .ZN(n3001) );
  NAND2_X1 U3813 ( .A1(n3176), .A2(n4330), .ZN(n4187) );
  INV_X1 U3814 ( .A(n3078), .ZN(n3077) );
  NAND2_X1 U3815 ( .A1(n3011), .A2(n3503), .ZN(n3078) );
  NAND2_X2 U3816 ( .A1(n4076), .A2(n4874), .ZN(n4083) );
  OR2_X1 U3817 ( .A1(n5736), .A2(n3044), .ZN(n3002) );
  NAND2_X1 U3818 ( .A1(n3250), .A2(n3017), .ZN(n3068) );
  INV_X1 U3819 ( .A(n3020), .ZN(n5554) );
  NAND2_X1 U3820 ( .A1(n3021), .A2(n3008), .ZN(n3020) );
  AND2_X1 U3821 ( .A1(n5263), .A2(n3852), .ZN(n5414) );
  AND2_X1 U3822 ( .A1(n3182), .A2(n3105), .ZN(n3003) );
  OR3_X1 U3823 ( .A1(n5736), .A2(n5737), .A3(n3045), .ZN(n3004) );
  AND3_X1 U3824 ( .A1(n4315), .A2(n4874), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3274) );
  AND2_X1 U3825 ( .A1(n3074), .A2(n3071), .ZN(n3005) );
  AND2_X1 U3826 ( .A1(n3493), .A2(n5237), .ZN(n3006) );
  OR2_X1 U3827 ( .A1(n3393), .A2(n3378), .ZN(n3007) );
  NAND2_X1 U3828 ( .A1(n5569), .A2(n5568), .ZN(n5391) );
  NAND2_X1 U3829 ( .A1(n3167), .A2(n3104), .ZN(n3210) );
  INV_X1 U3830 ( .A(n3210), .ZN(n3176) );
  NAND2_X1 U3831 ( .A1(n5635), .A2(n3077), .ZN(n5634) );
  NAND2_X1 U3832 ( .A1(n3338), .A2(n3401), .ZN(n3079) );
  NAND2_X1 U3833 ( .A1(n3493), .A2(n3511), .ZN(n3008) );
  INV_X1 U3834 ( .A(n3241), .ZN(n3203) );
  NAND2_X1 U3835 ( .A1(n4901), .A2(n3492), .ZN(n5106) );
  NAND2_X1 U3836 ( .A1(n3058), .A2(n3496), .ZN(n5230) );
  NAND2_X1 U3837 ( .A1(n3208), .A2(n4645), .ZN(n4049) );
  AND2_X1 U3838 ( .A1(n3008), .A2(n5575), .ZN(n3009) );
  INV_X1 U3839 ( .A(n3099), .ZN(n3098) );
  NAND2_X1 U3840 ( .A1(n3931), .A2(n5603), .ZN(n3099) );
  AND2_X1 U3841 ( .A1(n3493), .A2(n4201), .ZN(n3010) );
  NAND2_X1 U3842 ( .A1(n3493), .A2(n5948), .ZN(n3011) );
  INV_X1 U3843 ( .A(n3072), .ZN(n3071) );
  NAND2_X1 U3844 ( .A1(n5594), .A2(n3073), .ZN(n3072) );
  INV_X1 U3845 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3034) );
  AND2_X1 U3846 ( .A1(n3087), .A2(n3086), .ZN(n3012) );
  AND2_X1 U3847 ( .A1(n3075), .A2(n3001), .ZN(n3013) );
  NOR2_X1 U3848 ( .A1(n3460), .A2(n3458), .ZN(n3014) );
  NOR2_X1 U3849 ( .A1(n5189), .A2(n5132), .ZN(n3015) );
  AND2_X1 U3850 ( .A1(n4494), .A2(n4874), .ZN(n4227) );
  NAND2_X1 U3851 ( .A1(n3570), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3847) );
  INV_X1 U3852 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6669) );
  AND2_X1 U3853 ( .A1(n3085), .A2(n3083), .ZN(n3016) );
  INV_X1 U3854 ( .A(n5408), .ZN(n3046) );
  INV_X1 U3855 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3663) );
  NAND2_X1 U3856 ( .A1(n3017), .A2(n3280), .ZN(n3281) );
  NAND2_X1 U3857 ( .A1(n3249), .A2(n3248), .ZN(n3017) );
  NAND2_X1 U3858 ( .A1(n3509), .A2(n3508), .ZN(n5555) );
  INV_X1 U3859 ( .A(n3021), .ZN(n5584) );
  NAND2_X1 U3860 ( .A1(n3024), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3246) );
  NAND3_X1 U3861 ( .A1(n3026), .A2(n5976), .A3(n3025), .ZN(n3024) );
  INV_X1 U3862 ( .A(n4183), .ZN(n3025) );
  NAND2_X1 U3863 ( .A1(n5635), .A2(n3027), .ZN(n5605) );
  NAND2_X2 U3864 ( .A1(n5653), .A2(n3502), .ZN(n5635) );
  NOR2_X1 U3865 ( .A1(n3031), .A2(n3030), .ZN(n3029) );
  INV_X1 U3866 ( .A(n3169), .ZN(n3031) );
  NAND2_X1 U3867 ( .A1(n3033), .A2(n3032), .ZN(n3472) );
  AND2_X1 U3868 ( .A1(n3014), .A2(n3424), .ZN(n3032) );
  AND2_X2 U3869 ( .A1(n3114), .A2(n3035), .ZN(n5283) );
  AND2_X2 U3870 ( .A1(n3034), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3114)
         );
  AND2_X4 U3871 ( .A1(n4500), .A2(n3035), .ZN(n3188) );
  NOR2_X2 U3872 ( .A1(n6052), .A2(n4109), .ZN(n5131) );
  NAND2_X2 U3873 ( .A1(n3003), .A2(n3039), .ZN(n4323) );
  NAND3_X1 U3874 ( .A1(n3184), .A2(n3186), .A3(n3183), .ZN(n3040) );
  NOR2_X2 U3875 ( .A1(n5511), .A2(n5510), .ZN(n3043) );
  NAND2_X1 U3876 ( .A1(n4088), .A2(n3049), .ZN(n3048) );
  NAND2_X1 U3877 ( .A1(n4087), .A2(n4086), .ZN(n4433) );
  OAI21_X1 U3878 ( .B1(n5116), .B2(n3061), .A(n3059), .ZN(n5258) );
  NAND2_X1 U3879 ( .A1(n3068), .A2(n3065), .ZN(n3066) );
  NAND2_X1 U3880 ( .A1(n5628), .A2(n3013), .ZN(n3070) );
  NAND2_X1 U3881 ( .A1(n5628), .A2(n3075), .ZN(n3074) );
  NAND2_X1 U3882 ( .A1(n4557), .A2(n3076), .ZN(n4913) );
  NAND2_X1 U3883 ( .A1(n4900), .A2(n3490), .ZN(n4901) );
  NAND2_X1 U3884 ( .A1(n3080), .A2(n3341), .ZN(n6254) );
  NAND3_X1 U3885 ( .A1(n3338), .A2(n3401), .A3(n3519), .ZN(n3080) );
  AND2_X2 U3886 ( .A1(n4506), .A2(n4500), .ZN(n3267) );
  AND2_X2 U3887 ( .A1(n5340), .A2(n4506), .ZN(n3157) );
  AND2_X2 U3888 ( .A1(n3107), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4506)
         );
  NAND2_X1 U3889 ( .A1(n5228), .A2(n3082), .ZN(n3081) );
  INV_X1 U3890 ( .A(n3733), .ZN(n3085) );
  NOR2_X2 U3891 ( .A1(n4781), .A2(n3625), .ZN(n4803) );
  CLKBUF_X1 U3892 ( .A(n5263), .Z(n5458) );
  AND4_X2 U3893 ( .A1(n3120), .A2(n3119), .A3(n3118), .A4(n3117), .ZN(n3121)
         );
  NAND2_X1 U3894 ( .A1(n3339), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3379) );
  NAND2_X1 U3895 ( .A1(n3339), .A2(n4323), .ZN(n4186) );
  AND2_X1 U3896 ( .A1(n3157), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3137) );
  AND2_X1 U3897 ( .A1(n3523), .A2(n4874), .ZN(n3224) );
  INV_X1 U3898 ( .A(n4645), .ZN(n4303) );
  OR2_X1 U3899 ( .A1(n5395), .A2(n4179), .ZN(n3100) );
  NOR2_X1 U3900 ( .A1(n4323), .A2(n4047), .ZN(n3101) );
  XNOR2_X1 U3901 ( .A(n3401), .B(n4284), .ZN(n3590) );
  NAND2_X1 U3902 ( .A1(n5544), .A2(n4643), .ZN(n5890) );
  AND3_X1 U3903 ( .A1(n5917), .A2(n5744), .A3(n6692), .ZN(n3103) );
  AND4_X1 U3904 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3104)
         );
  AND3_X1 U3905 ( .A1(n3181), .A2(n3180), .A3(n3179), .ZN(n3105) );
  NAND2_X1 U3906 ( .A1(n3444), .A2(n3443), .ZN(n4557) );
  INV_X1 U3907 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3627) );
  INV_X1 U3908 ( .A(n5582), .ZN(n3510) );
  NOR2_X1 U3909 ( .A1(n4645), .A2(n5007), .ZN(n3593) );
  AND2_X1 U3910 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3106) );
  INV_X1 U3911 ( .A(n3559), .ZN(n3527) );
  OAI21_X1 U3912 ( .B1(n3527), .B2(n3523), .A(n3155), .ZN(n3535) );
  AND2_X1 U3913 ( .A1(n5005), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3525)
         );
  INV_X1 U3914 ( .A(n4187), .ZN(n3177) );
  AND3_X1 U3915 ( .A1(n3329), .A2(n3328), .A3(n3327), .ZN(n3330) );
  OR2_X1 U3916 ( .A1(n3434), .A2(n3433), .ZN(n3463) );
  AND2_X1 U3917 ( .A1(n3232), .A2(n3231), .ZN(n3233) );
  AOI22_X1 U3918 ( .A1(n2988), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n2974), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3175) );
  NOR2_X1 U3919 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3115) );
  XNOR2_X1 U3920 ( .A(n3472), .B(n3471), .ZN(n3626) );
  OR2_X1 U3921 ( .A1(n3390), .A2(n3389), .ZN(n3416) );
  OR3_X1 U3922 ( .A1(n3556), .A2(n6365), .A3(INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .ZN(n4061) );
  NAND2_X1 U3923 ( .A1(n3415), .A2(n3414), .ZN(n3424) );
  AND2_X1 U3924 ( .A1(n3849), .A2(n5439), .ZN(n5440) );
  NAND2_X1 U3925 ( .A1(n3713), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3714)
         );
  NAND2_X1 U3926 ( .A1(n3626), .A2(n3732), .ZN(n3633) );
  AND2_X1 U3927 ( .A1(n4095), .A2(n4094), .ZN(n4311) );
  NAND2_X1 U3928 ( .A1(n2981), .A2(n3519), .ZN(n3563) );
  INV_X1 U3929 ( .A(n3593), .ZN(n3594) );
  OR2_X1 U3930 ( .A1(n3932), .A2(n5406), .ZN(n3933) );
  AND2_X1 U3931 ( .A1(n3850), .A2(n5440), .ZN(n5426) );
  INV_X1 U3932 ( .A(n3847), .ZN(n3732) );
  NAND2_X1 U3933 ( .A1(n3442), .A2(n3441), .ZN(n3445) );
  NAND2_X1 U3934 ( .A1(n5606), .A2(n3493), .ZN(n5607) );
  OR2_X1 U3935 ( .A1(n3563), .A2(n3562), .ZN(n3564) );
  NAND2_X1 U3936 ( .A1(n3885), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3886)
         );
  NAND2_X1 U3937 ( .A1(n3843), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3818)
         );
  INV_X1 U3938 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5195) );
  INV_X1 U3939 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4896) );
  INV_X1 U3940 ( .A(n6053), .ZN(n6093) );
  NAND2_X1 U3941 ( .A1(n5359), .A2(n4870), .ZN(n5448) );
  INV_X1 U3942 ( .A(n3926), .ZN(n5350) );
  NOR2_X1 U3943 ( .A1(n3853), .A2(n5622), .ZN(n3885) );
  OR2_X1 U3944 ( .A1(n5507), .A2(n5506), .ZN(n5508) );
  INV_X1 U3945 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3604) );
  INV_X1 U3946 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U3947 ( .A1(n5615), .A2(n5595), .ZN(n5596) );
  INV_X1 U3948 ( .A(n6340), .ZN(n6358) );
  OAI21_X1 U3949 ( .B1(n6617), .B2(n4528), .A(n6497), .ZN(n4271) );
  AND2_X1 U3950 ( .A1(n5016), .A2(n5015), .ZN(n5046) );
  AND2_X1 U3951 ( .A1(n3079), .A2(n4817), .ZN(n4806) );
  INV_X1 U3952 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4704) );
  OR2_X1 U3953 ( .A1(n4389), .A2(n5008), .ZN(n6787) );
  NAND2_X1 U3954 ( .A1(n4296), .A2(n5008), .ZN(n4690) );
  INV_X1 U3955 ( .A(n4034), .ZN(n6613) );
  AND2_X1 U3956 ( .A1(n3969), .A2(n3968), .ZN(n3988) );
  NOR2_X1 U3957 ( .A1(n6563), .A2(n5834), .ZN(n5823) );
  INV_X1 U3958 ( .A(n5872), .ZN(n6064) );
  INV_X1 U3959 ( .A(n6055), .ZN(n6070) );
  AND2_X1 U3960 ( .A1(n6084), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6053) );
  INV_X1 U3961 ( .A(n5885), .ZN(n6115) );
  INV_X1 U3962 ( .A(n5890), .ZN(n6123) );
  INV_X1 U3963 ( .A(n5544), .ZN(n6125) );
  NAND2_X1 U3964 ( .A1(n6149), .A2(n4640), .ZN(n6226) );
  AOI21_X1 U3965 ( .B1(n5442), .B2(n5509), .A(n5441), .ZN(n6119) );
  INV_X1 U3966 ( .A(n3591), .ZN(n3592) );
  OR2_X1 U3967 ( .A1(n4222), .A2(n4045), .ZN(n4223) );
  OAI21_X1 U3968 ( .B1(n5615), .B2(n3103), .A(n5596), .ZN(n5597) );
  NOR2_X1 U3969 ( .A1(n6282), .A2(n4208), .ZN(n5935) );
  NAND2_X1 U3970 ( .A1(n5118), .A2(n5123), .ZN(n5789) );
  NOR3_X1 U3971 ( .A1(n4198), .A2(n5123), .A3(n5125), .ZN(n5952) );
  NAND2_X1 U3972 ( .A1(n4204), .A2(n4232), .ZN(n5123) );
  INV_X1 U3973 ( .A(n5123), .ZN(n6341) );
  AND2_X1 U3974 ( .A1(n4204), .A2(n4075), .ZN(n6354) );
  INV_X1 U3975 ( .A(n4807), .ZN(n5799) );
  OR2_X1 U3976 ( .A1(n4662), .A2(n4661), .ZN(n4689) );
  AND2_X1 U3977 ( .A1(n4657), .A2(n4656), .ZN(n5009) );
  INV_X1 U3978 ( .A(n6387), .ZN(n5179) );
  INV_X1 U3979 ( .A(n4793), .ZN(n4787) );
  INV_X1 U3980 ( .A(n4635), .ZN(n6401) );
  INV_X1 U3981 ( .A(n4966), .ZN(n4993) );
  AND2_X1 U3982 ( .A1(n4818), .A2(n4817), .ZN(n6459) );
  INV_X1 U3983 ( .A(n4703), .ZN(n5008) );
  AND2_X1 U3984 ( .A1(n4296), .A2(n4703), .ZN(n4468) );
  NOR2_X1 U3985 ( .A1(n6689), .A2(n4742), .ZN(n6430) );
  NOR2_X1 U3986 ( .A1(n6161), .A2(n4742), .ZN(n6422) );
  INV_X1 U3987 ( .A(n6091), .ZN(n6080) );
  OR2_X1 U3988 ( .A1(n5369), .A2(n4867), .ZN(n5872) );
  NAND2_X1 U3989 ( .A1(n6118), .A2(n4645), .ZN(n5886) );
  INV_X1 U3990 ( .A(n4908), .ZN(n4910) );
  NOR2_X1 U3991 ( .A1(n6609), .A2(n6129), .ZN(n5802) );
  INV_X1 U3992 ( .A(n6129), .ZN(n6147) );
  OR2_X1 U3993 ( .A1(n5604), .A2(n5495), .ZN(n5843) );
  OR2_X1 U3994 ( .A1(n5461), .A2(n5507), .ZN(n5652) );
  INV_X1 U3995 ( .A(n6257), .ZN(n6273) );
  OR2_X1 U3996 ( .A1(n6509), .A2(n5799), .ZN(n6271) );
  AND2_X1 U3997 ( .A1(n5754), .A2(n4215), .ZN(n5745) );
  NOR2_X1 U3998 ( .A1(n5952), .A2(n5232), .ZN(n6282) );
  INV_X1 U3999 ( .A(n6354), .ZN(n6313) );
  INV_X1 U4000 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U4001 ( .A1(n5009), .A2(n4703), .ZN(n5052) );
  NAND2_X1 U4002 ( .A1(n5009), .A2(n5008), .ZN(n5182) );
  NAND2_X1 U4003 ( .A1(n4816), .A2(n4657), .ZN(n6387) );
  NOR2_X1 U4004 ( .A1(n4572), .A2(n4571), .ZN(n4783) );
  INV_X1 U4005 ( .A(n4265), .ZN(n4374) );
  OR2_X1 U4006 ( .A1(n4616), .A2(n4615), .ZN(n6426) );
  NAND2_X1 U4007 ( .A1(n4710), .A2(n4703), .ZN(n4779) );
  INV_X1 U4008 ( .A(n6461), .ZN(n5174) );
  NAND2_X1 U4009 ( .A1(n4816), .A2(n4817), .ZN(n6465) );
  AND2_X1 U4010 ( .A1(n5057), .A2(n5056), .ZN(n5105) );
  NAND2_X1 U4011 ( .A1(n4383), .A2(n5008), .ZN(n6793) );
  AND2_X1 U4012 ( .A1(n4440), .A2(n4439), .ZN(n4540) );
  INV_X1 U4013 ( .A(n6784), .ZN(n5070) );
  INV_X1 U4014 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6589) );
  NOR2_X4 U4015 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U4016 ( .A1(n5283), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3113) );
  INV_X1 U4017 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3107) );
  AOI22_X1 U4018 ( .A1(n3193), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3112) );
  AOI22_X1 U4019 ( .A1(n3000), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3111) );
  AND4_X2 U4020 ( .A1(n3113), .A2(n3112), .A3(n3111), .A4(n3110), .ZN(n3122)
         );
  AOI22_X1 U4021 ( .A1(n3296), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U4022 ( .A1(n2974), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U4023 ( .A1(n3307), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U4024 ( .A1(n2995), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3117) );
  AOI22_X1 U4025 ( .A1(n3193), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U4026 ( .A1(n2986), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U4027 ( .A1(n5283), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3124) );
  AOI22_X1 U4028 ( .A1(n3000), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U4029 ( .A1(n3296), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U4030 ( .A1(n3307), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U4031 ( .A1(n2975), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4032 ( .A1(n2995), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U4033 ( .A1(n2975), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3136) );
  AOI22_X1 U4034 ( .A1(n3259), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4035 ( .A1(n3000), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4036 ( .A1(n5283), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3133) );
  NAND4_X1 U4037 ( .A1(n3136), .A2(n3135), .A3(n3134), .A4(n3133), .ZN(n3143)
         );
  AOI22_X1 U4038 ( .A1(n2992), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2982), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U4039 ( .A1(n3307), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4040 ( .A1(n3296), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3138) );
  NAND4_X1 U4041 ( .A1(n3141), .A2(n3140), .A3(n3139), .A4(n3138), .ZN(n3142)
         );
  NAND2_X1 U4042 ( .A1(n3241), .A2(n4645), .ZN(n3154) );
  AOI22_X1 U4043 ( .A1(n2974), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4044 ( .A1(n3266), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4045 ( .A1(n3193), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3145) );
  NAND4_X1 U4046 ( .A1(n3147), .A2(n3146), .A3(n3145), .A4(n3144), .ZN(n3153)
         );
  AOI22_X1 U4047 ( .A1(n3307), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4048 ( .A1(n3265), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U4049 ( .A1(n2995), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4050 ( .A1(n3296), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3148) );
  NAND4_X1 U4051 ( .A1(n3151), .A2(n3150), .A3(n3149), .A4(n3148), .ZN(n3152)
         );
  OR2_X2 U4052 ( .A1(n3153), .A2(n3152), .ZN(n4319) );
  NAND2_X1 U4053 ( .A1(n3154), .A2(n3239), .ZN(n3156) );
  NAND2_X1 U4054 ( .A1(n3156), .A2(n3209), .ZN(n3228) );
  INV_X1 U4055 ( .A(n3228), .ZN(n3178) );
  AOI22_X1 U4056 ( .A1(n3193), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4057 ( .A1(n3380), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4058 ( .A1(n2979), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4059 ( .A1(n3296), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4060 ( .A1(n2995), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4061 ( .A1(n2992), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4062 ( .A1(n3259), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4063 ( .A1(n5283), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4064 ( .A1(n3193), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4065 ( .A1(n3380), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4066 ( .A1(n5283), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4067 ( .A1(n2982), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4068 ( .A1(n3307), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4069 ( .A1(n3296), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4070 ( .A1(n2995), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3172) );
  NAND2_X1 U4071 ( .A1(n3178), .A2(n3177), .ZN(n3567) );
  AOI22_X1 U4072 ( .A1(n5283), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4073 ( .A1(n2986), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5284), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4074 ( .A1(n3380), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U4075 ( .A1(n2980), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4076 ( .A1(n3307), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4077 ( .A1(n2995), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4078 ( .A1(n3296), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3185) );
  XNOR2_X1 U4079 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4054) );
  NAND2_X1 U4080 ( .A1(n3523), .A2(n4054), .ZN(n3240) );
  NAND2_X1 U4081 ( .A1(n3240), .A2(n3214), .ZN(n3201) );
  AOI22_X1 U4082 ( .A1(n2995), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U4083 ( .A1(n3000), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4084 ( .A1(n3307), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3190) );
  AOI22_X1 U4085 ( .A1(n5283), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3189) );
  NAND4_X1 U4086 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n3200)
         );
  AOI22_X1 U4087 ( .A1(n3193), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3157), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4088 ( .A1(n3296), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4089 ( .A1(n2979), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3196) );
  NAND4_X1 U4090 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3199)
         );
  NAND2_X1 U4091 ( .A1(n3201), .A2(n4186), .ZN(n3202) );
  NOR2_X1 U4092 ( .A1(n3567), .A2(n3202), .ZN(n3206) );
  NAND2_X1 U4094 ( .A1(n4049), .A2(n3224), .ZN(n3205) );
  NAND2_X1 U4095 ( .A1(n3204), .A2(n3203), .ZN(n4195) );
  NAND2_X1 U4096 ( .A1(n3206), .A2(n3231), .ZN(n3207) );
  NAND2_X1 U4097 ( .A1(n3207), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3218) );
  NAND3_X1 U4098 ( .A1(n3208), .A2(n3223), .A3(n3210), .ZN(n3213) );
  OAI21_X1 U4099 ( .B1(n4304), .B2(n4319), .A(n3209), .ZN(n3211) );
  NAND2_X1 U4100 ( .A1(n3213), .A2(n3212), .ZN(n3215) );
  NAND2_X1 U4101 ( .A1(n4642), .A2(n4330), .ZN(n3225) );
  NAND2_X1 U4102 ( .A1(n3218), .A2(n3217), .ZN(n3251) );
  NAND2_X1 U4103 ( .A1(n3251), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4104 ( .A1(n6592), .A2(n6589), .ZN(n6597) );
  MUX2_X1 U4105 ( .A(n3255), .B(n6613), .S(n5005), .Z(n3219) );
  INV_X1 U4106 ( .A(n3219), .ZN(n3220) );
  INV_X1 U4107 ( .A(n4186), .ZN(n4923) );
  AND2_X1 U4108 ( .A1(n3210), .A2(n4874), .ZN(n3222) );
  OR2_X1 U4109 ( .A1(n6597), .A2(n6669), .ZN(n6503) );
  INV_X1 U4110 ( .A(n6503), .ZN(n3227) );
  NAND4_X1 U4111 ( .A1(n3339), .A2(n3575), .A3(n4305), .A4(n4315), .ZN(n4515)
         );
  NAND2_X1 U4112 ( .A1(n3225), .A2(n3224), .ZN(n3226) );
  INV_X1 U4113 ( .A(n3237), .ZN(n4922) );
  NAND2_X1 U4114 ( .A1(n4048), .A2(n3237), .ZN(n4192) );
  NAND2_X1 U4115 ( .A1(n4642), .A2(n4315), .ZN(n3229) );
  NAND2_X1 U4116 ( .A1(n3229), .A2(n4330), .ZN(n3230) );
  OAI21_X1 U4117 ( .B1(n3228), .B2(n3230), .A(n4323), .ZN(n3232) );
  INV_X1 U4118 ( .A(n3294), .ZN(n3235) );
  INV_X1 U4119 ( .A(n4330), .ZN(n4076) );
  AND3_X1 U4120 ( .A1(n3214), .A2(n3176), .A3(n4076), .ZN(n3238) );
  NAND2_X1 U4121 ( .A1(n3238), .A2(n3237), .ZN(n4492) );
  NOR2_X1 U4122 ( .A1(n4492), .A2(n3239), .ZN(n4183) );
  XNOR2_X1 U4123 ( .A(n4704), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5141)
         );
  NAND2_X1 U4124 ( .A1(n6613), .A2(n5141), .ZN(n3244) );
  NAND2_X1 U4125 ( .A1(n3255), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3243) );
  NAND2_X1 U4126 ( .A1(n3244), .A2(n3243), .ZN(n3247) );
  AOI21_X1 U4127 ( .B1(n3251), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3247), 
        .ZN(n3245) );
  NAND2_X1 U4128 ( .A1(n3246), .A2(n3245), .ZN(n3280) );
  NAND2_X1 U4129 ( .A1(n3279), .A2(n3280), .ZN(n3250) );
  INV_X1 U4130 ( .A(n3246), .ZN(n3249) );
  NAND2_X1 U4131 ( .A1(n3251), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3257) );
  AND2_X1 U4132 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3252) );
  NAND2_X1 U4133 ( .A1(n3252), .A2(n6478), .ZN(n4810) );
  INV_X1 U4134 ( .A(n3252), .ZN(n3253) );
  NAND2_X1 U4135 ( .A1(n3253), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3254) );
  NAND2_X1 U4136 ( .A1(n4810), .A2(n3254), .ZN(n4443) );
  AOI22_X1 U4137 ( .A1(n6613), .A2(n4443), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3255), .ZN(n3256) );
  AOI22_X1 U4138 ( .A1(n2994), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4139 ( .A1(n3380), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4140 ( .A1(n5283), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4141 ( .A1(n2982), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3261) );
  NAND4_X1 U4142 ( .A1(n3264), .A2(n3263), .A3(n3262), .A4(n3261), .ZN(n3273)
         );
  AOI22_X1 U4143 ( .A1(n3308), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4144 ( .A1(n5285), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3270) );
  INV_X1 U4145 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6722) );
  AOI22_X1 U4146 ( .A1(n2980), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4147 ( .A1(n2995), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3268) );
  NAND4_X1 U4148 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), .ZN(n3272)
         );
  AOI22_X1 U4149 ( .A1(n3276), .A2(n3275), .B1(n2981), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3277) );
  INV_X1 U4150 ( .A(n3337), .ZN(n3335) );
  NAND2_X1 U4151 ( .A1(n4262), .A2(n6669), .ZN(n3293) );
  AOI22_X1 U4152 ( .A1(n2975), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4153 ( .A1(n4014), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4154 ( .A1(n3308), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4155 ( .A1(n3000), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3282) );
  NAND4_X1 U4156 ( .A1(n3285), .A2(n3284), .A3(n3283), .A4(n3282), .ZN(n3291)
         );
  AOI22_X1 U4157 ( .A1(n3259), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4158 ( .A1(n2994), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4159 ( .A1(n3267), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4160 ( .A1(n3992), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3286) );
  NAND4_X1 U4161 ( .A1(n3289), .A2(n3288), .A3(n3287), .A4(n3286), .ZN(n3290)
         );
  OR2_X1 U4162 ( .A1(n3378), .A2(n3326), .ZN(n3292) );
  NAND2_X1 U4163 ( .A1(n3293), .A2(n3292), .ZN(n3344) );
  INV_X1 U4164 ( .A(n3344), .ZN(n3333) );
  AOI22_X1 U4165 ( .A1(n2994), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4166 ( .A1(n3308), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4167 ( .A1(n2975), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4168 ( .A1(n3267), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3297) );
  NAND4_X1 U4169 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3306)
         );
  AOI22_X1 U4170 ( .A1(n3000), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3259), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4171 ( .A1(n2991), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4172 ( .A1(n4014), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4173 ( .A1(n2982), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3301) );
  NAND4_X1 U4174 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3305)
         );
  AOI22_X1 U4175 ( .A1(n4014), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4176 ( .A1(n2994), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4177 ( .A1(n2974), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4178 ( .A1(n3308), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3309) );
  NAND4_X1 U4179 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3318)
         );
  AOI22_X1 U4180 ( .A1(n2995), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2986), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4181 ( .A1(n3265), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4182 ( .A1(n3259), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4183 ( .A1(n3157), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3313) );
  NAND4_X1 U4184 ( .A1(n3316), .A2(n3315), .A3(n3314), .A4(n3313), .ZN(n3317)
         );
  XNOR2_X1 U4185 ( .A(n3484), .B(n3360), .ZN(n3319) );
  NOR2_X1 U4186 ( .A1(n3319), .A2(n3378), .ZN(n3355) );
  INV_X1 U4187 ( .A(n3360), .ZN(n3322) );
  NAND2_X1 U4188 ( .A1(n2981), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3321) );
  AOI21_X1 U4189 ( .B1(n4304), .B2(n3484), .A(n6669), .ZN(n3320) );
  OAI211_X1 U4190 ( .C1(n3322), .C2(n4874), .A(n3321), .B(n3320), .ZN(n3354)
         );
  INV_X1 U4191 ( .A(n3484), .ZN(n3324) );
  OR2_X1 U4192 ( .A1(n3378), .A2(n3324), .ZN(n3325) );
  OR2_X1 U4193 ( .A1(n3378), .A2(n3484), .ZN(n3329) );
  OR2_X1 U4194 ( .A1(n3379), .A2(n3326), .ZN(n3328) );
  NAND2_X1 U4195 ( .A1(n2981), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3327) );
  OR2_X2 U4196 ( .A1(n3331), .A2(n3330), .ZN(n3343) );
  AOI21_X2 U4197 ( .B1(n3333), .B2(n3343), .A(n3332), .ZN(n3336) );
  INV_X1 U4198 ( .A(n3336), .ZN(n3334) );
  NAND2_X1 U4199 ( .A1(n3335), .A2(n3334), .ZN(n3338) );
  NAND2_X1 U4200 ( .A1(n3348), .A2(n3360), .ZN(n3394) );
  XNOR2_X1 U4201 ( .A(n3394), .B(n3393), .ZN(n3340) );
  AND2_X1 U4202 ( .A1(n3339), .A2(n4330), .ZN(n3358) );
  AOI21_X1 U4203 ( .B1(n3340), .B2(n6152), .A(n3358), .ZN(n3341) );
  NAND2_X1 U4204 ( .A1(n3343), .A2(n3342), .ZN(n3345) );
  NAND2_X1 U4205 ( .A1(n3345), .A2(n3344), .ZN(n3346) );
  NAND2_X1 U4206 ( .A1(n4259), .A2(n3519), .ZN(n3352) );
  OAI21_X1 U4207 ( .B1(n3360), .B2(n3348), .A(n3394), .ZN(n3349) );
  INV_X1 U4208 ( .A(n6152), .ZN(n6616) );
  OAI211_X1 U4209 ( .C1(n3349), .C2(n6616), .A(n3177), .B(n3155), .ZN(n3350)
         );
  INV_X1 U4210 ( .A(n3350), .ZN(n3351) );
  NAND2_X1 U4211 ( .A1(n3352), .A2(n3351), .ZN(n4277) );
  INV_X1 U4212 ( .A(n3353), .ZN(n3357) );
  NOR2_X1 U4213 ( .A1(n3355), .A2(n3354), .ZN(n3356) );
  INV_X1 U4214 ( .A(n3519), .ZN(n3363) );
  INV_X1 U4215 ( .A(n3358), .ZN(n3359) );
  OAI21_X1 U4216 ( .B1(n6616), .B2(n3360), .A(n3359), .ZN(n3361) );
  INV_X1 U4217 ( .A(n3361), .ZN(n3362) );
  NAND2_X1 U4218 ( .A1(n6269), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3364)
         );
  INV_X1 U4219 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U4220 ( .A1(n3364), .A2(n5324), .ZN(n3366) );
  AND2_X1 U4221 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U4222 ( .A1(n6269), .A2(n3365), .ZN(n3367) );
  AND2_X1 U4223 ( .A1(n3366), .A2(n3367), .ZN(n4276) );
  INV_X1 U4224 ( .A(n3367), .ZN(n3368) );
  NAND2_X1 U4225 ( .A1(n3369), .A2(n6255), .ZN(n3373) );
  INV_X1 U4226 ( .A(n6254), .ZN(n3371) );
  INV_X1 U4227 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U4228 ( .A1(n3371), .A2(n3370), .ZN(n3372) );
  AND2_X1 U4229 ( .A1(n3373), .A2(n3372), .ZN(n6247) );
  NAND2_X1 U4230 ( .A1(n3251), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3377) );
  NOR3_X1 U4231 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6478), .A3(n4704), 
        .ZN(n4844) );
  NAND2_X1 U4232 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4844), .ZN(n6417) );
  NAND2_X1 U4233 ( .A1(n6768), .A2(n6417), .ZN(n3374) );
  NAND3_X1 U4234 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4441) );
  INV_X1 U4235 ( .A(n4441), .ZN(n4293) );
  NAND2_X1 U4236 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4293), .ZN(n4338) );
  NAND2_X1 U4237 ( .A1(n3374), .A2(n4338), .ZN(n4741) );
  OAI22_X1 U4238 ( .A1(n4034), .A2(n4741), .B1(n3566), .B2(n6768), .ZN(n3375)
         );
  INV_X1 U4239 ( .A(n3375), .ZN(n3376) );
  XNOR2_X1 U4240 ( .A(n4487), .B(n4263), .ZN(n4286) );
  AOI22_X1 U4241 ( .A1(n2974), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4242 ( .A1(n3308), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4243 ( .A1(n5283), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4244 ( .A1(n2995), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3381) );
  NAND4_X1 U4245 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3390)
         );
  AOI22_X1 U4246 ( .A1(n3157), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4247 ( .A1(n3265), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4248 ( .A1(n5282), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4249 ( .A1(n2994), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3385) );
  NAND4_X1 U4250 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), .ZN(n3389)
         );
  AOI22_X1 U4251 ( .A1(n3559), .A2(n3416), .B1(n2981), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4252 ( .A1(n3590), .A2(n3519), .ZN(n3398) );
  NAND2_X1 U4253 ( .A1(n3394), .A2(n3393), .ZN(n3417) );
  INV_X1 U4254 ( .A(n3416), .ZN(n3395) );
  XNOR2_X1 U4255 ( .A(n3417), .B(n3395), .ZN(n3396) );
  NAND2_X1 U4256 ( .A1(n3396), .A2(n6152), .ZN(n3397) );
  INV_X1 U4257 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6336) );
  XNOR2_X1 U4258 ( .A(n3399), .B(n6336), .ZN(n6248) );
  NAND2_X1 U4259 ( .A1(n6247), .A2(n6248), .ZN(n6246) );
  NAND2_X1 U4260 ( .A1(n3399), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3400)
         );
  NAND2_X1 U4261 ( .A1(n6246), .A2(n3400), .ZN(n4828) );
  INV_X1 U4262 ( .A(n3401), .ZN(n3402) );
  AOI22_X1 U4263 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3308), .B1(n3265), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4264 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3873), .B1(n3403), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4265 ( .A1(n3267), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4266 ( .A1(n5282), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3404) );
  NAND4_X1 U4267 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(n3413)
         );
  AOI22_X1 U4268 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4014), .B1(n3380), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4269 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n2994), .B1(n2984), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4270 ( .A1(n2975), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4271 ( .A1(n5285), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3408) );
  NAND4_X1 U4272 ( .A1(n3411), .A2(n3410), .A3(n3409), .A4(n3408), .ZN(n3412)
         );
  NAND2_X1 U4273 ( .A1(n3559), .A2(n3437), .ZN(n3415) );
  NAND2_X1 U4274 ( .A1(n2981), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3414) );
  NAND2_X1 U4275 ( .A1(n3609), .A2(n3519), .ZN(n3420) );
  NAND2_X1 U4276 ( .A1(n3417), .A2(n3416), .ZN(n3439) );
  XNOR2_X1 U4277 ( .A(n3439), .B(n3437), .ZN(n3418) );
  NAND2_X1 U4278 ( .A1(n3418), .A2(n6152), .ZN(n3419) );
  NAND2_X1 U4279 ( .A1(n3420), .A2(n3419), .ZN(n3421) );
  INV_X1 U4280 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6328) );
  XNOR2_X1 U4281 ( .A(n3421), .B(n6328), .ZN(n4827) );
  NAND2_X1 U4282 ( .A1(n4828), .A2(n4827), .ZN(n4826) );
  NAND2_X1 U4283 ( .A1(n3421), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3422)
         );
  INV_X1 U4284 ( .A(n4559), .ZN(n3444) );
  AOI22_X1 U4285 ( .A1(n2994), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4286 ( .A1(n3380), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4287 ( .A1(n4014), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4288 ( .A1(n3403), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3425) );
  NAND4_X1 U4289 ( .A1(n3428), .A2(n3427), .A3(n3426), .A4(n3425), .ZN(n3434)
         );
  AOI22_X1 U4290 ( .A1(n3308), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4291 ( .A1(n5285), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4292 ( .A1(n2979), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4293 ( .A1(n3267), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3429) );
  NAND4_X1 U4294 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3433)
         );
  NAND2_X1 U4295 ( .A1(n3559), .A2(n3463), .ZN(n3436) );
  NAND2_X1 U4296 ( .A1(n2981), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U4297 ( .A1(n3436), .A2(n3435), .ZN(n3457) );
  NAND2_X1 U4298 ( .A1(n3610), .A2(n3519), .ZN(n3442) );
  INV_X1 U4299 ( .A(n3437), .ZN(n3438) );
  OR2_X1 U4300 ( .A1(n3439), .A2(n3438), .ZN(n3462) );
  XNOR2_X1 U4301 ( .A(n3462), .B(n3463), .ZN(n3440) );
  NAND2_X1 U4302 ( .A1(n3440), .A2(n6152), .ZN(n3441) );
  INV_X1 U4303 ( .A(n4558), .ZN(n3443) );
  OR2_X1 U4304 ( .A1(n3445), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3446)
         );
  AOI22_X1 U4305 ( .A1(n2994), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4306 ( .A1(n3000), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4307 ( .A1(n4014), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4308 ( .A1(n3403), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3447) );
  NAND4_X1 U4309 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3456)
         );
  AOI22_X1 U4310 ( .A1(n3308), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4311 ( .A1(n5285), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4312 ( .A1(n2974), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4313 ( .A1(n2995), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3451) );
  NAND4_X1 U4314 ( .A1(n3454), .A2(n3453), .A3(n3452), .A4(n3451), .ZN(n3455)
         );
  AOI22_X1 U4315 ( .A1(n3559), .A2(n3474), .B1(n2981), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3460) );
  INV_X1 U4316 ( .A(n3457), .ZN(n3458) );
  NAND2_X1 U4317 ( .A1(n3461), .A2(n3460), .ZN(n3618) );
  NAND3_X1 U4318 ( .A1(n3472), .A2(n3519), .A3(n3618), .ZN(n3467) );
  INV_X1 U4319 ( .A(n3462), .ZN(n3464) );
  NAND2_X1 U4320 ( .A1(n3464), .A2(n3463), .ZN(n3473) );
  XNOR2_X1 U4321 ( .A(n3473), .B(n3474), .ZN(n3465) );
  NAND2_X1 U4322 ( .A1(n3465), .A2(n6152), .ZN(n3466) );
  INV_X1 U4323 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U4324 ( .A1(n3468), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6232)
         );
  NAND2_X1 U4325 ( .A1(n3559), .A2(n3484), .ZN(n3470) );
  NAND2_X1 U4326 ( .A1(n2981), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U4327 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  NAND2_X1 U4328 ( .A1(n3626), .A2(n3519), .ZN(n3478) );
  INV_X1 U4329 ( .A(n3473), .ZN(n3475) );
  NAND2_X1 U4330 ( .A1(n3475), .A2(n3474), .ZN(n3486) );
  XNOR2_X1 U4331 ( .A(n3486), .B(n3484), .ZN(n3476) );
  NAND2_X1 U4332 ( .A1(n3476), .A2(n6152), .ZN(n3477) );
  NAND2_X1 U4333 ( .A1(n3478), .A2(n3477), .ZN(n3480) );
  NAND2_X1 U4334 ( .A1(n3480), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3481)
         );
  AND2_X1 U4335 ( .A1(n6232), .A2(n3481), .ZN(n3479) );
  INV_X1 U4336 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6305) );
  XNOR2_X1 U4337 ( .A(n3480), .B(n6305), .ZN(n6233) );
  INV_X1 U4338 ( .A(n3481), .ZN(n3482) );
  AND2_X1 U4339 ( .A1(n3519), .A2(n3484), .ZN(n3483) );
  NAND2_X4 U4340 ( .A1(n3472), .A2(n3483), .ZN(n3493) );
  NAND2_X1 U4341 ( .A1(n6152), .A2(n3484), .ZN(n3485) );
  OR2_X1 U4342 ( .A1(n3486), .A2(n3485), .ZN(n3487) );
  NAND2_X1 U4343 ( .A1(n3493), .A2(n3487), .ZN(n3491) );
  INV_X1 U4344 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6299) );
  XNOR2_X1 U4345 ( .A(n3491), .B(n6299), .ZN(n4902) );
  INV_X1 U4346 ( .A(n4902), .ZN(n3488) );
  NOR2_X1 U4347 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  NAND2_X1 U4348 ( .A1(n3491), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3492)
         );
  INV_X1 U4349 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U4350 ( .A1(n3493), .A2(n5126), .ZN(n5107) );
  NAND2_X1 U4351 ( .A1(n5917), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5108)
         );
  INV_X1 U4352 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3494) );
  NAND2_X1 U4353 ( .A1(n3493), .A2(n3494), .ZN(n5115) );
  INV_X1 U4354 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5209) );
  AND2_X1 U4355 ( .A1(n3493), .A2(n5209), .ZN(n3497) );
  NAND2_X1 U4356 ( .A1(n5917), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U4357 ( .A1(n5917), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3495) );
  INV_X1 U4358 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5237) );
  XNOR2_X1 U4359 ( .A(n3493), .B(n5237), .ZN(n5231) );
  XNOR2_X1 U4360 ( .A(n3493), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5257)
         );
  INV_X1 U4361 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U4362 ( .A1(n3493), .A2(n5974), .ZN(n3498) );
  NAND2_X1 U4363 ( .A1(n5256), .A2(n3498), .ZN(n5659) );
  NAND2_X1 U4364 ( .A1(n5917), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3499) );
  NAND2_X1 U4365 ( .A1(n5659), .A2(n3499), .ZN(n3501) );
  INV_X1 U4366 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6653) );
  NAND2_X1 U4367 ( .A1(n3493), .A2(n6653), .ZN(n3500) );
  NAND2_X1 U4368 ( .A1(n3501), .A2(n3500), .ZN(n5653) );
  NAND2_X1 U4369 ( .A1(n5917), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3502) );
  INV_X1 U4370 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U4371 ( .A1(n3493), .A2(n5942), .ZN(n3503) );
  INV_X1 U4372 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U4373 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4201) );
  INV_X1 U4374 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5764) );
  INV_X1 U4375 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5939) );
  NAND3_X1 U4376 ( .A1(n5764), .A2(n5948), .A3(n5939), .ZN(n3504) );
  NAND2_X1 U4377 ( .A1(n5917), .A2(n3504), .ZN(n3505) );
  NOR2_X1 U4378 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5768) );
  NOR2_X1 U4379 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3506) );
  INV_X1 U4380 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6692) );
  INV_X1 U4381 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5746) );
  NAND4_X1 U4382 ( .A1(n5768), .A2(n3506), .A3(n6692), .A4(n5746), .ZN(n3507)
         );
  OAI21_X1 U4383 ( .B1(n5592), .B2(n3507), .A(n5917), .ZN(n3509) );
  AND2_X1 U4384 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5767) );
  AND2_X1 U4385 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4213) );
  NAND2_X1 U4386 ( .A1(n5767), .A2(n4213), .ZN(n5738) );
  NAND2_X1 U4387 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4216) );
  NOR2_X1 U4388 ( .A1(n5738), .A2(n4216), .ZN(n4202) );
  NAND2_X1 U4389 ( .A1(n5592), .A2(n4202), .ZN(n3508) );
  XNOR2_X1 U4390 ( .A(n3493), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5582)
         );
  INV_X1 U4391 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3511) );
  AND2_X1 U4392 ( .A1(n3493), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5575)
         );
  NAND2_X1 U4393 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4221) );
  NOR2_X2 U4394 ( .A1(n5566), .A2(n4221), .ZN(n5545) );
  INV_X1 U4395 ( .A(n5545), .ZN(n3512) );
  INV_X1 U4396 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U4397 ( .A1(n5917), .A2(n5557), .ZN(n5574) );
  NOR3_X1 U4398 ( .A1(n5574), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4042) );
  NAND2_X1 U4399 ( .A1(n3020), .A2(n4042), .ZN(n5547) );
  NAND2_X1 U4400 ( .A1(n3512), .A2(n5547), .ZN(n3513) );
  XNOR2_X1 U4401 ( .A(n3513), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5685)
         );
  XNOR2_X1 U4402 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3526) );
  NAND2_X1 U4403 ( .A1(n3526), .A2(n3525), .ZN(n3524) );
  NAND2_X1 U4404 ( .A1(n4704), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U4405 ( .A1(n3524), .A2(n3514), .ZN(n3540) );
  XNOR2_X1 U4406 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3538) );
  NAND2_X1 U4407 ( .A1(n3540), .A2(n3538), .ZN(n3516) );
  NAND2_X1 U4408 ( .A1(n6478), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3515) );
  NAND2_X1 U4409 ( .A1(n3516), .A2(n3515), .ZN(n3522) );
  XNOR2_X1 U4410 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4411 ( .A1(n3522), .A2(n3520), .ZN(n3518) );
  NAND2_X1 U4412 ( .A1(n6768), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U4413 ( .A1(n3518), .A2(n3517), .ZN(n3556) );
  INV_X1 U4414 ( .A(n3520), .ZN(n3521) );
  XNOR2_X1 U4415 ( .A(n3522), .B(n3521), .ZN(n4058) );
  OAI21_X1 U4416 ( .B1(n3526), .B2(n3525), .A(n3524), .ZN(n3536) );
  INV_X1 U4417 ( .A(n3536), .ZN(n4056) );
  XNOR2_X1 U4418 ( .A(n3034), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3529)
         );
  NOR2_X1 U4419 ( .A1(n3527), .A2(n3529), .ZN(n3531) );
  AND2_X1 U4420 ( .A1(n3523), .A2(n3155), .ZN(n3528) );
  OAI21_X1 U4421 ( .B1(n3203), .B2(n3529), .A(n4874), .ZN(n3530) );
  NAND2_X1 U4422 ( .A1(n3547), .A2(n3530), .ZN(n3532) );
  OAI211_X1 U4423 ( .C1(n3535), .C2(n4056), .A(n3531), .B(n3532), .ZN(n3534)
         );
  INV_X1 U4424 ( .A(n3532), .ZN(n3533) );
  AOI22_X1 U4425 ( .A1(n3563), .A2(n3534), .B1(n3533), .B2(n4056), .ZN(n3546)
         );
  INV_X1 U4426 ( .A(n3535), .ZN(n3537) );
  NOR3_X1 U4427 ( .A1(n3537), .A2(n6669), .A3(n3536), .ZN(n3545) );
  INV_X1 U4428 ( .A(n3538), .ZN(n3539) );
  XNOR2_X1 U4429 ( .A(n3540), .B(n3539), .ZN(n4057) );
  NAND2_X1 U4430 ( .A1(n3559), .A2(n4057), .ZN(n3542) );
  INV_X1 U4431 ( .A(n4058), .ZN(n3541) );
  AOI21_X1 U4432 ( .B1(n3547), .B2(n3542), .A(n3541), .ZN(n3549) );
  NOR2_X1 U4433 ( .A1(n3543), .A2(n4057), .ZN(n3544) );
  OAI22_X1 U4434 ( .A1(n3546), .A2(n3545), .B1(n3549), .B2(n3544), .ZN(n3551)
         );
  INV_X1 U4435 ( .A(n3547), .ZN(n3548) );
  NAND4_X1 U4436 ( .A1(n3549), .A2(n4057), .A3(n3559), .A4(n3548), .ZN(n3550)
         );
  OAI211_X1 U4437 ( .C1(n4058), .C2(n3563), .A(n3551), .B(n3550), .ZN(n3552)
         );
  OAI21_X1 U4438 ( .B1(n2981), .B2(n4061), .A(n3552), .ZN(n3553) );
  AND2_X1 U4439 ( .A1(n6365), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3555)
         );
  INV_X1 U4440 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U4441 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5980), .ZN(n3557) );
  NAND2_X1 U4442 ( .A1(n4060), .A2(n3559), .ZN(n3560) );
  INV_X1 U4443 ( .A(n4060), .ZN(n3562) );
  NAND2_X1 U4444 ( .A1(n4645), .A2(n4315), .ZN(n3568) );
  OR2_X1 U4445 ( .A1(n4642), .A2(n3568), .ZN(n5334) );
  AND2_X1 U4446 ( .A1(n5334), .A2(n3339), .ZN(n3569) );
  NOR2_X1 U4447 ( .A1(n3567), .A2(n3569), .ZN(n4072) );
  AND2_X1 U4448 ( .A1(n4072), .A2(n3203), .ZN(n4229) );
  INV_X2 U4449 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U4450 ( .A1(n5007), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3926) );
  NAND2_X1 U4451 ( .A1(n4259), .A2(n3732), .ZN(n3574) );
  NOR2_X1 U4452 ( .A1(n3239), .A2(n5007), .ZN(n3601) );
  NAND2_X1 U4453 ( .A1(n3601), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4454 ( .A1(n3593), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5007), .ZN(n3571) );
  AND2_X1 U4455 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  NAND2_X1 U4456 ( .A1(n3574), .A2(n3573), .ZN(n4376) );
  AOI21_X1 U4457 ( .B1(n4703), .B2(n3575), .A(n5007), .ZN(n4348) );
  NAND2_X1 U4458 ( .A1(n2985), .A2(n3732), .ZN(n3581) );
  INV_X1 U4459 ( .A(n3601), .ZN(n3597) );
  NAND2_X1 U4460 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5007), .ZN(n3578)
         );
  NAND2_X1 U4461 ( .A1(n3593), .A2(EAX_REG_0__SCAN_IN), .ZN(n3577) );
  OAI211_X1 U4462 ( .C1(n3597), .C2(n3034), .A(n3578), .B(n3577), .ZN(n3579)
         );
  INV_X1 U4463 ( .A(n3579), .ZN(n3580) );
  NAND2_X1 U4464 ( .A1(n3581), .A2(n3580), .ZN(n4347) );
  NAND2_X1 U4465 ( .A1(n4348), .A2(n4347), .ZN(n4350) );
  INV_X1 U4466 ( .A(n4347), .ZN(n3582) );
  NAND2_X1 U4467 ( .A1(n3582), .A2(n4028), .ZN(n3583) );
  NAND2_X1 U4468 ( .A1(n4350), .A2(n3583), .ZN(n4375) );
  INV_X1 U4469 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3586) );
  NAND2_X1 U4470 ( .A1(n3601), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3585) );
  OAI21_X1 U4471 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3591), .ZN(n6262) );
  AOI22_X1 U4472 ( .A1(n4028), .A2(n6262), .B1(n5350), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3584) );
  OAI211_X1 U4473 ( .C1(n3594), .C2(n3586), .A(n3585), .B(n3584), .ZN(n4435)
         );
  NAND2_X1 U4474 ( .A1(n4436), .A2(n4435), .ZN(n3589) );
  NAND2_X1 U4475 ( .A1(n3587), .A2(n4378), .ZN(n3588) );
  NAND2_X1 U4476 ( .A1(n4817), .A2(n3732), .ZN(n3600) );
  OAI21_X1 U4477 ( .B1(n3592), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3605), 
        .ZN(n6253) );
  AOI22_X1 U4478 ( .A1(n6253), .A2(n4028), .B1(n5350), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4479 ( .A1(n5351), .A2(EAX_REG_3__SCAN_IN), .ZN(n3595) );
  OAI211_X1 U4480 ( .C1(n3597), .C2(n3109), .A(n3596), .B(n3595), .ZN(n3598)
         );
  INV_X1 U4481 ( .A(n3598), .ZN(n3599) );
  NAND2_X1 U4482 ( .A1(n3600), .A2(n3599), .ZN(n4650) );
  NAND2_X1 U4483 ( .A1(n3601), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3607) );
  INV_X1 U4484 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5987) );
  OAI21_X1 U4485 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n5987), .A(n5007), 
        .ZN(n3602) );
  INV_X1 U4486 ( .A(n3602), .ZN(n3603) );
  AOI21_X1 U4487 ( .B1(n5351), .B2(EAX_REG_4__SCAN_IN), .A(n3603), .ZN(n3606)
         );
  AOI21_X1 U4488 ( .B1(n3605), .B2(n3604), .A(n3611), .ZN(n4952) );
  AOI22_X1 U4489 ( .A1(n3607), .A2(n3606), .B1(n4028), .B2(n4952), .ZN(n3608)
         );
  NAND2_X1 U4490 ( .A1(n3610), .A2(n3732), .ZN(n3617) );
  INV_X1 U4491 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3614) );
  NAND2_X1 U4492 ( .A1(n5350), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3613)
         );
  OAI21_X1 U4493 ( .B1(n3611), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3628), 
        .ZN(n6245) );
  NAND2_X1 U4494 ( .A1(n6245), .A2(n4028), .ZN(n3612) );
  OAI211_X1 U4495 ( .C1(n3594), .C2(n3614), .A(n3613), .B(n3612), .ZN(n3615)
         );
  INV_X1 U4496 ( .A(n3615), .ZN(n3616) );
  NAND2_X1 U4497 ( .A1(n3618), .A2(n3732), .ZN(n3624) );
  INV_X1 U4498 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3620) );
  OAI21_X1 U4499 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n5987), .A(n5007), 
        .ZN(n3619) );
  OAI21_X1 U4500 ( .B1(n3594), .B2(n3620), .A(n3619), .ZN(n3622) );
  XNOR2_X1 U4501 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3628), .ZN(n4919) );
  NAND2_X1 U4502 ( .A1(n4919), .A2(n4028), .ZN(n3621) );
  NAND2_X1 U4503 ( .A1(n3622), .A2(n3621), .ZN(n3623) );
  NAND2_X1 U4504 ( .A1(n3624), .A2(n3623), .ZN(n4605) );
  OAI21_X1 U4505 ( .B1(n3629), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3647), 
        .ZN(n6240) );
  NAND2_X1 U4506 ( .A1(n6240), .A2(n4028), .ZN(n3631) );
  AOI22_X1 U4507 ( .A1(n5351), .A2(EAX_REG_7__SCAN_IN), .B1(n5350), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3630) );
  AND2_X1 U4508 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  XNOR2_X1 U4509 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3647), .ZN(n4904) );
  AOI22_X1 U4510 ( .A1(n2994), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4511 ( .A1(n3000), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4512 ( .A1(n3308), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4513 ( .A1(n4014), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4514 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3643)
         );
  AOI22_X1 U4515 ( .A1(n2975), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n2995), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4516 ( .A1(n2991), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4517 ( .A1(n3403), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4518 ( .A1(n5285), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4519 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3642)
         );
  OR2_X1 U4520 ( .A1(n3643), .A2(n3642), .ZN(n3644) );
  AOI22_X1 U4521 ( .A1(n3732), .A2(n3644), .B1(n5350), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3646) );
  NAND2_X1 U4522 ( .A1(n5351), .A2(EAX_REG_8__SCAN_IN), .ZN(n3645) );
  OAI211_X1 U4523 ( .C1(n4904), .C2(n5279), .A(n3646), .B(n3645), .ZN(n4832)
         );
  XNOR2_X1 U4524 ( .A(n3664), .B(n3663), .ZN(n5110) );
  AOI22_X1 U4525 ( .A1(n4014), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4526 ( .A1(n3000), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4527 ( .A1(n2992), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4528 ( .A1(n5285), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3648) );
  NAND4_X1 U4529 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3657)
         );
  AOI22_X1 U4530 ( .A1(n2994), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4531 ( .A1(n3308), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4532 ( .A1(n2980), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4533 ( .A1(n3267), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3652) );
  NAND4_X1 U4534 ( .A1(n3655), .A2(n3654), .A3(n3653), .A4(n3652), .ZN(n3656)
         );
  NOR2_X1 U4535 ( .A1(n3657), .A2(n3656), .ZN(n3660) );
  NAND2_X1 U4536 ( .A1(n5351), .A2(EAX_REG_9__SCAN_IN), .ZN(n3659) );
  NAND2_X1 U4537 ( .A1(n5350), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3658)
         );
  OAI211_X1 U4538 ( .C1(n3847), .C2(n3660), .A(n3659), .B(n3658), .ZN(n3661)
         );
  AOI21_X1 U4539 ( .B1(n5110), .B2(n4864), .A(n3661), .ZN(n4931) );
  XOR2_X1 U4540 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3690), .Z(n6044) );
  INV_X1 U4541 ( .A(n6044), .ZN(n3679) );
  AOI22_X1 U4542 ( .A1(n2979), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4543 ( .A1(n2991), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4544 ( .A1(n5285), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4545 ( .A1(n3157), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3665) );
  NAND4_X1 U4546 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(n3674)
         );
  AOI22_X1 U4547 ( .A1(n4014), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4548 ( .A1(n5282), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4549 ( .A1(n3000), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4550 ( .A1(n3267), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4551 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3673)
         );
  NOR2_X1 U4552 ( .A1(n3674), .A2(n3673), .ZN(n3677) );
  NAND2_X1 U4553 ( .A1(n5351), .A2(EAX_REG_10__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4554 ( .A1(n5350), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3675)
         );
  OAI211_X1 U4555 ( .C1(n3847), .C2(n3677), .A(n3676), .B(n3675), .ZN(n3678)
         );
  AOI21_X1 U4556 ( .B1(n3679), .B2(n4864), .A(n3678), .ZN(n5218) );
  AOI22_X1 U4557 ( .A1(n2975), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4558 ( .A1(n2994), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4559 ( .A1(n4014), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4560 ( .A1(n5285), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3680) );
  NAND4_X1 U4561 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), .ZN(n3689)
         );
  AOI22_X1 U4562 ( .A1(n2991), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4563 ( .A1(n3308), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4564 ( .A1(n3260), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5284), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4565 ( .A1(n2995), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4566 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3688)
         );
  NOR2_X1 U4567 ( .A1(n3689), .A2(n3688), .ZN(n3693) );
  XNOR2_X1 U4568 ( .A(n3694), .B(n5195), .ZN(n5213) );
  NAND2_X1 U4569 ( .A1(n5213), .A2(n4028), .ZN(n3692) );
  AOI22_X1 U4570 ( .A1(n5351), .A2(EAX_REG_11__SCAN_IN), .B1(n5350), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3691) );
  OAI211_X1 U4571 ( .C1(n3693), .C2(n3847), .A(n3692), .B(n3691), .ZN(n5183)
         );
  NAND2_X1 U4572 ( .A1(n5184), .A2(n5183), .ZN(n5185) );
  INV_X1 U4573 ( .A(n5185), .ZN(n3712) );
  XOR2_X1 U4574 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3713), .Z(n6038) );
  NAND2_X1 U4575 ( .A1(n6038), .A2(n4028), .ZN(n3710) );
  INV_X1 U4576 ( .A(EAX_REG_12__SCAN_IN), .ZN(n3696) );
  OAI21_X1 U4577 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5987), .A(n5007), 
        .ZN(n3695) );
  OAI21_X1 U4578 ( .B1(n3594), .B2(n3696), .A(n3695), .ZN(n3709) );
  AOI22_X1 U4579 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n2994), .B1(n3873), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4580 ( .A1(n2974), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4581 ( .A1(n2991), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4582 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n5282), .B1(n2984), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3697) );
  NAND4_X1 U4583 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3706)
         );
  AOI22_X1 U4584 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4014), .B1(n3403), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4585 ( .A1(n3000), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4586 ( .A1(n3267), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4587 ( .A1(n3308), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3701) );
  NAND4_X1 U4588 ( .A1(n3704), .A2(n3703), .A3(n3702), .A4(n3701), .ZN(n3705)
         );
  NOR2_X1 U4589 ( .A1(n3706), .A2(n3705), .ZN(n3707) );
  NOR2_X1 U4590 ( .A1(n3847), .A2(n3707), .ZN(n3708) );
  AOI21_X1 U4591 ( .B1(n3710), .B2(n3709), .A(n3708), .ZN(n5227) );
  INV_X1 U4592 ( .A(n5227), .ZN(n3711) );
  INV_X1 U4593 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3717) );
  NAND2_X1 U4594 ( .A1(n3714), .A2(n3717), .ZN(n3716) );
  INV_X1 U4595 ( .A(n3843), .ZN(n3715) );
  NAND2_X1 U4596 ( .A1(n3716), .A2(n3715), .ZN(n6024) );
  NAND2_X1 U4597 ( .A1(n6024), .A2(n4028), .ZN(n3720) );
  NOR2_X1 U4598 ( .A1(n3926), .A2(n3717), .ZN(n3718) );
  AOI21_X1 U4599 ( .B1(n5351), .B2(EAX_REG_13__SCAN_IN), .A(n3718), .ZN(n3719)
         );
  NAND2_X1 U4600 ( .A1(n3720), .A2(n3719), .ZN(n3733) );
  AOI22_X1 U4601 ( .A1(n2994), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4602 ( .A1(n3380), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4603 ( .A1(n4014), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4604 ( .A1(n3403), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3721) );
  NAND4_X1 U4605 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3730)
         );
  AOI22_X1 U4606 ( .A1(n3308), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4607 ( .A1(n5285), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4608 ( .A1(n2975), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4609 ( .A1(n3267), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3725) );
  NAND4_X1 U4610 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3729)
         );
  OR2_X1 U4611 ( .A1(n3730), .A2(n3729), .ZN(n3731) );
  AND2_X1 U4612 ( .A1(n3732), .A2(n3731), .ZN(n5250) );
  INV_X1 U4613 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3734) );
  INV_X1 U4614 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5451) );
  OAI21_X1 U4615 ( .B1(n3751), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n3853), 
        .ZN(n5629) );
  OR2_X1 U4616 ( .A1(n5629), .A2(n5279), .ZN(n3750) );
  AOI22_X1 U4617 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n2994), .B1(n3873), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4618 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4014), .B1(n3403), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4619 ( .A1(n3992), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4620 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5282), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3735) );
  NAND4_X1 U4621 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(n3746)
         );
  AOI22_X1 U4622 ( .A1(n2975), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4623 ( .A1(n2995), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4624 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3308), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3742) );
  AOI21_X1 U4625 ( .B1(n2989), .B2(INSTQUEUE_REG_9__4__SCAN_IN), .A(n4864), 
        .ZN(n3740) );
  NAND2_X1 U4626 ( .A1(n2983), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3739)
         );
  AND2_X1 U4627 ( .A1(n3740), .A2(n3739), .ZN(n3741) );
  NAND4_X1 U4628 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3745)
         );
  INV_X1 U4629 ( .A(n5334), .ZN(n6467) );
  NAND2_X1 U4630 ( .A1(n6467), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U4631 ( .A1(n4023), .A2(n5279), .ZN(n3880) );
  OAI21_X1 U4632 ( .B1(n3746), .B2(n3745), .A(n3880), .ZN(n3748) );
  AOI22_X1 U4633 ( .A1(n5351), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5007), .ZN(n3747) );
  NAND2_X1 U4634 ( .A1(n3748), .A2(n3747), .ZN(n3749) );
  NAND2_X1 U4635 ( .A1(n3750), .A2(n3749), .ZN(n5427) );
  INV_X1 U4636 ( .A(n5427), .ZN(n3851) );
  INV_X1 U4637 ( .A(n3751), .ZN(n3754) );
  OR2_X1 U4638 ( .A1(n3752), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3753)
         );
  NAND2_X1 U4639 ( .A1(n3754), .A2(n3753), .ZN(n5916) );
  AOI22_X1 U4640 ( .A1(n2995), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4641 ( .A1(n4014), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4642 ( .A1(n5285), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4643 ( .A1(n2994), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3755) );
  NAND4_X1 U4644 ( .A1(n3758), .A2(n3757), .A3(n3756), .A4(n3755), .ZN(n3764)
         );
  AOI22_X1 U4645 ( .A1(n3873), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4646 ( .A1(n3308), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4647 ( .A1(n3380), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4648 ( .A1(n2979), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3759) );
  NAND4_X1 U4649 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(n3763)
         );
  NOR2_X1 U4650 ( .A1(n3764), .A2(n3763), .ZN(n3767) );
  OAI21_X1 U4651 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5987), .A(n5007), 
        .ZN(n3766) );
  NAND2_X1 U4652 ( .A1(n5351), .A2(EAX_REG_19__SCAN_IN), .ZN(n3765) );
  OAI211_X1 U4653 ( .C1(n4023), .C2(n3767), .A(n3766), .B(n3765), .ZN(n3768)
         );
  OAI21_X1 U4654 ( .B1(n5916), .B2(n5279), .A(n3768), .ZN(n5861) );
  INV_X1 U4655 ( .A(n5861), .ZN(n3850) );
  AOI22_X1 U4656 ( .A1(n3267), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4657 ( .A1(n3308), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4658 ( .A1(n4014), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4659 ( .A1(n2980), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3769) );
  NAND4_X1 U4660 ( .A1(n3772), .A2(n3771), .A3(n3770), .A4(n3769), .ZN(n3780)
         );
  AOI22_X1 U4661 ( .A1(n2991), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4662 ( .A1(n5282), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4663 ( .A1(n3873), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3776) );
  NAND2_X1 U4664 ( .A1(n2994), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3774)
         );
  AOI21_X1 U4665 ( .B1(n2987), .B2(INSTQUEUE_REG_9__2__SCAN_IN), .A(n4864), 
        .ZN(n3773) );
  AND2_X1 U4666 ( .A1(n3774), .A2(n3773), .ZN(n3775) );
  NAND4_X1 U4667 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3779)
         );
  OAI21_X1 U4668 ( .B1(n3780), .B2(n3779), .A(n3880), .ZN(n3782) );
  AOI22_X1 U4669 ( .A1(n5351), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5007), .ZN(n3781) );
  NAND2_X1 U4670 ( .A1(n3782), .A2(n3781), .ZN(n3784) );
  XNOR2_X1 U4671 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3799), .ZN(n5637)
         );
  NAND2_X1 U4672 ( .A1(n4864), .A2(n5637), .ZN(n3783) );
  NAND2_X1 U4673 ( .A1(n3784), .A2(n3783), .ZN(n5442) );
  INV_X1 U4674 ( .A(n5442), .ZN(n3849) );
  AOI22_X1 U4675 ( .A1(n3308), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4676 ( .A1(n3380), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4677 ( .A1(n3267), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4678 ( .A1(n4014), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4679 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3794)
         );
  AOI22_X1 U4680 ( .A1(n2994), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4681 ( .A1(n2980), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4682 ( .A1(n3403), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4683 ( .A1(n5285), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4684 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3793)
         );
  NOR2_X1 U4685 ( .A1(n3794), .A2(n3793), .ZN(n3798) );
  OAI21_X1 U4686 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n5987), .A(n5007), 
        .ZN(n3795) );
  INV_X1 U4687 ( .A(n3795), .ZN(n3796) );
  AOI21_X1 U4688 ( .B1(n5351), .B2(EAX_REG_17__SCAN_IN), .A(n3796), .ZN(n3797)
         );
  OAI21_X1 U4689 ( .B1(n4023), .B2(n3798), .A(n3797), .ZN(n3802) );
  OAI21_X1 U4690 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3800), .A(n3799), 
        .ZN(n6014) );
  OR2_X1 U4691 ( .A1(n5279), .A2(n6014), .ZN(n3801) );
  AND2_X1 U4692 ( .A1(n3802), .A2(n3801), .ZN(n5506) );
  XNOR2_X1 U4693 ( .A(n3803), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5462)
         );
  AOI22_X1 U4694 ( .A1(n3308), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4695 ( .A1(n4014), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n2994), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4696 ( .A1(n3380), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4697 ( .A1(n2984), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4698 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3813)
         );
  AOI22_X1 U4699 ( .A1(n2995), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4700 ( .A1(n2974), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4701 ( .A1(n3873), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4702 ( .A1(n5285), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4703 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812)
         );
  NOR2_X1 U4704 ( .A1(n3813), .A2(n3812), .ZN(n3816) );
  INV_X1 U4705 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5645) );
  NOR2_X1 U4706 ( .A1(n3926), .A2(n5645), .ZN(n3814) );
  AOI21_X1 U4707 ( .B1(n5351), .B2(EAX_REG_16__SCAN_IN), .A(n3814), .ZN(n3815)
         );
  OAI21_X1 U4708 ( .B1(n4023), .B2(n3816), .A(n3815), .ZN(n3817) );
  AOI21_X1 U4709 ( .B1(n5462), .B2(n4864), .A(n3817), .ZN(n5456) );
  XNOR2_X1 U4710 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3818), .ZN(n6020)
         );
  INV_X1 U4711 ( .A(n6020), .ZN(n5656) );
  AOI22_X1 U4712 ( .A1(n2974), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4713 ( .A1(n2994), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4714 ( .A1(n2995), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4715 ( .A1(n5282), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4716 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3828)
         );
  AOI22_X1 U4717 ( .A1(n3873), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4718 ( .A1(n4014), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4719 ( .A1(n5285), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4720 ( .A1(n3308), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4721 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3827)
         );
  NOR2_X1 U4722 ( .A1(n3828), .A2(n3827), .ZN(n3831) );
  NAND2_X1 U4723 ( .A1(n5351), .A2(EAX_REG_15__SCAN_IN), .ZN(n3830) );
  NAND2_X1 U4724 ( .A1(n5350), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3829)
         );
  OAI211_X1 U4725 ( .C1(n3847), .C2(n3831), .A(n3830), .B(n3829), .ZN(n3832)
         );
  AOI21_X1 U4726 ( .B1(n5656), .B2(n4864), .A(n3832), .ZN(n5537) );
  NOR2_X1 U4727 ( .A1(n5456), .A2(n5537), .ZN(n5459) );
  AND2_X1 U4728 ( .A1(n5506), .A2(n5459), .ZN(n3848) );
  AOI22_X1 U4729 ( .A1(n3308), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4730 ( .A1(n3265), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4731 ( .A1(n3873), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4732 ( .A1(n2995), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3833) );
  NAND4_X1 U4733 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(n3842)
         );
  AOI22_X1 U4734 ( .A1(n5282), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4735 ( .A1(n4014), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4736 ( .A1(n2994), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4737 ( .A1(n2979), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3837) );
  NAND4_X1 U4738 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3841)
         );
  NOR2_X1 U4739 ( .A1(n3842), .A2(n3841), .ZN(n3846) );
  XNOR2_X1 U4740 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3843), .ZN(n5663)
         );
  AOI22_X1 U4741 ( .A1(n4864), .A2(n5663), .B1(n5350), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3845) );
  NAND2_X1 U4742 ( .A1(n5351), .A2(EAX_REG_14__SCAN_IN), .ZN(n3844) );
  OAI211_X1 U4743 ( .C1(n3847), .C2(n3846), .A(n3845), .B(n3844), .ZN(n5457)
         );
  AND2_X1 U4744 ( .A1(n3848), .A2(n5457), .ZN(n5439) );
  INV_X1 U4745 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5622) );
  AND2_X1 U4746 ( .A1(n3853), .A2(n5622), .ZN(n3854) );
  OR2_X1 U4747 ( .A1(n3854), .A2(n3885), .ZN(n5422) );
  INV_X1 U4748 ( .A(n5422), .ZN(n5625) );
  INV_X1 U4749 ( .A(n4023), .ZN(n5298) );
  AOI22_X1 U4750 ( .A1(n3265), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4751 ( .A1(n4014), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4752 ( .A1(n2980), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4753 ( .A1(n2994), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3855) );
  NAND4_X1 U4754 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n3864)
         );
  AOI22_X1 U4755 ( .A1(n3873), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4756 ( .A1(n3308), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4757 ( .A1(n5285), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4758 ( .A1(n2995), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3859) );
  NAND4_X1 U4759 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3863)
         );
  OR2_X1 U4760 ( .A1(n3864), .A2(n3863), .ZN(n3867) );
  NAND2_X1 U4761 ( .A1(n5351), .A2(EAX_REG_21__SCAN_IN), .ZN(n3865) );
  OAI211_X1 U4762 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n5622), .A(n3865), .B(
        n5279), .ZN(n3866) );
  AOI21_X1 U4763 ( .B1(n5298), .B2(n3867), .A(n3866), .ZN(n3868) );
  AOI21_X1 U4764 ( .B1(n5625), .B2(n4864), .A(n3868), .ZN(n5415) );
  AND2_X2 U4765 ( .A1(n5414), .A2(n5415), .ZN(n5494) );
  INV_X1 U4766 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5616) );
  XNOR2_X1 U4767 ( .A(n3885), .B(n5616), .ZN(n5845) );
  AOI22_X1 U4768 ( .A1(n5351), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5007), .ZN(n3884) );
  AOI22_X1 U4769 ( .A1(n2974), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4770 ( .A1(n5283), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3296), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4771 ( .A1(n2994), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4772 ( .A1(n3267), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5284), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4773 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3882)
         );
  AOI22_X1 U4774 ( .A1(n3000), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4775 ( .A1(n3992), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4776 ( .A1(n5282), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3877) );
  NAND2_X1 U4777 ( .A1(n3873), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3875)
         );
  AOI21_X1 U4778 ( .B1(n2989), .B2(INSTQUEUE_REG_9__6__SCAN_IN), .A(n4864), 
        .ZN(n3874) );
  AND2_X1 U4779 ( .A1(n3875), .A2(n3874), .ZN(n3876) );
  NAND4_X1 U4780 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3881)
         );
  OAI21_X1 U4781 ( .B1(n3882), .B2(n3881), .A(n3880), .ZN(n3883) );
  AOI22_X1 U4782 ( .A1(n5845), .A2(n4028), .B1(n3884), .B2(n3883), .ZN(n5493)
         );
  AND2_X2 U4783 ( .A1(n5494), .A2(n5493), .ZN(n5604) );
  INV_X1 U4784 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3908) );
  NAND2_X1 U4785 ( .A1(n3886), .A2(n3908), .ZN(n3887) );
  NAND2_X1 U4786 ( .A1(n3932), .A2(n3887), .ZN(n5841) );
  AOI22_X1 U4787 ( .A1(n4014), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4788 ( .A1(n2994), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4789 ( .A1(n2975), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4790 ( .A1(n5285), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3888) );
  NAND4_X1 U4791 ( .A1(n3891), .A2(n3890), .A3(n3889), .A4(n3888), .ZN(n3897)
         );
  AOI22_X1 U4792 ( .A1(n3308), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4793 ( .A1(n3873), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4794 ( .A1(n3267), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4795 ( .A1(n3380), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3892) );
  NAND4_X1 U4796 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3896)
         );
  NOR2_X1 U4797 ( .A1(n3897), .A2(n3896), .ZN(n3914) );
  AOI22_X1 U4798 ( .A1(n3308), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4799 ( .A1(n2994), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4800 ( .A1(n2975), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4801 ( .A1(n2995), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3898) );
  NAND4_X1 U4802 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3907)
         );
  AOI22_X1 U4803 ( .A1(n3000), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4804 ( .A1(n4014), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3260), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4805 ( .A1(n3873), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4806 ( .A1(n5285), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4807 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3906)
         );
  NOR2_X1 U4808 ( .A1(n3907), .A2(n3906), .ZN(n3915) );
  XNOR2_X1 U4809 ( .A(n3914), .B(n3915), .ZN(n3911) );
  OAI21_X1 U4810 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3908), .A(n5279), .ZN(
        n3909) );
  AOI21_X1 U4811 ( .B1(n5351), .B2(EAX_REG_23__SCAN_IN), .A(n3909), .ZN(n3910)
         );
  OAI21_X1 U4812 ( .B1(n4023), .B2(n3911), .A(n3910), .ZN(n3912) );
  INV_X1 U4813 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5406) );
  XNOR2_X1 U4814 ( .A(n3932), .B(n5406), .ZN(n5599) );
  NOR2_X1 U4815 ( .A1(n3915), .A2(n3914), .ZN(n3946) );
  AOI22_X1 U4816 ( .A1(n2994), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4817 ( .A1(n3380), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4818 ( .A1(n4014), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4819 ( .A1(n3403), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5284), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3916) );
  NAND4_X1 U4820 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3925)
         );
  AOI22_X1 U4821 ( .A1(n3308), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4822 ( .A1(n5285), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4823 ( .A1(n2974), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4824 ( .A1(n3267), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3920) );
  NAND4_X1 U4825 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3920), .ZN(n3924)
         );
  OR2_X1 U4826 ( .A1(n3925), .A2(n3924), .ZN(n3945) );
  XNOR2_X1 U4827 ( .A(n3946), .B(n3945), .ZN(n3929) );
  NOR2_X1 U4828 ( .A1(n3926), .A2(n5406), .ZN(n3927) );
  AOI21_X1 U4829 ( .B1(n5351), .B2(EAX_REG_24__SCAN_IN), .A(n3927), .ZN(n3928)
         );
  OAI21_X1 U4830 ( .B1(n3929), .B2(n4023), .A(n3928), .ZN(n3930) );
  AOI21_X1 U4831 ( .B1(n5599), .B2(n4028), .A(n3930), .ZN(n5404) );
  INV_X1 U4832 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5827) );
  AND2_X1 U4833 ( .A1(n3933), .A2(n5827), .ZN(n3934) );
  OR2_X1 U4834 ( .A1(n3934), .A2(n3969), .ZN(n5824) );
  AOI22_X1 U4835 ( .A1(n3308), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4836 ( .A1(n5282), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4837 ( .A1(n5285), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4838 ( .A1(n2994), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5284), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3935) );
  NAND4_X1 U4839 ( .A1(n3938), .A2(n3937), .A3(n3936), .A4(n3935), .ZN(n3944)
         );
  AOI22_X1 U4840 ( .A1(n4014), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4841 ( .A1(n2974), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4842 ( .A1(n3000), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4843 ( .A1(n2995), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3939) );
  NAND4_X1 U4844 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3943)
         );
  NOR2_X1 U4845 ( .A1(n3944), .A2(n3943), .ZN(n3952) );
  NAND2_X1 U4846 ( .A1(n3946), .A2(n3945), .ZN(n3951) );
  XNOR2_X1 U4847 ( .A(n3952), .B(n3951), .ZN(n3949) );
  AOI21_X1 U4848 ( .B1(n5827), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3947) );
  AOI21_X1 U4849 ( .B1(n5351), .B2(EAX_REG_25__SCAN_IN), .A(n3947), .ZN(n3948)
         );
  OAI21_X1 U4850 ( .B1(n3949), .B2(n4023), .A(n3948), .ZN(n3950) );
  OAI21_X1 U4851 ( .B1(n5824), .B2(n5279), .A(n3950), .ZN(n5585) );
  INV_X1 U4852 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5578) );
  XNOR2_X1 U4853 ( .A(n3969), .B(n5578), .ZN(n5814) );
  OR2_X1 U4854 ( .A1(n3952), .A2(n3951), .ZN(n3971) );
  AOI22_X1 U4855 ( .A1(n2994), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4856 ( .A1(n5282), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4857 ( .A1(n4014), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4858 ( .A1(n5285), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n2970), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4859 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3962)
         );
  AOI22_X1 U4860 ( .A1(n3308), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4861 ( .A1(n3380), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4862 ( .A1(n2974), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4863 ( .A1(n3267), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3957) );
  NAND4_X1 U4864 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n3961)
         );
  NOR2_X1 U4865 ( .A1(n3962), .A2(n3961), .ZN(n3972) );
  XOR2_X1 U4866 ( .A(n3971), .B(n3972), .Z(n3966) );
  INV_X1 U4867 ( .A(EAX_REG_26__SCAN_IN), .ZN(n3964) );
  NAND2_X1 U4868 ( .A1(n5007), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3963)
         );
  OAI211_X1 U4869 ( .C1(n3594), .C2(n3964), .A(n5279), .B(n3963), .ZN(n3965)
         );
  AOI21_X1 U4870 ( .B1(n3966), .B2(n5298), .A(n3965), .ZN(n3967) );
  AOI21_X1 U4871 ( .B1(n5814), .B2(n4028), .A(n3967), .ZN(n5485) );
  AND2_X2 U4872 ( .A1(n5588), .A2(n5485), .ZN(n5569) );
  AND2_X1 U4873 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3968) );
  AOI21_X1 U4874 ( .B1(n3969), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3970) );
  OR2_X1 U4875 ( .A1(n3988), .A2(n3970), .ZN(n5813) );
  OR2_X1 U4876 ( .A1(n3972), .A2(n3971), .ZN(n3990) );
  AOI22_X1 U4877 ( .A1(n3308), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4878 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n2994), .B1(n3403), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4879 ( .A1(n5285), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n2989), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4880 ( .A1(n3267), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3973) );
  NAND4_X1 U4881 ( .A1(n3976), .A2(n3975), .A3(n3974), .A4(n3973), .ZN(n3982)
         );
  AOI22_X1 U4882 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3000), .B1(n5282), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4883 ( .A1(n2975), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4884 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4014), .B1(n3260), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4885 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3873), .B1(n5284), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3977) );
  NAND4_X1 U4886 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n3977), .ZN(n3981)
         );
  NOR2_X1 U4887 ( .A1(n3982), .A2(n3981), .ZN(n3991) );
  XNOR2_X1 U4888 ( .A(n3990), .B(n3991), .ZN(n3985) );
  INV_X1 U4889 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5807) );
  AOI21_X1 U4890 ( .B1(n5807), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3983) );
  AOI21_X1 U4891 ( .B1(n5351), .B2(EAX_REG_27__SCAN_IN), .A(n3983), .ZN(n3984)
         );
  OAI21_X1 U4892 ( .B1(n3985), .B2(n4023), .A(n3984), .ZN(n3986) );
  OAI21_X1 U4893 ( .B1(n5813), .B2(n5279), .A(n3986), .ZN(n3987) );
  INV_X1 U4894 ( .A(n3987), .ZN(n5568) );
  OR2_X1 U4895 ( .A1(n3988), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3989)
         );
  NAND2_X1 U4896 ( .A1(n4008), .A2(n3989), .ZN(n5561) );
  INV_X1 U4897 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4006) );
  NOR2_X1 U4898 ( .A1(n3991), .A2(n3990), .ZN(n4022) );
  AOI22_X1 U4899 ( .A1(n3308), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2992), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4900 ( .A1(n4014), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4901 ( .A1(n3992), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4902 ( .A1(n3403), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U4903 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4002)
         );
  AOI22_X1 U4904 ( .A1(n2994), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4905 ( .A1(n2974), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4906 ( .A1(n5285), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4907 ( .A1(n3000), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U4908 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4001)
         );
  OR2_X1 U4909 ( .A1(n4002), .A2(n4001), .ZN(n4021) );
  XOR2_X1 U4910 ( .A(n4022), .B(n4021), .Z(n4003) );
  NAND2_X1 U4911 ( .A1(n4003), .A2(n5298), .ZN(n4005) );
  OAI21_X1 U4912 ( .B1(n5987), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5007), 
        .ZN(n4004) );
  OAI211_X1 U4913 ( .C1(n3594), .C2(n4006), .A(n4005), .B(n4004), .ZN(n4007)
         );
  OAI21_X1 U4914 ( .B1(n5561), .B2(n5279), .A(n4007), .ZN(n5392) );
  INV_X1 U4915 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U4916 ( .A1(n4008), .A2(n4035), .ZN(n4009) );
  AOI21_X1 U4917 ( .B1(n4035), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4918 ( .A1(n3296), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4919 ( .A1(n3380), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4920 ( .A1(n3403), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n2983), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4921 ( .A1(n2970), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n2988), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4922 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4020)
         );
  AOI22_X1 U4923 ( .A1(n2979), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5285), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4924 ( .A1(n2995), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n2991), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4925 ( .A1(n2994), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3873), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4926 ( .A1(n4014), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4015) );
  NAND4_X1 U4927 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4019)
         );
  NOR2_X1 U4928 ( .A1(n4020), .A2(n4019), .ZN(n5281) );
  NAND2_X1 U4929 ( .A1(n4022), .A2(n4021), .ZN(n5280) );
  XNOR2_X1 U4930 ( .A(n5281), .B(n5280), .ZN(n4024) );
  NOR2_X1 U4931 ( .A1(n4024), .A2(n4023), .ZN(n4025) );
  AOI211_X1 U4932 ( .C1(n5351), .C2(EAX_REG_29__SCAN_IN), .A(n4026), .B(n4025), 
        .ZN(n4027) );
  AOI21_X1 U4933 ( .B1(n5382), .B2(n4028), .A(n4027), .ZN(n4030) );
  AND2_X1 U4934 ( .A1(n6669), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U4935 ( .A1(n4865), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6509) );
  NOR2_X1 U4936 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n4807) );
  NOR2_X1 U4937 ( .A1(n5380), .A2(n6271), .ZN(n4040) );
  AOI21_X1 U4938 ( .B1(n5799), .B2(n4034), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n4031) );
  NAND2_X1 U4939 ( .A1(n6669), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4033) );
  NAND2_X1 U4940 ( .A1(n5987), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4032) );
  NAND2_X1 U4941 ( .A1(n4033), .A2(n4032), .ZN(n6275) );
  NAND2_X1 U4942 ( .A1(n5649), .A2(n5382), .ZN(n4038) );
  OR2_X1 U4943 ( .A1(n4034), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U4944 ( .A1(n6338), .A2(REIP_REG_29__SCAN_IN), .ZN(n5677) );
  OAI21_X1 U4945 ( .B1(n5646), .B2(n4035), .A(n5677), .ZN(n4036) );
  INV_X1 U4946 ( .A(n4036), .ZN(n4037) );
  OAI21_X1 U4947 ( .B1(n5685), .B2(n6273), .A(n4041), .ZN(U2957) );
  NAND2_X1 U4948 ( .A1(n5545), .A2(n3106), .ZN(n4044) );
  INV_X1 U4949 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5668) );
  INV_X1 U4950 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5682) );
  NAND3_X1 U4951 ( .A1(n4042), .A2(n5668), .A3(n5682), .ZN(n4043) );
  NAND2_X1 U4952 ( .A1(n4044), .A2(n3102), .ZN(n4046) );
  XNOR2_X1 U4953 ( .A(n4046), .B(n4045), .ZN(n5368) );
  NOR2_X1 U4954 ( .A1(n5334), .A2(n3523), .ZN(n4197) );
  INV_X1 U4955 ( .A(n4197), .ZN(n4065) );
  NOR2_X1 U4956 ( .A1(n4048), .A2(n4047), .ZN(n4234) );
  INV_X1 U4957 ( .A(n4234), .ZN(n4053) );
  NAND2_X1 U4958 ( .A1(n4049), .A2(n4874), .ZN(n4051) );
  MUX2_X1 U4959 ( .A(n4051), .B(n6616), .S(n4050), .Z(n4194) );
  NAND2_X1 U4960 ( .A1(n4194), .A2(n4072), .ZN(n4052) );
  NAND2_X1 U4961 ( .A1(n4053), .A2(n4052), .ZN(n4474) );
  INV_X1 U4962 ( .A(n4054), .ZN(n4055) );
  INV_X1 U4963 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U4964 ( .A1(n4055), .A2(n6519), .ZN(n6517) );
  NAND2_X1 U4965 ( .A1(n4323), .A2(n6517), .ZN(n4063) );
  AND3_X1 U4966 ( .A1(n4058), .A2(n4057), .A3(n4056), .ZN(n4059) );
  OR2_X1 U4967 ( .A1(n4060), .A2(n4059), .ZN(n4062) );
  NAND2_X1 U4968 ( .A1(n4062), .A2(n4061), .ZN(n4228) );
  INV_X1 U4969 ( .A(n4228), .ZN(n4233) );
  NOR2_X1 U4970 ( .A1(n4233), .A2(READY_N), .ZN(n4481) );
  NAND3_X1 U4971 ( .A1(n4063), .A2(n4481), .A3(n3210), .ZN(n4064) );
  OAI211_X1 U4972 ( .C1(n4480), .C2(n4065), .A(n4474), .B(n4064), .ZN(n4066)
         );
  NAND2_X1 U4973 ( .A1(n4066), .A2(n6490), .ZN(n4071) );
  INV_X1 U4974 ( .A(READY_N), .ZN(n6610) );
  NAND2_X1 U4975 ( .A1(n3523), .A2(n6517), .ZN(n4869) );
  NAND3_X1 U4976 ( .A1(n4494), .A2(n6610), .A3(n4869), .ZN(n4068) );
  AND2_X1 U4977 ( .A1(n3239), .A2(n4874), .ZN(n4067) );
  AOI21_X1 U4978 ( .B1(n4068), .B2(n4067), .A(n3210), .ZN(n4069) );
  NAND2_X1 U4979 ( .A1(n6149), .A2(n4069), .ZN(n4070) );
  INV_X1 U4980 ( .A(n4229), .ZN(n6484) );
  AND2_X1 U4981 ( .A1(n4072), .A2(n3237), .ZN(n4479) );
  INV_X1 U4982 ( .A(n4479), .ZN(n4498) );
  NAND2_X1 U4983 ( .A1(n4494), .A2(n4307), .ZN(n4639) );
  NAND2_X1 U4984 ( .A1(n4183), .A2(n4315), .ZN(n4073) );
  AND2_X1 U4985 ( .A1(n4639), .A2(n4073), .ZN(n4074) );
  NAND4_X1 U4986 ( .A1(n5976), .A2(n6484), .A3(n4498), .A4(n4074), .ZN(n4075)
         );
  NAND2_X1 U4987 ( .A1(n5368), .A2(n6354), .ZN(n4226) );
  CLKBUF_X3 U4988 ( .A(n4077), .Z(n5444) );
  INV_X2 U4989 ( .A(n4158), .ZN(n4174) );
  MUX2_X1 U4990 ( .A(n4174), .B(n5444), .S(EBX_REG_2__SCAN_IN), .Z(n4078) );
  OAI21_X1 U4991 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n4344), .A(n4078), 
        .ZN(n4432) );
  INV_X1 U4992 ( .A(n4432), .ZN(n4088) );
  INV_X1 U4993 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4079) );
  NAND2_X1 U4994 ( .A1(n4158), .A2(n4079), .ZN(n4082) );
  INV_X2 U4995 ( .A(n4307), .ZN(n4880) );
  NAND2_X1 U4996 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4080)
         );
  OAI211_X1 U4997 ( .C1(n4880), .C2(EBX_REG_1__SCAN_IN), .A(n4083), .B(n4080), 
        .ZN(n4081) );
  NAND2_X1 U4998 ( .A1(n4082), .A2(n4081), .ZN(n4085) );
  INV_X1 U4999 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4084) );
  OAI22_X1 U5000 ( .A1(n4083), .A2(n4084), .B1(n5444), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4345) );
  XNOR2_X1 U5001 ( .A(n4085), .B(n4345), .ZN(n4281) );
  NAND2_X1 U5002 ( .A1(n4281), .A2(n4307), .ZN(n4087) );
  INV_X1 U5003 ( .A(n4085), .ZN(n4086) );
  NAND2_X1 U5004 ( .A1(n4083), .A2(n6336), .ZN(n4090) );
  INV_X1 U5005 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6753) );
  NAND2_X1 U5006 ( .A1(n4307), .A2(n6753), .ZN(n4089) );
  NAND3_X1 U5007 ( .A1(n4090), .A2(n5444), .A3(n4089), .ZN(n4092) );
  NAND2_X1 U5008 ( .A1(n2977), .A2(n6753), .ZN(n4091) );
  INV_X1 U5009 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4950) );
  NAND2_X1 U5010 ( .A1(n4158), .A2(n4950), .ZN(n4095) );
  NAND2_X1 U5011 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4093)
         );
  OAI211_X1 U5012 ( .C1(n4880), .C2(EBX_REG_4__SCAN_IN), .A(n4083), .B(n4093), 
        .ZN(n4094) );
  NAND2_X1 U5013 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4096)
         );
  NAND2_X1 U5014 ( .A1(n4083), .A2(n4096), .ZN(n4098) );
  INV_X1 U5015 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4799) );
  NAND2_X1 U5016 ( .A1(n4307), .A2(n4799), .ZN(n4097) );
  NAND2_X1 U5017 ( .A1(n4098), .A2(n4097), .ZN(n4100) );
  NAND2_X1 U5018 ( .A1(n2977), .A2(n4799), .ZN(n4099) );
  NAND2_X1 U5019 ( .A1(n4100), .A2(n4099), .ZN(n4561) );
  NAND2_X1 U5020 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4101)
         );
  OAI211_X1 U5021 ( .C1(n4880), .C2(EBX_REG_6__SCAN_IN), .A(n4083), .B(n4101), 
        .ZN(n4102) );
  OAI21_X1 U5022 ( .B1(n4174), .B2(EBX_REG_6__SCAN_IN), .A(n4102), .ZN(n4607)
         );
  MUX2_X1 U5023 ( .A(n4174), .B(n5444), .S(EBX_REG_8__SCAN_IN), .Z(n4103) );
  OAI21_X1 U5024 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n4344), .A(n4103), 
        .ZN(n4891) );
  INV_X1 U5025 ( .A(n4891), .ZN(n4108) );
  NAND2_X1 U5026 ( .A1(n4083), .A2(n6305), .ZN(n4105) );
  INV_X1 U5027 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U5028 ( .A1(n4307), .A2(n6735), .ZN(n4104) );
  NAND3_X1 U5029 ( .A1(n4105), .A2(n5444), .A3(n4104), .ZN(n4107) );
  NAND2_X1 U5030 ( .A1(n2977), .A2(n6735), .ZN(n4106) );
  NAND2_X1 U5031 ( .A1(n4107), .A2(n4106), .ZN(n6051) );
  NAND2_X1 U5032 ( .A1(n4108), .A2(n6051), .ZN(n4109) );
  NAND2_X1 U5033 ( .A1(n4083), .A2(n5126), .ZN(n4111) );
  INV_X1 U5034 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U5035 ( .A1(n4307), .A2(n6671), .ZN(n4110) );
  NAND3_X1 U5036 ( .A1(n4111), .A2(n5444), .A3(n4110), .ZN(n4113) );
  NAND2_X1 U5037 ( .A1(n2977), .A2(n6671), .ZN(n4112) );
  AND2_X1 U5038 ( .A1(n4113), .A2(n4112), .ZN(n4935) );
  NAND2_X1 U5039 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4114) );
  OAI211_X1 U5040 ( .C1(n4880), .C2(EBX_REG_10__SCAN_IN), .A(n4083), .B(n4114), 
        .ZN(n4115) );
  OAI21_X1 U5041 ( .B1(n4174), .B2(EBX_REG_10__SCAN_IN), .A(n4115), .ZN(n5128)
         );
  NOR2_X1 U5042 ( .A1(n4935), .A2(n5128), .ZN(n4116) );
  NAND2_X1 U5043 ( .A1(n4083), .A2(n5209), .ZN(n4118) );
  INV_X1 U5044 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U5045 ( .A1(n4307), .A2(n5191), .ZN(n4117) );
  NAND3_X1 U5046 ( .A1(n4118), .A2(n5444), .A3(n4117), .ZN(n4120) );
  NAND2_X1 U5047 ( .A1(n2977), .A2(n5191), .ZN(n4119) );
  NAND2_X1 U5048 ( .A1(n4120), .A2(n4119), .ZN(n5188) );
  NAND2_X1 U5049 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4121) );
  OAI211_X1 U5050 ( .C1(n4880), .C2(EBX_REG_12__SCAN_IN), .A(n4083), .B(n4121), 
        .ZN(n4122) );
  OAI21_X1 U5051 ( .B1(n4174), .B2(EBX_REG_12__SCAN_IN), .A(n4122), .ZN(n5234)
         );
  NAND2_X1 U5052 ( .A1(n4083), .A2(n5974), .ZN(n4124) );
  INV_X1 U5053 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U5054 ( .A1(n4307), .A2(n6752), .ZN(n4123) );
  NAND3_X1 U5055 ( .A1(n4124), .A2(n5444), .A3(n4123), .ZN(n4126) );
  NAND2_X1 U5056 ( .A1(n2977), .A2(n6752), .ZN(n4125) );
  AND2_X1 U5057 ( .A1(n4126), .A2(n4125), .ZN(n5251) );
  MUX2_X1 U5058 ( .A(n4174), .B(n5444), .S(EBX_REG_14__SCAN_IN), .Z(n4127) );
  OAI21_X1 U5059 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n4344), .A(n4127), 
        .ZN(n4128) );
  INV_X1 U5060 ( .A(n4128), .ZN(n5265) );
  AND2_X2 U5061 ( .A1(n5266), .A2(n5265), .ZN(n5786) );
  MUX2_X1 U5062 ( .A(n4174), .B(n5444), .S(EBX_REG_16__SCAN_IN), .Z(n4130) );
  OR2_X1 U5063 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4129)
         );
  NAND2_X1 U5064 ( .A1(n4130), .A2(n4129), .ZN(n5464) );
  NAND2_X1 U5065 ( .A1(n4083), .A2(n5942), .ZN(n4132) );
  INV_X1 U5066 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U5067 ( .A1(n4307), .A2(n6107), .ZN(n4131) );
  NAND3_X1 U5068 ( .A1(n4132), .A2(n5444), .A3(n4131), .ZN(n4134) );
  NAND2_X1 U5069 ( .A1(n2977), .A2(n6107), .ZN(n4133) );
  AND2_X1 U5070 ( .A1(n4134), .A2(n4133), .ZN(n5785) );
  NOR2_X1 U5071 ( .A1(n5464), .A2(n5785), .ZN(n4135) );
  NAND2_X1 U5072 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4136) );
  NAND2_X1 U5073 ( .A1(n4083), .A2(n4136), .ZN(n4138) );
  INV_X1 U5074 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U5075 ( .A1(n4307), .A2(n5515), .ZN(n4137) );
  AOI22_X1 U5076 ( .A1(n4138), .A2(n4137), .B1(n2977), .B2(n5515), .ZN(n5510)
         );
  INV_X1 U5077 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U5078 ( .A1(n4158), .A2(n5889), .ZN(n4141) );
  NAND2_X1 U5079 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4139) );
  OAI211_X1 U5080 ( .C1(n4880), .C2(EBX_REG_19__SCAN_IN), .A(n4083), .B(n4139), 
        .ZN(n4140) );
  NAND2_X1 U5081 ( .A1(n4141), .A2(n4140), .ZN(n5867) );
  OR2_X1 U5082 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4143)
         );
  INV_X1 U5083 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U5084 ( .A1(n4307), .A2(n5503), .ZN(n4142) );
  OAI22_X1 U5085 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4880), .ZN(n5430) );
  NAND2_X1 U5086 ( .A1(n5445), .A2(n5430), .ZN(n4145) );
  NAND2_X1 U5087 ( .A1(n2977), .A2(EBX_REG_20__SCAN_IN), .ZN(n4144) );
  OAI211_X1 U5088 ( .C1(n5445), .C2(n2977), .A(n4145), .B(n4144), .ZN(n4146)
         );
  MUX2_X1 U5089 ( .A(n4174), .B(n5444), .S(EBX_REG_21__SCAN_IN), .Z(n4147) );
  OAI21_X1 U5090 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4344), .A(n4147), 
        .ZN(n4148) );
  INV_X1 U5091 ( .A(n4148), .ZN(n5417) );
  NAND2_X1 U5092 ( .A1(n4083), .A2(n6692), .ZN(n4150) );
  INV_X1 U5093 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U5094 ( .A1(n4307), .A2(n5499), .ZN(n4149) );
  NAND3_X1 U5095 ( .A1(n4150), .A2(n5444), .A3(n4149), .ZN(n4152) );
  NAND2_X1 U5096 ( .A1(n2977), .A2(n5499), .ZN(n4151) );
  AND2_X1 U5097 ( .A1(n4152), .A2(n4151), .ZN(n5496) );
  OR2_X2 U5098 ( .A1(n5497), .A2(n5496), .ZN(n5736) );
  MUX2_X1 U5099 ( .A(n4174), .B(n5444), .S(EBX_REG_23__SCAN_IN), .Z(n4153) );
  OAI21_X1 U5100 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n4344), .A(n4153), 
        .ZN(n5737) );
  INV_X1 U5101 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U5102 ( .A1(n4083), .A2(n5728), .ZN(n4155) );
  INV_X1 U5103 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U5104 ( .A1(n4307), .A2(n5489), .ZN(n4154) );
  NAND3_X1 U5105 ( .A1(n4155), .A2(n5444), .A3(n4154), .ZN(n4157) );
  NAND2_X1 U5106 ( .A1(n2977), .A2(n5489), .ZN(n4156) );
  NAND2_X1 U5107 ( .A1(n4157), .A2(n4156), .ZN(n5408) );
  INV_X1 U5108 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U5109 ( .A1(n4158), .A2(n5882), .ZN(n4161) );
  NAND2_X1 U5110 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4159) );
  OAI211_X1 U5111 ( .C1(n4880), .C2(EBX_REG_25__SCAN_IN), .A(n4083), .B(n4159), 
        .ZN(n4160) );
  AND2_X1 U5112 ( .A1(n4161), .A2(n4160), .ZN(n5716) );
  NAND2_X1 U5113 ( .A1(n4083), .A2(n5557), .ZN(n4163) );
  INV_X1 U5114 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U5115 ( .A1(n4307), .A2(n5822), .ZN(n4162) );
  NAND3_X1 U5116 ( .A1(n4163), .A2(n5444), .A3(n4162), .ZN(n4165) );
  NAND2_X1 U5117 ( .A1(n2977), .A2(n5822), .ZN(n4164) );
  AND2_X1 U5118 ( .A1(n4165), .A2(n4164), .ZN(n5486) );
  NAND2_X1 U5119 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4166) );
  OAI211_X1 U5120 ( .C1(n4880), .C2(EBX_REG_27__SCAN_IN), .A(n4083), .B(n4166), 
        .ZN(n4167) );
  OAI21_X1 U5121 ( .B1(n4174), .B2(EBX_REG_27__SCAN_IN), .A(n4167), .ZN(n5698)
         );
  INV_X1 U5122 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U5123 ( .A1(n4083), .A2(n5689), .ZN(n4169) );
  INV_X1 U5124 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U5125 ( .A1(n4307), .A2(n5481), .ZN(n4168) );
  NAND3_X1 U5126 ( .A1(n4169), .A2(n5444), .A3(n4168), .ZN(n4171) );
  NAND2_X1 U5127 ( .A1(n2977), .A2(n5481), .ZN(n4170) );
  NAND2_X1 U5128 ( .A1(n4171), .A2(n4170), .ZN(n5393) );
  NOR2_X1 U5129 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4173)
         );
  NOR2_X1 U5130 ( .A1(n4880), .A2(EBX_REG_29__SCAN_IN), .ZN(n4172) );
  OR3_X2 U5131 ( .A1(n5395), .A2(n4173), .A3(n4172), .ZN(n5318) );
  NAND2_X1 U5132 ( .A1(n5318), .A2(n5444), .ZN(n5315) );
  MUX2_X1 U5133 ( .A(EBX_REG_29__SCAN_IN), .B(n4173), .S(n5444), .Z(n4176) );
  NOR2_X1 U5134 ( .A1(n4174), .A2(EBX_REG_29__SCAN_IN), .ZN(n4175) );
  NOR2_X1 U5135 ( .A1(n4176), .A2(n4175), .ZN(n5375) );
  NAND2_X1 U5136 ( .A1(n4344), .A2(EBX_REG_30__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U5137 ( .A1(n4880), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4177) );
  AND2_X1 U5138 ( .A1(n4178), .A2(n4177), .ZN(n5317) );
  NAND2_X1 U5139 ( .A1(n5375), .A2(n5317), .ZN(n4179) );
  NAND2_X1 U5140 ( .A1(n5315), .A2(n3100), .ZN(n4182) );
  OAI22_X1 U5141 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4880), .ZN(n4180) );
  INV_X1 U5142 ( .A(n4180), .ZN(n4181) );
  NAND2_X1 U5143 ( .A1(n4494), .A2(n6152), .ZN(n6493) );
  NAND2_X1 U5144 ( .A1(n4183), .A2(n4304), .ZN(n4184) );
  NAND2_X1 U5145 ( .A1(n6493), .A2(n4184), .ZN(n4185) );
  INV_X1 U5146 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6701) );
  NOR2_X1 U5147 ( .A1(n5966), .A2(n6701), .ZN(n5371) );
  NOR2_X1 U5148 ( .A1(n6305), .A2(n6299), .ZN(n6294) );
  NAND3_X1 U5149 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6294), .ZN(n4198) );
  NOR2_X1 U5150 ( .A1(n4186), .A2(n3210), .ZN(n4472) );
  OAI21_X1 U5151 ( .B1(n4472), .B2(n4344), .A(n4187), .ZN(n4190) );
  NAND2_X1 U5152 ( .A1(n3228), .A2(n2977), .ZN(n4189) );
  NAND2_X1 U5153 ( .A1(n3239), .A2(n3210), .ZN(n4188) );
  AND4_X1 U5154 ( .A1(n4191), .A2(n4190), .A3(n4189), .A4(n4188), .ZN(n4193)
         );
  NAND3_X1 U5155 ( .A1(n4194), .A2(n4193), .A3(n4192), .ZN(n4496) );
  OAI21_X1 U5156 ( .B1(n4195), .B2(n4874), .A(n4515), .ZN(n4196) );
  NOR2_X1 U5157 ( .A1(n4496), .A2(n4196), .ZN(n4199) );
  NAND2_X1 U5158 ( .A1(n4199), .A2(n4197), .ZN(n4499) );
  INV_X1 U5159 ( .A(n4499), .ZN(n4232) );
  AOI21_X1 U5160 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6343) );
  NAND2_X1 U5161 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6324) );
  NOR2_X1 U5162 ( .A1(n6343), .A2(n6324), .ZN(n6307) );
  NAND3_X1 U5163 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6307), .ZN(n5125) );
  NAND2_X1 U5164 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4550) );
  NOR2_X1 U5165 ( .A1(n4550), .A2(n6324), .ZN(n4555) );
  NAND3_X1 U5166 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4555), .ZN(n5119) );
  NOR2_X1 U5167 ( .A1(n5119), .A2(n4198), .ZN(n4207) );
  INV_X1 U5168 ( .A(n4207), .ZN(n5965) );
  AND2_X1 U5169 ( .A1(n4234), .A2(n4323), .ZN(n6469) );
  NAND2_X1 U5170 ( .A1(n4204), .A2(n6469), .ZN(n6362) );
  INV_X1 U5171 ( .A(n4199), .ZN(n4200) );
  NAND2_X1 U5172 ( .A1(n4204), .A2(n4200), .ZN(n5950) );
  INV_X1 U5173 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6363) );
  AND2_X1 U5174 ( .A1(n6362), .A2(n6363), .ZN(n4278) );
  NOR2_X1 U5175 ( .A1(n5965), .A2(n4554), .ZN(n5232) );
  NOR3_X1 U5176 ( .A1(n5209), .A2(n5237), .A3(n5974), .ZN(n5957) );
  NAND2_X1 U5177 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5957), .ZN(n5788) );
  INV_X1 U5178 ( .A(n5788), .ZN(n5787) );
  NAND3_X1 U5179 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5787), .ZN(n4208) );
  INV_X1 U5180 ( .A(n4201), .ZN(n4210) );
  NAND2_X1 U5181 ( .A1(n5926), .A2(n4202), .ZN(n5715) );
  NAND2_X1 U5182 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4219) );
  NOR2_X1 U5183 ( .A1(n5686), .A2(n4221), .ZN(n5683) );
  AND4_X1 U5184 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n4045), .ZN(n4203) );
  AOI211_X1 U5185 ( .C1(n5477), .C2(n6340), .A(n5371), .B(n4203), .ZN(n4224)
         );
  INV_X1 U5186 ( .A(n5789), .ZN(n5124) );
  NAND2_X1 U5187 ( .A1(n5950), .A2(n5123), .ZN(n5956) );
  NAND2_X1 U5188 ( .A1(n6363), .A2(n5956), .ZN(n6356) );
  INV_X1 U5189 ( .A(n4204), .ZN(n4205) );
  NAND2_X1 U5190 ( .A1(n4205), .A2(n5966), .ZN(n6361) );
  NAND2_X1 U5191 ( .A1(n6356), .A2(n6361), .ZN(n5122) );
  NOR2_X1 U5192 ( .A1(n6341), .A2(n5122), .ZN(n4206) );
  OAI22_X1 U5193 ( .A1(n5118), .A2(n4207), .B1(n5952), .B2(n4206), .ZN(n5954)
         );
  AND2_X1 U5194 ( .A1(n5789), .A2(n4208), .ZN(n4209) );
  OR2_X1 U5195 ( .A1(n5954), .A2(n4209), .ZN(n5934) );
  NAND2_X1 U5196 ( .A1(n4210), .A2(n5767), .ZN(n4211) );
  AND2_X1 U5197 ( .A1(n5789), .A2(n4211), .ZN(n4212) );
  NOR2_X1 U5198 ( .A1(n5934), .A2(n4212), .ZN(n5754) );
  INV_X1 U5199 ( .A(n4213), .ZN(n4214) );
  NAND2_X1 U5200 ( .A1(n5789), .A2(n4214), .ZN(n4215) );
  NAND2_X1 U5201 ( .A1(n4554), .A2(n5123), .ZN(n4217) );
  NAND2_X1 U5202 ( .A1(n4217), .A2(n4216), .ZN(n4218) );
  NAND2_X1 U5203 ( .A1(n5789), .A2(n4219), .ZN(n4220) );
  NAND2_X1 U5204 ( .A1(n5726), .A2(n4220), .ZN(n5705) );
  AOI21_X1 U5205 ( .B1(n5789), .B2(n4221), .A(n5705), .ZN(n5679) );
  OAI21_X1 U5206 ( .B1(n5124), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5679), 
        .ZN(n5673) );
  AOI21_X1 U5207 ( .B1(n5789), .B2(n5668), .A(n5673), .ZN(n4222) );
  AND2_X1 U5208 ( .A1(n4224), .A2(n4223), .ZN(n4225) );
  NAND2_X1 U5209 ( .A1(n4226), .A2(n4225), .ZN(U2987) );
  AND2_X1 U5210 ( .A1(n4234), .A2(n4228), .ZN(n4242) );
  OAI22_X1 U5211 ( .A1(n4480), .A2(n3237), .B1(n4227), .B2(n4242), .ZN(n5982)
         );
  NAND2_X1 U5212 ( .A1(n6616), .A2(n4186), .ZN(n4244) );
  AOI21_X1 U5213 ( .B1(n4244), .B2(n6517), .A(READY_N), .ZN(n6615) );
  NOR2_X1 U5214 ( .A1(n5982), .A2(n6615), .ZN(n6483) );
  INV_X1 U5215 ( .A(n6490), .ZN(n6502) );
  OR2_X1 U5216 ( .A1(n6483), .A2(n6502), .ZN(n5988) );
  INV_X1 U5217 ( .A(n5988), .ZN(n4240) );
  INV_X1 U5218 ( .A(MORE_REG_SCAN_IN), .ZN(n4239) );
  OR2_X1 U5219 ( .A1(n4229), .A2(n4227), .ZN(n4230) );
  NOR2_X1 U5220 ( .A1(n4230), .A2(n4479), .ZN(n4231) );
  OR2_X1 U5221 ( .A1(n4480), .A2(n4231), .ZN(n4237) );
  NAND2_X1 U5222 ( .A1(n4480), .A2(n4232), .ZN(n4236) );
  NAND2_X1 U5223 ( .A1(n4234), .A2(n4233), .ZN(n4235) );
  AND3_X1 U5224 ( .A1(n4237), .A2(n4236), .A3(n4235), .ZN(n6485) );
  OR2_X1 U5225 ( .A1(n5988), .A2(n6485), .ZN(n4238) );
  OAI21_X1 U5226 ( .B1(n4240), .B2(n4239), .A(n4238), .ZN(U3471) );
  AND2_X1 U5227 ( .A1(n4807), .A2(n6592), .ZN(n4883) );
  INV_X1 U5228 ( .A(n4883), .ZN(n4241) );
  NAND2_X1 U5229 ( .A1(n6150), .A2(n4241), .ZN(n5803) );
  NAND2_X1 U5230 ( .A1(n4242), .A2(n6490), .ZN(n5804) );
  INV_X1 U5231 ( .A(n5804), .ZN(n4243) );
  OR3_X1 U5232 ( .A1(n5803), .A2(n4243), .A3(READREQUEST_REG_SCAN_IN), .ZN(
        n4246) );
  NAND2_X1 U5233 ( .A1(n6614), .A2(n4244), .ZN(n4245) );
  AND2_X1 U5234 ( .A1(n4246), .A2(n4245), .ZN(U3474) );
  INV_X1 U5235 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6163) );
  INV_X1 U5236 ( .A(n6517), .ZN(n4872) );
  OAI21_X1 U5237 ( .B1(n6469), .B2(n4494), .A(n4872), .ZN(n4471) );
  NOR2_X1 U5238 ( .A1(n6469), .A2(n6152), .ZN(n4247) );
  NOR2_X1 U5239 ( .A1(n4471), .A2(n4247), .ZN(n4248) );
  NAND2_X1 U5240 ( .A1(n6129), .A2(n4874), .ZN(n4602) );
  NOR2_X1 U5241 ( .A1(n6592), .A2(n5007), .ZN(n4528) );
  INV_X1 U5242 ( .A(n4528), .ZN(n4530) );
  NOR2_X1 U5243 ( .A1(n4530), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4600) );
  AOI22_X1 U5244 ( .A1(n6609), .A2(UWORD_REG_4__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4249) );
  OAI21_X1 U5245 ( .B1(n6163), .B2(n4602), .A(n4249), .ZN(U2903) );
  INV_X1 U5246 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6158) );
  AOI22_X1 U5247 ( .A1(n6609), .A2(UWORD_REG_2__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4250) );
  OAI21_X1 U5248 ( .B1(n6158), .B2(n4602), .A(n4250), .ZN(U2905) );
  INV_X1 U5249 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6160) );
  AOI22_X1 U5250 ( .A1(n6609), .A2(UWORD_REG_3__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4251) );
  OAI21_X1 U5251 ( .B1(n6160), .B2(n4602), .A(n4251), .ZN(U2904) );
  INV_X1 U5252 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6174) );
  AOI22_X1 U5253 ( .A1(n4600), .A2(UWORD_REG_8__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4252) );
  OAI21_X1 U5254 ( .B1(n6174), .B2(n4602), .A(n4252), .ZN(U2899) );
  AOI22_X1 U5255 ( .A1(n4600), .A2(UWORD_REG_12__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4253) );
  OAI21_X1 U5256 ( .B1(n4006), .B2(n4602), .A(n4253), .ZN(U2895) );
  INV_X1 U5257 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6182) );
  AOI22_X1 U5258 ( .A1(n4600), .A2(UWORD_REG_13__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4254) );
  OAI21_X1 U5259 ( .B1(n6182), .B2(n4602), .A(n4254), .ZN(U2894) );
  INV_X1 U5260 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6168) );
  AOI22_X1 U5261 ( .A1(n4600), .A2(UWORD_REG_6__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4255) );
  OAI21_X1 U5262 ( .B1(n6168), .B2(n4602), .A(n4255), .ZN(U2901) );
  INV_X1 U5263 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6165) );
  AOI22_X1 U5264 ( .A1(n4600), .A2(UWORD_REG_5__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4256) );
  OAI21_X1 U5265 ( .B1(n6165), .B2(n4602), .A(n4256), .ZN(U2902) );
  INV_X1 U5266 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6764) );
  AOI22_X1 U5267 ( .A1(n4600), .A2(UWORD_REG_9__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4257) );
  OAI21_X1 U5268 ( .B1(n6764), .B2(n4602), .A(n4257), .ZN(U2898) );
  AOI22_X1 U5269 ( .A1(n4600), .A2(UWORD_REG_10__SCAN_IN), .B1(n5802), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4258) );
  OAI21_X1 U5270 ( .B1(n3964), .B2(n4602), .A(n4258), .ZN(U2897) );
  INV_X1 U5271 ( .A(n4284), .ZN(n4381) );
  NAND2_X1 U5272 ( .A1(n4655), .A2(n4381), .ZN(n4616) );
  NOR3_X1 U5273 ( .A1(n4616), .A2(n4259), .A3(n5987), .ZN(n4260) );
  NOR2_X1 U5274 ( .A1(n4260), .A2(n5799), .ZN(n4267) );
  INV_X1 U5275 ( .A(n4267), .ZN(n4264) );
  NOR2_X1 U5276 ( .A1(n4261), .A2(n4262), .ZN(n5058) );
  INV_X1 U5277 ( .A(n4263), .ZN(n5060) );
  AND2_X1 U5278 ( .A1(n5058), .A2(n5060), .ZN(n4567) );
  NAND3_X1 U5279 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6768), .A3(n4704), .ZN(n4569) );
  NOR2_X1 U5280 ( .A1(n5005), .A2(n4569), .ZN(n4369) );
  AOI21_X1 U5281 ( .B1(n4567), .B2(n2985), .A(n4369), .ZN(n4266) );
  OAI22_X1 U5282 ( .A1(n4264), .A2(n4266), .B1(n4569), .B2(n5007), .ZN(n4265)
         );
  NAND2_X1 U5283 ( .A1(n6592), .A2(n5007), .ZN(n6508) );
  INV_X1 U5284 ( .A(n6508), .ZN(n6617) );
  AND2_X1 U5285 ( .A1(DATAI_7_), .A2(n4442), .ZN(n6461) );
  INV_X1 U5286 ( .A(n5799), .ZN(n6612) );
  INV_X1 U5287 ( .A(n4569), .ZN(n4269) );
  NAND2_X1 U5288 ( .A1(n4267), .A2(n4266), .ZN(n4268) );
  OAI21_X1 U5289 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6589), .A(n4442), 
        .ZN(n4812) );
  OAI211_X1 U5290 ( .C1(n6612), .C2(n4269), .A(n4268), .B(n5016), .ZN(n4372)
         );
  NAND2_X1 U5291 ( .A1(n4372), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U5292 ( .A1(n6258), .A2(DATAI_23_), .ZN(n4976) );
  INV_X1 U5293 ( .A(n4976), .ZN(n6458) );
  NOR2_X1 U5294 ( .A1(n4616), .A2(n4703), .ZN(n4739) );
  NAND2_X1 U5295 ( .A1(n4739), .A2(n4702), .ZN(n4635) );
  INV_X1 U5296 ( .A(n4616), .ZN(n4270) );
  NAND3_X1 U5297 ( .A1(n4270), .A2(n4702), .A3(n4703), .ZN(n4793) );
  NAND2_X1 U5298 ( .A1(n6258), .A2(DATAI_31_), .ZN(n6466) );
  NOR2_X1 U5299 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6589), .ZN(n5329) );
  NAND2_X1 U5300 ( .A1(n4337), .A2(n4645), .ZN(n5177) );
  INV_X1 U5301 ( .A(n4369), .ZN(n4272) );
  OAI22_X1 U5302 ( .A1(n4793), .A2(n6466), .B1(n5177), .B2(n4272), .ZN(n4273)
         );
  AOI21_X1 U5303 ( .B1(n6458), .B2(n6401), .A(n4273), .ZN(n4274) );
  OAI211_X1 U5304 ( .C1(n4374), .C2(n5174), .A(n4275), .B(n4274), .ZN(U3067)
         );
  XNOR2_X1 U5305 ( .A(n4277), .B(n4276), .ZN(n6263) );
  INV_X1 U5306 ( .A(n5122), .ZN(n4280) );
  OR2_X1 U5307 ( .A1(n5124), .A2(n4278), .ZN(n4279) );
  MUX2_X1 U5308 ( .A(n4280), .B(n4279), .S(n5324), .Z(n4283) );
  XNOR2_X1 U5309 ( .A(n4281), .B(n4880), .ZN(n4924) );
  INV_X1 U5310 ( .A(n4924), .ZN(n4379) );
  INV_X1 U5311 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6599) );
  NOR2_X1 U5312 ( .A1(n5966), .A2(n6599), .ZN(n6266) );
  AOI21_X1 U5313 ( .B1(n6340), .B2(n4379), .A(n6266), .ZN(n4282) );
  OAI211_X1 U5314 ( .C1(n6263), .C2(n6313), .A(n4283), .B(n4282), .ZN(U3017)
         );
  AND2_X1 U5315 ( .A1(n4259), .A2(n4284), .ZN(n4285) );
  AND2_X1 U5316 ( .A1(n4655), .A2(n4285), .ZN(n4296) );
  NAND2_X1 U5317 ( .A1(n6612), .A2(n5987), .ZN(n5136) );
  OAI21_X1 U5318 ( .B1(n4296), .B2(n6271), .A(n5136), .ZN(n4289) );
  AND2_X1 U5319 ( .A1(n2990), .A2(n2985), .ZN(n4705) );
  INV_X1 U5320 ( .A(n4261), .ZN(n4287) );
  AND2_X1 U5321 ( .A1(n4262), .A2(n4287), .ZN(n4617) );
  INV_X1 U5322 ( .A(n4338), .ZN(n4288) );
  AOI21_X1 U5323 ( .B1(n4705), .B2(n4617), .A(n4288), .ZN(n4291) );
  NAND2_X1 U5324 ( .A1(n4289), .A2(n4291), .ZN(n4290) );
  OAI211_X1 U5325 ( .C1(n6612), .C2(n4293), .A(n4290), .B(n5016), .ZN(n4341)
         );
  INV_X1 U5326 ( .A(n4291), .ZN(n4292) );
  NAND2_X1 U5327 ( .A1(n4292), .A2(n6612), .ZN(n4295) );
  NAND2_X1 U5328 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4293), .ZN(n4294) );
  AND2_X1 U5329 ( .A1(n4295), .A2(n4294), .ZN(n4343) );
  OAI22_X1 U5330 ( .A1(n5177), .A2(n4338), .B1(n4343), .B2(n5174), .ZN(n4298)
         );
  OAI22_X1 U5331 ( .A1(n4542), .A2(n6466), .B1(n4976), .B2(n4690), .ZN(n4297)
         );
  AOI211_X1 U5332 ( .C1(INSTQUEUE_REG_15__7__SCAN_IN), .C2(n4341), .A(n4298), 
        .B(n4297), .ZN(n4299) );
  INV_X1 U5333 ( .A(n4299), .ZN(U3147) );
  NAND2_X1 U5334 ( .A1(n4301), .A2(n4300), .ZN(n4302) );
  NAND2_X1 U5335 ( .A1(n4781), .A2(n4302), .ZN(n4955) );
  OR2_X1 U5336 ( .A1(n4480), .A2(n4499), .ZN(n4477) );
  NAND3_X1 U5337 ( .A1(n4305), .A2(n4304), .A3(n4303), .ZN(n4306) );
  OR2_X1 U5338 ( .A1(n4306), .A2(n3209), .ZN(n4636) );
  INV_X1 U5339 ( .A(n4636), .ZN(n4308) );
  NAND2_X1 U5340 ( .A1(n4308), .A2(n4307), .ZN(n4309) );
  NAND2_X1 U5341 ( .A1(n4477), .A2(n4309), .ZN(n4310) );
  NOR2_X1 U5342 ( .A1(n4698), .A2(n4311), .ZN(n4312) );
  OR2_X1 U5343 ( .A1(n4562), .A2(n4312), .ZN(n4945) );
  OAI22_X1 U5344 ( .A1(n5885), .A2(n4945), .B1(n4950), .B2(n6118), .ZN(n4313)
         );
  INV_X1 U5345 ( .A(n4313), .ZN(n4314) );
  OAI21_X1 U5346 ( .B1(n4955), .B2(n5886), .A(n4314), .ZN(U2855) );
  NAND2_X1 U5347 ( .A1(n4337), .A2(n4315), .ZN(n6416) );
  NAND2_X1 U5348 ( .A1(n6258), .A2(DATAI_20_), .ZN(n6418) );
  OAI22_X1 U5349 ( .A1(n6416), .A2(n4338), .B1(n4690), .B2(n6418), .ZN(n4317)
         );
  NAND2_X1 U5350 ( .A1(n6258), .A2(DATAI_28_), .ZN(n6427) );
  NOR2_X1 U5351 ( .A1(n4542), .A2(n6427), .ZN(n4316) );
  AOI211_X1 U5352 ( .C1(INSTQUEUE_REG_15__4__SCAN_IN), .C2(n4341), .A(n4317), 
        .B(n4316), .ZN(n4318) );
  OAI21_X1 U5353 ( .B1(n4343), .B2(n5089), .A(n4318), .ZN(U3144) );
  INV_X1 U5354 ( .A(DATAI_6_), .ZN(n4654) );
  NAND2_X1 U5355 ( .A1(n4337), .A2(n4319), .ZN(n5164) );
  NAND2_X1 U5356 ( .A1(n6258), .A2(DATAI_22_), .ZN(n5165) );
  OAI22_X1 U5357 ( .A1(n5164), .A2(n4338), .B1(n4690), .B2(n5165), .ZN(n4321)
         );
  NAND2_X1 U5358 ( .A1(n6258), .A2(DATAI_30_), .ZN(n6386) );
  NOR2_X1 U5359 ( .A1(n4542), .A2(n6386), .ZN(n4320) );
  AOI211_X1 U5360 ( .C1(INSTQUEUE_REG_15__6__SCAN_IN), .C2(n4341), .A(n4321), 
        .B(n4320), .ZN(n4322) );
  OAI21_X1 U5361 ( .B1(n4343), .B2(n5084), .A(n4322), .ZN(U3146) );
  INV_X1 U5362 ( .A(DATAI_1_), .ZN(n4653) );
  INV_X1 U5363 ( .A(n6436), .ZN(n5093) );
  NAND2_X1 U5364 ( .A1(n4337), .A2(n4323), .ZN(n5146) );
  NAND2_X1 U5365 ( .A1(n6258), .A2(DATAI_17_), .ZN(n6395) );
  OAI22_X1 U5366 ( .A1(n5146), .A2(n4338), .B1(n4690), .B2(n6395), .ZN(n4325)
         );
  NAND2_X1 U5367 ( .A1(n6258), .A2(DATAI_25_), .ZN(n6439) );
  NOR2_X1 U5368 ( .A1(n4542), .A2(n6439), .ZN(n4324) );
  AOI211_X1 U5369 ( .C1(INSTQUEUE_REG_15__1__SCAN_IN), .C2(n4341), .A(n4325), 
        .B(n4324), .ZN(n4326) );
  OAI21_X1 U5370 ( .B1(n4343), .B2(n5093), .A(n4326), .ZN(U3141) );
  INV_X1 U5371 ( .A(DATAI_0_), .ZN(n6689) );
  NAND2_X1 U5372 ( .A1(n4337), .A2(n4874), .ZN(n6406) );
  NAND2_X1 U5373 ( .A1(n6258), .A2(DATAI_16_), .ZN(n6407) );
  OAI22_X1 U5374 ( .A1(n6406), .A2(n4338), .B1(n4690), .B2(n6407), .ZN(n4328)
         );
  NAND2_X1 U5375 ( .A1(n6258), .A2(DATAI_24_), .ZN(n6433) );
  NOR2_X1 U5376 ( .A1(n4542), .A2(n6433), .ZN(n4327) );
  AOI211_X1 U5377 ( .C1(INSTQUEUE_REG_15__0__SCAN_IN), .C2(n4341), .A(n4328), 
        .B(n4327), .ZN(n4329) );
  OAI21_X1 U5378 ( .B1(n4343), .B2(n5097), .A(n4329), .ZN(U3140) );
  INV_X1 U5379 ( .A(DATAI_3_), .ZN(n4651) );
  INV_X1 U5380 ( .A(n6446), .ZN(n5074) );
  NAND2_X1 U5381 ( .A1(n4337), .A2(n4330), .ZN(n6411) );
  NAND2_X1 U5382 ( .A1(n6258), .A2(DATAI_19_), .ZN(n6412) );
  OAI22_X1 U5383 ( .A1(n6411), .A2(n4338), .B1(n4690), .B2(n6412), .ZN(n4332)
         );
  NAND2_X1 U5384 ( .A1(n6258), .A2(DATAI_27_), .ZN(n6449) );
  NOR2_X1 U5385 ( .A1(n4542), .A2(n6449), .ZN(n4331) );
  AOI211_X1 U5386 ( .C1(INSTQUEUE_REG_15__3__SCAN_IN), .C2(n4341), .A(n4332), 
        .B(n4331), .ZN(n4333) );
  OAI21_X1 U5387 ( .B1(n4343), .B2(n5074), .A(n4333), .ZN(U3143) );
  INV_X1 U5388 ( .A(DATAI_5_), .ZN(n4782) );
  INV_X1 U5389 ( .A(n6452), .ZN(n5104) );
  NAND2_X1 U5390 ( .A1(n4337), .A2(n3155), .ZN(n5156) );
  NAND2_X1 U5391 ( .A1(n6258), .A2(DATAI_21_), .ZN(n5157) );
  OAI22_X1 U5392 ( .A1(n5156), .A2(n4338), .B1(n4690), .B2(n5157), .ZN(n4335)
         );
  NAND2_X1 U5393 ( .A1(n6258), .A2(DATAI_29_), .ZN(n6455) );
  NOR2_X1 U5394 ( .A1(n4542), .A2(n6455), .ZN(n4334) );
  AOI211_X1 U5395 ( .C1(INSTQUEUE_REG_15__5__SCAN_IN), .C2(n4341), .A(n4335), 
        .B(n4334), .ZN(n4336) );
  OAI21_X1 U5396 ( .B1(n4343), .B2(n5104), .A(n4336), .ZN(U3145) );
  INV_X1 U5397 ( .A(DATAI_2_), .ZN(n4647) );
  NAND2_X1 U5398 ( .A1(n4337), .A2(n3210), .ZN(n6789) );
  NAND2_X1 U5399 ( .A1(n6258), .A2(DATAI_18_), .ZN(n6794) );
  OAI22_X1 U5400 ( .A1(n6789), .A2(n4338), .B1(n4690), .B2(n6794), .ZN(n4340)
         );
  NAND2_X1 U5401 ( .A1(n6258), .A2(DATAI_26_), .ZN(n6786) );
  NOR2_X1 U5402 ( .A1(n4542), .A2(n6786), .ZN(n4339) );
  AOI211_X1 U5403 ( .C1(INSTQUEUE_REG_15__2__SCAN_IN), .C2(n4341), .A(n4340), 
        .B(n4339), .ZN(n4342) );
  OAI21_X1 U5404 ( .B1(n4343), .B2(n5070), .A(n4342), .ZN(U3142) );
  NOR2_X1 U5405 ( .A1(n4344), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4346)
         );
  OR2_X1 U5406 ( .A1(n4346), .A2(n4345), .ZN(n6357) );
  OR2_X1 U5407 ( .A1(n4348), .A2(n4347), .ZN(n4349) );
  NAND2_X1 U5408 ( .A1(n4350), .A2(n4349), .ZN(n6270) );
  OAI222_X1 U5409 ( .A1(n6357), .A2(n5885), .B1(n4084), .B2(n6118), .C1(n6270), 
        .C2(n5886), .ZN(U2859) );
  INV_X1 U5410 ( .A(n6786), .ZN(n6396) );
  INV_X1 U5411 ( .A(n6789), .ZN(n6440) );
  AOI22_X1 U5412 ( .A1(n4787), .A2(n6396), .B1(n6440), .B2(n4369), .ZN(n4351)
         );
  OAI21_X1 U5413 ( .B1(n6794), .B2(n4635), .A(n4351), .ZN(n4352) );
  AOI21_X1 U5414 ( .B1(INSTQUEUE_REG_5__2__SCAN_IN), .B2(n4372), .A(n4352), 
        .ZN(n4353) );
  OAI21_X1 U5415 ( .B1(n4374), .B2(n5070), .A(n4353), .ZN(U3062) );
  INV_X1 U5416 ( .A(n6455), .ZN(n5101) );
  INV_X1 U5417 ( .A(n5156), .ZN(n6450) );
  AOI22_X1 U5418 ( .A1(n4787), .A2(n5101), .B1(n6450), .B2(n4369), .ZN(n4354)
         );
  OAI21_X1 U5419 ( .B1(n5157), .B2(n4635), .A(n4354), .ZN(n4355) );
  AOI21_X1 U5420 ( .B1(INSTQUEUE_REG_5__5__SCAN_IN), .B2(n4372), .A(n4355), 
        .ZN(n4356) );
  OAI21_X1 U5421 ( .B1(n4374), .B2(n5104), .A(n4356), .ZN(U3065) );
  INV_X1 U5422 ( .A(n6386), .ZN(n5081) );
  INV_X1 U5423 ( .A(n5164), .ZN(n6378) );
  AOI22_X1 U5424 ( .A1(n4787), .A2(n5081), .B1(n6378), .B2(n4369), .ZN(n4357)
         );
  OAI21_X1 U5425 ( .B1(n5165), .B2(n4635), .A(n4357), .ZN(n4358) );
  AOI21_X1 U5426 ( .B1(INSTQUEUE_REG_5__6__SCAN_IN), .B2(n4372), .A(n4358), 
        .ZN(n4359) );
  OAI21_X1 U5427 ( .B1(n4374), .B2(n5084), .A(n4359), .ZN(U3066) );
  INV_X1 U5428 ( .A(n6449), .ZN(n6402) );
  INV_X1 U5429 ( .A(n6411), .ZN(n6444) );
  AOI22_X1 U5430 ( .A1(n4787), .A2(n6402), .B1(n6444), .B2(n4369), .ZN(n4360)
         );
  OAI21_X1 U5431 ( .B1(n6412), .B2(n4635), .A(n4360), .ZN(n4361) );
  AOI21_X1 U5432 ( .B1(INSTQUEUE_REG_5__3__SCAN_IN), .B2(n4372), .A(n4361), 
        .ZN(n4362) );
  OAI21_X1 U5433 ( .B1(n4374), .B2(n5074), .A(n4362), .ZN(U3063) );
  INV_X1 U5434 ( .A(n6433), .ZN(n6389) );
  INV_X1 U5435 ( .A(n6406), .ZN(n6428) );
  AOI22_X1 U5436 ( .A1(n4787), .A2(n6389), .B1(n6428), .B2(n4369), .ZN(n4363)
         );
  OAI21_X1 U5437 ( .B1(n6407), .B2(n4635), .A(n4363), .ZN(n4364) );
  AOI21_X1 U5438 ( .B1(INSTQUEUE_REG_5__0__SCAN_IN), .B2(n4372), .A(n4364), 
        .ZN(n4365) );
  OAI21_X1 U5439 ( .B1(n4374), .B2(n5097), .A(n4365), .ZN(U3060) );
  INV_X1 U5440 ( .A(n6439), .ZN(n6392) );
  INV_X1 U5441 ( .A(n5146), .ZN(n6434) );
  AOI22_X1 U5442 ( .A1(n4787), .A2(n6392), .B1(n6434), .B2(n4369), .ZN(n4366)
         );
  OAI21_X1 U5443 ( .B1(n6395), .B2(n4635), .A(n4366), .ZN(n4367) );
  AOI21_X1 U5444 ( .B1(INSTQUEUE_REG_5__1__SCAN_IN), .B2(n4372), .A(n4367), 
        .ZN(n4368) );
  OAI21_X1 U5445 ( .B1(n4374), .B2(n5093), .A(n4368), .ZN(U3061) );
  INV_X1 U5446 ( .A(n6427), .ZN(n5086) );
  INV_X1 U5447 ( .A(n6416), .ZN(n6371) );
  AOI22_X1 U5448 ( .A1(n4787), .A2(n5086), .B1(n6371), .B2(n4369), .ZN(n4370)
         );
  OAI21_X1 U5449 ( .B1(n6418), .B2(n4635), .A(n4370), .ZN(n4371) );
  AOI21_X1 U5450 ( .B1(INSTQUEUE_REG_5__4__SCAN_IN), .B2(n4372), .A(n4371), 
        .ZN(n4373) );
  OAI21_X1 U5451 ( .B1(n4374), .B2(n5089), .A(n4373), .ZN(U3064) );
  NOR2_X1 U5452 ( .A1(n4376), .A2(n4375), .ZN(n4377) );
  OR2_X1 U5453 ( .A1(n4378), .A2(n4377), .ZN(n6268) );
  INV_X1 U5454 ( .A(n6118), .ZN(n5517) );
  AOI22_X1 U5455 ( .A1(n6115), .A2(n4379), .B1(EBX_REG_1__SCAN_IN), .B2(n5517), 
        .ZN(n4380) );
  OAI21_X1 U5456 ( .B1(n5886), .B2(n6268), .A(n4380), .ZN(U2858) );
  NOR2_X1 U5457 ( .A1(n4259), .A2(n4381), .ZN(n4382) );
  NAND2_X1 U5458 ( .A1(n4655), .A2(n4382), .ZN(n4389) );
  INV_X1 U5459 ( .A(n4389), .ZN(n4383) );
  NAND3_X1 U5460 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n4704), .ZN(n5063) );
  INV_X1 U5461 ( .A(n5063), .ZN(n4385) );
  NOR2_X1 U5462 ( .A1(n5005), .A2(n5063), .ZN(n4388) );
  AOI21_X1 U5463 ( .B1(n4705), .B2(n5058), .A(n4388), .ZN(n4387) );
  NAND2_X1 U5464 ( .A1(n4383), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4411) );
  NAND3_X1 U5465 ( .A1(n6612), .A2(n4387), .A3(n4411), .ZN(n4384) );
  OAI211_X1 U5466 ( .C1(n6612), .C2(n4385), .A(n5016), .B(n4384), .ZN(n6785)
         );
  NAND2_X1 U5467 ( .A1(n6612), .A2(n4411), .ZN(n4386) );
  OAI22_X1 U5468 ( .A1(n4387), .A2(n4386), .B1(n5007), .B2(n5063), .ZN(n6783)
         );
  AOI22_X1 U5469 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6785), .B1(n6452), 
        .B2(n6783), .ZN(n4392) );
  INV_X1 U5470 ( .A(n4388), .ZN(n6788) );
  OAI22_X1 U5471 ( .A1(n5156), .A2(n6788), .B1(n6787), .B2(n6455), .ZN(n4390)
         );
  INV_X1 U5472 ( .A(n4390), .ZN(n4391) );
  OAI211_X1 U5473 ( .C1(n5157), .C2(n6793), .A(n4392), .B(n4391), .ZN(U3129)
         );
  AOI22_X1 U5474 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6785), .B1(n6436), 
        .B2(n6783), .ZN(n4395) );
  OAI22_X1 U5475 ( .A1(n5146), .A2(n6788), .B1(n6787), .B2(n6439), .ZN(n4393)
         );
  INV_X1 U5476 ( .A(n4393), .ZN(n4394) );
  OAI211_X1 U5477 ( .C1(n6395), .C2(n6793), .A(n4395), .B(n4394), .ZN(U3125)
         );
  AOI22_X1 U5478 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6785), .B1(n6430), 
        .B2(n6783), .ZN(n4398) );
  OAI22_X1 U5479 ( .A1(n6406), .A2(n6788), .B1(n6787), .B2(n6433), .ZN(n4396)
         );
  INV_X1 U5480 ( .A(n4396), .ZN(n4397) );
  OAI211_X1 U5481 ( .C1(n6407), .C2(n6793), .A(n4398), .B(n4397), .ZN(U3124)
         );
  AOI22_X1 U5482 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6785), .B1(n6382), 
        .B2(n6783), .ZN(n4401) );
  OAI22_X1 U5483 ( .A1(n5164), .A2(n6788), .B1(n6787), .B2(n6386), .ZN(n4399)
         );
  INV_X1 U5484 ( .A(n4399), .ZN(n4400) );
  OAI211_X1 U5485 ( .C1(n5165), .C2(n6793), .A(n4401), .B(n4400), .ZN(U3130)
         );
  AOI22_X1 U5486 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6785), .B1(n6461), 
        .B2(n6783), .ZN(n4404) );
  OAI22_X1 U5487 ( .A1(n5177), .A2(n6788), .B1(n6787), .B2(n6466), .ZN(n4402)
         );
  INV_X1 U5488 ( .A(n4402), .ZN(n4403) );
  OAI211_X1 U5489 ( .C1(n4976), .C2(n6793), .A(n4404), .B(n4403), .ZN(U3131)
         );
  AOI22_X1 U5490 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6785), .B1(n6446), 
        .B2(n6783), .ZN(n4407) );
  OAI22_X1 U5491 ( .A1(n6411), .A2(n6788), .B1(n6787), .B2(n6449), .ZN(n4405)
         );
  INV_X1 U5492 ( .A(n4405), .ZN(n4406) );
  OAI211_X1 U5493 ( .C1(n6412), .C2(n6793), .A(n4407), .B(n4406), .ZN(U3127)
         );
  AOI22_X1 U5494 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6785), .B1(n6422), 
        .B2(n6783), .ZN(n4410) );
  OAI22_X1 U5495 ( .A1(n6416), .A2(n6788), .B1(n6787), .B2(n6427), .ZN(n4408)
         );
  INV_X1 U5496 ( .A(n4408), .ZN(n4409) );
  OAI211_X1 U5497 ( .C1(n6418), .C2(n6793), .A(n4410), .B(n4409), .ZN(U3128)
         );
  INV_X1 U5498 ( .A(n4411), .ZN(n4412) );
  NOR2_X1 U5499 ( .A1(n4412), .A2(n4806), .ZN(n4534) );
  NAND2_X1 U5500 ( .A1(n4259), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5797) );
  INV_X1 U5501 ( .A(n5797), .ZN(n4413) );
  NAND3_X1 U5502 ( .A1(n4534), .A2(n4413), .A3(n3079), .ZN(n4414) );
  NAND2_X1 U5503 ( .A1(n4414), .A2(n6612), .ZN(n4422) );
  INV_X1 U5504 ( .A(n2990), .ZN(n6077) );
  AND2_X1 U5505 ( .A1(n4262), .A2(n4261), .ZN(n4809) );
  NAND2_X1 U5506 ( .A1(n6077), .A2(n4809), .ZN(n5144) );
  INV_X1 U5507 ( .A(n2985), .ZN(n4938) );
  OR2_X1 U5508 ( .A1(n5144), .A2(n4938), .ZN(n4416) );
  INV_X1 U5509 ( .A(n4810), .ZN(n4415) );
  NAND2_X1 U5510 ( .A1(n4415), .A2(n6768), .ZN(n6366) );
  NAND2_X1 U5511 ( .A1(n4416), .A2(n6366), .ZN(n4421) );
  INV_X1 U5512 ( .A(n4421), .ZN(n4417) );
  NAND3_X1 U5513 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6768), .A3(n6478), .ZN(n5135) );
  OAI22_X1 U5514 ( .A1(n4422), .A2(n4417), .B1(n5135), .B2(n5007), .ZN(n6381)
         );
  INV_X1 U5515 ( .A(n6381), .ZN(n4431) );
  INV_X1 U5516 ( .A(n6466), .ZN(n4978) );
  OR2_X1 U5517 ( .A1(n4655), .A2(n4702), .ZN(n4418) );
  NOR2_X1 U5518 ( .A1(n4418), .A2(n5008), .ZN(n4816) );
  NOR2_X1 U5519 ( .A1(n4418), .A2(n4703), .ZN(n4818) );
  NAND2_X1 U5520 ( .A1(n4818), .A2(n4657), .ZN(n4791) );
  OAI22_X1 U5521 ( .A1(n4791), .A2(n4976), .B1(n5177), .B2(n6366), .ZN(n4419)
         );
  AOI21_X1 U5522 ( .B1(n4978), .B2(n5179), .A(n4419), .ZN(n4424) );
  AOI21_X1 U5523 ( .B1(n5799), .B2(n5135), .A(n4812), .ZN(n4420) );
  OAI21_X1 U5524 ( .B1(n4422), .B2(n4421), .A(n4420), .ZN(n6383) );
  NAND2_X1 U5525 ( .A1(n6383), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4423) );
  OAI211_X1 U5526 ( .C1(n4431), .C2(n5174), .A(n4424), .B(n4423), .ZN(U3051)
         );
  OAI22_X1 U5527 ( .A1(n4791), .A2(n6395), .B1(n5146), .B2(n6366), .ZN(n4425)
         );
  AOI21_X1 U5528 ( .B1(n6392), .B2(n5179), .A(n4425), .ZN(n4427) );
  NAND2_X1 U5529 ( .A1(n6383), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4426) );
  OAI211_X1 U5530 ( .C1(n4431), .C2(n5093), .A(n4427), .B(n4426), .ZN(U3045)
         );
  OAI22_X1 U5531 ( .A1(n4791), .A2(n6407), .B1(n6406), .B2(n6366), .ZN(n4428)
         );
  AOI21_X1 U5532 ( .B1(n6389), .B2(n5179), .A(n4428), .ZN(n4430) );
  NAND2_X1 U5533 ( .A1(n6383), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4429) );
  OAI211_X1 U5534 ( .C1(n4431), .C2(n5097), .A(n4430), .B(n4429), .ZN(U3044)
         );
  NAND2_X1 U5535 ( .A1(n4433), .A2(n4432), .ZN(n4434) );
  NAND2_X1 U5536 ( .A1(n4697), .A2(n4434), .ZN(n6089) );
  INV_X1 U5537 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4438) );
  NOR2_X1 U5538 ( .A1(n4436), .A2(n4435), .ZN(n4437) );
  NOR2_X1 U5539 ( .A1(n4649), .A2(n4437), .ZN(n6259) );
  INV_X1 U5540 ( .A(n6259), .ZN(n4648) );
  OAI222_X1 U5541 ( .A1(n6089), .A2(n5885), .B1(n4438), .B2(n6118), .C1(n4648), 
        .C2(n5886), .ZN(U2857) );
  AND2_X1 U5542 ( .A1(n2990), .A2(n4807), .ZN(n5053) );
  NAND2_X1 U5543 ( .A1(n5053), .A2(n4617), .ZN(n4440) );
  AND2_X1 U5544 ( .A1(n4443), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5054) );
  NAND3_X1 U5545 ( .A1(n5054), .A2(n5141), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4439) );
  NOR2_X1 U5546 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4441), .ZN(n4448)
         );
  OAI21_X1 U5547 ( .B1(n5141), .B2(n5007), .A(n4442), .ZN(n4960) );
  NOR2_X1 U5548 ( .A1(n4443), .A2(n5007), .ZN(n5142) );
  NOR3_X1 U5549 ( .A1(n4960), .A2(n6768), .A3(n5142), .ZN(n4447) );
  INV_X1 U5550 ( .A(n4617), .ZN(n4612) );
  INV_X1 U5551 ( .A(n6793), .ZN(n4444) );
  OAI21_X1 U5552 ( .B1(n4444), .B2(n4468), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4445) );
  NAND3_X1 U5553 ( .A1(n4612), .A2(n6612), .A3(n4445), .ZN(n4446) );
  OAI211_X1 U5554 ( .C1(n4448), .C2(n6589), .A(n4447), .B(n4446), .ZN(n4545)
         );
  NAND2_X1 U5555 ( .A1(n4545), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4451)
         );
  INV_X1 U5556 ( .A(n6412), .ZN(n6445) );
  INV_X1 U5557 ( .A(n4448), .ZN(n4541) );
  OAI22_X1 U5558 ( .A1(n6411), .A2(n4541), .B1(n6793), .B2(n6449), .ZN(n4449)
         );
  AOI21_X1 U5559 ( .B1(n6445), .B2(n4468), .A(n4449), .ZN(n4450) );
  OAI211_X1 U5560 ( .C1(n4540), .C2(n5074), .A(n4451), .B(n4450), .ZN(U3135)
         );
  NAND2_X1 U5561 ( .A1(n4545), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4454)
         );
  INV_X1 U5562 ( .A(n5165), .ZN(n6379) );
  OAI22_X1 U5563 ( .A1(n5164), .A2(n4541), .B1(n6793), .B2(n6386), .ZN(n4452)
         );
  AOI21_X1 U5564 ( .B1(n6379), .B2(n4468), .A(n4452), .ZN(n4453) );
  OAI211_X1 U5565 ( .C1(n4540), .C2(n5084), .A(n4454), .B(n4453), .ZN(U3138)
         );
  NAND2_X1 U5566 ( .A1(n4545), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4457)
         );
  INV_X1 U5567 ( .A(n6794), .ZN(n6441) );
  OAI22_X1 U5568 ( .A1(n6789), .A2(n4541), .B1(n6793), .B2(n6786), .ZN(n4455)
         );
  AOI21_X1 U5569 ( .B1(n6441), .B2(n4468), .A(n4455), .ZN(n4456) );
  OAI211_X1 U5570 ( .C1(n4540), .C2(n5070), .A(n4457), .B(n4456), .ZN(U3134)
         );
  NAND2_X1 U5571 ( .A1(n4545), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4460)
         );
  INV_X1 U5572 ( .A(n5157), .ZN(n6451) );
  OAI22_X1 U5573 ( .A1(n5156), .A2(n4541), .B1(n6793), .B2(n6455), .ZN(n4458)
         );
  AOI21_X1 U5574 ( .B1(n6451), .B2(n4468), .A(n4458), .ZN(n4459) );
  OAI211_X1 U5575 ( .C1(n4540), .C2(n5104), .A(n4460), .B(n4459), .ZN(U3137)
         );
  NAND2_X1 U5576 ( .A1(n4545), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4463)
         );
  INV_X1 U5577 ( .A(n6418), .ZN(n6372) );
  OAI22_X1 U5578 ( .A1(n6416), .A2(n4541), .B1(n6793), .B2(n6427), .ZN(n4461)
         );
  AOI21_X1 U5579 ( .B1(n6372), .B2(n4468), .A(n4461), .ZN(n4462) );
  OAI211_X1 U5580 ( .C1(n4540), .C2(n5089), .A(n4463), .B(n4462), .ZN(U3136)
         );
  NAND2_X1 U5581 ( .A1(n4545), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4466)
         );
  INV_X1 U5582 ( .A(n6407), .ZN(n6429) );
  OAI22_X1 U5583 ( .A1(n6406), .A2(n4541), .B1(n6793), .B2(n6433), .ZN(n4464)
         );
  AOI21_X1 U5584 ( .B1(n6429), .B2(n4468), .A(n4464), .ZN(n4465) );
  OAI211_X1 U5585 ( .C1(n4540), .C2(n5097), .A(n4466), .B(n4465), .ZN(U3132)
         );
  NAND2_X1 U5586 ( .A1(n4545), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4470)
         );
  INV_X1 U5587 ( .A(n6395), .ZN(n6435) );
  OAI22_X1 U5588 ( .A1(n5146), .A2(n4541), .B1(n6793), .B2(n6439), .ZN(n4467)
         );
  AOI21_X1 U5589 ( .B1(n6435), .B2(n4468), .A(n4467), .ZN(n4469) );
  OAI211_X1 U5590 ( .C1(n4540), .C2(n5093), .A(n4470), .B(n4469), .ZN(U3133)
         );
  AOI21_X1 U5591 ( .B1(n4471), .B2(n4639), .A(READY_N), .ZN(n4476) );
  INV_X1 U5592 ( .A(n4472), .ZN(n4473) );
  NAND2_X1 U5593 ( .A1(n4474), .A2(n4473), .ZN(n4475) );
  AOI21_X1 U5594 ( .B1(n4480), .B2(n4476), .A(n4475), .ZN(n4478) );
  AND2_X1 U5595 ( .A1(n4478), .A2(n4477), .ZN(n4486) );
  NAND2_X1 U5596 ( .A1(n4480), .A2(n4479), .ZN(n4484) );
  INV_X1 U5597 ( .A(n5976), .ZN(n4482) );
  NAND2_X1 U5598 ( .A1(n4482), .A2(n4481), .ZN(n4483) );
  NAND2_X1 U5599 ( .A1(n4484), .A2(n4483), .ZN(n4638) );
  INV_X1 U5600 ( .A(n4638), .ZN(n4485) );
  NAND2_X1 U5601 ( .A1(n4486), .A2(n4485), .ZN(n6470) );
  OR2_X1 U5602 ( .A1(n4487), .A2(n5060), .ZN(n4488) );
  XNOR2_X1 U5603 ( .A(n4488), .B(n5980), .ZN(n5978) );
  OAI22_X1 U5604 ( .A1(n6470), .A2(n5980), .B1(n5976), .B2(n5978), .ZN(n4489)
         );
  NOR2_X1 U5605 ( .A1(n6592), .A2(FLUSH_REG_SCAN_IN), .ZN(n4491) );
  AOI22_X1 U5606 ( .A1(n4489), .A2(n6592), .B1(n4491), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4527) );
  INV_X1 U5607 ( .A(n4491), .ZN(n4525) );
  NAND2_X1 U5608 ( .A1(n4492), .A2(n4195), .ZN(n4493) );
  OR2_X1 U5609 ( .A1(n4494), .A2(n4493), .ZN(n4495) );
  NOR2_X1 U5610 ( .A1(n4496), .A2(n4495), .ZN(n4497) );
  AND2_X1 U5611 ( .A1(n4497), .A2(n5976), .ZN(n5337) );
  NAND2_X1 U5612 ( .A1(n4499), .A2(n4498), .ZN(n4518) );
  XNOR2_X1 U5613 ( .A(n4500), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4504)
         );
  XNOR2_X1 U5614 ( .A(n3108), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4501)
         );
  NAND2_X1 U5615 ( .A1(n6469), .A2(n4501), .ZN(n4502) );
  OAI21_X1 U5616 ( .B1(n4504), .B2(n4515), .A(n4502), .ZN(n4503) );
  AOI21_X1 U5617 ( .B1(n4518), .B2(n4504), .A(n4503), .ZN(n4505) );
  OAI21_X1 U5618 ( .B1(n4261), .B2(n5337), .A(n4505), .ZN(n5327) );
  MUX2_X1 U5619 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5327), .S(n6470), 
        .Z(n6477) );
  OR2_X1 U5620 ( .A1(n6470), .A2(n3109), .ZN(n4522) );
  INV_X1 U5621 ( .A(n5337), .ZN(n6468) );
  NAND2_X1 U5622 ( .A1(n2990), .A2(n6468), .ZN(n4520) );
  INV_X1 U5623 ( .A(n4506), .ZN(n4510) );
  MUX2_X1 U5624 ( .A(n4510), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4500), 
        .Z(n4509) );
  INV_X1 U5625 ( .A(n4507), .ZN(n4508) );
  NAND2_X1 U5626 ( .A1(n4509), .A2(n4508), .ZN(n4517) );
  OAI21_X1 U5627 ( .B1(n4500), .B2(n3109), .A(n4510), .ZN(n4511) );
  NOR2_X1 U5628 ( .A1(n4511), .A2(n3403), .ZN(n5344) );
  XNOR2_X1 U5629 ( .A(n4512), .B(n3109), .ZN(n4513) );
  NAND2_X1 U5630 ( .A1(n6469), .A2(n4513), .ZN(n4514) );
  OAI21_X1 U5631 ( .B1(n5344), .B2(n4515), .A(n4514), .ZN(n4516) );
  AOI21_X1 U5632 ( .B1(n4518), .B2(n4517), .A(n4516), .ZN(n4519) );
  NAND2_X1 U5633 ( .A1(n4520), .A2(n4519), .ZN(n5347) );
  NAND2_X1 U5634 ( .A1(n6470), .A2(n5347), .ZN(n4521) );
  NAND2_X1 U5635 ( .A1(n4522), .A2(n4521), .ZN(n6479) );
  NAND3_X1 U5636 ( .A1(n6477), .A2(n6592), .A3(n6479), .ZN(n4523) );
  OAI211_X1 U5637 ( .C1(n4525), .C2(n4524), .A(n4523), .B(n4527), .ZN(n6488)
         );
  INV_X1 U5638 ( .A(n6488), .ZN(n4526) );
  AOI21_X1 U5639 ( .B1(n4527), .B2(n4490), .A(n4526), .ZN(n4531) );
  NAND2_X1 U5640 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4528), .ZN(n6586) );
  INV_X1 U5641 ( .A(n6586), .ZN(n5328) );
  OAI21_X1 U5642 ( .B1(n4531), .B2(FLUSH_REG_SCAN_IN), .A(n5328), .ZN(n4529)
         );
  NAND2_X1 U5643 ( .A1(n4529), .A2(n4742), .ZN(n6364) );
  NOR2_X1 U5644 ( .A1(n4531), .A2(n4530), .ZN(n6496) );
  AND2_X1 U5645 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6589), .ZN(n5798) );
  OAI22_X1 U5646 ( .A1(n4703), .A2(n5799), .B1(n4938), .B2(n5798), .ZN(n4532)
         );
  OAI21_X1 U5647 ( .B1(n6496), .B2(n4532), .A(n6364), .ZN(n4533) );
  OAI21_X1 U5648 ( .B1(n6364), .B2(n5005), .A(n4533), .ZN(U3465) );
  OR2_X1 U5649 ( .A1(n4616), .A2(n5797), .ZN(n4836) );
  AOI21_X1 U5650 ( .B1(n4534), .B2(n4836), .A(n5799), .ZN(n4536) );
  OAI22_X1 U5651 ( .A1(n4657), .A2(n5136), .B1(n6077), .B2(n5798), .ZN(n4535)
         );
  OAI21_X1 U5652 ( .B1(n4536), .B2(n4535), .A(n6364), .ZN(n4537) );
  OAI21_X1 U5653 ( .B1(n6364), .B2(n6768), .A(n4537), .ZN(U3462) );
  INV_X1 U5654 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6156) );
  AOI22_X1 U5655 ( .A1(n6609), .A2(UWORD_REG_1__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4538) );
  OAI21_X1 U5656 ( .B1(n6156), .B2(n4602), .A(n4538), .ZN(U2906) );
  INV_X1 U5657 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6154) );
  AOI22_X1 U5658 ( .A1(n6609), .A2(UWORD_REG_0__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4539) );
  OAI21_X1 U5659 ( .B1(n6154), .B2(n4602), .A(n4539), .ZN(U2907) );
  OAI22_X1 U5660 ( .A1(n5177), .A2(n4541), .B1(n4540), .B2(n5174), .ZN(n4544)
         );
  OAI22_X1 U5661 ( .A1(n4542), .A2(n4976), .B1(n6466), .B2(n6793), .ZN(n4543)
         );
  AOI211_X1 U5662 ( .C1(n4545), .C2(INSTQUEUE_REG_14__7__SCAN_IN), .A(n4544), 
        .B(n4543), .ZN(n4546) );
  INV_X1 U5663 ( .A(n4546), .ZN(U3139) );
  INV_X1 U5664 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6185) );
  AOI22_X1 U5665 ( .A1(n4600), .A2(UWORD_REG_14__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4547) );
  OAI21_X1 U5666 ( .B1(n6185), .B2(n4602), .A(n4547), .ZN(U2893) );
  INV_X1 U5667 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6179) );
  AOI22_X1 U5668 ( .A1(n4600), .A2(UWORD_REG_11__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4548) );
  OAI21_X1 U5669 ( .B1(n6179), .B2(n4602), .A(n4548), .ZN(U2896) );
  NAND2_X1 U5670 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6307), .ZN(n4549)
         );
  AND2_X1 U5671 ( .A1(n5789), .A2(n4549), .ZN(n4553) );
  INV_X1 U5672 ( .A(n4550), .ZN(n6342) );
  OR2_X1 U5673 ( .A1(n5118), .A2(n6342), .ZN(n4552) );
  NAND2_X1 U5674 ( .A1(n5123), .A2(n5122), .ZN(n4551) );
  NAND2_X1 U5675 ( .A1(n4552), .A2(n4551), .ZN(n6344) );
  NOR2_X1 U5676 ( .A1(n4553), .A2(n6344), .ZN(n6312) );
  INV_X1 U5677 ( .A(n4554), .ZN(n6346) );
  AOI22_X1 U5678 ( .A1(n4555), .A2(n6346), .B1(n6341), .B2(n6307), .ZN(n4556)
         );
  INV_X1 U5679 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6738) );
  AND2_X1 U5680 ( .A1(n4556), .A2(n6738), .ZN(n4566) );
  NAND2_X1 U5681 ( .A1(n4559), .A2(n4558), .ZN(n4560) );
  NAND2_X1 U5682 ( .A1(n4557), .A2(n4560), .ZN(n6242) );
  NAND2_X1 U5683 ( .A1(n6242), .A2(n6354), .ZN(n4565) );
  OR2_X1 U5684 ( .A1(n4562), .A2(n4561), .ZN(n4563) );
  AND2_X1 U5685 ( .A1(n4608), .A2(n4563), .ZN(n4798) );
  AOI22_X1 U5686 ( .A1(n6340), .A2(n4798), .B1(n6338), .B2(REIP_REG_5__SCAN_IN), .ZN(n4564) );
  OAI211_X1 U5687 ( .C1(n6312), .C2(n4566), .A(n4565), .B(n4564), .ZN(U3013)
         );
  AOI21_X1 U5688 ( .B1(n4791), .B2(n4793), .A(n5987), .ZN(n4568) );
  NOR3_X1 U5689 ( .A1(n4568), .A2(n4567), .A3(n5799), .ZN(n4572) );
  NOR2_X1 U5690 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4569), .ZN(n4784)
         );
  INV_X1 U5691 ( .A(n4741), .ZN(n4570) );
  OR2_X1 U5692 ( .A1(n5141), .A2(n4570), .ZN(n4663) );
  AOI21_X1 U5693 ( .B1(n4663), .B2(STATE2_REG_2__SCAN_IN), .A(n4742), .ZN(
        n4659) );
  INV_X1 U5694 ( .A(n5142), .ZN(n4958) );
  OAI211_X1 U5695 ( .C1(n4784), .C2(n6589), .A(n4659), .B(n4958), .ZN(n4571)
         );
  INV_X1 U5696 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4579) );
  NAND3_X1 U5697 ( .A1(n6077), .A2(n4807), .A3(n5058), .ZN(n4575) );
  INV_X1 U5698 ( .A(n4663), .ZN(n4573) );
  NAND2_X1 U5699 ( .A1(n4573), .A2(n5054), .ZN(n4574) );
  NAND2_X1 U5700 ( .A1(n4575), .A2(n4574), .ZN(n4785) );
  AOI22_X1 U5701 ( .A1(n4787), .A2(n6435), .B1(n6434), .B2(n4784), .ZN(n4576)
         );
  OAI21_X1 U5702 ( .B1(n6439), .B2(n4791), .A(n4576), .ZN(n4577) );
  AOI21_X1 U5703 ( .B1(n6436), .B2(n4785), .A(n4577), .ZN(n4578) );
  OAI21_X1 U5704 ( .B1(n4783), .B2(n4579), .A(n4578), .ZN(U3053) );
  INV_X1 U5705 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4583) );
  AOI22_X1 U5706 ( .A1(n4787), .A2(n6451), .B1(n6450), .B2(n4784), .ZN(n4580)
         );
  OAI21_X1 U5707 ( .B1(n6455), .B2(n4791), .A(n4580), .ZN(n4581) );
  AOI21_X1 U5708 ( .B1(n6452), .B2(n4785), .A(n4581), .ZN(n4582) );
  OAI21_X1 U5709 ( .B1(n4783), .B2(n4583), .A(n4582), .ZN(U3057) );
  INV_X1 U5710 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4587) );
  AOI22_X1 U5711 ( .A1(n4787), .A2(n6379), .B1(n6378), .B2(n4784), .ZN(n4584)
         );
  OAI21_X1 U5712 ( .B1(n6386), .B2(n4791), .A(n4584), .ZN(n4585) );
  AOI21_X1 U5713 ( .B1(n6382), .B2(n4785), .A(n4585), .ZN(n4586) );
  OAI21_X1 U5714 ( .B1(n4783), .B2(n4587), .A(n4586), .ZN(U3058) );
  INV_X1 U5715 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4591) );
  AOI22_X1 U5716 ( .A1(n4787), .A2(n6441), .B1(n6440), .B2(n4784), .ZN(n4588)
         );
  OAI21_X1 U5717 ( .B1(n6786), .B2(n4791), .A(n4588), .ZN(n4589) );
  AOI21_X1 U5718 ( .B1(n6784), .B2(n4785), .A(n4589), .ZN(n4590) );
  OAI21_X1 U5719 ( .B1(n4783), .B2(n4591), .A(n4590), .ZN(U3054) );
  INV_X1 U5720 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4595) );
  AOI22_X1 U5721 ( .A1(n4787), .A2(n6445), .B1(n6444), .B2(n4784), .ZN(n4592)
         );
  OAI21_X1 U5722 ( .B1(n6449), .B2(n4791), .A(n4592), .ZN(n4593) );
  AOI21_X1 U5723 ( .B1(n6446), .B2(n4785), .A(n4593), .ZN(n4594) );
  OAI21_X1 U5724 ( .B1(n4783), .B2(n4595), .A(n4594), .ZN(U3055) );
  INV_X1 U5725 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4599) );
  AOI22_X1 U5726 ( .A1(n4787), .A2(n6372), .B1(n6371), .B2(n4784), .ZN(n4596)
         );
  OAI21_X1 U5727 ( .B1(n6427), .B2(n4791), .A(n4596), .ZN(n4597) );
  AOI21_X1 U5728 ( .B1(n6422), .B2(n4785), .A(n4597), .ZN(n4598) );
  OAI21_X1 U5729 ( .B1(n4783), .B2(n4599), .A(n4598), .ZN(U3056) );
  INV_X1 U5730 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6171) );
  AOI22_X1 U5731 ( .A1(n4600), .A2(UWORD_REG_7__SCAN_IN), .B1(
        DATAO_REG_23__SCAN_IN), .B2(n6145), .ZN(n4601) );
  OAI21_X1 U5732 ( .B1(n6171), .B2(n4602), .A(n4601), .ZN(U2900) );
  INV_X1 U5733 ( .A(n4780), .ZN(n4603) );
  NOR2_X1 U5734 ( .A1(n4781), .A2(n4603), .ZN(n4606) );
  INV_X1 U5735 ( .A(n4803), .ZN(n4604) );
  OAI21_X1 U5736 ( .B1(n4606), .B2(n4605), .A(n4604), .ZN(n4916) );
  NAND2_X1 U5737 ( .A1(n4608), .A2(n4607), .ZN(n4609) );
  NAND2_X1 U5738 ( .A1(n6052), .A2(n4609), .ZN(n4882) );
  INV_X1 U5739 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4885) );
  OAI22_X1 U5740 ( .A1(n5885), .A2(n4882), .B1(n4885), .B2(n6118), .ZN(n4610)
         );
  INV_X1 U5741 ( .A(n4610), .ZN(n4611) );
  OAI21_X1 U5742 ( .B1(n4916), .B2(n5886), .A(n4611), .ZN(U2853) );
  INV_X1 U5743 ( .A(n5054), .ZN(n4660) );
  NOR2_X1 U5744 ( .A1(n4660), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4614)
         );
  NOR3_X1 U5745 ( .A1(n4612), .A2(n2990), .A3(n5799), .ZN(n4613) );
  AOI21_X1 U5746 ( .B1(n5141), .B2(n4614), .A(n4613), .ZN(n6388) );
  NAND2_X1 U5747 ( .A1(n4259), .A2(n4703), .ZN(n4615) );
  AOI21_X1 U5748 ( .B1(n4635), .B2(n6426), .A(n5987), .ZN(n4620) );
  NAND2_X1 U5749 ( .A1(n4617), .A2(n5060), .ZN(n4837) );
  NAND2_X1 U5750 ( .A1(n4837), .A2(n6612), .ZN(n4619) );
  INV_X1 U5751 ( .A(n4844), .ZN(n4839) );
  NOR2_X1 U5752 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4839), .ZN(n6399)
         );
  INV_X1 U5753 ( .A(n6399), .ZN(n4630) );
  AOI211_X1 U5754 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4630), .A(n5142), .B(
        n4960), .ZN(n4618) );
  OAI211_X1 U5755 ( .C1(n4620), .C2(n4619), .A(n4618), .B(n6768), .ZN(n6403)
         );
  NAND2_X1 U5756 ( .A1(n6403), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4623) );
  OAI22_X1 U5757 ( .A1(n5164), .A2(n4630), .B1(n6426), .B2(n5165), .ZN(n4621)
         );
  AOI21_X1 U5758 ( .B1(n5081), .B2(n6401), .A(n4621), .ZN(n4622) );
  OAI211_X1 U5759 ( .C1(n6388), .C2(n5084), .A(n4623), .B(n4622), .ZN(U3074)
         );
  NAND2_X1 U5760 ( .A1(n6403), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4626) );
  OAI22_X1 U5761 ( .A1(n6416), .A2(n4630), .B1(n6426), .B2(n6418), .ZN(n4624)
         );
  AOI21_X1 U5762 ( .B1(n5086), .B2(n6401), .A(n4624), .ZN(n4625) );
  OAI211_X1 U5763 ( .C1(n6388), .C2(n5089), .A(n4626), .B(n4625), .ZN(U3072)
         );
  NAND2_X1 U5764 ( .A1(n6403), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4629) );
  OAI22_X1 U5765 ( .A1(n5156), .A2(n4630), .B1(n6426), .B2(n5157), .ZN(n4627)
         );
  AOI21_X1 U5766 ( .B1(n5101), .B2(n6401), .A(n4627), .ZN(n4628) );
  OAI211_X1 U5767 ( .C1(n6388), .C2(n5104), .A(n4629), .B(n4628), .ZN(U3073)
         );
  NAND2_X1 U5768 ( .A1(n6403), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4634) );
  INV_X1 U5769 ( .A(n6426), .ZN(n4632) );
  OAI22_X1 U5770 ( .A1(n5177), .A2(n4630), .B1(n6388), .B2(n5174), .ZN(n4631)
         );
  AOI21_X1 U5771 ( .B1(n6458), .B2(n4632), .A(n4631), .ZN(n4633) );
  OAI211_X1 U5772 ( .C1(n4635), .C2(n6466), .A(n4634), .B(n4633), .ZN(U3075)
         );
  NOR2_X1 U5773 ( .A1(n4636), .A2(n4922), .ZN(n4637) );
  NOR2_X1 U5774 ( .A1(n4639), .A2(READY_N), .ZN(n4640) );
  NAND2_X1 U5775 ( .A1(n4642), .A2(n4645), .ZN(n4643) );
  INV_X1 U5776 ( .A(n3239), .ZN(n4644) );
  AND2_X1 U5777 ( .A1(n3214), .A2(n4645), .ZN(n4646) );
  INV_X1 U5778 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6188) );
  OAI222_X1 U5779 ( .A1(n6270), .A2(n5890), .B1(n5543), .B2(n6689), .C1(n5544), 
        .C2(n6188), .ZN(U2891) );
  INV_X1 U5780 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6199) );
  OAI222_X1 U5781 ( .A1(n4955), .A2(n5890), .B1(n5543), .B2(n6161), .C1(n5544), 
        .C2(n6199), .ZN(U2887) );
  OAI222_X1 U5782 ( .A1(n4648), .A2(n5890), .B1(n5543), .B2(n4647), .C1(n5544), 
        .C2(n3586), .ZN(U2889) );
  XOR2_X1 U5783 ( .A(n4650), .B(n4649), .Z(n6250) );
  INV_X1 U5784 ( .A(n6250), .ZN(n4652) );
  INV_X1 U5785 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6196) );
  OAI222_X1 U5786 ( .A1(n4652), .A2(n5890), .B1(n5543), .B2(n4651), .C1(n5544), 
        .C2(n6196), .ZN(U2888) );
  INV_X1 U5787 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6191) );
  OAI222_X1 U5788 ( .A1(n6268), .A2(n5890), .B1(n5543), .B2(n4653), .C1(n5544), 
        .C2(n6191), .ZN(U2890) );
  OAI222_X1 U5789 ( .A1(n4916), .A2(n5890), .B1(n5543), .B2(n4654), .C1(n5544), 
        .C2(n3620), .ZN(U2885) );
  NOR2_X1 U5790 ( .A1(n4655), .A2(n4259), .ZN(n4656) );
  AOI21_X1 U5791 ( .B1(n5052), .B2(n4690), .A(n5987), .ZN(n4658) );
  INV_X1 U5792 ( .A(n4262), .ZN(n5795) );
  NAND2_X1 U5793 ( .A1(n5795), .A2(n4261), .ZN(n4740) );
  NOR2_X1 U5794 ( .A1(n4740), .A2(n2990), .ZN(n5006) );
  NOR3_X1 U5795 ( .A1(n4658), .A2(n5006), .A3(n5799), .ZN(n4662) );
  NAND3_X1 U5796 ( .A1(n6768), .A2(n6478), .A3(n4704), .ZN(n5012) );
  NOR2_X1 U5797 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5012), .ZN(n4665)
         );
  OAI211_X1 U5798 ( .C1(n6589), .C2(n4665), .A(n4660), .B(n4659), .ZN(n4661)
         );
  NAND2_X1 U5799 ( .A1(n4689), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4668) );
  INV_X1 U5800 ( .A(n5006), .ZN(n4664) );
  OAI22_X1 U5801 ( .A1(n4664), .A2(n5799), .B1(n4958), .B2(n4663), .ZN(n4693)
         );
  INV_X1 U5802 ( .A(n4665), .ZN(n4691) );
  OAI22_X1 U5803 ( .A1(n5146), .A2(n4691), .B1(n4690), .B2(n6439), .ZN(n4666)
         );
  AOI21_X1 U5804 ( .B1(n6436), .B2(n4693), .A(n4666), .ZN(n4667) );
  OAI211_X1 U5805 ( .C1(n5052), .C2(n6395), .A(n4668), .B(n4667), .ZN(U3021)
         );
  NAND2_X1 U5806 ( .A1(n4689), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4671) );
  OAI22_X1 U5807 ( .A1(n6789), .A2(n4691), .B1(n4690), .B2(n6786), .ZN(n4669)
         );
  AOI21_X1 U5808 ( .B1(n6784), .B2(n4693), .A(n4669), .ZN(n4670) );
  OAI211_X1 U5809 ( .C1(n5052), .C2(n6794), .A(n4671), .B(n4670), .ZN(U3022)
         );
  NAND2_X1 U5810 ( .A1(n4689), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4674) );
  OAI22_X1 U5811 ( .A1(n6406), .A2(n4691), .B1(n4690), .B2(n6433), .ZN(n4672)
         );
  AOI21_X1 U5812 ( .B1(n6430), .B2(n4693), .A(n4672), .ZN(n4673) );
  OAI211_X1 U5813 ( .C1(n5052), .C2(n6407), .A(n4674), .B(n4673), .ZN(U3020)
         );
  NAND2_X1 U5814 ( .A1(n4689), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4677) );
  OAI22_X1 U5815 ( .A1(n6416), .A2(n4691), .B1(n4690), .B2(n6427), .ZN(n4675)
         );
  AOI21_X1 U5816 ( .B1(n6422), .B2(n4693), .A(n4675), .ZN(n4676) );
  OAI211_X1 U5817 ( .C1(n5052), .C2(n6418), .A(n4677), .B(n4676), .ZN(U3024)
         );
  NAND2_X1 U5818 ( .A1(n4689), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4680) );
  OAI22_X1 U5819 ( .A1(n5156), .A2(n4691), .B1(n4690), .B2(n6455), .ZN(n4678)
         );
  AOI21_X1 U5820 ( .B1(n6452), .B2(n4693), .A(n4678), .ZN(n4679) );
  OAI211_X1 U5821 ( .C1(n5052), .C2(n5157), .A(n4680), .B(n4679), .ZN(U3025)
         );
  NAND2_X1 U5822 ( .A1(n4689), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4683) );
  OAI22_X1 U5823 ( .A1(n5164), .A2(n4691), .B1(n4690), .B2(n6386), .ZN(n4681)
         );
  AOI21_X1 U5824 ( .B1(n6382), .B2(n4693), .A(n4681), .ZN(n4682) );
  OAI211_X1 U5825 ( .C1(n5052), .C2(n5165), .A(n4683), .B(n4682), .ZN(U3026)
         );
  NAND2_X1 U5826 ( .A1(n4689), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4688) );
  INV_X1 U5827 ( .A(n4690), .ZN(n4686) );
  INV_X1 U5828 ( .A(n4693), .ZN(n4684) );
  OAI22_X1 U5829 ( .A1(n5177), .A2(n4691), .B1(n4684), .B2(n5174), .ZN(n4685)
         );
  AOI21_X1 U5830 ( .B1(n4978), .B2(n4686), .A(n4685), .ZN(n4687) );
  OAI211_X1 U5831 ( .C1(n5052), .C2(n4976), .A(n4688), .B(n4687), .ZN(U3027)
         );
  NAND2_X1 U5832 ( .A1(n4689), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4695) );
  OAI22_X1 U5833 ( .A1(n6411), .A2(n4691), .B1(n4690), .B2(n6449), .ZN(n4692)
         );
  AOI21_X1 U5834 ( .B1(n6446), .B2(n4693), .A(n4692), .ZN(n4694) );
  OAI211_X1 U5835 ( .C1(n5052), .C2(n6412), .A(n4695), .B(n4694), .ZN(U3023)
         );
  AND2_X1 U5836 ( .A1(n4697), .A2(n4696), .ZN(n4699) );
  OR2_X1 U5837 ( .A1(n4699), .A2(n4698), .ZN(n6329) );
  OAI22_X1 U5838 ( .A1(n5885), .A2(n6329), .B1(n6753), .B2(n6118), .ZN(n4700)
         );
  AOI21_X1 U5839 ( .B1(n6250), .B2(n6116), .A(n4700), .ZN(n4701) );
  INV_X1 U5840 ( .A(n4701), .ZN(U2856) );
  AOI21_X1 U5841 ( .B1(n4710), .B2(STATEBS16_REG_SCAN_IN), .A(n5799), .ZN(
        n4707) );
  INV_X1 U5842 ( .A(n4740), .ZN(n4747) );
  NAND3_X1 U5843 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6478), .A3(n4704), .ZN(n4743) );
  NOR2_X1 U5844 ( .A1(n5005), .A2(n4743), .ZN(n4711) );
  AOI21_X1 U5845 ( .B1(n4705), .B2(n4747), .A(n4711), .ZN(n4709) );
  AOI22_X1 U5846 ( .A1(n4707), .A2(n4709), .B1(n5799), .B2(n4743), .ZN(n4706)
         );
  NAND2_X1 U5847 ( .A1(n5016), .A2(n4706), .ZN(n4734) );
  INV_X1 U5848 ( .A(n4707), .ZN(n4708) );
  OAI22_X1 U5849 ( .A1(n4709), .A2(n4708), .B1(n5007), .B2(n4743), .ZN(n4733)
         );
  AOI22_X1 U5850 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4734), .B1(n6422), 
        .B2(n4733), .ZN(n4714) );
  INV_X1 U5851 ( .A(n4711), .ZN(n4735) );
  OAI22_X1 U5852 ( .A1(n4966), .A2(n6418), .B1(n6416), .B2(n4735), .ZN(n4712)
         );
  INV_X1 U5853 ( .A(n4712), .ZN(n4713) );
  OAI211_X1 U5854 ( .C1(n6427), .C2(n4779), .A(n4714), .B(n4713), .ZN(U3096)
         );
  AOI22_X1 U5855 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4734), .B1(n6446), 
        .B2(n4733), .ZN(n4717) );
  OAI22_X1 U5856 ( .A1(n4966), .A2(n6412), .B1(n6411), .B2(n4735), .ZN(n4715)
         );
  INV_X1 U5857 ( .A(n4715), .ZN(n4716) );
  OAI211_X1 U5858 ( .C1(n6449), .C2(n4779), .A(n4717), .B(n4716), .ZN(U3095)
         );
  AOI22_X1 U5859 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4734), .B1(n6461), 
        .B2(n4733), .ZN(n4720) );
  OAI22_X1 U5860 ( .A1(n4966), .A2(n4976), .B1(n5177), .B2(n4735), .ZN(n4718)
         );
  INV_X1 U5861 ( .A(n4718), .ZN(n4719) );
  OAI211_X1 U5862 ( .C1(n6466), .C2(n4779), .A(n4720), .B(n4719), .ZN(U3099)
         );
  AOI22_X1 U5863 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4734), .B1(n6436), 
        .B2(n4733), .ZN(n4723) );
  OAI22_X1 U5864 ( .A1(n4966), .A2(n6395), .B1(n5146), .B2(n4735), .ZN(n4721)
         );
  INV_X1 U5865 ( .A(n4721), .ZN(n4722) );
  OAI211_X1 U5866 ( .C1(n6439), .C2(n4779), .A(n4723), .B(n4722), .ZN(U3093)
         );
  AOI22_X1 U5867 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4734), .B1(n6382), 
        .B2(n4733), .ZN(n4726) );
  OAI22_X1 U5868 ( .A1(n4966), .A2(n5165), .B1(n5164), .B2(n4735), .ZN(n4724)
         );
  INV_X1 U5869 ( .A(n4724), .ZN(n4725) );
  OAI211_X1 U5870 ( .C1(n6386), .C2(n4779), .A(n4726), .B(n4725), .ZN(U3098)
         );
  AOI22_X1 U5871 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4734), .B1(n6784), 
        .B2(n4733), .ZN(n4729) );
  OAI22_X1 U5872 ( .A1(n4966), .A2(n6794), .B1(n6789), .B2(n4735), .ZN(n4727)
         );
  INV_X1 U5873 ( .A(n4727), .ZN(n4728) );
  OAI211_X1 U5874 ( .C1(n6786), .C2(n4779), .A(n4729), .B(n4728), .ZN(U3094)
         );
  AOI22_X1 U5875 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4734), .B1(n6430), 
        .B2(n4733), .ZN(n4732) );
  OAI22_X1 U5876 ( .A1(n4966), .A2(n6407), .B1(n6406), .B2(n4735), .ZN(n4730)
         );
  INV_X1 U5877 ( .A(n4730), .ZN(n4731) );
  OAI211_X1 U5878 ( .C1(n6433), .C2(n4779), .A(n4732), .B(n4731), .ZN(U3092)
         );
  AOI22_X1 U5879 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4734), .B1(n6452), 
        .B2(n4733), .ZN(n4738) );
  OAI22_X1 U5880 ( .A1(n4966), .A2(n5157), .B1(n5156), .B2(n4735), .ZN(n4736)
         );
  INV_X1 U5881 ( .A(n4736), .ZN(n4737) );
  OAI211_X1 U5882 ( .C1(n6455), .C2(n4779), .A(n4738), .B(n4737), .ZN(U3097)
         );
  NAND2_X1 U5883 ( .A1(n4739), .A2(n4259), .ZN(n6419) );
  AOI21_X1 U5884 ( .B1(n4779), .B2(n6419), .A(n5987), .ZN(n4746) );
  OAI21_X1 U5885 ( .B1(n6077), .B2(n4740), .A(n6612), .ZN(n4745) );
  OR2_X1 U5886 ( .A1(n5141), .A2(n4741), .ZN(n4748) );
  AOI21_X1 U5887 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4748), .A(n4742), .ZN(
        n5065) );
  OR2_X1 U5888 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4743), .ZN(n4774)
         );
  AOI21_X1 U5889 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4774), .A(n5054), .ZN(
        n4744) );
  OAI211_X1 U5890 ( .C1(n4746), .C2(n4745), .A(n5065), .B(n4744), .ZN(n4773)
         );
  NAND2_X1 U5891 ( .A1(n4773), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4753) );
  NAND2_X1 U5892 ( .A1(n5053), .A2(n4747), .ZN(n4750) );
  INV_X1 U5893 ( .A(n4748), .ZN(n5055) );
  NAND2_X1 U5894 ( .A1(n5142), .A2(n5055), .ZN(n4749) );
  NAND2_X1 U5895 ( .A1(n4750), .A2(n4749), .ZN(n4776) );
  OAI22_X1 U5896 ( .A1(n6419), .A2(n6427), .B1(n6416), .B2(n4774), .ZN(n4751)
         );
  AOI21_X1 U5897 ( .B1(n6422), .B2(n4776), .A(n4751), .ZN(n4752) );
  OAI211_X1 U5898 ( .C1(n4779), .C2(n6418), .A(n4753), .B(n4752), .ZN(U3088)
         );
  NAND2_X1 U5899 ( .A1(n4773), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4756) );
  OAI22_X1 U5900 ( .A1(n6419), .A2(n6386), .B1(n5164), .B2(n4774), .ZN(n4754)
         );
  AOI21_X1 U5901 ( .B1(n6382), .B2(n4776), .A(n4754), .ZN(n4755) );
  OAI211_X1 U5902 ( .C1(n4779), .C2(n5165), .A(n4756), .B(n4755), .ZN(U3090)
         );
  NAND2_X1 U5903 ( .A1(n4773), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4760) );
  INV_X1 U5904 ( .A(n6419), .ZN(n4860) );
  INV_X1 U5905 ( .A(n4776), .ZN(n4757) );
  OAI22_X1 U5906 ( .A1(n5177), .A2(n4774), .B1(n4757), .B2(n5174), .ZN(n4758)
         );
  AOI21_X1 U5907 ( .B1(n4978), .B2(n4860), .A(n4758), .ZN(n4759) );
  OAI211_X1 U5908 ( .C1(n4779), .C2(n4976), .A(n4760), .B(n4759), .ZN(U3091)
         );
  NAND2_X1 U5909 ( .A1(n4773), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4763) );
  OAI22_X1 U5910 ( .A1(n6419), .A2(n6786), .B1(n6789), .B2(n4774), .ZN(n4761)
         );
  AOI21_X1 U5911 ( .B1(n6784), .B2(n4776), .A(n4761), .ZN(n4762) );
  OAI211_X1 U5912 ( .C1(n4779), .C2(n6794), .A(n4763), .B(n4762), .ZN(U3086)
         );
  NAND2_X1 U5913 ( .A1(n4773), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4766) );
  OAI22_X1 U5914 ( .A1(n6419), .A2(n6455), .B1(n5156), .B2(n4774), .ZN(n4764)
         );
  AOI21_X1 U5915 ( .B1(n6452), .B2(n4776), .A(n4764), .ZN(n4765) );
  OAI211_X1 U5916 ( .C1(n4779), .C2(n5157), .A(n4766), .B(n4765), .ZN(U3089)
         );
  NAND2_X1 U5917 ( .A1(n4773), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4769) );
  OAI22_X1 U5918 ( .A1(n6419), .A2(n6449), .B1(n6411), .B2(n4774), .ZN(n4767)
         );
  AOI21_X1 U5919 ( .B1(n6446), .B2(n4776), .A(n4767), .ZN(n4768) );
  OAI211_X1 U5920 ( .C1(n4779), .C2(n6412), .A(n4769), .B(n4768), .ZN(U3087)
         );
  NAND2_X1 U5921 ( .A1(n4773), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4772) );
  OAI22_X1 U5922 ( .A1(n6419), .A2(n6439), .B1(n5146), .B2(n4774), .ZN(n4770)
         );
  AOI21_X1 U5923 ( .B1(n6436), .B2(n4776), .A(n4770), .ZN(n4771) );
  OAI211_X1 U5924 ( .C1(n4779), .C2(n6395), .A(n4772), .B(n4771), .ZN(U3085)
         );
  NAND2_X1 U5925 ( .A1(n4773), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4778) );
  OAI22_X1 U5926 ( .A1(n6419), .A2(n6433), .B1(n6406), .B2(n4774), .ZN(n4775)
         );
  AOI21_X1 U5927 ( .B1(n6430), .B2(n4776), .A(n4775), .ZN(n4777) );
  OAI211_X1 U5928 ( .C1(n4779), .C2(n6407), .A(n4778), .B(n4777), .ZN(U3084)
         );
  XNOR2_X1 U5929 ( .A(n4781), .B(n4780), .ZN(n6241) );
  INV_X1 U5930 ( .A(n6241), .ZN(n4800) );
  OAI222_X1 U5931 ( .A1(n5890), .A2(n4800), .B1(n5544), .B2(n3614), .C1(n4782), 
        .C2(n5543), .ZN(U2886) );
  INV_X1 U5932 ( .A(n4783), .ZN(n4790) );
  NAND2_X1 U5933 ( .A1(n4790), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4789) );
  INV_X1 U5934 ( .A(n4784), .ZN(n4792) );
  INV_X1 U5935 ( .A(n4785), .ZN(n4797) );
  OAI22_X1 U5936 ( .A1(n5177), .A2(n4792), .B1(n4797), .B2(n5174), .ZN(n4786)
         );
  AOI21_X1 U5937 ( .B1(n6458), .B2(n4787), .A(n4786), .ZN(n4788) );
  OAI211_X1 U5938 ( .C1(n4791), .C2(n6466), .A(n4789), .B(n4788), .ZN(U3059)
         );
  NAND2_X1 U5939 ( .A1(n4790), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4796) );
  INV_X1 U5940 ( .A(n4791), .ZN(n6380) );
  OAI22_X1 U5941 ( .A1(n4793), .A2(n6407), .B1(n6406), .B2(n4792), .ZN(n4794)
         );
  AOI21_X1 U5942 ( .B1(n6389), .B2(n6380), .A(n4794), .ZN(n4795) );
  OAI211_X1 U5943 ( .C1(n4797), .C2(n5097), .A(n4796), .B(n4795), .ZN(U3052)
         );
  INV_X1 U5944 ( .A(n4798), .ZN(n6068) );
  OAI222_X1 U5945 ( .A1(n6068), .A2(n5885), .B1(n5886), .B2(n4800), .C1(n4799), 
        .C2(n6118), .ZN(U2854) );
  INV_X1 U5946 ( .A(n4801), .ZN(n4802) );
  XNOR2_X1 U5947 ( .A(n4803), .B(n4802), .ZN(n6237) );
  INV_X1 U5948 ( .A(n6237), .ZN(n4805) );
  AOI22_X1 U5949 ( .A1(n5538), .A2(DATAI_7_), .B1(EAX_REG_7__SCAN_IN), .B2(
        n6125), .ZN(n4804) );
  OAI21_X1 U5950 ( .B1(n4805), .B2(n5890), .A(n4804), .ZN(U2884) );
  INV_X1 U5951 ( .A(n4806), .ZN(n4808) );
  OAI21_X1 U5952 ( .B1(n4808), .B2(n5797), .A(n4807), .ZN(n4815) );
  AND2_X1 U5953 ( .A1(n4809), .A2(n2990), .ZN(n4961) );
  NOR2_X1 U5954 ( .A1(n4810), .A2(n6768), .ZN(n6456) );
  AOI21_X1 U5955 ( .B1(n4961), .B2(n2985), .A(n6456), .ZN(n4811) );
  NAND3_X1 U5956 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6478), .ZN(n4962) );
  OAI22_X1 U5957 ( .A1(n4815), .A2(n4811), .B1(n4962), .B2(n5007), .ZN(n6460)
         );
  INV_X1 U5958 ( .A(n6460), .ZN(n4825) );
  INV_X1 U5959 ( .A(n4811), .ZN(n4814) );
  AOI21_X1 U5960 ( .B1(n5799), .B2(n4962), .A(n4812), .ZN(n4813) );
  OAI21_X1 U5961 ( .B1(n4815), .B2(n4814), .A(n4813), .ZN(n6462) );
  AOI22_X1 U5962 ( .A1(n6459), .A2(n6372), .B1(n6371), .B2(n6456), .ZN(n4819)
         );
  OAI21_X1 U5963 ( .B1(n6465), .B2(n6427), .A(n4819), .ZN(n4820) );
  AOI21_X1 U5964 ( .B1(n6462), .B2(INSTQUEUE_REG_11__4__SCAN_IN), .A(n4820), 
        .ZN(n4821) );
  OAI21_X1 U5965 ( .B1(n4825), .B2(n5089), .A(n4821), .ZN(U3112) );
  AOI22_X1 U5966 ( .A1(n6459), .A2(n6379), .B1(n6378), .B2(n6456), .ZN(n4822)
         );
  OAI21_X1 U5967 ( .B1(n6465), .B2(n6386), .A(n4822), .ZN(n4823) );
  AOI21_X1 U5968 ( .B1(n6462), .B2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n4823), 
        .ZN(n4824) );
  OAI21_X1 U5969 ( .B1(n4825), .B2(n5084), .A(n4824), .ZN(U3114) );
  OAI21_X1 U5970 ( .B1(n4828), .B2(n4827), .A(n4826), .ZN(n6322) );
  NAND2_X1 U5971 ( .A1(n6338), .A2(REIP_REG_4__SCAN_IN), .ZN(n6319) );
  OAI21_X1 U5972 ( .B1(n5646), .B2(n3604), .A(n6319), .ZN(n4830) );
  NOR2_X1 U5973 ( .A1(n4955), .A2(n6271), .ZN(n4829) );
  AOI211_X1 U5974 ( .C1(n5649), .C2(n4952), .A(n4830), .B(n4829), .ZN(n4831)
         );
  OAI21_X1 U5975 ( .B1(n6273), .B2(n6322), .A(n4831), .ZN(U2982) );
  OR2_X1 U5976 ( .A1(n4833), .A2(n4832), .ZN(n4834) );
  AND2_X1 U5977 ( .A1(n4834), .A2(n4932), .ZN(n4908) );
  AOI22_X1 U5978 ( .A1(n5538), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6125), .ZN(n4835) );
  OAI21_X1 U5979 ( .B1(n4910), .B2(n5890), .A(n4835), .ZN(U2883) );
  NAND2_X1 U5980 ( .A1(n4836), .A2(n6612), .ZN(n4840) );
  INV_X1 U5981 ( .A(n4837), .ZN(n4838) );
  INV_X1 U5982 ( .A(n6417), .ZN(n4857) );
  AOI21_X1 U5983 ( .B1(n4838), .B2(n2985), .A(n4857), .ZN(n4842) );
  OAI22_X1 U5984 ( .A1(n4840), .A2(n4842), .B1(n5007), .B2(n4839), .ZN(n6421)
         );
  INV_X1 U5985 ( .A(n6421), .ZN(n4862) );
  INV_X1 U5986 ( .A(n4840), .ZN(n4841) );
  NAND2_X1 U5987 ( .A1(n4842), .A2(n4841), .ZN(n4843) );
  OAI211_X1 U5988 ( .C1(n4844), .C2(n6612), .A(n5016), .B(n4843), .ZN(n6423)
         );
  AOI22_X1 U5989 ( .A1(n6434), .A2(n4857), .B1(INSTQUEUE_REG_7__1__SCAN_IN), 
        .B2(n6423), .ZN(n4845) );
  OAI21_X1 U5990 ( .B1(n6439), .B2(n6426), .A(n4845), .ZN(n4846) );
  AOI21_X1 U5991 ( .B1(n6435), .B2(n4860), .A(n4846), .ZN(n4847) );
  OAI21_X1 U5992 ( .B1(n4862), .B2(n5093), .A(n4847), .ZN(U3077) );
  AOI22_X1 U5993 ( .A1(n6440), .A2(n4857), .B1(INSTQUEUE_REG_7__2__SCAN_IN), 
        .B2(n6423), .ZN(n4848) );
  OAI21_X1 U5994 ( .B1(n6786), .B2(n6426), .A(n4848), .ZN(n4849) );
  AOI21_X1 U5995 ( .B1(n6441), .B2(n4860), .A(n4849), .ZN(n4850) );
  OAI21_X1 U5996 ( .B1(n4862), .B2(n5070), .A(n4850), .ZN(U3078) );
  AOI22_X1 U5997 ( .A1(n6450), .A2(n4857), .B1(INSTQUEUE_REG_7__5__SCAN_IN), 
        .B2(n6423), .ZN(n4851) );
  OAI21_X1 U5998 ( .B1(n6455), .B2(n6426), .A(n4851), .ZN(n4852) );
  AOI21_X1 U5999 ( .B1(n6451), .B2(n4860), .A(n4852), .ZN(n4853) );
  OAI21_X1 U6000 ( .B1(n4862), .B2(n5104), .A(n4853), .ZN(U3081) );
  AOI22_X1 U6001 ( .A1(n6378), .A2(n4857), .B1(INSTQUEUE_REG_7__6__SCAN_IN), 
        .B2(n6423), .ZN(n4854) );
  OAI21_X1 U6002 ( .B1(n6386), .B2(n6426), .A(n4854), .ZN(n4855) );
  AOI21_X1 U6003 ( .B1(n6379), .B2(n4860), .A(n4855), .ZN(n4856) );
  OAI21_X1 U6004 ( .B1(n4862), .B2(n5084), .A(n4856), .ZN(U3082) );
  INV_X1 U6005 ( .A(n5177), .ZN(n6457) );
  AOI22_X1 U6006 ( .A1(n6457), .A2(n4857), .B1(INSTQUEUE_REG_7__7__SCAN_IN), 
        .B2(n6423), .ZN(n4858) );
  OAI21_X1 U6007 ( .B1(n6466), .B2(n6426), .A(n4858), .ZN(n4859) );
  AOI21_X1 U6008 ( .B1(n6458), .B2(n4860), .A(n4859), .ZN(n4861) );
  OAI21_X1 U6009 ( .B1(n4862), .B2(n5174), .A(n4861), .ZN(U3083) );
  INV_X1 U6010 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5321) );
  XNOR2_X1 U6011 ( .A(n4863), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5369)
         );
  NOR3_X1 U6012 ( .A1(n6669), .A2(n6589), .A3(n6508), .ZN(n6495) );
  INV_X2 U6013 ( .A(n5966), .ZN(n6338) );
  AND2_X1 U6014 ( .A1(n4865), .A2(n4864), .ZN(n6504) );
  OR2_X1 U6015 ( .A1(n6338), .A2(n6504), .ZN(n4866) );
  NAND2_X1 U6016 ( .A1(n6084), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4867) );
  INV_X1 U6017 ( .A(n4867), .ZN(n4868) );
  INV_X1 U6018 ( .A(n6084), .ZN(n5305) );
  INV_X1 U6019 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6534) );
  NAND3_X1 U6020 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n4946) );
  NOR2_X1 U6021 ( .A1(n6534), .A2(n4946), .ZN(n4871) );
  NAND2_X1 U6022 ( .A1(REIP_REG_5__SCAN_IN), .A2(n4871), .ZN(n4889) );
  NOR2_X1 U6023 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4873) );
  AND3_X1 U6024 ( .A1(n4869), .A2(n4873), .A3(n4874), .ZN(n4870) );
  NAND2_X1 U6025 ( .A1(n5448), .A2(n6084), .ZN(n5847) );
  OAI21_X1 U6026 ( .B1(n5305), .B2(n4889), .A(n5847), .ZN(n6075) );
  NAND2_X1 U6027 ( .A1(n6066), .A2(REIP_REG_5__SCAN_IN), .ZN(n6059) );
  INV_X1 U6028 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6536) );
  AOI22_X1 U6029 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6075), .B1(n6059), .B2(n6536), .ZN(n4887) );
  NAND2_X1 U6030 ( .A1(n4872), .A2(n4873), .ZN(n6494) );
  NAND2_X1 U6031 ( .A1(n6152), .A2(n6494), .ZN(n4876) );
  INV_X1 U6032 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5478) );
  INV_X1 U6033 ( .A(n4873), .ZN(n4878) );
  NAND3_X1 U6034 ( .A1(n4874), .A2(n5478), .A3(n4878), .ZN(n4875) );
  NAND2_X1 U6035 ( .A1(n4876), .A2(n4875), .ZN(n4877) );
  NAND2_X1 U6036 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4878), .ZN(n4879) );
  NOR2_X1 U6037 ( .A1(n4880), .A2(n4879), .ZN(n4881) );
  INV_X1 U6038 ( .A(n4882), .ZN(n6310) );
  AOI22_X1 U6039 ( .A1(n6090), .A2(n6310), .B1(n6053), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U6040 ( .A1(n6084), .A2(n4883), .ZN(n6055) );
  OAI211_X1 U6041 ( .C1(n6080), .C2(n4885), .A(n4884), .B(n6055), .ZN(n4886)
         );
  AOI211_X1 U6042 ( .C1(n4919), .C2(n6072), .A(n4887), .B(n4886), .ZN(n4888)
         );
  OAI21_X1 U6043 ( .B1(n5872), .B2(n4916), .A(n4888), .ZN(U2821) );
  INV_X1 U6044 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6541) );
  NAND2_X1 U6045 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n6057) );
  NOR3_X1 U6046 ( .A1(n6541), .A2(n4889), .A3(n6057), .ZN(n5269) );
  NAND2_X1 U6047 ( .A1(n5269), .A2(n6084), .ZN(n5197) );
  AND2_X1 U6048 ( .A1(n5847), .A2(n5197), .ZN(n6046) );
  OAI21_X1 U6049 ( .B1(n6057), .B2(n6059), .A(n6541), .ZN(n4890) );
  AOI22_X1 U6050 ( .A1(n4904), .A2(n6072), .B1(n6046), .B2(n4890), .ZN(n4899)
         );
  INV_X1 U6051 ( .A(n6051), .ZN(n4892) );
  OAI21_X1 U6052 ( .B1(n6052), .B2(n4892), .A(n4891), .ZN(n4893) );
  INV_X1 U6053 ( .A(n4893), .ZN(n4894) );
  OR2_X1 U6054 ( .A1(n4894), .A2(n5131), .ZN(n4912) );
  INV_X1 U6055 ( .A(n4912), .ZN(n6292) );
  NAND2_X1 U6056 ( .A1(n6090), .A2(n6292), .ZN(n4895) );
  OAI211_X1 U6057 ( .C1(n4896), .C2(n6093), .A(n4895), .B(n6055), .ZN(n4897)
         );
  AOI21_X1 U6058 ( .B1(EBX_REG_8__SCAN_IN), .B2(n6091), .A(n4897), .ZN(n4898)
         );
  OAI211_X1 U6059 ( .C1(n5872), .C2(n4910), .A(n4899), .B(n4898), .ZN(U2819)
         );
  OAI21_X1 U6060 ( .B1(n4903), .B2(n4902), .A(n4901), .ZN(n6293) );
  INV_X1 U6061 ( .A(n4904), .ZN(n4906) );
  NAND2_X1 U6062 ( .A1(n6338), .A2(REIP_REG_8__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U6063 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4905)
         );
  OAI211_X1 U6064 ( .C1(n6264), .C2(n4906), .A(n6290), .B(n4905), .ZN(n4907)
         );
  AOI21_X1 U6065 ( .B1(n4908), .B2(n6258), .A(n4907), .ZN(n4909) );
  OAI21_X1 U6066 ( .B1(n6293), .B2(n6273), .A(n4909), .ZN(U2978) );
  INV_X1 U6067 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4911) );
  OAI222_X1 U6068 ( .A1(n4912), .A2(n5885), .B1(n6118), .B2(n4911), .C1(n4910), 
        .C2(n5886), .ZN(U2851) );
  OAI21_X1 U6069 ( .B1(n4915), .B2(n4914), .A(n4913), .ZN(n6314) );
  NAND2_X1 U6070 ( .A1(n6338), .A2(REIP_REG_6__SCAN_IN), .ZN(n6308) );
  OAI21_X1 U6071 ( .B1(n5646), .B2(n3627), .A(n6308), .ZN(n4918) );
  NOR2_X1 U6072 ( .A1(n4916), .A2(n6271), .ZN(n4917) );
  AOI211_X1 U6073 ( .C1(n5649), .C2(n4919), .A(n4918), .B(n4917), .ZN(n4920)
         );
  OAI21_X1 U6074 ( .B1(n6273), .B2(n6314), .A(n4920), .ZN(U2980) );
  INV_X1 U6075 ( .A(n5359), .ZN(n4921) );
  OAI21_X1 U6076 ( .B1(n4922), .B2(n4921), .A(n5872), .ZN(n6100) );
  INV_X1 U6077 ( .A(n6100), .ZN(n4956) );
  INV_X1 U6078 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4929) );
  NAND2_X1 U6079 ( .A1(n5359), .A2(n4923), .ZN(n6092) );
  OAI22_X1 U6080 ( .A1(n6079), .A2(n4924), .B1(n5795), .B2(n6092), .ZN(n4928)
         );
  NAND2_X1 U6081 ( .A1(n6091), .A2(EBX_REG_1__SCAN_IN), .ZN(n4926) );
  AOI22_X1 U6082 ( .A1(n6053), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5305), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4925) );
  OAI211_X1 U6083 ( .C1(REIP_REG_1__SCAN_IN), .C2(n5448), .A(n4926), .B(n4925), 
        .ZN(n4927) );
  AOI211_X1 U6084 ( .C1(n6072), .C2(n4929), .A(n4928), .B(n4927), .ZN(n4930)
         );
  OAI21_X1 U6085 ( .B1(n4956), .B2(n6268), .A(n4930), .ZN(U2826) );
  NAND2_X1 U6086 ( .A1(n4932), .A2(n4931), .ZN(n4933) );
  NAND2_X1 U6087 ( .A1(n5219), .A2(n4933), .ZN(n5114) );
  AOI22_X1 U6088 ( .A1(n5538), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6125), .ZN(n4934) );
  OAI21_X1 U6089 ( .B1(n5114), .B2(n5890), .A(n4934), .ZN(U2882) );
  INV_X1 U6090 ( .A(n4935), .ZN(n5130) );
  XNOR2_X1 U6091 ( .A(n5131), .B(n5130), .ZN(n4997) );
  OAI22_X1 U6092 ( .A1(n5885), .A2(n4997), .B1(n6671), .B2(n6118), .ZN(n4936)
         );
  INV_X1 U6093 ( .A(n4936), .ZN(n4937) );
  OAI21_X1 U6094 ( .B1(n5114), .B2(n5886), .A(n4937), .ZN(U2850) );
  NOR2_X1 U6095 ( .A1(n6080), .A2(n4084), .ZN(n4940) );
  OAI22_X1 U6096 ( .A1(n6079), .A2(n6357), .B1(n4938), .B2(n6092), .ZN(n4939)
         );
  AOI211_X1 U6097 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5847), .A(n4940), .B(n4939), 
        .ZN(n4942) );
  OAI21_X1 U6098 ( .B1(n6072), .B2(n6053), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4941) );
  OAI211_X1 U6099 ( .C1(n4956), .C2(n6270), .A(n4942), .B(n4941), .ZN(U2827)
         );
  INV_X1 U6100 ( .A(n4946), .ZN(n4943) );
  OAI21_X1 U6101 ( .B1(n5448), .B2(n4943), .A(n6084), .ZN(n6086) );
  NOR2_X1 U6102 ( .A1(n6092), .A2(n5978), .ZN(n4944) );
  AOI211_X1 U6103 ( .C1(n6053), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6070), 
        .B(n4944), .ZN(n4949) );
  INV_X1 U6104 ( .A(n4945), .ZN(n6321) );
  NOR3_X1 U6105 ( .A1(n5448), .A2(REIP_REG_4__SCAN_IN), .A3(n4946), .ZN(n4947)
         );
  AOI21_X1 U6106 ( .B1(n6321), .B2(n6090), .A(n4947), .ZN(n4948) );
  OAI211_X1 U6107 ( .C1(n4950), .C2(n6080), .A(n4949), .B(n4948), .ZN(n4951)
         );
  AOI21_X1 U6108 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6086), .A(n4951), .ZN(n4954)
         );
  NAND2_X1 U6109 ( .A1(n6072), .A2(n4952), .ZN(n4953) );
  OAI211_X1 U6110 ( .C1(n4956), .C2(n4955), .A(n4954), .B(n4953), .ZN(U2823)
         );
  NAND2_X1 U6111 ( .A1(n4966), .A2(n6465), .ZN(n4957) );
  AOI21_X1 U6112 ( .B1(n4957), .B2(STATEBS16_REG_SCAN_IN), .A(n5799), .ZN(
        n4964) );
  NOR2_X1 U6113 ( .A1(n4958), .A2(n6768), .ZN(n4959) );
  AOI22_X1 U6114 ( .A1(n4964), .A2(n4961), .B1(n5141), .B2(n4959), .ZN(n4996)
         );
  NOR2_X1 U6115 ( .A1(n5054), .A2(n4960), .ZN(n5139) );
  INV_X1 U6116 ( .A(n4961), .ZN(n4963) );
  OR2_X1 U6117 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4962), .ZN(n4991)
         );
  AOI22_X1 U6118 ( .A1(n4964), .A2(n4963), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4991), .ZN(n4965) );
  OAI211_X1 U6119 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n5007), .A(n5139), .B(n4965), .ZN(n4990) );
  NAND2_X1 U6120 ( .A1(n4990), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4969)
         );
  OAI22_X1 U6121 ( .A1(n6465), .A2(n6794), .B1(n4991), .B2(n6789), .ZN(n4967)
         );
  AOI21_X1 U6122 ( .B1(n4993), .B2(n6396), .A(n4967), .ZN(n4968) );
  OAI211_X1 U6123 ( .C1(n4996), .C2(n5070), .A(n4969), .B(n4968), .ZN(U3102)
         );
  NAND2_X1 U6124 ( .A1(n4990), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4972)
         );
  OAI22_X1 U6125 ( .A1(n6465), .A2(n6412), .B1(n4991), .B2(n6411), .ZN(n4970)
         );
  AOI21_X1 U6126 ( .B1(n4993), .B2(n6402), .A(n4970), .ZN(n4971) );
  OAI211_X1 U6127 ( .C1(n4996), .C2(n5074), .A(n4972), .B(n4971), .ZN(U3103)
         );
  NAND2_X1 U6128 ( .A1(n4990), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4975)
         );
  OAI22_X1 U6129 ( .A1(n6465), .A2(n6407), .B1(n6406), .B2(n4991), .ZN(n4973)
         );
  AOI21_X1 U6130 ( .B1(n4993), .B2(n6389), .A(n4973), .ZN(n4974) );
  OAI211_X1 U6131 ( .C1(n4996), .C2(n5097), .A(n4975), .B(n4974), .ZN(U3100)
         );
  NAND2_X1 U6132 ( .A1(n4990), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4980)
         );
  OAI22_X1 U6133 ( .A1(n6465), .A2(n4976), .B1(n4991), .B2(n5177), .ZN(n4977)
         );
  AOI21_X1 U6134 ( .B1(n4993), .B2(n4978), .A(n4977), .ZN(n4979) );
  OAI211_X1 U6135 ( .C1(n4996), .C2(n5174), .A(n4980), .B(n4979), .ZN(U3107)
         );
  NAND2_X1 U6136 ( .A1(n4990), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4983)
         );
  OAI22_X1 U6137 ( .A1(n6465), .A2(n5157), .B1(n4991), .B2(n5156), .ZN(n4981)
         );
  AOI21_X1 U6138 ( .B1(n4993), .B2(n5101), .A(n4981), .ZN(n4982) );
  OAI211_X1 U6139 ( .C1(n4996), .C2(n5104), .A(n4983), .B(n4982), .ZN(U3105)
         );
  NAND2_X1 U6140 ( .A1(n4990), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4986)
         );
  OAI22_X1 U6141 ( .A1(n6465), .A2(n6418), .B1(n4991), .B2(n6416), .ZN(n4984)
         );
  AOI21_X1 U6142 ( .B1(n4993), .B2(n5086), .A(n4984), .ZN(n4985) );
  OAI211_X1 U6143 ( .C1(n4996), .C2(n5089), .A(n4986), .B(n4985), .ZN(U3104)
         );
  NAND2_X1 U6144 ( .A1(n4990), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4989)
         );
  OAI22_X1 U6145 ( .A1(n6465), .A2(n5165), .B1(n4991), .B2(n5164), .ZN(n4987)
         );
  AOI21_X1 U6146 ( .B1(n4993), .B2(n5081), .A(n4987), .ZN(n4988) );
  OAI211_X1 U6147 ( .C1(n4996), .C2(n5084), .A(n4989), .B(n4988), .ZN(U3106)
         );
  NAND2_X1 U6148 ( .A1(n4990), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4995)
         );
  OAI22_X1 U6149 ( .A1(n6465), .A2(n6395), .B1(n4991), .B2(n5146), .ZN(n4992)
         );
  AOI21_X1 U6150 ( .B1(n4993), .B2(n6392), .A(n4992), .ZN(n4994) );
  OAI211_X1 U6151 ( .C1(n4996), .C2(n5093), .A(n4995), .B(n4994), .ZN(U3101)
         );
  NOR3_X1 U6152 ( .A1(n6541), .A2(n6057), .A3(n6059), .ZN(n6026) );
  INV_X1 U6153 ( .A(n6026), .ZN(n6042) );
  NOR2_X1 U6154 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6042), .ZN(n6045) );
  INV_X1 U6155 ( .A(n6045), .ZN(n5003) );
  INV_X1 U6156 ( .A(n5110), .ZN(n5001) );
  AOI21_X1 U6157 ( .B1(n6053), .B2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6070), 
        .ZN(n4999) );
  INV_X1 U6158 ( .A(n4997), .ZN(n6284) );
  AOI22_X1 U6159 ( .A1(n6046), .A2(REIP_REG_9__SCAN_IN), .B1(n6090), .B2(n6284), .ZN(n4998) );
  OAI211_X1 U6160 ( .C1(n6671), .C2(n6080), .A(n4999), .B(n4998), .ZN(n5000)
         );
  AOI21_X1 U6161 ( .B1(n6072), .B2(n5001), .A(n5000), .ZN(n5002) );
  OAI211_X1 U6162 ( .C1(n5114), .C2(n5872), .A(n5003), .B(n5002), .ZN(U2818)
         );
  INV_X1 U6163 ( .A(n5009), .ZN(n5004) );
  INV_X1 U6164 ( .A(n5136), .ZN(n5061) );
  AOI21_X1 U6165 ( .B1(n5004), .B2(n6612), .A(n5061), .ZN(n5011) );
  NOR2_X1 U6166 ( .A1(n5005), .A2(n5012), .ZN(n5010) );
  AOI21_X1 U6167 ( .B1(n5006), .B2(n2985), .A(n5010), .ZN(n5014) );
  OAI22_X1 U6168 ( .A1(n5011), .A2(n5014), .B1(n5012), .B2(n5007), .ZN(n5045)
         );
  NAND2_X1 U6169 ( .A1(n5045), .A2(n6784), .ZN(n5020) );
  INV_X1 U6170 ( .A(n5010), .ZN(n5048) );
  INV_X1 U6171 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5017) );
  INV_X1 U6172 ( .A(n5011), .ZN(n5013) );
  AOI22_X1 U6173 ( .A1(n5014), .A2(n5013), .B1(n5012), .B2(n5799), .ZN(n5015)
         );
  OAI22_X1 U6174 ( .A1(n6789), .A2(n5048), .B1(n5017), .B2(n5046), .ZN(n5018)
         );
  AOI21_X1 U6175 ( .B1(n5137), .B2(n6441), .A(n5018), .ZN(n5019) );
  OAI211_X1 U6176 ( .C1(n5052), .C2(n6786), .A(n5020), .B(n5019), .ZN(U3030)
         );
  NAND2_X1 U6177 ( .A1(n5045), .A2(n6382), .ZN(n5024) );
  INV_X1 U6178 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5021) );
  OAI22_X1 U6179 ( .A1(n5164), .A2(n5048), .B1(n5021), .B2(n5046), .ZN(n5022)
         );
  AOI21_X1 U6180 ( .B1(n5137), .B2(n6379), .A(n5022), .ZN(n5023) );
  OAI211_X1 U6181 ( .C1(n5052), .C2(n6386), .A(n5024), .B(n5023), .ZN(U3034)
         );
  NAND2_X1 U6182 ( .A1(n5045), .A2(n6446), .ZN(n5028) );
  INV_X1 U6183 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5025) );
  OAI22_X1 U6184 ( .A1(n6411), .A2(n5048), .B1(n5025), .B2(n5046), .ZN(n5026)
         );
  AOI21_X1 U6185 ( .B1(n5137), .B2(n6445), .A(n5026), .ZN(n5027) );
  OAI211_X1 U6186 ( .C1(n5052), .C2(n6449), .A(n5028), .B(n5027), .ZN(U3031)
         );
  NAND2_X1 U6187 ( .A1(n5045), .A2(n6436), .ZN(n5032) );
  INV_X1 U6188 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5029) );
  OAI22_X1 U6189 ( .A1(n5146), .A2(n5048), .B1(n5029), .B2(n5046), .ZN(n5030)
         );
  AOI21_X1 U6190 ( .B1(n5137), .B2(n6435), .A(n5030), .ZN(n5031) );
  OAI211_X1 U6191 ( .C1(n5052), .C2(n6439), .A(n5032), .B(n5031), .ZN(U3029)
         );
  NAND2_X1 U6192 ( .A1(n5045), .A2(n6452), .ZN(n5036) );
  INV_X1 U6193 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5033) );
  OAI22_X1 U6194 ( .A1(n5156), .A2(n5048), .B1(n5033), .B2(n5046), .ZN(n5034)
         );
  AOI21_X1 U6195 ( .B1(n5137), .B2(n6451), .A(n5034), .ZN(n5035) );
  OAI211_X1 U6196 ( .C1(n5052), .C2(n6455), .A(n5036), .B(n5035), .ZN(U3033)
         );
  NAND2_X1 U6197 ( .A1(n5045), .A2(n6422), .ZN(n5040) );
  INV_X1 U6198 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5037) );
  OAI22_X1 U6199 ( .A1(n6416), .A2(n5048), .B1(n5037), .B2(n5046), .ZN(n5038)
         );
  AOI21_X1 U6200 ( .B1(n5137), .B2(n6372), .A(n5038), .ZN(n5039) );
  OAI211_X1 U6201 ( .C1(n5052), .C2(n6427), .A(n5040), .B(n5039), .ZN(U3032)
         );
  NAND2_X1 U6202 ( .A1(n5045), .A2(n6430), .ZN(n5044) );
  INV_X1 U6203 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5041) );
  OAI22_X1 U6204 ( .A1(n6406), .A2(n5048), .B1(n5041), .B2(n5046), .ZN(n5042)
         );
  AOI21_X1 U6205 ( .B1(n5137), .B2(n6429), .A(n5042), .ZN(n5043) );
  OAI211_X1 U6206 ( .C1(n5052), .C2(n6433), .A(n5044), .B(n5043), .ZN(U3028)
         );
  NAND2_X1 U6207 ( .A1(n5045), .A2(n6461), .ZN(n5051) );
  INV_X1 U6208 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5047) );
  OAI22_X1 U6209 ( .A1(n5177), .A2(n5048), .B1(n5047), .B2(n5046), .ZN(n5049)
         );
  AOI21_X1 U6210 ( .B1(n5137), .B2(n6458), .A(n5049), .ZN(n5050) );
  OAI211_X1 U6211 ( .C1(n5052), .C2(n6466), .A(n5051), .B(n5050), .ZN(U3035)
         );
  NAND2_X1 U6212 ( .A1(n5053), .A2(n5058), .ZN(n5057) );
  NAND2_X1 U6213 ( .A1(n5055), .A2(n5054), .ZN(n5056) );
  INV_X1 U6214 ( .A(n6787), .ZN(n5076) );
  NOR3_X1 U6215 ( .A1(n6459), .A2(n5076), .A3(n5799), .ZN(n5062) );
  INV_X1 U6216 ( .A(n5058), .ZN(n5059) );
  OAI22_X1 U6217 ( .A1(n5062), .A2(n5061), .B1(n5060), .B2(n5059), .ZN(n5066)
         );
  OR2_X1 U6218 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5063), .ZN(n5099)
         );
  AOI21_X1 U6219 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5099), .A(n5142), .ZN(
        n5064) );
  NAND3_X1 U6220 ( .A1(n5066), .A2(n5065), .A3(n5064), .ZN(n5098) );
  NAND2_X1 U6221 ( .A1(n5098), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5069)
         );
  OAI22_X1 U6222 ( .A1(n6789), .A2(n5099), .B1(n6787), .B2(n6794), .ZN(n5067)
         );
  AOI21_X1 U6223 ( .B1(n6396), .B2(n6459), .A(n5067), .ZN(n5068) );
  OAI211_X1 U6224 ( .C1(n5105), .C2(n5070), .A(n5069), .B(n5068), .ZN(U3118)
         );
  NAND2_X1 U6225 ( .A1(n5098), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5073)
         );
  OAI22_X1 U6226 ( .A1(n6411), .A2(n5099), .B1(n6787), .B2(n6412), .ZN(n5071)
         );
  AOI21_X1 U6227 ( .B1(n6402), .B2(n6459), .A(n5071), .ZN(n5072) );
  OAI211_X1 U6228 ( .C1(n5105), .C2(n5074), .A(n5073), .B(n5072), .ZN(U3119)
         );
  INV_X1 U6229 ( .A(n6459), .ZN(n5079) );
  NAND2_X1 U6230 ( .A1(n5098), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5078)
         );
  OAI22_X1 U6231 ( .A1(n5177), .A2(n5099), .B1(n5105), .B2(n5174), .ZN(n5075)
         );
  AOI21_X1 U6232 ( .B1(n6458), .B2(n5076), .A(n5075), .ZN(n5077) );
  OAI211_X1 U6233 ( .C1(n5079), .C2(n6466), .A(n5078), .B(n5077), .ZN(U3123)
         );
  NAND2_X1 U6234 ( .A1(n5098), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5083)
         );
  OAI22_X1 U6235 ( .A1(n5164), .A2(n5099), .B1(n6787), .B2(n5165), .ZN(n5080)
         );
  AOI21_X1 U6236 ( .B1(n5081), .B2(n6459), .A(n5080), .ZN(n5082) );
  OAI211_X1 U6237 ( .C1(n5105), .C2(n5084), .A(n5083), .B(n5082), .ZN(U3122)
         );
  NAND2_X1 U6238 ( .A1(n5098), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5088)
         );
  OAI22_X1 U6239 ( .A1(n6416), .A2(n5099), .B1(n6787), .B2(n6418), .ZN(n5085)
         );
  AOI21_X1 U6240 ( .B1(n5086), .B2(n6459), .A(n5085), .ZN(n5087) );
  OAI211_X1 U6241 ( .C1(n5105), .C2(n5089), .A(n5088), .B(n5087), .ZN(U3120)
         );
  NAND2_X1 U6242 ( .A1(n5098), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5092)
         );
  OAI22_X1 U6243 ( .A1(n5146), .A2(n5099), .B1(n6787), .B2(n6395), .ZN(n5090)
         );
  AOI21_X1 U6244 ( .B1(n6392), .B2(n6459), .A(n5090), .ZN(n5091) );
  OAI211_X1 U6245 ( .C1(n5105), .C2(n5093), .A(n5092), .B(n5091), .ZN(U3117)
         );
  NAND2_X1 U6246 ( .A1(n5098), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5096)
         );
  OAI22_X1 U6247 ( .A1(n6406), .A2(n5099), .B1(n6787), .B2(n6407), .ZN(n5094)
         );
  AOI21_X1 U6248 ( .B1(n6389), .B2(n6459), .A(n5094), .ZN(n5095) );
  OAI211_X1 U6249 ( .C1(n5105), .C2(n5097), .A(n5096), .B(n5095), .ZN(U3116)
         );
  NAND2_X1 U6250 ( .A1(n5098), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5103)
         );
  OAI22_X1 U6251 ( .A1(n5156), .A2(n5099), .B1(n6787), .B2(n5157), .ZN(n5100)
         );
  AOI21_X1 U6252 ( .B1(n5101), .B2(n6459), .A(n5100), .ZN(n5102) );
  OAI211_X1 U6253 ( .C1(n5105), .C2(n5104), .A(n5103), .B(n5102), .ZN(U3121)
         );
  NAND2_X1 U6254 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  XNOR2_X1 U6255 ( .A(n5106), .B(n5109), .ZN(n6286) );
  NAND2_X1 U6256 ( .A1(n6286), .A2(n6257), .ZN(n5113) );
  AND2_X1 U6257 ( .A1(n6338), .A2(REIP_REG_9__SCAN_IN), .ZN(n6283) );
  NOR2_X1 U6258 ( .A1(n6264), .A2(n5110), .ZN(n5111) );
  AOI211_X1 U6259 ( .C1(n6276), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6283), 
        .B(n5111), .ZN(n5112) );
  OAI211_X1 U6260 ( .C1(n6271), .C2(n5114), .A(n5113), .B(n5112), .ZN(U2977)
         );
  NAND2_X1 U6261 ( .A1(n5207), .A2(n5115), .ZN(n5117) );
  XOR2_X1 U6262 ( .A(n5117), .B(n5116), .Z(n5226) );
  INV_X1 U6263 ( .A(n5118), .ZN(n5120) );
  AND2_X1 U6264 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  AOI221_X1 U6265 ( .B1(n6341), .B2(n5125), .C1(n5123), .C2(n5122), .A(n5121), 
        .ZN(n6306) );
  OAI21_X1 U6266 ( .B1(n5124), .B2(n6294), .A(n6306), .ZN(n6285) );
  AOI21_X1 U6267 ( .B1(n6342), .B2(n6346), .A(n6341), .ZN(n6331) );
  NOR2_X1 U6268 ( .A1(n6331), .A2(n5125), .ZN(n6301) );
  NAND2_X1 U6269 ( .A1(n6294), .A2(n6301), .ZN(n6289) );
  AOI221_X1 U6270 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5126), .C2(n3494), .A(n6289), 
        .ZN(n5127) );
  AOI21_X1 U6271 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6285), .A(n5127), 
        .ZN(n5134) );
  INV_X1 U6272 ( .A(n5128), .ZN(n5129) );
  AOI21_X1 U6273 ( .B1(n5131), .B2(n5130), .A(n5129), .ZN(n5132) );
  AND2_X1 U6274 ( .A1(n6338), .A2(REIP_REG_10__SCAN_IN), .ZN(n5223) );
  AOI21_X1 U6275 ( .B1(n6340), .B2(n3015), .A(n5223), .ZN(n5133) );
  OAI211_X1 U6276 ( .C1(n5226), .C2(n6313), .A(n5134), .B(n5133), .ZN(U3008)
         );
  NOR2_X1 U6277 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5135), .ZN(n5145)
         );
  OAI21_X1 U6278 ( .B1(n5137), .B2(n5179), .A(n5136), .ZN(n5138) );
  NAND2_X1 U6279 ( .A1(n5138), .A2(n5144), .ZN(n5140) );
  OAI221_X1 U6280 ( .B1(n5145), .B2(n6589), .C1(n5145), .C2(n5140), .A(n5139), 
        .ZN(n5172) );
  NAND2_X1 U6281 ( .A1(n5172), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5149) );
  NAND3_X1 U6282 ( .A1(n5142), .A2(n5141), .A3(n6768), .ZN(n5143) );
  OAI21_X1 U6283 ( .B1(n5144), .B2(n5799), .A(n5143), .ZN(n5173) );
  INV_X1 U6284 ( .A(n5145), .ZN(n5176) );
  OAI22_X1 U6285 ( .A1(n6387), .A2(n6395), .B1(n5146), .B2(n5176), .ZN(n5147)
         );
  AOI21_X1 U6286 ( .B1(n6436), .B2(n5173), .A(n5147), .ZN(n5148) );
  OAI211_X1 U6287 ( .C1(n5182), .C2(n6439), .A(n5149), .B(n5148), .ZN(U3037)
         );
  NAND2_X1 U6288 ( .A1(n5172), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5152) );
  OAI22_X1 U6289 ( .A1(n6387), .A2(n6407), .B1(n6406), .B2(n5176), .ZN(n5150)
         );
  AOI21_X1 U6290 ( .B1(n6430), .B2(n5173), .A(n5150), .ZN(n5151) );
  OAI211_X1 U6291 ( .C1(n6433), .C2(n5182), .A(n5152), .B(n5151), .ZN(U3036)
         );
  NAND2_X1 U6292 ( .A1(n5172), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5155) );
  OAI22_X1 U6293 ( .A1(n6387), .A2(n6794), .B1(n6789), .B2(n5176), .ZN(n5153)
         );
  AOI21_X1 U6294 ( .B1(n6784), .B2(n5173), .A(n5153), .ZN(n5154) );
  OAI211_X1 U6295 ( .C1(n5182), .C2(n6786), .A(n5155), .B(n5154), .ZN(U3038)
         );
  NAND2_X1 U6296 ( .A1(n5172), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5160) );
  OAI22_X1 U6297 ( .A1(n6387), .A2(n5157), .B1(n5156), .B2(n5176), .ZN(n5158)
         );
  AOI21_X1 U6298 ( .B1(n6452), .B2(n5173), .A(n5158), .ZN(n5159) );
  OAI211_X1 U6299 ( .C1(n5182), .C2(n6455), .A(n5160), .B(n5159), .ZN(U3041)
         );
  NAND2_X1 U6300 ( .A1(n5172), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5163) );
  OAI22_X1 U6301 ( .A1(n6387), .A2(n6418), .B1(n6416), .B2(n5176), .ZN(n5161)
         );
  AOI21_X1 U6302 ( .B1(n6422), .B2(n5173), .A(n5161), .ZN(n5162) );
  OAI211_X1 U6303 ( .C1(n5182), .C2(n6427), .A(n5163), .B(n5162), .ZN(U3040)
         );
  NAND2_X1 U6304 ( .A1(n5172), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5168) );
  OAI22_X1 U6305 ( .A1(n6387), .A2(n5165), .B1(n5164), .B2(n5176), .ZN(n5166)
         );
  AOI21_X1 U6306 ( .B1(n6382), .B2(n5173), .A(n5166), .ZN(n5167) );
  OAI211_X1 U6307 ( .C1(n5182), .C2(n6386), .A(n5168), .B(n5167), .ZN(U3042)
         );
  NAND2_X1 U6308 ( .A1(n5172), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5171) );
  OAI22_X1 U6309 ( .A1(n6387), .A2(n6412), .B1(n6411), .B2(n5176), .ZN(n5169)
         );
  AOI21_X1 U6310 ( .B1(n6446), .B2(n5173), .A(n5169), .ZN(n5170) );
  OAI211_X1 U6311 ( .C1(n5182), .C2(n6449), .A(n5171), .B(n5170), .ZN(U3039)
         );
  NAND2_X1 U6312 ( .A1(n5172), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5181) );
  INV_X1 U6313 ( .A(n5173), .ZN(n5175) );
  OAI22_X1 U6314 ( .A1(n5177), .A2(n5176), .B1(n5175), .B2(n5174), .ZN(n5178)
         );
  AOI21_X1 U6315 ( .B1(n5179), .B2(n6458), .A(n5178), .ZN(n5180) );
  OAI211_X1 U6316 ( .C1(n5182), .C2(n6466), .A(n5181), .B(n5180), .ZN(U3043)
         );
  INV_X1 U6317 ( .A(n5183), .ZN(n5187) );
  INV_X1 U6318 ( .A(n5184), .ZN(n5186) );
  INV_X1 U6319 ( .A(n5185), .ZN(n5229) );
  AOI21_X1 U6320 ( .B1(n5187), .B2(n5186), .A(n5229), .ZN(n5215) );
  OR2_X1 U6321 ( .A1(n5189), .A2(n5188), .ZN(n5190) );
  AND2_X1 U6322 ( .A1(n5235), .A2(n5190), .ZN(n6278) );
  INV_X1 U6323 ( .A(n6278), .ZN(n5192) );
  OAI22_X1 U6324 ( .A1(n5885), .A2(n5192), .B1(n5191), .B2(n6118), .ZN(n5193)
         );
  AOI21_X1 U6325 ( .B1(n5215), .B2(n6116), .A(n5193), .ZN(n5194) );
  INV_X1 U6326 ( .A(n5194), .ZN(U2848) );
  INV_X1 U6327 ( .A(n5215), .ZN(n5206) );
  INV_X1 U6328 ( .A(n5213), .ZN(n5201) );
  OAI21_X1 U6329 ( .B1(n6093), .B2(n5195), .A(n6055), .ZN(n5200) );
  INV_X1 U6330 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U6331 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5202) );
  NOR2_X1 U6332 ( .A1(n6546), .A2(n5202), .ZN(n6027) );
  INV_X1 U6333 ( .A(n6027), .ZN(n5196) );
  OAI21_X1 U6334 ( .B1(n5197), .B2(n5196), .A(n5847), .ZN(n6035) );
  AOI22_X1 U6335 ( .A1(n6091), .A2(EBX_REG_11__SCAN_IN), .B1(n6090), .B2(n6278), .ZN(n5198) );
  OAI21_X1 U6336 ( .B1(n6035), .B2(n6546), .A(n5198), .ZN(n5199) );
  AOI211_X1 U6337 ( .C1(n6072), .C2(n5201), .A(n5200), .B(n5199), .ZN(n5205)
         );
  NOR2_X1 U6338 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5202), .ZN(n5203) );
  NAND2_X1 U6339 ( .A1(n6026), .A2(n5203), .ZN(n5204) );
  OAI211_X1 U6340 ( .C1(n5206), .C2(n5872), .A(n5205), .B(n5204), .ZN(U2816)
         );
  INV_X1 U6341 ( .A(DATAI_11_), .ZN(n6656) );
  INV_X1 U6342 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6217) );
  OAI222_X1 U6343 ( .A1(n5206), .A2(n5890), .B1(n5543), .B2(n6656), .C1(n5544), 
        .C2(n6217), .ZN(U2880) );
  NAND2_X1 U6344 ( .A1(n5208), .A2(n5207), .ZN(n5211) );
  XNOR2_X1 U6345 ( .A(n3493), .B(n5209), .ZN(n5210) );
  XNOR2_X1 U6346 ( .A(n5211), .B(n5210), .ZN(n6279) );
  INV_X1 U6347 ( .A(n6279), .ZN(n5217) );
  AOI22_X1 U6348 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n6338), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n5212) );
  OAI21_X1 U6349 ( .B1(n5213), .B2(n6264), .A(n5212), .ZN(n5214) );
  AOI21_X1 U6350 ( .B1(n5215), .B2(n6258), .A(n5214), .ZN(n5216) );
  OAI21_X1 U6351 ( .B1(n5217), .B2(n6273), .A(n5216), .ZN(U2975) );
  AND2_X1 U6352 ( .A1(n5219), .A2(n5218), .ZN(n5220) );
  NOR2_X1 U6353 ( .A1(n5184), .A2(n5220), .ZN(n6112) );
  INV_X1 U6354 ( .A(n6112), .ZN(n5221) );
  INV_X1 U6355 ( .A(DATAI_10_), .ZN(n6750) );
  INV_X1 U6356 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6214) );
  OAI222_X1 U6357 ( .A1(n5221), .A2(n5890), .B1(n5543), .B2(n6750), .C1(n5544), 
        .C2(n6214), .ZN(U2881) );
  AND2_X1 U6358 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5222)
         );
  AOI211_X1 U6359 ( .C1(n5649), .C2(n6044), .A(n5223), .B(n5222), .ZN(n5225)
         );
  NAND2_X1 U6360 ( .A1(n6112), .A2(n6258), .ZN(n5224) );
  OAI211_X1 U6361 ( .C1(n5226), .C2(n6273), .A(n5225), .B(n5224), .ZN(U2976)
         );
  OAI21_X1 U6362 ( .B1(n5229), .B2(n3711), .A(n5228), .ZN(n6037) );
  INV_X1 U6363 ( .A(DATAI_12_), .ZN(n6668) );
  OAI222_X1 U6364 ( .A1(n6037), .A2(n5890), .B1(n5543), .B2(n6668), .C1(n5544), 
        .C2(n3696), .ZN(U2879) );
  XNOR2_X1 U6365 ( .A(n5230), .B(n5231), .ZN(n5243) );
  INV_X1 U6366 ( .A(n5954), .ZN(n6281) );
  OR2_X1 U6367 ( .A1(n5232), .A2(n6341), .ZN(n5762) );
  INV_X1 U6368 ( .A(n5762), .ZN(n5233) );
  AOI221_X1 U6369 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6281), .C1(
        n5233), .C2(n6281), .A(n5237), .ZN(n5241) );
  NAND2_X1 U6370 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  NAND2_X1 U6371 ( .A1(n5252), .A2(n5236), .ZN(n6033) );
  INV_X1 U6372 ( .A(n6282), .ZN(n5958) );
  NAND3_X1 U6373 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5237), .A3(n5958), .ZN(n5239) );
  NAND2_X1 U6374 ( .A1(n6338), .A2(REIP_REG_12__SCAN_IN), .ZN(n5238) );
  OAI211_X1 U6375 ( .C1(n6358), .C2(n6033), .A(n5239), .B(n5238), .ZN(n5240)
         );
  AOI211_X1 U6376 ( .C1(n5243), .C2(n6354), .A(n5241), .B(n5240), .ZN(n5242)
         );
  INV_X1 U6377 ( .A(n5242), .ZN(U3006) );
  NAND2_X1 U6378 ( .A1(n5243), .A2(n6257), .ZN(n5248) );
  INV_X1 U6379 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5245) );
  INV_X1 U6380 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5244) );
  OAI22_X1 U6381 ( .A1(n5646), .A2(n5245), .B1(n5966), .B2(n5244), .ZN(n5246)
         );
  AOI21_X1 U6382 ( .B1(n5649), .B2(n6038), .A(n5246), .ZN(n5247) );
  OAI211_X1 U6383 ( .C1(n6271), .C2(n6037), .A(n5248), .B(n5247), .ZN(U2974)
         );
  XOR2_X1 U6384 ( .A(n5250), .B(n5249), .Z(n6030) );
  AND2_X1 U6385 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  OR2_X1 U6386 ( .A1(n5266), .A2(n5253), .ZN(n6023) );
  OAI22_X1 U6387 ( .A1(n5885), .A2(n6023), .B1(n6752), .B2(n6118), .ZN(n5254)
         );
  AOI21_X1 U6388 ( .B1(n6030), .B2(n6116), .A(n5254), .ZN(n5255) );
  INV_X1 U6389 ( .A(n5255), .ZN(U2846) );
  OAI21_X1 U6390 ( .B1(n5258), .B2(n5257), .A(n5256), .ZN(n5259) );
  INV_X1 U6391 ( .A(n5259), .ZN(n5967) );
  AOI22_X1 U6392 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n6338), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n5260) );
  OAI21_X1 U6393 ( .B1(n6024), .B2(n6264), .A(n5260), .ZN(n5261) );
  AOI21_X1 U6394 ( .B1(n6030), .B2(n6258), .A(n5261), .ZN(n5262) );
  OAI21_X1 U6395 ( .B1(n5967), .B2(n6273), .A(n5262), .ZN(U2973) );
  NAND2_X1 U6396 ( .A1(n5458), .A2(n5457), .ZN(n5536) );
  OAI21_X1 U6397 ( .B1(n5458), .B2(n5457), .A(n5536), .ZN(n5661) );
  AOI22_X1 U6398 ( .A1(n5538), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6125), .ZN(n5264) );
  OAI21_X1 U6399 ( .B1(n5661), .B2(n5890), .A(n5264), .ZN(U2877) );
  INV_X1 U6400 ( .A(n5663), .ZN(n5276) );
  NOR2_X1 U6401 ( .A1(n5266), .A2(n5265), .ZN(n5267) );
  OR2_X1 U6402 ( .A1(n5786), .A2(n5267), .ZN(n5960) );
  AOI21_X1 U6403 ( .B1(n6053), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6070), 
        .ZN(n5268) );
  OAI21_X1 U6404 ( .B1(n6079), .B2(n5960), .A(n5268), .ZN(n5275) );
  NAND4_X1 U6405 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        n5269), .A4(n6027), .ZN(n5273) );
  INV_X1 U6406 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6728) );
  NOR2_X1 U6407 ( .A1(n6728), .A2(n5273), .ZN(n5469) );
  INV_X1 U6408 ( .A(n5469), .ZN(n5270) );
  NAND2_X1 U6409 ( .A1(n6095), .A2(n5270), .ZN(n5272) );
  NAND2_X1 U6410 ( .A1(n5272), .A2(n6084), .ZN(n6015) );
  AOI22_X1 U6411 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6091), .B1(
        REIP_REG_14__SCAN_IN), .B2(n6015), .ZN(n5271) );
  OAI21_X1 U6412 ( .B1(n5273), .B2(n5272), .A(n5271), .ZN(n5274) );
  AOI211_X1 U6413 ( .C1(n6072), .C2(n5276), .A(n5275), .B(n5274), .ZN(n5277)
         );
  OAI21_X1 U6414 ( .B1(n5661), .B2(n5872), .A(n5277), .ZN(U2813) );
  XNOR2_X1 U6415 ( .A(n5278), .B(n5321), .ZN(n5550) );
  NOR2_X1 U6416 ( .A1(n5281), .A2(n5280), .ZN(n5297) );
  AOI22_X1 U6417 ( .A1(n2975), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5282), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5289) );
  AOI22_X1 U6418 ( .A1(n5283), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n2997), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5288) );
  AOI22_X1 U6419 ( .A1(n3157), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n2984), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5287) );
  AOI22_X1 U6420 ( .A1(n5285), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n2987), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5286) );
  NAND4_X1 U6421 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n5286), .ZN(n5295)
         );
  AOI22_X1 U6422 ( .A1(n3265), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5293) );
  AOI22_X1 U6423 ( .A1(n2994), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5292) );
  AOI22_X1 U6424 ( .A1(n3296), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3992), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5291) );
  AOI22_X1 U6425 ( .A1(n2995), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5290) );
  NAND4_X1 U6426 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n5294)
         );
  NOR2_X1 U6427 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  XNOR2_X1 U6428 ( .A(n5297), .B(n5296), .ZN(n5299) );
  NAND2_X1 U6429 ( .A1(n5299), .A2(n5298), .ZN(n5302) );
  AOI21_X1 U6430 ( .B1(n5321), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n5300) );
  AOI21_X1 U6431 ( .B1(n5351), .B2(EAX_REG_30__SCAN_IN), .A(n5300), .ZN(n5301)
         );
  NAND2_X1 U6432 ( .A1(n5302), .A2(n5301), .ZN(n5303) );
  NAND2_X1 U6433 ( .A1(n5304), .A2(n5303), .ZN(n5352) );
  XOR2_X1 U6434 ( .A(n5352), .B(n5353), .Z(n5552) );
  INV_X1 U6435 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6563) );
  INV_X1 U6436 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6705) );
  NAND4_X1 U6437 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5469), .ZN(n5447) );
  NOR2_X1 U6438 ( .A1(n6705), .A2(n5447), .ZN(n5432) );
  NAND3_X1 U6439 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        n5432), .ZN(n5310) );
  OR2_X1 U6440 ( .A1(n5310), .A2(n5305), .ZN(n5846) );
  NAND2_X1 U6441 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5848) );
  NOR3_X1 U6442 ( .A1(n6563), .A2(n5846), .A3(n5848), .ZN(n5405) );
  INV_X1 U6443 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6565) );
  INV_X1 U6444 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6569) );
  INV_X1 U6445 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5825) );
  NOR3_X1 U6446 ( .A1(n6565), .A2(n6569), .A3(n5825), .ZN(n5306) );
  NAND2_X1 U6447 ( .A1(n5405), .A2(n5306), .ZN(n5307) );
  AND2_X1 U6448 ( .A1(n5307), .A2(n5847), .ZN(n5819) );
  NAND2_X1 U6449 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5311) );
  INV_X1 U6450 ( .A(n5311), .ZN(n5308) );
  NOR2_X1 U6451 ( .A1(n5448), .A2(n5308), .ZN(n5309) );
  NOR2_X1 U6452 ( .A1(n5819), .A2(n5309), .ZN(n5398) );
  NOR2_X1 U6453 ( .A1(n5448), .A2(n5310), .ZN(n5849) );
  NAND3_X1 U6454 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        n5849), .ZN(n5834) );
  NAND4_X1 U6455 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .A4(n5823), .ZN(n5806) );
  NOR2_X1 U6456 ( .A1(n5311), .A2(n5806), .ZN(n5358) );
  INV_X1 U6457 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6575) );
  NAND2_X1 U6458 ( .A1(n5358), .A2(n6575), .ZN(n5383) );
  NAND2_X1 U6459 ( .A1(n5398), .A2(n5383), .ZN(n5364) );
  INV_X1 U6460 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6573) );
  AND3_X1 U6461 ( .A1(n5358), .A2(REIP_REG_29__SCAN_IN), .A3(n6573), .ZN(n5365) );
  INV_X1 U6462 ( .A(n5395), .ZN(n5312) );
  NAND2_X1 U6463 ( .A1(n5318), .A2(n5312), .ZN(n5314) );
  INV_X1 U6464 ( .A(n5317), .ZN(n5313) );
  NAND3_X1 U6465 ( .A1(n5315), .A2(n5314), .A3(n5313), .ZN(n5320) );
  NAND2_X1 U6466 ( .A1(n5395), .A2(n2977), .ZN(n5316) );
  NAND3_X1 U6467 ( .A1(n5318), .A2(n5317), .A3(n5316), .ZN(n5319) );
  OAI22_X1 U6468 ( .A1(n5321), .A2(n6093), .B1(n5550), .B2(n6103), .ZN(n5322)
         );
  AOI21_X1 U6469 ( .B1(n6091), .B2(EBX_REG_30__SCAN_IN), .A(n5322), .ZN(n5323)
         );
  INV_X1 U6470 ( .A(n6597), .ZN(n5346) );
  NAND2_X1 U6471 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5333) );
  AOI22_X1 U6472 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4045), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5324), .ZN(n5338) );
  NOR2_X1 U6473 ( .A1(n5333), .A2(n5338), .ZN(n5326) );
  INV_X1 U6474 ( .A(n4500), .ZN(n5330) );
  NOR3_X1 U6475 ( .A1(n5330), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6497), 
        .ZN(n5325) );
  AOI211_X1 U6476 ( .C1(n5327), .C2(n5346), .A(n5326), .B(n5325), .ZN(n5332)
         );
  AOI22_X1 U6477 ( .A1(n6490), .A2(n6470), .B1(FLUSH_REG_SCAN_IN), .B2(n5328), 
        .ZN(n5977) );
  INV_X1 U6478 ( .A(n5329), .ZN(n6587) );
  NAND2_X1 U6479 ( .A1(n5977), .A2(n6587), .ZN(n6593) );
  INV_X1 U6480 ( .A(n6593), .ZN(n5348) );
  INV_X1 U6481 ( .A(n6497), .ZN(n5341) );
  AOI21_X1 U6482 ( .B1(n5330), .B2(n5341), .A(n5348), .ZN(n5331) );
  OAI22_X1 U6483 ( .A1(n5332), .A2(n5348), .B1(n5331), .B2(n3107), .ZN(U3459)
         );
  OAI21_X1 U6484 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6497), .A(n6593), 
        .ZN(n6594) );
  INV_X1 U6485 ( .A(n6594), .ZN(n5343) );
  INV_X1 U6486 ( .A(n5333), .ZN(n5339) );
  NOR3_X1 U6487 ( .A1(n5334), .A2(n4500), .A3(n4490), .ZN(n5335) );
  AOI21_X1 U6488 ( .B1(n6469), .B2(n3108), .A(n5335), .ZN(n5336) );
  OAI21_X1 U6489 ( .B1(n5795), .B2(n5337), .A(n5336), .ZN(n6473) );
  AOI222_X1 U6490 ( .A1(n5341), .A2(n5340), .B1(n5339), .B2(n5338), .C1(n6473), 
        .C2(n5346), .ZN(n5342) );
  OAI22_X1 U6491 ( .A1(n5343), .A2(n3108), .B1(n5348), .B2(n5342), .ZN(U3460)
         );
  NOR2_X1 U6492 ( .A1(n5344), .A2(n6497), .ZN(n5345) );
  AOI21_X1 U6493 ( .B1(n5347), .B2(n5346), .A(n5345), .ZN(n5349) );
  AOI22_X1 U6494 ( .A1(n6593), .A2(n5349), .B1(n5348), .B2(n3109), .ZN(U3456)
         );
  AOI22_X1 U6495 ( .A1(n5351), .A2(EAX_REG_31__SCAN_IN), .B1(n5350), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6496 ( .A1(n5544), .A2(n4303), .ZN(n5357) );
  AOI22_X1 U6497 ( .A1(n6122), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6125), .ZN(n5356) );
  OAI21_X1 U6498 ( .B1(n5374), .B2(n5357), .A(n5356), .ZN(U2860) );
  AND4_X1 U6499 ( .A1(n5358), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n6701), .ZN(n5363) );
  INV_X1 U6500 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5361) );
  NAND4_X1 U6501 ( .A1(n5359), .A2(n6152), .A3(EBX_REG_31__SCAN_IN), .A4(n6494), .ZN(n5360) );
  OAI21_X1 U6502 ( .B1(n6093), .B2(n5361), .A(n5360), .ZN(n5362) );
  AOI211_X1 U6503 ( .C1(n5477), .C2(n6090), .A(n5363), .B(n5362), .ZN(n5367)
         );
  OAI21_X1 U6504 ( .B1(n5365), .B2(n5364), .A(REIP_REG_31__SCAN_IN), .ZN(n5366) );
  OAI211_X1 U6505 ( .C1(n5374), .C2(n5872), .A(n5367), .B(n5366), .ZN(U2796)
         );
  NAND2_X1 U6506 ( .A1(n5368), .A2(n6257), .ZN(n5373) );
  NOR2_X1 U6507 ( .A1(n5369), .A2(n6264), .ZN(n5370) );
  AOI211_X1 U6508 ( .C1(n6276), .C2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5371), 
        .B(n5370), .ZN(n5372) );
  OAI211_X1 U6509 ( .C1(n5374), .C2(n6271), .A(n5373), .B(n5372), .ZN(U2955)
         );
  XNOR2_X1 U6510 ( .A(n5395), .B(n5375), .ZN(n5676) );
  INV_X1 U6511 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5387) );
  NOR2_X1 U6512 ( .A1(n6118), .A2(n5387), .ZN(n5376) );
  AOI21_X1 U6513 ( .B1(n5676), .B2(n6115), .A(n5376), .ZN(n5377) );
  OAI21_X1 U6514 ( .B1(n5380), .B2(n5886), .A(n5377), .ZN(U2830) );
  AOI22_X1 U6515 ( .A1(n6122), .A2(DATAI_29_), .B1(n6125), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6516 ( .A1(n6126), .A2(DATAI_13_), .ZN(n5378) );
  OAI211_X1 U6517 ( .C1(n5380), .C2(n5890), .A(n5379), .B(n5378), .ZN(U2862)
         );
  INV_X1 U6518 ( .A(n5380), .ZN(n5381) );
  NAND2_X1 U6519 ( .A1(n5381), .A2(n6064), .ZN(n5390) );
  NAND2_X1 U6520 ( .A1(n6072), .A2(n5382), .ZN(n5386) );
  INV_X1 U6521 ( .A(n5383), .ZN(n5384) );
  AOI21_X1 U6522 ( .B1(n6053), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5384), 
        .ZN(n5385) );
  OAI211_X1 U6523 ( .C1(n5387), .C2(n6080), .A(n5386), .B(n5385), .ZN(n5388)
         );
  AOI21_X1 U6524 ( .B1(n5676), .B2(n6090), .A(n5388), .ZN(n5389) );
  OAI211_X1 U6525 ( .C1(n5398), .C2(n6575), .A(n5390), .B(n5389), .ZN(U2798)
         );
  AOI21_X1 U6526 ( .B1(n5392), .B2(n5391), .A(n4029), .ZN(n5563) );
  INV_X1 U6527 ( .A(n5563), .ZN(n5525) );
  OR2_X1 U6528 ( .A1(n5700), .A2(n5393), .ZN(n5394) );
  NAND2_X1 U6529 ( .A1(n5395), .A2(n5394), .ZN(n5693) );
  INV_X1 U6530 ( .A(n5561), .ZN(n5396) );
  AOI22_X1 U6531 ( .A1(n6072), .A2(n5396), .B1(n6091), .B2(EBX_REG_28__SCAN_IN), .ZN(n5397) );
  OAI21_X1 U6532 ( .B1(n5693), .B2(n6079), .A(n5397), .ZN(n5401) );
  INV_X1 U6533 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5809) );
  NOR3_X1 U6534 ( .A1(REIP_REG_28__SCAN_IN), .A2(n5809), .A3(n5806), .ZN(n5400) );
  INV_X1 U6535 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6572) );
  INV_X1 U6536 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6741) );
  OAI22_X1 U6537 ( .A1(n5398), .A2(n6572), .B1(n6741), .B2(n6093), .ZN(n5399)
         );
  NOR3_X1 U6538 ( .A1(n5401), .A2(n5400), .A3(n5399), .ZN(n5402) );
  OAI21_X1 U6539 ( .B1(n5525), .B2(n5872), .A(n5402), .ZN(U2799) );
  INV_X1 U6540 ( .A(n5586), .ZN(n5403) );
  AOI21_X1 U6541 ( .B1(n5404), .B2(n5602), .A(n5403), .ZN(n5897) );
  INV_X1 U6542 ( .A(n5897), .ZN(n5413) );
  INV_X1 U6543 ( .A(n5847), .ZN(n6083) );
  NOR2_X1 U6544 ( .A1(n6083), .A2(n5405), .ZN(n5837) );
  OAI22_X1 U6545 ( .A1(n5489), .A2(n6080), .B1(n5406), .B2(n6093), .ZN(n5407)
         );
  AOI221_X1 U6546 ( .B1(n5837), .B2(REIP_REG_24__SCAN_IN), .C1(n5823), .C2(
        n6565), .A(n5407), .ZN(n5412) );
  NOR2_X1 U6547 ( .A1(n5735), .A2(n5408), .ZN(n5409) );
  OR2_X1 U6548 ( .A1(n5717), .A2(n5409), .ZN(n5490) );
  INV_X1 U6549 ( .A(n5490), .ZN(n5731) );
  INV_X1 U6550 ( .A(n5599), .ZN(n5410) );
  AOI22_X1 U6551 ( .A1(n5731), .A2(n6090), .B1(n5410), .B2(n6072), .ZN(n5411)
         );
  OAI211_X1 U6552 ( .C1(n5413), .C2(n5872), .A(n5412), .B(n5411), .ZN(U2803)
         );
  NOR2_X1 U6553 ( .A1(n5414), .A2(n5415), .ZN(n5416) );
  OR2_X1 U6554 ( .A1(n5494), .A2(n5416), .ZN(n5903) );
  NAND2_X1 U6555 ( .A1(n5847), .A2(n5846), .ZN(n5433) );
  INV_X1 U6556 ( .A(n5433), .ZN(n5424) );
  INV_X1 U6557 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6560) );
  INV_X1 U6558 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6675) );
  OAI22_X1 U6559 ( .A1(n6675), .A2(n6080), .B1(n5622), .B2(n6093), .ZN(n5420)
         );
  XNOR2_X1 U6560 ( .A(n5418), .B(n5417), .ZN(n5757) );
  NOR2_X1 U6561 ( .A1(n5757), .A2(n6079), .ZN(n5419) );
  AOI211_X1 U6562 ( .C1(n5849), .C2(n6560), .A(n5420), .B(n5419), .ZN(n5421)
         );
  OAI21_X1 U6563 ( .B1(n5422), .B2(n6103), .A(n5421), .ZN(n5423) );
  AOI21_X1 U6564 ( .B1(REIP_REG_21__SCAN_IN), .B2(n5424), .A(n5423), .ZN(n5425) );
  OAI21_X1 U6565 ( .B1(n5903), .B2(n5872), .A(n5425), .ZN(U2806) );
  NAND2_X1 U6566 ( .A1(n5458), .A2(n5426), .ZN(n5864) );
  AND2_X1 U6567 ( .A1(n5864), .A2(n5427), .ZN(n5428) );
  INV_X1 U6568 ( .A(n5629), .ZN(n5437) );
  INV_X1 U6569 ( .A(n5445), .ZN(n5429) );
  MUX2_X1 U6570 ( .A(n5429), .B(n5444), .S(n5870), .Z(n5431) );
  XNOR2_X1 U6571 ( .A(n5431), .B(n5430), .ZN(n5771) );
  INV_X1 U6572 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5502) );
  OAI22_X1 U6573 ( .A1(n5771), .A2(n6079), .B1(n5502), .B2(n6080), .ZN(n5436)
         );
  AND2_X1 U6574 ( .A1(n6095), .A2(n5432), .ZN(n5854) );
  AOI21_X1 U6575 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5854), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5434) );
  INV_X1 U6576 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6661) );
  OAI22_X1 U6577 ( .A1(n5434), .A2(n5433), .B1(n6661), .B2(n6093), .ZN(n5435)
         );
  AOI211_X1 U6578 ( .C1(n6072), .C2(n5437), .A(n5436), .B(n5435), .ZN(n5438)
         );
  OAI21_X1 U6579 ( .B1(n5633), .B2(n5872), .A(n5438), .ZN(U2807) );
  NAND2_X1 U6580 ( .A1(n5458), .A2(n5439), .ZN(n5509) );
  NAND2_X1 U6581 ( .A1(n5458), .A2(n5440), .ZN(n5862) );
  INV_X1 U6582 ( .A(n5862), .ZN(n5441) );
  INV_X1 U6583 ( .A(n6119), .ZN(n5455) );
  NOR2_X1 U6584 ( .A1(n5444), .A2(EBX_REG_18__SCAN_IN), .ZN(n5443) );
  AOI21_X1 U6585 ( .B1(n5445), .B2(n5444), .A(n5443), .ZN(n5866) );
  OR2_X1 U6586 ( .A1(n5513), .A2(n5866), .ZN(n5865) );
  NAND2_X1 U6587 ( .A1(n5513), .A2(n5866), .ZN(n5446) );
  NAND2_X1 U6588 ( .A1(n5865), .A2(n5446), .ZN(n5780) );
  OAI22_X1 U6589 ( .A1(n6080), .A2(n5503), .B1(n6079), .B2(n5780), .ZN(n5453)
         );
  INV_X1 U6590 ( .A(n5447), .ZN(n5449) );
  OAI21_X1 U6591 ( .B1(n5448), .B2(n5449), .A(n6084), .ZN(n6007) );
  NOR2_X1 U6592 ( .A1(n5448), .A2(REIP_REG_18__SCAN_IN), .ZN(n5855) );
  AOI22_X1 U6593 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6007), .B1(n5449), .B2(
        n5855), .ZN(n5450) );
  OAI211_X1 U6594 ( .C1(n6093), .C2(n5451), .A(n5450), .B(n6055), .ZN(n5452)
         );
  AOI211_X1 U6595 ( .C1(n6072), .C2(n5637), .A(n5453), .B(n5452), .ZN(n5454)
         );
  OAI21_X1 U6596 ( .B1(n5455), .B2(n5872), .A(n5454), .ZN(U2809) );
  AND2_X1 U6597 ( .A1(n5458), .A2(n5457), .ZN(n5460) );
  INV_X1 U6598 ( .A(n5462), .ZN(n5648) );
  INV_X1 U6599 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5468) );
  INV_X1 U6600 ( .A(n5785), .ZN(n5463) );
  NAND2_X1 U6601 ( .A1(n5786), .A2(n5463), .ZN(n5465) );
  NAND2_X1 U6602 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  AND2_X1 U6603 ( .A1(n5466), .A2(n5511), .ZN(n5944) );
  INV_X1 U6604 ( .A(n5944), .ZN(n5467) );
  OAI22_X1 U6605 ( .A1(n6080), .A2(n5468), .B1(n6079), .B2(n5467), .ZN(n5475)
         );
  INV_X1 U6606 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U6607 ( .A1(n6095), .A2(n5469), .ZN(n5470) );
  NOR2_X1 U6608 ( .A1(n6552), .A2(n5470), .ZN(n6005) );
  INV_X1 U6609 ( .A(n6005), .ZN(n5472) );
  NOR2_X1 U6610 ( .A1(n5470), .A2(REIP_REG_15__SCAN_IN), .ZN(n6016) );
  NOR2_X1 U6611 ( .A1(n6016), .A2(n6015), .ZN(n5471) );
  MUX2_X1 U6612 ( .A(n5472), .B(n5471), .S(REIP_REG_16__SCAN_IN), .Z(n5473) );
  OAI211_X1 U6613 ( .C1(n6093), .C2(n5645), .A(n5473), .B(n6055), .ZN(n5474)
         );
  AOI211_X1 U6614 ( .C1(n6072), .C2(n5648), .A(n5475), .B(n5474), .ZN(n5476)
         );
  OAI21_X1 U6615 ( .B1(n5652), .B2(n5872), .A(n5476), .ZN(U2811) );
  INV_X1 U6616 ( .A(n5477), .ZN(n5479) );
  OAI22_X1 U6617 ( .A1(n5479), .A2(n5885), .B1(n6118), .B2(n5478), .ZN(U2828)
         );
  INV_X1 U6618 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5480) );
  OAI222_X1 U6619 ( .A1(n5886), .A2(n5522), .B1(n5480), .B2(n6118), .C1(n5671), 
        .C2(n5885), .ZN(U2829) );
  OAI22_X1 U6620 ( .A1(n5693), .A2(n5885), .B1(n5481), .B2(n6118), .ZN(n5482)
         );
  AOI21_X1 U6621 ( .B1(n5563), .B2(n6116), .A(n5482), .ZN(n5483) );
  INV_X1 U6622 ( .A(n5483), .ZN(U2831) );
  INV_X1 U6623 ( .A(n5569), .ZN(n5484) );
  OAI21_X1 U6624 ( .B1(n5485), .B2(n5588), .A(n5484), .ZN(n5816) );
  NAND2_X1 U6625 ( .A1(n3004), .A2(n5486), .ZN(n5487) );
  NAND2_X1 U6626 ( .A1(n3002), .A2(n5487), .ZN(n5815) );
  INV_X1 U6627 ( .A(n5815), .ZN(n5708) );
  AOI22_X1 U6628 ( .A1(n5708), .A2(n6115), .B1(EBX_REG_26__SCAN_IN), .B2(n5517), .ZN(n5488) );
  OAI21_X1 U6629 ( .B1(n5816), .B2(n5886), .A(n5488), .ZN(U2833) );
  OAI22_X1 U6630 ( .A1(n5490), .A2(n5885), .B1(n5489), .B2(n6118), .ZN(n5491)
         );
  AOI21_X1 U6631 ( .B1(n5897), .B2(n6116), .A(n5491), .ZN(n5492) );
  INV_X1 U6632 ( .A(n5492), .ZN(U2835) );
  NOR2_X1 U6633 ( .A1(n5494), .A2(n5493), .ZN(n5495) );
  NAND2_X1 U6634 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  NAND2_X1 U6635 ( .A1(n5736), .A2(n5498), .ZN(n5842) );
  OAI22_X1 U6636 ( .A1(n5842), .A2(n5885), .B1(n5499), .B2(n6118), .ZN(n5500)
         );
  INV_X1 U6637 ( .A(n5500), .ZN(n5501) );
  OAI21_X1 U6638 ( .B1(n5843), .B2(n5886), .A(n5501), .ZN(U2837) );
  OAI222_X1 U6639 ( .A1(n5885), .A2(n5757), .B1(n6118), .B2(n6675), .C1(n5903), 
        .C2(n5886), .ZN(U2838) );
  OAI222_X1 U6640 ( .A1(n5885), .A2(n5771), .B1(n5502), .B2(n6118), .C1(n5633), 
        .C2(n5886), .ZN(U2839) );
  OAI22_X1 U6641 ( .A1(n5780), .A2(n5885), .B1(n5503), .B2(n6118), .ZN(n5504)
         );
  AOI21_X1 U6642 ( .B1(n6119), .B2(n6116), .A(n5504), .ZN(n5505) );
  INV_X1 U6643 ( .A(n5505), .ZN(U2841) );
  INV_X1 U6644 ( .A(n6124), .ZN(n5516) );
  NAND2_X1 U6645 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  AND2_X1 U6646 ( .A1(n5513), .A2(n5512), .ZN(n6011) );
  INV_X1 U6647 ( .A(n6011), .ZN(n5514) );
  OAI222_X1 U6648 ( .A1(n5516), .A2(n5886), .B1(n5515), .B2(n6118), .C1(n5885), 
        .C2(n5514), .ZN(U2842) );
  AOI22_X1 U6649 ( .A1(n5944), .A2(n6115), .B1(EBX_REG_16__SCAN_IN), .B2(n5517), .ZN(n5518) );
  OAI21_X1 U6650 ( .B1(n5652), .B2(n5886), .A(n5518), .ZN(U2843) );
  INV_X1 U6651 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5519) );
  OAI222_X1 U6652 ( .A1(n5661), .A2(n5886), .B1(n5519), .B2(n6118), .C1(n5885), 
        .C2(n5960), .ZN(U2845) );
  AOI22_X1 U6653 ( .A1(n6122), .A2(DATAI_30_), .B1(n6125), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U6654 ( .A1(n6126), .A2(DATAI_14_), .ZN(n5520) );
  OAI211_X1 U6655 ( .C1(n5522), .C2(n5890), .A(n5521), .B(n5520), .ZN(U2861)
         );
  AOI22_X1 U6656 ( .A1(n6122), .A2(DATAI_28_), .B1(n6125), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U6657 ( .A1(n6126), .A2(DATAI_12_), .ZN(n5523) );
  OAI211_X1 U6658 ( .C1(n5525), .C2(n5890), .A(n5524), .B(n5523), .ZN(U2863)
         );
  AOI22_X1 U6659 ( .A1(n6126), .A2(DATAI_10_), .B1(n6125), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6660 ( .A1(n6122), .A2(DATAI_26_), .ZN(n5526) );
  OAI211_X1 U6661 ( .C1(n5816), .C2(n5890), .A(n5527), .B(n5526), .ZN(U2865)
         );
  AOI22_X1 U6662 ( .A1(n6126), .A2(DATAI_6_), .B1(n6125), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U6663 ( .A1(n6122), .A2(DATAI_22_), .ZN(n5528) );
  OAI211_X1 U6664 ( .C1(n5843), .C2(n5890), .A(n5529), .B(n5528), .ZN(U2869)
         );
  AOI22_X1 U6665 ( .A1(n6122), .A2(DATAI_20_), .B1(n6125), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U6666 ( .A1(n6126), .A2(DATAI_4_), .ZN(n5530) );
  OAI211_X1 U6667 ( .C1(n5633), .C2(n5890), .A(n5531), .B(n5530), .ZN(U2871)
         );
  AOI22_X1 U6668 ( .A1(n6122), .A2(DATAI_16_), .B1(n6125), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U6669 ( .A1(n6126), .A2(DATAI_0_), .ZN(n5532) );
  OAI211_X1 U6670 ( .C1(n5652), .C2(n5890), .A(n5533), .B(n5532), .ZN(U2875)
         );
  INV_X1 U6671 ( .A(n5534), .ZN(n5535) );
  INV_X1 U6672 ( .A(n6105), .ZN(n5540) );
  AOI22_X1 U6673 ( .A1(n5538), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6125), .ZN(n5539) );
  OAI21_X1 U6674 ( .B1(n5540), .B2(n5890), .A(n5539), .ZN(U2876) );
  INV_X1 U6675 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6222) );
  INV_X1 U6676 ( .A(DATAI_13_), .ZN(n5542) );
  INV_X1 U6677 ( .A(n6030), .ZN(n5541) );
  OAI222_X1 U6678 ( .A1(n5544), .A2(n6222), .B1(n5543), .B2(n5542), .C1(n5890), 
        .C2(n5541), .ZN(U2878) );
  NAND2_X1 U6679 ( .A1(n5545), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5546) );
  OAI21_X1 U6680 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5547), .A(n5546), 
        .ZN(n5548) );
  XNOR2_X1 U6681 ( .A(n5548), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5675)
         );
  NAND2_X1 U6682 ( .A1(n6338), .A2(REIP_REG_30__SCAN_IN), .ZN(n5670) );
  NAND2_X1 U6683 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5549)
         );
  OAI211_X1 U6684 ( .C1(n5550), .C2(n6264), .A(n5670), .B(n5549), .ZN(n5551)
         );
  AOI21_X1 U6685 ( .B1(n5552), .B2(n6258), .A(n5551), .ZN(n5553) );
  OAI21_X1 U6686 ( .B1(n5675), .B2(n6273), .A(n5553), .ZN(U2956) );
  NAND3_X1 U6687 ( .A1(n5554), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n3493), .ZN(n5558) );
  INV_X1 U6688 ( .A(n5555), .ZN(n5583) );
  NOR2_X1 U6689 ( .A1(n5574), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5556)
         );
  NAND2_X1 U6690 ( .A1(n5583), .A2(n5556), .ZN(n5565) );
  AOI22_X1 U6691 ( .A1(n5558), .A2(n5565), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5557), .ZN(n5559) );
  XNOR2_X1 U6692 ( .A(n5559), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5697)
         );
  NAND2_X1 U6693 ( .A1(n6338), .A2(REIP_REG_28__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U6694 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5560)
         );
  OAI211_X1 U6695 ( .C1(n5561), .C2(n6264), .A(n5691), .B(n5560), .ZN(n5562)
         );
  AOI21_X1 U6696 ( .B1(n5563), .B2(n6258), .A(n5562), .ZN(n5564) );
  OAI21_X1 U6697 ( .B1(n6273), .B2(n5697), .A(n5564), .ZN(U2958) );
  NAND2_X1 U6698 ( .A1(n5566), .A2(n5565), .ZN(n5567) );
  XNOR2_X1 U6699 ( .A(n5567), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5707)
         );
  OR2_X1 U6700 ( .A1(n5569), .A2(n5568), .ZN(n5570) );
  NAND2_X1 U6701 ( .A1(n6338), .A2(REIP_REG_27__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6702 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5571)
         );
  OAI211_X1 U6703 ( .C1(n5813), .C2(n6264), .A(n5702), .B(n5571), .ZN(n5572)
         );
  AOI21_X1 U6704 ( .B1(n5891), .B2(n6258), .A(n5572), .ZN(n5573) );
  OAI21_X1 U6705 ( .B1(n5707), .B2(n6273), .A(n5573), .ZN(U2959) );
  INV_X1 U6706 ( .A(n5574), .ZN(n5576) );
  NOR2_X1 U6707 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  XNOR2_X1 U6708 ( .A(n3020), .B(n5577), .ZN(n5714) );
  NAND2_X1 U6709 ( .A1(n6338), .A2(REIP_REG_26__SCAN_IN), .ZN(n5710) );
  OAI21_X1 U6710 ( .B1(n5646), .B2(n5578), .A(n5710), .ZN(n5580) );
  NOR2_X1 U6711 ( .A1(n5816), .A2(n6271), .ZN(n5579) );
  AOI211_X1 U6712 ( .C1(n5814), .C2(n5649), .A(n5580), .B(n5579), .ZN(n5581)
         );
  OAI21_X1 U6713 ( .B1(n5714), .B2(n6273), .A(n5581), .ZN(U2960) );
  AOI21_X1 U6714 ( .B1(n3510), .B2(n5555), .A(n5584), .ZN(n5724) );
  AND2_X1 U6715 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  NOR2_X1 U6716 ( .A1(n5588), .A2(n5587), .ZN(n5894) );
  NAND2_X1 U6717 ( .A1(n6338), .A2(REIP_REG_25__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U6718 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5589)
         );
  OAI211_X1 U6719 ( .C1(n5824), .C2(n6264), .A(n5719), .B(n5589), .ZN(n5590)
         );
  AOI21_X1 U6720 ( .B1(n5894), .B2(n6258), .A(n5590), .ZN(n5591) );
  OAI21_X1 U6721 ( .B1(n5724), .B2(n6273), .A(n5591), .ZN(U2961) );
  XNOR2_X1 U6722 ( .A(n3493), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5911)
         );
  INV_X1 U6723 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5932) );
  INV_X1 U6724 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6659) );
  XNOR2_X1 U6725 ( .A(n3493), .B(n5746), .ZN(n5621) );
  INV_X1 U6726 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5744) );
  NAND3_X1 U6727 ( .A1(n3493), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5595) );
  XNOR2_X1 U6728 ( .A(n5597), .B(n5728), .ZN(n5733) );
  AND2_X1 U6729 ( .A1(n6338), .A2(REIP_REG_24__SCAN_IN), .ZN(n5730) );
  AOI21_X1 U6730 ( .B1(n6276), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5730), 
        .ZN(n5598) );
  OAI21_X1 U6731 ( .B1(n6264), .B2(n5599), .A(n5598), .ZN(n5600) );
  AOI21_X1 U6732 ( .B1(n5897), .B2(n6258), .A(n5600), .ZN(n5601) );
  OAI21_X1 U6733 ( .B1(n5733), .B2(n6273), .A(n5601), .ZN(U2962) );
  OAI21_X1 U6734 ( .B1(n5604), .B2(n5603), .A(n5602), .ZN(n5838) );
  INV_X1 U6735 ( .A(n3005), .ZN(n5609) );
  NOR2_X1 U6736 ( .A1(n5605), .A2(n5738), .ZN(n5606) );
  XNOR2_X1 U6737 ( .A(n5610), .B(n5744), .ZN(n5734) );
  NAND2_X1 U6738 ( .A1(n5734), .A2(n6257), .ZN(n5613) );
  AND2_X1 U6739 ( .A1(n6338), .A2(REIP_REG_23__SCAN_IN), .ZN(n5741) );
  NOR2_X1 U6740 ( .A1(n6264), .A2(n5841), .ZN(n5611) );
  AOI211_X1 U6741 ( .C1(PHYADDRPOINTER_REG_23__SCAN_IN), .C2(n6276), .A(n5741), 
        .B(n5611), .ZN(n5612) );
  OAI211_X1 U6742 ( .C1(n6271), .C2(n5838), .A(n5613), .B(n5612), .ZN(U2963)
         );
  XNOR2_X1 U6743 ( .A(n3493), .B(n6692), .ZN(n5614) );
  XNOR2_X1 U6744 ( .A(n5615), .B(n5614), .ZN(n5752) );
  NAND2_X1 U6745 ( .A1(n5752), .A2(n6257), .ZN(n5619) );
  NAND2_X1 U6746 ( .A1(n6338), .A2(REIP_REG_22__SCAN_IN), .ZN(n5748) );
  OAI21_X1 U6747 ( .B1(n5646), .B2(n5616), .A(n5748), .ZN(n5617) );
  AOI21_X1 U6748 ( .B1(n5649), .B2(n5845), .A(n5617), .ZN(n5618) );
  OAI211_X1 U6749 ( .C1(n6271), .C2(n5843), .A(n5619), .B(n5618), .ZN(U2964)
         );
  AOI21_X1 U6750 ( .B1(n5621), .B2(n5620), .A(n3005), .ZN(n5761) );
  NAND2_X1 U6751 ( .A1(n6338), .A2(REIP_REG_21__SCAN_IN), .ZN(n5755) );
  OAI21_X1 U6752 ( .B1(n5646), .B2(n5622), .A(n5755), .ZN(n5624) );
  NOR2_X1 U6753 ( .A1(n5903), .A2(n6271), .ZN(n5623) );
  AOI211_X1 U6754 ( .C1(n5649), .C2(n5625), .A(n5624), .B(n5623), .ZN(n5626)
         );
  OAI21_X1 U6755 ( .B1(n5761), .B2(n6273), .A(n5626), .ZN(U2965) );
  XNOR2_X1 U6756 ( .A(n5917), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5627)
         );
  XNOR2_X1 U6757 ( .A(n5628), .B(n5627), .ZN(n5766) );
  NAND2_X1 U6758 ( .A1(n5766), .A2(n6257), .ZN(n5632) );
  AND2_X1 U6759 ( .A1(n6338), .A2(REIP_REG_20__SCAN_IN), .ZN(n5769) );
  NOR2_X1 U6760 ( .A1(n6264), .A2(n5629), .ZN(n5630) );
  AOI211_X1 U6761 ( .C1(n6276), .C2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5769), 
        .B(n5630), .ZN(n5631) );
  OAI211_X1 U6762 ( .C1(n6271), .C2(n5633), .A(n5632), .B(n5631), .ZN(U2966)
         );
  NOR3_X1 U6763 ( .A1(n5634), .A2(n5917), .A3(n5939), .ZN(n5922) );
  NAND2_X1 U6764 ( .A1(n5917), .A2(n5948), .ZN(n5919) );
  NOR3_X1 U6765 ( .A1(n5635), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5919), 
        .ZN(n5920) );
  NOR2_X1 U6766 ( .A1(n5922), .A2(n5920), .ZN(n5636) );
  XNOR2_X1 U6767 ( .A(n5636), .B(n5764), .ZN(n5784) );
  INV_X1 U6768 ( .A(n5637), .ZN(n5639) );
  NAND2_X1 U6769 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5638)
         );
  NAND2_X1 U6770 ( .A1(n6338), .A2(REIP_REG_18__SCAN_IN), .ZN(n5778) );
  OAI211_X1 U6771 ( .C1(n6264), .C2(n5639), .A(n5638), .B(n5778), .ZN(n5640)
         );
  AOI21_X1 U6772 ( .B1(n6119), .B2(n6258), .A(n5640), .ZN(n5641) );
  OAI21_X1 U6773 ( .B1(n5784), .B2(n6273), .A(n5641), .ZN(U2968) );
  OAI21_X1 U6774 ( .B1(n5917), .B2(n5948), .A(n5919), .ZN(n5642) );
  XNOR2_X1 U6775 ( .A(n5643), .B(n5642), .ZN(n5945) );
  NAND2_X1 U6776 ( .A1(n5945), .A2(n6257), .ZN(n5651) );
  INV_X1 U6777 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5644) );
  OAI22_X1 U6778 ( .A1(n5646), .A2(n5645), .B1(n5966), .B2(n5644), .ZN(n5647)
         );
  AOI21_X1 U6779 ( .B1(n5649), .B2(n5648), .A(n5647), .ZN(n5650) );
  OAI211_X1 U6780 ( .C1(n6271), .C2(n5652), .A(n5651), .B(n5650), .ZN(U2970)
         );
  XNOR2_X1 U6781 ( .A(n3493), .B(n5942), .ZN(n5654) );
  XNOR2_X1 U6782 ( .A(n5653), .B(n5654), .ZN(n5793) );
  AOI22_X1 U6783 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6338), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5655) );
  OAI21_X1 U6784 ( .B1(n6264), .B2(n5656), .A(n5655), .ZN(n5657) );
  AOI21_X1 U6785 ( .B1(n6105), .B2(n6258), .A(n5657), .ZN(n5658) );
  OAI21_X1 U6786 ( .B1(n5793), .B2(n6273), .A(n5658), .ZN(U2971) );
  XNOR2_X1 U6787 ( .A(n3493), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5660)
         );
  XNOR2_X1 U6788 ( .A(n5659), .B(n5660), .ZN(n5962) );
  INV_X1 U6789 ( .A(n5962), .ZN(n5667) );
  INV_X1 U6790 ( .A(n5661), .ZN(n5665) );
  AOI22_X1 U6791 ( .A1(n6276), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6338), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5662) );
  OAI21_X1 U6792 ( .B1(n5663), .B2(n6264), .A(n5662), .ZN(n5664) );
  AOI21_X1 U6793 ( .B1(n5665), .B2(n6258), .A(n5664), .ZN(n5666) );
  OAI21_X1 U6794 ( .B1(n5667), .B2(n6273), .A(n5666), .ZN(U2972) );
  NAND3_X1 U6795 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5668), .ZN(n5669) );
  OAI211_X1 U6796 ( .C1(n5671), .C2(n6358), .A(n5670), .B(n5669), .ZN(n5672)
         );
  AOI21_X1 U6797 ( .B1(n5673), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5672), 
        .ZN(n5674) );
  OAI21_X1 U6798 ( .B1(n5675), .B2(n6313), .A(n5674), .ZN(U2988) );
  INV_X1 U6799 ( .A(n5676), .ZN(n5678) );
  OAI21_X1 U6800 ( .B1(n5678), .B2(n6358), .A(n5677), .ZN(n5681) );
  NOR2_X1 U6801 ( .A1(n5679), .A2(n5682), .ZN(n5680) );
  AOI211_X1 U6802 ( .C1(n5683), .C2(n5682), .A(n5681), .B(n5680), .ZN(n5684)
         );
  OAI21_X1 U6803 ( .B1(n5685), .B2(n6313), .A(n5684), .ZN(U2989) );
  INV_X1 U6804 ( .A(n5705), .ZN(n5688) );
  INV_X1 U6805 ( .A(n5686), .ZN(n5690) );
  INV_X1 U6806 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U6807 ( .A1(n5690), .A2(n5687), .ZN(n5703) );
  AOI21_X1 U6808 ( .B1(n5688), .B2(n5703), .A(n5689), .ZN(n5695) );
  NAND3_X1 U6809 ( .A1(n5690), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5689), .ZN(n5692) );
  OAI211_X1 U6810 ( .C1(n6358), .C2(n5693), .A(n5692), .B(n5691), .ZN(n5694)
         );
  NOR2_X1 U6811 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  OAI21_X1 U6812 ( .B1(n5697), .B2(n6313), .A(n5696), .ZN(U2990) );
  AND2_X1 U6813 ( .A1(n3002), .A2(n5698), .ZN(n5699) );
  NOR2_X1 U6814 ( .A1(n5700), .A2(n5699), .ZN(n5876) );
  NAND2_X1 U6815 ( .A1(n5876), .A2(n6340), .ZN(n5701) );
  NAND3_X1 U6816 ( .A1(n5703), .A2(n5702), .A3(n5701), .ZN(n5704) );
  AOI21_X1 U6817 ( .B1(n5705), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5704), 
        .ZN(n5706) );
  OAI21_X1 U6818 ( .B1(n5707), .B2(n6313), .A(n5706), .ZN(U2991) );
  INV_X1 U6819 ( .A(n5726), .ZN(n5722) );
  XNOR2_X1 U6820 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6821 ( .A1(n5708), .A2(n6340), .ZN(n5709) );
  OAI211_X1 U6822 ( .C1(n5715), .C2(n5711), .A(n5710), .B(n5709), .ZN(n5712)
         );
  AOI21_X1 U6823 ( .B1(n5722), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5712), 
        .ZN(n5713) );
  OAI21_X1 U6824 ( .B1(n5714), .B2(n6313), .A(n5713), .ZN(U2992) );
  NOR2_X1 U6825 ( .A1(n5715), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5721)
         );
  OR2_X1 U6826 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  NAND2_X1 U6827 ( .A1(n3004), .A2(n5718), .ZN(n5879) );
  OAI21_X1 U6828 ( .B1(n5879), .B2(n6358), .A(n5719), .ZN(n5720) );
  AOI211_X1 U6829 ( .C1(n5722), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5721), .B(n5720), .ZN(n5723) );
  OAI21_X1 U6830 ( .B1(n5724), .B2(n6313), .A(n5723), .ZN(U2993) );
  INV_X1 U6831 ( .A(n5738), .ZN(n5725) );
  NAND3_X1 U6832 ( .A1(n5926), .A2(n5725), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5727) );
  AOI21_X1 U6833 ( .B1(n5728), .B2(n5727), .A(n5726), .ZN(n5729) );
  AOI211_X1 U6834 ( .C1(n6340), .C2(n5731), .A(n5730), .B(n5729), .ZN(n5732)
         );
  OAI21_X1 U6835 ( .B1(n5733), .B2(n6313), .A(n5732), .ZN(U2994) );
  NAND2_X1 U6836 ( .A1(n5734), .A2(n6354), .ZN(n5743) );
  AOI21_X1 U6837 ( .B1(n5737), .B2(n5736), .A(n5735), .ZN(n5883) );
  INV_X1 U6838 ( .A(n5926), .ZN(n5739) );
  NOR3_X1 U6839 ( .A1(n5739), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5738), 
        .ZN(n5740) );
  AOI211_X1 U6840 ( .C1(n6340), .C2(n5883), .A(n5741), .B(n5740), .ZN(n5742)
         );
  OAI211_X1 U6841 ( .C1(n5745), .C2(n5744), .A(n5743), .B(n5742), .ZN(U2995)
         );
  AND2_X1 U6842 ( .A1(n5767), .A2(n5746), .ZN(n5747) );
  NAND2_X1 U6843 ( .A1(n5926), .A2(n5747), .ZN(n5756) );
  AOI21_X1 U6844 ( .B1(n5754), .B2(n5756), .A(n6692), .ZN(n5751) );
  NAND4_X1 U6845 ( .A1(n5926), .A2(n5767), .A3(INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n6692), .ZN(n5749) );
  OAI211_X1 U6846 ( .C1(n6358), .C2(n5842), .A(n5749), .B(n5748), .ZN(n5750)
         );
  AOI211_X1 U6847 ( .C1(n5752), .C2(n6354), .A(n5751), .B(n5750), .ZN(n5753)
         );
  INV_X1 U6848 ( .A(n5753), .ZN(U2996) );
  INV_X1 U6849 ( .A(n5754), .ZN(n5759) );
  OAI211_X1 U6850 ( .C1(n6358), .C2(n5757), .A(n5756), .B(n5755), .ZN(n5758)
         );
  AOI21_X1 U6851 ( .B1(n5759), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5758), 
        .ZN(n5760) );
  OAI21_X1 U6852 ( .B1(n5761), .B2(n6313), .A(n5760), .ZN(U2997) );
  AND2_X1 U6853 ( .A1(n5762), .A2(n5939), .ZN(n5763) );
  NOR2_X1 U6854 ( .A1(n5934), .A2(n5763), .ZN(n5776) );
  NAND2_X1 U6855 ( .A1(n5789), .A2(n5764), .ZN(n5765) );
  AND2_X1 U6856 ( .A1(n5776), .A2(n5765), .ZN(n5933) );
  NAND2_X1 U6857 ( .A1(n5766), .A2(n6354), .ZN(n5775) );
  NOR2_X1 U6858 ( .A1(n5768), .A2(n5767), .ZN(n5773) );
  INV_X1 U6859 ( .A(n5769), .ZN(n5770) );
  OAI21_X1 U6860 ( .B1(n5771), .B2(n6358), .A(n5770), .ZN(n5772) );
  AOI21_X1 U6861 ( .B1(n5926), .B2(n5773), .A(n5772), .ZN(n5774) );
  OAI211_X1 U6862 ( .C1(n5933), .C2(n6659), .A(n5775), .B(n5774), .ZN(U2998)
         );
  INV_X1 U6863 ( .A(n5776), .ZN(n5782) );
  NOR2_X1 U6864 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5939), .ZN(n5777)
         );
  NAND2_X1 U6865 ( .A1(n5935), .A2(n5777), .ZN(n5779) );
  OAI211_X1 U6866 ( .C1(n6358), .C2(n5780), .A(n5779), .B(n5778), .ZN(n5781)
         );
  AOI21_X1 U6867 ( .B1(n5782), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5781), 
        .ZN(n5783) );
  OAI21_X1 U6868 ( .B1(n5784), .B2(n6313), .A(n5783), .ZN(U3000) );
  XNOR2_X1 U6869 ( .A(n5786), .B(n5785), .ZN(n6104) );
  NAND2_X1 U6870 ( .A1(n5787), .A2(n5958), .ZN(n5941) );
  AOI21_X1 U6871 ( .B1(n5789), .B2(n5788), .A(n5954), .ZN(n5949) );
  NAND2_X1 U6872 ( .A1(n6338), .A2(REIP_REG_15__SCAN_IN), .ZN(n5790) );
  OAI221_X1 U6873 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5941), .C1(
        n5942), .C2(n5949), .A(n5790), .ZN(n5791) );
  AOI21_X1 U6874 ( .B1(n6340), .B2(n6104), .A(n5791), .ZN(n5792) );
  OAI21_X1 U6875 ( .B1(n5793), .B2(n6313), .A(n5792), .ZN(U3003) );
  OAI211_X1 U6876 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4259), .A(n5797), .B(
        n6612), .ZN(n5794) );
  OAI21_X1 U6877 ( .B1(n5798), .B2(n5795), .A(n5794), .ZN(n5796) );
  MUX2_X1 U6878 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5796), .S(n6364), 
        .Z(U3464) );
  XNOR2_X1 U6879 ( .A(n3079), .B(n5797), .ZN(n5800) );
  OAI22_X1 U6880 ( .A1(n5800), .A2(n5799), .B1(n4261), .B2(n5798), .ZN(n5801)
         );
  MUX2_X1 U6881 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5801), .S(n6364), 
        .Z(U3463) );
  AND2_X1 U6882 ( .A1(n5802), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6883 ( .B1(n5804), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n5803), .ZN(
        n5805) );
  INV_X1 U6884 ( .A(n5805), .ZN(U2788) );
  INV_X1 U6885 ( .A(n5806), .ZN(n5810) );
  INV_X1 U6886 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5878) );
  OAI22_X1 U6887 ( .A1(n5878), .A2(n6080), .B1(n5807), .B2(n6093), .ZN(n5808)
         );
  AOI221_X1 U6888 ( .B1(n5819), .B2(REIP_REG_27__SCAN_IN), .C1(n5810), .C2(
        n5809), .A(n5808), .ZN(n5812) );
  AOI22_X1 U6889 ( .A1(n5891), .A2(n6064), .B1(n5876), .B2(n6090), .ZN(n5811)
         );
  OAI211_X1 U6890 ( .C1(n5813), .C2(n6103), .A(n5812), .B(n5811), .ZN(U2800)
         );
  AOI22_X1 U6891 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6053), .B1(n5814), 
        .B2(n6072), .ZN(n5821) );
  NAND2_X1 U6892 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5823), .ZN(n5828) );
  OAI21_X1 U6893 ( .B1(n5825), .B2(n5828), .A(n6569), .ZN(n5818) );
  OAI22_X1 U6894 ( .A1(n5816), .A2(n5872), .B1(n5815), .B2(n6079), .ZN(n5817)
         );
  AOI21_X1 U6895 ( .B1(n5819), .B2(n5818), .A(n5817), .ZN(n5820) );
  OAI211_X1 U6896 ( .C1(n5822), .C2(n6080), .A(n5821), .B(n5820), .ZN(U2801)
         );
  AOI21_X1 U6897 ( .B1(n5823), .B2(n6565), .A(n5837), .ZN(n5826) );
  OAI22_X1 U6898 ( .A1(n5826), .A2(n5825), .B1(n5824), .B2(n6103), .ZN(n5830)
         );
  OAI22_X1 U6899 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5828), .B1(n5827), .B2(
        n6093), .ZN(n5829) );
  AOI211_X1 U6900 ( .C1(EBX_REG_25__SCAN_IN), .C2(n6091), .A(n5830), .B(n5829), 
        .ZN(n5833) );
  NOR2_X1 U6901 ( .A1(n5879), .A2(n6079), .ZN(n5831) );
  AOI21_X1 U6902 ( .B1(n5894), .B2(n6064), .A(n5831), .ZN(n5832) );
  NAND2_X1 U6903 ( .A1(n5833), .A2(n5832), .ZN(U2802) );
  NAND2_X1 U6904 ( .A1(n5834), .A2(n6563), .ZN(n5836) );
  INV_X1 U6905 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6757) );
  OAI22_X1 U6906 ( .A1(n6757), .A2(n6080), .B1(n3908), .B2(n6093), .ZN(n5835)
         );
  AOI21_X1 U6907 ( .B1(n5837), .B2(n5836), .A(n5835), .ZN(n5840) );
  INV_X1 U6908 ( .A(n5838), .ZN(n5900) );
  AOI22_X1 U6909 ( .A1(n5900), .A2(n6064), .B1(n5883), .B2(n6090), .ZN(n5839)
         );
  OAI211_X1 U6910 ( .C1(n5841), .C2(n6103), .A(n5840), .B(n5839), .ZN(U2804)
         );
  AOI22_X1 U6911 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6091), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6053), .ZN(n5853) );
  OAI22_X1 U6912 ( .A1(n5843), .A2(n5872), .B1(n5842), .B2(n6079), .ZN(n5844)
         );
  AOI21_X1 U6913 ( .B1(n5845), .B2(n6072), .A(n5844), .ZN(n5852) );
  NAND3_X1 U6914 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5847), .A3(n5846), .ZN(
        n5851) );
  OAI211_X1 U6915 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5849), .B(n5848), .ZN(n5850) );
  NAND4_X1 U6916 ( .A1(n5853), .A2(n5852), .A3(n5851), .A4(n5850), .ZN(U2805)
         );
  INV_X1 U6917 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5859) );
  INV_X1 U6918 ( .A(n5854), .ZN(n5857) );
  NOR2_X1 U6919 ( .A1(n6007), .A2(n5855), .ZN(n5856) );
  MUX2_X1 U6920 ( .A(n5857), .B(n5856), .S(REIP_REG_19__SCAN_IN), .Z(n5858) );
  OAI211_X1 U6921 ( .C1(n6093), .C2(n5859), .A(n5858), .B(n6055), .ZN(n5860)
         );
  AOI21_X1 U6922 ( .B1(EBX_REG_19__SCAN_IN), .B2(n6091), .A(n5860), .ZN(n5875)
         );
  NAND2_X1 U6923 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  NAND2_X1 U6924 ( .A1(n5864), .A2(n5863), .ZN(n5912) );
  NAND2_X1 U6925 ( .A1(n5865), .A2(n5867), .ZN(n5871) );
  INV_X1 U6926 ( .A(n5866), .ZN(n5868) );
  NOR2_X1 U6927 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  AOI21_X1 U6928 ( .B1(n5871), .B2(n5870), .A(n5869), .ZN(n5927) );
  OAI22_X1 U6929 ( .A1(n5912), .A2(n5872), .B1(n5927), .B2(n6079), .ZN(n5873)
         );
  INV_X1 U6930 ( .A(n5873), .ZN(n5874) );
  OAI211_X1 U6931 ( .C1(n5916), .C2(n6103), .A(n5875), .B(n5874), .ZN(U2808)
         );
  AOI22_X1 U6932 ( .A1(n5891), .A2(n6116), .B1(n5876), .B2(n6115), .ZN(n5877)
         );
  OAI21_X1 U6933 ( .B1(n6118), .B2(n5878), .A(n5877), .ZN(U2832) );
  NOR2_X1 U6934 ( .A1(n5879), .A2(n5885), .ZN(n5880) );
  AOI21_X1 U6935 ( .B1(n5894), .B2(n6116), .A(n5880), .ZN(n5881) );
  OAI21_X1 U6936 ( .B1(n6118), .B2(n5882), .A(n5881), .ZN(U2834) );
  AOI22_X1 U6937 ( .A1(n5900), .A2(n6116), .B1(n5883), .B2(n6115), .ZN(n5884)
         );
  OAI21_X1 U6938 ( .B1(n6118), .B2(n6757), .A(n5884), .ZN(U2836) );
  OAI22_X1 U6939 ( .A1(n5912), .A2(n5886), .B1(n5927), .B2(n5885), .ZN(n5887)
         );
  INV_X1 U6940 ( .A(n5887), .ZN(n5888) );
  OAI21_X1 U6941 ( .B1(n6118), .B2(n5889), .A(n5888), .ZN(U2840) );
  AOI22_X1 U6942 ( .A1(n5891), .A2(n6123), .B1(n6122), .B2(DATAI_27_), .ZN(
        n5893) );
  AOI22_X1 U6943 ( .A1(n6126), .A2(DATAI_11_), .B1(n6125), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U6944 ( .A1(n5893), .A2(n5892), .ZN(U2864) );
  AOI22_X1 U6945 ( .A1(n5894), .A2(n6123), .B1(n6122), .B2(DATAI_25_), .ZN(
        n5896) );
  AOI22_X1 U6946 ( .A1(n6126), .A2(DATAI_9_), .B1(n6125), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U6947 ( .A1(n5896), .A2(n5895), .ZN(U2866) );
  AOI22_X1 U6948 ( .A1(n5897), .A2(n6123), .B1(n6122), .B2(DATAI_24_), .ZN(
        n5899) );
  AOI22_X1 U6949 ( .A1(n6126), .A2(DATAI_8_), .B1(n6125), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U6950 ( .A1(n5899), .A2(n5898), .ZN(U2867) );
  AOI22_X1 U6951 ( .A1(n5900), .A2(n6123), .B1(n6122), .B2(DATAI_23_), .ZN(
        n5902) );
  AOI22_X1 U6952 ( .A1(n6126), .A2(DATAI_7_), .B1(n6125), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U6953 ( .A1(n5902), .A2(n5901), .ZN(U2868) );
  INV_X1 U6954 ( .A(n5903), .ZN(n5904) );
  AOI22_X1 U6955 ( .A1(n5904), .A2(n6123), .B1(n6122), .B2(DATAI_21_), .ZN(
        n5906) );
  AOI22_X1 U6956 ( .A1(n6126), .A2(DATAI_5_), .B1(n6125), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U6957 ( .A1(n5906), .A2(n5905), .ZN(U2870) );
  INV_X1 U6958 ( .A(n5912), .ZN(n5907) );
  AOI22_X1 U6959 ( .A1(n5907), .A2(n6123), .B1(n6122), .B2(DATAI_19_), .ZN(
        n5909) );
  AOI22_X1 U6960 ( .A1(n6126), .A2(DATAI_3_), .B1(n6125), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U6961 ( .A1(n5909), .A2(n5908), .ZN(U2872) );
  AOI22_X1 U6962 ( .A1(n6338), .A2(REIP_REG_19__SCAN_IN), .B1(n6276), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5915) );
  OAI21_X1 U6963 ( .B1(n5592), .B2(n5911), .A(n5910), .ZN(n5928) );
  OAI22_X1 U6964 ( .A1(n5928), .A2(n6273), .B1(n6271), .B2(n5912), .ZN(n5913)
         );
  INV_X1 U6965 ( .A(n5913), .ZN(n5914) );
  OAI211_X1 U6966 ( .C1(n6264), .C2(n5916), .A(n5915), .B(n5914), .ZN(U2967)
         );
  AOI22_X1 U6967 ( .A1(n6338), .A2(REIP_REG_17__SCAN_IN), .B1(n6276), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5925) );
  AOI21_X1 U6968 ( .B1(n5917), .B2(n5939), .A(n5634), .ZN(n5918) );
  AOI21_X1 U6969 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5919), .A(n5918), 
        .ZN(n5923) );
  INV_X1 U6970 ( .A(n5920), .ZN(n5921) );
  OAI21_X1 U6971 ( .B1(n5923), .B2(n5922), .A(n5921), .ZN(n5936) );
  AOI22_X1 U6972 ( .A1(n5936), .A2(n6257), .B1(n6258), .B2(n6124), .ZN(n5924)
         );
  OAI211_X1 U6973 ( .C1(n6264), .C2(n6014), .A(n5925), .B(n5924), .ZN(U2969)
         );
  AOI22_X1 U6974 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6338), .B1(n5926), .B2(
        n5932), .ZN(n5931) );
  OAI22_X1 U6975 ( .A1(n5928), .A2(n6313), .B1(n5927), .B2(n6358), .ZN(n5929)
         );
  INV_X1 U6976 ( .A(n5929), .ZN(n5930) );
  OAI211_X1 U6977 ( .C1(n5933), .C2(n5932), .A(n5931), .B(n5930), .ZN(U2999)
         );
  INV_X1 U6978 ( .A(n5934), .ZN(n5940) );
  AOI22_X1 U6979 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6338), .B1(n5935), .B2(
        n5939), .ZN(n5938) );
  AOI22_X1 U6980 ( .A1(n5936), .A2(n6354), .B1(n6340), .B2(n6011), .ZN(n5937)
         );
  OAI211_X1 U6981 ( .C1(n5940), .C2(n5939), .A(n5938), .B(n5937), .ZN(U3001)
         );
  AOI221_X1 U6982 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n5942), .C2(n5948), .A(n5941), 
        .ZN(n5943) );
  AOI21_X1 U6983 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6338), .A(n5943), .ZN(n5947) );
  AOI22_X1 U6984 ( .A1(n5945), .A2(n6354), .B1(n6340), .B2(n5944), .ZN(n5946)
         );
  OAI211_X1 U6985 ( .C1(n5949), .C2(n5948), .A(n5947), .B(n5946), .ZN(U3002)
         );
  NAND2_X1 U6986 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5955) );
  NOR3_X1 U6987 ( .A1(n5950), .A2(n5965), .A3(n6363), .ZN(n5951) );
  NOR2_X1 U6988 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5955), .ZN(n5971)
         );
  OAI21_X1 U6989 ( .B1(n5952), .B2(n5951), .A(n5971), .ZN(n5973) );
  OAI21_X1 U6990 ( .B1(n5957), .B2(n6362), .A(n5973), .ZN(n5953) );
  AOI211_X1 U6991 ( .C1(n5956), .C2(n5955), .A(n5954), .B(n5953), .ZN(n5975)
         );
  AND3_X1 U6992 ( .A1(n6653), .A2(n5958), .A3(n5957), .ZN(n5959) );
  AOI21_X1 U6993 ( .B1(REIP_REG_14__SCAN_IN), .B2(n6338), .A(n5959), .ZN(n5964) );
  INV_X1 U6994 ( .A(n5960), .ZN(n5961) );
  AOI22_X1 U6995 ( .A1(n5962), .A2(n6354), .B1(n6340), .B2(n5961), .ZN(n5963)
         );
  OAI211_X1 U6996 ( .C1(n5975), .C2(n6653), .A(n5964), .B(n5963), .ZN(U3004)
         );
  NOR2_X1 U6997 ( .A1(n6362), .A2(n5965), .ZN(n5970) );
  INV_X1 U6998 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6548) );
  NOR2_X1 U6999 ( .A1(n5966), .A2(n6548), .ZN(n5969) );
  OAI22_X1 U7000 ( .A1(n5967), .A2(n6313), .B1(n6358), .B2(n6023), .ZN(n5968)
         );
  AOI211_X1 U7001 ( .C1(n5971), .C2(n5970), .A(n5969), .B(n5968), .ZN(n5972)
         );
  OAI211_X1 U7002 ( .C1(n5975), .C2(n5974), .A(n5973), .B(n5972), .ZN(U3005)
         );
  OR4_X1 U7003 ( .A1(n5978), .A2(n5977), .A3(n6597), .A4(n5976), .ZN(n5979) );
  OAI21_X1 U7004 ( .B1(n6593), .B2(n5980), .A(n5979), .ZN(U3455) );
  INV_X1 U7005 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6528) );
  AOI21_X1 U7006 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6528), .A(n6519), .ZN(n5985) );
  INV_X1 U7007 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5981) );
  INV_X1 U7008 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6518) );
  NOR2_X2 U7009 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6518), .ZN(n6622) );
  AOI21_X1 U7010 ( .B1(n5985), .B2(n5981), .A(n6622), .ZN(U2789) );
  OAI21_X1 U7011 ( .B1(n5982), .B2(n6502), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5983) );
  OAI21_X1 U7012 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6503), .A(n5983), .ZN(
        U2790) );
  NOR2_X1 U7013 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5986) );
  OAI21_X1 U7014 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5986), .A(n6608), .ZN(n5984)
         );
  OAI21_X1 U7015 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6608), .A(n5984), .ZN(
        U2791) );
  NOR2_X1 U7016 ( .A1(n6622), .A2(n5985), .ZN(n6585) );
  OAI21_X1 U7017 ( .B1(BS16_N), .B2(n5986), .A(n6585), .ZN(n6583) );
  OAI21_X1 U7018 ( .B1(n6585), .B2(n5987), .A(n6583), .ZN(U2792) );
  AOI21_X1 U7019 ( .B1(n5988), .B2(FLUSH_REG_SCAN_IN), .A(n6257), .ZN(n5989)
         );
  INV_X1 U7020 ( .A(n5989), .ZN(U2793) );
  NOR4_X1 U7021 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n5993) );
  NOR4_X1 U7022 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5992) );
  NOR4_X1 U7023 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5991) );
  NOR4_X1 U7024 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n5990) );
  NAND4_X1 U7025 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n5999)
         );
  NOR4_X1 U7026 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n5997) );
  AOI211_X1 U7027 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_21__SCAN_IN), .B(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n5996) );
  NOR4_X1 U7028 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5995) );
  NOR4_X1 U7029 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5994) );
  NAND4_X1 U7030 ( .A1(n5997), .A2(n5996), .A3(n5995), .A4(n5994), .ZN(n5998)
         );
  NOR2_X1 U7031 ( .A1(n5999), .A2(n5998), .ZN(n6606) );
  INV_X1 U7032 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6001) );
  NOR3_X1 U7033 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6002) );
  OAI21_X1 U7034 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6002), .A(n6606), .ZN(n6000)
         );
  OAI21_X1 U7035 ( .B1(n6606), .B2(n6001), .A(n6000), .ZN(U2794) );
  INV_X1 U7036 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6584) );
  AOI21_X1 U7037 ( .B1(n6599), .B2(n6584), .A(n6002), .ZN(n6004) );
  INV_X1 U7038 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6003) );
  INV_X1 U7039 ( .A(n6606), .ZN(n6601) );
  AOI22_X1 U7040 ( .A1(n6606), .A2(n6004), .B1(n6003), .B2(n6601), .ZN(U2795)
         );
  AOI21_X1 U7041 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6005), .A(
        REIP_REG_17__SCAN_IN), .ZN(n6006) );
  INV_X1 U7042 ( .A(n6006), .ZN(n6008) );
  AOI22_X1 U7043 ( .A1(n6008), .A2(n6007), .B1(PHYADDRPOINTER_REG_17__SCAN_IN), 
        .B2(n6053), .ZN(n6009) );
  OAI211_X1 U7044 ( .C1(n6080), .C2(n5515), .A(n6055), .B(n6009), .ZN(n6010)
         );
  INV_X1 U7045 ( .A(n6010), .ZN(n6013) );
  AOI22_X1 U7046 ( .A1(n6124), .A2(n6064), .B1(n6090), .B2(n6011), .ZN(n6012)
         );
  OAI211_X1 U7047 ( .C1(n6014), .C2(n6103), .A(n6013), .B(n6012), .ZN(U2810)
         );
  AOI22_X1 U7048 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6091), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6015), .ZN(n6018) );
  AOI211_X1 U7049 ( .C1(n6053), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6070), 
        .B(n6016), .ZN(n6017) );
  NAND2_X1 U7050 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  AOI21_X1 U7051 ( .B1(n6105), .B2(n6064), .A(n6019), .ZN(n6022) );
  AOI22_X1 U7052 ( .A1(n6072), .A2(n6020), .B1(n6090), .B2(n6104), .ZN(n6021)
         );
  NAND2_X1 U7053 ( .A1(n6022), .A2(n6021), .ZN(U2812) );
  OAI22_X1 U7054 ( .A1(n6103), .A2(n6024), .B1(n6079), .B2(n6023), .ZN(n6025)
         );
  AOI211_X1 U7055 ( .C1(n6053), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6070), 
        .B(n6025), .ZN(n6032) );
  NAND2_X1 U7056 ( .A1(n6027), .A2(n6026), .ZN(n6041) );
  XNOR2_X1 U7057 ( .A(n6548), .B(n5244), .ZN(n6028) );
  OAI22_X1 U7058 ( .A1(n6041), .A2(n6028), .B1(n6548), .B2(n6035), .ZN(n6029)
         );
  AOI21_X1 U7059 ( .B1(n6030), .B2(n6064), .A(n6029), .ZN(n6031) );
  OAI211_X1 U7060 ( .C1(n6752), .C2(n6080), .A(n6032), .B(n6031), .ZN(U2814)
         );
  INV_X1 U7061 ( .A(n6033), .ZN(n6108) );
  AOI22_X1 U7062 ( .A1(n6091), .A2(EBX_REG_12__SCAN_IN), .B1(n6090), .B2(n6108), .ZN(n6034) );
  OAI21_X1 U7063 ( .B1(n5244), .B2(n6035), .A(n6034), .ZN(n6036) );
  AOI211_X1 U7064 ( .C1(n6053), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6070), 
        .B(n6036), .ZN(n6040) );
  INV_X1 U7065 ( .A(n6037), .ZN(n6109) );
  AOI22_X1 U7066 ( .A1(n6109), .A2(n6064), .B1(n6038), .B2(n6072), .ZN(n6039)
         );
  OAI211_X1 U7067 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6041), .A(n6040), .B(n6039), .ZN(U2815) );
  AOI22_X1 U7068 ( .A1(n6091), .A2(EBX_REG_10__SCAN_IN), .B1(n6090), .B2(n3015), .ZN(n6050) );
  INV_X1 U7069 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6543) );
  NOR3_X1 U7070 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6543), .A3(n6042), .ZN(n6043) );
  AOI211_X1 U7071 ( .C1(n6053), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6070), 
        .B(n6043), .ZN(n6049) );
  AOI22_X1 U7072 ( .A1(n6112), .A2(n6064), .B1(n6072), .B2(n6044), .ZN(n6048)
         );
  OAI21_X1 U7073 ( .B1(n6046), .B2(n6045), .A(REIP_REG_10__SCAN_IN), .ZN(n6047) );
  NAND4_X1 U7074 ( .A1(n6050), .A2(n6049), .A3(n6048), .A4(n6047), .ZN(U2817)
         );
  INV_X1 U7075 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6538) );
  XNOR2_X1 U7076 ( .A(n6052), .B(n6051), .ZN(n6300) );
  NAND2_X1 U7077 ( .A1(n6090), .A2(n6300), .ZN(n6056) );
  NAND2_X1 U7078 ( .A1(n6053), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6054)
         );
  NAND3_X1 U7079 ( .A1(n6056), .A2(n6055), .A3(n6054), .ZN(n6061) );
  OAI21_X1 U7080 ( .B1(REIP_REG_7__SCAN_IN), .B2(REIP_REG_6__SCAN_IN), .A(
        n6057), .ZN(n6058) );
  NOR2_X1 U7081 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  AOI211_X1 U7082 ( .C1(n6091), .C2(EBX_REG_7__SCAN_IN), .A(n6061), .B(n6060), 
        .ZN(n6062) );
  OAI21_X1 U7083 ( .B1(n6538), .B2(n6075), .A(n6062), .ZN(n6063) );
  AOI21_X1 U7084 ( .B1(n6064), .B2(n6237), .A(n6063), .ZN(n6065) );
  OAI21_X1 U7085 ( .B1(n6240), .B2(n6103), .A(n6065), .ZN(U2820) );
  NOR2_X1 U7086 ( .A1(n6066), .A2(REIP_REG_5__SCAN_IN), .ZN(n6076) );
  INV_X1 U7087 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6067) );
  OAI22_X1 U7088 ( .A1(n6079), .A2(n6068), .B1(n6067), .B2(n6093), .ZN(n6069)
         );
  AOI211_X1 U7089 ( .C1(n6091), .C2(EBX_REG_5__SCAN_IN), .A(n6070), .B(n6069), 
        .ZN(n6074) );
  INV_X1 U7090 ( .A(n6245), .ZN(n6071) );
  AOI22_X1 U7091 ( .A1(n6100), .A2(n6241), .B1(n6072), .B2(n6071), .ZN(n6073)
         );
  OAI211_X1 U7092 ( .C1(n6076), .C2(n6075), .A(n6074), .B(n6073), .ZN(U2822)
         );
  INV_X1 U7093 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6078) );
  OAI22_X1 U7094 ( .A1(n6078), .A2(n6093), .B1(n6092), .B2(n6077), .ZN(n6082)
         );
  OAI22_X1 U7095 ( .A1(n6753), .A2(n6080), .B1(n6079), .B2(n6329), .ZN(n6081)
         );
  AOI211_X1 U7096 ( .C1(n6100), .C2(n6250), .A(n6082), .B(n6081), .ZN(n6088)
         );
  AOI21_X1 U7097 ( .B1(n6084), .B2(REIP_REG_1__SCAN_IN), .A(n6083), .ZN(n6085)
         );
  INV_X1 U7098 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6531) );
  NOR2_X1 U7099 ( .A1(n6085), .A2(n6531), .ZN(n6096) );
  OAI21_X1 U7100 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6096), .A(n6086), .ZN(n6087)
         );
  OAI211_X1 U7101 ( .C1(n6103), .C2(n6253), .A(n6088), .B(n6087), .ZN(U2824)
         );
  INV_X1 U7102 ( .A(n6089), .ZN(n6339) );
  AOI22_X1 U7103 ( .A1(n6091), .A2(EBX_REG_2__SCAN_IN), .B1(n6090), .B2(n6339), 
        .ZN(n6102) );
  INV_X1 U7104 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6094) );
  OAI22_X1 U7105 ( .A1(n6094), .A2(n6093), .B1(n6092), .B2(n4261), .ZN(n6099)
         );
  NAND2_X1 U7106 ( .A1(n6095), .A2(REIP_REG_1__SCAN_IN), .ZN(n6097) );
  AOI21_X1 U7107 ( .B1(n6531), .B2(n6097), .A(n6096), .ZN(n6098) );
  AOI211_X1 U7108 ( .C1(n6259), .C2(n6100), .A(n6099), .B(n6098), .ZN(n6101)
         );
  OAI211_X1 U7109 ( .C1(n6262), .C2(n6103), .A(n6102), .B(n6101), .ZN(U2825)
         );
  AOI22_X1 U7110 ( .A1(n6105), .A2(n6116), .B1(n6115), .B2(n6104), .ZN(n6106)
         );
  OAI21_X1 U7111 ( .B1(n6118), .B2(n6107), .A(n6106), .ZN(U2844) );
  INV_X1 U7112 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6111) );
  AOI22_X1 U7113 ( .A1(n6109), .A2(n6116), .B1(n6115), .B2(n6108), .ZN(n6110)
         );
  OAI21_X1 U7114 ( .B1(n6118), .B2(n6111), .A(n6110), .ZN(U2847) );
  INV_X1 U7115 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6114) );
  AOI22_X1 U7116 ( .A1(n6112), .A2(n6116), .B1(n6115), .B2(n3015), .ZN(n6113)
         );
  OAI21_X1 U7117 ( .B1(n6118), .B2(n6114), .A(n6113), .ZN(U2849) );
  AOI22_X1 U7118 ( .A1(n6237), .A2(n6116), .B1(n6115), .B2(n6300), .ZN(n6117)
         );
  OAI21_X1 U7119 ( .B1(n6118), .B2(n6735), .A(n6117), .ZN(U2852) );
  AOI22_X1 U7120 ( .A1(n6119), .A2(n6123), .B1(n6122), .B2(DATAI_18_), .ZN(
        n6121) );
  AOI22_X1 U7121 ( .A1(n6126), .A2(DATAI_2_), .B1(n6125), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7122 ( .A1(n6121), .A2(n6120), .ZN(U2873) );
  AOI22_X1 U7123 ( .A1(n6124), .A2(n6123), .B1(n6122), .B2(DATAI_17_), .ZN(
        n6128) );
  AOI22_X1 U7124 ( .A1(n6126), .A2(DATAI_1_), .B1(n6125), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7125 ( .A1(n6128), .A2(n6127), .ZN(U2874) );
  INV_X1 U7126 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6231) );
  AOI22_X1 U7127 ( .A1(n6609), .A2(LWORD_REG_15__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6130) );
  OAI21_X1 U7128 ( .B1(n6231), .B2(n6147), .A(n6130), .ZN(U2908) );
  INV_X1 U7129 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6225) );
  AOI22_X1 U7130 ( .A1(n6609), .A2(LWORD_REG_14__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6131) );
  OAI21_X1 U7131 ( .B1(n6225), .B2(n6147), .A(n6131), .ZN(U2909) );
  AOI22_X1 U7132 ( .A1(n6609), .A2(LWORD_REG_13__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6132) );
  OAI21_X1 U7133 ( .B1(n6222), .B2(n6147), .A(n6132), .ZN(U2910) );
  AOI22_X1 U7134 ( .A1(n6609), .A2(LWORD_REG_12__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6133) );
  OAI21_X1 U7135 ( .B1(n3696), .B2(n6147), .A(n6133), .ZN(U2911) );
  AOI22_X1 U7136 ( .A1(n6609), .A2(LWORD_REG_11__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6134) );
  OAI21_X1 U7137 ( .B1(n6217), .B2(n6147), .A(n6134), .ZN(U2912) );
  AOI22_X1 U7138 ( .A1(n6609), .A2(LWORD_REG_10__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6135) );
  OAI21_X1 U7139 ( .B1(n6214), .B2(n6147), .A(n6135), .ZN(U2913) );
  INV_X1 U7140 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6684) );
  AOI22_X1 U7141 ( .A1(n6609), .A2(LWORD_REG_9__SCAN_IN), .B1(
        DATAO_REG_9__SCAN_IN), .B2(n6145), .ZN(n6136) );
  OAI21_X1 U7142 ( .B1(n6684), .B2(n6147), .A(n6136), .ZN(U2914) );
  INV_X1 U7143 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6209) );
  AOI22_X1 U7144 ( .A1(n6609), .A2(LWORD_REG_8__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6137) );
  OAI21_X1 U7145 ( .B1(n6209), .B2(n6147), .A(n6137), .ZN(U2915) );
  INV_X1 U7146 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6206) );
  AOI22_X1 U7147 ( .A1(n6609), .A2(LWORD_REG_7__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U7148 ( .B1(n6206), .B2(n6147), .A(n6138), .ZN(U2916) );
  AOI22_X1 U7149 ( .A1(n6609), .A2(LWORD_REG_6__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6139) );
  OAI21_X1 U7150 ( .B1(n3620), .B2(n6147), .A(n6139), .ZN(U2917) );
  AOI22_X1 U7151 ( .A1(n6609), .A2(LWORD_REG_5__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7152 ( .B1(n3614), .B2(n6147), .A(n6140), .ZN(U2918) );
  AOI22_X1 U7153 ( .A1(n6609), .A2(LWORD_REG_4__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6141) );
  OAI21_X1 U7154 ( .B1(n6199), .B2(n6147), .A(n6141), .ZN(U2919) );
  AOI22_X1 U7155 ( .A1(n6609), .A2(LWORD_REG_3__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6142) );
  OAI21_X1 U7156 ( .B1(n6196), .B2(n6147), .A(n6142), .ZN(U2920) );
  AOI22_X1 U7157 ( .A1(n6609), .A2(LWORD_REG_2__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6143) );
  OAI21_X1 U7158 ( .B1(n3586), .B2(n6147), .A(n6143), .ZN(U2921) );
  AOI22_X1 U7159 ( .A1(n6609), .A2(LWORD_REG_1__SCAN_IN), .B1(
        DATAO_REG_1__SCAN_IN), .B2(n6145), .ZN(n6144) );
  OAI21_X1 U7160 ( .B1(n6191), .B2(n6147), .A(n6144), .ZN(U2922) );
  AOI22_X1 U7161 ( .A1(n6609), .A2(LWORD_REG_0__SCAN_IN), .B1(n6145), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6146) );
  OAI21_X1 U7162 ( .B1(n6188), .B2(n6147), .A(n6146), .ZN(U2923) );
  INV_X1 U7163 ( .A(n6493), .ZN(n6148) );
  NAND2_X2 U7164 ( .A1(n6149), .A2(n6148), .ZN(n6230) );
  INV_X1 U7165 ( .A(n6150), .ZN(n6151) );
  OAI21_X1 U7166 ( .B1(n6610), .B2(n6152), .A(n6151), .ZN(n6166) );
  NOR2_X1 U7167 ( .A1(n6226), .A2(n6689), .ZN(n6186) );
  AOI21_X1 U7168 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6166), .A(n6186), .ZN(n6153) );
  OAI21_X1 U7169 ( .B1(n6154), .B2(n6230), .A(n6153), .ZN(U2924) );
  NOR2_X1 U7170 ( .A1(n6226), .A2(n4653), .ZN(n6189) );
  AOI21_X1 U7171 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6166), .A(n6189), .ZN(n6155) );
  OAI21_X1 U7172 ( .B1(n6156), .B2(n6230), .A(n6155), .ZN(U2925) );
  NOR2_X1 U7173 ( .A1(n6226), .A2(n4647), .ZN(n6192) );
  AOI21_X1 U7174 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6166), .A(n6192), .ZN(n6157) );
  OAI21_X1 U7175 ( .B1(n6158), .B2(n6230), .A(n6157), .ZN(U2926) );
  NOR2_X1 U7176 ( .A1(n6226), .A2(n4651), .ZN(n6194) );
  AOI21_X1 U7177 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6166), .A(n6194), .ZN(n6159) );
  OAI21_X1 U7178 ( .B1(n6160), .B2(n6230), .A(n6159), .ZN(U2927) );
  INV_X1 U7179 ( .A(DATAI_4_), .ZN(n6161) );
  NOR2_X1 U7180 ( .A1(n6226), .A2(n6161), .ZN(n6197) );
  AOI21_X1 U7181 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6166), .A(n6197), .ZN(n6162) );
  OAI21_X1 U7182 ( .B1(n6163), .B2(n6230), .A(n6162), .ZN(U2928) );
  NOR2_X1 U7183 ( .A1(n6226), .A2(n4782), .ZN(n6200) );
  AOI21_X1 U7184 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6166), .A(n6200), .ZN(n6164) );
  OAI21_X1 U7185 ( .B1(n6165), .B2(n6230), .A(n6164), .ZN(U2929) );
  NOR2_X1 U7186 ( .A1(n6226), .A2(n4654), .ZN(n6202) );
  AOI21_X1 U7187 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6228), .A(n6202), .ZN(n6167) );
  OAI21_X1 U7188 ( .B1(n6168), .B2(n6230), .A(n6167), .ZN(U2930) );
  INV_X1 U7189 ( .A(DATAI_7_), .ZN(n6169) );
  NOR2_X1 U7190 ( .A1(n6226), .A2(n6169), .ZN(n6204) );
  AOI21_X1 U7191 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6228), .A(n6204), .ZN(n6170) );
  OAI21_X1 U7192 ( .B1(n6171), .B2(n6230), .A(n6170), .ZN(U2931) );
  INV_X1 U7193 ( .A(DATAI_8_), .ZN(n6172) );
  NOR2_X1 U7194 ( .A1(n6226), .A2(n6172), .ZN(n6207) );
  AOI21_X1 U7195 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6228), .A(n6207), .ZN(n6173) );
  OAI21_X1 U7196 ( .B1(n6174), .B2(n6230), .A(n6173), .ZN(U2932) );
  INV_X1 U7197 ( .A(DATAI_9_), .ZN(n6175) );
  NOR2_X1 U7198 ( .A1(n6226), .A2(n6175), .ZN(n6210) );
  AOI21_X1 U7199 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6228), .A(n6210), .ZN(n6176) );
  OAI21_X1 U7200 ( .B1(n6764), .B2(n6230), .A(n6176), .ZN(U2933) );
  NOR2_X1 U7201 ( .A1(n6226), .A2(n6750), .ZN(n6212) );
  AOI21_X1 U7202 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6228), .A(n6212), .ZN(
        n6177) );
  OAI21_X1 U7203 ( .B1(n3964), .B2(n6230), .A(n6177), .ZN(U2934) );
  NOR2_X1 U7204 ( .A1(n6226), .A2(n6656), .ZN(n6215) );
  AOI21_X1 U7205 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6228), .A(n6215), .ZN(
        n6178) );
  OAI21_X1 U7206 ( .B1(n6179), .B2(n6230), .A(n6178), .ZN(U2935) );
  NOR2_X1 U7207 ( .A1(n6226), .A2(n6668), .ZN(n6218) );
  AOI21_X1 U7208 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6228), .A(n6218), .ZN(
        n6180) );
  OAI21_X1 U7209 ( .B1(n4006), .B2(n6230), .A(n6180), .ZN(U2936) );
  NOR2_X1 U7210 ( .A1(n6226), .A2(n5542), .ZN(n6220) );
  AOI21_X1 U7211 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6228), .A(n6220), .ZN(
        n6181) );
  OAI21_X1 U7212 ( .B1(n6182), .B2(n6230), .A(n6181), .ZN(U2937) );
  INV_X1 U7213 ( .A(DATAI_14_), .ZN(n6183) );
  NOR2_X1 U7214 ( .A1(n6226), .A2(n6183), .ZN(n6223) );
  AOI21_X1 U7215 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6228), .A(n6223), .ZN(
        n6184) );
  OAI21_X1 U7216 ( .B1(n6185), .B2(n6230), .A(n6184), .ZN(U2938) );
  AOI21_X1 U7217 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6228), .A(n6186), .ZN(n6187) );
  OAI21_X1 U7218 ( .B1(n6188), .B2(n6230), .A(n6187), .ZN(U2939) );
  AOI21_X1 U7219 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6228), .A(n6189), .ZN(n6190) );
  OAI21_X1 U7220 ( .B1(n6191), .B2(n6230), .A(n6190), .ZN(U2940) );
  AOI21_X1 U7221 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6228), .A(n6192), .ZN(n6193) );
  OAI21_X1 U7222 ( .B1(n3586), .B2(n6230), .A(n6193), .ZN(U2941) );
  AOI21_X1 U7223 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6228), .A(n6194), .ZN(n6195) );
  OAI21_X1 U7224 ( .B1(n6196), .B2(n6230), .A(n6195), .ZN(U2942) );
  AOI21_X1 U7225 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6228), .A(n6197), .ZN(n6198) );
  OAI21_X1 U7226 ( .B1(n6199), .B2(n6230), .A(n6198), .ZN(U2943) );
  AOI21_X1 U7227 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6228), .A(n6200), .ZN(n6201) );
  OAI21_X1 U7228 ( .B1(n3614), .B2(n6230), .A(n6201), .ZN(U2944) );
  AOI21_X1 U7229 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6228), .A(n6202), .ZN(n6203) );
  OAI21_X1 U7230 ( .B1(n3620), .B2(n6230), .A(n6203), .ZN(U2945) );
  AOI21_X1 U7231 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6228), .A(n6204), .ZN(n6205) );
  OAI21_X1 U7232 ( .B1(n6206), .B2(n6230), .A(n6205), .ZN(U2946) );
  AOI21_X1 U7233 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6228), .A(n6207), .ZN(n6208) );
  OAI21_X1 U7234 ( .B1(n6209), .B2(n6230), .A(n6208), .ZN(U2947) );
  AOI21_X1 U7235 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6228), .A(n6210), .ZN(n6211) );
  OAI21_X1 U7236 ( .B1(n6684), .B2(n6230), .A(n6211), .ZN(U2948) );
  AOI21_X1 U7237 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6228), .A(n6212), .ZN(
        n6213) );
  OAI21_X1 U7238 ( .B1(n6214), .B2(n6230), .A(n6213), .ZN(U2949) );
  AOI21_X1 U7239 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6228), .A(n6215), .ZN(
        n6216) );
  OAI21_X1 U7240 ( .B1(n6217), .B2(n6230), .A(n6216), .ZN(U2950) );
  AOI21_X1 U7241 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6228), .A(n6218), .ZN(
        n6219) );
  OAI21_X1 U7242 ( .B1(n3696), .B2(n6230), .A(n6219), .ZN(U2951) );
  AOI21_X1 U7243 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6228), .A(n6220), .ZN(
        n6221) );
  OAI21_X1 U7244 ( .B1(n6222), .B2(n6230), .A(n6221), .ZN(U2952) );
  AOI21_X1 U7245 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6228), .A(n6223), .ZN(
        n6224) );
  OAI21_X1 U7246 ( .B1(n6225), .B2(n6230), .A(n6224), .ZN(U2953) );
  INV_X1 U7247 ( .A(n6226), .ZN(n6227) );
  AOI22_X1 U7248 ( .A1(n6228), .A2(LWORD_REG_15__SCAN_IN), .B1(n6227), .B2(
        DATAI_15_), .ZN(n6229) );
  OAI21_X1 U7249 ( .B1(n6231), .B2(n6230), .A(n6229), .ZN(U2954) );
  AOI22_X1 U7250 ( .A1(n6338), .A2(REIP_REG_7__SCAN_IN), .B1(n6276), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7251 ( .A1(n4913), .A2(n6232), .ZN(n6235) );
  NAND2_X1 U7252 ( .A1(n6235), .A2(n6233), .ZN(n6234) );
  OAI21_X1 U7253 ( .B1(n6235), .B2(n6233), .A(n6234), .ZN(n6236) );
  INV_X1 U7254 ( .A(n6236), .ZN(n6302) );
  AOI22_X1 U7255 ( .A1(n6302), .A2(n6257), .B1(n6258), .B2(n6237), .ZN(n6238)
         );
  OAI211_X1 U7256 ( .C1(n6264), .C2(n6240), .A(n6239), .B(n6238), .ZN(U2979)
         );
  AOI22_X1 U7257 ( .A1(n6338), .A2(REIP_REG_5__SCAN_IN), .B1(n6276), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6244) );
  AOI22_X1 U7258 ( .A1(n6242), .A2(n6257), .B1(n6258), .B2(n6241), .ZN(n6243)
         );
  OAI211_X1 U7259 ( .C1(n6264), .C2(n6245), .A(n6244), .B(n6243), .ZN(U2981)
         );
  AOI22_X1 U7260 ( .A1(n6338), .A2(REIP_REG_3__SCAN_IN), .B1(n6276), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6252) );
  OAI21_X1 U7261 ( .B1(n6248), .B2(n6247), .A(n6246), .ZN(n6249) );
  INV_X1 U7262 ( .A(n6249), .ZN(n6332) );
  AOI22_X1 U7263 ( .A1(n6250), .A2(n6258), .B1(n6332), .B2(n6257), .ZN(n6251)
         );
  OAI211_X1 U7264 ( .C1(n6264), .C2(n6253), .A(n6252), .B(n6251), .ZN(U2983)
         );
  AOI22_X1 U7265 ( .A1(n6338), .A2(REIP_REG_2__SCAN_IN), .B1(n6276), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6261) );
  XOR2_X1 U7266 ( .A(n6255), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6256) );
  XNOR2_X1 U7267 ( .A(n6254), .B(n6256), .ZN(n6345) );
  AOI22_X1 U7268 ( .A1(n6259), .A2(n6258), .B1(n6345), .B2(n6257), .ZN(n6260)
         );
  OAI211_X1 U7269 ( .C1(n6264), .C2(n6262), .A(n6261), .B(n6260), .ZN(U2984)
         );
  OAI22_X1 U7270 ( .A1(n6264), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6263), 
        .B2(n6273), .ZN(n6265) );
  AOI211_X1 U7271 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6276), .A(n6266), 
        .B(n6265), .ZN(n6267) );
  OAI21_X1 U7272 ( .B1(n6271), .B2(n6268), .A(n6267), .ZN(U2985) );
  XNOR2_X1 U7273 ( .A(n6269), .B(n6363), .ZN(n6353) );
  INV_X1 U7274 ( .A(n6353), .ZN(n6272) );
  OAI22_X1 U7275 ( .A1(n6273), .A2(n6272), .B1(n6271), .B2(n6270), .ZN(n6274)
         );
  AOI221_X1 U7276 ( .B1(n6276), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .C1(n6275), 
        .C2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n6274), .ZN(n6277) );
  NAND2_X1 U7277 ( .A1(n6338), .A2(REIP_REG_0__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U7278 ( .A1(n6277), .A2(n6351), .ZN(U2986) );
  AOI222_X1 U7279 ( .A1(n6279), .A2(n6354), .B1(n6340), .B2(n6278), .C1(
        REIP_REG_11__SCAN_IN), .C2(n6338), .ZN(n6280) );
  OAI221_X1 U7280 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6282), .C1(
        n5209), .C2(n6281), .A(n6280), .ZN(U3007) );
  AOI21_X1 U7281 ( .B1(n6340), .B2(n6284), .A(n6283), .ZN(n6288) );
  AOI22_X1 U7282 ( .A1(n6286), .A2(n6354), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6285), .ZN(n6287) );
  OAI211_X1 U7283 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6289), .A(n6288), 
        .B(n6287), .ZN(U3009) );
  INV_X1 U7284 ( .A(n6290), .ZN(n6291) );
  AOI21_X1 U7285 ( .B1(n6340), .B2(n6292), .A(n6291), .ZN(n6298) );
  INV_X1 U7286 ( .A(n6293), .ZN(n6296) );
  AOI21_X1 U7287 ( .B1(n6305), .B2(n6299), .A(n6294), .ZN(n6295) );
  AOI22_X1 U7288 ( .A1(n6296), .A2(n6354), .B1(n6301), .B2(n6295), .ZN(n6297)
         );
  OAI211_X1 U7289 ( .C1(n6306), .C2(n6299), .A(n6298), .B(n6297), .ZN(U3010)
         );
  AOI22_X1 U7290 ( .A1(n6340), .A2(n6300), .B1(n6338), .B2(REIP_REG_7__SCAN_IN), .ZN(n6304) );
  AOI22_X1 U7291 ( .A1(n6302), .A2(n6354), .B1(n6301), .B2(n6305), .ZN(n6303)
         );
  OAI211_X1 U7292 ( .C1(n6306), .C2(n6305), .A(n6304), .B(n6303), .ZN(U3011)
         );
  NAND3_X1 U7293 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6307), .A3(n6311), 
        .ZN(n6318) );
  INV_X1 U7294 ( .A(n6308), .ZN(n6309) );
  AOI21_X1 U7295 ( .B1(n6340), .B2(n6310), .A(n6309), .ZN(n6317) );
  OAI22_X1 U7296 ( .A1(n6314), .A2(n6313), .B1(n6312), .B2(n6311), .ZN(n6315)
         );
  INV_X1 U7297 ( .A(n6315), .ZN(n6316) );
  OAI211_X1 U7298 ( .C1(n6331), .C2(n6318), .A(n6317), .B(n6316), .ZN(U3012)
         );
  AOI21_X1 U7299 ( .B1(n6341), .B2(n6343), .A(n6344), .ZN(n6337) );
  INV_X1 U7300 ( .A(n6319), .ZN(n6320) );
  AOI21_X1 U7301 ( .B1(n6340), .B2(n6321), .A(n6320), .ZN(n6327) );
  AOI211_X1 U7302 ( .C1(n6336), .C2(n6328), .A(n6331), .B(n6343), .ZN(n6325)
         );
  INV_X1 U7303 ( .A(n6322), .ZN(n6323) );
  AOI22_X1 U7304 ( .A1(n6325), .A2(n6324), .B1(n6354), .B2(n6323), .ZN(n6326)
         );
  OAI211_X1 U7305 ( .C1(n6337), .C2(n6328), .A(n6327), .B(n6326), .ZN(U3014)
         );
  INV_X1 U7306 ( .A(n6329), .ZN(n6330) );
  AOI22_X1 U7307 ( .A1(n6340), .A2(n6330), .B1(n6338), .B2(REIP_REG_3__SCAN_IN), .ZN(n6335) );
  NOR2_X1 U7308 ( .A1(n6343), .A2(n6331), .ZN(n6333) );
  AOI22_X1 U7309 ( .A1(n6333), .A2(n6336), .B1(n6354), .B2(n6332), .ZN(n6334)
         );
  OAI211_X1 U7310 ( .C1(n6337), .C2(n6336), .A(n6335), .B(n6334), .ZN(U3015)
         );
  AOI22_X1 U7311 ( .A1(n6340), .A2(n6339), .B1(n6338), .B2(REIP_REG_2__SCAN_IN), .ZN(n6350) );
  OAI221_X1 U7312 ( .B1(n6343), .B2(n6342), .C1(n6343), .C2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6341), .ZN(n6349) );
  AOI22_X1 U7313 ( .A1(n6345), .A2(n6354), .B1(n6344), .B2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6348) );
  NAND3_X1 U7314 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6346), .A3(n3370), 
        .ZN(n6347) );
  NAND4_X1 U7315 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(U3016)
         );
  INV_X1 U7316 ( .A(n6351), .ZN(n6352) );
  AOI21_X1 U7317 ( .B1(n6354), .B2(n6353), .A(n6352), .ZN(n6355) );
  OAI211_X1 U7318 ( .C1(n6358), .C2(n6357), .A(n6356), .B(n6355), .ZN(n6359)
         );
  INV_X1 U7319 ( .A(n6359), .ZN(n6360) );
  OAI221_X1 U7320 ( .B1(n6363), .B2(n6362), .C1(n6363), .C2(n6361), .A(n6360), 
        .ZN(U3018) );
  NOR2_X1 U7321 ( .A1(n6365), .A2(n6364), .ZN(U3019) );
  INV_X1 U7322 ( .A(n6366), .ZN(n6377) );
  AOI22_X1 U7323 ( .A1(n6380), .A2(n6441), .B1(n6440), .B2(n6377), .ZN(n6368)
         );
  AOI22_X1 U7324 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6383), .B1(n6784), 
        .B2(n6381), .ZN(n6367) );
  OAI211_X1 U7325 ( .C1(n6387), .C2(n6786), .A(n6368), .B(n6367), .ZN(U3046)
         );
  AOI22_X1 U7326 ( .A1(n6380), .A2(n6445), .B1(n6444), .B2(n6377), .ZN(n6370)
         );
  AOI22_X1 U7327 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6383), .B1(n6446), 
        .B2(n6381), .ZN(n6369) );
  OAI211_X1 U7328 ( .C1(n6387), .C2(n6449), .A(n6370), .B(n6369), .ZN(U3047)
         );
  AOI22_X1 U7329 ( .A1(n6380), .A2(n6372), .B1(n6371), .B2(n6377), .ZN(n6374)
         );
  AOI22_X1 U7330 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6383), .B1(n6422), 
        .B2(n6381), .ZN(n6373) );
  OAI211_X1 U7331 ( .C1(n6387), .C2(n6427), .A(n6374), .B(n6373), .ZN(U3048)
         );
  AOI22_X1 U7332 ( .A1(n6380), .A2(n6451), .B1(n6450), .B2(n6377), .ZN(n6376)
         );
  AOI22_X1 U7333 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6383), .B1(n6452), 
        .B2(n6381), .ZN(n6375) );
  OAI211_X1 U7334 ( .C1(n6387), .C2(n6455), .A(n6376), .B(n6375), .ZN(U3049)
         );
  AOI22_X1 U7335 ( .A1(n6380), .A2(n6379), .B1(n6378), .B2(n6377), .ZN(n6385)
         );
  AOI22_X1 U7336 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6383), .B1(n6382), 
        .B2(n6381), .ZN(n6384) );
  OAI211_X1 U7337 ( .C1(n6387), .C2(n6386), .A(n6385), .B(n6384), .ZN(U3050)
         );
  INV_X1 U7338 ( .A(n6388), .ZN(n6400) );
  AOI22_X1 U7339 ( .A1(n6430), .A2(n6400), .B1(n6428), .B2(n6399), .ZN(n6391)
         );
  AOI22_X1 U7340 ( .A1(n6403), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6389), 
        .B2(n6401), .ZN(n6390) );
  OAI211_X1 U7341 ( .C1(n6407), .C2(n6426), .A(n6391), .B(n6390), .ZN(U3068)
         );
  AOI22_X1 U7342 ( .A1(n6436), .A2(n6400), .B1(n6434), .B2(n6399), .ZN(n6394)
         );
  AOI22_X1 U7343 ( .A1(n6403), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6392), 
        .B2(n6401), .ZN(n6393) );
  OAI211_X1 U7344 ( .C1(n6395), .C2(n6426), .A(n6394), .B(n6393), .ZN(U3069)
         );
  AOI22_X1 U7345 ( .A1(n6784), .A2(n6400), .B1(n6440), .B2(n6399), .ZN(n6398)
         );
  AOI22_X1 U7346 ( .A1(n6403), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6396), 
        .B2(n6401), .ZN(n6397) );
  OAI211_X1 U7347 ( .C1(n6794), .C2(n6426), .A(n6398), .B(n6397), .ZN(U3070)
         );
  AOI22_X1 U7348 ( .A1(n6446), .A2(n6400), .B1(n6444), .B2(n6399), .ZN(n6405)
         );
  AOI22_X1 U7349 ( .A1(n6403), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6402), 
        .B2(n6401), .ZN(n6404) );
  OAI211_X1 U7350 ( .C1(n6412), .C2(n6426), .A(n6405), .B(n6404), .ZN(U3071)
         );
  OAI22_X1 U7351 ( .A1(n6419), .A2(n6407), .B1(n6417), .B2(n6406), .ZN(n6408)
         );
  INV_X1 U7352 ( .A(n6408), .ZN(n6410) );
  AOI22_X1 U7353 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6423), .B1(n6430), 
        .B2(n6421), .ZN(n6409) );
  OAI211_X1 U7354 ( .C1(n6433), .C2(n6426), .A(n6410), .B(n6409), .ZN(U3076)
         );
  OAI22_X1 U7355 ( .A1(n6419), .A2(n6412), .B1(n6417), .B2(n6411), .ZN(n6413)
         );
  INV_X1 U7356 ( .A(n6413), .ZN(n6415) );
  AOI22_X1 U7357 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6423), .B1(n6446), 
        .B2(n6421), .ZN(n6414) );
  OAI211_X1 U7358 ( .C1(n6449), .C2(n6426), .A(n6415), .B(n6414), .ZN(U3079)
         );
  OAI22_X1 U7359 ( .A1(n6419), .A2(n6418), .B1(n6417), .B2(n6416), .ZN(n6420)
         );
  INV_X1 U7360 ( .A(n6420), .ZN(n6425) );
  AOI22_X1 U7361 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6423), .B1(n6422), 
        .B2(n6421), .ZN(n6424) );
  OAI211_X1 U7362 ( .C1(n6427), .C2(n6426), .A(n6425), .B(n6424), .ZN(U3080)
         );
  AOI22_X1 U7363 ( .A1(n6459), .A2(n6429), .B1(n6428), .B2(n6456), .ZN(n6432)
         );
  AOI22_X1 U7364 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6462), .B1(n6430), 
        .B2(n6460), .ZN(n6431) );
  OAI211_X1 U7365 ( .C1(n6433), .C2(n6465), .A(n6432), .B(n6431), .ZN(U3108)
         );
  AOI22_X1 U7366 ( .A1(n6459), .A2(n6435), .B1(n6434), .B2(n6456), .ZN(n6438)
         );
  AOI22_X1 U7367 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6462), .B1(n6436), 
        .B2(n6460), .ZN(n6437) );
  OAI211_X1 U7368 ( .C1(n6439), .C2(n6465), .A(n6438), .B(n6437), .ZN(U3109)
         );
  AOI22_X1 U7369 ( .A1(n6459), .A2(n6441), .B1(n6440), .B2(n6456), .ZN(n6443)
         );
  AOI22_X1 U7370 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6462), .B1(n6784), 
        .B2(n6460), .ZN(n6442) );
  OAI211_X1 U7371 ( .C1(n6786), .C2(n6465), .A(n6443), .B(n6442), .ZN(U3110)
         );
  AOI22_X1 U7372 ( .A1(n6459), .A2(n6445), .B1(n6444), .B2(n6456), .ZN(n6448)
         );
  AOI22_X1 U7373 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6462), .B1(n6446), 
        .B2(n6460), .ZN(n6447) );
  OAI211_X1 U7374 ( .C1(n6449), .C2(n6465), .A(n6448), .B(n6447), .ZN(U3111)
         );
  AOI22_X1 U7375 ( .A1(n6459), .A2(n6451), .B1(n6450), .B2(n6456), .ZN(n6454)
         );
  AOI22_X1 U7376 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6462), .B1(n6452), 
        .B2(n6460), .ZN(n6453) );
  OAI211_X1 U7377 ( .C1(n6455), .C2(n6465), .A(n6454), .B(n6453), .ZN(U3113)
         );
  AOI22_X1 U7378 ( .A1(n6459), .A2(n6458), .B1(n6457), .B2(n6456), .ZN(n6464)
         );
  AOI22_X1 U7379 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6462), .B1(n6461), 
        .B2(n6460), .ZN(n6463) );
  OAI211_X1 U7380 ( .C1(n6466), .C2(n6465), .A(n6464), .B(n6463), .ZN(U3115)
         );
  AOI22_X1 U7381 ( .A1(n2985), .A2(n6468), .B1(n6467), .B2(n3034), .ZN(n6590)
         );
  NAND2_X1 U7382 ( .A1(n6469), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6598) );
  AND3_X1 U7383 ( .A1(n6590), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6598), 
        .ZN(n6475) );
  INV_X1 U7384 ( .A(n6470), .ZN(n6471) );
  AOI21_X1 U7385 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6475), .A(n6471), 
        .ZN(n6472) );
  NAND2_X1 U7386 ( .A1(n6473), .A2(n6472), .ZN(n6474) );
  OAI21_X1 U7387 ( .B1(n6475), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6474), 
        .ZN(n6476) );
  AOI222_X1 U7388 ( .A1(n6478), .A2(n6477), .B1(n6478), .B2(n6476), .C1(n6477), 
        .C2(n6476), .ZN(n6482) );
  INV_X1 U7389 ( .A(n6482), .ZN(n6480) );
  AOI21_X1 U7390 ( .B1(n6480), .B2(n6768), .A(n6479), .ZN(n6481) );
  AOI211_X1 U7391 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6482), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n6481), .ZN(n6489) );
  OAI21_X1 U7392 ( .B1(MORE_REG_SCAN_IN), .B2(FLUSH_REG_SCAN_IN), .A(n6483), 
        .ZN(n6486) );
  NAND3_X1 U7393 ( .A1(n6486), .A2(n6485), .A3(n6484), .ZN(n6487) );
  NOR3_X1 U7394 ( .A1(n6489), .A2(n6488), .A3(n6487), .ZN(n6500) );
  AOI22_X1 U7395 ( .A1(n6500), .A2(n6490), .B1(READY_N), .B2(n6609), .ZN(n6491) );
  INV_X1 U7396 ( .A(n6491), .ZN(n6492) );
  OAI21_X1 U7397 ( .B1(n6494), .B2(n6493), .A(n6492), .ZN(n6588) );
  OAI21_X1 U7398 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6610), .A(n6588), .ZN(
        n6501) );
  AOI221_X1 U7399 ( .B1(n6496), .B2(STATE2_REG_0__SCAN_IN), .C1(n6501), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6495), .ZN(n6499) );
  OAI211_X1 U7400 ( .C1(n6508), .C2(n6497), .A(n6669), .B(n6588), .ZN(n6498)
         );
  OAI211_X1 U7401 ( .C1(n6500), .C2(n6502), .A(n6499), .B(n6498), .ZN(U3148)
         );
  NOR2_X1 U7402 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6511) );
  NAND2_X1 U7403 ( .A1(n6501), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6507) );
  OAI21_X1 U7404 ( .B1(READY_N), .B2(n6503), .A(n6502), .ZN(n6505) );
  AOI21_X1 U7405 ( .B1(n6588), .B2(n6505), .A(n6504), .ZN(n6506) );
  OAI21_X1 U7406 ( .B1(n6511), .B2(n6507), .A(n6506), .ZN(U3149) );
  OAI211_X1 U7407 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6610), .A(n6586), .B(
        n6508), .ZN(n6510) );
  OAI21_X1 U7408 ( .B1(n6511), .B2(n6510), .A(n6509), .ZN(U3150) );
  INV_X1 U7409 ( .A(n6585), .ZN(n6581) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6581), .ZN(U3151) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6581), .ZN(U3152) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6581), .ZN(U3153) );
  AND2_X1 U7413 ( .A1(n6581), .A2(DATAWIDTH_REG_28__SCAN_IN), .ZN(U3154) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6581), .ZN(U3155) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6581), .ZN(U3156) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6581), .ZN(U3157) );
  AND2_X1 U7417 ( .A1(n6581), .A2(DATAWIDTH_REG_24__SCAN_IN), .ZN(U3158) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6581), .ZN(U3159) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6581), .ZN(U3160) );
  AND2_X1 U7420 ( .A1(n6581), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6581), .ZN(U3162) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6581), .ZN(U3163) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6581), .ZN(U3164) );
  AND2_X1 U7424 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6581), .ZN(U3165) );
  AND2_X1 U7425 ( .A1(n6581), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  AND2_X1 U7426 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6581), .ZN(U3167) );
  AND2_X1 U7427 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6581), .ZN(U3168) );
  AND2_X1 U7428 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6581), .ZN(U3169) );
  AND2_X1 U7429 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6581), .ZN(U3170) );
  AND2_X1 U7430 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6581), .ZN(U3171) );
  AND2_X1 U7431 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6581), .ZN(U3172) );
  AND2_X1 U7432 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6581), .ZN(U3173) );
  AND2_X1 U7433 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6581), .ZN(U3174) );
  AND2_X1 U7434 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6581), .ZN(U3175) );
  AND2_X1 U7435 ( .A1(n6581), .A2(DATAWIDTH_REG_6__SCAN_IN), .ZN(U3176) );
  AND2_X1 U7436 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6581), .ZN(U3177) );
  AND2_X1 U7437 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6581), .ZN(U3178) );
  AND2_X1 U7438 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6581), .ZN(U3179) );
  AND2_X1 U7439 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6581), .ZN(U3180) );
  NOR2_X1 U7440 ( .A1(n6518), .A2(n6528), .ZN(n6521) );
  AOI22_X1 U7441 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6525) );
  AND2_X1 U7442 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6515) );
  INV_X1 U7443 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6513) );
  INV_X1 U7444 ( .A(NA_N), .ZN(n6522) );
  AOI211_X1 U7445 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6522), .A(
        STATE_REG_0__SCAN_IN), .B(n6521), .ZN(n6527) );
  AOI221_X1 U7446 ( .B1(n6515), .B2(n6608), .C1(n6513), .C2(n6608), .A(n6527), 
        .ZN(n6512) );
  OAI21_X1 U7447 ( .B1(n6521), .B2(n6525), .A(n6512), .ZN(U3181) );
  NOR2_X1 U7448 ( .A1(n6519), .A2(n6513), .ZN(n6523) );
  NAND2_X1 U7449 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6514) );
  OAI21_X1 U7450 ( .B1(n6523), .B2(n6515), .A(n6514), .ZN(n6516) );
  OAI211_X1 U7451 ( .C1(n6518), .C2(n6610), .A(n6517), .B(n6516), .ZN(U3182)
         );
  AOI221_X1 U7452 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6610), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6520) );
  AOI221_X1 U7453 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6520), .C2(HOLD), .A(n6519), .ZN(n6526) );
  AOI21_X1 U7454 ( .B1(n6523), .B2(n6522), .A(n6521), .ZN(n6524) );
  OAI22_X1 U7455 ( .A1(n6527), .A2(n6526), .B1(n6525), .B2(n6524), .ZN(U3183)
         );
  NAND2_X1 U7456 ( .A1(n6622), .A2(n6528), .ZN(n6579) );
  INV_X1 U7457 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U7458 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6622), .ZN(n6576) );
  OAI222_X1 U7459 ( .A1(n6579), .A2(n6531), .B1(n6529), .B2(n6622), .C1(n6599), 
        .C2(n6576), .ZN(U3184) );
  INV_X1 U7460 ( .A(n6579), .ZN(n6567) );
  AOI22_X1 U7461 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6608), .ZN(n6530) );
  OAI21_X1 U7462 ( .B1(n6531), .B2(n6576), .A(n6530), .ZN(U3185) );
  INV_X1 U7463 ( .A(n6576), .ZN(n6577) );
  AOI22_X1 U7464 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6608), .ZN(n6532) );
  OAI21_X1 U7465 ( .B1(n6534), .B2(n6579), .A(n6532), .ZN(U3186) );
  AOI22_X1 U7466 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6608), .ZN(n6533) );
  OAI21_X1 U7467 ( .B1(n6534), .B2(n6576), .A(n6533), .ZN(U3187) );
  AOI22_X1 U7468 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6608), .ZN(n6535) );
  OAI21_X1 U7469 ( .B1(n6536), .B2(n6579), .A(n6535), .ZN(U3188) );
  AOI22_X1 U7470 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6608), .ZN(n6537) );
  OAI21_X1 U7471 ( .B1(n6538), .B2(n6579), .A(n6537), .ZN(U3189) );
  AOI22_X1 U7472 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6608), .ZN(n6539) );
  OAI21_X1 U7473 ( .B1(n6541), .B2(n6579), .A(n6539), .ZN(U3190) );
  AOI22_X1 U7474 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6608), .ZN(n6540) );
  OAI21_X1 U7475 ( .B1(n6541), .B2(n6576), .A(n6540), .ZN(U3191) );
  AOI22_X1 U7476 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6608), .ZN(n6542) );
  OAI21_X1 U7477 ( .B1(n6543), .B2(n6576), .A(n6542), .ZN(U3192) );
  AOI22_X1 U7478 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6608), .ZN(n6544) );
  OAI21_X1 U7479 ( .B1(n6546), .B2(n6579), .A(n6544), .ZN(U3193) );
  INV_X1 U7480 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6545) );
  OAI222_X1 U7481 ( .A1(n6576), .A2(n6546), .B1(n6545), .B2(n6622), .C1(n5244), 
        .C2(n6579), .ZN(U3194) );
  INV_X1 U7482 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6547) );
  OAI222_X1 U7483 ( .A1(n6579), .A2(n6548), .B1(n6547), .B2(n6622), .C1(n5244), 
        .C2(n6576), .ZN(U3195) );
  AOI22_X1 U7484 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6608), .ZN(n6549) );
  OAI21_X1 U7485 ( .B1(n6728), .B2(n6579), .A(n6549), .ZN(U3196) );
  AOI22_X1 U7486 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6608), .ZN(n6550) );
  OAI21_X1 U7487 ( .B1(n6552), .B2(n6579), .A(n6550), .ZN(U3197) );
  AOI22_X1 U7488 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6608), .ZN(n6551) );
  OAI21_X1 U7489 ( .B1(n6552), .B2(n6576), .A(n6551), .ZN(U3198) );
  AOI22_X1 U7490 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6608), .ZN(n6553) );
  OAI21_X1 U7491 ( .B1(n5644), .B2(n6576), .A(n6553), .ZN(U3199) );
  AOI22_X1 U7492 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6608), .ZN(n6554) );
  OAI21_X1 U7493 ( .B1(n6705), .B2(n6579), .A(n6554), .ZN(U3200) );
  AOI22_X1 U7494 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6608), .ZN(n6555) );
  OAI21_X1 U7495 ( .B1(n6705), .B2(n6576), .A(n6555), .ZN(U3201) );
  INV_X1 U7496 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6557) );
  AOI22_X1 U7497 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6608), .ZN(n6556) );
  OAI21_X1 U7498 ( .B1(n6557), .B2(n6576), .A(n6556), .ZN(U3202) );
  AOI22_X1 U7499 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6608), .ZN(n6558) );
  OAI21_X1 U7500 ( .B1(n6560), .B2(n6579), .A(n6558), .ZN(U3203) );
  AOI22_X1 U7501 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6608), .ZN(n6559) );
  OAI21_X1 U7502 ( .B1(n6560), .B2(n6576), .A(n6559), .ZN(U3204) );
  AOI22_X1 U7503 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6608), .ZN(n6561) );
  OAI21_X1 U7504 ( .B1(n6563), .B2(n6579), .A(n6561), .ZN(U3205) );
  AOI22_X1 U7505 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6608), .ZN(n6562) );
  OAI21_X1 U7506 ( .B1(n6563), .B2(n6576), .A(n6562), .ZN(U3206) );
  AOI22_X1 U7507 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6608), .ZN(n6564) );
  OAI21_X1 U7508 ( .B1(n6565), .B2(n6576), .A(n6564), .ZN(U3207) );
  AOI22_X1 U7509 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6608), .ZN(n6566) );
  OAI21_X1 U7510 ( .B1(n6569), .B2(n6579), .A(n6566), .ZN(U3208) );
  AOI22_X1 U7511 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6567), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6608), .ZN(n6568) );
  OAI21_X1 U7512 ( .B1(n6569), .B2(n6576), .A(n6568), .ZN(U3209) );
  AOI22_X1 U7513 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6608), .ZN(n6570) );
  OAI21_X1 U7514 ( .B1(n6572), .B2(n6579), .A(n6570), .ZN(U3210) );
  INV_X1 U7515 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6571) );
  OAI222_X1 U7516 ( .A1(n6576), .A2(n6572), .B1(n6571), .B2(n6622), .C1(n6575), 
        .C2(n6579), .ZN(U3211) );
  INV_X1 U7517 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6574) );
  OAI222_X1 U7518 ( .A1(n6576), .A2(n6575), .B1(n6574), .B2(n6622), .C1(n6573), 
        .C2(n6579), .ZN(U3212) );
  AOI22_X1 U7519 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6577), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6608), .ZN(n6578) );
  OAI21_X1 U7520 ( .B1(n6701), .B2(n6579), .A(n6578), .ZN(U3213) );
  MUX2_X1 U7521 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6622), .Z(U3445) );
  MUX2_X1 U7522 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6622), .Z(U3446) );
  MUX2_X1 U7523 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6622), .Z(U3447) );
  MUX2_X1 U7524 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6622), .Z(U3448) );
  INV_X1 U7525 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6582) );
  INV_X1 U7526 ( .A(n6583), .ZN(n6580) );
  AOI21_X1 U7527 ( .B1(n6582), .B2(n6581), .A(n6580), .ZN(U3451) );
  OAI21_X1 U7528 ( .B1(n6585), .B2(n6584), .A(n6583), .ZN(U3452) );
  OAI211_X1 U7529 ( .C1(n6589), .C2(n6588), .A(n6587), .B(n6586), .ZN(U3453)
         );
  OR2_X1 U7530 ( .A1(n6590), .A2(n6597), .ZN(n6591) );
  OAI21_X1 U7531 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6592), .A(n6591), 
        .ZN(n6595) );
  OAI22_X1 U7532 ( .A1(n6595), .A2(n6594), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6593), .ZN(n6596) );
  OAI21_X1 U7533 ( .B1(n6598), .B2(n6597), .A(n6596), .ZN(U3461) );
  AOI21_X1 U7534 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6600) );
  AOI22_X1 U7535 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6600), .B2(n6599), .ZN(n6603) );
  INV_X1 U7536 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6602) );
  AOI22_X1 U7537 ( .A1(n6606), .A2(n6603), .B1(n6602), .B2(n6601), .ZN(U3468)
         );
  INV_X1 U7538 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6605) );
  OAI21_X1 U7539 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6606), .ZN(n6604) );
  OAI21_X1 U7540 ( .B1(n6606), .B2(n6605), .A(n6604), .ZN(U3469) );
  NAND2_X1 U7541 ( .A1(n6608), .A2(W_R_N_REG_SCAN_IN), .ZN(n6607) );
  OAI21_X1 U7542 ( .B1(n6608), .B2(READREQUEST_REG_SCAN_IN), .A(n6607), .ZN(
        U3470) );
  AND2_X1 U7543 ( .A1(n6610), .A2(n6609), .ZN(n6611) );
  NOR4_X1 U7544 ( .A1(n6614), .A2(n6613), .A3(n6612), .A4(n6611), .ZN(n6621)
         );
  OAI211_X1 U7545 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6616), .A(n6615), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6618) );
  AOI21_X1 U7546 ( .B1(n6618), .B2(STATE2_REG_0__SCAN_IN), .A(n6617), .ZN(
        n6620) );
  NAND2_X1 U7547 ( .A1(n6621), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6619) );
  OAI21_X1 U7548 ( .B1(n6621), .B2(n6620), .A(n6619), .ZN(U3472) );
  MUX2_X1 U7549 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6622), .Z(U3473) );
  NOR2_X1 U7550 ( .A1(keyinput26), .A2(keyinput30), .ZN(n6628) );
  NAND2_X1 U7551 ( .A1(keyinput47), .A2(keyinput15), .ZN(n6626) );
  NOR4_X1 U7552 ( .A1(keyinput37), .A2(keyinput61), .A3(keyinput45), .A4(
        keyinput33), .ZN(n6624) );
  NOR2_X1 U7553 ( .A1(keyinput23), .A2(keyinput42), .ZN(n6623) );
  NAND4_X1 U7554 ( .A1(n6624), .A2(keyinput39), .A3(keyinput50), .A4(n6623), 
        .ZN(n6625) );
  NOR4_X1 U7555 ( .A1(keyinput62), .A2(keyinput24), .A3(n6626), .A4(n6625), 
        .ZN(n6627) );
  NAND4_X1 U7556 ( .A1(keyinput1), .A2(keyinput22), .A3(n6628), .A4(n6627), 
        .ZN(n6650) );
  NAND2_X1 U7557 ( .A1(keyinput40), .A2(keyinput7), .ZN(n6629) );
  NOR3_X1 U7558 ( .A1(keyinput54), .A2(keyinput55), .A3(n6629), .ZN(n6648) );
  NOR4_X1 U7559 ( .A1(keyinput6), .A2(keyinput46), .A3(keyinput16), .A4(
        keyinput32), .ZN(n6647) );
  NAND4_X1 U7560 ( .A1(keyinput9), .A2(keyinput17), .A3(keyinput49), .A4(
        keyinput3), .ZN(n6631) );
  NAND2_X1 U7561 ( .A1(keyinput29), .A2(keyinput60), .ZN(n6630) );
  NOR4_X1 U7562 ( .A1(keyinput27), .A2(keyinput13), .A3(n6631), .A4(n6630), 
        .ZN(n6646) );
  NAND3_X1 U7563 ( .A1(keyinput41), .A2(keyinput58), .A3(keyinput63), .ZN(
        n6644) );
  INV_X1 U7564 ( .A(keyinput43), .ZN(n6635) );
  NOR3_X1 U7565 ( .A1(keyinput25), .A2(keyinput36), .A3(keyinput44), .ZN(n6633) );
  NOR3_X1 U7566 ( .A1(keyinput38), .A2(keyinput12), .A3(keyinput2), .ZN(n6632)
         );
  NAND4_X1 U7567 ( .A1(keyinput8), .A2(n6633), .A3(keyinput51), .A4(n6632), 
        .ZN(n6634) );
  OR4_X1 U7568 ( .A1(keyinput56), .A2(keyinput53), .A3(n6635), .A4(n6634), 
        .ZN(n6643) );
  NOR2_X1 U7569 ( .A1(keyinput48), .A2(keyinput20), .ZN(n6641) );
  NAND2_X1 U7570 ( .A1(keyinput59), .A2(keyinput14), .ZN(n6639) );
  NOR4_X1 U7571 ( .A1(keyinput35), .A2(keyinput5), .A3(keyinput31), .A4(
        keyinput57), .ZN(n6637) );
  NOR2_X1 U7572 ( .A1(keyinput34), .A2(keyinput10), .ZN(n6636) );
  NAND4_X1 U7573 ( .A1(n6637), .A2(keyinput0), .A3(keyinput19), .A4(n6636), 
        .ZN(n6638) );
  NOR4_X1 U7574 ( .A1(keyinput4), .A2(keyinput52), .A3(n6639), .A4(n6638), 
        .ZN(n6640) );
  NAND4_X1 U7575 ( .A1(keyinput28), .A2(keyinput21), .A3(n6641), .A4(n6640), 
        .ZN(n6642) );
  NOR4_X1 U7576 ( .A1(keyinput18), .A2(n6644), .A3(n6643), .A4(n6642), .ZN(
        n6645) );
  NAND4_X1 U7577 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n6649)
         );
  OAI21_X1 U7578 ( .B1(n6650), .B2(n6649), .A(keyinput11), .ZN(n6782) );
  INV_X1 U7579 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6651) );
  AOI22_X1 U7580 ( .A1(keyinput56), .A2(n6653), .B1(keyinput11), .B2(n6651), 
        .ZN(n6652) );
  OAI21_X1 U7581 ( .B1(n6653), .B2(keyinput56), .A(n6652), .ZN(n6666) );
  INV_X1 U7582 ( .A(keyinput53), .ZN(n6655) );
  AOI22_X1 U7583 ( .A1(n6656), .A2(keyinput25), .B1(DATAWIDTH_REG_21__SCAN_IN), 
        .B2(n6655), .ZN(n6654) );
  OAI221_X1 U7584 ( .B1(n6656), .B2(keyinput25), .C1(n6655), .C2(
        DATAWIDTH_REG_21__SCAN_IN), .A(n6654), .ZN(n6665) );
  INV_X1 U7585 ( .A(keyinput8), .ZN(n6658) );
  AOI22_X1 U7586 ( .A1(n6659), .A2(keyinput36), .B1(DATAWIDTH_REG_28__SCAN_IN), 
        .B2(n6658), .ZN(n6657) );
  OAI221_X1 U7587 ( .B1(n6659), .B2(keyinput36), .C1(n6658), .C2(
        DATAWIDTH_REG_28__SCAN_IN), .A(n6657), .ZN(n6664) );
  INV_X1 U7588 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6662) );
  AOI22_X1 U7589 ( .A1(n6662), .A2(keyinput44), .B1(keyinput38), .B2(n6661), 
        .ZN(n6660) );
  OAI221_X1 U7590 ( .B1(n6662), .B2(keyinput44), .C1(n6661), .C2(keyinput38), 
        .A(n6660), .ZN(n6663) );
  NOR4_X1 U7591 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n6716)
         );
  AOI22_X1 U7592 ( .A1(n6669), .A2(keyinput58), .B1(keyinput18), .B2(n6668), 
        .ZN(n6667) );
  OAI221_X1 U7593 ( .B1(n6669), .B2(keyinput58), .C1(n6668), .C2(keyinput18), 
        .A(n6667), .ZN(n6681) );
  INV_X1 U7594 ( .A(DATAI_26_), .ZN(n6672) );
  AOI22_X1 U7595 ( .A1(n6672), .A2(keyinput12), .B1(n6671), .B2(keyinput51), 
        .ZN(n6670) );
  OAI221_X1 U7596 ( .B1(n6672), .B2(keyinput12), .C1(n6671), .C2(keyinput51), 
        .A(n6670), .ZN(n6680) );
  INV_X1 U7597 ( .A(keyinput41), .ZN(n6674) );
  AOI22_X1 U7598 ( .A1(n6675), .A2(keyinput2), .B1(LWORD_REG_11__SCAN_IN), 
        .B2(n6674), .ZN(n6673) );
  OAI221_X1 U7599 ( .B1(n6675), .B2(keyinput2), .C1(n6674), .C2(
        LWORD_REG_11__SCAN_IN), .A(n6673), .ZN(n6679) );
  XNOR2_X1 U7600 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(keyinput1), .ZN(
        n6677) );
  XNOR2_X1 U7601 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput63), .ZN(
        n6676) );
  NAND2_X1 U7602 ( .A1(n6677), .A2(n6676), .ZN(n6678) );
  NOR4_X1 U7603 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6715)
         );
  INV_X1 U7604 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U7605 ( .A1(n6684), .A2(keyinput26), .B1(n6683), .B2(keyinput22), 
        .ZN(n6682) );
  OAI221_X1 U7606 ( .B1(n6684), .B2(keyinput26), .C1(n6683), .C2(keyinput22), 
        .A(n6682), .ZN(n6696) );
  INV_X1 U7607 ( .A(keyinput30), .ZN(n6686) );
  AOI22_X1 U7608 ( .A1(n5519), .A2(keyinput37), .B1(DATAWIDTH_REG_6__SCAN_IN), 
        .B2(n6686), .ZN(n6685) );
  OAI221_X1 U7609 ( .B1(n5519), .B2(keyinput37), .C1(n6686), .C2(
        DATAWIDTH_REG_6__SCAN_IN), .A(n6685), .ZN(n6695) );
  INV_X1 U7610 ( .A(keyinput61), .ZN(n6688) );
  AOI22_X1 U7611 ( .A1(n6689), .A2(keyinput45), .B1(DATAO_REG_1__SCAN_IN), 
        .B2(n6688), .ZN(n6687) );
  OAI221_X1 U7612 ( .B1(n6689), .B2(keyinput45), .C1(n6688), .C2(
        DATAO_REG_1__SCAN_IN), .A(n6687), .ZN(n6694) );
  INV_X1 U7613 ( .A(keyinput33), .ZN(n6691) );
  AOI22_X1 U7614 ( .A1(n6692), .A2(keyinput62), .B1(DATAO_REG_23__SCAN_IN), 
        .B2(n6691), .ZN(n6690) );
  OAI221_X1 U7615 ( .B1(n6692), .B2(keyinput62), .C1(n6691), .C2(
        DATAO_REG_23__SCAN_IN), .A(n6690), .ZN(n6693) );
  NOR4_X1 U7616 ( .A1(n6696), .A2(n6695), .A3(n6694), .A4(n6693), .ZN(n6714)
         );
  INV_X1 U7617 ( .A(keyinput47), .ZN(n6699) );
  INV_X1 U7618 ( .A(keyinput24), .ZN(n6698) );
  AOI22_X1 U7619 ( .A1(n6699), .A2(ADDRESS_REG_4__SCAN_IN), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6698), .ZN(n6697) );
  OAI221_X1 U7620 ( .B1(n6699), .B2(ADDRESS_REG_4__SCAN_IN), .C1(n6698), .C2(
        ADDRESS_REG_27__SCAN_IN), .A(n6697), .ZN(n6712) );
  INV_X1 U7621 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6702) );
  AOI22_X1 U7622 ( .A1(n6702), .A2(keyinput15), .B1(keyinput39), .B2(n6701), 
        .ZN(n6700) );
  OAI221_X1 U7623 ( .B1(n6702), .B2(keyinput15), .C1(n6701), .C2(keyinput39), 
        .A(n6700), .ZN(n6711) );
  INV_X1 U7624 ( .A(DATAI_19_), .ZN(n6704) );
  AOI22_X1 U7625 ( .A1(n6705), .A2(keyinput23), .B1(keyinput50), .B2(n6704), 
        .ZN(n6703) );
  OAI221_X1 U7626 ( .B1(n6705), .B2(keyinput23), .C1(n6704), .C2(keyinput50), 
        .A(n6703), .ZN(n6710) );
  INV_X1 U7627 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6708) );
  INV_X1 U7628 ( .A(keyinput28), .ZN(n6707) );
  AOI22_X1 U7629 ( .A1(n6708), .A2(keyinput42), .B1(UWORD_REG_10__SCAN_IN), 
        .B2(n6707), .ZN(n6706) );
  OAI221_X1 U7630 ( .B1(n6708), .B2(keyinput42), .C1(n6707), .C2(
        UWORD_REG_10__SCAN_IN), .A(n6706), .ZN(n6709) );
  NOR4_X1 U7631 ( .A1(n6712), .A2(n6711), .A3(n6710), .A4(n6709), .ZN(n6713)
         );
  NAND4_X1 U7632 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n6781)
         );
  INV_X1 U7633 ( .A(DATAI_25_), .ZN(n6719) );
  INV_X1 U7634 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6718) );
  AOI22_X1 U7635 ( .A1(n6719), .A2(keyinput57), .B1(n6718), .B2(keyinput0), 
        .ZN(n6717) );
  OAI221_X1 U7636 ( .B1(n6719), .B2(keyinput57), .C1(n6718), .C2(keyinput0), 
        .A(n6717), .ZN(n6732) );
  INV_X1 U7637 ( .A(keyinput31), .ZN(n6721) );
  AOI22_X1 U7638 ( .A1(n6722), .A2(keyinput5), .B1(DATAO_REG_9__SCAN_IN), .B2(
        n6721), .ZN(n6720) );
  OAI221_X1 U7639 ( .B1(n6722), .B2(keyinput5), .C1(n6721), .C2(
        DATAO_REG_9__SCAN_IN), .A(n6720), .ZN(n6731) );
  INV_X1 U7640 ( .A(DATAI_31_), .ZN(n6725) );
  INV_X1 U7641 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6724) );
  AOI22_X1 U7642 ( .A1(n6725), .A2(keyinput10), .B1(n6724), .B2(keyinput9), 
        .ZN(n6723) );
  OAI221_X1 U7643 ( .B1(n6725), .B2(keyinput10), .C1(n6724), .C2(keyinput9), 
        .A(n6723), .ZN(n6730) );
  INV_X1 U7644 ( .A(keyinput34), .ZN(n6727) );
  AOI22_X1 U7645 ( .A1(n6728), .A2(keyinput19), .B1(ADDRESS_REG_3__SCAN_IN), 
        .B2(n6727), .ZN(n6726) );
  OAI221_X1 U7646 ( .B1(n6728), .B2(keyinput19), .C1(n6727), .C2(
        ADDRESS_REG_3__SCAN_IN), .A(n6726), .ZN(n6729) );
  NOR4_X1 U7647 ( .A1(n6732), .A2(n6731), .A3(n6730), .A4(n6729), .ZN(n6779)
         );
  INV_X1 U7648 ( .A(keyinput14), .ZN(n6734) );
  AOI22_X1 U7649 ( .A1(n6735), .A2(keyinput59), .B1(ADDRESS_REG_11__SCAN_IN), 
        .B2(n6734), .ZN(n6733) );
  OAI221_X1 U7650 ( .B1(n6735), .B2(keyinput59), .C1(n6734), .C2(
        ADDRESS_REG_11__SCAN_IN), .A(n6733), .ZN(n6747) );
  INV_X1 U7651 ( .A(keyinput35), .ZN(n6737) );
  AOI22_X1 U7652 ( .A1(n6738), .A2(keyinput52), .B1(DATAWIDTH_REG_16__SCAN_IN), 
        .B2(n6737), .ZN(n6736) );
  OAI221_X1 U7653 ( .B1(n6738), .B2(keyinput52), .C1(n6737), .C2(
        DATAWIDTH_REG_16__SCAN_IN), .A(n6736), .ZN(n6746) );
  INV_X1 U7654 ( .A(keyinput4), .ZN(n6740) );
  AOI22_X1 U7655 ( .A1(n6741), .A2(keyinput20), .B1(ADDRESS_REG_0__SCAN_IN), 
        .B2(n6740), .ZN(n6739) );
  OAI221_X1 U7656 ( .B1(n6741), .B2(keyinput20), .C1(n6740), .C2(
        ADDRESS_REG_0__SCAN_IN), .A(n6739), .ZN(n6745) );
  XNOR2_X1 U7657 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(keyinput48), .ZN(
        n6743) );
  XNOR2_X1 U7658 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .B(keyinput21), .ZN(n6742)
         );
  NAND2_X1 U7659 ( .A1(n6743), .A2(n6742), .ZN(n6744) );
  NOR4_X1 U7660 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6778)
         );
  INV_X1 U7661 ( .A(keyinput6), .ZN(n6749) );
  AOI22_X1 U7662 ( .A1(n6750), .A2(keyinput60), .B1(DATAWIDTH_REG_24__SCAN_IN), 
        .B2(n6749), .ZN(n6748) );
  OAI221_X1 U7663 ( .B1(n6750), .B2(keyinput60), .C1(n6749), .C2(
        DATAWIDTH_REG_24__SCAN_IN), .A(n6748), .ZN(n6761) );
  AOI22_X1 U7664 ( .A1(n6753), .A2(keyinput13), .B1(keyinput27), .B2(n6752), 
        .ZN(n6751) );
  OAI221_X1 U7665 ( .B1(n6753), .B2(keyinput13), .C1(n6752), .C2(keyinput27), 
        .A(n6751), .ZN(n6760) );
  INV_X1 U7666 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6755) );
  AOI22_X1 U7667 ( .A1(n5244), .A2(keyinput43), .B1(n6755), .B2(keyinput32), 
        .ZN(n6754) );
  OAI221_X1 U7668 ( .B1(n5244), .B2(keyinput43), .C1(n6755), .C2(keyinput32), 
        .A(n6754), .ZN(n6759) );
  AOI22_X1 U7669 ( .A1(n3494), .A2(keyinput46), .B1(n6757), .B2(keyinput16), 
        .ZN(n6756) );
  OAI221_X1 U7670 ( .B1(n3494), .B2(keyinput46), .C1(n6757), .C2(keyinput16), 
        .A(n6756), .ZN(n6758) );
  NOR4_X1 U7671 ( .A1(n6761), .A2(n6760), .A3(n6759), .A4(n6758), .ZN(n6777)
         );
  INV_X1 U7672 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U7673 ( .A1(n6764), .A2(keyinput3), .B1(n6763), .B2(keyinput54), 
        .ZN(n6762) );
  OAI221_X1 U7674 ( .B1(n6764), .B2(keyinput3), .C1(n6763), .C2(keyinput54), 
        .A(n6762), .ZN(n6775) );
  AOI22_X1 U7675 ( .A1(n5041), .A2(keyinput17), .B1(keyinput49), .B2(n5515), 
        .ZN(n6765) );
  OAI221_X1 U7676 ( .B1(n5041), .B2(keyinput17), .C1(n5515), .C2(keyinput49), 
        .A(n6765), .ZN(n6774) );
  INV_X1 U7677 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6767) );
  AOI22_X1 U7678 ( .A1(n6768), .A2(keyinput55), .B1(keyinput29), .B2(n6767), 
        .ZN(n6766) );
  OAI221_X1 U7679 ( .B1(n6768), .B2(keyinput55), .C1(n6767), .C2(keyinput29), 
        .A(n6766), .ZN(n6773) );
  INV_X1 U7680 ( .A(keyinput7), .ZN(n6771) );
  INV_X1 U7681 ( .A(keyinput40), .ZN(n6770) );
  AOI22_X1 U7682 ( .A1(n6771), .A2(ADDRESS_REG_28__SCAN_IN), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6770), .ZN(n6769) );
  OAI221_X1 U7683 ( .B1(n6771), .B2(ADDRESS_REG_28__SCAN_IN), .C1(n6770), .C2(
        ADDRESS_REG_10__SCAN_IN), .A(n6769), .ZN(n6772) );
  NOR4_X1 U7684 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n6772), .ZN(n6776)
         );
  NAND4_X1 U7685 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n6780)
         );
  AOI211_X1 U7686 ( .C1(LWORD_REG_10__SCAN_IN), .C2(n6782), .A(n6781), .B(
        n6780), .ZN(n6796) );
  AOI22_X1 U7687 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6785), .B1(n6784), 
        .B2(n6783), .ZN(n6792) );
  OAI22_X1 U7688 ( .A1(n6789), .A2(n6788), .B1(n6787), .B2(n6786), .ZN(n6790)
         );
  INV_X1 U7689 ( .A(n6790), .ZN(n6791) );
  OAI211_X1 U7690 ( .C1(n6794), .C2(n6793), .A(n6792), .B(n6791), .ZN(n6795)
         );
  XOR2_X1 U7691 ( .A(n6796), .B(n6795), .Z(U3126) );
  AND2_X1 U4093 ( .A1(n3209), .A2(n4304), .ZN(n3208) );
  CLKBUF_X1 U3423 ( .A(n3158), .Z(n2980) );
  CLKBUF_X2 U3425 ( .A(n3296), .Z(n3308) );
  CLKBUF_X1 U3433 ( .A(n3274), .Z(n2981) );
  CLKBUF_X3 U3437 ( .A(n3194), .Z(n2988) );
  CLKBUF_X1 U3438 ( .A(n3204), .Z(n2977) );
  NAND2_X1 U3443 ( .A1(n4319), .A2(n4645), .ZN(n3239) );
  CLKBUF_X1 U34550 ( .A(n5802), .Z(n6145) );
  CLKBUF_X1 U3510 ( .A(n3590), .Z(n4817) );
endmodule

