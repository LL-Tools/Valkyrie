

module b20_C_SARLock_k_128_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345;

  INV_X4 U4935 ( .A(n10058), .ZN(n10100) );
  OR2_X1 U4936 ( .A1(n9697), .A2(n7451), .ZN(n7642) );
  NAND2_X1 U4937 ( .A1(n5574), .A2(n5573), .ZN(n8861) );
  NAND2_X1 U4938 ( .A1(n4870), .A2(n5607), .ZN(n5743) );
  XNOR2_X1 U4939 ( .A(n5478), .B(n5477), .ZN(n7337) );
  INV_X1 U4940 ( .A(n4428), .ZN(n4437) );
  AOI21_X1 U4941 ( .B1(n7510), .B2(n7511), .A(n7507), .ZN(n7462) );
  CLKBUF_X2 U4943 ( .A(n6268), .Z(n9127) );
  INV_X1 U4944 ( .A(n9075), .ZN(n9125) );
  CLKBUF_X2 U4945 ( .A(n5264), .Z(n7912) );
  CLKBUF_X2 U4946 ( .A(n7443), .Z(n4431) );
  AND4_X1 U4947 ( .A1(n4799), .A2(n4798), .A3(n4797), .A4(n4796), .ZN(n5880)
         );
  CLKBUF_X1 U4948 ( .A(n6143), .Z(n4433) );
  NAND3_X2 U4949 ( .A1(n6002), .A2(n5999), .A3(n5998), .ZN(n6171) );
  OR2_X1 U4950 ( .A1(n5978), .A2(n6492), .ZN(n5980) );
  NAND2_X1 U4952 ( .A1(n6033), .A2(n9759), .ZN(n9763) );
  OR2_X1 U4953 ( .A1(n5192), .A2(n5405), .ZN(n5163) );
  INV_X2 U4954 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6492) );
  NAND2_X2 U4955 ( .A1(n7278), .A2(n7277), .ZN(n9976) );
  OR2_X1 U4956 ( .A1(n8265), .A2(n8264), .ZN(n8288) );
  INV_X1 U4957 ( .A(n8103), .ZN(n8096) );
  OAI21_X1 U4958 ( .B1(n6135), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6017) );
  BUF_X1 U4959 ( .A(n9122), .Z(n4435) );
  INV_X1 U4960 ( .A(n7319), .ZN(n7450) );
  BUF_X1 U4961 ( .A(n7443), .Z(n4432) );
  NAND2_X1 U4962 ( .A1(n9697), .A2(n7451), .ZN(n9468) );
  NAND2_X1 U4963 ( .A1(n4538), .A2(n7258), .ZN(n7589) );
  NAND2_X1 U4964 ( .A1(n4987), .A2(n4985), .ZN(n6035) );
  NAND2_X1 U4965 ( .A1(n5568), .A2(n5567), .ZN(n5586) );
  NAND2_X1 U4966 ( .A1(n4878), .A2(n5141), .ZN(n5515) );
  NAND2_X1 U4967 ( .A1(n5609), .A2(n5608), .ZN(n7785) );
  AND4_X1 U4968 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n6591)
         );
  NOR2_X1 U4969 ( .A1(n5924), .A2(n5925), .ZN(n5923) );
  OAI21_X1 U4970 ( .B1(n5806), .B2(n6807), .A(n6803), .ZN(n6930) );
  NAND2_X2 U4971 ( .A1(n5408), .A2(n5407), .ZN(n7679) );
  NAND2_X1 U4972 ( .A1(n5199), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5195) );
  BUF_X1 U4973 ( .A(n10078), .Z(n4440) );
  CLKBUF_X3 U4974 ( .A(n10026), .Z(n4434) );
  NAND4_X1 U4975 ( .A1(n5399), .A2(n5398), .A3(n5397), .A4(n5396), .ZN(n8125)
         );
  AOI21_X1 U4976 ( .B1(n4449), .B2(n8148), .A(n4654), .ZN(n4653) );
  AND2_X1 U4977 ( .A1(n7290), .A2(n7289), .ZN(n4428) );
  AND2_X1 U4978 ( .A1(n5764), .A2(n5053), .ZN(n4429) );
  XNOR2_X1 U4979 ( .A(n6142), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10026) );
  AND2_X2 U4980 ( .A1(n5404), .A2(n5403), .ZN(n6992) );
  NOR2_X2 U4981 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n6575) );
  INV_X2 U4982 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5833) );
  OAI21_X2 U4983 ( .B1(n6963), .B2(n4783), .A(n4780), .ZN(n7049) );
  NAND2_X2 U4984 ( .A1(n5340), .A2(n5339), .ZN(n6963) );
  NAND2_X2 U4985 ( .A1(n7187), .A2(n4512), .ZN(n7209) );
  XNOR2_X2 U4986 ( .A(n7910), .B(n7946), .ZN(n5762) );
  NAND2_X2 U4987 ( .A1(n5753), .A2(n5752), .ZN(n7910) );
  AND2_X1 U4988 ( .A1(n4710), .A2(n4711), .ZN(n4430) );
  AND2_X2 U4989 ( .A1(n4710), .A2(n4711), .ZN(n7904) );
  AND2_X2 U4990 ( .A1(n5978), .A2(n5979), .ZN(n5964) );
  AND2_X2 U4992 ( .A1(n5043), .A2(n4795), .ZN(n6586) );
  OR2_X1 U4993 ( .A1(n5247), .A2(n5835), .ZN(n5043) );
  INV_X1 U4994 ( .A(n7360), .ZN(n7443) );
  XNOR2_X2 U4995 ( .A(n5061), .B(n4875), .ZN(n5060) );
  XNOR2_X1 U4996 ( .A(n6017), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6143) );
  INV_X2 U4997 ( .A(n5634), .ZN(n8116) );
  OAI21_X2 U4998 ( .B1(n5351), .B2(n5350), .A(n5087), .ZN(n5364) );
  NAND2_X2 U4999 ( .A1(n5081), .A2(n5080), .ZN(n5351) );
  AOI211_X2 U5000 ( .C1(n10097), .C2(n9691), .A(n9500), .B(n9499), .ZN(n9501)
         );
  NAND2_X2 U5001 ( .A1(n4573), .A2(n4935), .ZN(n6835) );
  OAI21_X2 U5002 ( .B1(n8318), .B2(n5604), .A(n5603), .ZN(n5741) );
  NAND2_X2 U5003 ( .A1(n5584), .A2(n5583), .ZN(n8318) );
  OAI21_X2 U5004 ( .B1(n9835), .B2(n9841), .A(n7625), .ZN(n9645) );
  NAND2_X2 U5005 ( .A1(n9665), .A2(n7531), .ZN(n9835) );
  AOI21_X2 U5006 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n9331), .A(n9324), .ZN(
        n9340) );
  INV_X2 U5007 ( .A(n5663), .ZN(n4575) );
  NAND2_X1 U5008 ( .A1(n7735), .A2(n8479), .ZN(n7736) );
  OAI21_X2 U5009 ( .B1(n5515), .B2(n5514), .A(n5146), .ZN(n5527) );
  XNOR2_X2 U5010 ( .A(n5743), .B(n5742), .ZN(n9770) );
  NAND2_X2 U5012 ( .A1(n7642), .A2(n9468), .ZN(n9508) );
  OAI22_X2 U5013 ( .A1(n7156), .A2(n7155), .B1(n7154), .B2(n7163), .ZN(n7158)
         );
  NAND2_X2 U5014 ( .A1(n4532), .A2(n5485), .ZN(n8819) );
  AOI22_X2 U5015 ( .A1(n7787), .A2(n7788), .B1(n8393), .B2(n7702), .ZN(n7862)
         );
  NAND2_X2 U5016 ( .A1(n4626), .A2(n4949), .ZN(n7787) );
  INV_X1 U5017 ( .A(n8125), .ZN(n7801) );
  NAND2_X2 U5018 ( .A1(n5496), .A2(n5495), .ZN(n8896) );
  XNOR2_X2 U5019 ( .A(n6035), .B(n6034), .ZN(n6039) );
  AOI21_X1 U5020 ( .B1(n6268), .B2(n10089), .A(n4934), .ZN(n6273) );
  XNOR2_X2 U5021 ( .A(n7185), .B(n7183), .ZN(n7087) );
  NAND2_X2 U5022 ( .A1(n4599), .A2(n4958), .ZN(n7185) );
  XNOR2_X2 U5023 ( .A(n5586), .B(n5585), .ZN(n8952) );
  AOI22_X2 U5024 ( .A1(n6930), .A2(n6931), .B1(n4659), .B2(n5808), .ZN(n6971)
         );
  OAI21_X2 U5025 ( .B1(n6035), .B2(n6029), .A(n6028), .ZN(n6033) );
  AOI22_X2 U5026 ( .A1(n6695), .A2(n7490), .B1(n6694), .B2(n6693), .ZN(n10049)
         );
  OAI22_X2 U5027 ( .A1(n10062), .A2(n10061), .B1(n10060), .B2(n9281), .ZN(
        n6695) );
  AOI21_X2 U5028 ( .B1(n8452), .B2(n8830), .A(n8439), .ZN(n8421) );
  OAI21_X2 U5029 ( .B1(n9509), .B2(n9508), .A(n9468), .ZN(n9492) );
  NOR2_X2 U5030 ( .A1(n9524), .A2(n9467), .ZN(n9509) );
  INV_X1 U5031 ( .A(n4428), .ZN(n4436) );
  INV_X1 U5032 ( .A(n4428), .ZN(n4438) );
  CLKBUF_X1 U5033 ( .A(n10078), .Z(n4439) );
  OAI211_X1 U5034 ( .C1(n6786), .C2(n6267), .A(n6266), .B(n6265), .ZN(n10078)
         );
  INV_X2 U5035 ( .A(n7678), .ZN(n5242) );
  AOI21_X2 U5036 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9345), .A(n9338), .ZN(
        n9799) );
  AOI211_X2 U5037 ( .C1(P1_ADDR_REG_19__SCAN_IN), .C2(n9883), .A(n9400), .B(
        n9399), .ZN(n9401) );
  NAND2_X1 U5038 ( .A1(n9194), .A2(n9056), .ZN(n9160) );
  INV_X1 U5039 ( .A(n7589), .ZN(n9684) );
  OAI21_X1 U5040 ( .B1(n9103), .B2(n9105), .A(n9104), .ZN(n9102) );
  NAND2_X2 U5041 ( .A1(n8007), .A2(n7991), .ZN(n7211) );
  CLKBUF_X1 U5042 ( .A(n8779), .Z(n4556) );
  AND4_X2 U5043 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n8134)
         );
  INV_X1 U5044 ( .A(n6656), .ZN(n10124) );
  CLKBUF_X2 U5045 ( .A(n5243), .Z(n5746) );
  CLKBUF_X1 U5046 ( .A(n5247), .Z(n7905) );
  NAND2_X2 U5047 ( .A1(n5242), .A2(n8942), .ZN(n5249) );
  NOR2_X1 U5048 ( .A1(n6507), .A2(n4433), .ZN(n7600) );
  CLKBUF_X2 U5050 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9779) );
  AOI21_X1 U5051 ( .B1(n4429), .B2(n4760), .A(n4529), .ZN(n4759) );
  OAI21_X1 U5052 ( .B1(n9131), .B2(n9086), .A(n9247), .ZN(n9090) );
  NAND2_X1 U5053 ( .A1(n9159), .A2(n9069), .ZN(n9246) );
  NAND2_X1 U5054 ( .A1(n4621), .A2(n7722), .ZN(n7725) );
  NAND2_X1 U5055 ( .A1(n8849), .A2(n8312), .ZN(n8101) );
  AOI21_X1 U5056 ( .B1(n9496), .B2(n10112), .A(n9495), .ZN(n9694) );
  NAND2_X1 U5057 ( .A1(n9160), .A2(n9161), .ZN(n9159) );
  NAND2_X1 U5058 ( .A1(n7906), .A2(n7905), .ZN(n8849) );
  NOR4_X1 U5059 ( .A1(n9470), .A2(n9484), .A3(n9508), .A4(n7481), .ZN(n7483)
         );
  NAND2_X1 U5060 ( .A1(n7255), .A2(n7254), .ZN(n7593) );
  NAND2_X1 U5061 ( .A1(n9689), .A2(n7453), .ZN(n7583) );
  NAND2_X1 U5062 ( .A1(n7903), .A2(n7902), .ZN(n8790) );
  NAND2_X1 U5063 ( .A1(n7714), .A2(n7713), .ZN(n7807) );
  NAND2_X1 U5064 ( .A1(n5748), .A2(n5747), .ZN(n7951) );
  OR2_X1 U5065 ( .A1(n8855), .A2(n7881), .ZN(n8088) );
  XNOR2_X1 U5066 ( .A(n7257), .B(n7256), .ZN(n7901) );
  OAI21_X1 U5067 ( .B1(n7246), .B2(n7245), .A(n7244), .ZN(n7257) );
  XNOR2_X1 U5068 ( .A(n7246), .B(SI_29_), .ZN(n7259) );
  XNOR2_X1 U5069 ( .A(n4656), .B(n8286), .ZN(n4655) );
  NAND2_X1 U5070 ( .A1(n7427), .A2(n7426), .ZN(n9697) );
  XNOR2_X1 U5071 ( .A(n7243), .B(n7242), .ZN(n7246) );
  NAND2_X1 U5072 ( .A1(n5525), .A2(n4793), .ZN(n8346) );
  AND2_X1 U5073 ( .A1(n7923), .A2(n7922), .ZN(n8337) );
  OR2_X1 U5074 ( .A1(n9703), .A2(n9454), .ZN(n7458) );
  NOR2_X1 U5075 ( .A1(n8248), .A2(n8249), .ZN(n8274) );
  XNOR2_X1 U5076 ( .A(n5606), .B(n5605), .ZN(n8947) );
  NAND2_X1 U5077 ( .A1(n7860), .A2(n7704), .ZN(n7709) );
  NAND2_X1 U5078 ( .A1(n9201), .A2(n9025), .ZN(n9141) );
  NAND2_X1 U5079 ( .A1(n5588), .A2(n5587), .ZN(n5606) );
  AOI21_X1 U5080 ( .B1(n8308), .B2(n8309), .A(n8307), .ZN(n4858) );
  OAI211_X1 U5081 ( .C1(n8367), .C2(n4814), .A(n4508), .B(n4547), .ZN(n5702)
         );
  NOR2_X1 U5082 ( .A1(n9544), .A2(n4845), .ZN(n4844) );
  OR2_X1 U5083 ( .A1(n9713), .A2(n9447), .ZN(n9465) );
  NAND2_X1 U5084 ( .A1(n7345), .A2(n7344), .ZN(n9713) );
  NAND2_X1 U5085 ( .A1(n5534), .A2(n5533), .ZN(n7839) );
  AOI22_X1 U5086 ( .A1(n9602), .A2(n9436), .B1(n9435), .B2(n9733), .ZN(n9588)
         );
  NAND2_X1 U5087 ( .A1(n5548), .A2(n5547), .ZN(n5566) );
  AOI21_X1 U5088 ( .B1(n4773), .B2(n4769), .A(n4768), .ZN(n4767) );
  AND2_X1 U5089 ( .A1(n5171), .A2(n5170), .ZN(n7706) );
  NAND2_X1 U5090 ( .A1(n5517), .A2(n5516), .ZN(n8884) );
  NAND2_X1 U5091 ( .A1(n4774), .A2(n8391), .ZN(n4773) );
  XNOR2_X1 U5092 ( .A(n5527), .B(n5526), .ZN(n7354) );
  OR2_X2 U5093 ( .A1(n9819), .A2(n9818), .ZN(n9821) );
  NAND2_X1 U5094 ( .A1(n7404), .A2(n7403), .ZN(n9728) );
  CLKBUF_X1 U5095 ( .A(n7734), .Z(n4574) );
  NAND2_X1 U5096 ( .A1(n5507), .A2(n5506), .ZN(n8890) );
  OR2_X1 U5097 ( .A1(n8896), .A2(n7791), .ZN(n8055) );
  NAND2_X1 U5098 ( .A1(n4906), .A2(n4905), .ZN(n9228) );
  AOI21_X1 U5099 ( .B1(n4566), .B2(n4456), .A(n4494), .ZN(n9650) );
  NAND2_X1 U5100 ( .A1(n7341), .A2(n7340), .ZN(n9737) );
  OR2_X1 U5101 ( .A1(n8999), .A2(n8998), .ZN(n4904) );
  XNOR2_X1 U5102 ( .A(n5493), .B(n5492), .ZN(n7415) );
  NAND2_X1 U5103 ( .A1(n7327), .A2(n7326), .ZN(n9641) );
  NAND2_X1 U5104 ( .A1(n4886), .A2(n5132), .ZN(n5493) );
  NAND2_X1 U5105 ( .A1(n5469), .A2(n5468), .ZN(n8903) );
  XNOR2_X1 U5106 ( .A(n8993), .B(n9125), .ZN(n9169) );
  OR2_X1 U5107 ( .A1(n5466), .A2(n4572), .ZN(n4885) );
  NAND2_X1 U5108 ( .A1(n7316), .A2(n7315), .ZN(n9825) );
  CLKBUF_X1 U5109 ( .A(n9656), .Z(n4578) );
  XNOR2_X1 U5110 ( .A(n5466), .B(n5465), .ZN(n7325) );
  NAND2_X1 U5111 ( .A1(n7305), .A2(n7304), .ZN(n9656) );
  NAND2_X1 U5112 ( .A1(n5232), .A2(n5231), .ZN(n8830) );
  NAND2_X1 U5113 ( .A1(n5455), .A2(n5454), .ZN(n8916) );
  AND2_X1 U5114 ( .A1(n6593), .A2(n6592), .ZN(n6598) );
  NAND2_X1 U5115 ( .A1(n6627), .A2(n6626), .ZN(n6736) );
  XNOR2_X1 U5116 ( .A(n5227), .B(n5226), .ZN(n7303) );
  NAND2_X1 U5117 ( .A1(n4856), .A2(n7062), .ZN(n5853) );
  NAND2_X1 U5118 ( .A1(n4887), .A2(n5117), .ZN(n5227) );
  NAND2_X1 U5119 ( .A1(n5442), .A2(n5441), .ZN(n8923) );
  NAND2_X1 U5120 ( .A1(n5451), .A2(n5116), .ZN(n4887) );
  NAND2_X1 U5121 ( .A1(n4914), .A2(n4911), .ZN(n6631) );
  NAND2_X1 U5122 ( .A1(n5848), .A2(n6983), .ZN(n6986) );
  NAND2_X1 U5123 ( .A1(n5393), .A2(n5392), .ZN(n8779) );
  OAI21_X1 U5124 ( .B1(n6715), .B2(n4459), .A(n4496), .ZN(n6892) );
  NAND2_X1 U5125 ( .A1(n4699), .A2(n4700), .ZN(n5402) );
  NAND2_X1 U5126 ( .A1(n6429), .A2(n6428), .ZN(n6459) );
  OAI21_X1 U5127 ( .B1(n5372), .B2(n5094), .A(n5097), .ZN(n5389) );
  NAND2_X1 U5128 ( .A1(n6851), .A2(n6850), .ZN(n10024) );
  AND2_X1 U5129 ( .A1(n6910), .A2(n7506), .ZN(n10032) );
  OAI211_X1 U5130 ( .C1(n7905), .C2(n6979), .A(n5354), .B(n5353), .ZN(n7086)
         );
  BUF_X4 U5131 ( .A(n5886), .Z(n7778) );
  INV_X2 U5132 ( .A(n6046), .ZN(n6197) );
  AND3_X1 U5133 ( .A1(n5306), .A2(n5305), .A3(n5304), .ZN(n10256) );
  NAND2_X1 U5134 ( .A1(n4862), .A2(n4863), .ZN(n5336) );
  CLKBUF_X1 U5135 ( .A(n5656), .Z(n5989) );
  NOR2_X1 U5136 ( .A1(n6285), .A2(n10082), .ZN(n7464) );
  OAI211_X2 U5137 ( .C1(n7319), .C2(n6289), .A(n6184), .B(n6183), .ZN(n9283)
         );
  NAND2_X1 U5138 ( .A1(n5072), .A2(n5071), .ZN(n5299) );
  INV_X1 U5139 ( .A(n5746), .ZN(n5484) );
  AND3_X1 U5140 ( .A1(n5261), .A2(n5260), .A3(n5259), .ZN(n6537) );
  INV_X2 U5141 ( .A(n5246), .ZN(n7900) );
  AND3_X1 U5142 ( .A1(n5233), .A2(n5236), .A3(n4959), .ZN(n6581) );
  NAND2_X1 U5143 ( .A1(n4435), .A2(n9075), .ZN(n6268) );
  AOI21_X1 U5144 ( .B1(n6239), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6229), .ZN(
        n9326) );
  AND2_X1 U5145 ( .A1(n5651), .A2(n5650), .ZN(n5663) );
  CLKBUF_X1 U5146 ( .A(n5652), .Z(n5653) );
  NAND2_X1 U5147 ( .A1(n4546), .A2(n5068), .ZN(n5287) );
  INV_X4 U5148 ( .A(n5045), .ZN(n9121) );
  INV_X2 U5149 ( .A(n6847), .ZN(n7425) );
  XNOR2_X1 U5150 ( .A(n5366), .B(n5365), .ZN(n6979) );
  INV_X1 U5151 ( .A(n5456), .ZN(n5756) );
  OR2_X1 U5152 ( .A1(n9763), .A2(n6037), .ZN(n6180) );
  CLKBUF_X1 U5153 ( .A(n6185), .Z(n9774) );
  NAND2_X2 U5154 ( .A1(n6185), .A2(n6225), .ZN(n6786) );
  CLKBUF_X2 U5155 ( .A(n6039), .Z(n6037) );
  AOI21_X1 U5156 ( .B1(n4865), .B2(n4867), .A(n4498), .ZN(n4863) );
  NAND2_X1 U5157 ( .A1(n5200), .A2(n5199), .ZN(n8942) );
  XNOR2_X1 U5158 ( .A(n6025), .B(n6013), .ZN(n6185) );
  NAND2_X1 U5159 ( .A1(n5198), .A2(n5197), .ZN(n5200) );
  OAI21_X1 U5160 ( .B1(n5298), .B2(n4867), .A(n5321), .ZN(n4866) );
  NAND2_X1 U5161 ( .A1(n6030), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U5162 ( .A1(n5196), .A2(n5193), .ZN(n5199) );
  XNOR2_X1 U5163 ( .A(n6018), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7599) );
  AND2_X1 U5164 ( .A1(n6012), .A2(n6011), .ZN(n6014) );
  OR2_X1 U5165 ( .A1(n6133), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6135) );
  AND2_X1 U5166 ( .A1(n4982), .A2(n5160), .ZN(n4830) );
  CLKBUF_X1 U5167 ( .A(n6345), .Z(n6346) );
  CLKBUF_X1 U5168 ( .A(n5967), .Z(n5983) );
  INV_X2 U5169 ( .A(n7904), .ZN(n5549) );
  AND2_X1 U5170 ( .A1(n5780), .A2(n5967), .ZN(n6345) );
  NOR2_X1 U5171 ( .A1(n4983), .A2(n4485), .ZN(n4982) );
  AND2_X1 U5172 ( .A1(n5964), .A2(n5779), .ZN(n5967) );
  OR2_X1 U5173 ( .A1(n4664), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U5174 ( .A1(n6574), .A2(n5057), .ZN(n4710) );
  AND4_X1 U5175 ( .A1(n5153), .A2(n5152), .A3(n5151), .A4(n5316), .ZN(n5154)
         );
  INV_X1 U5176 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5316) );
  AND2_X1 U5177 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n6574) );
  INV_X4 U5178 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5179 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5438) );
  NOR2_X1 U5180 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5781) );
  INV_X1 U5181 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6013) );
  NOR2_X1 U5182 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5793) );
  INV_X1 U5183 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8636) );
  NOR2_X1 U5184 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5775) );
  NOR2_X1 U5185 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5152) );
  INV_X1 U5186 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5773) );
  NOR2_X1 U5187 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5151) );
  INV_X4 U5188 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U5189 ( .A1(n5372), .A2(n4703), .ZN(n4699) );
  NOR2_X2 U5190 ( .A1(n9525), .A2(n9526), .ZN(n9524) );
  XNOR2_X1 U5191 ( .A(n5364), .B(n5363), .ZN(n6848) );
  NAND2_X2 U5192 ( .A1(n7087), .A2(n7088), .ZN(n7187) );
  MUX2_X2 U5193 ( .A(n9398), .B(n9397), .S(n6507), .Z(n9399) );
  INV_X1 U5194 ( .A(n4965), .ZN(n4963) );
  INV_X1 U5195 ( .A(n5249), .ZN(n4442) );
  CLKBUF_X1 U5196 ( .A(n5880), .Z(n6532) );
  INV_X1 U5197 ( .A(n5880), .ZN(n5248) );
  NAND2_X1 U5198 ( .A1(n6586), .A2(n5880), .ZN(n5687) );
  XNOR2_X2 U5199 ( .A(n7709), .B(n7707), .ZN(n7747) );
  OAI21_X2 U5200 ( .B1(n6553), .B2(n5291), .A(n5290), .ZN(n6715) );
  AOI21_X2 U5201 ( .B1(n7807), .B2(n7808), .A(n7717), .ZN(n7719) );
  OAI21_X2 U5202 ( .B1(n8485), .B2(n4820), .A(n4818), .ZN(n8448) );
  NAND2_X2 U5203 ( .A1(n5634), .A2(n5633), .ZN(n5247) );
  XNOR2_X2 U5204 ( .A(n5163), .B(n5191), .ZN(n5633) );
  INV_X2 U5205 ( .A(n4435), .ZN(n6421) );
  INV_X1 U5206 ( .A(n4664), .ZN(n5256) );
  NAND2_X1 U5207 ( .A1(n7699), .A2(n8394), .ZN(n4957) );
  NAND2_X1 U5208 ( .A1(n5931), .A2(n5820), .ZN(n5821) );
  AND2_X1 U5209 ( .A1(n4978), .A2(n4977), .ZN(n4976) );
  INV_X1 U5210 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4977) );
  INV_X1 U5211 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5213) );
  NAND3_X1 U5212 ( .A1(n6166), .A2(n4923), .A3(n7604), .ZN(n4921) );
  NAND2_X1 U5213 ( .A1(n4922), .A2(n4434), .ZN(n4923) );
  INV_X1 U5214 ( .A(n10032), .ZN(n5003) );
  NAND2_X1 U5215 ( .A1(n4430), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4876) );
  AND2_X1 U5216 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  AND2_X2 U5217 ( .A1(n7689), .A2(n7739), .ZN(n4973) );
  AOI21_X1 U5218 ( .B1(n7737), .B2(n7687), .A(n7686), .ZN(n7689) );
  AOI21_X1 U5219 ( .B1(n4900), .B2(n4897), .A(n4896), .ZN(n4895) );
  INV_X1 U5220 ( .A(n9237), .ZN(n4896) );
  NOR2_X1 U5221 ( .A1(n4901), .A2(n9236), .ZN(n4897) );
  NAND2_X1 U5222 ( .A1(n4726), .A2(n4482), .ZN(n7533) );
  OR2_X1 U5223 ( .A1(n7622), .A2(n4734), .ZN(n4724) );
  INV_X1 U5224 ( .A(n4872), .ZN(n4871) );
  OAI21_X1 U5225 ( .B1(n5605), .B2(n4873), .A(n5742), .ZN(n4872) );
  AOI21_X1 U5226 ( .B1(n4694), .B2(n4693), .A(n8082), .ZN(n4692) );
  INV_X1 U5227 ( .A(n4701), .ZN(n4700) );
  OAI21_X1 U5228 ( .B1(n5373), .B2(n4702), .A(n4488), .ZN(n4701) );
  AOI21_X1 U5229 ( .B1(n4444), .B2(n6836), .A(n4489), .ZN(n4958) );
  NAND2_X1 U5230 ( .A1(n6835), .A2(n4444), .ZN(n4599) );
  NOR2_X1 U5231 ( .A1(n8098), .A2(n8097), .ZN(n8109) );
  AND2_X1 U5232 ( .A1(n8104), .A2(n8096), .ZN(n8108) );
  AND2_X1 U5233 ( .A1(n5200), .A2(n5199), .ZN(n5241) );
  NAND2_X1 U5234 ( .A1(n4670), .A2(n4669), .ZN(n7232) );
  NAND2_X1 U5235 ( .A1(n7060), .A2(n4461), .ZN(n4669) );
  NAND2_X1 U5236 ( .A1(n4672), .A2(n4671), .ZN(n4670) );
  OR2_X1 U5237 ( .A1(n7951), .A2(n7953), .ZN(n8102) );
  OR2_X1 U5238 ( .A1(n8819), .A2(n8394), .ZN(n8047) );
  AND2_X1 U5239 ( .A1(n4632), .A2(n5156), .ZN(n4631) );
  AND2_X1 U5240 ( .A1(n4615), .A2(n4608), .ZN(n4607) );
  NAND2_X1 U5241 ( .A1(n4610), .A2(n4609), .ZN(n4608) );
  AOI21_X1 U5242 ( .B1(n9149), .B2(n4617), .A(n4499), .ZN(n4615) );
  INV_X1 U5243 ( .A(n9111), .ZN(n4892) );
  AND2_X1 U5244 ( .A1(n4739), .A2(n7596), .ZN(n4545) );
  AND2_X1 U5245 ( .A1(n6089), .A2(n6088), .ZN(n7293) );
  NAND2_X1 U5246 ( .A1(n10183), .A2(n9414), .ZN(n5031) );
  NAND2_X1 U5247 ( .A1(n5031), .A2(n5032), .ZN(n5020) );
  OR2_X1 U5248 ( .A1(n9156), .A2(n9414), .ZN(n7519) );
  AND2_X1 U5249 ( .A1(n9279), .A2(n10141), .ZN(n7615) );
  OR2_X1 U5250 ( .A1(n7243), .A2(n7242), .ZN(n7244) );
  NAND2_X1 U5251 ( .A1(n7209), .A2(n7208), .ZN(n4606) );
  INV_X1 U5252 ( .A(n7843), .ZN(n4950) );
  NAND2_X1 U5253 ( .A1(n4601), .A2(n4604), .ZN(n7734) );
  NAND2_X1 U5254 ( .A1(n7760), .A2(n7210), .ZN(n4604) );
  NOR2_X1 U5255 ( .A1(n4605), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U5256 ( .A1(n7696), .A2(n8440), .ZN(n4627) );
  INV_X1 U5257 ( .A(n7889), .ZN(n4969) );
  INV_X1 U5258 ( .A(n5192), .ZN(n5169) );
  AOI21_X1 U5259 ( .B1(n5167), .B2(n5166), .A(n5165), .ZN(n5168) );
  AND2_X1 U5260 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5166) );
  INV_X1 U5261 ( .A(n7912), .ZN(n5630) );
  NAND2_X1 U5262 ( .A1(n5822), .A2(n6814), .ZN(n6819) );
  OR2_X1 U5263 ( .A1(n8194), .A2(n8834), .ZN(n4637) );
  OR2_X1 U5264 ( .A1(n8830), .A2(n8423), .ZN(n8044) );
  AOI21_X1 U5265 ( .B1(n4782), .B2(n4781), .A(n4486), .ZN(n4780) );
  INV_X1 U5266 ( .A(n5356), .ZN(n4781) );
  INV_X1 U5267 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5056) );
  XNOR2_X1 U5268 ( .A(n7785), .B(n8320), .ZN(n7919) );
  OR2_X1 U5269 ( .A1(n8929), .A2(n8465), .ZN(n5430) );
  INV_X1 U5270 ( .A(n8477), .ZN(n8461) );
  AND2_X1 U5271 ( .A1(n4830), .A2(n5191), .ZN(n4829) );
  OAI21_X1 U5272 ( .B1(n5467), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5480) );
  INV_X1 U5273 ( .A(n9271), .ZN(n9454) );
  AND3_X1 U5274 ( .A1(n9170), .A2(n9169), .A3(n8994), .ZN(n8998) );
  NAND2_X1 U5275 ( .A1(n4570), .A2(n7597), .ZN(n4569) );
  OAI21_X1 U5276 ( .B1(n4540), .B2(n6190), .A(n4539), .ZN(n7658) );
  NAND2_X1 U5277 ( .A1(n4540), .A2(n7657), .ZN(n4539) );
  OAI21_X1 U5278 ( .B1(n7655), .B2(n7656), .A(n7654), .ZN(n4540) );
  AOI21_X1 U5279 ( .B1(n9515), .B2(n5036), .A(n5034), .ZN(n9459) );
  AND2_X1 U5280 ( .A1(n9458), .A2(n5038), .ZN(n5036) );
  OAI21_X1 U5281 ( .B1(n5037), .B2(n5035), .A(n4490), .ZN(n5034) );
  OR2_X1 U5282 ( .A1(n10002), .A2(n7009), .ZN(n7518) );
  OR2_X1 U5283 ( .A1(n10002), .A2(n8963), .ZN(n5032) );
  AOI21_X1 U5284 ( .B1(n5002), .B2(n4993), .A(n4992), .ZN(n4991) );
  NOR2_X1 U5285 ( .A1(n4995), .A2(n6913), .ZN(n4992) );
  AND2_X1 U5286 ( .A1(n4999), .A2(n5005), .ZN(n4993) );
  NOR2_X1 U5287 ( .A1(n4998), .A2(n4995), .ZN(n4994) );
  INV_X1 U5288 ( .A(n7439), .ZN(n7339) );
  INV_X1 U5289 ( .A(n6786), .ZN(n7338) );
  NAND2_X1 U5290 ( .A1(n4733), .A2(n4729), .ZN(n7500) );
  NAND2_X1 U5291 ( .A1(n4730), .A2(n7600), .ZN(n4729) );
  AOI21_X1 U5292 ( .B1(n8029), .B2(n8030), .A(n4721), .ZN(n4720) );
  INV_X1 U5293 ( .A(n8028), .ZN(n4721) );
  INV_X1 U5294 ( .A(n8484), .ZN(n4719) );
  MUX2_X1 U5295 ( .A(n7514), .B(n7513), .S(n4734), .Z(n7522) );
  NAND2_X1 U5296 ( .A1(n4560), .A2(n8039), .ZN(n8040) );
  AND2_X1 U5297 ( .A1(n8449), .A2(n8037), .ZN(n4561) );
  OAI21_X1 U5298 ( .B1(n4688), .B2(n8043), .A(n4687), .ZN(n4686) );
  AND2_X1 U5299 ( .A1(n8048), .A2(n8042), .ZN(n4687) );
  NAND2_X1 U5300 ( .A1(n4685), .A2(n4683), .ZN(n8050) );
  OR2_X1 U5301 ( .A1(n4688), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U5302 ( .A1(n4686), .A2(n8096), .ZN(n4685) );
  NAND2_X1 U5303 ( .A1(n8044), .A2(n8103), .ZN(n4684) );
  NAND2_X1 U5304 ( .A1(n4553), .A2(n4549), .ZN(n7556) );
  OR2_X1 U5305 ( .A1(n7548), .A2(n4554), .ZN(n4553) );
  NAND2_X1 U5306 ( .A1(n4552), .A2(n4550), .ZN(n4549) );
  NAND2_X1 U5307 ( .A1(n9431), .A2(n4734), .ZN(n4554) );
  AND2_X1 U5308 ( .A1(n7530), .A2(n7531), .ZN(n4723) );
  OAI21_X1 U5309 ( .B1(n4713), .B2(n4712), .A(n8069), .ZN(n8076) );
  NAND2_X1 U5310 ( .A1(n8366), .A2(n8062), .ZN(n4712) );
  AOI21_X1 U5311 ( .B1(n4716), .B2(n4715), .A(n4714), .ZN(n4713) );
  INV_X1 U5312 ( .A(n5607), .ZN(n4873) );
  INV_X1 U5313 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5041) );
  INV_X1 U5314 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5160) );
  AND2_X1 U5315 ( .A1(n4619), .A2(n4618), .ZN(n4617) );
  INV_X1 U5316 ( .A(n6783), .ZN(n4920) );
  AOI22_X1 U5317 ( .A1(n7583), .A2(n7587), .B1(n7582), .B2(n4734), .ZN(n7585)
         );
  NOR2_X1 U5318 ( .A1(n9156), .A2(n9984), .ZN(n4589) );
  NAND2_X1 U5319 ( .A1(n5401), .A2(n5103), .ZN(n4882) );
  INV_X1 U5320 ( .A(SI_14_), .ZN(n8606) );
  INV_X1 U5321 ( .A(n5097), .ZN(n4704) );
  AND2_X1 U5322 ( .A1(n7827), .A2(n7826), .ZN(n4629) );
  AOI21_X1 U5323 ( .B1(n8849), .B2(n8790), .A(n8094), .ZN(n4800) );
  NAND2_X1 U5324 ( .A1(n5664), .A2(n4981), .ZN(n5167) );
  INV_X1 U5325 ( .A(n4983), .ZN(n4981) );
  NAND2_X1 U5326 ( .A1(n6379), .A2(n5838), .ZN(n5839) );
  NAND2_X1 U5327 ( .A1(n4674), .A2(n4522), .ZN(n4672) );
  NAND2_X1 U5328 ( .A1(n8819), .A2(n8415), .ZN(n4779) );
  NAND2_X1 U5329 ( .A1(n5355), .A2(n5356), .ZN(n4784) );
  OR2_X1 U5330 ( .A1(n8861), .A2(n7718), .ZN(n8083) );
  OR2_X1 U5331 ( .A1(n8867), .A2(n8328), .ZN(n7922) );
  OR2_X1 U5332 ( .A1(n7839), .A2(n7750), .ZN(n8074) );
  OR2_X1 U5333 ( .A1(n8884), .A2(n8385), .ZN(n5524) );
  INV_X1 U5334 ( .A(n8382), .ZN(n4771) );
  NOR2_X1 U5335 ( .A1(n4467), .A2(n8382), .ZN(n4769) );
  OR2_X1 U5336 ( .A1(n8890), .A2(n8393), .ZN(n8061) );
  OR2_X1 U5337 ( .A1(n8903), .A2(n8424), .ZN(n8048) );
  AOI21_X1 U5338 ( .B1(n8032), .B2(n7938), .A(n4822), .ZN(n4821) );
  INV_X1 U5339 ( .A(n8037), .ZN(n4822) );
  INV_X1 U5340 ( .A(n7991), .ZN(n4813) );
  INV_X1 U5341 ( .A(n8020), .ZN(n4812) );
  INV_X1 U5342 ( .A(n4807), .ZN(n4806) );
  INV_X1 U5343 ( .A(n8007), .ZN(n4803) );
  NOR2_X1 U5344 ( .A1(n7052), .A2(n4808), .ZN(n4807) );
  INV_X1 U5345 ( .A(n8008), .ZN(n4808) );
  NAND2_X1 U5346 ( .A1(n8291), .A2(n8100), .ZN(n5876) );
  INV_X1 U5347 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5666) );
  INV_X1 U5348 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5161) );
  AND2_X1 U5349 ( .A1(n5215), .A2(n5213), .ZN(n4632) );
  AND2_X1 U5350 ( .A1(n5257), .A2(n4980), .ZN(n4633) );
  AND2_X1 U5351 ( .A1(n6285), .A2(n9121), .ZN(n4934) );
  AOI21_X1 U5352 ( .B1(n4890), .B2(n4898), .A(n4518), .ZN(n4889) );
  NOR2_X1 U5353 ( .A1(n4843), .A2(n9538), .ZN(n4842) );
  INV_X1 U5354 ( .A(n4844), .ZN(n4843) );
  NOR2_X1 U5355 ( .A1(n9728), .A2(n9733), .ZN(n4584) );
  NOR2_X1 U5356 ( .A1(n9723), .A2(n4583), .ZN(n4582) );
  INV_X1 U5357 ( .A(n4584), .ZN(n4583) );
  OR2_X1 U5358 ( .A1(n9728), .A2(n9438), .ZN(n9439) );
  OR2_X1 U5359 ( .A1(n9598), .A2(n9437), .ZN(n5047) );
  OR2_X1 U5360 ( .A1(n9733), .A2(n9434), .ZN(n7545) );
  NAND2_X1 U5361 ( .A1(n9674), .A2(n9418), .ZN(n5030) );
  NOR2_X1 U5362 ( .A1(n4468), .A2(n5020), .ZN(n5019) );
  NAND2_X1 U5363 ( .A1(n7388), .A2(n7387), .ZN(n9707) );
  XNOR2_X1 U5364 ( .A(n5134), .B(SI_20_), .ZN(n5492) );
  INV_X1 U5365 ( .A(n5401), .ZN(n4705) );
  AND2_X1 U5366 ( .A1(n5093), .A2(n5092), .ZN(n5363) );
  INV_X1 U5367 ( .A(n5075), .ZN(n4867) );
  INV_X1 U5368 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5779) );
  INV_X1 U5369 ( .A(n7698), .ZN(n4954) );
  OAI21_X1 U5370 ( .B1(n4947), .B2(n4944), .A(n4943), .ZN(n4942) );
  NOR2_X1 U5371 ( .A1(n4948), .A2(n4945), .ZN(n4944) );
  NAND2_X1 U5372 ( .A1(n4947), .A2(n7776), .ZN(n4943) );
  INV_X1 U5373 ( .A(n7776), .ZN(n4945) );
  INV_X1 U5374 ( .A(n8338), .ZN(n7718) );
  INV_X1 U5375 ( .A(n7190), .ZN(n4939) );
  NAND2_X1 U5376 ( .A1(n4955), .A2(n4957), .ZN(n4952) );
  NAND2_X1 U5377 ( .A1(n4956), .A2(n7700), .ZN(n4955) );
  OR2_X1 U5378 ( .A1(n7870), .A2(n7698), .ZN(n4956) );
  NAND2_X1 U5379 ( .A1(n4957), .A2(n4954), .ZN(n4953) );
  INV_X1 U5380 ( .A(n6835), .ZN(n6833) );
  NAND2_X1 U5381 ( .A1(n8105), .A2(n8106), .ZN(n4563) );
  INV_X1 U5382 ( .A(n8109), .ZN(n4562) );
  AOI21_X1 U5383 ( .B1(n8109), .B2(n8108), .A(n8107), .ZN(n4709) );
  AND4_X1 U5384 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n7084)
         );
  AND4_X1 U5385 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n6829)
         );
  NAND2_X1 U5386 ( .A1(n5819), .A2(n5934), .ZN(n5931) );
  NAND2_X1 U5387 ( .A1(n6819), .A2(n5823), .ZN(n5824) );
  NOR2_X1 U5388 ( .A1(n7062), .A2(n4645), .ZN(n4644) );
  AND2_X1 U5389 ( .A1(n5851), .A2(n5853), .ZN(n7060) );
  NAND2_X1 U5390 ( .A1(n6986), .A2(n4474), .ZN(n5851) );
  NAND2_X1 U5391 ( .A1(n4675), .A2(n4676), .ZN(n4674) );
  INV_X1 U5392 ( .A(n5853), .ZN(n4675) );
  OAI211_X1 U5393 ( .C1(n6978), .C2(n5850), .A(n4646), .B(n4643), .ZN(n7065)
         );
  AOI21_X1 U5394 ( .B1(n7062), .B2(n4645), .A(n7078), .ZN(n4643) );
  NAND2_X1 U5395 ( .A1(n4642), .A2(n7062), .ZN(n5829) );
  NOR2_X1 U5396 ( .A1(n8777), .A2(n7166), .ZN(n7231) );
  NAND2_X1 U5397 ( .A1(n4651), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U5398 ( .A1(n8176), .A2(n4651), .ZN(n4647) );
  INV_X1 U5399 ( .A(n8178), .ZN(n4651) );
  NOR2_X1 U5400 ( .A1(n8274), .A2(n8275), .ZN(n8278) );
  AND2_X1 U5401 ( .A1(n4816), .A2(n8065), .ZN(n4815) );
  NAND2_X1 U5402 ( .A1(n4776), .A2(n4779), .ZN(n4775) );
  NAND2_X1 U5403 ( .A1(n8402), .A2(n4778), .ZN(n4776) );
  NAND2_X1 U5404 ( .A1(n4465), .A2(n5476), .ZN(n4778) );
  INV_X1 U5405 ( .A(n8291), .ZN(n8296) );
  OR2_X1 U5406 ( .A1(n8435), .A2(n8043), .ZN(n4828) );
  AND2_X1 U5407 ( .A1(n8042), .A2(n8411), .ZN(n8428) );
  INV_X1 U5408 ( .A(n8405), .ZN(n8424) );
  AND2_X1 U5409 ( .A1(n8004), .A2(n7984), .ZN(n7929) );
  NAND2_X1 U5410 ( .A1(n6445), .A2(n5278), .ZN(n6553) );
  NAND2_X1 U5411 ( .A1(n4960), .A2(n5242), .ZN(n4959) );
  OAI21_X1 U5412 ( .B1(n8346), .B2(n5544), .A(n4493), .ZN(n8336) );
  AND2_X1 U5413 ( .A1(n5205), .A2(n5204), .ZN(n8349) );
  NAND2_X1 U5414 ( .A1(n8367), .A2(n8366), .ZN(n4817) );
  OR2_X1 U5415 ( .A1(n8890), .A2(n8371), .ZN(n5513) );
  NAND2_X1 U5416 ( .A1(n8414), .A2(n4467), .ZN(n4766) );
  NAND2_X1 U5417 ( .A1(n5218), .A2(n5217), .ZN(n8826) );
  INV_X1 U5418 ( .A(n5385), .ZN(n4764) );
  AND2_X1 U5419 ( .A1(n5636), .A2(n8103), .ZN(n8466) );
  NAND2_X1 U5420 ( .A1(n7045), .A2(n6969), .ZN(n10270) );
  AND2_X1 U5421 ( .A1(n5623), .A2(n5622), .ZN(n7961) );
  INV_X1 U5422 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5624) );
  NOR2_X1 U5423 ( .A1(n5158), .A2(n5157), .ZN(n5159) );
  INV_X1 U5424 ( .A(n5374), .ZN(n4979) );
  INV_X1 U5425 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5482) );
  INV_X1 U5426 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U5427 ( .A1(n5833), .A2(n4598), .ZN(n4664) );
  INV_X1 U5428 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4598) );
  INV_X1 U5429 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5257) );
  XNOR2_X1 U5430 ( .A(n4652), .B(P2_IR_REG_1__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U5431 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4652) );
  NAND2_X1 U5432 ( .A1(n6091), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6098) );
  AND2_X1 U5433 ( .A1(n9085), .A2(n9161), .ZN(n4931) );
  INV_X1 U5434 ( .A(n9272), .ZN(n9447) );
  NAND2_X1 U5435 ( .A1(n4624), .A2(n6463), .ZN(n4915) );
  INV_X1 U5436 ( .A(n6477), .ZN(n4624) );
  NAND2_X1 U5437 ( .A1(n9055), .A2(n9191), .ZN(n9194) );
  INV_X1 U5438 ( .A(n4915), .ZN(n4916) );
  OAI21_X1 U5439 ( .B1(n9141), .B2(n4927), .A(n4925), .ZN(n9036) );
  INV_X1 U5440 ( .A(n4926), .ZN(n4925) );
  NAND2_X1 U5441 ( .A1(n9141), .A2(n9142), .ZN(n9140) );
  OAI211_X1 U5442 ( .C1(n4433), .C2(n6509), .A(n6171), .B(n9660), .ZN(n9122)
         );
  NAND2_X1 U5443 ( .A1(n6171), .A2(n6137), .ZN(n5045) );
  AND2_X1 U5444 ( .A1(n8956), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U5445 ( .A1(n4909), .A2(n7123), .ZN(n4908) );
  OR2_X1 U5446 ( .A1(n8958), .A2(n8959), .ZN(n8956) );
  INV_X1 U5447 ( .A(n7108), .ZN(n4909) );
  INV_X1 U5448 ( .A(n9180), .ZN(n4903) );
  AOI21_X1 U5449 ( .B1(n4901), .B2(n4904), .A(n4527), .ZN(n4900) );
  AND2_X1 U5450 ( .A1(n9248), .A2(n9245), .ZN(n9069) );
  OAI22_X1 U5451 ( .A1(n6128), .A2(n7445), .B1(n7319), .B2(n10091), .ZN(n6129)
         );
  BUF_X1 U5452 ( .A(n6180), .Z(n7296) );
  XNOR2_X1 U5453 ( .A(n5797), .B(n8626), .ZN(n6020) );
  AOI21_X1 U5454 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9789), .A(n9784), .ZN(
        n9889) );
  NOR2_X1 U5455 ( .A1(n9689), .A2(n4535), .ZN(n9476) );
  NAND2_X1 U5456 ( .A1(n4592), .A2(n9533), .ZN(n4535) );
  AND2_X1 U5457 ( .A1(n7486), .A2(n9469), .ZN(n9493) );
  NAND2_X1 U5458 ( .A1(n9533), .A2(n4592), .ZN(n9486) );
  NAND2_X1 U5459 ( .A1(n4507), .A2(n4451), .ZN(n5037) );
  NAND2_X1 U5460 ( .A1(n4473), .A2(n9455), .ZN(n5039) );
  AND2_X1 U5461 ( .A1(n4451), .A2(n9455), .ZN(n5038) );
  NAND2_X1 U5462 ( .A1(n9564), .A2(n4844), .ZN(n4846) );
  AND2_X1 U5463 ( .A1(n7459), .A2(n9464), .ZN(n9566) );
  NAND2_X1 U5464 ( .A1(n9440), .A2(n9439), .ZN(n9572) );
  NOR2_X1 U5465 ( .A1(n9635), .A2(n4838), .ZN(n4837) );
  AND2_X1 U5466 ( .A1(n7635), .A2(n7640), .ZN(n9623) );
  NAND2_X1 U5467 ( .A1(n7293), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7329) );
  INV_X1 U5468 ( .A(n9840), .ZN(n4566) );
  NOR2_X1 U5469 ( .A1(n9984), .A2(n9417), .ZN(n5024) );
  NAND2_X1 U5470 ( .A1(n6087), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U5471 ( .A1(n4505), .A2(n5031), .ZN(n5026) );
  NAND2_X1 U5472 ( .A1(n9995), .A2(n5032), .ZN(n5029) );
  INV_X1 U5473 ( .A(n5020), .ZN(n5018) );
  AND2_X1 U5474 ( .A1(n7518), .A2(n7517), .ZN(n9995) );
  NAND2_X1 U5475 ( .A1(n4988), .A2(n5004), .ZN(n7017) );
  OR2_X1 U5476 ( .A1(n10024), .A2(n9276), .ZN(n5004) );
  NAND2_X1 U5477 ( .A1(n4555), .A2(n7599), .ZN(n9660) );
  NOR2_X1 U5478 ( .A1(n10013), .A2(n10024), .ZN(n10011) );
  NOR2_X1 U5479 ( .A1(n9277), .A2(n10038), .ZN(n5000) );
  NAND2_X1 U5480 ( .A1(n5003), .A2(n7469), .ZN(n5002) );
  OR2_X1 U5481 ( .A1(n4440), .A2(n10089), .ZN(n10080) );
  OR2_X1 U5482 ( .A1(n4434), .A2(n7601), .ZN(n6509) );
  OR2_X1 U5483 ( .A1(n6143), .A2(n7599), .ZN(n6166) );
  INV_X1 U5484 ( .A(n4849), .ZN(n4848) );
  NAND2_X1 U5485 ( .A1(n4851), .A2(n10112), .ZN(n4850) );
  OAI22_X1 U5486 ( .A1(n9474), .A2(n9475), .B1(n9473), .B2(n9472), .ZN(n4849)
         );
  NAND2_X1 U5487 ( .A1(n9689), .A2(n10148), .ZN(n4852) );
  AND2_X1 U5488 ( .A1(n5997), .A2(n6020), .ZN(n6502) );
  AND2_X1 U5489 ( .A1(n6171), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5997) );
  XNOR2_X1 U5490 ( .A(n7253), .B(n7252), .ZN(n8937) );
  OAI21_X1 U5491 ( .B1(n7257), .B2(n7256), .A(n7250), .ZN(n7253) );
  INV_X1 U5492 ( .A(n4986), .ZN(n4985) );
  OR2_X1 U5493 ( .A1(n6014), .A2(n6492), .ZN(n4987) );
  OAI21_X1 U5494 ( .B1(n6015), .B2(n6492), .A(n6024), .ZN(n4986) );
  XNOR2_X1 U5495 ( .A(n5745), .B(SI_28_), .ZN(n5742) );
  AND2_X1 U5496 ( .A1(n5607), .A2(n5591), .ZN(n5605) );
  XNOR2_X1 U5497 ( .A(n6016), .B(n6015), .ZN(n6225) );
  OR2_X1 U5498 ( .A1(n6014), .A2(n6492), .ZN(n6016) );
  XNOR2_X1 U5499 ( .A(n5786), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U5500 ( .A1(n5791), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5786) );
  AND2_X1 U5501 ( .A1(n5792), .A2(n5791), .ZN(n5998) );
  NAND2_X1 U5502 ( .A1(n4885), .A2(n5129), .ZN(n5478) );
  OAI21_X1 U5503 ( .B1(n6661), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6682) );
  XNOR2_X1 U5504 ( .A(n5418), .B(n5417), .ZN(n7273) );
  OAI21_X1 U5505 ( .B1(n5372), .B2(n4698), .A(n4695), .ZN(n5418) );
  AOI21_X1 U5506 ( .B1(n4697), .B2(n4702), .A(n4696), .ZN(n4695) );
  INV_X1 U5507 ( .A(n5103), .ZN(n4696) );
  OR2_X1 U5508 ( .A1(n6116), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6122) );
  INV_X1 U5509 ( .A(SI_5_), .ZN(n5073) );
  INV_X1 U5510 ( .A(n5060), .ZN(n5245) );
  INV_X1 U5511 ( .A(n7905), .ZN(n5800) );
  INV_X1 U5512 ( .A(n8360), .ZN(n7750) );
  INV_X1 U5513 ( .A(n7734), .ZN(n4964) );
  AOI21_X1 U5514 ( .B1(n4967), .B2(n4966), .A(n4484), .ZN(n4965) );
  AND4_X1 U5515 ( .A1(n5224), .A2(n5223), .A3(n5222), .A4(n5221), .ZN(n8423)
         );
  INV_X1 U5516 ( .A(n8328), .ZN(n8348) );
  AND2_X1 U5517 ( .A1(n6766), .A2(n6596), .ZN(n6597) );
  AND4_X1 U5518 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n8394)
         );
  NAND2_X1 U5519 ( .A1(n5616), .A2(n5615), .ZN(n8320) );
  INV_X1 U5520 ( .A(n7826), .ZN(n8440) );
  NAND4_X1 U5521 ( .A1(n5429), .A2(n5428), .A3(n5427), .A4(n5426), .ZN(n8465)
         );
  INV_X1 U5522 ( .A(n7084), .ZN(n8129) );
  INV_X1 U5523 ( .A(n6829), .ZN(n8131) );
  OR2_X1 U5524 ( .A1(n5249), .A2(n6548), .ZN(n5251) );
  NAND2_X1 U5525 ( .A1(n6932), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6976) );
  OR2_X1 U5526 ( .A1(n7220), .A2(n8842), .ZN(n4650) );
  NOR2_X1 U5527 ( .A1(n8454), .A2(n8186), .ZN(n8219) );
  INV_X1 U5528 ( .A(n8207), .ZN(n4635) );
  AND2_X1 U5529 ( .A1(n8280), .A2(n8287), .ZN(n4682) );
  NOR2_X1 U5530 ( .A1(n4680), .A2(n4679), .ZN(n4678) );
  INV_X1 U5531 ( .A(n8277), .ZN(n4680) );
  INV_X1 U5532 ( .A(n8278), .ZN(n4679) );
  NAND2_X1 U5533 ( .A1(n4762), .A2(n8461), .ZN(n4761) );
  INV_X1 U5534 ( .A(n7182), .ZN(n10227) );
  INV_X2 U5535 ( .A(n10233), .ZN(n8489) );
  NAND2_X1 U5536 ( .A1(n5762), .A2(n5763), .ZN(n5764) );
  INV_X1 U5537 ( .A(n7951), .ZN(n7672) );
  INV_X1 U5538 ( .A(n8909), .ZN(n8930) );
  NAND2_X1 U5539 ( .A1(n10275), .A2(n10244), .ZN(n8909) );
  AND2_X1 U5540 ( .A1(n5660), .A2(n5659), .ZN(n8936) );
  AND2_X1 U5541 ( .A1(n4612), .A2(n4472), .ZN(n9150) );
  NAND2_X1 U5542 ( .A1(n9228), .A2(n9227), .ZN(n4612) );
  NAND2_X1 U5543 ( .A1(n4917), .A2(n6463), .ZN(n6478) );
  AOI21_X1 U5544 ( .B1(n7660), .B2(n7659), .A(n7658), .ZN(n7661) );
  OR2_X1 U5545 ( .A1(n6074), .A2(n6073), .ZN(n8963) );
  OR2_X1 U5546 ( .A1(n6488), .A2(n6487), .ZN(n9279) );
  NAND2_X1 U5547 ( .A1(n9687), .A2(n10058), .ZN(n4534) );
  NAND2_X1 U5548 ( .A1(n7007), .A2(n7006), .ZN(n10002) );
  NAND2_X1 U5549 ( .A1(n10058), .A2(n10023), .ZN(n9621) );
  NAND2_X1 U5550 ( .A1(n4731), .A2(n7608), .ZN(n4730) );
  NAND2_X1 U5551 ( .A1(n4732), .A2(n4480), .ZN(n4731) );
  NAND2_X1 U5552 ( .A1(n10055), .A2(n7609), .ZN(n4732) );
  NOR2_X1 U5553 ( .A1(n8012), .A2(n7989), .ZN(n8005) );
  NOR2_X1 U5554 ( .A1(n4738), .A2(n4737), .ZN(n7512) );
  NOR2_X1 U5555 ( .A1(n7504), .A2(n7600), .ZN(n4738) );
  AND2_X1 U5556 ( .A1(n10016), .A2(n7506), .ZN(n4735) );
  INV_X1 U5557 ( .A(n8033), .ZN(n4722) );
  INV_X1 U5558 ( .A(n8473), .ZN(n4717) );
  OAI21_X1 U5559 ( .B1(n4728), .B2(n7619), .A(n7525), .ZN(n4727) );
  AOI21_X1 U5560 ( .B1(n7520), .B2(n7620), .A(n7619), .ZN(n4725) );
  NAND2_X1 U5561 ( .A1(n4689), .A2(n8428), .ZN(n4688) );
  NAND2_X1 U5562 ( .A1(n8040), .A2(n8103), .ZN(n4690) );
  NAND2_X1 U5563 ( .A1(n8041), .A2(n8096), .ZN(n4691) );
  INV_X1 U5564 ( .A(n4551), .ZN(n4550) );
  AOI21_X1 U5565 ( .B1(n7546), .B2(n9622), .A(n7600), .ZN(n4551) );
  NOR2_X1 U5566 ( .A1(n7547), .A2(n9589), .ZN(n4552) );
  NAND2_X1 U5567 ( .A1(n8053), .A2(n8103), .ZN(n4716) );
  INV_X1 U5568 ( .A(n8058), .ZN(n4714) );
  NOR2_X1 U5569 ( .A1(n9460), .A2(n4734), .ZN(n4748) );
  INV_X1 U5570 ( .A(n7557), .ZN(n4749) );
  NAND2_X1 U5571 ( .A1(n7549), .A2(n7556), .ZN(n4750) );
  AOI21_X1 U5572 ( .B1(n4753), .B2(n4752), .A(n9818), .ZN(n4751) );
  NAND2_X1 U5573 ( .A1(n7538), .A2(n7600), .ZN(n4752) );
  AOI21_X1 U5574 ( .B1(n8078), .B2(n8096), .A(n8337), .ZN(n4694) );
  AOI21_X1 U5575 ( .B1(n7566), .B2(n7400), .A(n7574), .ZN(n7424) );
  NAND2_X1 U5576 ( .A1(n4504), .A2(n5666), .ZN(n4983) );
  AND2_X1 U5577 ( .A1(n5624), .A2(n4980), .ZN(n4978) );
  INV_X1 U5578 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5419) );
  INV_X1 U5579 ( .A(n9213), .ZN(n4616) );
  INV_X1 U5580 ( .A(n9227), .ZN(n4609) );
  OR2_X1 U5581 ( .A1(n7570), .A2(n4742), .ZN(n4741) );
  OR2_X1 U5582 ( .A1(n7645), .A2(n4743), .ZN(n4742) );
  OR2_X1 U5583 ( .A1(n7569), .A2(n4734), .ZN(n4743) );
  NAND2_X1 U5584 ( .A1(n4861), .A2(n4859), .ZN(n7582) );
  NOR2_X1 U5585 ( .A1(n7453), .A2(n4860), .ZN(n4859) );
  INV_X1 U5586 ( .A(n7260), .ZN(n4860) );
  NOR2_X1 U5587 ( .A1(n9445), .A2(n5014), .ZN(n5013) );
  INV_X1 U5588 ( .A(n5016), .ZN(n5014) );
  NOR2_X1 U5589 ( .A1(n9674), .A2(n4588), .ZN(n4587) );
  INV_X1 U5590 ( .A(n4589), .ZN(n4588) );
  NAND2_X1 U5591 ( .A1(n4869), .A2(n4868), .ZN(n7243) );
  AOI21_X1 U5592 ( .B1(n4871), .B2(n4873), .A(n4530), .ZN(n4868) );
  AND2_X1 U5593 ( .A1(n6345), .A2(n4855), .ZN(n6012) );
  AND2_X1 U5594 ( .A1(n5040), .A2(n5049), .ZN(n4855) );
  AND2_X1 U5595 ( .A1(n4515), .A2(n5781), .ZN(n5040) );
  INV_X1 U5596 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5785) );
  NOR2_X1 U5597 ( .A1(n5477), .A2(n4884), .ZN(n4883) );
  INV_X1 U5598 ( .A(n5129), .ZN(n4884) );
  NOR2_X1 U5599 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5774) );
  INV_X1 U5600 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5082) );
  NOR2_X1 U5601 ( .A1(n7760), .A2(n7210), .ZN(n4605) );
  INV_X1 U5602 ( .A(n7208), .ZN(n4603) );
  NAND2_X1 U5603 ( .A1(n5256), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U5604 ( .A1(n5256), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U5605 ( .A1(n5930), .A2(n5842), .ZN(n5843) );
  OAI21_X1 U5606 ( .B1(n8219), .B2(n4666), .A(n4665), .ZN(n8272) );
  NAND2_X1 U5607 ( .A1(n8224), .A2(n8246), .ZN(n4665) );
  NAND2_X1 U5608 ( .A1(n4667), .A2(n8246), .ZN(n4666) );
  INV_X1 U5609 ( .A(n8220), .ZN(n4667) );
  INV_X1 U5610 ( .A(SI_17_), .ZN(n8629) );
  OR2_X1 U5611 ( .A1(n5378), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5394) );
  INV_X1 U5612 ( .A(n5308), .ZN(n4754) );
  NAND2_X1 U5613 ( .A1(n4755), .A2(n4478), .ZN(n4756) );
  INV_X1 U5614 ( .A(n5326), .ZN(n4755) );
  INV_X1 U5615 ( .A(n5307), .ZN(n4757) );
  INV_X1 U5616 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U5617 ( .A1(n4962), .A2(n4961), .ZN(n4960) );
  NAND2_X1 U5618 ( .A1(n5241), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4962) );
  NAND2_X1 U5619 ( .A1(n8942), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4961) );
  INV_X1 U5620 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5057) );
  NAND2_X1 U5621 ( .A1(n4506), .A2(n4446), .ZN(n4789) );
  AND2_X1 U5622 ( .A1(n4446), .A2(n4469), .ZN(n4790) );
  INV_X1 U5623 ( .A(n8465), .ZN(n5694) );
  INV_X1 U5624 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5647) );
  INV_X1 U5625 ( .A(n5167), .ZN(n5646) );
  AND2_X1 U5626 ( .A1(n5159), .A2(n4978), .ZN(n4975) );
  INV_X1 U5627 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U5628 ( .A1(n4600), .A2(n4918), .ZN(n7034) );
  AOI21_X1 U5629 ( .B1(n6737), .B2(n4919), .A(n4497), .ZN(n4918) );
  NAND2_X1 U5630 ( .A1(n6736), .A2(n4919), .ZN(n4600) );
  NOR2_X1 U5631 ( .A1(n7034), .A2(n7033), .ZN(n7099) );
  OR2_X1 U5632 ( .A1(n7593), .A2(n9407), .ZN(n7654) );
  INV_X1 U5633 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8626) );
  AOI21_X1 U5634 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9907), .A(n9902), .ZN(
        n9917) );
  AOI21_X1 U5635 ( .B1(n9911), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9916), .ZN(
        n9371) );
  NOR2_X1 U5636 ( .A1(n9928), .A2(n9361), .ZN(n9946) );
  INV_X1 U5637 ( .A(n6510), .ZN(n7485) );
  INV_X1 U5638 ( .A(n9458), .ZN(n5035) );
  NAND2_X1 U5639 ( .A1(n7259), .A2(n7425), .ZN(n4861) );
  OR2_X1 U5640 ( .A1(n9692), .A2(n9474), .ZN(n7486) );
  NOR2_X1 U5641 ( .A1(n9692), .A2(n4593), .ZN(n4592) );
  INV_X1 U5642 ( .A(n4594), .ZN(n4593) );
  NOR2_X1 U5643 ( .A1(n9697), .A2(n9703), .ZN(n4594) );
  NOR2_X1 U5644 ( .A1(n5012), .A2(n5009), .ZN(n5008) );
  INV_X1 U5645 ( .A(n9439), .ZN(n5009) );
  INV_X1 U5646 ( .A(n5013), .ZN(n5012) );
  NAND2_X1 U5647 ( .A1(n5013), .A2(n5011), .ZN(n5010) );
  INV_X1 U5648 ( .A(n5048), .ZN(n5011) );
  OR2_X1 U5649 ( .A1(n4578), .A2(n9423), .ZN(n7535) );
  INV_X1 U5650 ( .A(n10019), .ZN(n4989) );
  NAND2_X1 U5651 ( .A1(n10162), .A2(n6886), .ZN(n5005) );
  INV_X1 U5652 ( .A(n5005), .ZN(n4995) );
  AND2_X1 U5653 ( .A1(n4596), .A2(n10155), .ZN(n4595) );
  AND2_X1 U5654 ( .A1(n10141), .A2(n6884), .ZN(n4596) );
  AND2_X1 U5655 ( .A1(n10129), .A2(n10064), .ZN(n6512) );
  NAND2_X1 U5656 ( .A1(n6694), .A2(n10135), .ZN(n7496) );
  XNOR2_X1 U5657 ( .A(n4559), .B(n10124), .ZN(n7466) );
  INV_X1 U5658 ( .A(n9282), .ZN(n4559) );
  NAND2_X1 U5659 ( .A1(n9617), .A2(n9613), .ZN(n9607) );
  NOR2_X1 U5660 ( .A1(n9828), .A2(n9825), .ZN(n9829) );
  AND2_X1 U5661 ( .A1(n10004), .A2(n4586), .ZN(n9843) );
  AND2_X1 U5662 ( .A1(n4587), .A2(n9868), .ZN(n4586) );
  NAND2_X1 U5663 ( .A1(n10004), .A2(n4587), .ZN(n9842) );
  NAND2_X1 U5664 ( .A1(n10004), .A2(n10183), .ZN(n9985) );
  NOR2_X1 U5665 ( .A1(n10003), .A2(n10002), .ZN(n10004) );
  INV_X1 U5666 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6015) );
  AND2_X1 U5667 ( .A1(n5587), .A2(n5572), .ZN(n5585) );
  AND2_X1 U5668 ( .A1(n5547), .A2(n5532), .ZN(n5545) );
  INV_X1 U5669 ( .A(n5465), .ZN(n4572) );
  INV_X1 U5670 ( .A(SI_15_), .ZN(n5114) );
  INV_X1 U5671 ( .A(n4880), .ZN(n4879) );
  OAI21_X1 U5672 ( .B1(n4881), .B2(n5103), .A(n5109), .ZN(n4880) );
  NAND2_X1 U5673 ( .A1(n4882), .A2(n5108), .ZN(n4881) );
  AND2_X1 U5674 ( .A1(n5113), .A2(n5112), .ZN(n5432) );
  INV_X1 U5675 ( .A(n4866), .ZN(n4865) );
  INV_X1 U5676 ( .A(SI_1_), .ZN(n4875) );
  INV_X1 U5677 ( .A(n7724), .ZN(n4948) );
  INV_X1 U5678 ( .A(n4973), .ZN(n4966) );
  XNOR2_X1 U5679 ( .A(n6537), .B(n5886), .ZN(n5887) );
  NAND2_X1 U5680 ( .A1(n7869), .A2(n7870), .ZN(n7868) );
  INV_X1 U5681 ( .A(n7853), .ZN(n7891) );
  INV_X1 U5682 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5191) );
  AND4_X1 U5683 ( .A1(n5210), .A2(n5209), .A3(n5208), .A4(n5207), .ZN(n7826)
         );
  NAND2_X1 U5684 ( .A1(n6403), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U5685 ( .A1(n5839), .A2(n6400), .ZN(n5927) );
  AND2_X1 U5686 ( .A1(n4661), .A2(n6809), .ZN(n6751) );
  NAND2_X1 U5687 ( .A1(n4663), .A2(n4662), .ZN(n4661) );
  INV_X1 U5688 ( .A(n5843), .ZN(n4663) );
  AND2_X1 U5689 ( .A1(n6815), .A2(n4640), .ZN(n6747) );
  INV_X1 U5690 ( .A(n5821), .ZN(n4641) );
  NAND2_X1 U5691 ( .A1(n6751), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6811) );
  AND2_X1 U5692 ( .A1(n6982), .A2(n4658), .ZN(n6935) );
  INV_X1 U5693 ( .A(n5847), .ZN(n4660) );
  NAND2_X1 U5694 ( .A1(n6986), .A2(n5849), .ZN(n4856) );
  NAND2_X1 U5695 ( .A1(n7060), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7059) );
  AOI22_X1 U5696 ( .A1(n7057), .A2(n7058), .B1(n5850), .B2(n5811), .ZN(n7156)
         );
  AND2_X1 U5697 ( .A1(n4668), .A2(n4673), .ZN(n7164) );
  INV_X1 U5698 ( .A(n4672), .ZN(n4668) );
  OR2_X1 U5699 ( .A1(n7231), .A2(n7232), .ZN(n8144) );
  NAND2_X1 U5700 ( .A1(n8144), .A2(n8145), .ZN(n8143) );
  AND2_X1 U5701 ( .A1(n4450), .A2(n5213), .ZN(n5420) );
  NAND2_X1 U5702 ( .A1(n7223), .A2(n7224), .ZN(n8151) );
  XNOR2_X1 U5703 ( .A(n8158), .B(n8174), .ZN(n7234) );
  AND2_X1 U5704 ( .A1(n8143), .A2(n4857), .ZN(n8158) );
  NAND2_X1 U5705 ( .A1(n7233), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4857) );
  XNOR2_X1 U5706 ( .A(n8272), .B(n8273), .ZN(n8248) );
  AND2_X1 U5707 ( .A1(n8233), .A2(n8232), .ZN(n8256) );
  NAND2_X1 U5708 ( .A1(n5536), .A2(n5535), .ZN(n5558) );
  INV_X1 U5709 ( .A(n5537), .ZN(n5536) );
  OR2_X1 U5710 ( .A1(n5520), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U5711 ( .A1(n5187), .A2(n5186), .ZN(n5497) );
  INV_X1 U5712 ( .A(n5486), .ZN(n5187) );
  OR2_X1 U5713 ( .A1(n5497), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5508) );
  OAI21_X1 U5714 ( .B1(n8435), .B2(n4825), .A(n4824), .ZN(n4823) );
  AOI21_X1 U5715 ( .B1(n5699), .B2(n4827), .A(n5698), .ZN(n4824) );
  NAND2_X1 U5716 ( .A1(n5699), .A2(n5696), .ZN(n4825) );
  INV_X1 U5717 ( .A(n5220), .ZN(n5185) );
  OR2_X1 U5718 ( .A1(n5443), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U5719 ( .A1(n5416), .A2(n5415), .ZN(n8476) );
  NAND2_X1 U5720 ( .A1(n4763), .A2(n4483), .ZN(n5416) );
  NAND2_X1 U5721 ( .A1(n5181), .A2(n5180), .ZN(n5443) );
  INV_X1 U5722 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5180) );
  INV_X1 U5723 ( .A(n5424), .ZN(n5181) );
  OR2_X1 U5724 ( .A1(n5394), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U5725 ( .A1(n5179), .A2(n7799), .ZN(n5424) );
  INV_X1 U5726 ( .A(n5409), .ZN(n5179) );
  AND4_X1 U5727 ( .A1(n5362), .A2(n5361), .A3(n5360), .A4(n5359), .ZN(n7051)
         );
  NAND2_X1 U5728 ( .A1(n4811), .A2(n4810), .ZN(n4809) );
  INV_X1 U5729 ( .A(n7072), .ZN(n4811) );
  NAND2_X1 U5730 ( .A1(n5178), .A2(n5177), .ZN(n5378) );
  INV_X1 U5731 ( .A(n5357), .ZN(n5178) );
  NAND2_X1 U5732 ( .A1(n5176), .A2(n5175), .ZN(n5341) );
  INV_X1 U5733 ( .A(n5327), .ZN(n5176) );
  OR2_X1 U5734 ( .A1(n5341), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5357) );
  INV_X1 U5735 ( .A(n8128), .ZN(n7088) );
  OR2_X1 U5736 ( .A1(n5309), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U5737 ( .A1(n6716), .A2(n7930), .ZN(n6775) );
  AND2_X1 U5738 ( .A1(n7999), .A2(n7983), .ZN(n7930) );
  AND3_X1 U5739 ( .A1(n6367), .A2(n10270), .A3(n5705), .ZN(n6719) );
  OR2_X1 U5740 ( .A1(n8878), .A2(n8372), .ZN(n4793) );
  INV_X1 U5741 ( .A(n8381), .ZN(n4768) );
  NAND2_X1 U5742 ( .A1(n4828), .A2(n4826), .ZN(n8427) );
  NAND2_X1 U5743 ( .A1(n4785), .A2(n4789), .ZN(n8437) );
  NAND2_X1 U5744 ( .A1(n4792), .A2(n4790), .ZN(n4785) );
  OAI21_X1 U5745 ( .B1(n8460), .B2(n4788), .A(n4786), .ZN(n8439) );
  NAND2_X1 U5746 ( .A1(n8436), .A2(n4790), .ZN(n4788) );
  NAND2_X1 U5747 ( .A1(n4787), .A2(n8436), .ZN(n4786) );
  INV_X1 U5748 ( .A(n4789), .ZN(n4787) );
  AOI21_X1 U5749 ( .B1(n4821), .B2(n8031), .A(n4819), .ZN(n4818) );
  INV_X1 U5750 ( .A(n4821), .ZN(n4820) );
  INV_X1 U5751 ( .A(n8034), .ZN(n4819) );
  OR2_X1 U5752 ( .A1(n8032), .A2(n8031), .ZN(n8484) );
  INV_X1 U5753 ( .A(n4805), .ZN(n4804) );
  AOI21_X1 U5754 ( .B1(n4805), .B2(n4806), .A(n4803), .ZN(n4802) );
  AOI21_X1 U5755 ( .B1(n4807), .B2(n7933), .A(n4503), .ZN(n4805) );
  NAND2_X1 U5756 ( .A1(n4809), .A2(n4807), .ZN(n7144) );
  XNOR2_X1 U5757 ( .A(n5667), .B(n5666), .ZN(n5901) );
  NAND2_X1 U5758 ( .A1(n5193), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5197) );
  AND2_X1 U5759 ( .A1(n5230), .A2(n5467), .ZN(n8222) );
  NAND2_X1 U5760 ( .A1(n4450), .A2(n4632), .ZN(n5228) );
  OR2_X1 U5761 ( .A1(n5348), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5349) );
  OR2_X1 U5762 ( .A1(n5319), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5348) );
  INV_X1 U5763 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U5764 ( .A1(n4900), .A2(n4899), .ZN(n4898) );
  NOR2_X1 U5765 ( .A1(n7099), .A2(n7035), .ZN(n7036) );
  AND2_X1 U5766 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  AND2_X1 U5767 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  NAND2_X1 U5768 ( .A1(n4916), .A2(n4913), .ZN(n4912) );
  INV_X1 U5769 ( .A(n6458), .ZN(n4913) );
  AND2_X1 U5770 ( .A1(n9056), .A2(n9054), .ZN(n9191) );
  NAND2_X1 U5771 ( .A1(n4625), .A2(n6621), .ZN(n6477) );
  NAND2_X1 U5772 ( .A1(n6475), .A2(n6476), .ZN(n4625) );
  NAND2_X1 U5773 ( .A1(n6462), .A2(n6461), .ZN(n6463) );
  NAND2_X1 U5774 ( .A1(n7107), .A2(n7108), .ZN(n7124) );
  NAND2_X1 U5775 ( .A1(n6273), .A2(n6144), .ZN(n6149) );
  NAND2_X1 U5776 ( .A1(n6149), .A2(n6148), .ZN(n6275) );
  NAND2_X1 U5777 ( .A1(n4622), .A2(n4576), .ZN(n9202) );
  OR2_X1 U5778 ( .A1(n8972), .A2(n8971), .ZN(n4619) );
  NAND2_X1 U5779 ( .A1(n6625), .A2(n6624), .ZN(n6627) );
  NAND2_X1 U5780 ( .A1(n6734), .A2(n6733), .ZN(n6784) );
  INV_X1 U5781 ( .A(n9475), .ZN(n9251) );
  INV_X1 U5782 ( .A(n9406), .ZN(n9250) );
  AND2_X1 U5783 ( .A1(n8990), .A2(n8989), .ZN(n8994) );
  AOI21_X1 U5784 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9814), .A(n9806), .ZN(
        n6249) );
  AND2_X1 U5785 ( .A1(n9927), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U5786 ( .A1(n7295), .A2(n9932), .ZN(n9931) );
  AND2_X1 U5787 ( .A1(n9388), .A2(n4531), .ZN(n9964) );
  NAND2_X1 U5788 ( .A1(n7901), .A2(n7425), .ZN(n4538) );
  AND2_X1 U5789 ( .A1(n9533), .A2(n4594), .ZN(n9503) );
  INV_X1 U5790 ( .A(n4841), .ZN(n4840) );
  OAI21_X1 U5791 ( .B1(n9538), .B2(n9465), .A(n9466), .ZN(n4841) );
  NOR2_X1 U5792 ( .A1(n9550), .A2(n9707), .ZN(n9533) );
  OR2_X1 U5793 ( .A1(n9545), .A2(n9446), .ZN(n9449) );
  NAND2_X1 U5794 ( .A1(n7262), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7389) );
  AND2_X1 U5795 ( .A1(n9617), .A2(n4510), .ZN(n9560) );
  OR2_X1 U5796 ( .A1(n7407), .A2(n9221), .ZN(n7369) );
  NAND2_X1 U5797 ( .A1(n9617), .A2(n4582), .ZN(n9573) );
  INV_X1 U5798 ( .A(n7545), .ZN(n9589) );
  NAND2_X1 U5799 ( .A1(n7640), .A2(n7542), .ZN(n4832) );
  INV_X1 U5800 ( .A(n4835), .ZN(n4834) );
  OAI21_X1 U5801 ( .B1(n4837), .B2(n4836), .A(n9623), .ZN(n4835) );
  NOR2_X1 U5802 ( .A1(n9638), .A2(n9737), .ZN(n9617) );
  AOI22_X1 U5803 ( .A1(n9634), .A2(n9430), .B1(n9429), .B2(n9641), .ZN(n9616)
         );
  OR2_X1 U5804 ( .A1(n7329), .A2(n6090), .ZN(n7330) );
  INV_X1 U5805 ( .A(n5022), .ZN(n5021) );
  OAI21_X1 U5806 ( .B1(n4447), .B2(n4468), .A(n5030), .ZN(n5022) );
  OR2_X1 U5807 ( .A1(n6997), .A2(n6086), .ZN(n6998) );
  AND2_X1 U5808 ( .A1(n4831), .A2(n7516), .ZN(n9994) );
  NAND2_X1 U5809 ( .A1(n9994), .A2(n9995), .ZN(n9993) );
  OR2_X1 U5810 ( .A1(n6871), .A2(n8562), .ZN(n6997) );
  NAND3_X1 U5811 ( .A1(n10051), .A2(n4595), .A3(n10162), .ZN(n10013) );
  OR2_X1 U5812 ( .A1(n10043), .A2(n7615), .ZN(n6700) );
  NAND2_X1 U5813 ( .A1(n10051), .A2(n10141), .ZN(n10050) );
  AND2_X1 U5814 ( .A1(n6512), .A2(n6693), .ZN(n10051) );
  AND2_X1 U5815 ( .A1(n7492), .A2(n7609), .ZN(n10061) );
  NAND3_X1 U5816 ( .A1(n4853), .A2(n4558), .A3(n4557), .ZN(n6656) );
  OR2_X1 U5817 ( .A1(n6847), .A2(n6309), .ZN(n4557) );
  OR2_X1 U5818 ( .A1(n7439), .A2(n6308), .ZN(n4558) );
  NOR2_X1 U5819 ( .A1(n10080), .A2(n6656), .ZN(n10064) );
  INV_X1 U5820 ( .A(n7466), .ZN(n6649) );
  BUF_X1 U5821 ( .A(n6515), .Z(n10070) );
  NAND2_X1 U5822 ( .A1(n7415), .A2(n7425), .ZN(n7418) );
  INV_X1 U5823 ( .A(n9641), .ZN(n9851) );
  INV_X1 U5824 ( .A(n4578), .ZN(n9862) );
  INV_X1 U5825 ( .A(n10194), .ZN(n10148) );
  NAND2_X1 U5826 ( .A1(n10088), .A2(n6509), .ZN(n10194) );
  INV_X1 U5827 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6034) );
  AND2_X1 U5828 ( .A1(n5528), .A2(n5150), .ZN(n5526) );
  NAND2_X1 U5829 ( .A1(n6135), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6018) );
  AND2_X1 U5830 ( .A1(n4514), .A2(n4453), .ZN(n4933) );
  AND2_X1 U5831 ( .A1(n6346), .A2(n5781), .ZN(n6493) );
  XNOR2_X1 U5832 ( .A(n5451), .B(n5450), .ZN(n7288) );
  INV_X1 U5833 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U5834 ( .A1(n4699), .A2(n4697), .ZN(n5403) );
  XNOR2_X1 U5835 ( .A(n5079), .B(n5078), .ZN(n5335) );
  OR2_X1 U5836 ( .A1(n6215), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5994) );
  XNOR2_X1 U5837 ( .A(n5069), .B(SI_4_), .ZN(n5286) );
  INV_X1 U5838 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5984) );
  XNOR2_X1 U5839 ( .A(n5066), .B(SI_3_), .ZN(n5273) );
  INV_X1 U5840 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5979) );
  XNOR2_X1 U5841 ( .A(n5063), .B(SI_2_), .ZN(n5254) );
  NAND2_X1 U5842 ( .A1(n6947), .A2(n4444), .ZN(n7085) );
  AND2_X1 U5843 ( .A1(n6947), .A2(n6946), .ZN(n6950) );
  AND2_X1 U5844 ( .A1(n5593), .A2(n5592), .ZN(n7732) );
  OAI21_X1 U5845 ( .B1(n4574), .B2(n7690), .A(n4973), .ZN(n7738) );
  NAND2_X1 U5846 ( .A1(n4606), .A2(n8126), .ZN(n7759) );
  NAND2_X1 U5847 ( .A1(n7868), .A2(n4954), .ZN(n7769) );
  NAND2_X1 U5848 ( .A1(n4942), .A2(n4946), .ZN(n4941) );
  NAND2_X1 U5849 ( .A1(n7779), .A2(n7776), .ZN(n4946) );
  AOI21_X1 U5850 ( .B1(n4448), .B2(n4953), .A(n4502), .ZN(n4949) );
  NAND2_X1 U5851 ( .A1(n4448), .A2(n7869), .ZN(n4626) );
  NAND2_X1 U5852 ( .A1(n4937), .A2(n6765), .ZN(n6831) );
  NAND2_X1 U5853 ( .A1(n6764), .A2(n6766), .ZN(n4937) );
  NAND2_X1 U5854 ( .A1(n7815), .A2(n8423), .ZN(n7694) );
  OR2_X1 U5855 ( .A1(n7815), .A2(n8423), .ZN(n7693) );
  NAND2_X1 U5856 ( .A1(n4951), .A2(n4952), .ZN(n7842) );
  OR2_X1 U5857 ( .A1(n7869), .A2(n4953), .ZN(n4951) );
  INV_X1 U5858 ( .A(n4936), .ZN(n4935) );
  OAI21_X1 U5859 ( .B1(n4938), .B2(n6766), .A(n6830), .ZN(n4936) );
  AND2_X1 U5860 ( .A1(n5602), .A2(n5601), .ZN(n7881) );
  OR2_X1 U5861 ( .A1(n5916), .A2(n5915), .ZN(n7893) );
  NAND2_X1 U5862 ( .A1(n5911), .A2(n8444), .ZN(n7883) );
  NAND2_X1 U5863 ( .A1(n4970), .A2(n4971), .ZN(n7888) );
  AND2_X1 U5864 ( .A1(n4970), .A2(n4967), .ZN(n7886) );
  NAND2_X1 U5865 ( .A1(n4574), .A2(n4973), .ZN(n4970) );
  INV_X1 U5866 ( .A(n7821), .ZN(n7895) );
  AOI21_X1 U5867 ( .B1(n4567), .B2(n7950), .A(n4495), .ZN(n8112) );
  XNOR2_X1 U5868 ( .A(n5619), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8118) );
  INV_X1 U5869 ( .A(n7881), .ZN(n8329) );
  NAND2_X1 U5870 ( .A1(n5581), .A2(n5580), .ZN(n8338) );
  NAND2_X1 U5871 ( .A1(n5564), .A2(n5563), .ZN(n8328) );
  INV_X1 U5872 ( .A(n8349), .ZN(n8372) );
  OAI211_X1 U5873 ( .C1(n5249), .C2(n8591), .A(n5522), .B(n5521), .ZN(n8385)
         );
  INV_X1 U5874 ( .A(n8393), .ZN(n8371) );
  INV_X1 U5875 ( .A(n8394), .ZN(n8415) );
  INV_X1 U5876 ( .A(n7051), .ZN(n8127) );
  AND2_X1 U5877 ( .A1(n6974), .A2(n4638), .ZN(n6932) );
  INV_X1 U5878 ( .A(n5824), .ZN(n4639) );
  NAND2_X1 U5879 ( .A1(n5829), .A2(n4646), .ZN(n7063) );
  NOR2_X1 U5880 ( .A1(n7218), .A2(n4564), .ZN(n7162) );
  AND2_X1 U5881 ( .A1(n7161), .A2(n7167), .ZN(n4564) );
  NAND2_X1 U5882 ( .A1(n7162), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8139) );
  INV_X1 U5883 ( .A(n8176), .ZN(n4649) );
  OR2_X1 U5884 ( .A1(n8225), .A2(n8224), .ZN(n8247) );
  NOR2_X1 U5885 ( .A1(n8219), .A2(n8220), .ZN(n8225) );
  AND2_X1 U5886 ( .A1(n4637), .A2(n4471), .ZN(n8208) );
  OR2_X1 U5887 ( .A1(P2_U3150), .A2(n5861), .ZN(n8300) );
  OR2_X1 U5888 ( .A1(n8285), .A2(n8284), .ZN(n4656) );
  NAND2_X1 U5889 ( .A1(n4817), .A2(n4815), .ZN(n5054) );
  NAND2_X1 U5890 ( .A1(n8414), .A2(n4466), .ZN(n4772) );
  NAND2_X1 U5891 ( .A1(n7337), .A2(n7900), .ZN(n4532) );
  NAND2_X1 U5892 ( .A1(n4777), .A2(n4465), .ZN(n8403) );
  OR2_X1 U5893 ( .A1(n8414), .A2(n5476), .ZN(n4777) );
  NAND2_X1 U5894 ( .A1(n6715), .A2(n5307), .ZN(n4758) );
  INV_X1 U5895 ( .A(n8783), .ZN(n8486) );
  OAI22_X1 U5896 ( .A1(n5972), .A2(n5549), .B1(P1_DATAO_REG_1__SCAN_IN), .B2(
        n7904), .ZN(n4794) );
  INV_X1 U5897 ( .A(n8431), .ZN(n10226) );
  NAND2_X1 U5898 ( .A1(n8935), .A2(n5729), .ZN(n8444) );
  OAI22_X1 U5899 ( .A1(n5741), .A2(n5740), .B1(n8106), .B2(n8095), .ZN(n5749)
         );
  NOR2_X1 U5900 ( .A1(n5770), .A2(n8461), .ZN(n4760) );
  NAND2_X1 U5901 ( .A1(n4537), .A2(n4536), .ZN(n7906) );
  NAND2_X1 U5902 ( .A1(n4443), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n4536) );
  NAND2_X1 U5903 ( .A1(n8937), .A2(n7904), .ZN(n4537) );
  INV_X1 U5904 ( .A(n7732), .ZN(n8855) );
  OR2_X1 U5905 ( .A1(n5746), .A2(n8953), .ZN(n5573) );
  OR2_X1 U5906 ( .A1(n5746), .A2(n7176), .ZN(n5554) );
  INV_X1 U5907 ( .A(n7839), .ZN(n8872) );
  NAND2_X1 U5908 ( .A1(n4817), .A2(n8065), .ZN(n8357) );
  AND2_X1 U5909 ( .A1(n4791), .A2(n4470), .ZN(n8450) );
  NAND2_X1 U5910 ( .A1(n4792), .A2(n4469), .ZN(n4791) );
  NAND2_X1 U5911 ( .A1(n5423), .A2(n5422), .ZN(n8929) );
  NAND2_X1 U5912 ( .A1(n4763), .A2(n4464), .ZN(n7195) );
  AND2_X1 U5913 ( .A1(n5370), .A2(n5369), .ZN(n7182) );
  INV_X2 U5914 ( .A(n10277), .ZN(n10275) );
  AND2_X1 U5915 ( .A1(n5902), .A2(n5991), .ZN(n8935) );
  INV_X1 U5916 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U5917 ( .A1(n5642), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5644) );
  INV_X1 U5918 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8573) );
  INV_X1 U5919 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6968) );
  INV_X1 U5920 ( .A(n7961), .ZN(n6969) );
  XNOR2_X1 U5921 ( .A(n5625), .B(n5624), .ZN(n8100) );
  XNOR2_X1 U5922 ( .A(n5483), .B(n5482), .ZN(n8291) );
  INV_X1 U5923 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6119) );
  INV_X1 U5924 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5986) );
  INV_X1 U5925 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5971) );
  INV_X1 U5926 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U5927 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4664), .ZN(n5258) );
  NAND2_X1 U5928 ( .A1(n6784), .A2(n6783), .ZN(n7028) );
  NAND2_X1 U5929 ( .A1(n7124), .A2(n7123), .ZN(n8957) );
  NAND2_X1 U5930 ( .A1(n4893), .A2(n4895), .ZN(n9113) );
  OR2_X1 U5931 ( .A1(n9168), .A2(n4898), .ZN(n4893) );
  NAND2_X1 U5932 ( .A1(n9085), .A2(n4930), .ZN(n4929) );
  INV_X1 U5933 ( .A(n9069), .ZN(n4930) );
  INV_X1 U5934 ( .A(n10047), .ZN(n10141) );
  INV_X1 U5935 ( .A(n6736), .ZN(n6734) );
  AOI21_X1 U5936 ( .B1(n9168), .B2(n9000), .A(n4904), .ZN(n9182) );
  NAND2_X1 U5937 ( .A1(n4917), .A2(n4916), .ZN(n6622) );
  NAND2_X1 U5938 ( .A1(n4620), .A2(n4619), .ZN(n9214) );
  NAND2_X1 U5939 ( .A1(n4614), .A2(n4613), .ZN(n4620) );
  INV_X1 U5940 ( .A(n9149), .ZN(n4613) );
  INV_X1 U5941 ( .A(n9150), .ZN(n4614) );
  NAND2_X1 U5942 ( .A1(n9036), .A2(n4630), .ZN(n9219) );
  NAND2_X1 U5943 ( .A1(n9140), .A2(n4924), .ZN(n4630) );
  AND2_X1 U5944 ( .A1(n9035), .A2(n9032), .ZN(n4924) );
  AOI21_X1 U5946 ( .B1(n4907), .B2(n4910), .A(n4452), .ZN(n4905) );
  NAND2_X1 U5947 ( .A1(n4901), .A2(n9168), .ZN(n4894) );
  INV_X1 U5948 ( .A(n9222), .ZN(n9262) );
  OR2_X1 U5949 ( .A1(n6189), .A2(n6167), .ZN(n9268) );
  AND2_X1 U5950 ( .A1(n6176), .A2(n6175), .ZN(n9264) );
  INV_X1 U5951 ( .A(n8994), .ZN(n9260) );
  INV_X1 U5952 ( .A(n9258), .ZN(n9266) );
  AND3_X1 U5953 ( .A1(n6043), .A2(n6042), .A3(n6041), .ZN(n9472) );
  OR2_X1 U5954 ( .A1(n7313), .A2(n7312), .ZN(n9273) );
  OR2_X1 U5955 ( .A1(n6066), .A2(n6065), .ZN(n7111) );
  INV_X1 U5956 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5352) );
  OR2_X1 U5957 ( .A1(n7445), .A2(n6182), .ZN(n6183) );
  OR2_X1 U5958 ( .A1(n7443), .A2(n6127), .ZN(n6131) );
  NAND2_X1 U5959 ( .A1(n5798), .A2(n6020), .ZN(n9284) );
  AOI21_X1 U5960 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9802), .A(n9794), .ZN(
        n9808) );
  AND2_X1 U5961 ( .A1(n6194), .A2(n6125), .ZN(n9789) );
  AOI21_X1 U5962 ( .B1(n9968), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9957), .ZN(
        n9387) );
  INV_X1 U5963 ( .A(n7593), .ZN(n9678) );
  NAND2_X1 U5964 ( .A1(n5033), .A2(n5037), .ZN(n9485) );
  AND2_X1 U5965 ( .A1(n4846), .A2(n9465), .ZN(n9537) );
  INV_X1 U5966 ( .A(n9713), .ZN(n9556) );
  NAND2_X1 U5967 ( .A1(n5015), .A2(n5016), .ZN(n9559) );
  NAND2_X1 U5968 ( .A1(n9572), .A2(n5048), .ZN(n5015) );
  NAND2_X1 U5969 ( .A1(n4833), .A2(n7542), .ZN(n9624) );
  NAND2_X1 U5970 ( .A1(n9821), .A2(n4837), .ZN(n4833) );
  NAND2_X1 U5971 ( .A1(n9821), .A2(n7631), .ZN(n9631) );
  NAND2_X1 U5972 ( .A1(n5025), .A2(n5023), .ZN(n9659) );
  INV_X1 U5973 ( .A(n5024), .ZN(n5023) );
  NAND2_X1 U5974 ( .A1(n5027), .A2(n4447), .ZN(n5025) );
  NAND2_X1 U5975 ( .A1(n7275), .A2(n7274), .ZN(n9984) );
  NAND2_X1 U5976 ( .A1(n5027), .A2(n5026), .ZN(n9983) );
  NAND2_X1 U5977 ( .A1(n5028), .A2(n5032), .ZN(n9416) );
  OR2_X1 U5978 ( .A1(n9991), .A2(n9995), .ZN(n5028) );
  NAND2_X1 U5979 ( .A1(n6684), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U5980 ( .A1(n4990), .A2(n4991), .ZN(n10010) );
  NAND2_X1 U5981 ( .A1(n4997), .A2(n4999), .ZN(n6904) );
  NAND2_X1 U5982 ( .A1(n6885), .A2(n5001), .ZN(n4997) );
  INV_X1 U5983 ( .A(n5002), .ZN(n5001) );
  AOI21_X1 U5984 ( .B1(n6885), .B2(n7469), .A(n5006), .ZN(n10030) );
  NAND2_X1 U5985 ( .A1(n9679), .A2(n6502), .ZN(n10090) );
  OR2_X1 U5986 ( .A1(n7439), .A2(n4877), .ZN(n6266) );
  AND2_X1 U5987 ( .A1(n10058), .A2(n6507), .ZN(n10097) );
  AND3_X2 U5988 ( .A1(n9743), .A2(n9742), .A3(n9681), .ZN(n10221) );
  INV_X1 U5989 ( .A(n9688), .ZN(n4565) );
  AND3_X2 U5990 ( .A1(n9743), .A2(n9742), .A3(n9741), .ZN(n10201) );
  NAND2_X1 U5991 ( .A1(n6502), .A2(n6165), .ZN(n10110) );
  NAND2_X1 U5992 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6027), .ZN(n6028) );
  OR2_X1 U5993 ( .A1(n6026), .A2(n6027), .ZN(n6029) );
  INV_X1 U5994 ( .A(n6039), .ZN(n9767) );
  NAND2_X1 U5995 ( .A1(n5606), .A2(n5605), .ZN(n4870) );
  CLKBUF_X1 U5996 ( .A(n6225), .Z(n9404) );
  INV_X1 U5997 ( .A(n5998), .ZN(n7177) );
  INV_X1 U5998 ( .A(n4433), .ZN(n9685) );
  INV_X1 U5999 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7402) );
  INV_X1 U6000 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7416) );
  INV_X1 U6001 ( .A(n4434), .ZN(n6507) );
  XNOR2_X1 U6002 ( .A(n6195), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9895) );
  INV_X1 U6003 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U6004 ( .A1(n4864), .A2(n5075), .ZN(n5322) );
  NAND2_X1 U6005 ( .A1(n5299), .A2(n5298), .ZN(n4864) );
  INV_X1 U6006 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6464) );
  INV_X1 U6007 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6415) );
  NOR2_X2 U6008 ( .A1(n5858), .A2(P2_U3151), .ZN(P2_U3893) );
  INV_X1 U6009 ( .A(n4650), .ZN(n8175) );
  OAI211_X1 U6010 ( .C1(n8281), .C2(n8310), .A(n4681), .B(n4677), .ZN(P2_U3200) );
  OAI21_X1 U6011 ( .B1(n8303), .B2(n4678), .A(n8148), .ZN(n4677) );
  NOR2_X1 U6012 ( .A1(n4682), .A2(n8279), .ZN(n4681) );
  AND2_X1 U6013 ( .A1(n4761), .A2(n5053), .ZN(n7669) );
  INV_X1 U6014 ( .A(n5737), .ZN(n5738) );
  OAI21_X1 U6015 ( .B1(n5736), .B2(n8783), .A(n5735), .ZN(n5737) );
  INV_X1 U6016 ( .A(n5707), .ZN(n5708) );
  OAI21_X1 U6017 ( .B1(n5736), .B2(n8837), .A(n5706), .ZN(n5707) );
  NOR2_X1 U6018 ( .A1(n5765), .A2(n5767), .ZN(n5768) );
  INV_X1 U6019 ( .A(n5723), .ZN(n5724) );
  OAI21_X1 U6020 ( .B1(n5736), .B2(n8919), .A(n5722), .ZN(n5723) );
  OR2_X1 U6021 ( .A1(n7666), .A2(n7665), .ZN(n4541) );
  OAI21_X1 U6022 ( .B1(n9483), .B2(n9630), .A(n4534), .ZN(n4533) );
  AND2_X1 U6023 ( .A1(n6949), .A2(n6946), .ZN(n4444) );
  OR2_X1 U6024 ( .A1(n4454), .A2(n7887), .ZN(n4445) );
  NAND2_X1 U6025 ( .A1(n6788), .A2(n6787), .ZN(n10038) );
  AOI21_X1 U6026 ( .B1(n5003), .B2(n5006), .A(n5000), .ZN(n4999) );
  OR2_X1 U6027 ( .A1(n8916), .A2(n8464), .ZN(n4446) );
  INV_X1 U6028 ( .A(n8451), .ZN(n4972) );
  AND2_X1 U6029 ( .A1(n5049), .A2(n5781), .ZN(n5042) );
  INV_X2 U6030 ( .A(n5235), .ZN(n5343) );
  AND2_X1 U6031 ( .A1(n5026), .A2(n9973), .ZN(n4447) );
  INV_X1 U6032 ( .A(n5827), .ZN(n4645) );
  AND2_X1 U6033 ( .A1(n4952), .A2(n4950), .ZN(n4448) );
  XOR2_X1 U6034 ( .A(n8305), .B(n8304), .Z(n4449) );
  AND3_X1 U6035 ( .A1(n5154), .A2(n5256), .A3(n4633), .ZN(n4450) );
  OR2_X1 U6036 ( .A1(n9697), .A2(n9456), .ZN(n4451) );
  AND2_X1 U6037 ( .A1(n8958), .A2(n8959), .ZN(n4452) );
  AND2_X1 U6038 ( .A1(n5781), .A2(n8557), .ZN(n4453) );
  INV_X1 U6039 ( .A(n6836), .ZN(n6832) );
  INV_X1 U6040 ( .A(n7933), .ZN(n4810) );
  AND2_X1 U6041 ( .A1(n4942), .A2(n4487), .ZN(n4454) );
  AND2_X1 U6042 ( .A1(n8101), .A2(n4800), .ZN(n4455) );
  NAND2_X1 U6043 ( .A1(n4438), .A2(n9421), .ZN(n4456) );
  OR2_X1 U6044 ( .A1(n9464), .A2(n4734), .ZN(n4457) );
  INV_X1 U6045 ( .A(n9674), .ZN(n10195) );
  NAND2_X1 U6046 ( .A1(n7281), .A2(n7280), .ZN(n9674) );
  NAND2_X1 U6047 ( .A1(n4773), .A2(n4766), .ZN(n8380) );
  AND2_X1 U6048 ( .A1(n8942), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4458) );
  OR2_X1 U6049 ( .A1(n5326), .A2(n4754), .ZN(n4459) );
  INV_X1 U6050 ( .A(n4783), .ZN(n4782) );
  INV_X1 U6051 ( .A(n7791), .ZN(n8404) );
  AND4_X1 U6052 ( .A1(n5502), .A2(n5501), .A3(n5500), .A4(n5499), .ZN(n7791)
         );
  AND2_X1 U6053 ( .A1(n4676), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4460) );
  AND2_X1 U6054 ( .A1(n4460), .A2(n4671), .ZN(n4461) );
  INV_X1 U6055 ( .A(n7599), .ZN(n4922) );
  INV_X1 U6056 ( .A(n6190), .ZN(n4555) );
  AND2_X1 U6057 ( .A1(n10051), .A2(n4596), .ZN(n4462) );
  NAND2_X1 U6058 ( .A1(n7920), .A2(n8083), .ZN(n4463) );
  OR2_X1 U6059 ( .A1(n4556), .A2(n8125), .ZN(n4464) );
  INV_X1 U6060 ( .A(n6281), .ZN(n7360) );
  OR2_X1 U6061 ( .A1(n7877), .A2(n8424), .ZN(n4465) );
  INV_X1 U6062 ( .A(n7706), .ZN(n8878) );
  INV_X2 U6063 ( .A(n5756), .ZN(n7913) );
  NAND2_X1 U6064 ( .A1(n6581), .A2(n6298), .ZN(n5884) );
  AND2_X1 U6065 ( .A1(n4779), .A2(n4465), .ZN(n4466) );
  AND2_X1 U6066 ( .A1(n8391), .A2(n4466), .ZN(n4467) );
  NOR2_X1 U6067 ( .A1(n5098), .A2(n4704), .ZN(n4703) );
  OR2_X1 U6068 ( .A1(n9420), .A2(n5024), .ZN(n4468) );
  INV_X1 U6069 ( .A(n5850), .ZN(n7062) );
  OR2_X1 U6070 ( .A1(n8923), .A2(n8451), .ZN(n4469) );
  INV_X1 U6071 ( .A(n9464), .ZN(n4845) );
  NAND2_X1 U6072 ( .A1(n8923), .A2(n8451), .ZN(n4470) );
  NAND2_X1 U6073 ( .A1(n5639), .A2(n5161), .ZN(n5642) );
  OR2_X1 U6074 ( .A1(n8218), .A2(n8203), .ZN(n4471) );
  NAND2_X1 U6075 ( .A1(n8966), .A2(n8965), .ZN(n4472) );
  NOR2_X1 U6076 ( .A1(n9519), .A2(n9454), .ZN(n4473) );
  AND2_X1 U6077 ( .A1(n5849), .A2(n5850), .ZN(n4474) );
  NAND2_X1 U6078 ( .A1(n7357), .A2(n7356), .ZN(n9717) );
  INV_X1 U6079 ( .A(n9717), .ZN(n4581) );
  AND3_X1 U6080 ( .A1(n8104), .A2(n8103), .A3(n8102), .ZN(n4475) );
  NAND2_X1 U6081 ( .A1(n9091), .A2(n8985), .ZN(n9168) );
  AND2_X1 U6082 ( .A1(n7462), .A2(n7502), .ZN(n4476) );
  AND2_X1 U6083 ( .A1(n9564), .A2(n9464), .ZN(n4477) );
  AND2_X1 U6084 ( .A1(n5308), .A2(n4757), .ZN(n4478) );
  NAND2_X1 U6085 ( .A1(n4975), .A2(n4979), .ZN(n5620) );
  OR2_X1 U6086 ( .A1(n8861), .A2(n8338), .ZN(n4479) );
  INV_X1 U6087 ( .A(n7542), .ZN(n4836) );
  NAND2_X1 U6088 ( .A1(n7367), .A2(n7366), .ZN(n9723) );
  INV_X1 U6089 ( .A(n9156), .ZN(n10183) );
  NAND2_X1 U6090 ( .A1(n6994), .A2(n6993), .ZN(n9156) );
  INV_X1 U6091 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5405) );
  INV_X1 U6092 ( .A(n9733), .ZN(n9613) );
  NAND2_X1 U6093 ( .A1(n7418), .A2(n7417), .ZN(n9733) );
  AND2_X1 U6094 ( .A1(n7496), .A2(n7492), .ZN(n4480) );
  NOR2_X1 U6095 ( .A1(n7027), .A2(n4920), .ZN(n4919) );
  AND2_X1 U6096 ( .A1(n8786), .A2(n7947), .ZN(n4481) );
  INV_X1 U6097 ( .A(n4703), .ZN(n4702) );
  AND2_X1 U6098 ( .A1(n7526), .A2(n7529), .ZN(n9982) );
  OR2_X1 U6099 ( .A1(n4725), .A2(n4724), .ZN(n4482) );
  INV_X1 U6100 ( .A(n4827), .ZN(n4826) );
  NAND2_X1 U6101 ( .A1(n8428), .A2(n8044), .ZN(n4827) );
  AND2_X1 U6102 ( .A1(n5050), .A2(n4464), .ZN(n4483) );
  AND2_X1 U6103 ( .A1(n7692), .A2(n8464), .ZN(n4484) );
  NAND2_X1 U6104 ( .A1(n5647), .A2(n5162), .ZN(n4485) );
  AND2_X1 U6105 ( .A1(n8127), .A2(n10227), .ZN(n4486) );
  NAND2_X1 U6106 ( .A1(n4861), .A2(n7260), .ZN(n9689) );
  INV_X1 U6107 ( .A(n9689), .ZN(n4591) );
  NAND2_X1 U6108 ( .A1(n4947), .A2(n4948), .ZN(n4487) );
  INV_X1 U6109 ( .A(n7779), .ZN(n4947) );
  OR2_X1 U6110 ( .A1(n5387), .A2(SI_11_), .ZN(n4488) );
  AND2_X1 U6111 ( .A1(n7084), .A2(n7083), .ZN(n4489) );
  NAND2_X1 U6112 ( .A1(n9692), .A2(n9457), .ZN(n4490) );
  NAND3_X1 U6113 ( .A1(n4979), .A2(n5159), .A3(n4980), .ZN(n4491) );
  NAND2_X1 U6114 ( .A1(n6346), .A2(n5042), .ZN(n4492) );
  OR2_X1 U6115 ( .A1(n8872), .A2(n7750), .ZN(n4493) );
  AND2_X1 U6116 ( .A1(n9868), .A2(n9422), .ZN(n4494) );
  AND2_X1 U6117 ( .A1(n8786), .A2(n7949), .ZN(n4495) );
  AND2_X1 U6118 ( .A1(n4756), .A2(n5325), .ZN(n4496) );
  INV_X1 U6119 ( .A(n4698), .ZN(n4697) );
  NAND2_X1 U6120 ( .A1(n4700), .A2(n4705), .ZN(n4698) );
  AND2_X1 U6121 ( .A1(n7026), .A2(n7025), .ZN(n4497) );
  AND2_X1 U6122 ( .A1(n5077), .A2(SI_6_), .ZN(n4498) );
  INV_X1 U6123 ( .A(n4611), .ZN(n4610) );
  NAND2_X1 U6124 ( .A1(n4472), .A2(n4617), .ZN(n4611) );
  AND2_X1 U6125 ( .A1(n4616), .A2(n4618), .ZN(n4499) );
  AND2_X1 U6126 ( .A1(n7688), .A2(n4972), .ZN(n4500) );
  OR2_X1 U6127 ( .A1(n4581), .A2(n9444), .ZN(n4501) );
  INV_X1 U6128 ( .A(n8370), .ZN(n8366) );
  AND2_X1 U6129 ( .A1(n5524), .A2(n5523), .ZN(n8370) );
  AND2_X1 U6130 ( .A1(n7701), .A2(n7791), .ZN(n4502) );
  OR2_X1 U6131 ( .A1(n4813), .A2(n4812), .ZN(n4503) );
  AND2_X1 U6132 ( .A1(n5161), .A2(n4984), .ZN(n4504) );
  NAND2_X1 U6133 ( .A1(n9415), .A2(n5029), .ZN(n4505) );
  INV_X1 U6134 ( .A(n6765), .ZN(n4938) );
  NAND2_X1 U6135 ( .A1(n5464), .A2(n4470), .ZN(n4506) );
  NAND2_X1 U6136 ( .A1(n9508), .A2(n5039), .ZN(n4507) );
  NAND2_X1 U6137 ( .A1(n6136), .A2(n6135), .ZN(n10092) );
  NAND2_X1 U6138 ( .A1(n7583), .A2(n7582), .ZN(n9470) );
  INV_X1 U6139 ( .A(n9470), .ZN(n4745) );
  AND2_X1 U6140 ( .A1(n8352), .A2(n8071), .ZN(n4508) );
  AND2_X1 U6141 ( .A1(n4991), .A2(n4989), .ZN(n4509) );
  AND2_X1 U6142 ( .A1(n4582), .A2(n4581), .ZN(n4510) );
  NOR2_X1 U6143 ( .A1(n5400), .A2(n4764), .ZN(n4511) );
  AND2_X1 U6144 ( .A1(n7186), .A2(n4939), .ZN(n4512) );
  AND2_X1 U6145 ( .A1(n7706), .A2(n8372), .ZN(n8070) );
  INV_X1 U6146 ( .A(n8070), .ZN(n4816) );
  AND2_X1 U6147 ( .A1(n9690), .A2(n4852), .ZN(n4513) );
  NOR2_X1 U6148 ( .A1(n5794), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n4514) );
  AND2_X1 U6149 ( .A1(n5785), .A2(n5041), .ZN(n4515) );
  AND2_X1 U6150 ( .A1(n4941), .A2(n7871), .ZN(n4516) );
  AND2_X1 U6151 ( .A1(n4501), .A2(n5010), .ZN(n4517) );
  INV_X1 U6152 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4980) );
  AND2_X1 U6153 ( .A1(n5618), .A2(n4830), .ZN(n5192) );
  INV_X1 U6154 ( .A(n6004), .ZN(n4659) );
  NAND2_X1 U6155 ( .A1(n9991), .A2(n5018), .ZN(n5027) );
  INV_X1 U6156 ( .A(n8126), .ZN(n7210) );
  INV_X1 U6157 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4877) );
  INV_X1 U6158 ( .A(n4823), .ZN(n8401) );
  NAND2_X1 U6159 ( .A1(n5386), .A2(n5385), .ZN(n7146) );
  NAND2_X1 U6160 ( .A1(n4894), .A2(n4900), .ZN(n9235) );
  INV_X1 U6161 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4984) );
  AND2_X1 U6162 ( .A1(n9016), .A2(n9015), .ZN(n4518) );
  NAND2_X1 U6163 ( .A1(n7187), .A2(n7186), .ZN(n7188) );
  OR2_X1 U6164 ( .A1(n9825), .A2(n9427), .ZN(n7631) );
  INV_X1 U6165 ( .A(n7631), .ZN(n4838) );
  AND2_X1 U6166 ( .A1(n4809), .A2(n8008), .ZN(n4519) );
  NAND2_X1 U6167 ( .A1(n9617), .A2(n4584), .ZN(n4585) );
  AND2_X1 U6168 ( .A1(n4772), .A2(n4775), .ZN(n4520) );
  INV_X1 U6169 ( .A(n9236), .ZN(n4899) );
  INV_X1 U6170 ( .A(n9418), .ZN(n9419) );
  OR2_X1 U6171 ( .A1(n7286), .A2(n7285), .ZN(n9418) );
  AND2_X1 U6172 ( .A1(n4650), .A2(n4649), .ZN(n4521) );
  OR2_X1 U6173 ( .A1(n5864), .A2(n5852), .ZN(n4522) );
  NAND2_X1 U6174 ( .A1(n5225), .A2(SI_16_), .ZN(n4523) );
  INV_X1 U6175 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5193) );
  AND2_X1 U6176 ( .A1(n4523), .A2(n5117), .ZN(n4524) );
  AND2_X1 U6177 ( .A1(n4828), .A2(n8044), .ZN(n4525) );
  OR2_X1 U6178 ( .A1(n4606), .A2(n8126), .ZN(n4526) );
  INV_X1 U6179 ( .A(n7167), .ZN(n4671) );
  INV_X1 U6180 ( .A(n7887), .ZN(n7871) );
  NAND2_X1 U6181 ( .A1(n6597), .A2(n6598), .ZN(n6764) );
  AND2_X1 U6182 ( .A1(n8118), .A2(n7961), .ZN(n8103) );
  OR2_X1 U6183 ( .A1(n6899), .A2(n7989), .ZN(n6898) );
  NAND2_X1 U6184 ( .A1(n4758), .A2(n5308), .ZN(n6777) );
  XNOR2_X1 U6185 ( .A(n5644), .B(n4984), .ZN(n5658) );
  AND2_X1 U6186 ( .A1(n9006), .A2(n9005), .ZN(n4527) );
  NAND2_X1 U6187 ( .A1(n6833), .A2(n6832), .ZN(n6947) );
  AND2_X1 U6188 ( .A1(n4674), .A2(n4673), .ZN(n4528) );
  NOR2_X1 U6189 ( .A1(n10289), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4529) );
  AND2_X1 U6190 ( .A1(n5745), .A2(n5744), .ZN(n4530) );
  NAND2_X1 U6191 ( .A1(n10051), .A2(n4595), .ZN(n4597) );
  NAND2_X1 U6192 ( .A1(n10004), .A2(n4589), .ZN(n4590) );
  INV_X1 U6193 ( .A(n7123), .ZN(n4910) );
  AND2_X1 U6194 ( .A1(n5713), .A2(n8113), .ZN(n8477) );
  OR2_X1 U6195 ( .A1(n9389), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4531) );
  AND2_X1 U6196 ( .A1(n5885), .A2(n5882), .ZN(n5051) );
  AND2_X2 U6197 ( .A1(n5727), .A2(n5684), .ZN(n10289) );
  XNOR2_X1 U6198 ( .A(n5272), .B(n5271), .ZN(n6400) );
  INV_X1 U6199 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5175) );
  NAND2_X1 U6200 ( .A1(n10026), .A2(n10092), .ZN(n6190) );
  NAND2_X1 U6201 ( .A1(n6805), .A2(n6804), .ZN(n6803) );
  AOI21_X1 U6202 ( .B1(n5805), .B2(n6754), .A(n6744), .ZN(n6805) );
  INV_X1 U6203 ( .A(n6754), .ZN(n4662) );
  NAND2_X1 U6204 ( .A1(n5124), .A2(n5123), .ZN(n5466) );
  NAND2_X1 U6205 ( .A1(n4759), .A2(n4544), .ZN(n5772) );
  OAI21_X2 U6206 ( .B1(n5402), .B2(n4881), .A(n4879), .ZN(n5433) );
  NAND2_X1 U6207 ( .A1(n5434), .A2(n5113), .ZN(n5451) );
  OR2_X1 U6208 ( .A1(n9482), .A2(n4533), .ZN(P1_U3356) );
  NAND2_X1 U6209 ( .A1(n5433), .A2(n5432), .ZN(n5434) );
  NAND2_X1 U6210 ( .A1(n5529), .A2(n5528), .ZN(n5546) );
  OAI21_X1 U6211 ( .B1(n7649), .B2(n9407), .A(n7593), .ZN(n7596) );
  AOI21_X1 U6212 ( .B1(n7484), .B2(n7485), .A(n4434), .ZN(n4570) );
  AOI21_X1 U6213 ( .B1(n4801), .B2(n4455), .A(n4481), .ZN(n8114) );
  OR2_X1 U6214 ( .A1(n8114), .A2(n8113), .ZN(n4706) );
  NAND2_X1 U6215 ( .A1(n4888), .A2(n5120), .ZN(n5212) );
  NAND2_X1 U6216 ( .A1(n5060), .A2(n5244), .ZN(n4568) );
  NAND2_X1 U6217 ( .A1(n5606), .A2(n4871), .ZN(n4869) );
  OAI21_X1 U6218 ( .B1(n9000), .B2(n4904), .A(n4903), .ZN(n4902) );
  NAND2_X1 U6219 ( .A1(n4542), .A2(n4541), .ZN(P1_U3242) );
  NAND2_X1 U6220 ( .A1(n4543), .A2(n6174), .ZN(n4542) );
  OAI21_X1 U6221 ( .B1(n7663), .B2(n7662), .A(n7661), .ZN(n4543) );
  AOI21_X1 U6222 ( .B1(n7648), .B2(n7647), .A(n7646), .ZN(n7652) );
  AOI21_X1 U6223 ( .B1(n7640), .B2(n7639), .A(n7638), .ZN(n7644) );
  NAND2_X1 U6224 ( .A1(n7572), .A2(n7571), .ZN(n4746) );
  NAND2_X1 U6225 ( .A1(n5586), .A2(n5585), .ZN(n5588) );
  OAI21_X2 U6226 ( .B1(n8335), .B2(n8081), .A(n8079), .ZN(n8326) );
  NAND3_X1 U6227 ( .A1(n5761), .A2(n4429), .A3(n10289), .ZN(n4544) );
  AOI21_X2 U6228 ( .B1(n4740), .B2(n4545), .A(n7595), .ZN(n7603) );
  NAND2_X1 U6229 ( .A1(n5364), .A2(n5363), .ZN(n4874) );
  NAND2_X1 U6230 ( .A1(n5274), .A2(n5273), .ZN(n4546) );
  NAND2_X1 U6231 ( .A1(n8370), .A2(n4815), .ZN(n4547) );
  OAI211_X1 U6232 ( .C1(n8111), .C2(n8110), .A(n4709), .B(n4708), .ZN(n4707)
         );
  NAND2_X1 U6233 ( .A1(n4850), .A2(n4848), .ZN(n9687) );
  OAI21_X2 U6234 ( .B1(n9604), .B2(n9461), .A(n9460), .ZN(n9580) );
  AND2_X1 U6235 ( .A1(n7515), .A2(n10016), .ZN(n7510) );
  NAND2_X1 U6236 ( .A1(n9565), .A2(n9566), .ZN(n9564) );
  NAND2_X1 U6237 ( .A1(n4568), .A2(n5062), .ZN(n5255) );
  NAND2_X1 U6238 ( .A1(n4548), .A2(n5065), .ZN(n5274) );
  NAND2_X1 U6239 ( .A1(n9645), .A2(n9646), .ZN(n9644) );
  NAND2_X1 U6240 ( .A1(n4839), .A2(n4840), .ZN(n9525) );
  INV_X1 U6241 ( .A(n9687), .ZN(n4847) );
  NOR2_X1 U6242 ( .A1(n10024), .A2(n6916), .ZN(n6887) );
  NAND2_X1 U6243 ( .A1(n6909), .A2(n4476), .ZN(n7612) );
  NOR2_X1 U6244 ( .A1(n9584), .A2(n9463), .ZN(n9565) );
  NAND2_X1 U6245 ( .A1(n5255), .A2(n5254), .ZN(n4548) );
  NAND2_X1 U6246 ( .A1(n4579), .A2(n7567), .ZN(n7573) );
  NOR2_X1 U6247 ( .A1(n4749), .A2(n4748), .ZN(n4747) );
  OR4_X2 U6248 ( .A1(n4463), .A2(n8337), .A3(n8354), .A4(n7944), .ZN(n7945) );
  NAND2_X1 U6249 ( .A1(n9202), .A2(n9203), .ZN(n9201) );
  NAND2_X1 U6250 ( .A1(n6682), .A2(n8593), .ZN(n6684) );
  NAND2_X1 U6251 ( .A1(n7107), .A2(n4907), .ZN(n4906) );
  OAI21_X2 U6252 ( .B1(n9228), .B2(n4611), .A(n4607), .ZN(n8984) );
  INV_X1 U6253 ( .A(n4891), .ZN(n4890) );
  NOR2_X1 U6254 ( .A1(n9219), .A2(n9220), .ZN(n9103) );
  NAND2_X1 U6255 ( .A1(n7598), .A2(n4434), .ZN(n4571) );
  INV_X1 U6256 ( .A(n4775), .ZN(n4774) );
  NAND2_X1 U6257 ( .A1(n4761), .A2(n4429), .ZN(n5771) );
  NAND2_X1 U6258 ( .A1(n4773), .A2(n4771), .ZN(n4770) );
  OAI21_X1 U6259 ( .B1(n8336), .B2(n7921), .A(n7922), .ZN(n8327) );
  NAND2_X1 U6260 ( .A1(n4571), .A2(n4569), .ZN(n7663) );
  NAND3_X1 U6261 ( .A1(n4706), .A2(n8112), .A3(n4707), .ZN(n8115) );
  AOI21_X2 U6262 ( .B1(n4964), .B2(n4967), .A(n4963), .ZN(n7817) );
  INV_X1 U6263 ( .A(n4968), .ZN(n4967) );
  NAND2_X1 U6264 ( .A1(n6813), .A2(n5846), .ZN(n5847) );
  NAND2_X1 U6265 ( .A1(n4660), .A2(n4659), .ZN(n4658) );
  NAND2_X1 U6266 ( .A1(n6646), .A2(n7466), .ZN(n4854) );
  XNOR2_X1 U6267 ( .A(n9471), .B(n4745), .ZN(n4851) );
  OAI22_X2 U6268 ( .A1(n9821), .A2(n4832), .B1(n4834), .B2(n7550), .ZN(n9604)
         );
  NAND3_X1 U6269 ( .A1(n8024), .A2(n8025), .A3(n8023), .ZN(n8030) );
  NAND2_X1 U6270 ( .A1(n8038), .A2(n4561), .ZN(n4560) );
  NAND2_X1 U6271 ( .A1(n8077), .A2(n8103), .ZN(n4693) );
  NAND2_X1 U6272 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  AOI21_X1 U6273 ( .B1(n8054), .B2(n8096), .A(n8059), .ZN(n4715) );
  OAI21_X1 U6274 ( .B1(n4692), .B2(n4463), .A(n8087), .ZN(n8091) );
  NAND3_X1 U6275 ( .A1(n4563), .A2(n4562), .A3(n4475), .ZN(n4708) );
  OR2_X2 U6276 ( .A1(n7725), .A2(n7724), .ZN(n7777) );
  NAND2_X1 U6277 ( .A1(n4971), .A2(n4969), .ZN(n4968) );
  XNOR2_X2 U6278 ( .A(n7211), .B(n7778), .ZN(n7682) );
  NAND2_X1 U6279 ( .A1(n4639), .A2(n4659), .ZN(n4638) );
  NAND2_X1 U6280 ( .A1(n4641), .A2(n4662), .ZN(n4640) );
  INV_X1 U6281 ( .A(n8208), .ZN(n4636) );
  NOR2_X1 U6282 ( .A1(n8257), .A2(n8258), .ZN(n8260) );
  OAI21_X1 U6283 ( .B1(n7220), .B2(n4648), .A(n4647), .ZN(n8192) );
  NAND2_X4 U6284 ( .A1(n6786), .A2(n7904), .ZN(n7439) );
  NAND3_X1 U6285 ( .A1(n4513), .A2(n4847), .A3(n4565), .ZN(n9746) );
  NAND2_X1 U6286 ( .A1(n4509), .A2(n4990), .ZN(n4988) );
  AOI21_X1 U6287 ( .B1(n6650), .B2(n6649), .A(n6499), .ZN(n10062) );
  XNOR2_X2 U6288 ( .A(n5982), .B(n5981), .ZN(n6267) );
  AOI22_X2 U6289 ( .A1(n7017), .A2(n7016), .B1(n7015), .B2(n10172), .ZN(n9991)
         );
  NAND4_X1 U6290 ( .A1(n7948), .A2(n8101), .A3(n8104), .A4(n8099), .ZN(n4567)
         );
  NAND2_X1 U6291 ( .A1(n6575), .A2(n5056), .ZN(n4711) );
  NAND2_X1 U6292 ( .A1(n5136), .A2(n5135), .ZN(n5505) );
  NAND2_X1 U6293 ( .A1(n5139), .A2(n5138), .ZN(n4878) );
  OR4_X1 U6294 ( .A1(n9526), .A2(n7480), .A3(n9538), .A4(n9544), .ZN(n7481) );
  NAND2_X1 U6295 ( .A1(n7585), .A2(n7584), .ZN(n4739) );
  NAND2_X1 U6296 ( .A1(n7878), .A2(n7718), .ZN(n4621) );
  NAND2_X1 U6297 ( .A1(n7158), .A2(n7157), .ZN(n7223) );
  AOI21_X1 U6298 ( .B1(n7725), .B2(n7724), .A(n7887), .ZN(n7726) );
  NAND3_X1 U6299 ( .A1(n6598), .A2(n6597), .A3(n6765), .ZN(n4573) );
  OAI22_X2 U6300 ( .A1(n6971), .A2(n6972), .B1(n5809), .B2(n6979), .ZN(n7057)
         );
  AND2_X2 U6301 ( .A1(n5664), .A2(n5666), .ZN(n5639) );
  INV_X1 U6302 ( .A(n5154), .ZN(n4634) );
  INV_X1 U6303 ( .A(n5897), .ZN(n5893) );
  INV_X1 U6304 ( .A(n4858), .ZN(n4654) );
  AOI21_X2 U6305 ( .B1(n5645), .B2(n5658), .A(n4575), .ZN(n5656) );
  INV_X1 U6306 ( .A(n4577), .ZN(n4576) );
  NOR2_X1 U6307 ( .A1(n4891), .A2(n9091), .ZN(n4577) );
  INV_X1 U6308 ( .A(n4902), .ZN(n4901) );
  OAI21_X1 U6309 ( .B1(n8985), .B2(n4891), .A(n4889), .ZN(n4623) );
  NAND2_X1 U6310 ( .A1(n4727), .A2(n4734), .ZN(n4726) );
  OAI21_X1 U6311 ( .B1(n7505), .B2(n4734), .A(n10032), .ZN(n4737) );
  NAND3_X1 U6312 ( .A1(n7565), .A2(n9546), .A3(n4457), .ZN(n4579) );
  AOI21_X1 U6313 ( .B1(n7533), .B2(n7532), .A(n4723), .ZN(n7536) );
  AOI22_X1 U6314 ( .A1(n7537), .A2(n4734), .B1(n7539), .B2(n7540), .ZN(n4753)
         );
  AOI21_X1 U6315 ( .B1(n7524), .B2(n7617), .A(n7523), .ZN(n4728) );
  OAI21_X1 U6316 ( .B1(n4751), .B2(n4750), .A(n4747), .ZN(n7558) );
  INV_X1 U6317 ( .A(n7512), .ZN(n4736) );
  NAND2_X1 U6318 ( .A1(n4736), .A2(n4735), .ZN(n7509) );
  NAND2_X1 U6319 ( .A1(n7493), .A2(n4734), .ZN(n4733) );
  NAND2_X1 U6320 ( .A1(n5845), .A2(n6808), .ZN(n6813) );
  XNOR2_X1 U6321 ( .A(n5839), .B(n4657), .ZN(n6399) );
  OAI21_X1 U6322 ( .B1(n4655), .B2(n8310), .A(n4653), .ZN(P2_U3201) );
  NAND2_X1 U6323 ( .A1(n4895), .A2(n4892), .ZN(n4891) );
  INV_X1 U6324 ( .A(n4623), .ZN(n4622) );
  NAND2_X1 U6325 ( .A1(n4996), .A2(n4994), .ZN(n4990) );
  INV_X1 U6326 ( .A(n4999), .ZN(n4998) );
  NAND2_X2 U6327 ( .A1(n9453), .A2(n9452), .ZN(n9515) );
  AOI21_X2 U6328 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n9802), .A(n9797), .ZN(
        n9811) );
  AOI21_X2 U6329 ( .B1(n9789), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9781), .ZN(
        n9892) );
  AOI21_X2 U6330 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9895), .A(n9890), .ZN(
        n6675) );
  AOI21_X2 U6331 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9814), .A(n9809), .ZN(
        n6233) );
  AOI21_X2 U6332 ( .B1(n9907), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9899), .ZN(
        n9914) );
  INV_X1 U6333 ( .A(n4585), .ZN(n9594) );
  INV_X1 U6334 ( .A(n4590), .ZN(n9986) );
  NAND2_X1 U6335 ( .A1(n9533), .A2(n9519), .ZN(n9516) );
  INV_X1 U6336 ( .A(n4597), .ZN(n10039) );
  NAND2_X1 U6337 ( .A1(n7209), .A2(n4602), .ZN(n4601) );
  XNOR2_X2 U6338 ( .A(n8984), .B(n8982), .ZN(n9093) );
  NAND2_X1 U6339 ( .A1(n8978), .A2(n8977), .ZN(n4618) );
  AND2_X2 U6340 ( .A1(n4628), .A2(n4627), .ZN(n7869) );
  OR2_X2 U6341 ( .A1(n7825), .A2(n4629), .ZN(n4628) );
  NAND2_X1 U6342 ( .A1(n4450), .A2(n4631), .ZN(n5467) );
  OR2_X2 U6343 ( .A1(n5284), .A2(n4634), .ZN(n5374) );
  INV_X1 U6344 ( .A(n4637), .ZN(n8204) );
  NAND2_X1 U6345 ( .A1(n4636), .A2(n4635), .ZN(n8233) );
  XNOR2_X1 U6346 ( .A(n8203), .B(n8218), .ZN(n8194) );
  NAND2_X1 U6347 ( .A1(n6978), .A2(n4644), .ZN(n4646) );
  NAND2_X1 U6348 ( .A1(n6978), .A2(n5827), .ZN(n4642) );
  XNOR2_X1 U6349 ( .A(n8173), .B(n8174), .ZN(n7220) );
  INV_X1 U6350 ( .A(n6400), .ZN(n4657) );
  NAND2_X1 U6351 ( .A1(n6399), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U6352 ( .A1(n6398), .A2(n5927), .ZN(n5841) );
  NAND2_X1 U6353 ( .A1(n7060), .A2(n4460), .ZN(n4673) );
  INV_X1 U6354 ( .A(n5854), .ZN(n4676) );
  NAND3_X1 U6355 ( .A1(n4691), .A2(n4690), .A3(n5696), .ZN(n4689) );
  INV_X2 U6356 ( .A(n7904), .ZN(n5963) );
  MUX2_X1 U6357 ( .A(n6308), .B(n5961), .S(n4430), .Z(n5063) );
  NAND3_X1 U6358 ( .A1(n4722), .A2(n4718), .A3(n4717), .ZN(n8038) );
  INV_X2 U6359 ( .A(n7600), .ZN(n4734) );
  NAND3_X1 U6360 ( .A1(n7586), .A2(n4744), .A3(n4741), .ZN(n4740) );
  AND2_X1 U6361 ( .A1(n4746), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U6362 ( .A1(n6892), .A2(n7989), .ZN(n5340) );
  INV_X1 U6363 ( .A(n5761), .ZN(n4762) );
  NAND2_X1 U6364 ( .A1(n5386), .A2(n4511), .ZN(n4763) );
  OR2_X1 U6365 ( .A1(n8414), .A2(n4770), .ZN(n4765) );
  NAND2_X1 U6366 ( .A1(n4765), .A2(n4767), .ZN(n8384) );
  OAI21_X1 U6367 ( .B1(n6963), .B2(n5355), .A(n5356), .ZN(n7073) );
  NAND2_X1 U6368 ( .A1(n4784), .A2(n5371), .ZN(n4783) );
  AND2_X2 U6369 ( .A1(n5618), .A2(n5160), .ZN(n5664) );
  INV_X1 U6370 ( .A(n8460), .ZN(n4792) );
  NAND2_X1 U6371 ( .A1(n5247), .A2(n4794), .ZN(n4795) );
  NAND2_X1 U6372 ( .A1(n5247), .A2(n4443), .ZN(n5243) );
  NAND2_X1 U6373 ( .A1(n5247), .A2(n7904), .ZN(n5246) );
  NAND3_X1 U6374 ( .A1(n5242), .A2(n5241), .A3(P2_REG3_REG_1__SCAN_IN), .ZN(
        n4796) );
  AND2_X2 U6375 ( .A1(n5241), .A2(n7678), .ZN(n5264) );
  AND2_X2 U6376 ( .A1(n8942), .A2(n7678), .ZN(n5456) );
  NAND3_X1 U6377 ( .A1(n7678), .A2(P2_REG0_REG_1__SCAN_IN), .A3(n8942), .ZN(
        n4797) );
  NAND2_X1 U6378 ( .A1(n5242), .A2(n4458), .ZN(n4798) );
  NAND2_X1 U6379 ( .A1(n5264), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4799) );
  OR2_X1 U6380 ( .A1(n7910), .A2(n7909), .ZN(n4801) );
  OAI21_X2 U6381 ( .B1(n7072), .B2(n4804), .A(n4802), .ZN(n7194) );
  INV_X1 U6382 ( .A(n4815), .ZN(n4814) );
  OAI21_X1 U6383 ( .B1(n8485), .B2(n8032), .A(n7938), .ZN(n8472) );
  AND2_X1 U6384 ( .A1(n5618), .A2(n4829), .ZN(n5196) );
  OAI21_X2 U6385 ( .B1(n8326), .B2(n8085), .A(n8083), .ZN(n8317) );
  NAND2_X1 U6386 ( .A1(n8369), .A2(n8370), .ZN(n8368) );
  NAND2_X1 U6387 ( .A1(n5701), .A2(n8061), .ZN(n8367) );
  NAND2_X1 U6388 ( .A1(n5702), .A2(n8074), .ZN(n8335) );
  NAND2_X1 U6389 ( .A1(n5169), .A2(n5168), .ZN(n5634) );
  NAND2_X1 U6390 ( .A1(n5248), .A2(n10235), .ZN(n7964) );
  NAND3_X1 U6391 ( .A1(n7612), .A2(n7473), .A3(n7616), .ZN(n4831) );
  NAND2_X1 U6392 ( .A1(n6867), .A2(n7462), .ZN(n7616) );
  NAND2_X1 U6393 ( .A1(n9564), .A2(n4842), .ZN(n4839) );
  INV_X1 U6394 ( .A(n4846), .ZN(n9548) );
  OR2_X1 U6395 ( .A1(n6786), .A2(n6310), .ZN(n4853) );
  NAND2_X2 U6396 ( .A1(n6786), .A2(n5963), .ZN(n6847) );
  OAI21_X2 U6397 ( .B1(n10055), .B2(n6521), .A(n7609), .ZN(n7491) );
  NAND2_X1 U6399 ( .A1(n5299), .A2(n4865), .ZN(n4862) );
  NAND2_X2 U6400 ( .A1(n4874), .A2(n5093), .ZN(n5372) );
  OAI21_X2 U6401 ( .B1(n4430), .B2(n4877), .A(n4876), .ZN(n5061) );
  NAND2_X1 U6402 ( .A1(n4885), .A2(n4883), .ZN(n4886) );
  NAND2_X1 U6403 ( .A1(n4887), .A2(n4524), .ZN(n4888) );
  NAND2_X1 U6404 ( .A1(n6459), .A2(n6458), .ZN(n4917) );
  AND2_X1 U6405 ( .A1(n6618), .A2(n4912), .ZN(n4911) );
  OR2_X1 U6406 ( .A1(n6459), .A2(n4915), .ZN(n4914) );
  NAND2_X4 U6407 ( .A1(n4921), .A2(n6171), .ZN(n9075) );
  OAI21_X1 U6408 ( .B1(n9142), .B2(n4927), .A(n9034), .ZN(n4926) );
  INV_X1 U6409 ( .A(n9032), .ZN(n4927) );
  NAND2_X1 U6410 ( .A1(n9160), .A2(n4931), .ZN(n4928) );
  NAND2_X1 U6411 ( .A1(n4928), .A2(n4929), .ZN(n9131) );
  NAND2_X1 U6412 ( .A1(n9131), .A2(n4932), .ZN(n9138) );
  AND2_X1 U6413 ( .A1(n9135), .A2(n9247), .ZN(n4932) );
  NAND2_X1 U6414 ( .A1(n6345), .A2(n4453), .ZN(n6661) );
  NAND2_X1 U6415 ( .A1(n6345), .A2(n4933), .ZN(n6133) );
  OAI211_X1 U6416 ( .C1(n7725), .C2(n4445), .A(n4940), .B(n7786), .ZN(P2_U3160) );
  NAND2_X1 U6417 ( .A1(n7725), .A2(n4516), .ZN(n4940) );
  NAND2_X1 U6418 ( .A1(n5242), .A2(n5241), .ZN(n5235) );
  AOI21_X2 U6419 ( .B1(n4973), .B2(n7690), .A(n4500), .ZN(n4971) );
  AND3_X2 U6420 ( .A1(n4974), .A2(n4976), .A3(n5159), .ZN(n5618) );
  INV_X1 U6421 ( .A(n5374), .ZN(n4974) );
  NAND2_X1 U6422 ( .A1(n6014), .A2(n6015), .ZN(n6030) );
  INV_X1 U6423 ( .A(n6885), .ZN(n4996) );
  AND2_X1 U6424 ( .A1(n6883), .A2(n6884), .ZN(n5006) );
  NAND2_X1 U6425 ( .A1(n9440), .A2(n5008), .ZN(n5007) );
  NAND2_X1 U6426 ( .A1(n5007), .A2(n4517), .ZN(n9545) );
  OR2_X1 U6427 ( .A1(n9723), .A2(n9442), .ZN(n5016) );
  NAND2_X1 U6428 ( .A1(n5017), .A2(n5021), .ZN(n9840) );
  NAND2_X1 U6429 ( .A1(n9991), .A2(n5019), .ZN(n5017) );
  NAND2_X1 U6430 ( .A1(n9515), .A2(n5038), .ZN(n5033) );
  OAI21_X1 U6431 ( .B1(n9515), .B2(n4473), .A(n9455), .ZN(n9502) );
  NAND3_X1 U6432 ( .A1(n6346), .A2(n5042), .A3(n5785), .ZN(n5787) );
  XNOR2_X2 U6433 ( .A(n5258), .B(n5257), .ZN(n6391) );
  NAND2_X1 U6434 ( .A1(n6277), .A2(n6276), .ZN(n6307) );
  NAND2_X1 U6435 ( .A1(n5771), .A2(n10275), .ZN(n5769) );
  NOR2_X1 U6436 ( .A1(n6214), .A2(n5778), .ZN(n5780) );
  NAND2_X1 U6437 ( .A1(n9093), .A2(n9092), .ZN(n9091) );
  INV_X1 U6438 ( .A(n6129), .ZN(n6130) );
  NAND2_X1 U6439 ( .A1(n7600), .A2(n7599), .ZN(n7602) );
  OR2_X1 U6440 ( .A1(n5243), .A2(n5961), .ZN(n5261) );
  XNOR2_X1 U6441 ( .A(n9283), .B(n4439), .ZN(n6515) );
  NOR2_X1 U6442 ( .A1(n6498), .A2(n10082), .ZN(n10069) );
  OAI211_X2 U6443 ( .C1(n7296), .C2(n6132), .A(n6131), .B(n6130), .ZN(n6285)
         );
  AOI21_X2 U6444 ( .B1(n8440), .B2(n8826), .A(n8422), .ZN(n8414) );
  OR2_X1 U6445 ( .A1(n7672), .A2(n8831), .ZN(n5044) );
  NAND2_X2 U6446 ( .A1(n6506), .A2(n10090), .ZN(n10058) );
  OR2_X1 U6447 ( .A1(n9862), .A2(n9423), .ZN(n5046) );
  OR2_X1 U6448 ( .A1(n9441), .A2(n9575), .ZN(n5048) );
  INV_X1 U6449 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n5494) );
  INV_X1 U6450 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5177) );
  OR2_X1 U6451 ( .A1(n4443), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9769) );
  AND4_X1 U6452 ( .A1(n5793), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n5049)
         );
  NAND2_X1 U6453 ( .A1(n5914), .A2(n8103), .ZN(n8481) );
  INV_X1 U6454 ( .A(n10236), .ZN(n5763) );
  OR2_X1 U6455 ( .A1(n7679), .A2(n8124), .ZN(n5050) );
  OR2_X1 U6456 ( .A1(n9707), .A2(n9451), .ZN(n5052) );
  AND2_X1 U6457 ( .A1(n5760), .A2(n5759), .ZN(n5053) );
  INV_X1 U6458 ( .A(n7919), .ZN(n5617) );
  OR2_X1 U6459 ( .A1(n7706), .A2(n8349), .ZN(n5055) );
  INV_X1 U6460 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5156) );
  INV_X1 U6461 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5162) );
  INV_X1 U6462 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5777) );
  OR2_X1 U6463 ( .A1(n7703), .A2(n8063), .ZN(n7704) );
  NAND2_X1 U6464 ( .A1(n5263), .A2(n7927), .ZN(n6446) );
  INV_X1 U6465 ( .A(n5558), .ZN(n5557) );
  NAND2_X1 U6466 ( .A1(n5582), .A2(n4479), .ZN(n5584) );
  INV_X1 U6467 ( .A(n7330), .ZN(n6091) );
  OR2_X1 U6468 ( .A1(n9031), .A2(n9030), .ZN(n9032) );
  INV_X1 U6469 ( .A(n7405), .ZN(n7261) );
  INV_X1 U6470 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U6471 ( .A1(n9856), .A2(n9427), .ZN(n9425) );
  INV_X1 U6472 ( .A(SI_22_), .ZN(n5142) );
  INV_X1 U6473 ( .A(SI_16_), .ZN(n5118) );
  INV_X1 U6474 ( .A(SI_9_), .ZN(n5089) );
  INV_X1 U6475 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5173) );
  NAND2_X2 U6476 ( .A1(n5878), .A2(n5877), .ZN(n5886) );
  OR2_X1 U6477 ( .A1(n5610), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U6478 ( .A1(n5557), .A2(n5556), .ZN(n5575) );
  INV_X1 U6479 ( .A(n5508), .ZN(n5189) );
  INV_X1 U6480 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5182) );
  INV_X1 U6481 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5172) );
  AND2_X1 U6482 ( .A1(n5679), .A2(n8096), .ZN(n5726) );
  AND2_X1 U6483 ( .A1(n8861), .A2(n7718), .ZN(n8085) );
  INV_X1 U6484 ( .A(n7369), .ZN(n7262) );
  OR2_X1 U6485 ( .A1(n6098), .A2(n9208), .ZN(n7405) );
  INV_X1 U6486 ( .A(n10092), .ZN(n7601) );
  OR3_X1 U6487 ( .A1(n7389), .A2(n9197), .A3(n9163), .ZN(n7390) );
  NAND2_X1 U6488 ( .A1(n7261), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n7407) );
  INV_X1 U6489 ( .A(n6677), .ZN(n9368) );
  INV_X1 U6490 ( .A(n6187), .ZN(n10023) );
  INV_X1 U6491 ( .A(n9424), .ZN(n9427) );
  INV_X1 U6492 ( .A(n7111), .ZN(n6886) );
  AND2_X1 U6493 ( .A1(n6519), .A2(n10124), .ZN(n6499) );
  INV_X1 U6494 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6027) );
  INV_X1 U6495 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8593) );
  INV_X1 U6496 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U6497 ( .A1(n5185), .A2(n5184), .ZN(n5470) );
  OR2_X1 U6498 ( .A1(n5713), .A2(n5873), .ZN(n5905) );
  INV_X1 U6499 ( .A(n5626), .ZN(n7670) );
  INV_X1 U6500 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U6501 ( .A1(n5595), .A2(n5594), .ZN(n5610) );
  OR2_X1 U6502 ( .A1(n5575), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U6503 ( .A1(n5189), .A2(n5188), .ZN(n5518) );
  OR2_X1 U6504 ( .A1(n5470), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6505 ( .A1(n5183), .A2(n5182), .ZN(n5459) );
  INV_X1 U6506 ( .A(n7927), .ZN(n7971) );
  OR2_X1 U6507 ( .A1(n5876), .A2(n8096), .ZN(n6367) );
  INV_X1 U6508 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5766) );
  INV_X1 U6509 ( .A(n8481), .ZN(n8463) );
  INV_X1 U6510 ( .A(n8466), .ZN(n8480) );
  OR2_X1 U6511 ( .A1(n5732), .A2(n8118), .ZN(n10236) );
  INV_X1 U6512 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9208) );
  OR2_X1 U6513 ( .A1(n6189), .A2(n7664), .ZN(n9222) );
  OR2_X1 U6514 ( .A1(n7428), .A2(n9087), .ZN(n9478) );
  NAND2_X1 U6515 ( .A1(n9450), .A2(n5052), .ZN(n9453) );
  INV_X1 U6516 ( .A(n9723), .ZN(n9575) );
  INV_X1 U6517 ( .A(n9273), .ZN(n9423) );
  INV_X1 U6518 ( .A(n9274), .ZN(n9414) );
  NAND2_X1 U6519 ( .A1(n10088), .A2(n10092), .ZN(n10012) );
  INV_X1 U6520 ( .A(n6165), .ZN(n6164) );
  AND2_X1 U6521 ( .A1(n6522), .A2(n7604), .ZN(n10072) );
  AND2_X1 U6522 ( .A1(n10088), .A2(n4555), .ZN(n9679) );
  AND2_X1 U6523 ( .A1(n5567), .A2(n5553), .ZN(n5565) );
  AND2_X1 U6524 ( .A1(n5129), .A2(n5128), .ZN(n5465) );
  INV_X1 U6525 ( .A(n7893), .ZN(n7850) );
  AND2_X1 U6526 ( .A1(n5909), .A2(n5908), .ZN(n7821) );
  AND3_X1 U6527 ( .A1(n5512), .A2(n5511), .A3(n5510), .ZN(n8393) );
  INV_X1 U6528 ( .A(n8297), .ZN(n8266) );
  INV_X1 U6529 ( .A(n5633), .ZN(n5856) );
  AND2_X1 U6530 ( .A1(P2_U3893), .A2(n5633), .ZN(n8309) );
  INV_X1 U6531 ( .A(n8444), .ZN(n10228) );
  INV_X1 U6532 ( .A(n8831), .ZN(n8843) );
  AND2_X1 U6533 ( .A1(n8026), .A2(n8027), .ZN(n8029) );
  OR2_X1 U6534 ( .A1(n6719), .A2(n5763), .ZN(n10274) );
  OR2_X1 U6535 ( .A1(n5916), .A2(n5898), .ZN(n5719) );
  AND2_X1 U6536 ( .A1(n5901), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5991) );
  INV_X1 U6537 ( .A(n8954), .ZN(n8946) );
  INV_X1 U6538 ( .A(n9268), .ZN(n9247) );
  NAND2_X1 U6539 ( .A1(n6286), .A2(n7485), .ZN(n9475) );
  OR2_X1 U6540 ( .A1(n6095), .A2(n6094), .ZN(n9435) );
  INV_X1 U6541 ( .A(n9774), .ZN(n6286) );
  INV_X1 U6542 ( .A(n9958), .ZN(n9948) );
  INV_X1 U6543 ( .A(n9930), .ZN(n9961) );
  INV_X1 U6544 ( .A(n10012), .ZN(n10081) );
  INV_X1 U6545 ( .A(n9493), .ZN(n9484) );
  INV_X1 U6546 ( .A(n9462), .ZN(n9581) );
  INV_X1 U6547 ( .A(n10072), .ZN(n10112) );
  INV_X1 U6548 ( .A(n9621), .ZN(n10077) );
  AOI21_X1 U6549 ( .B1(n6164), .B2(n6161), .A(n6160), .ZN(n9681) );
  INV_X1 U6550 ( .A(n10190), .ZN(n10150) );
  NAND2_X1 U6551 ( .A1(n9992), .A2(n10116), .ZN(n10190) );
  AOI21_X1 U6552 ( .B1(n10110), .B2(n6505), .A(n6504), .ZN(n9742) );
  AND2_X1 U6553 ( .A1(n9775), .A2(n7177), .ZN(n6162) );
  AND2_X1 U6554 ( .A1(n6348), .A2(n6347), .ZN(n9907) );
  OR2_X1 U6555 ( .A1(n5902), .A2(n7121), .ZN(n5858) );
  AND2_X1 U6556 ( .A1(n5892), .A2(n5891), .ZN(n7887) );
  AND2_X1 U6557 ( .A1(n7918), .A2(n5632), .ZN(n7953) );
  NAND2_X1 U6558 ( .A1(n5543), .A2(n5542), .ZN(n8360) );
  INV_X1 U6559 ( .A(n8309), .ZN(n7070) );
  NAND2_X1 U6560 ( .A1(n6259), .A2(n8292), .ZN(n8310) );
  NAND2_X1 U6561 ( .A1(n5734), .A2(n8482), .ZN(n8431) );
  NAND2_X2 U6562 ( .A1(n5733), .A2(n8444), .ZN(n10233) );
  NAND2_X1 U6563 ( .A1(n10233), .A2(n10222), .ZN(n8783) );
  NAND2_X1 U6564 ( .A1(n10289), .A2(n10274), .ZN(n8837) );
  NAND2_X1 U6565 ( .A1(n10289), .A2(n10244), .ZN(n8831) );
  INV_X1 U6566 ( .A(n8790), .ZN(n8852) );
  NAND2_X1 U6567 ( .A1(n10275), .A2(n10274), .ZN(n8919) );
  AND2_X1 U6568 ( .A1(n5720), .A2(n5719), .ZN(n10277) );
  INV_X1 U6569 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8945) );
  INV_X1 U6570 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7047) );
  INV_X1 U6571 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6121) );
  OR2_X1 U6572 ( .A1(n4443), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8954) );
  AND2_X1 U6573 ( .A1(n6023), .A2(n6224), .ZN(n9883) );
  AND2_X1 U6574 ( .A1(n6191), .A2(n10090), .ZN(n9258) );
  INV_X1 U6575 ( .A(n9703), .ZN(n9519) );
  NAND2_X1 U6576 ( .A1(n7438), .A2(n7437), .ZN(n9456) );
  OR2_X1 U6577 ( .A1(n7324), .A2(n7323), .ZN(n9424) );
  OR2_X1 U6578 ( .A1(n9885), .A2(n6286), .ZN(n9952) );
  OR2_X1 U6579 ( .A1(n9885), .A2(n9875), .ZN(n9958) );
  INV_X1 U6580 ( .A(n10097), .ZN(n9671) );
  NAND2_X1 U6581 ( .A1(n10058), .A2(n10028), .ZN(n9630) );
  INV_X1 U6582 ( .A(n10221), .ZN(n10219) );
  INV_X1 U6583 ( .A(n10201), .ZN(n10200) );
  INV_X1 U6584 ( .A(n10110), .ZN(n10109) );
  INV_X1 U6585 ( .A(n5999), .ZN(n7175) );
  INV_X1 U6586 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8607) );
  INV_X2 U6587 ( .A(n9284), .ZN(P1_U3973) );
  INV_X1 U6588 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5685) );
  AND2_X1 U6589 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6590 ( .A1(n7904), .A2(n5058), .ZN(n5240) );
  AND2_X1 U6591 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6592 ( .A1(n5549), .A2(n5059), .ZN(n6140) );
  NAND2_X1 U6593 ( .A1(n5240), .A2(n6140), .ZN(n5244) );
  NAND2_X1 U6594 ( .A1(n5061), .A2(SI_1_), .ZN(n5062) );
  INV_X1 U6595 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5961) );
  INV_X1 U6596 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6308) );
  INV_X1 U6597 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U6598 ( .A1(n5064), .A2(SI_2_), .ZN(n5065) );
  MUX2_X1 U6599 ( .A(n5962), .B(n6415), .S(n5963), .Z(n5066) );
  INV_X1 U6600 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6601 ( .A1(n5067), .A2(SI_3_), .ZN(n5068) );
  MUX2_X1 U6602 ( .A(n5971), .B(n6464), .S(n5963), .Z(n5069) );
  NAND2_X1 U6603 ( .A1(n5287), .A2(n5286), .ZN(n5072) );
  INV_X1 U6604 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6605 ( .A1(n5070), .A2(SI_4_), .ZN(n5071) );
  MUX2_X1 U6606 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5963), .Z(n5074) );
  XNOR2_X1 U6607 ( .A(n5074), .B(n5073), .ZN(n5298) );
  NAND2_X1 U6608 ( .A1(n5074), .A2(SI_5_), .ZN(n5075) );
  MUX2_X1 U6609 ( .A(n5986), .B(n6689), .S(n5549), .Z(n5076) );
  XNOR2_X1 U6610 ( .A(n5076), .B(SI_6_), .ZN(n5321) );
  INV_X1 U6611 ( .A(n5076), .ZN(n5077) );
  MUX2_X1 U6612 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5549), .Z(n5079) );
  INV_X1 U6613 ( .A(SI_7_), .ZN(n5078) );
  NAND2_X1 U6614 ( .A1(n5336), .A2(n5335), .ZN(n5081) );
  NAND2_X1 U6615 ( .A1(n5079), .A2(SI_7_), .ZN(n5080) );
  MUX2_X1 U6616 ( .A(n5352), .B(n5082), .S(n5549), .Z(n5084) );
  INV_X1 U6617 ( .A(SI_8_), .ZN(n5083) );
  NAND2_X1 U6618 ( .A1(n5084), .A2(n5083), .ZN(n5087) );
  INV_X1 U6619 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6620 ( .A1(n5085), .A2(SI_8_), .ZN(n5086) );
  NAND2_X1 U6621 ( .A1(n5087), .A2(n5086), .ZN(n5350) );
  INV_X1 U6622 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5088) );
  MUX2_X1 U6623 ( .A(n6119), .B(n5088), .S(n5963), .Z(n5090) );
  NAND2_X1 U6624 ( .A1(n5090), .A2(n5089), .ZN(n5093) );
  INV_X1 U6625 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U6626 ( .A1(n5091), .A2(SI_9_), .ZN(n5092) );
  MUX2_X1 U6627 ( .A(n6121), .B(n8607), .S(n5963), .Z(n5095) );
  XNOR2_X1 U6628 ( .A(n5095), .B(SI_10_), .ZN(n5373) );
  INV_X1 U6629 ( .A(n5373), .ZN(n5094) );
  INV_X1 U6630 ( .A(n5095), .ZN(n5096) );
  NAND2_X1 U6631 ( .A1(n5096), .A2(SI_10_), .ZN(n5097) );
  MUX2_X1 U6632 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5963), .Z(n5387) );
  AND2_X1 U6633 ( .A1(n5387), .A2(SI_11_), .ZN(n5098) );
  MUX2_X1 U6634 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5549), .Z(n5099) );
  NAND2_X1 U6635 ( .A1(n5099), .A2(SI_12_), .ZN(n5103) );
  INV_X1 U6636 ( .A(n5099), .ZN(n5101) );
  INV_X1 U6637 ( .A(SI_12_), .ZN(n5100) );
  NAND2_X1 U6638 ( .A1(n5101), .A2(n5100), .ZN(n5102) );
  NAND2_X1 U6639 ( .A1(n5103), .A2(n5102), .ZN(n5401) );
  MUX2_X1 U6640 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5549), .Z(n5104) );
  NAND2_X1 U6641 ( .A1(n5104), .A2(SI_13_), .ZN(n5109) );
  INV_X1 U6642 ( .A(n5104), .ZN(n5106) );
  INV_X1 U6643 ( .A(SI_13_), .ZN(n5105) );
  NAND2_X1 U6644 ( .A1(n5106), .A2(n5105), .ZN(n5107) );
  NAND2_X1 U6645 ( .A1(n5109), .A2(n5107), .ZN(n5417) );
  INV_X1 U6646 ( .A(n5417), .ZN(n5108) );
  MUX2_X1 U6647 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4443), .Z(n5110) );
  NAND2_X1 U6648 ( .A1(n5110), .A2(SI_14_), .ZN(n5113) );
  INV_X1 U6649 ( .A(n5110), .ZN(n5111) );
  NAND2_X1 U6650 ( .A1(n5111), .A2(n8606), .ZN(n5112) );
  MUX2_X1 U6651 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4443), .Z(n5449) );
  INV_X1 U6652 ( .A(n5449), .ZN(n5115) );
  NAND2_X1 U6653 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  NAND2_X1 U6654 ( .A1(n5449), .A2(SI_15_), .ZN(n5117) );
  MUX2_X1 U6655 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4443), .Z(n5225) );
  INV_X1 U6656 ( .A(n5225), .ZN(n5119) );
  NAND2_X1 U6657 ( .A1(n5119), .A2(n5118), .ZN(n5120) );
  MUX2_X1 U6658 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4443), .Z(n5121) );
  XNOR2_X1 U6659 ( .A(n5121), .B(n8629), .ZN(n5211) );
  NAND2_X1 U6660 ( .A1(n5212), .A2(n5211), .ZN(n5124) );
  INV_X1 U6661 ( .A(n5121), .ZN(n5122) );
  NAND2_X1 U6662 ( .A1(n5122), .A2(n8629), .ZN(n5123) );
  MUX2_X1 U6663 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4443), .Z(n5125) );
  NAND2_X1 U6664 ( .A1(n5125), .A2(SI_18_), .ZN(n5129) );
  INV_X1 U6665 ( .A(n5125), .ZN(n5127) );
  INV_X1 U6666 ( .A(SI_18_), .ZN(n5126) );
  NAND2_X1 U6667 ( .A1(n5127), .A2(n5126), .ZN(n5128) );
  MUX2_X1 U6668 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4443), .Z(n5130) );
  XNOR2_X1 U6669 ( .A(n5130), .B(SI_19_), .ZN(n5477) );
  INV_X1 U6670 ( .A(n5130), .ZN(n5131) );
  INV_X1 U6671 ( .A(SI_19_), .ZN(n8746) );
  NAND2_X1 U6672 ( .A1(n5131), .A2(n8746), .ZN(n5132) );
  MUX2_X1 U6673 ( .A(n5494), .B(n7416), .S(n4443), .Z(n5134) );
  NAND2_X1 U6674 ( .A1(n5493), .A2(n5492), .ZN(n5136) );
  INV_X1 U6675 ( .A(SI_20_), .ZN(n5133) );
  NAND2_X1 U6676 ( .A1(n5134), .A2(n5133), .ZN(n5135) );
  INV_X1 U6677 ( .A(n5505), .ZN(n5139) );
  MUX2_X1 U6678 ( .A(n6968), .B(n7402), .S(n4443), .Z(n5503) );
  INV_X1 U6679 ( .A(SI_21_), .ZN(n5137) );
  NAND2_X1 U6680 ( .A1(n5503), .A2(n5137), .ZN(n5138) );
  INV_X1 U6681 ( .A(n5503), .ZN(n5140) );
  NAND2_X1 U6682 ( .A1(n5140), .A2(SI_21_), .ZN(n5141) );
  INV_X1 U6683 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7365) );
  MUX2_X1 U6684 ( .A(n7047), .B(n7365), .S(n4443), .Z(n5143) );
  NAND2_X1 U6685 ( .A1(n5143), .A2(n5142), .ZN(n5146) );
  INV_X1 U6686 ( .A(n5143), .ZN(n5144) );
  NAND2_X1 U6687 ( .A1(n5144), .A2(SI_22_), .ZN(n5145) );
  NAND2_X1 U6688 ( .A1(n5146), .A2(n5145), .ZN(n5514) );
  INV_X1 U6689 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7355) );
  MUX2_X1 U6690 ( .A(n8573), .B(n7355), .S(n4443), .Z(n5148) );
  INV_X1 U6691 ( .A(SI_23_), .ZN(n5147) );
  NAND2_X1 U6692 ( .A1(n5148), .A2(n5147), .ZN(n5528) );
  INV_X1 U6693 ( .A(n5148), .ZN(n5149) );
  NAND2_X1 U6694 ( .A1(n5149), .A2(SI_23_), .ZN(n5150) );
  NOR2_X1 U6695 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5153) );
  NOR2_X1 U6696 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5155) );
  NAND4_X1 U6697 ( .A1(n5155), .A2(n5479), .A3(n5438), .A4(n8636), .ZN(n5158)
         );
  NAND4_X1 U6698 ( .A1(n5156), .A2(n5213), .A3(n5214), .A4(n5482), .ZN(n5157)
         );
  NAND2_X1 U6699 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n5164) );
  AOI22_X1 U6700 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n5405), .B1(n5164), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6701 ( .A1(n7354), .A2(n7900), .ZN(n5171) );
  OR2_X1 U6702 ( .A1(n5746), .A2(n8573), .ZN(n5170) );
  NAND2_X1 U6703 ( .A1(n5265), .A2(n5172), .ZN(n5292) );
  INV_X1 U6704 ( .A(n5292), .ZN(n5174) );
  NAND2_X1 U6705 ( .A1(n5174), .A2(n5173), .ZN(n5309) );
  INV_X1 U6706 ( .A(n5457), .ZN(n5183) );
  OR2_X2 U6707 ( .A1(n5459), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5220) );
  INV_X1 U6708 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5184) );
  INV_X1 U6709 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5186) );
  INV_X1 U6710 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5188) );
  OR2_X2 U6711 ( .A1(n5518), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U6712 ( .A1(n5520), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6713 ( .A1(n5537), .A2(n5190), .ZN(n8363) );
  XNOR2_X2 U6714 ( .A(n5195), .B(n5194), .ZN(n7678) );
  OAI21_X1 U6715 ( .B1(n5196), .B2(n5405), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n5198) );
  INV_X1 U6716 ( .A(n5235), .ZN(n5266) );
  NAND2_X1 U6717 ( .A1(n8363), .A2(n5266), .ZN(n5205) );
  INV_X1 U6718 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8877) );
  INV_X2 U6719 ( .A(n5249), .ZN(n7911) );
  NAND2_X1 U6720 ( .A1(n7911), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U6721 ( .A1(n7912), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5201) );
  OAI211_X1 U6722 ( .C1(n5756), .C2(n8877), .A(n5202), .B(n5201), .ZN(n5203)
         );
  INV_X1 U6723 ( .A(n5203), .ZN(n5204) );
  NAND2_X1 U6724 ( .A1(n7912), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6725 ( .A1(n5456), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6726 ( .A1(n5220), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5206) );
  NAND2_X1 U6727 ( .A1(n5470), .A2(n5206), .ZN(n8429) );
  NAND2_X1 U6728 ( .A1(n5343), .A2(n8429), .ZN(n5208) );
  INV_X1 U6729 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8249) );
  OR2_X1 U6730 ( .A1(n5249), .A2(n8249), .ZN(n5207) );
  XNOR2_X1 U6731 ( .A(n5212), .B(n5211), .ZN(n7314) );
  NAND2_X1 U6732 ( .A1(n7314), .A2(n7900), .ZN(n5218) );
  AND4_X1 U6733 ( .A1(n5419), .A2(n5438), .A3(n8636), .A4(n5214), .ZN(n5215)
         );
  NAND2_X1 U6734 ( .A1(n5467), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5216) );
  XNOR2_X1 U6735 ( .A(n5216), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8273) );
  AOI22_X1 U6736 ( .A1(n5484), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5800), .B2(
        n8273), .ZN(n5217) );
  NAND2_X1 U6737 ( .A1(n7912), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6738 ( .A1(n5456), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6739 ( .A1(n5459), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6740 ( .A1(n5220), .A2(n5219), .ZN(n7818) );
  NAND2_X1 U6741 ( .A1(n5343), .A2(n7818), .ZN(n5222) );
  NAND2_X1 U6742 ( .A1(n7911), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5221) );
  INV_X1 U6743 ( .A(n8423), .ZN(n8452) );
  XNOR2_X1 U6744 ( .A(n5225), .B(SI_16_), .ZN(n5226) );
  NAND2_X1 U6745 ( .A1(n7303), .A2(n7900), .ZN(n5232) );
  NAND2_X1 U6746 ( .A1(n5228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5229) );
  MUX2_X1 U6747 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5229), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5230) );
  AOI22_X1 U6748 ( .A1(n5484), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5800), .B2(
        n8222), .ZN(n5231) );
  NAND2_X1 U6749 ( .A1(n5456), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5233) );
  INV_X1 U6750 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6751 ( .A1(n5264), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5236) );
  INV_X1 U6752 ( .A(n6581), .ZN(n8136) );
  INV_X1 U6753 ( .A(SI_0_), .ZN(n5238) );
  INV_X1 U6754 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5237) );
  OAI21_X1 U6755 ( .B1(n4443), .B2(n5238), .A(n5237), .ZN(n5239) );
  AND2_X1 U6756 ( .A1(n5240), .A2(n5239), .ZN(n8955) );
  MUX2_X1 U6757 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8955), .S(n5247), .Z(n6298) );
  NAND2_X1 U6758 ( .A1(n8136), .A2(n6298), .ZN(n6580) );
  XNOR2_X1 U6759 ( .A(n5245), .B(n5244), .ZN(n5972) );
  INV_X1 U6760 ( .A(n6586), .ZN(n10235) );
  NAND2_X1 U6761 ( .A1(n7964), .A2(n5687), .ZN(n5686) );
  NAND2_X1 U6762 ( .A1(n6580), .A2(n5686), .ZN(n6529) );
  NAND2_X1 U6763 ( .A1(n6532), .A2(n10235), .ZN(n6530) );
  NAND2_X1 U6764 ( .A1(n6529), .A2(n6530), .ZN(n5263) );
  NAND2_X1 U6765 ( .A1(n5456), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6766 ( .A1(n5266), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6767 ( .A1(n5264), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5250) );
  XNOR2_X1 U6768 ( .A(n5255), .B(n5254), .ZN(n6309) );
  OR2_X1 U6769 ( .A1(n5246), .A2(n6309), .ZN(n5260) );
  OR2_X1 U6770 ( .A1(n5247), .A2(n6391), .ZN(n5259) );
  NAND2_X1 U6771 ( .A1(n8134), .A2(n6537), .ZN(n6447) );
  OR2_X1 U6772 ( .A1(n8134), .A2(n6537), .ZN(n5262) );
  AND2_X1 U6773 ( .A1(n6447), .A2(n5262), .ZN(n7927) );
  NAND2_X1 U6774 ( .A1(n6446), .A2(n6447), .ZN(n5277) );
  NAND2_X1 U6775 ( .A1(n5264), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6776 ( .A1(n5456), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6777 ( .A1(n5266), .A2(n5265), .ZN(n5268) );
  NAND2_X1 U6778 ( .A1(n4442), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6779 ( .A1(n5284), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5272) );
  INV_X1 U6780 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5271) );
  XNOR2_X1 U6781 ( .A(n5274), .B(n5273), .ZN(n6414) );
  OR2_X1 U6782 ( .A1(n5246), .A2(n6414), .ZN(n5276) );
  OR2_X1 U6783 ( .A1(n5243), .A2(n5962), .ZN(n5275) );
  OAI211_X1 U6784 ( .C1(n5247), .C2(n6400), .A(n5276), .B(n5275), .ZN(n10245)
         );
  NAND2_X1 U6785 ( .A1(n6591), .A2(n10245), .ZN(n7982) );
  INV_X1 U6786 ( .A(n6591), .ZN(n8133) );
  INV_X1 U6787 ( .A(n10245), .ZN(n6452) );
  NAND2_X1 U6788 ( .A1(n8133), .A2(n6452), .ZN(n7997) );
  NAND2_X1 U6789 ( .A1(n7982), .A2(n7997), .ZN(n7926) );
  NAND2_X1 U6790 ( .A1(n5277), .A2(n7926), .ZN(n6445) );
  NAND2_X1 U6791 ( .A1(n6591), .A2(n6452), .ZN(n5278) );
  NAND2_X1 U6792 ( .A1(n7912), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6793 ( .A1(n5456), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6794 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5279) );
  NAND2_X1 U6795 ( .A1(n5292), .A2(n5279), .ZN(n6599) );
  NAND2_X1 U6796 ( .A1(n5343), .A2(n6599), .ZN(n5281) );
  NAND2_X1 U6797 ( .A1(n7911), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5280) );
  NAND4_X1 U6798 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n8132)
         );
  OR2_X1 U6799 ( .A1(n5284), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6800 ( .A1(n5300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5285) );
  XNOR2_X1 U6801 ( .A(n5285), .B(n5301), .ZN(n5970) );
  XNOR2_X1 U6802 ( .A(n5287), .B(n5286), .ZN(n6465) );
  OR2_X1 U6803 ( .A1(n5246), .A2(n6465), .ZN(n5289) );
  OR2_X1 U6804 ( .A1(n5746), .A2(n5971), .ZN(n5288) );
  OAI211_X1 U6805 ( .C1(n7905), .C2(n5970), .A(n5289), .B(n5288), .ZN(n6602)
         );
  NOR2_X1 U6806 ( .A1(n8132), .A2(n6602), .ZN(n5291) );
  NAND2_X1 U6807 ( .A1(n8132), .A2(n6602), .ZN(n5290) );
  NAND2_X1 U6808 ( .A1(n7912), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6809 ( .A1(n5456), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6810 ( .A1(n5292), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6811 ( .A1(n5309), .A2(n5293), .ZN(n6770) );
  NAND2_X1 U6812 ( .A1(n5343), .A2(n6770), .ZN(n5295) );
  NAND2_X1 U6813 ( .A1(n7911), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5294) );
  XNOR2_X1 U6814 ( .A(n5299), .B(n5298), .ZN(n6610) );
  OR2_X1 U6815 ( .A1(n5246), .A2(n6610), .ZN(n5306) );
  INV_X1 U6816 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5977) );
  OR2_X1 U6817 ( .A1(n5746), .A2(n5977), .ZN(n5305) );
  INV_X1 U6818 ( .A(n5300), .ZN(n5302) );
  NAND2_X1 U6819 ( .A1(n5302), .A2(n5301), .ZN(n5315) );
  NAND2_X1 U6820 ( .A1(n5315), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5303) );
  XNOR2_X1 U6821 ( .A(n5303), .B(n5316), .ZN(n6754) );
  OR2_X1 U6822 ( .A1(n7905), .A2(n6754), .ZN(n5304) );
  NAND2_X1 U6823 ( .A1(n6829), .A2(n10256), .ZN(n5307) );
  INV_X1 U6824 ( .A(n10256), .ZN(n6722) );
  NAND2_X1 U6825 ( .A1(n8131), .A2(n6722), .ZN(n5308) );
  NAND2_X1 U6826 ( .A1(n7912), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6827 ( .A1(n5456), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6828 ( .A1(n5309), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6829 ( .A1(n5327), .A2(n5310), .ZN(n6837) );
  NAND2_X1 U6830 ( .A1(n5343), .A2(n6837), .ZN(n5312) );
  NAND2_X1 U6831 ( .A1(n7911), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5311) );
  NAND4_X1 U6832 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n8130)
         );
  INV_X1 U6833 ( .A(n5315), .ZN(n5317) );
  NAND2_X1 U6834 ( .A1(n5317), .A2(n5316), .ZN(n5319) );
  NAND2_X1 U6835 ( .A1(n5319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5318) );
  MUX2_X1 U6836 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5318), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5320) );
  NAND2_X1 U6837 ( .A1(n5320), .A2(n5348), .ZN(n6807) );
  XNOR2_X1 U6838 ( .A(n5322), .B(n5321), .ZN(n6688) );
  OR2_X1 U6839 ( .A1(n5246), .A2(n6688), .ZN(n5324) );
  OR2_X1 U6840 ( .A1(n5746), .A2(n5986), .ZN(n5323) );
  OAI211_X1 U6841 ( .C1(n7905), .C2(n6807), .A(n5324), .B(n5323), .ZN(n6840)
         );
  AND2_X1 U6842 ( .A1(n8130), .A2(n6840), .ZN(n5326) );
  INV_X1 U6843 ( .A(n8130), .ZN(n6894) );
  INV_X1 U6844 ( .A(n6840), .ZN(n10262) );
  NAND2_X1 U6845 ( .A1(n6894), .A2(n10262), .ZN(n5325) );
  NAND2_X1 U6846 ( .A1(n7912), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6847 ( .A1(n5456), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6848 ( .A1(n5327), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6849 ( .A1(n5341), .A2(n5328), .ZN(n6895) );
  NAND2_X1 U6850 ( .A1(n5343), .A2(n6895), .ZN(n5330) );
  NAND2_X1 U6851 ( .A1(n7911), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6852 ( .A1(n5348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5334) );
  INV_X1 U6853 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5333) );
  XNOR2_X1 U6854 ( .A(n5334), .B(n5333), .ZN(n6004) );
  XNOR2_X1 U6855 ( .A(n5336), .B(n5335), .ZN(n6785) );
  OR2_X1 U6856 ( .A1(n5246), .A2(n6785), .ZN(n5338) );
  INV_X1 U6857 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6005) );
  OR2_X1 U6858 ( .A1(n5746), .A2(n6005), .ZN(n5337) );
  OAI211_X1 U6859 ( .C1(n7905), .C2(n6004), .A(n5338), .B(n5337), .ZN(n6948)
         );
  NAND2_X1 U6860 ( .A1(n7084), .A2(n6948), .ZN(n7956) );
  INV_X1 U6861 ( .A(n6948), .ZN(n6960) );
  NAND2_X1 U6862 ( .A1(n8129), .A2(n6960), .ZN(n6961) );
  NAND2_X1 U6863 ( .A1(n7956), .A2(n6961), .ZN(n7989) );
  NAND2_X1 U6864 ( .A1(n7084), .A2(n6960), .ZN(n5339) );
  NAND2_X1 U6865 ( .A1(n7912), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6866 ( .A1(n5456), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6867 ( .A1(n5341), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6868 ( .A1(n5357), .A2(n5342), .ZN(n7089) );
  NAND2_X1 U6869 ( .A1(n5343), .A2(n7089), .ZN(n5345) );
  NAND2_X1 U6870 ( .A1(n7911), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5344) );
  NAND4_X1 U6871 ( .A1(n5347), .A2(n5346), .A3(n5345), .A4(n5344), .ZN(n8128)
         );
  NAND2_X1 U6872 ( .A1(n5349), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5366) );
  INV_X1 U6873 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5365) );
  XNOR2_X1 U6874 ( .A(n5351), .B(n5350), .ZN(n6862) );
  NAND2_X1 U6875 ( .A1(n6862), .A2(n7900), .ZN(n5354) );
  OR2_X1 U6876 ( .A1(n5746), .A2(n5352), .ZN(n5353) );
  NOR2_X1 U6877 ( .A1(n8128), .A2(n7086), .ZN(n5355) );
  NAND2_X1 U6878 ( .A1(n8128), .A2(n7086), .ZN(n5356) );
  NAND2_X1 U6879 ( .A1(n7912), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6880 ( .A1(n7913), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6881 ( .A1(n5357), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6882 ( .A1(n5378), .A2(n5358), .ZN(n10229) );
  NAND2_X1 U6883 ( .A1(n5343), .A2(n10229), .ZN(n5360) );
  NAND2_X1 U6884 ( .A1(n7911), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6885 ( .A1(n6848), .A2(n7900), .ZN(n5370) );
  NAND2_X1 U6886 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  NAND2_X1 U6887 ( .A1(n5367), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5368) );
  XNOR2_X1 U6888 ( .A(n5368), .B(P2_IR_REG_9__SCAN_IN), .ZN(n5850) );
  AOI22_X1 U6889 ( .A1(n5484), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5800), .B2(
        n5850), .ZN(n5369) );
  NAND2_X1 U6890 ( .A1(n7051), .A2(n7182), .ZN(n5371) );
  XNOR2_X1 U6891 ( .A(n5372), .B(n5373), .ZN(n6868) );
  NAND2_X1 U6892 ( .A1(n6868), .A2(n7900), .ZN(n5377) );
  NAND2_X1 U6893 ( .A1(n5374), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5375) );
  XNOR2_X1 U6894 ( .A(n5375), .B(P2_IR_REG_10__SCAN_IN), .ZN(n5864) );
  AOI22_X1 U6895 ( .A1(n5484), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5800), .B2(
        n5864), .ZN(n5376) );
  NAND2_X1 U6896 ( .A1(n5377), .A2(n5376), .ZN(n7765) );
  NAND2_X1 U6897 ( .A1(n7912), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6898 ( .A1(n5456), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6899 ( .A1(n5378), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6900 ( .A1(n5394), .A2(n5379), .ZN(n7754) );
  NAND2_X1 U6901 ( .A1(n5343), .A2(n7754), .ZN(n5381) );
  NAND2_X1 U6902 ( .A1(n7911), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5380) );
  NAND4_X1 U6903 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n8126)
         );
  OR2_X1 U6904 ( .A1(n7765), .A2(n8126), .ZN(n5384) );
  NAND2_X1 U6905 ( .A1(n7049), .A2(n5384), .ZN(n5386) );
  NAND2_X1 U6906 ( .A1(n7765), .A2(n8126), .ZN(n5385) );
  XNOR2_X1 U6907 ( .A(n5387), .B(SI_11_), .ZN(n5388) );
  XNOR2_X1 U6908 ( .A(n5389), .B(n5388), .ZN(n7005) );
  NAND2_X1 U6909 ( .A1(n7005), .A2(n7900), .ZN(n5393) );
  NOR2_X1 U6910 ( .A1(n4450), .A2(n5405), .ZN(n5390) );
  MUX2_X1 U6911 ( .A(n5405), .B(n5390), .S(P2_IR_REG_11__SCAN_IN), .Z(n5391)
         );
  NOR2_X1 U6912 ( .A1(n5391), .A2(n5420), .ZN(n7167) );
  AOI22_X1 U6913 ( .A1(n5484), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5800), .B2(
        n7167), .ZN(n5392) );
  NAND2_X1 U6914 ( .A1(n7912), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6915 ( .A1(n7913), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6916 ( .A1(n5394), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6917 ( .A1(n5409), .A2(n5395), .ZN(n8778) );
  NAND2_X1 U6918 ( .A1(n5343), .A2(n8778), .ZN(n5397) );
  NAND2_X1 U6919 ( .A1(n7911), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5396) );
  AND2_X1 U6920 ( .A1(n4556), .A2(n8125), .ZN(n5400) );
  NAND2_X1 U6921 ( .A1(n5402), .A2(n5401), .ZN(n5404) );
  NAND2_X1 U6922 ( .A1(n6992), .A2(n7900), .ZN(n5408) );
  OR2_X1 U6923 ( .A1(n5420), .A2(n5405), .ZN(n5406) );
  XNOR2_X1 U6924 ( .A(n5406), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8149) );
  AOI22_X1 U6925 ( .A1(n5484), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5800), .B2(
        n8149), .ZN(n5407) );
  NAND2_X1 U6926 ( .A1(n7912), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6927 ( .A1(n7913), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6928 ( .A1(n5409), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6929 ( .A1(n5424), .A2(n5410), .ZN(n7803) );
  NAND2_X1 U6930 ( .A1(n5343), .A2(n7803), .ZN(n5412) );
  NAND2_X1 U6931 ( .A1(n7911), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5411) );
  NAND4_X1 U6932 ( .A1(n5414), .A2(n5413), .A3(n5412), .A4(n5411), .ZN(n8124)
         );
  NAND2_X1 U6933 ( .A1(n7679), .A2(n8124), .ZN(n5415) );
  NAND2_X1 U6934 ( .A1(n7273), .A2(n7900), .ZN(n5423) );
  NAND2_X1 U6935 ( .A1(n5420), .A2(n5419), .ZN(n5421) );
  NAND2_X1 U6936 ( .A1(n5421), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5436) );
  XNOR2_X1 U6937 ( .A(n5436), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8174) );
  AOI22_X1 U6938 ( .A1(n5484), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5800), .B2(
        n8174), .ZN(n5422) );
  NAND2_X1 U6939 ( .A1(n7913), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6940 ( .A1(n7912), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6941 ( .A1(n5424), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6942 ( .A1(n5443), .A2(n5425), .ZN(n8483) );
  NAND2_X1 U6943 ( .A1(n5343), .A2(n8483), .ZN(n5427) );
  NAND2_X1 U6944 ( .A1(n7911), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5426) );
  AND2_X1 U6945 ( .A1(n8929), .A2(n8465), .ZN(n5431) );
  OAI21_X2 U6946 ( .B1(n8476), .B2(n5431), .A(n5430), .ZN(n8460) );
  OR2_X1 U6947 ( .A1(n5433), .A2(n5432), .ZN(n5435) );
  AND2_X1 U6948 ( .A1(n5434), .A2(n5435), .ZN(n7279) );
  NAND2_X1 U6949 ( .A1(n7279), .A2(n7900), .ZN(n5442) );
  NAND2_X1 U6950 ( .A1(n5436), .A2(n8636), .ZN(n5437) );
  NAND2_X1 U6951 ( .A1(n5437), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6952 ( .A1(n5439), .A2(n5438), .ZN(n5452) );
  OR2_X1 U6953 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  AND2_X1 U6954 ( .A1(n5452), .A2(n5440), .ZN(n8177) );
  AOI22_X1 U6955 ( .A1(n5484), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5800), .B2(
        n8177), .ZN(n5441) );
  NAND2_X1 U6956 ( .A1(n7912), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U6957 ( .A1(n7913), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6958 ( .A1(n5443), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6959 ( .A1(n5457), .A2(n5444), .ZN(n8471) );
  NAND2_X1 U6960 ( .A1(n5343), .A2(n8471), .ZN(n5446) );
  NAND2_X1 U6961 ( .A1(n7911), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5445) );
  NAND4_X1 U6962 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(n8451)
         );
  XNOR2_X1 U6963 ( .A(n5449), .B(SI_15_), .ZN(n5450) );
  NAND2_X1 U6964 ( .A1(n7288), .A2(n7900), .ZN(n5455) );
  NAND2_X1 U6965 ( .A1(n5452), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5453) );
  XNOR2_X1 U6966 ( .A(n5453), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8218) );
  AOI22_X1 U6967 ( .A1(n5484), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5800), .B2(
        n8218), .ZN(n5454) );
  NAND2_X1 U6968 ( .A1(n5456), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6969 ( .A1(n7912), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6970 ( .A1(n5457), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6971 ( .A1(n5459), .A2(n5458), .ZN(n8455) );
  NAND2_X1 U6972 ( .A1(n5343), .A2(n8455), .ZN(n5461) );
  NAND2_X1 U6973 ( .A1(n7911), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5460) );
  NAND4_X1 U6974 ( .A1(n5463), .A2(n5462), .A3(n5461), .A4(n5460), .ZN(n8464)
         );
  NAND2_X1 U6975 ( .A1(n8916), .A2(n8464), .ZN(n5464) );
  NAND2_X1 U6976 ( .A1(n8830), .A2(n8423), .ZN(n5696) );
  NAND2_X1 U6977 ( .A1(n8044), .A2(n5696), .ZN(n8436) );
  OR2_X1 U6978 ( .A1(n8826), .A2(n7826), .ZN(n8042) );
  NAND2_X1 U6979 ( .A1(n8826), .A2(n7826), .ZN(n8411) );
  NOR2_X1 U6980 ( .A1(n8421), .A2(n8428), .ZN(n8422) );
  NAND2_X1 U6981 ( .A1(n7325), .A2(n7900), .ZN(n5469) );
  XNOR2_X1 U6982 ( .A(n5480), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8287) );
  AOI22_X1 U6983 ( .A1(n5484), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5800), .B2(
        n8287), .ZN(n5468) );
  NAND2_X1 U6984 ( .A1(n7913), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U6985 ( .A1(n7912), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6986 ( .A1(n5470), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6987 ( .A1(n5486), .A2(n5471), .ZN(n8418) );
  NAND2_X1 U6988 ( .A1(n5343), .A2(n8418), .ZN(n5473) );
  NAND2_X1 U6989 ( .A1(n7911), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5472) );
  NAND4_X1 U6990 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n8405)
         );
  NOR2_X1 U6991 ( .A1(n8903), .A2(n8405), .ZN(n5476) );
  INV_X1 U6992 ( .A(n8903), .ZN(n7877) );
  NAND2_X1 U6993 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  NAND2_X1 U6994 ( .A1(n5481), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5483) );
  AOI22_X1 U6995 ( .A1(n5484), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8296), .B2(
        n5800), .ZN(n5485) );
  NAND2_X1 U6996 ( .A1(n7913), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6997 ( .A1(n7911), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U6998 ( .A1(n5486), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6999 ( .A1(n5497), .A2(n5487), .ZN(n7770) );
  NAND2_X1 U7000 ( .A1(n5343), .A2(n7770), .ZN(n5489) );
  NAND2_X1 U7001 ( .A1(n7912), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7002 ( .A1(n8819), .A2(n8394), .ZN(n8051) );
  NAND2_X1 U7003 ( .A1(n8047), .A2(n8051), .ZN(n8402) );
  NAND2_X1 U7004 ( .A1(n7415), .A2(n7900), .ZN(n5496) );
  OR2_X1 U7005 ( .A1(n5746), .A2(n5494), .ZN(n5495) );
  NAND2_X1 U7006 ( .A1(n5497), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7007 ( .A1(n5508), .A2(n5498), .ZN(n8395) );
  NAND2_X1 U7008 ( .A1(n8395), .A2(n5343), .ZN(n5502) );
  NAND2_X1 U7009 ( .A1(n7913), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7010 ( .A1(n7912), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7011 ( .A1(n7911), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7012 ( .A1(n8896), .A2(n7791), .ZN(n8377) );
  NAND2_X1 U7013 ( .A1(n8055), .A2(n8377), .ZN(n8391) );
  NOR2_X1 U7014 ( .A1(n8896), .A2(n8404), .ZN(n8382) );
  XNOR2_X1 U7015 ( .A(n5503), .B(SI_21_), .ZN(n5504) );
  XNOR2_X1 U7016 ( .A(n5505), .B(n5504), .ZN(n7401) );
  NAND2_X1 U7017 ( .A1(n7401), .A2(n7900), .ZN(n5507) );
  OR2_X1 U7018 ( .A1(n5746), .A2(n6968), .ZN(n5506) );
  NAND2_X1 U7019 ( .A1(n5508), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7020 ( .A1(n5518), .A2(n5509), .ZN(n8388) );
  NAND2_X1 U7021 ( .A1(n8388), .A2(n5343), .ZN(n5512) );
  AOI22_X1 U7022 ( .A1(n7912), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5456), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7023 ( .A1(n4442), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7024 ( .A1(n8890), .A2(n8393), .ZN(n8060) );
  NAND2_X1 U7025 ( .A1(n8061), .A2(n8060), .ZN(n8381) );
  NAND2_X1 U7026 ( .A1(n8384), .A2(n5513), .ZN(n8369) );
  XNOR2_X1 U7027 ( .A(n5515), .B(n5514), .ZN(n7364) );
  NAND2_X1 U7028 ( .A1(n7364), .A2(n7900), .ZN(n5517) );
  OR2_X1 U7029 ( .A1(n5746), .A2(n7047), .ZN(n5516) );
  INV_X1 U7030 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U7031 ( .A1(n5518), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7032 ( .A1(n5520), .A2(n5519), .ZN(n8374) );
  NAND2_X1 U7033 ( .A1(n8374), .A2(n5266), .ZN(n5522) );
  AOI22_X1 U7034 ( .A1(n7912), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n5456), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7035 ( .A1(n8884), .A2(n8385), .ZN(n5523) );
  NAND2_X1 U7036 ( .A1(n8368), .A2(n5524), .ZN(n8359) );
  NAND2_X1 U7037 ( .A1(n8359), .A2(n5055), .ZN(n5525) );
  NAND2_X1 U7038 ( .A1(n5527), .A2(n5526), .ZN(n5529) );
  INV_X1 U7039 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7676) );
  INV_X1 U7040 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7343) );
  MUX2_X1 U7041 ( .A(n7676), .B(n7343), .S(n4443), .Z(n5530) );
  INV_X1 U7042 ( .A(SI_24_), .ZN(n8589) );
  NAND2_X1 U7043 ( .A1(n5530), .A2(n8589), .ZN(n5547) );
  INV_X1 U7044 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7045 ( .A1(n5531), .A2(SI_24_), .ZN(n5532) );
  XNOR2_X1 U7046 ( .A(n5546), .B(n5545), .ZN(n7342) );
  NAND2_X1 U7047 ( .A1(n7342), .A2(n7900), .ZN(n5534) );
  OR2_X1 U7048 ( .A1(n5746), .A2(n7676), .ZN(n5533) );
  INV_X1 U7049 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7050 ( .A1(n5537), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7051 ( .A1(n5558), .A2(n5538), .ZN(n8351) );
  NAND2_X1 U7052 ( .A1(n8351), .A2(n5343), .ZN(n5543) );
  INV_X1 U7053 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U7054 ( .A1(n7913), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U7055 ( .A1(n7912), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5539) );
  OAI211_X1 U7056 ( .C1(n8693), .C2(n5249), .A(n5540), .B(n5539), .ZN(n5541)
         );
  INV_X1 U7057 ( .A(n5541), .ZN(n5542) );
  NOR2_X1 U7058 ( .A1(n7839), .A2(n8360), .ZN(n5544) );
  NAND2_X1 U7059 ( .A1(n5546), .A2(n5545), .ZN(n5548) );
  INV_X1 U7060 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7176) );
  INV_X1 U7061 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8762) );
  MUX2_X1 U7062 ( .A(n7176), .B(n8762), .S(n4443), .Z(n5551) );
  INV_X1 U7063 ( .A(SI_25_), .ZN(n5550) );
  NAND2_X1 U7064 ( .A1(n5551), .A2(n5550), .ZN(n5567) );
  INV_X1 U7065 ( .A(n5551), .ZN(n5552) );
  NAND2_X1 U7066 ( .A1(n5552), .A2(SI_25_), .ZN(n5553) );
  XNOR2_X1 U7067 ( .A(n5566), .B(n5565), .ZN(n7386) );
  NAND2_X1 U7068 ( .A1(n7386), .A2(n7900), .ZN(n5555) );
  NAND2_X2 U7069 ( .A1(n5555), .A2(n5554), .ZN(n8867) );
  INV_X1 U7070 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7071 ( .A1(n5558), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7072 ( .A1(n5575), .A2(n5559), .ZN(n7809) );
  NAND2_X1 U7073 ( .A1(n7809), .A2(n5343), .ZN(n5564) );
  INV_X1 U7074 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U7075 ( .A1(n7913), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7076 ( .A1(n4442), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5560) );
  OAI211_X1 U7077 ( .C1(n5630), .C2(n8800), .A(n5561), .B(n5560), .ZN(n5562)
         );
  INV_X1 U7078 ( .A(n5562), .ZN(n5563) );
  AND2_X1 U7079 ( .A1(n8867), .A2(n8328), .ZN(n7921) );
  INV_X1 U7080 ( .A(n8327), .ZN(n5582) );
  NAND2_X1 U7081 ( .A1(n5566), .A2(n5565), .ZN(n5568) );
  INV_X1 U7082 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8953) );
  INV_X1 U7083 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9778) );
  MUX2_X1 U7084 ( .A(n8953), .B(n9778), .S(n4443), .Z(n5570) );
  INV_X1 U7085 ( .A(SI_26_), .ZN(n5569) );
  NAND2_X1 U7086 ( .A1(n5570), .A2(n5569), .ZN(n5587) );
  INV_X1 U7087 ( .A(n5570), .ZN(n5571) );
  NAND2_X1 U7088 ( .A1(n5571), .A2(SI_26_), .ZN(n5572) );
  NAND2_X1 U7089 ( .A1(n8952), .A2(n7900), .ZN(n5574) );
  NAND2_X1 U7090 ( .A1(n5575), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7091 ( .A1(n5596), .A2(n5576), .ZN(n8332) );
  NAND2_X1 U7092 ( .A1(n8332), .A2(n5343), .ZN(n5581) );
  INV_X1 U7093 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U7094 ( .A1(n7911), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7095 ( .A1(n7913), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5577) );
  OAI211_X1 U7096 ( .C1(n5630), .C2(n8797), .A(n5578), .B(n5577), .ZN(n5579)
         );
  INV_X1 U7097 ( .A(n5579), .ZN(n5580) );
  NAND2_X1 U7098 ( .A1(n8861), .A2(n8338), .ZN(n5583) );
  INV_X1 U7099 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8950) );
  INV_X1 U7100 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8764) );
  MUX2_X1 U7101 ( .A(n8950), .B(n8764), .S(n4443), .Z(n5589) );
  INV_X1 U7102 ( .A(SI_27_), .ZN(n8759) );
  NAND2_X1 U7103 ( .A1(n5589), .A2(n8759), .ZN(n5607) );
  INV_X1 U7104 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7105 ( .A1(n5590), .A2(SI_27_), .ZN(n5591) );
  NAND2_X1 U7106 ( .A1(n8947), .A2(n7900), .ZN(n5593) );
  OR2_X1 U7107 ( .A1(n5746), .A2(n8950), .ZN(n5592) );
  INV_X1 U7108 ( .A(n5596), .ZN(n5595) );
  INV_X1 U7109 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7110 ( .A1(n5596), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7111 ( .A1(n5610), .A2(n5597), .ZN(n8323) );
  NAND2_X1 U7112 ( .A1(n8323), .A2(n5343), .ZN(n5602) );
  INV_X1 U7113 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U7114 ( .A1(n7912), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7115 ( .A1(n7911), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5598) );
  OAI211_X1 U7116 ( .C1(n5756), .C2(n8854), .A(n5599), .B(n5598), .ZN(n5600)
         );
  INV_X1 U7117 ( .A(n5600), .ZN(n5601) );
  NOR2_X1 U7118 ( .A1(n7732), .A2(n7881), .ZN(n5604) );
  NAND2_X1 U7119 ( .A1(n7732), .A2(n7881), .ZN(n5603) );
  INV_X1 U7120 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9771) );
  MUX2_X1 U7121 ( .A(n8945), .B(n9771), .S(n4443), .Z(n5745) );
  NAND2_X1 U7122 ( .A1(n9770), .A2(n7900), .ZN(n5609) );
  OR2_X1 U7123 ( .A1(n5746), .A2(n8945), .ZN(n5608) );
  NAND2_X1 U7124 ( .A1(n5610), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7125 ( .A1(n5626), .A2(n5611), .ZN(n7780) );
  NAND2_X1 U7126 ( .A1(n7780), .A2(n5266), .ZN(n5616) );
  NAND2_X1 U7127 ( .A1(n7911), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7128 ( .A1(n7913), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5612) );
  OAI211_X1 U7129 ( .C1(n5630), .C2(n5685), .A(n5613), .B(n5612), .ZN(n5614)
         );
  INV_X1 U7130 ( .A(n5614), .ZN(n5615) );
  XNOR2_X1 U7131 ( .A(n5741), .B(n5617), .ZN(n5638) );
  INV_X1 U7132 ( .A(n5618), .ZN(n5622) );
  NAND2_X1 U7133 ( .A1(n5622), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7134 ( .A1(n8296), .A2(n8118), .ZN(n5713) );
  NAND2_X1 U7135 ( .A1(n5620), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5621) );
  MUX2_X1 U7136 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5621), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5623) );
  NAND2_X1 U7137 ( .A1(n4491), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5625) );
  INV_X1 U7138 ( .A(n8100), .ZN(n5712) );
  NAND2_X1 U7139 ( .A1(n7961), .A2(n5712), .ZN(n8113) );
  NAND2_X1 U7140 ( .A1(n7670), .A2(n5343), .ZN(n7918) );
  INV_X1 U7141 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7142 ( .A1(n4442), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7143 ( .A1(n5456), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5627) );
  OAI211_X1 U7144 ( .C1(n5630), .C2(n5629), .A(n5628), .B(n5627), .ZN(n5631)
         );
  INV_X1 U7145 ( .A(n5631), .ZN(n5632) );
  NAND2_X1 U7146 ( .A1(n5856), .A2(n8116), .ZN(n5635) );
  NAND2_X1 U7147 ( .A1(n7905), .A2(n5635), .ZN(n5914) );
  INV_X1 U7148 ( .A(n5914), .ZN(n5636) );
  OAI22_X1 U7149 ( .A1(n7953), .A2(n8481), .B1(n7881), .B2(n8480), .ZN(n5637)
         );
  AOI21_X1 U7150 ( .B1(n5638), .B2(n8461), .A(n5637), .ZN(n5730) );
  INV_X1 U7151 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7152 ( .A1(n5640), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5641) );
  MUX2_X1 U7153 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5641), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n5643) );
  NAND2_X1 U7154 ( .A1(n5643), .A2(n5642), .ZN(n5652) );
  XNOR2_X1 U7155 ( .A(n5652), .B(P2_B_REG_SCAN_IN), .ZN(n5645) );
  NOR2_X1 U7156 ( .A1(n5646), .A2(n5405), .ZN(n5649) );
  INV_X1 U7157 ( .A(n5649), .ZN(n5648) );
  NAND2_X1 U7158 ( .A1(n5648), .A2(n5647), .ZN(n5651) );
  NAND2_X1 U7159 ( .A1(n5649), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5650) );
  INV_X1 U7160 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7161 ( .A1(n5656), .A2(n5993), .ZN(n5655) );
  NAND2_X1 U7162 ( .A1(n4575), .A2(n5653), .ZN(n5654) );
  AND2_X2 U7163 ( .A1(n5655), .A2(n5654), .ZN(n5874) );
  INV_X1 U7164 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7165 ( .A1(n5989), .A2(n5657), .ZN(n5660) );
  NAND2_X1 U7166 ( .A1(n4575), .A2(n5658), .ZN(n5659) );
  NAND2_X1 U7167 ( .A1(n5874), .A2(n8936), .ZN(n5711) );
  INV_X1 U7168 ( .A(n5658), .ZN(n5662) );
  INV_X1 U7169 ( .A(n5653), .ZN(n5661) );
  NAND3_X1 U7170 ( .A1(n5663), .A2(n5662), .A3(n5661), .ZN(n5902) );
  INV_X1 U7171 ( .A(n5664), .ZN(n5665) );
  NAND2_X1 U7172 ( .A1(n5665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5667) );
  NOR2_X1 U7173 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .ZN(
        n5671) );
  NOR4_X1 U7174 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5670) );
  NOR4_X1 U7175 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5669) );
  NOR4_X1 U7176 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n5668) );
  NAND4_X1 U7177 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n5677)
         );
  NOR4_X1 U7178 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5675) );
  NOR4_X1 U7179 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5674) );
  NOR4_X1 U7180 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5673) );
  NOR4_X1 U7181 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5672) );
  NAND4_X1 U7182 ( .A1(n5675), .A2(n5674), .A3(n5673), .A4(n5672), .ZN(n5676)
         );
  OAI21_X1 U7183 ( .B1(n5677), .B2(n5676), .A(n5989), .ZN(n5710) );
  NAND2_X1 U7184 ( .A1(n5876), .A2(n8103), .ZN(n5900) );
  AND3_X1 U7185 ( .A1(n8935), .A2(n5710), .A3(n5900), .ZN(n5678) );
  AND2_X1 U7186 ( .A1(n5711), .A2(n5678), .ZN(n5727) );
  INV_X1 U7187 ( .A(n5874), .ZN(n5680) );
  NAND2_X1 U7188 ( .A1(n8296), .A2(n8100), .ZN(n5732) );
  NOR2_X1 U7189 ( .A1(n10236), .A2(n7961), .ZN(n5729) );
  NAND2_X1 U7190 ( .A1(n8291), .A2(n8118), .ZN(n5704) );
  OR2_X1 U7191 ( .A1(n5704), .A2(n8100), .ZN(n5679) );
  OAI21_X1 U7192 ( .B1(n5680), .B2(n5729), .A(n5726), .ZN(n5683) );
  INV_X1 U7193 ( .A(n8936), .ZN(n5716) );
  INV_X1 U7194 ( .A(n5726), .ZN(n5681) );
  NAND2_X1 U7195 ( .A1(n5716), .A2(n5681), .ZN(n5682) );
  AND2_X1 U7196 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  MUX2_X1 U7197 ( .A(n5685), .B(n5730), .S(n10289), .Z(n5709) );
  OR2_X1 U7198 ( .A1(n5686), .A2(n5884), .ZN(n6578) );
  NAND2_X1 U7199 ( .A1(n6578), .A2(n5687), .ZN(n6528) );
  NAND2_X1 U7200 ( .A1(n6528), .A2(n7971), .ZN(n5688) );
  INV_X1 U7201 ( .A(n6537), .ZN(n7973) );
  NAND2_X1 U7202 ( .A1(n8134), .A2(n7973), .ZN(n7974) );
  NAND2_X1 U7203 ( .A1(n5688), .A2(n7974), .ZN(n6454) );
  INV_X1 U7204 ( .A(n7926), .ZN(n6455) );
  NAND2_X1 U7205 ( .A1(n6454), .A2(n6455), .ZN(n5689) );
  NAND2_X1 U7206 ( .A1(n5689), .A2(n7982), .ZN(n6552) );
  INV_X1 U7207 ( .A(n6602), .ZN(n10251) );
  NAND2_X1 U7208 ( .A1(n8132), .A2(n10251), .ZN(n7985) );
  NAND2_X1 U7209 ( .A1(n6552), .A2(n7985), .ZN(n5690) );
  INV_X1 U7210 ( .A(n8132), .ZN(n6760) );
  NAND2_X1 U7211 ( .A1(n6760), .A2(n6602), .ZN(n7998) );
  NAND2_X1 U7212 ( .A1(n5690), .A2(n7998), .ZN(n6716) );
  NAND2_X1 U7213 ( .A1(n6829), .A2(n6722), .ZN(n7999) );
  NAND2_X1 U7214 ( .A1(n8131), .A2(n10256), .ZN(n7983) );
  NAND2_X1 U7215 ( .A1(n6775), .A2(n7999), .ZN(n5691) );
  NAND2_X1 U7216 ( .A1(n6894), .A2(n6840), .ZN(n8004) );
  NAND2_X1 U7217 ( .A1(n8130), .A2(n10262), .ZN(n7984) );
  NAND2_X1 U7218 ( .A1(n5691), .A2(n7929), .ZN(n6773) );
  NAND2_X1 U7219 ( .A1(n6773), .A2(n8004), .ZN(n6899) );
  INV_X1 U7220 ( .A(n7086), .ZN(n10271) );
  NAND2_X1 U7221 ( .A1(n8128), .A2(n10271), .ZN(n7957) );
  AND2_X1 U7222 ( .A1(n6961), .A2(n7957), .ZN(n8013) );
  NAND2_X1 U7223 ( .A1(n6898), .A2(n8013), .ZN(n5692) );
  NAND2_X1 U7224 ( .A1(n7088), .A2(n7086), .ZN(n7958) );
  NAND2_X1 U7225 ( .A1(n5692), .A2(n7958), .ZN(n7072) );
  NAND2_X1 U7226 ( .A1(n7051), .A2(n10227), .ZN(n7992) );
  NAND2_X1 U7227 ( .A1(n7182), .A2(n8127), .ZN(n8008) );
  NAND2_X1 U7228 ( .A1(n7992), .A2(n8008), .ZN(n7933) );
  OR2_X1 U7229 ( .A1(n7765), .A2(n7210), .ZN(n8014) );
  NAND2_X1 U7230 ( .A1(n7765), .A2(n7210), .ZN(n8020) );
  NAND2_X1 U7231 ( .A1(n8014), .A2(n8020), .ZN(n7052) );
  NAND2_X1 U7232 ( .A1(n8779), .A2(n7801), .ZN(n7991) );
  OR2_X2 U7233 ( .A1(n8779), .A2(n7801), .ZN(n8007) );
  INV_X1 U7234 ( .A(n7679), .ZN(n7806) );
  NAND2_X1 U7235 ( .A1(n7806), .A2(n8124), .ZN(n8026) );
  INV_X1 U7236 ( .A(n8124), .ZN(n8479) );
  NAND2_X1 U7237 ( .A1(n7679), .A2(n8479), .ZN(n8027) );
  NAND2_X1 U7238 ( .A1(n7194), .A2(n8029), .ZN(n5693) );
  NAND2_X1 U7239 ( .A1(n5693), .A2(n8026), .ZN(n8485) );
  NOR2_X1 U7240 ( .A1(n8929), .A2(n5694), .ZN(n8032) );
  NAND2_X1 U7241 ( .A1(n8929), .A2(n5694), .ZN(n7938) );
  INV_X1 U7242 ( .A(n8923), .ZN(n8459) );
  NAND2_X1 U7243 ( .A1(n8459), .A2(n8451), .ZN(n8037) );
  NAND2_X1 U7244 ( .A1(n8923), .A2(n4972), .ZN(n8034) );
  INV_X1 U7245 ( .A(n8464), .ZN(n7743) );
  OR2_X1 U7246 ( .A1(n8916), .A2(n7743), .ZN(n8035) );
  NAND2_X1 U7247 ( .A1(n8448), .A2(n8035), .ZN(n5695) );
  NAND2_X1 U7248 ( .A1(n8916), .A2(n7743), .ZN(n8039) );
  NAND2_X1 U7249 ( .A1(n5695), .A2(n8039), .ZN(n8435) );
  INV_X1 U7250 ( .A(n5696), .ZN(n8043) );
  NAND2_X1 U7251 ( .A1(n8903), .A2(n8424), .ZN(n8046) );
  NAND2_X1 U7252 ( .A1(n8048), .A2(n8046), .ZN(n8413) );
  INV_X1 U7253 ( .A(n8411), .ZN(n5697) );
  NOR2_X1 U7254 ( .A1(n8413), .A2(n5697), .ZN(n5699) );
  INV_X1 U7255 ( .A(n8048), .ZN(n5698) );
  NAND2_X1 U7256 ( .A1(n8401), .A2(n8047), .ZN(n5700) );
  NAND2_X1 U7257 ( .A1(n5700), .A2(n8051), .ZN(n8396) );
  NAND2_X1 U7258 ( .A1(n8396), .A2(n8055), .ZN(n8378) );
  AND2_X1 U7259 ( .A1(n8060), .A2(n8377), .ZN(n8056) );
  NAND2_X1 U7260 ( .A1(n8378), .A2(n8056), .ZN(n5701) );
  INV_X1 U7261 ( .A(n8385), .ZN(n8063) );
  OR2_X1 U7262 ( .A1(n8884), .A2(n8063), .ZN(n8065) );
  NAND2_X1 U7263 ( .A1(n7839), .A2(n7750), .ZN(n8071) );
  NAND2_X1 U7264 ( .A1(n8878), .A2(n8349), .ZN(n8352) );
  NOR2_X1 U7265 ( .A1(n8867), .A2(n8348), .ZN(n8081) );
  NAND2_X1 U7266 ( .A1(n8867), .A2(n8348), .ZN(n8079) );
  NAND2_X1 U7267 ( .A1(n8855), .A2(n7881), .ZN(n8089) );
  NAND2_X1 U7268 ( .A1(n8317), .A2(n8089), .ZN(n5703) );
  NAND2_X1 U7269 ( .A1(n5703), .A2(n8088), .ZN(n5751) );
  XNOR2_X1 U7270 ( .A(n5751), .B(n7919), .ZN(n5736) );
  INV_X1 U7271 ( .A(n8118), .ZN(n7045) );
  NAND2_X1 U7272 ( .A1(n5876), .A2(n5704), .ZN(n5705) );
  INV_X1 U7273 ( .A(n10270), .ZN(n10244) );
  NAND2_X1 U7274 ( .A1(n7785), .A2(n8843), .ZN(n5706) );
  NAND2_X1 U7275 ( .A1(n5709), .A2(n5708), .ZN(P2_U3487) );
  INV_X1 U7276 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5721) );
  INV_X1 U7277 ( .A(n5710), .ZN(n5715) );
  NOR2_X1 U7278 ( .A1(n5711), .A2(n5715), .ZN(n5899) );
  NAND2_X1 U7279 ( .A1(n5899), .A2(n8935), .ZN(n5910) );
  NAND2_X1 U7280 ( .A1(n6969), .A2(n5712), .ZN(n5873) );
  AND2_X1 U7281 ( .A1(n6367), .A2(n5905), .ZN(n5714) );
  OR2_X1 U7282 ( .A1(n5910), .A2(n5714), .ZN(n5720) );
  NOR2_X1 U7283 ( .A1(n5874), .A2(n5715), .ZN(n5717) );
  AND2_X1 U7284 ( .A1(n5717), .A2(n5716), .ZN(n5907) );
  NAND2_X1 U7285 ( .A1(n5907), .A2(n8935), .ZN(n5916) );
  NOR2_X1 U7286 ( .A1(n10244), .A2(n8103), .ZN(n5718) );
  NAND2_X1 U7287 ( .A1(n5905), .A2(n5718), .ZN(n5890) );
  NAND2_X1 U7288 ( .A1(n5732), .A2(n10244), .ZN(n8458) );
  AND2_X1 U7289 ( .A1(n5890), .A2(n8458), .ZN(n5898) );
  MUX2_X1 U7290 ( .A(n5721), .B(n5730), .S(n10275), .Z(n5725) );
  NAND2_X1 U7291 ( .A1(n7785), .A2(n8930), .ZN(n5722) );
  NAND2_X1 U7292 ( .A1(n5725), .A2(n5724), .ZN(P2_U3455) );
  INV_X1 U7293 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5731) );
  MUX2_X1 U7294 ( .A(n5874), .B(n8936), .S(n5726), .Z(n5728) );
  NAND2_X1 U7295 ( .A1(n5728), .A2(n5727), .ZN(n5733) );
  MUX2_X1 U7296 ( .A(n5731), .B(n5730), .S(n10233), .Z(n5739) );
  NOR2_X1 U7297 ( .A1(n5732), .A2(n6969), .ZN(n6545) );
  OR2_X1 U7298 ( .A1(n6719), .A2(n6545), .ZN(n10222) );
  INV_X1 U7299 ( .A(n5733), .ZN(n5734) );
  INV_X1 U7300 ( .A(n8458), .ZN(n8482) );
  AOI22_X1 U7301 ( .A1(n7785), .A2(n10226), .B1(n10228), .B2(n7780), .ZN(n5735) );
  NAND2_X1 U7302 ( .A1(n5739), .A2(n5738), .ZN(P2_U3205) );
  NOR2_X1 U7303 ( .A1(n7785), .A2(n8320), .ZN(n5740) );
  INV_X1 U7304 ( .A(n7785), .ZN(n8106) );
  INV_X1 U7305 ( .A(n8320), .ZN(n8095) );
  INV_X1 U7306 ( .A(SI_28_), .ZN(n5744) );
  INV_X1 U7307 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8941) );
  INV_X1 U7308 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9768) );
  MUX2_X1 U7309 ( .A(n8941), .B(n9768), .S(n4443), .Z(n7242) );
  NAND2_X1 U7310 ( .A1(n7259), .A2(n7900), .ZN(n5748) );
  OR2_X1 U7311 ( .A1(n5746), .A2(n8941), .ZN(n5747) );
  NAND2_X1 U7312 ( .A1(n7951), .A2(n7953), .ZN(n7908) );
  NAND2_X1 U7313 ( .A1(n8102), .A2(n7908), .ZN(n7946) );
  XNOR2_X1 U7314 ( .A(n5749), .B(n7946), .ZN(n5761) );
  NAND2_X1 U7315 ( .A1(n7785), .A2(n8095), .ZN(n5750) );
  NAND2_X1 U7316 ( .A1(n5751), .A2(n5750), .ZN(n5753) );
  OR2_X1 U7317 ( .A1(n7785), .A2(n8095), .ZN(n5752) );
  NAND2_X1 U7318 ( .A1(n5762), .A2(n6719), .ZN(n5760) );
  INV_X1 U7319 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U7320 ( .A1(n7912), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U7321 ( .A1(n7911), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5754) );
  OAI211_X1 U7322 ( .C1(n5756), .C2(n8638), .A(n5755), .B(n5754), .ZN(n5757)
         );
  INV_X1 U7323 ( .A(n5757), .ZN(n5758) );
  NAND2_X1 U7324 ( .A1(n7918), .A2(n5758), .ZN(n8123) );
  AOI21_X1 U7325 ( .B1(P2_B_REG_SCAN_IN), .B2(n7905), .A(n8481), .ZN(n8311) );
  AOI22_X1 U7326 ( .A1(n8466), .A2(n8320), .B1(n8123), .B2(n8311), .ZN(n5759)
         );
  NOR2_X1 U7327 ( .A1(n7672), .A2(n8909), .ZN(n5765) );
  NOR2_X1 U7328 ( .A1(n10275), .A2(n5766), .ZN(n5767) );
  NAND2_X1 U7329 ( .A1(n5769), .A2(n5768), .ZN(P2_U3456) );
  INV_X1 U7330 ( .A(n10289), .ZN(n5770) );
  NAND2_X1 U7331 ( .A1(n5772), .A2(n5044), .ZN(P2_U3488) );
  NOR2_X1 U7332 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5776) );
  NAND4_X1 U7333 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n6214)
         );
  NAND3_X1 U7334 ( .A1(n5984), .A2(n6218), .A3(n5777), .ZN(n5778) );
  NOR2_X1 U7335 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5784) );
  NOR2_X1 U7336 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5783) );
  NOR2_X1 U7337 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5782) );
  INV_X1 U7338 ( .A(n6012), .ZN(n5791) );
  NAND2_X1 U7339 ( .A1(n4492), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5788) );
  MUX2_X1 U7340 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5788), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5789) );
  AND2_X1 U7341 ( .A1(n5787), .A2(n5789), .ZN(n5999) );
  NAND2_X1 U7342 ( .A1(n5787), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5790) );
  MUX2_X1 U7343 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5790), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5792) );
  NOR2_X1 U7344 ( .A1(n6171), .A2(P1_U3086), .ZN(n5798) );
  INV_X1 U7345 ( .A(n5793), .ZN(n5794) );
  INV_X1 U7346 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7347 ( .A1(n6017), .A2(n5795), .ZN(n5796) );
  NAND2_X1 U7348 ( .A1(n5796), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5797) );
  INV_X1 U7349 ( .A(n5901), .ZN(n7121) );
  NAND2_X1 U7350 ( .A1(n5901), .A2(n8103), .ZN(n5799) );
  NAND2_X1 U7351 ( .A1(n5858), .A2(n5799), .ZN(n5855) );
  OAI21_X1 U7352 ( .B1(n5855), .B2(n5800), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  INV_X4 U7353 ( .A(n8116), .ZN(n8292) );
  MUX2_X1 U7354 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8292), .Z(n7154) );
  INV_X1 U7355 ( .A(n5864), .ZN(n7163) );
  XNOR2_X1 U7356 ( .A(n7154), .B(n7163), .ZN(n7155) );
  MUX2_X1 U7357 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8292), .Z(n5806) );
  MUX2_X1 U7358 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8292), .Z(n5805) );
  MUX2_X1 U7359 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8292), .Z(n5804) );
  MUX2_X1 U7360 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8292), .Z(n5803) );
  MUX2_X1 U7361 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8292), .Z(n5802) );
  MUX2_X1 U7362 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n5634), .Z(n5801) );
  INV_X1 U7363 ( .A(n5835), .ZN(n5973) );
  XOR2_X1 U7364 ( .A(n5835), .B(n5801), .Z(n5945) );
  INV_X1 U7365 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6371) );
  INV_X1 U7366 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8704) );
  MUX2_X1 U7367 ( .A(n6371), .B(n8704), .S(n8292), .Z(n6256) );
  AND2_X1 U7368 ( .A1(n6256), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6258) );
  NOR2_X1 U7369 ( .A1(n5945), .A2(n6258), .ZN(n5944) );
  AOI21_X1 U7370 ( .B1(n5801), .B2(n5973), .A(n5944), .ZN(n6377) );
  XNOR2_X1 U7371 ( .A(n5802), .B(n6391), .ZN(n6378) );
  NOR2_X1 U7372 ( .A1(n6377), .A2(n6378), .ZN(n6376) );
  AOI21_X1 U7373 ( .B1(n5802), .B2(n6391), .A(n6376), .ZN(n6397) );
  XOR2_X1 U7374 ( .A(n5803), .B(n6400), .Z(n6396) );
  NAND2_X1 U7375 ( .A1(n6397), .A2(n6396), .ZN(n6395) );
  OAI21_X1 U7376 ( .B1(n5803), .B2(n6400), .A(n6395), .ZN(n5924) );
  XNOR2_X1 U7377 ( .A(n5804), .B(n5970), .ZN(n5925) );
  AOI21_X1 U7378 ( .B1(n5804), .B2(n5970), .A(n5923), .ZN(n6745) );
  XNOR2_X1 U7379 ( .A(n5805), .B(n6754), .ZN(n6746) );
  NOR2_X1 U7380 ( .A1(n6745), .A2(n6746), .ZN(n6744) );
  XOR2_X1 U7381 ( .A(n6807), .B(n5806), .Z(n6804) );
  MUX2_X1 U7382 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8292), .Z(n5807) );
  XOR2_X1 U7383 ( .A(n6004), .B(n5807), .Z(n6931) );
  INV_X1 U7384 ( .A(n5807), .ZN(n5808) );
  MUX2_X1 U7385 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8292), .Z(n5809) );
  XNOR2_X1 U7386 ( .A(n5809), .B(n6979), .ZN(n6972) );
  MUX2_X1 U7387 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8292), .Z(n5810) );
  XNOR2_X1 U7388 ( .A(n5810), .B(n5850), .ZN(n7058) );
  INV_X1 U7389 ( .A(n5810), .ZN(n5811) );
  XOR2_X1 U7390 ( .A(n7155), .B(n7156), .Z(n5812) );
  NOR2_X1 U7391 ( .A1(n5812), .A2(n7070), .ZN(n5872) );
  INV_X1 U7392 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6540) );
  XNOR2_X1 U7393 ( .A(n6391), .B(n6540), .ZN(n6387) );
  NAND2_X1 U7394 ( .A1(n5833), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7395 ( .A1(n5835), .A2(n5813), .ZN(n5814) );
  NAND2_X1 U7396 ( .A1(n5814), .A2(n5815), .ZN(n5954) );
  INV_X1 U7397 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10278) );
  OR2_X1 U7398 ( .A1(n5954), .A2(n10278), .ZN(n5952) );
  NAND2_X1 U7399 ( .A1(n5952), .A2(n5815), .ZN(n6386) );
  NAND2_X1 U7400 ( .A1(n6387), .A2(n6386), .ZN(n6385) );
  NAND2_X1 U7401 ( .A1(n6391), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7402 ( .A1(n6385), .A2(n5816), .ZN(n5817) );
  NAND2_X1 U7403 ( .A1(n5817), .A2(n6400), .ZN(n5932) );
  OR2_X1 U7404 ( .A1(n5817), .A2(n6400), .ZN(n5818) );
  AND2_X1 U7405 ( .A1(n5932), .A2(n5818), .ZN(n6403) );
  NAND2_X1 U7406 ( .A1(n6402), .A2(n5932), .ZN(n5819) );
  INV_X1 U7407 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10282) );
  MUX2_X1 U7408 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10282), .S(n5970), .Z(n5934)
         );
  NAND2_X1 U7409 ( .A1(n5970), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7410 ( .A1(n5821), .A2(n6754), .ZN(n6815) );
  NAND2_X1 U7411 ( .A1(n6747), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U7412 ( .A1(n6817), .A2(n6815), .ZN(n5822) );
  INV_X1 U7413 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10286) );
  MUX2_X1 U7414 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10286), .S(n6807), .Z(n6814)
         );
  NAND2_X1 U7415 ( .A1(n6807), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7416 ( .A1(n5824), .A2(n6004), .ZN(n6974) );
  NAND2_X1 U7417 ( .A1(n6976), .A2(n6974), .ZN(n5826) );
  INV_X1 U7418 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5825) );
  XNOR2_X1 U7419 ( .A(n6979), .B(n5825), .ZN(n6973) );
  NAND2_X1 U7420 ( .A1(n5826), .A2(n6973), .ZN(n6978) );
  NAND2_X1 U7421 ( .A1(n6979), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5827) );
  INV_X1 U7422 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7078) );
  INV_X1 U7423 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5828) );
  XNOR2_X1 U7424 ( .A(n5864), .B(n5828), .ZN(n5830) );
  AOI21_X1 U7425 ( .B1(n7065), .B2(n5829), .A(n5830), .ZN(n7160) );
  INV_X1 U7426 ( .A(n7160), .ZN(n5832) );
  NAND3_X1 U7427 ( .A1(n7065), .A2(n5830), .A3(n5829), .ZN(n5831) );
  OR2_X1 U7428 ( .A1(n5633), .A2(P2_U3151), .ZN(n8943) );
  NOR2_X1 U7429 ( .A1(n5855), .A2(n8943), .ZN(n6259) );
  AOI21_X1 U7430 ( .B1(n5832), .B2(n5831), .A(n8310), .ZN(n5871) );
  INV_X1 U7431 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6548) );
  XNOR2_X1 U7432 ( .A(n6391), .B(n6548), .ZN(n6381) );
  NAND2_X1 U7433 ( .A1(n5833), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7434 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  NAND2_X1 U7435 ( .A1(n5836), .A2(n5837), .ZN(n5948) );
  INV_X1 U7436 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5949) );
  OR2_X1 U7437 ( .A1(n5948), .A2(n5949), .ZN(n5946) );
  NAND2_X1 U7438 ( .A1(n5946), .A2(n5837), .ZN(n6380) );
  NAND2_X1 U7439 ( .A1(n6381), .A2(n6380), .ZN(n6379) );
  NAND2_X1 U7440 ( .A1(n6391), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5838) );
  INV_X1 U7441 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5840) );
  MUX2_X1 U7442 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n5840), .S(n5970), .Z(n5926)
         );
  NAND2_X1 U7443 ( .A1(n5841), .A2(n5926), .ZN(n5930) );
  NAND2_X1 U7444 ( .A1(n5970), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7445 ( .A1(n5843), .A2(n6754), .ZN(n6809) );
  NAND2_X1 U7446 ( .A1(n6811), .A2(n6809), .ZN(n5845) );
  INV_X1 U7447 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5844) );
  MUX2_X1 U7448 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n5844), .S(n6807), .Z(n6808)
         );
  NAND2_X1 U7449 ( .A1(n6807), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U7450 ( .A1(n5847), .A2(n6004), .ZN(n6982) );
  NAND2_X1 U7451 ( .A1(n6935), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U7452 ( .A1(n6936), .A2(n6982), .ZN(n5848) );
  INV_X1 U7453 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6965) );
  XNOR2_X1 U7454 ( .A(n6979), .B(n6965), .ZN(n6983) );
  NAND2_X1 U7455 ( .A1(n6979), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5849) );
  INV_X1 U7456 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5852) );
  XNOR2_X1 U7457 ( .A(n5864), .B(n5852), .ZN(n5854) );
  NAND3_X1 U7458 ( .A1(n7059), .A2(n5854), .A3(n5853), .ZN(n5857) );
  OR2_X1 U7459 ( .A1(n8292), .A2(P2_U3151), .ZN(n8948) );
  NOR2_X1 U7460 ( .A1(n5855), .A2(n8948), .ZN(n5859) );
  NAND2_X1 U7461 ( .A1(n5859), .A2(n5856), .ZN(n8306) );
  AOI21_X1 U7462 ( .B1(n4528), .B2(n5857), .A(n8306), .ZN(n5870) );
  INV_X1 U7463 ( .A(n5858), .ZN(n5861) );
  INV_X1 U7464 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7465 ( .A1(n5859), .A2(n5633), .ZN(n5863) );
  INV_X1 U7466 ( .A(n8943), .ZN(n5860) );
  NAND2_X1 U7467 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  NAND2_X1 U7468 ( .A1(n5863), .A2(n5862), .ZN(n8297) );
  NAND2_X1 U7469 ( .A1(n8297), .A2(n5864), .ZN(n5867) );
  INV_X1 U7470 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5865) );
  NOR2_X1 U7471 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5865), .ZN(n7755) );
  INV_X1 U7472 ( .A(n7755), .ZN(n5866) );
  OAI211_X1 U7473 ( .C1(n8300), .C2(n5868), .A(n5867), .B(n5866), .ZN(n5869)
         );
  OR4_X1 U7474 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(P2_U3192)
         );
  INV_X1 U7475 ( .A(n5873), .ZN(n7950) );
  NAND2_X1 U7476 ( .A1(n5874), .A2(n7950), .ZN(n5878) );
  NAND2_X1 U7477 ( .A1(n7961), .A2(n8100), .ZN(n5875) );
  XNOR2_X1 U7478 ( .A(n10245), .B(n7778), .ZN(n6590) );
  XNOR2_X1 U7479 ( .A(n6591), .B(n6590), .ZN(n5897) );
  XNOR2_X1 U7480 ( .A(n6586), .B(n5886), .ZN(n5879) );
  NAND2_X1 U7481 ( .A1(n5880), .A2(n5879), .ZN(n5885) );
  INV_X1 U7482 ( .A(n5879), .ZN(n5881) );
  NAND2_X1 U7483 ( .A1(n5881), .A2(n5248), .ZN(n5882) );
  OR2_X1 U7484 ( .A1(n5886), .A2(n6298), .ZN(n5883) );
  NAND2_X1 U7485 ( .A1(n5884), .A2(n5883), .ZN(n6293) );
  NAND2_X1 U7486 ( .A1(n5051), .A2(n6293), .ZN(n6292) );
  NAND2_X1 U7487 ( .A1(n6292), .A2(n5885), .ZN(n6359) );
  XNOR2_X1 U7488 ( .A(n5887), .B(n8134), .ZN(n6360) );
  NAND2_X1 U7489 ( .A1(n6359), .A2(n6360), .ZN(n6358) );
  INV_X1 U7490 ( .A(n5887), .ZN(n5888) );
  NAND2_X1 U7491 ( .A1(n8134), .A2(n5888), .ZN(n5889) );
  NAND2_X1 U7492 ( .A1(n6358), .A2(n5889), .ZN(n5896) );
  OR2_X1 U7493 ( .A1(n5910), .A2(n5890), .ZN(n5892) );
  OR2_X1 U7494 ( .A1(n5916), .A2(n5905), .ZN(n5891) );
  INV_X1 U7495 ( .A(n5896), .ZN(n5894) );
  NAND2_X1 U7496 ( .A1(n5894), .A2(n5893), .ZN(n6593) );
  INV_X1 U7497 ( .A(n6593), .ZN(n5895) );
  AOI211_X1 U7498 ( .C1(n5897), .C2(n5896), .A(n7887), .B(n5895), .ZN(n5922)
         );
  OR2_X1 U7499 ( .A1(n5899), .A2(n5898), .ZN(n5904) );
  AND3_X1 U7500 ( .A1(n5902), .A2(n5901), .A3(n5900), .ZN(n5903) );
  OAI211_X1 U7501 ( .C1(n5907), .C2(n5905), .A(n5904), .B(n5903), .ZN(n5906)
         );
  NAND2_X1 U7502 ( .A1(n5906), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5909) );
  INV_X1 U7503 ( .A(n6367), .ZN(n5913) );
  NAND2_X1 U7504 ( .A1(n8935), .A2(n5913), .ZN(n8117) );
  OR2_X1 U7505 ( .A1(n5907), .A2(n8117), .ZN(n5908) );
  NOR2_X1 U7506 ( .A1(n7821), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5921) );
  OR2_X1 U7507 ( .A1(n5910), .A2(n10270), .ZN(n5911) );
  AND2_X1 U7508 ( .A1(n7883), .A2(n10245), .ZN(n5920) );
  OR2_X1 U7509 ( .A1(n5914), .A2(n6367), .ZN(n5912) );
  OR2_X1 U7510 ( .A1(n5916), .A2(n5912), .ZN(n7853) );
  NAND2_X1 U7511 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  NAND2_X1 U7512 ( .A1(n7850), .A2(n8132), .ZN(n5918) );
  AND2_X1 U7513 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6404) );
  INV_X1 U7514 ( .A(n6404), .ZN(n5917) );
  OAI211_X1 U7515 ( .C1(n8134), .C2(n7853), .A(n5918), .B(n5917), .ZN(n5919)
         );
  OR4_X1 U7516 ( .A1(n5922), .A2(n5921), .A3(n5920), .A4(n5919), .ZN(P2_U3158)
         );
  AOI211_X1 U7517 ( .C1(n5925), .C2(n5924), .A(n7070), .B(n5923), .ZN(n5943)
         );
  NOR2_X1 U7518 ( .A1(n8266), .A2(n5970), .ZN(n5942) );
  INV_X1 U7519 ( .A(n5926), .ZN(n5928) );
  NAND3_X1 U7520 ( .A1(n6398), .A2(n5928), .A3(n5927), .ZN(n5929) );
  AOI21_X1 U7521 ( .B1(n5930), .B2(n5929), .A(n8306), .ZN(n5941) );
  INV_X1 U7522 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n5939) );
  INV_X1 U7523 ( .A(n5931), .ZN(n5937) );
  INV_X1 U7524 ( .A(n6402), .ZN(n5935) );
  INV_X1 U7525 ( .A(n5932), .ZN(n5933) );
  NOR3_X1 U7526 ( .A1(n5935), .A2(n5934), .A3(n5933), .ZN(n5936) );
  INV_X1 U7527 ( .A(n8310), .ZN(n8140) );
  OAI21_X1 U7528 ( .B1(n5937), .B2(n5936), .A(n8140), .ZN(n5938) );
  NAND2_X1 U7529 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6600) );
  OAI211_X1 U7530 ( .C1(n5939), .C2(n8300), .A(n5938), .B(n6600), .ZN(n5940)
         );
  OR4_X1 U7531 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(P2_U3186)
         );
  AOI211_X1 U7532 ( .C1(n5945), .C2(n6258), .A(n7070), .B(n5944), .ZN(n5959)
         );
  INV_X1 U7533 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n5951) );
  INV_X1 U7534 ( .A(n5946), .ZN(n5947) );
  AOI21_X1 U7535 ( .B1(n5949), .B2(n5948), .A(n5947), .ZN(n5950) );
  OAI22_X1 U7536 ( .A1(n8300), .A2(n5951), .B1(n8306), .B2(n5950), .ZN(n5958)
         );
  NOR2_X1 U7537 ( .A1(n8266), .A2(n5973), .ZN(n5957) );
  INV_X1 U7538 ( .A(n5952), .ZN(n5953) );
  AOI21_X1 U7539 ( .B1(n10278), .B2(n5954), .A(n5953), .ZN(n5955) );
  INV_X1 U7540 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6297) );
  OAI22_X1 U7541 ( .A1(n8310), .A2(n5955), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6297), .ZN(n5956) );
  OR4_X1 U7542 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(P2_U3183)
         );
  XNOR2_X1 U7543 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U7544 ( .A1(n4443), .A2(P2_U3151), .ZN(n8939) );
  INV_X2 U7545 ( .A(n8939), .ZN(n8951) );
  OAI222_X1 U7546 ( .A1(n8951), .A2(n5961), .B1(n8954), .B2(n6309), .C1(
        P2_U3151), .C2(n6391), .ZN(P2_U3293) );
  OAI222_X1 U7547 ( .A1(n8951), .A2(n5962), .B1(n8954), .B2(n6414), .C1(
        P2_U3151), .C2(n6400), .ZN(P2_U3292) );
  NAND2_X1 U7548 ( .A1(n4443), .A2(P1_U3086), .ZN(n9773) );
  NOR2_X1 U7549 ( .A1(n5964), .A2(n6492), .ZN(n5965) );
  MUX2_X1 U7550 ( .A(n6492), .B(n5965), .S(P1_IR_REG_3__SCAN_IN), .Z(n5966) );
  INV_X1 U7551 ( .A(n5966), .ZN(n5969) );
  INV_X1 U7552 ( .A(n5983), .ZN(n5968) );
  NAND2_X1 U7553 ( .A1(n5969), .A2(n5968), .ZN(n9296) );
  OAI222_X1 U7554 ( .A1(n9769), .A2(n6415), .B1(n9773), .B2(n6414), .C1(
        P1_U3086), .C2(n9296), .ZN(P1_U3352) );
  OAI222_X1 U7555 ( .A1(n8951), .A2(n5971), .B1(n8954), .B2(n6465), .C1(
        P2_U3151), .C2(n5970), .ZN(P2_U3291) );
  INV_X1 U7556 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5974) );
  INV_X1 U7557 ( .A(n8946), .ZN(n7046) );
  INV_X1 U7558 ( .A(n5972), .ZN(n6264) );
  OAI222_X1 U7559 ( .A1(n8951), .A2(n5974), .B1(n7046), .B2(n6264), .C1(
        P2_U3151), .C2(n5973), .ZN(P2_U3294) );
  INV_X1 U7560 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U7561 ( .A1(n5983), .A2(n5984), .ZN(n6215) );
  NAND2_X1 U7562 ( .A1(n6215), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5975) );
  MUX2_X1 U7563 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5975), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5976) );
  NAND2_X1 U7564 ( .A1(n5976), .A2(n5994), .ZN(n6614) );
  OAI222_X1 U7565 ( .A1(n9769), .A2(n6611), .B1(n9773), .B2(n6610), .C1(
        P1_U3086), .C2(n6614), .ZN(P1_U3350) );
  OAI222_X1 U7566 ( .A1(n8951), .A2(n5977), .B1(n8954), .B2(n6610), .C1(
        P2_U3151), .C2(n6754), .ZN(P2_U3290) );
  INV_X1 U7567 ( .A(n9773), .ZN(n7119) );
  INV_X1 U7568 ( .A(n7119), .ZN(n9777) );
  XNOR2_X1 U7569 ( .A(n5980), .B(n5979), .ZN(n6310) );
  OAI222_X1 U7570 ( .A1(n9769), .A2(n6308), .B1(n9777), .B2(n6309), .C1(
        P1_U3086), .C2(n6310), .ZN(P1_U3353) );
  INV_X1 U7571 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7572 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9779), .ZN(n5981) );
  OAI222_X1 U7573 ( .A1(n9769), .A2(n4877), .B1(n9777), .B2(n6264), .C1(
        P1_U3086), .C2(n6267), .ZN(P1_U3354) );
  OR2_X1 U7574 ( .A1(n5983), .A2(n6492), .ZN(n5985) );
  OAI222_X1 U7575 ( .A1(n9769), .A2(n6464), .B1(n9777), .B2(n6465), .C1(
        P1_U3086), .C2(n9312), .ZN(P1_U3351) );
  OAI222_X1 U7576 ( .A1(n8951), .A2(n5986), .B1(n7046), .B2(n6688), .C1(
        P2_U3151), .C2(n6807), .ZN(P2_U3289) );
  NAND2_X1 U7577 ( .A1(n5994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5988) );
  INV_X1 U7578 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5987) );
  XNOR2_X1 U7579 ( .A(n5988), .B(n5987), .ZN(n6692) );
  OAI222_X1 U7580 ( .A1(n9769), .A2(n6689), .B1(n9777), .B2(n6688), .C1(
        P1_U3086), .C2(n6692), .ZN(P1_U3349) );
  INV_X1 U7581 ( .A(n5989), .ZN(n5990) );
  NAND2_X1 U7582 ( .A1(n8935), .A2(n5990), .ZN(n6046) );
  AND3_X1 U7583 ( .A1(n4575), .A2(n5991), .A3(n5653), .ZN(n5992) );
  AOI21_X1 U7584 ( .B1(n6046), .B2(n5993), .A(n5992), .ZN(P2_U3376) );
  NOR2_X1 U7585 ( .A1(n5994), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6008) );
  OR2_X1 U7586 ( .A1(n6008), .A2(n6492), .ZN(n5995) );
  XNOR2_X1 U7587 ( .A(n5995), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9802) );
  INV_X1 U7588 ( .A(n9769), .ZN(n6686) );
  AOI22_X1 U7589 ( .A1(n9802), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n6686), .ZN(n5996) );
  OAI21_X1 U7590 ( .B1(n6785), .B2(n9773), .A(n5996), .ZN(P1_U3348) );
  NAND2_X1 U7591 ( .A1(n7177), .A2(P1_B_REG_SCAN_IN), .ZN(n6000) );
  MUX2_X1 U7592 ( .A(P1_B_REG_SCAN_IN), .B(n6000), .S(n7175), .Z(n6001) );
  NAND2_X1 U7593 ( .A1(n6001), .A2(n6002), .ZN(n6165) );
  INV_X1 U7594 ( .A(n6002), .ZN(n9775) );
  AND2_X1 U7595 ( .A1(n9775), .A2(n7175), .ZN(n6160) );
  NAND2_X1 U7596 ( .A1(n10110), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6003) );
  OAI21_X1 U7597 ( .B1(n10110), .B2(n6160), .A(n6003), .ZN(P1_U3439) );
  OAI222_X1 U7598 ( .A1(n8951), .A2(n6005), .B1(n8954), .B2(n6785), .C1(
        P2_U3151), .C2(n6004), .ZN(P2_U3288) );
  INV_X1 U7599 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6163) );
  OR2_X1 U7600 ( .A1(n10110), .A2(n6162), .ZN(n6006) );
  OAI21_X1 U7601 ( .B1(n10109), .B2(n6163), .A(n6006), .ZN(P1_U3440) );
  INV_X1 U7602 ( .A(n6862), .ZN(n6045) );
  INV_X1 U7603 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7604 ( .A1(n6008), .A2(n6007), .ZN(n6116) );
  NAND2_X1 U7605 ( .A1(n6116), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6009) );
  XNOR2_X1 U7606 ( .A(n6009), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U7607 ( .A1(n9814), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n6686), .ZN(n6010) );
  OAI21_X1 U7608 ( .B1(n6045), .B2(n9773), .A(n6010), .ZN(P1_U3347) );
  INV_X1 U7609 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7610 ( .A1(n4433), .A2(n7599), .ZN(n6510) );
  NAND2_X1 U7611 ( .A1(n7485), .A2(n6020), .ZN(n6019) );
  AND2_X1 U7612 ( .A1(n6786), .A2(n6019), .ZN(n6223) );
  INV_X1 U7613 ( .A(n6223), .ZN(n6023) );
  INV_X1 U7614 ( .A(n6502), .ZN(n6022) );
  INV_X1 U7615 ( .A(n6020), .ZN(n6021) );
  AND2_X1 U7616 ( .A1(n6021), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6174) );
  INV_X1 U7617 ( .A(n6174), .ZN(n7667) );
  NAND2_X1 U7618 ( .A1(n6022), .A2(n7667), .ZN(n6224) );
  NOR2_X1 U7619 ( .A1(n9883), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U7620 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n6024) );
  AND2_X1 U7621 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6026) );
  INV_X1 U7622 ( .A(n6030), .ZN(n6032) );
  NOR3_X1 U7623 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .A3(
        P1_IR_REG_30__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7624 ( .A1(n6032), .A2(n6031), .ZN(n9759) );
  BUF_X4 U7625 ( .A(n6180), .Z(n7448) );
  INV_X1 U7626 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n6036) );
  OR2_X1 U7627 ( .A1(n7448), .A2(n6036), .ZN(n6043) );
  NAND2_X4 U7628 ( .A1(n9763), .A2(n6037), .ZN(n7445) );
  INV_X1 U7629 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6038) );
  OR2_X1 U7630 ( .A1(n7445), .A2(n6038), .ZN(n6042) );
  NAND2_X1 U7631 ( .A1(n9763), .A2(n9767), .ZN(n6281) );
  INV_X1 U7632 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6040) );
  OR2_X1 U7633 ( .A1(n4432), .A2(n6040), .ZN(n6041) );
  NAND2_X1 U7634 ( .A1(n9284), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6044) );
  OAI21_X1 U7635 ( .B1(n9472), .B2(n9284), .A(n6044), .ZN(P1_U3584) );
  OAI222_X1 U7636 ( .A1(n6979), .A2(P2_U3151), .B1(n8954), .B2(n6045), .C1(
        n8951), .C2(n5352), .ZN(P2_U3287) );
  INV_X1 U7637 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6047) );
  NOR2_X1 U7638 ( .A1(n6197), .A2(n6047), .ZN(P2_U3255) );
  INV_X1 U7639 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6048) );
  NOR2_X1 U7640 ( .A1(n6197), .A2(n6048), .ZN(P2_U3246) );
  INV_X1 U7641 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n6049) );
  NOR2_X1 U7642 ( .A1(n6197), .A2(n6049), .ZN(P2_U3250) );
  INV_X1 U7643 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n8614) );
  NOR2_X1 U7644 ( .A1(n6197), .A2(n8614), .ZN(P2_U3251) );
  INV_X1 U7645 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6050) );
  NOR2_X1 U7646 ( .A1(n6197), .A2(n6050), .ZN(P2_U3248) );
  INV_X1 U7647 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6051) );
  NOR2_X1 U7648 ( .A1(n6197), .A2(n6051), .ZN(P2_U3249) );
  INV_X1 U7649 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6052) );
  NOR2_X1 U7650 ( .A1(n6197), .A2(n6052), .ZN(P2_U3254) );
  INV_X1 U7651 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n6053) );
  NOR2_X1 U7652 ( .A1(n6197), .A2(n6053), .ZN(P2_U3247) );
  INV_X1 U7653 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6054) );
  NOR2_X1 U7654 ( .A1(n6197), .A2(n6054), .ZN(P2_U3252) );
  INV_X1 U7655 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6055) );
  NOR2_X1 U7656 ( .A1(n6197), .A2(n6055), .ZN(P2_U3257) );
  INV_X1 U7657 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n8753) );
  NOR2_X1 U7658 ( .A1(n6197), .A2(n8753), .ZN(P2_U3253) );
  INV_X1 U7659 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6056) );
  NOR2_X1 U7660 ( .A1(n6197), .A2(n6056), .ZN(P2_U3256) );
  INV_X1 U7661 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6906) );
  INV_X1 U7662 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6057) );
  OR2_X1 U7663 ( .A1(n7445), .A2(n6057), .ZN(n6058) );
  OAI21_X1 U7664 ( .B1(n7448), .B2(n6906), .A(n6058), .ZN(n6066) );
  OR2_X2 U7665 ( .A1(n9763), .A2(n9767), .ZN(n7319) );
  NAND3_X1 U7666 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6633) );
  INV_X1 U7667 ( .A(n6633), .ZN(n6059) );
  NAND2_X1 U7668 ( .A1(n6059), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6702) );
  INV_X1 U7669 ( .A(n6702), .ZN(n6060) );
  NAND2_X1 U7670 ( .A1(n6060), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6704) );
  INV_X1 U7671 ( .A(n6704), .ZN(n6061) );
  NAND2_X1 U7672 ( .A1(n6061), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6853) );
  INV_X1 U7673 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U7674 ( .A1(n6704), .A2(n8680), .ZN(n6062) );
  NAND2_X1 U7675 ( .A1(n6853), .A2(n6062), .ZN(n7039) );
  INV_X1 U7676 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6063) );
  OR2_X1 U7677 ( .A1(n4432), .A2(n6063), .ZN(n6064) );
  OAI21_X1 U7678 ( .B1(n7319), .B2(n7039), .A(n6064), .ZN(n6065) );
  NAND2_X1 U7679 ( .A1(n7111), .A2(P1_U3973), .ZN(n6067) );
  OAI21_X1 U7680 ( .B1(P1_U3973), .B2(n5352), .A(n6067), .ZN(P1_U3562) );
  INV_X1 U7681 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6211) );
  INV_X1 U7682 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6069) );
  INV_X1 U7683 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6673) );
  OR2_X1 U7684 ( .A1(n7445), .A2(n6673), .ZN(n6068) );
  OAI21_X1 U7685 ( .B1(n7448), .B2(n6069), .A(n6068), .ZN(n6074) );
  INV_X1 U7686 ( .A(n6853), .ZN(n6070) );
  NAND2_X1 U7687 ( .A1(n6070), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6871) );
  INV_X1 U7688 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6996) );
  XNOR2_X1 U7689 ( .A(n6997), .B(n6996), .ZN(n9999) );
  INV_X1 U7690 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6071) );
  OR2_X1 U7691 ( .A1(n4432), .A2(n6071), .ZN(n6072) );
  OAI21_X1 U7692 ( .B1(n7319), .B2(n9999), .A(n6072), .ZN(n6073) );
  NAND2_X1 U7693 ( .A1(n8963), .A2(P1_U3973), .ZN(n6075) );
  OAI21_X1 U7694 ( .B1(n6211), .B2(P1_U3973), .A(n6075), .ZN(P1_U3565) );
  INV_X1 U7695 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6082) );
  INV_X1 U7696 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6080) );
  INV_X1 U7697 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6076) );
  OR2_X1 U7698 ( .A1(n7296), .A2(n6076), .ZN(n6079) );
  INV_X1 U7699 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6077) );
  OR2_X1 U7700 ( .A1(n7445), .A2(n6077), .ZN(n6078) );
  OAI211_X1 U7701 ( .C1(n4431), .C2(n6080), .A(n6079), .B(n6078), .ZN(n7588)
         );
  NAND2_X1 U7702 ( .A1(n7588), .A2(P1_U3973), .ZN(n6081) );
  OAI21_X1 U7703 ( .B1(P1_U3973), .B2(n6082), .A(n6081), .ZN(P1_U3585) );
  INV_X1 U7704 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6085) );
  INV_X1 U7705 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6083) );
  OR2_X1 U7706 ( .A1(n7445), .A2(n6083), .ZN(n6084) );
  OAI21_X1 U7707 ( .B1(n7448), .B2(n6085), .A(n6084), .ZN(n6095) );
  NAND2_X1 U7708 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n6086) );
  INV_X1 U7709 ( .A(n6998), .ZN(n6087) );
  INV_X1 U7710 ( .A(n7292), .ZN(n6089) );
  AND2_X1 U7711 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n6088) );
  NAND2_X1 U7712 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n6090) );
  NAND2_X1 U7713 ( .A1(n6098), .A2(n9208), .ZN(n6092) );
  NAND2_X1 U7714 ( .A1(n7405), .A2(n6092), .ZN(n9205) );
  INV_X1 U7715 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8561) );
  OR2_X1 U7716 ( .A1(n4432), .A2(n8561), .ZN(n6093) );
  OAI21_X1 U7717 ( .B1(n7319), .B2(n9205), .A(n6093), .ZN(n6094) );
  NAND2_X1 U7718 ( .A1(n9435), .A2(P1_U3973), .ZN(n6096) );
  OAI21_X1 U7719 ( .B1(n5494), .B2(P1_U3973), .A(n6096), .ZN(P1_U3574) );
  INV_X1 U7720 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8603) );
  INV_X2 U7721 ( .A(n7450), .ZN(n7430) );
  INV_X1 U7722 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U7723 ( .A1(n7330), .A2(n9116), .ZN(n6097) );
  NAND2_X1 U7724 ( .A1(n6098), .A2(n6097), .ZN(n9618) );
  OR2_X1 U7725 ( .A1(n7430), .A2(n9618), .ZN(n6105) );
  INV_X1 U7726 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6099) );
  OR2_X1 U7727 ( .A1(n7448), .A2(n6099), .ZN(n6104) );
  INV_X1 U7728 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6100) );
  OR2_X1 U7729 ( .A1(n7445), .A2(n6100), .ZN(n6103) );
  INV_X1 U7730 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n6101) );
  OR2_X1 U7731 ( .A1(n4431), .A2(n6101), .ZN(n6102) );
  NAND4_X1 U7732 ( .A1(n6105), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(n9431)
         );
  NAND2_X1 U7733 ( .A1(n9431), .A2(P1_U3973), .ZN(n6106) );
  OAI21_X1 U7734 ( .B1(n8603), .B2(P1_U3973), .A(n6106), .ZN(P1_U3573) );
  INV_X1 U7735 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6350) );
  INV_X1 U7736 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U7737 ( .A1(n6998), .A2(n8748), .ZN(n6107) );
  NAND2_X1 U7738 ( .A1(n7292), .A2(n6107), .ZN(n9980) );
  OR2_X1 U7739 ( .A1(n7430), .A2(n9980), .ZN(n6114) );
  INV_X1 U7740 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6108) );
  OR2_X1 U7741 ( .A1(n7448), .A2(n6108), .ZN(n6113) );
  INV_X1 U7742 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6109) );
  OR2_X1 U7743 ( .A1(n4432), .A2(n6109), .ZN(n6112) );
  INV_X1 U7744 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6110) );
  OR2_X1 U7745 ( .A1(n7445), .A2(n6110), .ZN(n6111) );
  NAND4_X1 U7746 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(n9417)
         );
  NAND2_X1 U7747 ( .A1(n9417), .A2(P1_U3973), .ZN(n6115) );
  OAI21_X1 U7748 ( .B1(n6350), .B2(P1_U3973), .A(n6115), .ZN(P1_U3567) );
  INV_X1 U7749 ( .A(n6848), .ZN(n6120) );
  NAND2_X1 U7750 ( .A1(n6122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6117) );
  XNOR2_X1 U7751 ( .A(n6117), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6849) );
  AOI22_X1 U7752 ( .A1(n6849), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n6686), .ZN(n6118) );
  OAI21_X1 U7753 ( .B1(n6120), .B2(n9773), .A(n6118), .ZN(P1_U3346) );
  OAI222_X1 U7754 ( .A1(n7046), .A2(n6120), .B1(n7062), .B2(P2_U3151), .C1(
        n6119), .C2(n8951), .ZN(P2_U3286) );
  INV_X1 U7755 ( .A(n6868), .ZN(n6126) );
  OAI222_X1 U7756 ( .A1(n7046), .A2(n6126), .B1(n7163), .B2(P2_U3151), .C1(
        n6121), .C2(n8951), .ZN(P2_U3285) );
  OAI21_X1 U7757 ( .B1(n6122), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6124) );
  INV_X1 U7758 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7759 ( .A1(n6124), .A2(n6123), .ZN(n6194) );
  OR2_X1 U7760 ( .A1(n6124), .A2(n6123), .ZN(n6125) );
  INV_X1 U7761 ( .A(n9789), .ZN(n6666) );
  OAI222_X1 U7762 ( .A1(n9769), .A2(n8607), .B1(n9777), .B2(n6126), .C1(n6666), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U7763 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6132) );
  INV_X1 U7764 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6127) );
  INV_X1 U7765 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6128) );
  INV_X1 U7766 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U7767 ( .A1(n6133), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6134) );
  MUX2_X1 U7768 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6134), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n6136) );
  AND2_X1 U7769 ( .A1(n7599), .A2(n10092), .ZN(n6137) );
  NAND2_X1 U7770 ( .A1(n5549), .A2(SI_0_), .ZN(n6139) );
  INV_X1 U7771 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7772 ( .A1(n6139), .A2(n6138), .ZN(n6141) );
  AND2_X1 U7773 ( .A1(n6141), .A2(n6140), .ZN(n9780) );
  MUX2_X1 U7774 ( .A(n9779), .B(n9780), .S(n6786), .Z(n10089) );
  NAND2_X1 U7775 ( .A1(n7599), .A2(n7601), .ZN(n7604) );
  INV_X1 U7776 ( .A(n6171), .ZN(n6145) );
  NAND2_X1 U7777 ( .A1(n6145), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7778 ( .A1(n6285), .A2(n6421), .ZN(n6147) );
  AOI22_X1 U7779 ( .A1(n10089), .A2(n9121), .B1(n6145), .B2(n9779), .ZN(n6146)
         );
  NAND2_X1 U7780 ( .A1(n6147), .A2(n6146), .ZN(n6148) );
  OAI21_X1 U7781 ( .B1(n6149), .B2(n6148), .A(n6275), .ZN(n6325) );
  NOR2_X1 U7782 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .ZN(
        n6153) );
  NOR4_X1 U7783 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6152) );
  NOR4_X1 U7784 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6151) );
  NOR4_X1 U7785 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6150) );
  NAND4_X1 U7786 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n6159)
         );
  NOR4_X1 U7787 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6157) );
  NOR4_X1 U7788 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6156) );
  NOR4_X1 U7789 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6155) );
  NOR4_X1 U7790 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6154) );
  NAND4_X1 U7791 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(n6158)
         );
  NOR2_X1 U7792 ( .A1(n6159), .A2(n6158), .ZN(n6501) );
  INV_X1 U7793 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6161) );
  AOI21_X1 U7794 ( .B1(n6164), .B2(n6163), .A(n6162), .ZN(n9680) );
  OAI211_X1 U7795 ( .C1(n6501), .C2(n6165), .A(n9681), .B(n9680), .ZN(n6189)
         );
  INV_X1 U7796 ( .A(n6166), .ZN(n10088) );
  AND2_X1 U7797 ( .A1(n10194), .A2(n6510), .ZN(n6168) );
  NAND2_X1 U7798 ( .A1(n6168), .A2(n6502), .ZN(n6167) );
  INV_X1 U7799 ( .A(n6168), .ZN(n6169) );
  NAND2_X1 U7800 ( .A1(n10088), .A2(n7601), .ZN(n6187) );
  NAND2_X1 U7801 ( .A1(n6169), .A2(n6187), .ZN(n6170) );
  NAND2_X1 U7802 ( .A1(n6189), .A2(n6170), .ZN(n6172) );
  NAND2_X1 U7803 ( .A1(n7485), .A2(n6509), .ZN(n6503) );
  NAND3_X1 U7804 ( .A1(n6172), .A2(n6171), .A3(n6503), .ZN(n6173) );
  NAND2_X1 U7805 ( .A1(n6173), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6176) );
  INV_X1 U7806 ( .A(n6509), .ZN(n7657) );
  AND2_X1 U7807 ( .A1(n6502), .A2(n7657), .ZN(n6186) );
  AOI21_X1 U7808 ( .B1(n6189), .B2(n6186), .A(n6174), .ZN(n6175) );
  NAND2_X1 U7809 ( .A1(n9264), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6322) );
  INV_X1 U7810 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6289) );
  INV_X1 U7811 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6179) );
  INV_X1 U7812 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6177) );
  OR2_X1 U7813 ( .A1(n6281), .A2(n6177), .ZN(n6178) );
  OAI21_X1 U7814 ( .B1(n6180), .B2(n6179), .A(n6178), .ZN(n6181) );
  INV_X1 U7815 ( .A(n6181), .ZN(n6184) );
  INV_X1 U7816 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7817 ( .A1(n9774), .A2(n7485), .ZN(n9406) );
  NAND2_X1 U7818 ( .A1(n9283), .A2(n9250), .ZN(n10114) );
  INV_X1 U7819 ( .A(n6186), .ZN(n7664) );
  NAND2_X1 U7820 ( .A1(n10023), .A2(n6502), .ZN(n6188) );
  OR2_X1 U7821 ( .A1(n6189), .A2(n6188), .ZN(n6191) );
  INV_X1 U7822 ( .A(n10089), .ZN(n10082) );
  OAI22_X1 U7823 ( .A1(n10114), .A2(n9222), .B1(n9258), .B2(n10082), .ZN(n6192) );
  AOI21_X1 U7824 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6322), .A(n6192), .ZN(
        n6193) );
  OAI21_X1 U7825 ( .B1(n6325), .B2(n9268), .A(n6193), .ZN(P1_U3232) );
  INV_X1 U7826 ( .A(n7005), .ZN(n6212) );
  NAND2_X1 U7827 ( .A1(n6194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6195) );
  AOI22_X1 U7828 ( .A1(n9895), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n6686), .ZN(n6196) );
  OAI21_X1 U7829 ( .B1(n6212), .B2(n9773), .A(n6196), .ZN(P1_U3344) );
  INV_X1 U7830 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n8569) );
  NOR2_X1 U7831 ( .A1(n6197), .A2(n8569), .ZN(P2_U3245) );
  INV_X1 U7832 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n8616) );
  NOR2_X1 U7833 ( .A1(n6197), .A2(n8616), .ZN(P2_U3263) );
  INV_X1 U7834 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6198) );
  NOR2_X1 U7835 ( .A1(n6197), .A2(n6198), .ZN(P2_U3237) );
  INV_X1 U7836 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6199) );
  NOR2_X1 U7837 ( .A1(n6197), .A2(n6199), .ZN(P2_U3259) );
  INV_X1 U7838 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6200) );
  NOR2_X1 U7839 ( .A1(n6197), .A2(n6200), .ZN(P2_U3238) );
  INV_X1 U7840 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n8604) );
  NOR2_X1 U7841 ( .A1(n6197), .A2(n8604), .ZN(P2_U3243) );
  INV_X1 U7842 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n8646) );
  NOR2_X1 U7843 ( .A1(n6197), .A2(n8646), .ZN(P2_U3262) );
  INV_X1 U7844 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n8588) );
  NOR2_X1 U7845 ( .A1(n6197), .A2(n8588), .ZN(P2_U3261) );
  INV_X1 U7846 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6201) );
  NOR2_X1 U7847 ( .A1(n6197), .A2(n6201), .ZN(P2_U3240) );
  INV_X1 U7848 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6202) );
  NOR2_X1 U7849 ( .A1(n6197), .A2(n6202), .ZN(P2_U3234) );
  INV_X1 U7850 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n6203) );
  NOR2_X1 U7851 ( .A1(n6197), .A2(n6203), .ZN(P2_U3244) );
  INV_X1 U7852 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6204) );
  NOR2_X1 U7853 ( .A1(n6197), .A2(n6204), .ZN(P2_U3241) );
  INV_X1 U7854 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6205) );
  NOR2_X1 U7855 ( .A1(n6197), .A2(n6205), .ZN(P2_U3260) );
  INV_X1 U7856 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6206) );
  NOR2_X1 U7857 ( .A1(n6197), .A2(n6206), .ZN(P2_U3235) );
  INV_X1 U7858 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6207) );
  NOR2_X1 U7859 ( .A1(n6197), .A2(n6207), .ZN(P2_U3258) );
  INV_X1 U7860 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n6208) );
  NOR2_X1 U7861 ( .A1(n6197), .A2(n6208), .ZN(P2_U3239) );
  INV_X1 U7862 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6209) );
  NOR2_X1 U7863 ( .A1(n6197), .A2(n6209), .ZN(P2_U3242) );
  INV_X1 U7864 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6210) );
  NOR2_X1 U7865 ( .A1(n6197), .A2(n6210), .ZN(P2_U3236) );
  OAI222_X1 U7866 ( .A1(n4671), .A2(P2_U3151), .B1(n7046), .B2(n6212), .C1(
        n8951), .C2(n6211), .ZN(P2_U3284) );
  INV_X1 U7867 ( .A(n6992), .ZN(n6221) );
  INV_X1 U7868 ( .A(n8149), .ZN(n7233) );
  INV_X1 U7869 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6213) );
  OAI222_X1 U7870 ( .A1(n7046), .A2(n6221), .B1(n7233), .B2(P2_U3151), .C1(
        n6213), .C2(n8951), .ZN(P2_U3283) );
  INV_X1 U7871 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6222) );
  OR2_X1 U7872 ( .A1(n6215), .A2(n6214), .ZN(n6217) );
  NAND2_X1 U7873 ( .A1(n6217), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6216) );
  MUX2_X1 U7874 ( .A(n6216), .B(P1_IR_REG_31__SCAN_IN), .S(n6218), .Z(n6220)
         );
  INV_X1 U7875 ( .A(n6217), .ZN(n6219) );
  NAND2_X1 U7876 ( .A1(n6219), .A2(n6218), .ZN(n6343) );
  NAND2_X1 U7877 ( .A1(n6220), .A2(n6343), .ZN(n6677) );
  OAI222_X1 U7878 ( .A1(n9769), .A2(n6222), .B1(n9777), .B2(n6221), .C1(n6677), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U7879 ( .A(n6849), .ZN(n6255) );
  NAND2_X1 U7880 ( .A1(n6224), .A2(n6223), .ZN(n9885) );
  INV_X1 U7881 ( .A(n9404), .ZN(n9875) );
  INV_X1 U7882 ( .A(n6692), .ZN(n9345) );
  INV_X1 U7883 ( .A(n6614), .ZN(n9331) );
  INV_X1 U7884 ( .A(n9312), .ZN(n6239) );
  MUX2_X1 U7885 ( .A(n6182), .B(P1_REG1_REG_1__SCAN_IN), .S(n6267), .Z(n9290)
         );
  AND2_X1 U7886 ( .A1(n9779), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U7887 ( .A1(n9290), .A2(n9289), .ZN(n9288) );
  INV_X1 U7888 ( .A(n6267), .ZN(n9291) );
  NAND2_X1 U7889 ( .A1(n9291), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7890 ( .A1(n9288), .A2(n6226), .ZN(n6331) );
  INV_X1 U7891 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10204) );
  MUX2_X1 U7892 ( .A(n10204), .B(P1_REG1_REG_2__SCAN_IN), .S(n6310), .Z(n6332)
         );
  NAND2_X1 U7893 ( .A1(n6331), .A2(n6332), .ZN(n6330) );
  INV_X1 U7894 ( .A(n6310), .ZN(n6336) );
  NAND2_X1 U7895 ( .A1(n6336), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7896 ( .A1(n6330), .A2(n6227), .ZN(n9302) );
  XNOR2_X1 U7897 ( .A(n9296), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U7898 ( .A1(n9302), .A2(n9303), .ZN(n9301) );
  INV_X1 U7899 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6315) );
  OR2_X1 U7900 ( .A1(n9296), .A2(n6315), .ZN(n6228) );
  NAND2_X1 U7901 ( .A1(n9301), .A2(n6228), .ZN(n9318) );
  INV_X1 U7902 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10207) );
  MUX2_X1 U7903 ( .A(n10207), .B(P1_REG1_REG_4__SCAN_IN), .S(n9312), .Z(n9319)
         );
  NAND2_X1 U7904 ( .A1(n9318), .A2(n9319), .ZN(n9317) );
  INV_X1 U7905 ( .A(n9317), .ZN(n6229) );
  XNOR2_X1 U7906 ( .A(n9331), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9325) );
  NOR2_X1 U7907 ( .A1(n9326), .A2(n9325), .ZN(n9324) );
  INV_X1 U7908 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6636) );
  MUX2_X1 U7909 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6636), .S(n6692), .Z(n9339)
         );
  NOR2_X1 U7910 ( .A1(n9340), .A2(n9339), .ZN(n9338) );
  NAND2_X1 U7911 ( .A1(n9802), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6230) );
  OAI21_X1 U7912 ( .B1(n9802), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6230), .ZN(
        n9798) );
  NOR2_X1 U7913 ( .A1(n9799), .A2(n9798), .ZN(n9797) );
  NAND2_X1 U7914 ( .A1(n9814), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6231) );
  OAI21_X1 U7915 ( .B1(n9814), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6231), .ZN(
        n9810) );
  NOR2_X1 U7916 ( .A1(n9811), .A2(n9810), .ZN(n9809) );
  INV_X1 U7917 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6857) );
  MUX2_X1 U7918 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6857), .S(n6849), .Z(n6232)
         );
  NAND2_X1 U7919 ( .A1(n6232), .A2(n6233), .ZN(n6672) );
  OAI21_X1 U7920 ( .B1(n6233), .B2(n6232), .A(n6672), .ZN(n6251) );
  OR2_X1 U7921 ( .A1(n9774), .A2(n9404), .ZN(n6234) );
  OR2_X1 U7922 ( .A1(n9885), .A2(n6234), .ZN(n9930) );
  INV_X1 U7923 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n8639) );
  MUX2_X1 U7924 ( .A(n8639), .B(P1_REG2_REG_3__SCAN_IN), .S(n9296), .Z(n9306)
         );
  MUX2_X1 U7925 ( .A(n6179), .B(P1_REG2_REG_1__SCAN_IN), .S(n6267), .Z(n9287)
         );
  NAND2_X1 U7926 ( .A1(n9779), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6327) );
  INV_X1 U7927 ( .A(n6327), .ZN(n9286) );
  NAND2_X1 U7928 ( .A1(n9287), .A2(n9286), .ZN(n9285) );
  NAND2_X1 U7929 ( .A1(n9291), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U7930 ( .A1(n9285), .A2(n6235), .ZN(n6334) );
  INV_X1 U7931 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6654) );
  MUX2_X1 U7932 ( .A(n6654), .B(P1_REG2_REG_2__SCAN_IN), .S(n6310), .Z(n6335)
         );
  NAND2_X1 U7933 ( .A1(n6334), .A2(n6335), .ZN(n6333) );
  NAND2_X1 U7934 ( .A1(n6336), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7935 ( .A1(n6333), .A2(n6236), .ZN(n9305) );
  NAND2_X1 U7936 ( .A1(n9306), .A2(n9305), .ZN(n9304) );
  OR2_X1 U7937 ( .A1(n9296), .A2(n8639), .ZN(n6237) );
  NAND2_X1 U7938 ( .A1(n9304), .A2(n6237), .ZN(n9315) );
  INV_X1 U7939 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6238) );
  MUX2_X1 U7940 ( .A(n6238), .B(P1_REG2_REG_4__SCAN_IN), .S(n9312), .Z(n9316)
         );
  NAND2_X1 U7941 ( .A1(n9315), .A2(n9316), .ZN(n9314) );
  NAND2_X1 U7942 ( .A1(n6239), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7943 ( .A1(n9314), .A2(n6240), .ZN(n9333) );
  INV_X1 U7944 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n8695) );
  MUX2_X1 U7945 ( .A(n8695), .B(P1_REG2_REG_5__SCAN_IN), .S(n6614), .Z(n9334)
         );
  NAND2_X1 U7946 ( .A1(n9333), .A2(n9334), .ZN(n9332) );
  NAND2_X1 U7947 ( .A1(n9331), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7948 ( .A1(n9332), .A2(n6241), .ZN(n9347) );
  INV_X1 U7949 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6242) );
  MUX2_X1 U7950 ( .A(n6242), .B(P1_REG2_REG_6__SCAN_IN), .S(n6692), .Z(n9348)
         );
  NAND2_X1 U7951 ( .A1(n9347), .A2(n9348), .ZN(n9346) );
  OR2_X1 U7952 ( .A1(n6692), .A2(n6242), .ZN(n6243) );
  NAND2_X1 U7953 ( .A1(n9346), .A2(n6243), .ZN(n9793) );
  OR2_X1 U7954 ( .A1(n9802), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7955 ( .A1(n9802), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7956 ( .A1(n6245), .A2(n6244), .ZN(n9795) );
  INV_X1 U7957 ( .A(n9795), .ZN(n6246) );
  AND2_X1 U7958 ( .A1(n9793), .A2(n6246), .ZN(n9794) );
  NAND2_X1 U7959 ( .A1(n9814), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6247) );
  OAI21_X1 U7960 ( .B1(n9814), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6247), .ZN(
        n9807) );
  NOR2_X1 U7961 ( .A1(n9808), .A2(n9807), .ZN(n9806) );
  INV_X1 U7962 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6855) );
  MUX2_X1 U7963 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n6855), .S(n6849), .Z(n6248)
         );
  NAND2_X1 U7964 ( .A1(n6248), .A2(n6249), .ZN(n6667) );
  OAI21_X1 U7965 ( .B1(n6249), .B2(n6248), .A(n6667), .ZN(n6250) );
  AOI22_X1 U7966 ( .A1(n9948), .A2(n6251), .B1(n9961), .B2(n6250), .ZN(n6254)
         );
  NAND2_X1 U7967 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7114) );
  INV_X1 U7968 ( .A(n7114), .ZN(n6252) );
  AOI21_X1 U7969 ( .B1(n9883), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n6252), .ZN(
        n6253) );
  OAI211_X1 U7970 ( .C1(n6255), .C2(n9952), .A(n6254), .B(n6253), .ZN(P1_U3252) );
  INV_X1 U7971 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6263) );
  NOR2_X1 U7972 ( .A1(n6256), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6257) );
  OAI22_X1 U7973 ( .A1(n8309), .A2(n6259), .B1(n6258), .B2(n6257), .ZN(n6260)
         );
  OAI21_X1 U7974 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n5234), .A(n6260), .ZN(n6261) );
  AOI21_X1 U7975 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n8297), .A(n6261), .ZN(n6262) );
  OAI21_X1 U7976 ( .B1(n8300), .B2(n6263), .A(n6262), .ZN(P2_U3182) );
  INV_X1 U7977 ( .A(n6322), .ZN(n6290) );
  NAND2_X1 U7978 ( .A1(n9283), .A2(n9121), .ZN(n6270) );
  OR2_X1 U7979 ( .A1(n6847), .A2(n6264), .ZN(n6265) );
  NAND2_X1 U7980 ( .A1(n4440), .A2(n6268), .ZN(n6269) );
  NAND2_X1 U7981 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  XNOR2_X1 U7982 ( .A(n6271), .B(n9075), .ZN(n6303) );
  AND2_X1 U7983 ( .A1(n4440), .A2(n9121), .ZN(n6272) );
  AOI21_X1 U7984 ( .B1(n9283), .B2(n6421), .A(n6272), .ZN(n6304) );
  XNOR2_X1 U7985 ( .A(n6303), .B(n6304), .ZN(n6277) );
  NAND2_X1 U7986 ( .A1(n6273), .A2(n9125), .ZN(n6274) );
  OAI21_X1 U7987 ( .B1(n6277), .B2(n6276), .A(n6307), .ZN(n6278) );
  NAND2_X1 U7988 ( .A1(n6278), .A2(n9247), .ZN(n6288) );
  INV_X1 U7989 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6653) );
  OR2_X1 U7990 ( .A1(n7445), .A2(n10204), .ZN(n6279) );
  OAI21_X1 U7991 ( .B1(n7319), .B2(n6653), .A(n6279), .ZN(n6284) );
  INV_X1 U7992 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6280) );
  OR2_X1 U7993 ( .A1(n6281), .A2(n6280), .ZN(n6282) );
  OAI21_X1 U7994 ( .B1(n7448), .B2(n6654), .A(n6282), .ZN(n6283) );
  OR2_X2 U7995 ( .A1(n6284), .A2(n6283), .ZN(n9282) );
  INV_X1 U7996 ( .A(n9282), .ZN(n6519) );
  INV_X1 U7997 ( .A(n6285), .ZN(n6498) );
  OAI22_X1 U7998 ( .A1(n6519), .A2(n9406), .B1(n6498), .B2(n9475), .ZN(n10075)
         );
  AOI22_X1 U7999 ( .A1(n10075), .A2(n9262), .B1(n4440), .B2(n9266), .ZN(n6287)
         );
  OAI211_X1 U8000 ( .C1(n6290), .C2(n6289), .A(n6288), .B(n6287), .ZN(P1_U3222) );
  NOR2_X1 U8001 ( .A1(n7895), .A2(P2_U3151), .ZN(n6366) );
  OAI22_X1 U8002 ( .A1(n6581), .A2(n7853), .B1(n7893), .B2(n8134), .ZN(n6291)
         );
  AOI21_X1 U8003 ( .B1(n6586), .B2(n7883), .A(n6291), .ZN(n6296) );
  OAI21_X1 U8004 ( .B1(n5051), .B2(n6293), .A(n6292), .ZN(n6294) );
  NAND2_X1 U8005 ( .A1(n6294), .A2(n7871), .ZN(n6295) );
  OAI211_X1 U8006 ( .C1(n6366), .C2(n6297), .A(n6296), .B(n6295), .ZN(P2_U3162) );
  INV_X1 U8007 ( .A(n5884), .ZN(n6300) );
  INV_X1 U8008 ( .A(n6298), .ZN(n6372) );
  NAND2_X1 U8009 ( .A1(n8136), .A2(n6372), .ZN(n7968) );
  INV_X1 U8010 ( .A(n7968), .ZN(n6299) );
  NOR2_X1 U8011 ( .A1(n6300), .A2(n6299), .ZN(n7928) );
  INV_X1 U8012 ( .A(n7928), .ZN(n6368) );
  INV_X1 U8013 ( .A(n7883), .ZN(n7898) );
  OAI22_X1 U8014 ( .A1(n7898), .A2(n6372), .B1(n6532), .B2(n7893), .ZN(n6301)
         );
  AOI21_X1 U8015 ( .B1(n6368), .B2(n7871), .A(n6301), .ZN(n6302) );
  OAI21_X1 U8016 ( .B1(n6366), .B2(n5234), .A(n6302), .ZN(P2_U3172) );
  INV_X1 U8017 ( .A(n6303), .ZN(n6305) );
  NAND2_X1 U8018 ( .A1(n6305), .A2(n6304), .ZN(n6306) );
  NAND2_X1 U8019 ( .A1(n6307), .A2(n6306), .ZN(n6424) );
  NAND2_X1 U8020 ( .A1(n9282), .A2(n9121), .ZN(n6312) );
  NAND2_X1 U8021 ( .A1(n6656), .A2(n6268), .ZN(n6311) );
  NAND2_X1 U8022 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  XNOR2_X1 U8023 ( .A(n6313), .B(n9075), .ZN(n6425) );
  AND2_X1 U8024 ( .A1(n6656), .A2(n9121), .ZN(n6314) );
  AOI21_X1 U8025 ( .B1(n9282), .B2(n6421), .A(n6314), .ZN(n6426) );
  XNOR2_X1 U8026 ( .A(n6425), .B(n6426), .ZN(n6423) );
  XOR2_X1 U8027 ( .A(n6424), .B(n6423), .Z(n6324) );
  OR2_X1 U8028 ( .A1(n7445), .A2(n6315), .ZN(n6316) );
  OAI21_X1 U8029 ( .B1(n7448), .B2(n8639), .A(n6316), .ZN(n6320) );
  INV_X1 U8030 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6317) );
  OR2_X1 U8031 ( .A1(n4431), .A2(n6317), .ZN(n6318) );
  OAI21_X1 U8032 ( .B1(n7319), .B2(P1_REG3_REG_3__SCAN_IN), .A(n6318), .ZN(
        n6319) );
  OR2_X2 U8033 ( .A1(n6320), .A2(n6319), .ZN(n9281) );
  AOI22_X1 U8034 ( .A1(n9250), .A2(n9281), .B1(n9283), .B2(n9251), .ZN(n6647)
         );
  OAI22_X1 U8035 ( .A1(n6647), .A2(n9222), .B1(n10124), .B2(n9258), .ZN(n6321)
         );
  AOI21_X1 U8036 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6322), .A(n6321), .ZN(
        n6323) );
  OAI21_X1 U8037 ( .B1(n6324), .B2(n9268), .A(n6323), .ZN(P1_U3237) );
  INV_X1 U8038 ( .A(n6325), .ZN(n6326) );
  MUX2_X1 U8039 ( .A(n6327), .B(n6326), .S(n9404), .Z(n6329) );
  NOR2_X1 U8040 ( .A1(n9404), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6328) );
  OR2_X1 U8041 ( .A1(n9774), .A2(n6328), .ZN(n9876) );
  INV_X1 U8042 ( .A(n9779), .ZN(n9878) );
  NAND2_X1 U8043 ( .A1(n9876), .A2(n9878), .ZN(n9881) );
  OAI211_X1 U8044 ( .C1(n6329), .C2(n9774), .A(P1_U3973), .B(n9881), .ZN(n9323) );
  INV_X1 U8045 ( .A(n9323), .ZN(n6342) );
  OAI211_X1 U8046 ( .C1(n6332), .C2(n6331), .A(n9948), .B(n6330), .ZN(n6340)
         );
  OAI211_X1 U8047 ( .C1(n6335), .C2(n6334), .A(n9961), .B(n6333), .ZN(n6339)
         );
  AOI22_X1 U8048 ( .A1(n9883), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6338) );
  INV_X1 U8049 ( .A(n9952), .ZN(n9969) );
  NAND2_X1 U8050 ( .A1(n9969), .A2(n6336), .ZN(n6337) );
  NAND4_X1 U8051 ( .A1(n6340), .A2(n6339), .A3(n6338), .A4(n6337), .ZN(n6341)
         );
  OR2_X1 U8052 ( .A1(n6342), .A2(n6341), .ZN(P1_U3245) );
  INV_X1 U8053 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6349) );
  INV_X1 U8054 ( .A(n7273), .ZN(n6351) );
  NAND2_X1 U8055 ( .A1(n6343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6344) );
  MUX2_X1 U8056 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6344), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n6348) );
  INV_X1 U8057 ( .A(n6346), .ZN(n6347) );
  INV_X1 U8058 ( .A(n9907), .ZN(n9355) );
  OAI222_X1 U8059 ( .A1(n9769), .A2(n6349), .B1(n9777), .B2(n6351), .C1(
        P1_U3086), .C2(n9355), .ZN(P1_U3342) );
  INV_X1 U8060 ( .A(n8174), .ZN(n8164) );
  OAI222_X1 U8061 ( .A1(n8164), .A2(P2_U3151), .B1(n7046), .B2(n6351), .C1(
        n8951), .C2(n6350), .ZN(P2_U3282) );
  OAI21_X1 U8062 ( .B1(n8461), .B2(n10274), .A(n6368), .ZN(n6352) );
  NAND2_X1 U8063 ( .A1(n5248), .A2(n8463), .ZN(n6369) );
  OAI211_X1 U8064 ( .C1(n6372), .C2(n10270), .A(n6352), .B(n6369), .ZN(n6354)
         );
  NAND2_X1 U8065 ( .A1(n6354), .A2(n10289), .ZN(n6353) );
  OAI21_X1 U8066 ( .B1(n10289), .B2(n8704), .A(n6353), .ZN(P2_U3459) );
  INV_X1 U8067 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8068 ( .A1(n6354), .A2(n10275), .ZN(n6355) );
  OAI21_X1 U8069 ( .B1(n6356), .B2(n10275), .A(n6355), .ZN(P2_U3390) );
  INV_X1 U8070 ( .A(n7279), .ZN(n6413) );
  OR2_X1 U8071 ( .A1(n6346), .A2(n6492), .ZN(n6440) );
  XNOR2_X1 U8072 ( .A(n6440), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U8073 ( .A1(n9911), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n6686), .ZN(n6357) );
  OAI21_X1 U8074 ( .B1(n6413), .B2(n9773), .A(n6357), .ZN(P1_U3341) );
  INV_X1 U8075 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6365) );
  OAI21_X1 U8076 ( .B1(n6360), .B2(n6359), .A(n6358), .ZN(n6361) );
  NAND2_X1 U8077 ( .A1(n6361), .A2(n7871), .ZN(n6364) );
  OAI22_X1 U8078 ( .A1(n6532), .A2(n7853), .B1(n7893), .B2(n6591), .ZN(n6362)
         );
  AOI21_X1 U8079 ( .B1(n7973), .B2(n7883), .A(n6362), .ZN(n6363) );
  OAI211_X1 U8080 ( .C1(n6366), .C2(n6365), .A(n6364), .B(n6363), .ZN(P2_U3177) );
  NAND3_X1 U8081 ( .A1(n6368), .A2(n10270), .A3(n6367), .ZN(n6370) );
  AOI21_X1 U8082 ( .B1(n6370), .B2(n6369), .A(n8489), .ZN(n6375) );
  NOR2_X1 U8083 ( .A1(n10233), .A2(n6371), .ZN(n6374) );
  OAI22_X1 U8084 ( .A1(n8431), .A2(n6372), .B1(n5234), .B2(n8444), .ZN(n6373)
         );
  OR3_X1 U8085 ( .A1(n6375), .A2(n6374), .A3(n6373), .ZN(P2_U3233) );
  AOI211_X1 U8086 ( .C1(n6378), .C2(n6377), .A(n7070), .B(n6376), .ZN(n6394)
         );
  INV_X1 U8087 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6384) );
  OAI21_X1 U8088 ( .B1(n6381), .B2(n6380), .A(n6379), .ZN(n6382) );
  INV_X1 U8089 ( .A(n6382), .ZN(n6383) );
  OAI22_X1 U8090 ( .A1(n6384), .A2(n8300), .B1(n8306), .B2(n6383), .ZN(n6393)
         );
  OAI21_X1 U8091 ( .B1(n6387), .B2(n6386), .A(n6385), .ZN(n6389) );
  NOR2_X1 U8092 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6365), .ZN(n6388) );
  AOI21_X1 U8093 ( .B1(n8140), .B2(n6389), .A(n6388), .ZN(n6390) );
  OAI21_X1 U8094 ( .B1(n8266), .B2(n6391), .A(n6390), .ZN(n6392) );
  OR3_X1 U8095 ( .A1(n6394), .A2(n6393), .A3(n6392), .ZN(P2_U3184) );
  OAI21_X1 U8096 ( .B1(n6397), .B2(n6396), .A(n6395), .ZN(n6410) );
  INV_X1 U8097 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6408) );
  INV_X1 U8098 ( .A(n8306), .ZN(n8148) );
  OAI21_X1 U8099 ( .B1(n6399), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6398), .ZN(
        n6401) );
  AOI22_X1 U8100 ( .A1(n8148), .A2(n6401), .B1(n8297), .B2(n4657), .ZN(n6407)
         );
  OAI21_X1 U8101 ( .B1(n6403), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6402), .ZN(
        n6405) );
  AOI21_X1 U8102 ( .B1(n8140), .B2(n6405), .A(n6404), .ZN(n6406) );
  OAI211_X1 U8103 ( .C1(n6408), .C2(n8300), .A(n6407), .B(n6406), .ZN(n6409)
         );
  AOI21_X1 U8104 ( .B1(n6410), .B2(n8309), .A(n6409), .ZN(n6411) );
  INV_X1 U8105 ( .A(n6411), .ZN(P2_U3185) );
  INV_X1 U8106 ( .A(n8177), .ZN(n8193) );
  INV_X1 U8107 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6412) );
  OAI222_X1 U8108 ( .A1(n7046), .A2(n6413), .B1(n8193), .B2(P2_U3151), .C1(
        n6412), .C2(n8951), .ZN(P2_U3281) );
  NAND2_X1 U8109 ( .A1(n9281), .A2(n9121), .ZN(n6419) );
  OR2_X1 U8110 ( .A1(n6847), .A2(n6414), .ZN(n6417) );
  OR2_X1 U8111 ( .A1(n7439), .A2(n6415), .ZN(n6416) );
  OAI211_X1 U8112 ( .C1(n6786), .C2(n9296), .A(n6417), .B(n6416), .ZN(n10060)
         );
  NAND2_X1 U8113 ( .A1(n10060), .A2(n6268), .ZN(n6418) );
  NAND2_X1 U8114 ( .A1(n6419), .A2(n6418), .ZN(n6420) );
  XNOR2_X1 U8115 ( .A(n6420), .B(n9075), .ZN(n6460) );
  AND2_X1 U8116 ( .A1(n10060), .A2(n9121), .ZN(n6422) );
  AOI21_X1 U8117 ( .B1(n9281), .B2(n6421), .A(n6422), .ZN(n6461) );
  XNOR2_X1 U8118 ( .A(n6460), .B(n6461), .ZN(n6458) );
  NAND2_X1 U8119 ( .A1(n6424), .A2(n6423), .ZN(n6429) );
  INV_X1 U8120 ( .A(n6425), .ZN(n6427) );
  NAND2_X1 U8121 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  XOR2_X1 U8122 ( .A(n6458), .B(n6459), .Z(n6437) );
  XNOR2_X1 U8123 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6513) );
  OR2_X1 U8124 ( .A1(n7319), .A2(n6513), .ZN(n6434) );
  OR2_X1 U8125 ( .A1(n7448), .A2(n6238), .ZN(n6433) );
  INV_X1 U8126 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6430) );
  OR2_X1 U8127 ( .A1(n4431), .A2(n6430), .ZN(n6432) );
  OR2_X1 U8128 ( .A1(n7445), .A2(n10207), .ZN(n6431) );
  NAND4_X1 U8129 ( .A1(n6434), .A2(n6433), .A3(n6432), .A4(n6431), .ZN(n9280)
         );
  INV_X1 U8130 ( .A(n9280), .ZN(n6694) );
  OAI22_X1 U8131 ( .A1(n6519), .A2(n9475), .B1(n6694), .B2(n9406), .ZN(n10056)
         );
  AOI22_X1 U8132 ( .A1(n10056), .A2(n9262), .B1(n10060), .B2(n9266), .ZN(n6436) );
  MUX2_X1 U8133 ( .A(n9264), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6435) );
  OAI211_X1 U8134 ( .C1(n6437), .C2(n9268), .A(n6436), .B(n6435), .ZN(P1_U3218) );
  INV_X1 U8135 ( .A(n7288), .ZN(n6444) );
  AOI22_X1 U8136 ( .A1(n8218), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8939), .ZN(n6438) );
  OAI21_X1 U8137 ( .B1(n6444), .B2(n8954), .A(n6438), .ZN(P2_U3280) );
  INV_X1 U8138 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8139 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  NAND2_X1 U8140 ( .A1(n6441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6442) );
  XNOR2_X1 U8141 ( .A(n6442), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U8142 ( .A1(n9935), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n6686), .ZN(n6443) );
  OAI21_X1 U8143 ( .B1(n6444), .B2(n9773), .A(n6443), .ZN(P1_U3340) );
  NAND3_X1 U8144 ( .A1(n6446), .A2(n6455), .A3(n6447), .ZN(n6448) );
  NAND2_X1 U8145 ( .A1(n6445), .A2(n6448), .ZN(n6451) );
  NAND2_X1 U8146 ( .A1(n8132), .A2(n8463), .ZN(n6449) );
  OAI21_X1 U8147 ( .B1(n8134), .B2(n8480), .A(n6449), .ZN(n6450) );
  AOI21_X1 U8148 ( .B1(n6451), .B2(n8461), .A(n6450), .ZN(n10248) );
  OAI22_X1 U8149 ( .A1(n8431), .A2(n6452), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8444), .ZN(n6453) );
  AOI21_X1 U8150 ( .B1(n8489), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6453), .ZN(
        n6457) );
  XNOR2_X1 U8151 ( .A(n6454), .B(n6455), .ZN(n10243) );
  NAND2_X1 U8152 ( .A1(n10243), .A2(n8486), .ZN(n6456) );
  OAI211_X1 U8153 ( .C1(n10248), .C2(n8489), .A(n6457), .B(n6456), .ZN(
        P2_U3230) );
  INV_X1 U8154 ( .A(n6460), .ZN(n6462) );
  NAND2_X1 U8155 ( .A1(n9280), .A2(n9121), .ZN(n6469) );
  OR2_X1 U8156 ( .A1(n7439), .A2(n6464), .ZN(n6467) );
  OR2_X1 U8157 ( .A1(n6847), .A2(n6465), .ZN(n6466) );
  OAI211_X1 U8158 ( .C1(n6786), .C2(n9312), .A(n6467), .B(n6466), .ZN(n10135)
         );
  NAND2_X1 U8159 ( .A1(n10135), .A2(n6268), .ZN(n6468) );
  NAND2_X1 U8160 ( .A1(n6469), .A2(n6468), .ZN(n6470) );
  XNOR2_X1 U8161 ( .A(n6470), .B(n9075), .ZN(n6473) );
  NAND2_X1 U8162 ( .A1(n9280), .A2(n6421), .ZN(n6472) );
  NAND2_X1 U8163 ( .A1(n10135), .A2(n9121), .ZN(n6471) );
  NAND2_X1 U8164 ( .A1(n6472), .A2(n6471), .ZN(n6474) );
  NAND2_X1 U8165 ( .A1(n6473), .A2(n6474), .ZN(n6621) );
  INV_X1 U8166 ( .A(n6473), .ZN(n6476) );
  INV_X1 U8167 ( .A(n6474), .ZN(n6475) );
  AOI21_X1 U8168 ( .B1(n6478), .B2(n6477), .A(n9268), .ZN(n6479) );
  NAND2_X1 U8169 ( .A1(n6479), .A2(n6622), .ZN(n6491) );
  INV_X1 U8170 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6480) );
  OR2_X1 U8171 ( .A1(n7445), .A2(n6480), .ZN(n6481) );
  OAI21_X1 U8172 ( .B1(n7448), .B2(n8695), .A(n6481), .ZN(n6488) );
  INV_X1 U8173 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8174 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6482) );
  NAND2_X1 U8175 ( .A1(n6483), .A2(n6482), .ZN(n6484) );
  NAND2_X1 U8176 ( .A1(n6633), .A2(n6484), .ZN(n6632) );
  INV_X1 U8177 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6485) );
  OR2_X1 U8178 ( .A1(n4431), .A2(n6485), .ZN(n6486) );
  OAI21_X1 U8179 ( .B1(n7319), .B2(n6632), .A(n6486), .ZN(n6487) );
  AOI22_X1 U8180 ( .A1(n9250), .A2(n9279), .B1(n9281), .B2(n9251), .ZN(n6523)
         );
  NAND2_X1 U8181 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9311) );
  OAI21_X1 U8182 ( .B1(n6523), .B2(n9222), .A(n9311), .ZN(n6489) );
  AOI21_X1 U8183 ( .B1(n10135), .B2(n9266), .A(n6489), .ZN(n6490) );
  OAI211_X1 U8184 ( .C1(n9264), .C2(n6513), .A(n6491), .B(n6490), .ZN(P1_U3230) );
  INV_X1 U8185 ( .A(n7303), .ZN(n6542) );
  NOR2_X1 U8186 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  MUX2_X1 U8187 ( .A(n6492), .B(n6494), .S(P1_IR_REG_16__SCAN_IN), .Z(n6495)
         );
  INV_X1 U8188 ( .A(n6495), .ZN(n6496) );
  AND2_X1 U8189 ( .A1(n6496), .A2(n6661), .ZN(n9939) );
  AOI22_X1 U8190 ( .A1(n9939), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n6686), .ZN(n6497) );
  OAI21_X1 U8191 ( .B1(n6542), .B2(n9773), .A(n6497), .ZN(P1_U3339) );
  INV_X1 U8192 ( .A(n10135), .ZN(n6693) );
  NAND2_X1 U8193 ( .A1(n9280), .A2(n6693), .ZN(n7608) );
  NAND2_X1 U8194 ( .A1(n7496), .A2(n7608), .ZN(n7490) );
  OAI22_X1 U8195 ( .A1(n10069), .A2(n10070), .B1(n9283), .B2(n4440), .ZN(n6650) );
  INV_X1 U8196 ( .A(n9281), .ZN(n6500) );
  NAND2_X1 U8197 ( .A1(n6500), .A2(n10060), .ZN(n7492) );
  INV_X1 U8198 ( .A(n10060), .ZN(n10129) );
  NAND2_X1 U8199 ( .A1(n9281), .A2(n10129), .ZN(n7609) );
  XOR2_X1 U8200 ( .A(n7490), .B(n6695), .Z(n10138) );
  NAND2_X1 U8201 ( .A1(n6502), .A2(n6501), .ZN(n6505) );
  INV_X1 U8202 ( .A(n6503), .ZN(n6504) );
  INV_X1 U8203 ( .A(n9681), .ZN(n9741) );
  NAND3_X1 U8204 ( .A1(n9742), .A2(n9680), .A3(n9741), .ZN(n6506) );
  NAND2_X1 U8205 ( .A1(n6507), .A2(n4433), .ZN(n6508) );
  AND2_X1 U8206 ( .A1(n6508), .A2(n6509), .ZN(n6511) );
  OAI21_X1 U8207 ( .B1(n6510), .B2(n6509), .A(n6166), .ZN(n10087) );
  OR2_X1 U8208 ( .A1(n6511), .A2(n10087), .ZN(n9992) );
  NAND2_X1 U8209 ( .A1(n9992), .A2(n9660), .ZN(n10028) );
  INV_X1 U8210 ( .A(n6512), .ZN(n10063) );
  AOI211_X1 U8211 ( .C1(n10135), .C2(n10063), .A(n10012), .B(n10051), .ZN(
        n10134) );
  OAI22_X1 U8212 ( .A1(n9621), .A2(n6693), .B1(n6513), .B2(n10090), .ZN(n6514)
         );
  AOI21_X1 U8213 ( .B1(n10134), .B2(n10097), .A(n6514), .ZN(n6527) );
  NAND2_X1 U8214 ( .A1(n6515), .A2(n7464), .ZN(n6518) );
  INV_X1 U8215 ( .A(n9283), .ZN(n6516) );
  NAND2_X1 U8216 ( .A1(n6516), .A2(n4440), .ZN(n6517) );
  NAND2_X1 U8217 ( .A1(n6518), .A2(n6517), .ZN(n6646) );
  NAND2_X1 U8218 ( .A1(n6519), .A2(n6656), .ZN(n6520) );
  INV_X1 U8219 ( .A(n7492), .ZN(n6521) );
  XNOR2_X1 U8220 ( .A(n7491), .B(n7490), .ZN(n6525) );
  NAND2_X1 U8221 ( .A1(n4433), .A2(n4434), .ZN(n6522) );
  INV_X1 U8222 ( .A(n6523), .ZN(n6524) );
  AOI21_X1 U8223 ( .B1(n6525), .B2(n10112), .A(n6524), .ZN(n10137) );
  MUX2_X1 U8224 ( .A(n10137), .B(n6238), .S(n10100), .Z(n6526) );
  OAI211_X1 U8225 ( .C1(n10138), .C2(n9630), .A(n6527), .B(n6526), .ZN(
        P1_U3289) );
  XNOR2_X1 U8226 ( .A(n6528), .B(n7971), .ZN(n6544) );
  NAND2_X1 U8227 ( .A1(n6544), .A2(n6719), .ZN(n6536) );
  NAND3_X1 U8228 ( .A1(n7971), .A2(n6530), .A3(n6529), .ZN(n6531) );
  NAND2_X1 U8229 ( .A1(n6446), .A2(n6531), .ZN(n6534) );
  OAI22_X1 U8230 ( .A1(n6532), .A2(n8480), .B1(n6591), .B2(n8481), .ZN(n6533)
         );
  AOI21_X1 U8231 ( .B1(n6534), .B2(n8461), .A(n6533), .ZN(n6535) );
  AND2_X1 U8232 ( .A1(n6536), .A2(n6535), .ZN(n6547) );
  NOR2_X1 U8233 ( .A1(n6537), .A2(n10270), .ZN(n6538) );
  AOI21_X1 U8234 ( .B1(n6544), .B2(n5763), .A(n6538), .ZN(n6539) );
  AND2_X1 U8235 ( .A1(n6547), .A2(n6539), .ZN(n10241) );
  MUX2_X1 U8236 ( .A(n10241), .B(n6540), .S(n5770), .Z(n6541) );
  INV_X1 U8237 ( .A(n6541), .ZN(P2_U3461) );
  INV_X1 U8238 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6543) );
  INV_X1 U8239 ( .A(n8222), .ZN(n8237) );
  OAI222_X1 U8240 ( .A1(n8951), .A2(n6543), .B1(n7046), .B2(n6542), .C1(
        P2_U3151), .C2(n8237), .ZN(P2_U3279) );
  INV_X1 U8241 ( .A(n6544), .ZN(n6551) );
  AND2_X1 U8242 ( .A1(n10233), .A2(n6545), .ZN(n7674) );
  INV_X1 U8243 ( .A(n7674), .ZN(n6589) );
  AOI22_X1 U8244 ( .A1(n7973), .A2(n8482), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n10228), .ZN(n6546) );
  AND2_X1 U8245 ( .A1(n6547), .A2(n6546), .ZN(n6549) );
  MUX2_X1 U8246 ( .A(n6549), .B(n6548), .S(n8489), .Z(n6550) );
  OAI21_X1 U8247 ( .B1(n6551), .B2(n6589), .A(n6550), .ZN(P2_U3231) );
  AND2_X1 U8248 ( .A1(n7998), .A2(n7985), .ZN(n7980) );
  INV_X1 U8249 ( .A(n7980), .ZN(n7925) );
  XNOR2_X1 U8250 ( .A(n6552), .B(n7925), .ZN(n10252) );
  XNOR2_X1 U8251 ( .A(n6553), .B(n7925), .ZN(n6554) );
  AOI222_X1 U8252 ( .A1(n8461), .A2(n6554), .B1(n8131), .B2(n8463), .C1(n8133), 
        .C2(n8466), .ZN(n10250) );
  MUX2_X1 U8253 ( .A(n5840), .B(n10250), .S(n10233), .Z(n6556) );
  AOI22_X1 U8254 ( .A1(n10226), .A2(n6602), .B1(n10228), .B2(n6599), .ZN(n6555) );
  OAI211_X1 U8255 ( .C1(n8783), .C2(n10252), .A(n6556), .B(n6555), .ZN(
        P2_U3229) );
  INV_X1 U8256 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10295) );
  NOR2_X1 U8257 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6557) );
  AOI21_X1 U8258 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6557), .ZN(n10300) );
  NOR2_X1 U8259 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6558) );
  AOI21_X1 U8260 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6558), .ZN(n10303) );
  NOR2_X1 U8261 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6559) );
  AOI21_X1 U8262 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6559), .ZN(n10306) );
  NOR2_X1 U8263 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6560) );
  AOI21_X1 U8264 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6560), .ZN(n10309) );
  NOR2_X1 U8265 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6561) );
  AOI21_X1 U8266 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6561), .ZN(n10312) );
  NOR2_X1 U8267 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6562) );
  AOI21_X1 U8268 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6562), .ZN(n10315) );
  NOR2_X1 U8269 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6563) );
  AOI21_X1 U8270 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6563), .ZN(n10318) );
  NOR2_X1 U8271 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6564) );
  AOI21_X1 U8272 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6564), .ZN(n10321) );
  NOR2_X1 U8273 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n6565) );
  AOI21_X1 U8274 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n6565), .ZN(n10330) );
  NOR2_X1 U8275 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n6566) );
  AOI21_X1 U8276 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n6566), .ZN(n10336) );
  NOR2_X1 U8277 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6567) );
  AOI21_X1 U8278 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6567), .ZN(n10333) );
  NOR2_X1 U8279 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6568) );
  AOI21_X1 U8280 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6568), .ZN(n10324) );
  INV_X1 U8281 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6750) );
  INV_X1 U8282 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9329) );
  AOI22_X1 U8283 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .B1(n6750), .B2(n9329), .ZN(n10327) );
  INV_X1 U8284 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U8285 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n6569) );
  NAND2_X1 U8286 ( .A1(n8674), .A2(n6569), .ZN(n10292) );
  NAND3_X1 U8287 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U8288 ( .A1(n5951), .A2(n10293), .ZN(n10290) );
  NAND2_X1 U8289 ( .A1(n10292), .A2(n10290), .ZN(n10339) );
  NAND2_X1 U8290 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n6570) );
  OAI21_X1 U8291 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n6570), .ZN(n10338) );
  NOR2_X1 U8292 ( .A1(n10339), .A2(n10338), .ZN(n10337) );
  AOI21_X1 U8293 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10337), .ZN(n10342) );
  NAND2_X1 U8294 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6571) );
  OAI21_X1 U8295 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6571), .ZN(n10341) );
  NOR2_X1 U8296 ( .A1(n10342), .A2(n10341), .ZN(n10340) );
  AOI21_X1 U8297 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10340), .ZN(n10345) );
  NOR2_X1 U8298 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n6572) );
  AOI21_X1 U8299 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n6572), .ZN(n10344) );
  NAND2_X1 U8300 ( .A1(n10345), .A2(n10344), .ZN(n10343) );
  OAI21_X1 U8301 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10343), .ZN(n10326) );
  NAND2_X1 U8302 ( .A1(n10327), .A2(n10326), .ZN(n10325) );
  OAI21_X1 U8303 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10325), .ZN(n10323) );
  NAND2_X1 U8304 ( .A1(n10324), .A2(n10323), .ZN(n10322) );
  OAI21_X1 U8305 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10322), .ZN(n10332) );
  NAND2_X1 U8306 ( .A1(n10333), .A2(n10332), .ZN(n10331) );
  OAI21_X1 U8307 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10331), .ZN(n10335) );
  NAND2_X1 U8308 ( .A1(n10336), .A2(n10335), .ZN(n10334) );
  OAI21_X1 U8309 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10334), .ZN(n10329) );
  NAND2_X1 U8310 ( .A1(n10330), .A2(n10329), .ZN(n10328) );
  OAI21_X1 U8311 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10328), .ZN(n10320) );
  NAND2_X1 U8312 ( .A1(n10321), .A2(n10320), .ZN(n10319) );
  OAI21_X1 U8313 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10319), .ZN(n10317) );
  NAND2_X1 U8314 ( .A1(n10318), .A2(n10317), .ZN(n10316) );
  OAI21_X1 U8315 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10316), .ZN(n10314) );
  NAND2_X1 U8316 ( .A1(n10315), .A2(n10314), .ZN(n10313) );
  OAI21_X1 U8317 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10313), .ZN(n10311) );
  NAND2_X1 U8318 ( .A1(n10312), .A2(n10311), .ZN(n10310) );
  OAI21_X1 U8319 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10310), .ZN(n10308) );
  NAND2_X1 U8320 ( .A1(n10309), .A2(n10308), .ZN(n10307) );
  OAI21_X1 U8321 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10307), .ZN(n10305) );
  NAND2_X1 U8322 ( .A1(n10306), .A2(n10305), .ZN(n10304) );
  OAI21_X1 U8323 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10304), .ZN(n10302) );
  NAND2_X1 U8324 ( .A1(n10303), .A2(n10302), .ZN(n10301) );
  OAI21_X1 U8325 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10301), .ZN(n10299) );
  NAND2_X1 U8326 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  OAI21_X1 U8327 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10298), .ZN(n10296) );
  NAND2_X1 U8328 ( .A1(n10295), .A2(n10296), .ZN(n6573) );
  NOR2_X1 U8329 ( .A1(n10295), .A2(n10296), .ZN(n10294) );
  AOI21_X1 U8330 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n6573), .A(n10294), .ZN(
        n6577) );
  NOR2_X1 U8331 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  XNOR2_X1 U8332 ( .A(n6577), .B(n6576), .ZN(ADD_1068_U4) );
  INV_X1 U8333 ( .A(n6578), .ZN(n6579) );
  AOI21_X1 U8334 ( .B1(n5884), .B2(n5686), .A(n6579), .ZN(n10237) );
  OAI21_X1 U8335 ( .B1(n6580), .B2(n5686), .A(n6529), .ZN(n6585) );
  OAI22_X1 U8336 ( .A1(n6581), .A2(n8480), .B1(n8134), .B2(n8481), .ZN(n6584)
         );
  INV_X1 U8337 ( .A(n6719), .ZN(n6582) );
  NOR2_X1 U8338 ( .A1(n10237), .A2(n6582), .ZN(n6583) );
  AOI211_X1 U8339 ( .C1(n8461), .C2(n6585), .A(n6584), .B(n6583), .ZN(n10234)
         );
  MUX2_X1 U8340 ( .A(n5949), .B(n10234), .S(n10233), .Z(n6588) );
  AOI22_X1 U8341 ( .A1(n10226), .A2(n6586), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10228), .ZN(n6587) );
  OAI211_X1 U8342 ( .C1(n10237), .C2(n6589), .A(n6588), .B(n6587), .ZN(
        P2_U3232) );
  OR2_X1 U8343 ( .A1(n6591), .A2(n6590), .ZN(n6592) );
  XNOR2_X1 U8344 ( .A(n6602), .B(n7778), .ZN(n6594) );
  NAND2_X1 U8345 ( .A1(n6760), .A2(n6594), .ZN(n6766) );
  INV_X1 U8346 ( .A(n6594), .ZN(n6595) );
  NAND2_X1 U8347 ( .A1(n6595), .A2(n8132), .ZN(n6596) );
  OAI21_X1 U8348 ( .B1(n6598), .B2(n6597), .A(n6764), .ZN(n6608) );
  NAND2_X1 U8349 ( .A1(n7895), .A2(n6599), .ZN(n6606) );
  INV_X1 U8350 ( .A(n6600), .ZN(n6601) );
  AOI21_X1 U8351 ( .B1(n7850), .B2(n8131), .A(n6601), .ZN(n6605) );
  NAND2_X1 U8352 ( .A1(n7883), .A2(n6602), .ZN(n6604) );
  NAND2_X1 U8353 ( .A1(n7891), .A2(n8133), .ZN(n6603) );
  NAND4_X1 U8354 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n6607)
         );
  AOI21_X1 U8355 ( .B1(n6608), .B2(n7871), .A(n6607), .ZN(n6609) );
  INV_X1 U8356 ( .A(n6609), .ZN(P2_U3170) );
  NAND2_X1 U8357 ( .A1(n9279), .A2(n9121), .ZN(n6616) );
  OR2_X1 U8358 ( .A1(n6847), .A2(n6610), .ZN(n6613) );
  OR2_X1 U8359 ( .A1(n7439), .A2(n6611), .ZN(n6612) );
  OAI211_X1 U8360 ( .C1(n6786), .C2(n6614), .A(n6613), .B(n6612), .ZN(n10047)
         );
  NAND2_X1 U8361 ( .A1(n10047), .A2(n9127), .ZN(n6615) );
  NAND2_X1 U8362 ( .A1(n6616), .A2(n6615), .ZN(n6617) );
  XNOR2_X1 U8363 ( .A(n6617), .B(n9125), .ZN(n6623) );
  AND2_X1 U8364 ( .A1(n6621), .A2(n6623), .ZN(n6618) );
  NAND2_X1 U8365 ( .A1(n9279), .A2(n6421), .ZN(n6620) );
  NAND2_X1 U8366 ( .A1(n10047), .A2(n9121), .ZN(n6619) );
  NAND2_X1 U8367 ( .A1(n6620), .A2(n6619), .ZN(n6629) );
  NAND2_X1 U8368 ( .A1(n6631), .A2(n6629), .ZN(n6626) );
  NAND2_X1 U8369 ( .A1(n6622), .A2(n6621), .ZN(n6625) );
  INV_X1 U8370 ( .A(n6623), .ZN(n6624) );
  INV_X1 U8371 ( .A(n6626), .ZN(n6628) );
  NAND2_X1 U8372 ( .A1(n6628), .A2(n6627), .ZN(n6630) );
  AOI22_X1 U8373 ( .A1(n6734), .A2(n6631), .B1(n6630), .B2(n6629), .ZN(n6644)
         );
  INV_X1 U8374 ( .A(n6632), .ZN(n10046) );
  INV_X1 U8375 ( .A(n9264), .ZN(n9210) );
  INV_X1 U8376 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U8377 ( .A1(n6633), .A2(n8643), .ZN(n6634) );
  NAND2_X1 U8378 ( .A1(n6702), .A2(n6634), .ZN(n6738) );
  OR2_X1 U8379 ( .A1(n7430), .A2(n6738), .ZN(n6640) );
  OR2_X1 U8380 ( .A1(n7448), .A2(n6242), .ZN(n6639) );
  INV_X1 U8381 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6635) );
  OR2_X1 U8382 ( .A1(n4431), .A2(n6635), .ZN(n6638) );
  OR2_X1 U8383 ( .A1(n7445), .A2(n6636), .ZN(n6637) );
  NAND4_X1 U8384 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n9278)
         );
  INV_X1 U8385 ( .A(n9278), .ZN(n6883) );
  OAI22_X1 U8386 ( .A1(n6694), .A2(n9475), .B1(n6883), .B2(n9406), .ZN(n10044)
         );
  AOI22_X1 U8387 ( .A1(n10044), .A2(n9262), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n6641) );
  OAI21_X1 U8388 ( .B1(n10141), .B2(n9258), .A(n6641), .ZN(n6642) );
  AOI21_X1 U8389 ( .B1(n10046), .B2(n9210), .A(n6642), .ZN(n6643) );
  OAI21_X1 U8390 ( .B1(n6644), .B2(n9268), .A(n6643), .ZN(P1_U3227) );
  INV_X1 U8391 ( .A(n7314), .ZN(n6663) );
  INV_X1 U8392 ( .A(n8273), .ZN(n8236) );
  INV_X1 U8393 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6645) );
  OAI222_X1 U8394 ( .A1(n7046), .A2(n6663), .B1(n8236), .B2(P2_U3151), .C1(
        n6645), .C2(n8951), .ZN(P2_U3278) );
  XNOR2_X1 U8395 ( .A(n6646), .B(n6649), .ZN(n6648) );
  OAI21_X1 U8396 ( .B1(n6648), .B2(n10072), .A(n6647), .ZN(n10125) );
  INV_X1 U8397 ( .A(n10125), .ZN(n6660) );
  XNOR2_X1 U8398 ( .A(n6650), .B(n6649), .ZN(n10127) );
  INV_X1 U8399 ( .A(n9630), .ZN(n10066) );
  INV_X1 U8400 ( .A(n10080), .ZN(n6652) );
  INV_X1 U8401 ( .A(n10064), .ZN(n6651) );
  OAI211_X1 U8402 ( .C1(n10124), .C2(n6652), .A(n6651), .B(n10081), .ZN(n10123) );
  OAI22_X1 U8403 ( .A1(n10058), .A2(n6654), .B1(n6653), .B2(n10090), .ZN(n6655) );
  AOI21_X1 U8404 ( .B1(n10077), .B2(n6656), .A(n6655), .ZN(n6657) );
  OAI21_X1 U8405 ( .B1(n10123), .B2(n9671), .A(n6657), .ZN(n6658) );
  AOI21_X1 U8406 ( .B1(n10127), .B2(n10066), .A(n6658), .ZN(n6659) );
  OAI21_X1 U8407 ( .B1(n6660), .B2(n10100), .A(n6659), .ZN(P1_U3291) );
  INV_X1 U8408 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U8409 ( .A1(n6661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6662) );
  XNOR2_X1 U8410 ( .A(n6662), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9389) );
  INV_X1 U8411 ( .A(n9389), .ZN(n9378) );
  OAI222_X1 U8412 ( .A1(n9769), .A2(n6664), .B1(n9777), .B2(n6663), .C1(n9378), 
        .C2(P1_U3086), .ZN(P1_U3338) );
  NOR2_X1 U8413 ( .A1(n9368), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6665) );
  AOI21_X1 U8414 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9368), .A(n6665), .ZN(
        n6670) );
  INV_X1 U8415 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8568) );
  AOI22_X1 U8416 ( .A1(n9789), .A2(n8568), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n6666), .ZN(n9786) );
  OAI21_X1 U8417 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6849), .A(n6667), .ZN(
        n9785) );
  NOR2_X1 U8418 ( .A1(n9786), .A2(n9785), .ZN(n9784) );
  NAND2_X1 U8419 ( .A1(n9895), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6668) );
  OAI21_X1 U8420 ( .B1(n9895), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6668), .ZN(
        n9888) );
  NOR2_X1 U8421 ( .A1(n9889), .A2(n9888), .ZN(n9887) );
  AOI21_X1 U8422 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9895), .A(n9887), .ZN(
        n6669) );
  NAND2_X1 U8423 ( .A1(n6670), .A2(n6669), .ZN(n9367) );
  OAI21_X1 U8424 ( .B1(n6670), .B2(n6669), .A(n9367), .ZN(n6671) );
  NAND2_X1 U8425 ( .A1(n6671), .A2(n9961), .ZN(n6681) );
  OAI21_X1 U8426 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n6849), .A(n6672), .ZN(
        n9782) );
  INV_X1 U8427 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6874) );
  MUX2_X1 U8428 ( .A(n6874), .B(P1_REG1_REG_10__SCAN_IN), .S(n9789), .Z(n9783)
         );
  NOR2_X1 U8429 ( .A1(n9782), .A2(n9783), .ZN(n9781) );
  MUX2_X1 U8430 ( .A(n6673), .B(P1_REG1_REG_11__SCAN_IN), .S(n9895), .Z(n9891)
         );
  NOR2_X1 U8431 ( .A1(n9892), .A2(n9891), .ZN(n9890) );
  INV_X1 U8432 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U8433 ( .A1(n9368), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n10216), .B2(
        n6677), .ZN(n6674) );
  NAND2_X1 U8434 ( .A1(n6675), .A2(n6674), .ZN(n9356) );
  OAI21_X1 U8435 ( .B1(n6675), .B2(n6674), .A(n9356), .ZN(n6679) );
  NAND2_X1 U8436 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9152) );
  NAND2_X1 U8437 ( .A1(n9883), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6676) );
  OAI211_X1 U8438 ( .C1(n9952), .C2(n6677), .A(n9152), .B(n6676), .ZN(n6678)
         );
  AOI21_X1 U8439 ( .B1(n6679), .B2(n9948), .A(n6678), .ZN(n6680) );
  NAND2_X1 U8440 ( .A1(n6681), .A2(n6680), .ZN(P1_U3255) );
  INV_X1 U8441 ( .A(n7325), .ZN(n6729) );
  INV_X1 U8442 ( .A(n6682), .ZN(n6683) );
  NAND2_X1 U8443 ( .A1(n6683), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6685) );
  AND2_X1 U8444 ( .A1(n6685), .A2(n6684), .ZN(n9968) );
  AOI22_X1 U8445 ( .A1(n9968), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n6686), .ZN(n6687) );
  OAI21_X1 U8446 ( .B1(n6729), .B2(n9773), .A(n6687), .ZN(P1_U3337) );
  OR2_X1 U8447 ( .A1(n6688), .A2(n6847), .ZN(n6691) );
  OR2_X1 U8448 ( .A1(n7439), .A2(n6689), .ZN(n6690) );
  OAI211_X1 U8449 ( .C1(n6786), .C2(n6692), .A(n6691), .B(n6690), .ZN(n10147)
         );
  NAND2_X1 U8450 ( .A1(n6883), .A2(n10147), .ZN(n7502) );
  INV_X1 U8451 ( .A(n10147), .ZN(n6884) );
  NAND2_X1 U8452 ( .A1(n9278), .A2(n6884), .ZN(n7494) );
  NAND2_X1 U8453 ( .A1(n7502), .A2(n7494), .ZN(n7469) );
  NOR2_X1 U8454 ( .A1(n9279), .A2(n10141), .ZN(n6699) );
  NOR2_X1 U8455 ( .A1(n6699), .A2(n7615), .ZN(n10048) );
  OAI22_X2 U8456 ( .A1(n10049), .A2(n10048), .B1(n10047), .B2(n9279), .ZN(
        n6885) );
  XOR2_X1 U8457 ( .A(n7469), .B(n6885), .Z(n10151) );
  AOI211_X1 U8458 ( .C1(n10147), .C2(n10050), .A(n10012), .B(n4462), .ZN(
        n10146) );
  NOR2_X1 U8459 ( .A1(n9621), .A2(n6884), .ZN(n6697) );
  OAI22_X1 U8460 ( .A1(n10058), .A2(n6242), .B1(n6738), .B2(n10090), .ZN(n6696) );
  AOI211_X1 U8461 ( .C1(n10146), .C2(n10097), .A(n6697), .B(n6696), .ZN(n6714)
         );
  NAND2_X1 U8462 ( .A1(n7491), .A2(n7496), .ZN(n6698) );
  NAND2_X1 U8463 ( .A1(n6698), .A2(n7608), .ZN(n10043) );
  INV_X1 U8464 ( .A(n6699), .ZN(n7497) );
  AND2_X2 U8465 ( .A1(n6700), .A2(n7497), .ZN(n6909) );
  XOR2_X1 U8466 ( .A(n7469), .B(n6909), .Z(n6712) );
  INV_X1 U8467 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6701) );
  NAND2_X1 U8468 ( .A1(n6702), .A2(n6701), .ZN(n6703) );
  NAND2_X1 U8469 ( .A1(n6704), .A2(n6703), .ZN(n10036) );
  OR2_X1 U8470 ( .A1(n7430), .A2(n10036), .ZN(n6711) );
  INV_X1 U8471 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6705) );
  OR2_X1 U8472 ( .A1(n7448), .A2(n6705), .ZN(n6710) );
  INV_X1 U8473 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6706) );
  OR2_X1 U8474 ( .A1(n7445), .A2(n6706), .ZN(n6709) );
  INV_X1 U8475 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6707) );
  OR2_X1 U8476 ( .A1(n4431), .A2(n6707), .ZN(n6708) );
  NAND4_X1 U8477 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n9277)
         );
  AOI22_X1 U8478 ( .A1(n9251), .A2(n9279), .B1(n9277), .B2(n9250), .ZN(n6739)
         );
  OAI21_X1 U8479 ( .B1(n6712), .B2(n10072), .A(n6739), .ZN(n10152) );
  NAND2_X1 U8480 ( .A1(n10152), .A2(n10058), .ZN(n6713) );
  OAI211_X1 U8481 ( .C1(n10151), .C2(n9630), .A(n6714), .B(n6713), .ZN(
        P1_U3287) );
  XOR2_X1 U8482 ( .A(n6715), .B(n7930), .Z(n6721) );
  OR2_X1 U8483 ( .A1(n6716), .A2(n7930), .ZN(n6717) );
  NAND2_X1 U8484 ( .A1(n6775), .A2(n6717), .ZN(n10259) );
  OAI22_X1 U8485 ( .A1(n6760), .A2(n8480), .B1(n6894), .B2(n8481), .ZN(n6718)
         );
  AOI21_X1 U8486 ( .B1(n10259), .B2(n6719), .A(n6718), .ZN(n6720) );
  OAI21_X1 U8487 ( .B1(n6721), .B2(n8477), .A(n6720), .ZN(n10257) );
  INV_X1 U8488 ( .A(n10257), .ZN(n6727) );
  INV_X1 U8489 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6724) );
  AOI22_X1 U8490 ( .A1(n10226), .A2(n6722), .B1(n10228), .B2(n6770), .ZN(n6723) );
  OAI21_X1 U8491 ( .B1(n6724), .B2(n10233), .A(n6723), .ZN(n6725) );
  AOI21_X1 U8492 ( .B1(n10259), .B2(n7674), .A(n6725), .ZN(n6726) );
  OAI21_X1 U8493 ( .B1(n6727), .B2(n8489), .A(n6726), .ZN(P2_U3228) );
  INV_X1 U8494 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6728) );
  INV_X1 U8495 ( .A(n8287), .ZN(n8276) );
  OAI222_X1 U8496 ( .A1(n8954), .A2(n6729), .B1(n8951), .B2(n6728), .C1(
        P2_U3151), .C2(n8276), .ZN(P2_U3277) );
  NAND2_X1 U8497 ( .A1(n9278), .A2(n9121), .ZN(n6731) );
  NAND2_X1 U8498 ( .A1(n10147), .A2(n9127), .ZN(n6730) );
  NAND2_X1 U8499 ( .A1(n6731), .A2(n6730), .ZN(n6732) );
  XNOR2_X1 U8500 ( .A(n6732), .B(n9125), .ZN(n6782) );
  AOI22_X1 U8501 ( .A1(n9278), .A2(n6421), .B1(n9121), .B2(n10147), .ZN(n6781)
         );
  XNOR2_X1 U8502 ( .A(n6782), .B(n6781), .ZN(n6737) );
  INV_X1 U8503 ( .A(n6737), .ZN(n6733) );
  INV_X1 U8504 ( .A(n6784), .ZN(n6735) );
  AOI21_X1 U8505 ( .B1(n6737), .B2(n6736), .A(n6735), .ZN(n6743) );
  NOR2_X1 U8506 ( .A1(n9264), .A2(n6738), .ZN(n6741) );
  OAI22_X1 U8507 ( .A1(n6739), .A2(n9222), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8643), .ZN(n6740) );
  AOI211_X1 U8508 ( .C1(n10147), .C2(n9266), .A(n6741), .B(n6740), .ZN(n6742)
         );
  OAI21_X1 U8509 ( .B1(n6743), .B2(n9268), .A(n6742), .ZN(P1_U3239) );
  AOI211_X1 U8510 ( .C1(n6746), .C2(n6745), .A(n7070), .B(n6744), .ZN(n6757)
         );
  OAI21_X1 U8511 ( .B1(n6747), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6817), .ZN(
        n6748) );
  INV_X1 U8512 ( .A(n6748), .ZN(n6749) );
  OAI22_X1 U8513 ( .A1(n6750), .A2(n8300), .B1(n8310), .B2(n6749), .ZN(n6756)
         );
  NAND2_X1 U8514 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6759) );
  OAI21_X1 U8515 ( .B1(n6751), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6811), .ZN(
        n6752) );
  NAND2_X1 U8516 ( .A1(n8148), .A2(n6752), .ZN(n6753) );
  OAI211_X1 U8517 ( .C1(n8266), .C2(n6754), .A(n6759), .B(n6753), .ZN(n6755)
         );
  OR3_X1 U8518 ( .A1(n6757), .A2(n6756), .A3(n6755), .ZN(P2_U3187) );
  INV_X1 U8519 ( .A(P2_U3893), .ZN(n8267) );
  NAND2_X1 U8520 ( .A1(n8267), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6758) );
  OAI21_X1 U8521 ( .B1(n7953), .B2(n8267), .A(n6758), .ZN(P2_U3520) );
  INV_X1 U8522 ( .A(n6759), .ZN(n6762) );
  NOR2_X1 U8523 ( .A1(n7853), .A2(n6760), .ZN(n6761) );
  AOI211_X1 U8524 ( .C1(n7850), .C2(n8130), .A(n6762), .B(n6761), .ZN(n6763)
         );
  OAI21_X1 U8525 ( .B1(n10256), .B2(n7898), .A(n6763), .ZN(n6769) );
  XNOR2_X1 U8526 ( .A(n10256), .B(n7778), .ZN(n6827) );
  XNOR2_X1 U8527 ( .A(n6829), .B(n6827), .ZN(n6765) );
  NAND3_X1 U8528 ( .A1(n6764), .A2(n4938), .A3(n6766), .ZN(n6767) );
  AOI21_X1 U8529 ( .B1(n6831), .B2(n6767), .A(n7887), .ZN(n6768) );
  AOI211_X1 U8530 ( .C1(n6770), .C2(n7895), .A(n6769), .B(n6768), .ZN(n6771)
         );
  INV_X1 U8531 ( .A(n6771), .ZN(P2_U3167) );
  INV_X1 U8532 ( .A(n7999), .ZN(n6772) );
  NOR2_X1 U8533 ( .A1(n7929), .A2(n6772), .ZN(n6776) );
  INV_X1 U8534 ( .A(n6773), .ZN(n6774) );
  AOI21_X1 U8535 ( .B1(n6776), .B2(n6775), .A(n6774), .ZN(n10264) );
  XNOR2_X1 U8536 ( .A(n6777), .B(n7929), .ZN(n6778) );
  AOI222_X1 U8537 ( .A1(n8461), .A2(n6778), .B1(n8129), .B2(n8463), .C1(n8131), 
        .C2(n8466), .ZN(n10261) );
  MUX2_X1 U8538 ( .A(n5844), .B(n10261), .S(n10233), .Z(n6780) );
  AOI22_X1 U8539 ( .A1(n10226), .A2(n6840), .B1(n10228), .B2(n6837), .ZN(n6779) );
  OAI211_X1 U8540 ( .C1(n10264), .C2(n8783), .A(n6780), .B(n6779), .ZN(
        P2_U3227) );
  NAND2_X1 U8541 ( .A1(n6782), .A2(n6781), .ZN(n6783) );
  NAND2_X1 U8542 ( .A1(n9277), .A2(n9121), .ZN(n6790) );
  OR2_X1 U8543 ( .A1(n6785), .A2(n6847), .ZN(n6788) );
  AOI22_X1 U8544 ( .A1(n7339), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7338), .B2(
        n9802), .ZN(n6787) );
  NAND2_X1 U8545 ( .A1(n10038), .A2(n9127), .ZN(n6789) );
  NAND2_X1 U8546 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  XNOR2_X1 U8547 ( .A(n6791), .B(n9125), .ZN(n7023) );
  NAND2_X1 U8548 ( .A1(n9277), .A2(n6421), .ZN(n6793) );
  NAND2_X1 U8549 ( .A1(n10038), .A2(n9121), .ZN(n6792) );
  AND2_X1 U8550 ( .A1(n6793), .A2(n6792), .ZN(n7024) );
  XNOR2_X1 U8551 ( .A(n7023), .B(n7024), .ZN(n6794) );
  XNOR2_X1 U8552 ( .A(n7028), .B(n6794), .ZN(n6800) );
  NAND2_X1 U8553 ( .A1(n7111), .A2(n9250), .ZN(n6796) );
  NAND2_X1 U8554 ( .A1(n9278), .A2(n9251), .ZN(n6795) );
  NAND2_X1 U8555 ( .A1(n6796), .A2(n6795), .ZN(n10035) );
  AOI22_X1 U8556 ( .A1(n10035), .A2(n9262), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n6797) );
  OAI21_X1 U8557 ( .B1(n9264), .B2(n10036), .A(n6797), .ZN(n6798) );
  AOI21_X1 U8558 ( .B1(n10038), .B2(n9266), .A(n6798), .ZN(n6799) );
  OAI21_X1 U8559 ( .B1(n6800), .B2(n9268), .A(n6799), .ZN(P1_U3213) );
  INV_X1 U8560 ( .A(n7337), .ZN(n6801) );
  OAI222_X1 U8561 ( .A1(P2_U3151), .A2(n8291), .B1(n7046), .B2(n6801), .C1(
        n8951), .C2(n8603), .ZN(P2_U3276) );
  INV_X1 U8562 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6802) );
  OAI222_X1 U8563 ( .A1(n9769), .A2(n6802), .B1(n9777), .B2(n6801), .C1(
        P1_U3086), .C2(n6507), .ZN(P1_U3336) );
  OAI21_X1 U8564 ( .B1(n6805), .B2(n6804), .A(n6803), .ZN(n6806) );
  NAND2_X1 U8565 ( .A1(n6806), .A2(n8309), .ZN(n6826) );
  NAND2_X1 U8566 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8567 ( .B1(n8266), .B2(n6807), .A(n6838), .ZN(n6824) );
  INV_X1 U8568 ( .A(n6808), .ZN(n6810) );
  NAND3_X1 U8569 ( .A1(n6811), .A2(n6810), .A3(n6809), .ZN(n6812) );
  AOI21_X1 U8570 ( .B1(n6813), .B2(n6812), .A(n8306), .ZN(n6823) );
  INV_X1 U8571 ( .A(n6814), .ZN(n6816) );
  NAND3_X1 U8572 ( .A1(n6817), .A2(n6816), .A3(n6815), .ZN(n6818) );
  AOI21_X1 U8573 ( .B1(n6819), .B2(n6818), .A(n8310), .ZN(n6822) );
  INV_X1 U8574 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6820) );
  NOR2_X1 U8575 ( .A1(n8300), .A2(n6820), .ZN(n6821) );
  NOR4_X1 U8576 ( .A1(n6824), .A2(n6823), .A3(n6822), .A4(n6821), .ZN(n6825)
         );
  NAND2_X1 U8577 ( .A1(n6826), .A2(n6825), .ZN(P2_U3188) );
  XNOR2_X1 U8578 ( .A(n7705), .B(n6840), .ZN(n6945) );
  XNOR2_X1 U8579 ( .A(n6945), .B(n8130), .ZN(n6836) );
  INV_X1 U8580 ( .A(n6827), .ZN(n6828) );
  NAND2_X1 U8581 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  INV_X1 U8582 ( .A(n6947), .ZN(n6834) );
  AOI211_X1 U8583 ( .C1(n6836), .C2(n6835), .A(n7887), .B(n6834), .ZN(n6846)
         );
  NAND2_X1 U8584 ( .A1(n7895), .A2(n6837), .ZN(n6844) );
  INV_X1 U8585 ( .A(n6838), .ZN(n6839) );
  AOI21_X1 U8586 ( .B1(n7850), .B2(n8129), .A(n6839), .ZN(n6843) );
  NAND2_X1 U8587 ( .A1(n7883), .A2(n6840), .ZN(n6842) );
  NAND2_X1 U8588 ( .A1(n7891), .A2(n8131), .ZN(n6841) );
  NAND4_X1 U8589 ( .A1(n6844), .A2(n6843), .A3(n6842), .A4(n6841), .ZN(n6845)
         );
  OR2_X1 U8590 ( .A1(n6846), .A2(n6845), .ZN(P2_U3179) );
  NAND2_X1 U8591 ( .A1(n6848), .A2(n7425), .ZN(n6851) );
  AOI22_X1 U8592 ( .A1(n7339), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7338), .B2(
        n6849), .ZN(n6850) );
  INV_X1 U8593 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U8594 ( .A1(n6853), .A2(n6852), .ZN(n6854) );
  NAND2_X1 U8595 ( .A1(n6871), .A2(n6854), .ZN(n10021) );
  OR2_X1 U8596 ( .A1(n7430), .A2(n10021), .ZN(n6861) );
  OR2_X1 U8597 ( .A1(n7296), .A2(n6855), .ZN(n6860) );
  INV_X1 U8598 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n6856) );
  OR2_X1 U8599 ( .A1(n4431), .A2(n6856), .ZN(n6859) );
  OR2_X1 U8600 ( .A1(n7445), .A2(n6857), .ZN(n6858) );
  NAND4_X1 U8601 ( .A1(n6861), .A2(n6860), .A3(n6859), .A4(n6858), .ZN(n9276)
         );
  INV_X1 U8602 ( .A(n9276), .ZN(n6916) );
  INV_X1 U8603 ( .A(n6887), .ZN(n7515) );
  NAND2_X1 U8604 ( .A1(n6862), .A2(n7425), .ZN(n6864) );
  AOI22_X1 U8605 ( .A1(n7339), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7338), .B2(
        n9814), .ZN(n6863) );
  NAND2_X1 U8606 ( .A1(n6864), .A2(n6863), .ZN(n7029) );
  OR2_X1 U8607 ( .A1(n6886), .A2(n7029), .ZN(n10016) );
  NAND2_X1 U8608 ( .A1(n7029), .A2(n6886), .ZN(n7508) );
  INV_X1 U8609 ( .A(n9277), .ZN(n6917) );
  NAND2_X1 U8610 ( .A1(n6917), .A2(n10038), .ZN(n6910) );
  NAND2_X1 U8611 ( .A1(n7508), .A2(n6910), .ZN(n7511) );
  AND2_X1 U8612 ( .A1(n10024), .A2(n6916), .ZN(n7507) );
  INV_X1 U8613 ( .A(n7510), .ZN(n6866) );
  INV_X1 U8614 ( .A(n10038), .ZN(n10155) );
  NAND2_X1 U8615 ( .A1(n10155), .A2(n9277), .ZN(n7506) );
  INV_X1 U8616 ( .A(n7506), .ZN(n6865) );
  NOR2_X1 U8617 ( .A1(n6866), .A2(n6865), .ZN(n7463) );
  NAND2_X1 U8618 ( .A1(n7463), .A2(n7494), .ZN(n6867) );
  NAND2_X1 U8619 ( .A1(n7612), .A2(n7616), .ZN(n6879) );
  NAND2_X1 U8620 ( .A1(n6868), .A2(n7425), .ZN(n6870) );
  AOI22_X1 U8621 ( .A1(n7339), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7338), .B2(
        n9789), .ZN(n6869) );
  NAND2_X1 U8622 ( .A1(n6870), .A2(n6869), .ZN(n7134) );
  NAND2_X1 U8623 ( .A1(n6871), .A2(n8562), .ZN(n6872) );
  NAND2_X1 U8624 ( .A1(n6997), .A2(n6872), .ZN(n7132) );
  OR2_X1 U8625 ( .A1(n7430), .A2(n7132), .ZN(n6878) );
  OR2_X1 U8626 ( .A1(n7296), .A2(n8568), .ZN(n6877) );
  INV_X1 U8627 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6873) );
  OR2_X1 U8628 ( .A1(n4432), .A2(n6873), .ZN(n6876) );
  OR2_X1 U8629 ( .A1(n7445), .A2(n6874), .ZN(n6875) );
  NAND4_X1 U8630 ( .A1(n6878), .A2(n6877), .A3(n6876), .A4(n6875), .ZN(n9275)
         );
  INV_X1 U8631 ( .A(n9275), .ZN(n7015) );
  OR2_X1 U8632 ( .A1(n7134), .A2(n7015), .ZN(n7617) );
  NAND2_X1 U8633 ( .A1(n7134), .A2(n7015), .ZN(n7516) );
  NAND2_X1 U8634 ( .A1(n7617), .A2(n7516), .ZN(n7016) );
  XNOR2_X1 U8635 ( .A(n6879), .B(n7016), .ZN(n6882) );
  NAND2_X1 U8636 ( .A1(n8963), .A2(n9250), .ZN(n6881) );
  NAND2_X1 U8637 ( .A1(n9276), .A2(n9251), .ZN(n6880) );
  NAND2_X1 U8638 ( .A1(n6881), .A2(n6880), .ZN(n7130) );
  AOI21_X1 U8639 ( .B1(n6882), .B2(n10112), .A(n7130), .ZN(n10171) );
  NAND2_X1 U8640 ( .A1(n10016), .A2(n7508), .ZN(n6913) );
  INV_X1 U8641 ( .A(n7029), .ZN(n10162) );
  NOR2_X1 U8642 ( .A1(n6887), .A2(n7507), .ZN(n10019) );
  XNOR2_X1 U8643 ( .A(n7017), .B(n7016), .ZN(n10174) );
  NAND2_X1 U8644 ( .A1(n10174), .A2(n10066), .ZN(n6891) );
  OAI22_X1 U8645 ( .A1(n10058), .A2(n8568), .B1(n7132), .B2(n10090), .ZN(n6889) );
  INV_X1 U8646 ( .A(n7134), .ZN(n10172) );
  NAND2_X1 U8647 ( .A1(n10011), .A2(n10172), .ZN(n10003) );
  OAI211_X1 U8648 ( .C1(n10011), .C2(n10172), .A(n10003), .B(n10081), .ZN(
        n10170) );
  NOR2_X1 U8649 ( .A1(n10170), .A2(n9671), .ZN(n6888) );
  AOI211_X1 U8650 ( .C1(n10077), .C2(n7134), .A(n6889), .B(n6888), .ZN(n6890)
         );
  OAI211_X1 U8651 ( .C1(n10100), .C2(n10171), .A(n6891), .B(n6890), .ZN(
        P1_U3283) );
  XOR2_X1 U8652 ( .A(n6892), .B(n7989), .Z(n6893) );
  OAI222_X1 U8653 ( .A1(n8480), .A2(n6894), .B1(n8481), .B2(n7088), .C1(n8477), 
        .C2(n6893), .ZN(n6922) );
  INV_X1 U8654 ( .A(n6922), .ZN(n6903) );
  NOR2_X1 U8655 ( .A1(n8431), .A2(n6960), .ZN(n6897) );
  INV_X1 U8656 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6938) );
  INV_X1 U8657 ( .A(n6895), .ZN(n6956) );
  OAI22_X1 U8658 ( .A1(n10233), .A2(n6938), .B1(n6956), .B2(n8444), .ZN(n6896)
         );
  NOR2_X1 U8659 ( .A1(n6897), .A2(n6896), .ZN(n6902) );
  NAND2_X1 U8660 ( .A1(n6899), .A2(n7989), .ZN(n6900) );
  AND2_X1 U8661 ( .A1(n6898), .A2(n6900), .ZN(n6923) );
  NAND2_X1 U8662 ( .A1(n6923), .A2(n8486), .ZN(n6901) );
  OAI211_X1 U8663 ( .C1(n6903), .C2(n8489), .A(n6902), .B(n6901), .ZN(P2_U3226) );
  INV_X1 U8664 ( .A(n7415), .ZN(n6929) );
  OAI222_X1 U8665 ( .A1(n8954), .A2(n6929), .B1(n8951), .B2(n5494), .C1(n8100), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  XNOR2_X1 U8666 ( .A(n6904), .B(n6913), .ZN(n10164) );
  XNOR2_X1 U8667 ( .A(n10039), .B(n7029), .ZN(n6905) );
  NAND2_X1 U8668 ( .A1(n6905), .A2(n10081), .ZN(n10160) );
  OAI22_X1 U8669 ( .A1(n10058), .A2(n6906), .B1(n7039), .B2(n10090), .ZN(n6907) );
  AOI21_X1 U8670 ( .B1(n10077), .B2(n7029), .A(n6907), .ZN(n6908) );
  OAI21_X1 U8671 ( .B1(n10160), .B2(n9671), .A(n6908), .ZN(n6920) );
  INV_X1 U8672 ( .A(n7494), .ZN(n7501) );
  OAI21_X1 U8673 ( .B1(n6909), .B2(n7501), .A(n7502), .ZN(n10031) );
  INV_X1 U8674 ( .A(n6910), .ZN(n6911) );
  AOI21_X1 U8675 ( .B1(n10031), .B2(n10032), .A(n6911), .ZN(n6915) );
  INV_X1 U8676 ( .A(n6915), .ZN(n6912) );
  AOI21_X1 U8677 ( .B1(n6912), .B2(n6913), .A(n10072), .ZN(n6918) );
  INV_X1 U8678 ( .A(n6913), .ZN(n6914) );
  NAND2_X1 U8679 ( .A1(n6915), .A2(n6914), .ZN(n10017) );
  OAI22_X1 U8680 ( .A1(n6917), .A2(n9475), .B1(n6916), .B2(n9406), .ZN(n7042)
         );
  AOI21_X1 U8681 ( .B1(n6918), .B2(n10017), .A(n7042), .ZN(n10161) );
  NOR2_X1 U8682 ( .A1(n10161), .A2(n10100), .ZN(n6919) );
  AOI211_X1 U8683 ( .C1(n10066), .C2(n10164), .A(n6920), .B(n6919), .ZN(n6921)
         );
  INV_X1 U8684 ( .A(n6921), .ZN(P1_U3285) );
  AOI21_X1 U8685 ( .B1(n6923), .B2(n10274), .A(n6922), .ZN(n6928) );
  AOI22_X1 U8686 ( .A1(n8843), .A2(n6948), .B1(n5770), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n6924) );
  OAI21_X1 U8687 ( .B1(n6928), .B2(n5770), .A(n6924), .ZN(P2_U3466) );
  INV_X1 U8688 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6925) );
  OAI22_X1 U8689 ( .A1(n8909), .A2(n6960), .B1(n6925), .B2(n10275), .ZN(n6926)
         );
  INV_X1 U8690 ( .A(n6926), .ZN(n6927) );
  OAI21_X1 U8691 ( .B1(n6928), .B2(n10277), .A(n6927), .ZN(P2_U3411) );
  OAI222_X1 U8692 ( .A1(n9769), .A2(n7416), .B1(n9777), .B2(n6929), .C1(n10092), .C2(P1_U3086), .ZN(P1_U3335) );
  XOR2_X1 U8693 ( .A(n6931), .B(n6930), .Z(n6944) );
  OAI21_X1 U8694 ( .B1(n6932), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6976), .ZN(
        n6942) );
  INV_X1 U8695 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U8696 ( .A1(n8297), .A2(n4659), .ZN(n6933) );
  NAND2_X1 U8697 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6952) );
  OAI211_X1 U8698 ( .C1(n6934), .C2(n8300), .A(n6933), .B(n6952), .ZN(n6941)
         );
  INV_X1 U8699 ( .A(n6935), .ZN(n6937) );
  INV_X1 U8700 ( .A(n6936), .ZN(n6985) );
  AOI21_X1 U8701 ( .B1(n6938), .B2(n6937), .A(n6985), .ZN(n6939) );
  NOR2_X1 U8702 ( .A1(n6939), .A2(n8306), .ZN(n6940) );
  AOI211_X1 U8703 ( .C1(n8140), .C2(n6942), .A(n6941), .B(n6940), .ZN(n6943)
         );
  OAI21_X1 U8704 ( .B1(n6944), .B2(n7070), .A(n6943), .ZN(P2_U3189) );
  NAND2_X1 U8705 ( .A1(n6945), .A2(n8130), .ZN(n6946) );
  XNOR2_X1 U8706 ( .A(n7705), .B(n6948), .ZN(n7082) );
  XNOR2_X1 U8707 ( .A(n7084), .B(n7082), .ZN(n6949) );
  OAI21_X1 U8708 ( .B1(n6950), .B2(n6949), .A(n7085), .ZN(n6951) );
  NAND2_X1 U8709 ( .A1(n6951), .A2(n7871), .ZN(n6959) );
  INV_X1 U8710 ( .A(n6952), .ZN(n6953) );
  AOI21_X1 U8711 ( .B1(n7850), .B2(n8128), .A(n6953), .ZN(n6955) );
  NAND2_X1 U8712 ( .A1(n7891), .A2(n8130), .ZN(n6954) );
  OAI211_X1 U8713 ( .C1(n7821), .C2(n6956), .A(n6955), .B(n6954), .ZN(n6957)
         );
  INV_X1 U8714 ( .A(n6957), .ZN(n6958) );
  OAI211_X1 U8715 ( .C1(n6960), .C2(n7898), .A(n6959), .B(n6958), .ZN(P2_U3153) );
  NAND2_X1 U8716 ( .A1(n7958), .A2(n7957), .ZN(n7932) );
  NAND2_X1 U8717 ( .A1(n6898), .A2(n6961), .ZN(n6962) );
  XOR2_X1 U8718 ( .A(n7932), .B(n6962), .Z(n10268) );
  XNOR2_X1 U8719 ( .A(n6963), .B(n7932), .ZN(n6964) );
  AOI222_X1 U8720 ( .A1(n8461), .A2(n6964), .B1(n8127), .B2(n8463), .C1(n8129), 
        .C2(n8466), .ZN(n10269) );
  MUX2_X1 U8721 ( .A(n6965), .B(n10269), .S(n10233), .Z(n6967) );
  AOI22_X1 U8722 ( .A1(n10226), .A2(n7086), .B1(n10228), .B2(n7089), .ZN(n6966) );
  OAI211_X1 U8723 ( .C1(n10268), .C2(n8783), .A(n6967), .B(n6966), .ZN(
        P2_U3225) );
  INV_X1 U8724 ( .A(n7401), .ZN(n6970) );
  OAI222_X1 U8725 ( .A1(n8954), .A2(n6970), .B1(P2_U3151), .B2(n6969), .C1(
        n6968), .C2(n8951), .ZN(P2_U3274) );
  OAI222_X1 U8726 ( .A1(n9769), .A2(n7402), .B1(n9777), .B2(n6970), .C1(n4922), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  XOR2_X1 U8727 ( .A(n6972), .B(n6971), .Z(n6991) );
  INV_X1 U8728 ( .A(n8300), .ZN(n8195) );
  INV_X1 U8729 ( .A(n6973), .ZN(n6975) );
  NAND3_X1 U8730 ( .A1(n6976), .A2(n6975), .A3(n6974), .ZN(n6977) );
  AOI21_X1 U8731 ( .B1(n6978), .B2(n6977), .A(n8310), .ZN(n6981) );
  NAND2_X1 U8732 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7090) );
  OAI21_X1 U8733 ( .B1(n8266), .B2(n6979), .A(n7090), .ZN(n6980) );
  AOI211_X1 U8734 ( .C1(n8195), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6981), .B(
        n6980), .ZN(n6990) );
  INV_X1 U8735 ( .A(n6982), .ZN(n6984) );
  NOR3_X1 U8736 ( .A1(n6985), .A2(n6984), .A3(n6983), .ZN(n6988) );
  INV_X1 U8737 ( .A(n6986), .ZN(n6987) );
  OAI21_X1 U8738 ( .B1(n6988), .B2(n6987), .A(n8148), .ZN(n6989) );
  OAI211_X1 U8739 ( .C1(n6991), .C2(n7070), .A(n6990), .B(n6989), .ZN(P2_U3190) );
  NAND2_X1 U8740 ( .A1(n6992), .A2(n7425), .ZN(n6994) );
  AOI22_X1 U8741 ( .A1(n7339), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7338), .B2(
        n9368), .ZN(n6993) );
  INV_X1 U8742 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6995) );
  OAI21_X1 U8743 ( .B1(n6997), .B2(n6996), .A(n6995), .ZN(n6999) );
  NAND2_X1 U8744 ( .A1(n6999), .A2(n6998), .ZN(n9154) );
  OR2_X1 U8745 ( .A1(n7430), .A2(n9154), .ZN(n7004) );
  INV_X1 U8746 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7018) );
  OR2_X1 U8747 ( .A1(n7296), .A2(n7018), .ZN(n7003) );
  OR2_X1 U8748 ( .A1(n7445), .A2(n10216), .ZN(n7002) );
  INV_X1 U8749 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7000) );
  OR2_X1 U8750 ( .A1(n4432), .A2(n7000), .ZN(n7001) );
  NAND4_X1 U8751 ( .A1(n7004), .A2(n7003), .A3(n7002), .A4(n7001), .ZN(n9274)
         );
  NAND2_X1 U8752 ( .A1(n9156), .A2(n9414), .ZN(n7525) );
  NAND2_X1 U8753 ( .A1(n7519), .A2(n7525), .ZN(n9415) );
  INV_X1 U8754 ( .A(n9415), .ZN(n7474) );
  NAND2_X1 U8755 ( .A1(n7005), .A2(n7425), .ZN(n7007) );
  AOI22_X1 U8756 ( .A1(n7339), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7338), .B2(
        n9895), .ZN(n7006) );
  INV_X1 U8757 ( .A(n8963), .ZN(n7009) );
  INV_X1 U8758 ( .A(n7518), .ZN(n7008) );
  NOR2_X1 U8759 ( .A1(n7474), .A2(n7008), .ZN(n7011) );
  INV_X1 U8760 ( .A(n7016), .ZN(n7473) );
  NAND2_X1 U8761 ( .A1(n10002), .A2(n7009), .ZN(n7517) );
  NAND2_X1 U8762 ( .A1(n9993), .A2(n7518), .ZN(n7010) );
  NAND2_X1 U8763 ( .A1(n7010), .A2(n7474), .ZN(n7278) );
  INV_X1 U8764 ( .A(n7278), .ZN(n9975) );
  AOI211_X1 U8765 ( .C1(n7011), .C2(n9993), .A(n10072), .B(n9975), .ZN(n7014)
         );
  NAND2_X1 U8766 ( .A1(n8963), .A2(n9251), .ZN(n7013) );
  NAND2_X1 U8767 ( .A1(n9417), .A2(n9250), .ZN(n7012) );
  NAND2_X1 U8768 ( .A1(n7013), .A2(n7012), .ZN(n9151) );
  NOR2_X1 U8769 ( .A1(n7014), .A2(n9151), .ZN(n10182) );
  XNOR2_X1 U8770 ( .A(n9416), .B(n9415), .ZN(n10185) );
  NAND2_X1 U8771 ( .A1(n10185), .A2(n10066), .ZN(n7022) );
  OAI22_X1 U8772 ( .A1(n10058), .A2(n7018), .B1(n9154), .B2(n10090), .ZN(n7020) );
  OAI211_X1 U8773 ( .C1(n10004), .C2(n10183), .A(n9985), .B(n10081), .ZN(
        n10181) );
  NOR2_X1 U8774 ( .A1(n10181), .A2(n9671), .ZN(n7019) );
  AOI211_X1 U8775 ( .C1(n10077), .C2(n9156), .A(n7020), .B(n7019), .ZN(n7021)
         );
  OAI211_X1 U8776 ( .C1(n10100), .C2(n10182), .A(n7022), .B(n7021), .ZN(
        P1_U3281) );
  AOI22_X1 U8777 ( .A1(n7029), .A2(n9121), .B1(n6421), .B2(n7111), .ZN(n7037)
         );
  AND2_X1 U8778 ( .A1(n7023), .A2(n7024), .ZN(n7027) );
  INV_X1 U8779 ( .A(n7023), .ZN(n7026) );
  INV_X1 U8780 ( .A(n7024), .ZN(n7025) );
  NAND2_X1 U8781 ( .A1(n7029), .A2(n9127), .ZN(n7031) );
  NAND2_X1 U8782 ( .A1(n7111), .A2(n9121), .ZN(n7030) );
  NAND2_X1 U8783 ( .A1(n7031), .A2(n7030), .ZN(n7032) );
  XNOR2_X1 U8784 ( .A(n7032), .B(n9075), .ZN(n7033) );
  NAND2_X1 U8785 ( .A1(n7036), .A2(n7037), .ZN(n7101) );
  OAI21_X1 U8786 ( .B1(n7037), .B2(n7036), .A(n7101), .ZN(n7038) );
  NAND2_X1 U8787 ( .A1(n7038), .A2(n9247), .ZN(n7044) );
  NAND2_X1 U8788 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9815) );
  INV_X1 U8789 ( .A(n9815), .ZN(n7041) );
  NOR2_X1 U8790 ( .A1(n9264), .A2(n7039), .ZN(n7040) );
  AOI211_X1 U8791 ( .C1(n9262), .C2(n7042), .A(n7041), .B(n7040), .ZN(n7043)
         );
  OAI211_X1 U8792 ( .C1(n10162), .C2(n9258), .A(n7044), .B(n7043), .ZN(
        P1_U3221) );
  INV_X1 U8793 ( .A(n7364), .ZN(n7048) );
  OAI222_X1 U8794 ( .A1(n8951), .A2(n7047), .B1(n7046), .B2(n7048), .C1(n7045), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U8795 ( .A1(n9769), .A2(n7365), .B1(n9777), .B2(n7048), .C1(
        P1_U3086), .C2(n9685), .ZN(P1_U3333) );
  XNOR2_X1 U8796 ( .A(n7049), .B(n7052), .ZN(n7050) );
  OAI222_X1 U8797 ( .A1(n8480), .A2(n7051), .B1(n8481), .B2(n7801), .C1(n7050), 
        .C2(n8477), .ZN(n7137) );
  INV_X1 U8798 ( .A(n7137), .ZN(n7056) );
  INV_X1 U8799 ( .A(n7052), .ZN(n7935) );
  OAI21_X1 U8800 ( .B1(n4519), .B2(n7935), .A(n7144), .ZN(n7138) );
  INV_X1 U8801 ( .A(n7765), .ZN(n7143) );
  AOI22_X1 U8802 ( .A1(n8489), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10228), .B2(
        n7754), .ZN(n7053) );
  OAI21_X1 U8803 ( .B1(n7143), .B2(n8431), .A(n7053), .ZN(n7054) );
  AOI21_X1 U8804 ( .B1(n7138), .B2(n8486), .A(n7054), .ZN(n7055) );
  OAI21_X1 U8805 ( .B1(n7056), .B2(n8489), .A(n7055), .ZN(P2_U3223) );
  XOR2_X1 U8806 ( .A(n7058), .B(n7057), .Z(n7071) );
  OAI21_X1 U8807 ( .B1(n7060), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7059), .ZN(
        n7068) );
  NOR2_X1 U8808 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5177), .ZN(n7179) );
  AOI21_X1 U8809 ( .B1(n8195), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7179), .ZN(
        n7061) );
  OAI21_X1 U8810 ( .B1(n8266), .B2(n7062), .A(n7061), .ZN(n7067) );
  NAND2_X1 U8811 ( .A1(n7063), .A2(n7078), .ZN(n7064) );
  AOI21_X1 U8812 ( .B1(n7065), .B2(n7064), .A(n8310), .ZN(n7066) );
  AOI211_X1 U8813 ( .C1(n8148), .C2(n7068), .A(n7067), .B(n7066), .ZN(n7069)
         );
  OAI21_X1 U8814 ( .B1(n7071), .B2(n7070), .A(n7069), .ZN(P2_U3191) );
  INV_X1 U8815 ( .A(n10274), .ZN(n10263) );
  XNOR2_X1 U8816 ( .A(n7072), .B(n7933), .ZN(n10224) );
  XOR2_X1 U8817 ( .A(n7073), .B(n7933), .Z(n7074) );
  AOI222_X1 U8818 ( .A1(n8461), .A2(n7074), .B1(n8126), .B2(n8463), .C1(n8128), 
        .C2(n8466), .ZN(n10223) );
  OAI21_X1 U8819 ( .B1(n10263), .B2(n10224), .A(n10223), .ZN(n7080) );
  INV_X1 U8820 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7075) );
  OAI22_X1 U8821 ( .A1(n8909), .A2(n7182), .B1(n7075), .B2(n10275), .ZN(n7076)
         );
  AOI21_X1 U8822 ( .B1(n7080), .B2(n10275), .A(n7076), .ZN(n7077) );
  INV_X1 U8823 ( .A(n7077), .ZN(P2_U3417) );
  OAI22_X1 U8824 ( .A1(n8831), .A2(n7182), .B1(n10289), .B2(n7078), .ZN(n7079)
         );
  AOI21_X1 U8825 ( .B1(n7080), .B2(n10289), .A(n7079), .ZN(n7081) );
  INV_X1 U8826 ( .A(n7081), .ZN(P2_U3468) );
  INV_X1 U8827 ( .A(n7082), .ZN(n7083) );
  XNOR2_X1 U8828 ( .A(n7086), .B(n7705), .ZN(n7183) );
  OAI21_X1 U8829 ( .B1(n7088), .B2(n7087), .A(n7187), .ZN(n7097) );
  NOR2_X1 U8830 ( .A1(n7898), .A2(n10271), .ZN(n7096) );
  INV_X1 U8831 ( .A(n7089), .ZN(n7094) );
  INV_X1 U8832 ( .A(n7090), .ZN(n7091) );
  AOI21_X1 U8833 ( .B1(n7850), .B2(n8127), .A(n7091), .ZN(n7093) );
  NAND2_X1 U8834 ( .A1(n7891), .A2(n8129), .ZN(n7092) );
  OAI211_X1 U8835 ( .C1(n7821), .C2(n7094), .A(n7093), .B(n7092), .ZN(n7095)
         );
  AOI211_X1 U8836 ( .C1(n7097), .C2(n7871), .A(n7096), .B(n7095), .ZN(n7098)
         );
  INV_X1 U8837 ( .A(n7098), .ZN(P2_U3161) );
  INV_X1 U8838 ( .A(n10024), .ZN(n10167) );
  INV_X1 U8839 ( .A(n7099), .ZN(n7100) );
  NAND2_X1 U8840 ( .A1(n7101), .A2(n7100), .ZN(n7107) );
  NAND2_X1 U8841 ( .A1(n10024), .A2(n9127), .ZN(n7103) );
  NAND2_X1 U8842 ( .A1(n9276), .A2(n9121), .ZN(n7102) );
  NAND2_X1 U8843 ( .A1(n7103), .A2(n7102), .ZN(n7104) );
  XNOR2_X1 U8844 ( .A(n7104), .B(n9125), .ZN(n7106) );
  AOI22_X1 U8845 ( .A1(n10024), .A2(n9121), .B1(n6421), .B2(n9276), .ZN(n7105)
         );
  OR2_X1 U8846 ( .A1(n7106), .A2(n7105), .ZN(n7108) );
  NAND2_X1 U8847 ( .A1(n7106), .A2(n7105), .ZN(n7123) );
  NOR2_X1 U8848 ( .A1(n7124), .A2(n4910), .ZN(n7110) );
  AOI21_X1 U8849 ( .B1(n7108), .B2(n7123), .A(n7107), .ZN(n7109) );
  OAI21_X1 U8850 ( .B1(n7110), .B2(n7109), .A(n9247), .ZN(n7118) );
  NAND2_X1 U8851 ( .A1(n7111), .A2(n9251), .ZN(n7113) );
  NAND2_X1 U8852 ( .A1(n9275), .A2(n9250), .ZN(n7112) );
  NAND2_X1 U8853 ( .A1(n7113), .A2(n7112), .ZN(n10014) );
  NAND2_X1 U8854 ( .A1(n10014), .A2(n9262), .ZN(n7115) );
  OAI211_X1 U8855 ( .C1(n9264), .C2(n10021), .A(n7115), .B(n7114), .ZN(n7116)
         );
  INV_X1 U8856 ( .A(n7116), .ZN(n7117) );
  OAI211_X1 U8857 ( .C1(n10167), .C2(n9258), .A(n7118), .B(n7117), .ZN(
        P1_U3231) );
  NAND2_X1 U8858 ( .A1(n7354), .A2(n7119), .ZN(n7120) );
  OAI211_X1 U8859 ( .C1(n7355), .C2(n9769), .A(n7120), .B(n7667), .ZN(P1_U3332) );
  NAND2_X1 U8860 ( .A1(n7354), .A2(n8946), .ZN(n7122) );
  NAND2_X1 U8861 ( .A1(n7121), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8121) );
  OAI211_X1 U8862 ( .C1(n8573), .C2(n8951), .A(n7122), .B(n8121), .ZN(P2_U3272) );
  NAND2_X1 U8863 ( .A1(n7134), .A2(n9127), .ZN(n7126) );
  NAND2_X1 U8864 ( .A1(n9275), .A2(n9121), .ZN(n7125) );
  NAND2_X1 U8865 ( .A1(n7126), .A2(n7125), .ZN(n7127) );
  XNOR2_X1 U8866 ( .A(n7127), .B(n9125), .ZN(n8958) );
  AND2_X1 U8867 ( .A1(n9275), .A2(n6421), .ZN(n7128) );
  AOI21_X1 U8868 ( .B1(n7134), .B2(n9121), .A(n7128), .ZN(n8959) );
  XNOR2_X1 U8869 ( .A(n8958), .B(n8959), .ZN(n7129) );
  XNOR2_X1 U8870 ( .A(n8957), .B(n7129), .ZN(n7136) );
  AOI22_X1 U8871 ( .A1(n7130), .A2(n9262), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n7131) );
  OAI21_X1 U8872 ( .B1(n9264), .B2(n7132), .A(n7131), .ZN(n7133) );
  AOI21_X1 U8873 ( .B1(n7134), .B2(n9266), .A(n7133), .ZN(n7135) );
  OAI21_X1 U8874 ( .B1(n7136), .B2(n9268), .A(n7135), .ZN(P1_U3217) );
  INV_X1 U8875 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7139) );
  AOI21_X1 U8876 ( .B1(n10274), .B2(n7138), .A(n7137), .ZN(n7141) );
  MUX2_X1 U8877 ( .A(n7139), .B(n7141), .S(n10275), .Z(n7140) );
  OAI21_X1 U8878 ( .B1(n7143), .B2(n8909), .A(n7140), .ZN(P2_U3420) );
  MUX2_X1 U8879 ( .A(n5828), .B(n7141), .S(n10289), .Z(n7142) );
  OAI21_X1 U8880 ( .B1(n7143), .B2(n8831), .A(n7142), .ZN(P2_U3469) );
  NAND2_X1 U8881 ( .A1(n7144), .A2(n8020), .ZN(n7145) );
  XNOR2_X1 U8882 ( .A(n7211), .B(n7145), .ZN(n8782) );
  INV_X1 U8883 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7148) );
  INV_X1 U8884 ( .A(n7211), .ZN(n7936) );
  XNOR2_X1 U8885 ( .A(n7146), .B(n7936), .ZN(n7147) );
  AOI222_X1 U8886 ( .A1(n8461), .A2(n7147), .B1(n8126), .B2(n8466), .C1(n8124), 
        .C2(n8463), .ZN(n8776) );
  MUX2_X1 U8887 ( .A(n7148), .B(n8776), .S(n10275), .Z(n7150) );
  NAND2_X1 U8888 ( .A1(n8930), .A2(n4556), .ZN(n7149) );
  OAI211_X1 U8889 ( .C1(n8782), .C2(n8919), .A(n7150), .B(n7149), .ZN(P2_U3423) );
  INV_X1 U8890 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7151) );
  MUX2_X1 U8891 ( .A(n7151), .B(n8776), .S(n10289), .Z(n7153) );
  NAND2_X1 U8892 ( .A1(n4556), .A2(n8843), .ZN(n7152) );
  OAI211_X1 U8893 ( .C1(n8782), .C2(n8837), .A(n7153), .B(n7152), .ZN(P2_U3470) );
  MUX2_X1 U8894 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8292), .Z(n7222) );
  XNOR2_X1 U8895 ( .A(n7222), .B(n7167), .ZN(n7157) );
  OAI21_X1 U8896 ( .B1(n7158), .B2(n7157), .A(n7223), .ZN(n7159) );
  NAND2_X1 U8897 ( .A1(n7159), .A2(n8309), .ZN(n7174) );
  AOI21_X1 U8898 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7163), .A(n7160), .ZN(
        n7161) );
  NOR2_X1 U8899 ( .A1(n7161), .A2(n7167), .ZN(n7218) );
  OAI21_X1 U8900 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7162), .A(n8139), .ZN(
        n7172) );
  AOI21_X1 U8901 ( .B1(n7164), .B2(n7167), .A(n7232), .ZN(n7165) );
  INV_X1 U8902 ( .A(n7165), .ZN(n7166) );
  INV_X1 U8903 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8777) );
  AOI21_X1 U8904 ( .B1(n7166), .B2(n8777), .A(n7231), .ZN(n7170) );
  AND2_X1 U8905 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7212) );
  AOI21_X1 U8906 ( .B1(n8195), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7212), .ZN(
        n7169) );
  NAND2_X1 U8907 ( .A1(n8297), .A2(n7167), .ZN(n7168) );
  OAI211_X1 U8908 ( .C1(n7170), .C2(n8306), .A(n7169), .B(n7168), .ZN(n7171)
         );
  AOI21_X1 U8909 ( .B1(n8140), .B2(n7172), .A(n7171), .ZN(n7173) );
  NAND2_X1 U8910 ( .A1(n7174), .A2(n7173), .ZN(P2_U3193) );
  INV_X1 U8911 ( .A(n7342), .ZN(n7677) );
  OAI222_X1 U8912 ( .A1(n9769), .A2(n7343), .B1(n9777), .B2(n7677), .C1(n7175), 
        .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U8913 ( .A(n7386), .ZN(n7178) );
  OAI222_X1 U8914 ( .A1(n8954), .A2(n7178), .B1(P2_U3151), .B2(n5658), .C1(
        n7176), .C2(n8951), .ZN(P2_U3270) );
  OAI222_X1 U8915 ( .A1(n9769), .A2(n8762), .B1(n9773), .B2(n7178), .C1(n7177), 
        .C2(P1_U3086), .ZN(P1_U3330) );
  NAND2_X1 U8916 ( .A1(n7895), .A2(n10229), .ZN(n7181) );
  AOI21_X1 U8917 ( .B1(n7891), .B2(n8128), .A(n7179), .ZN(n7180) );
  OAI211_X1 U8918 ( .C1(n7210), .C2(n7893), .A(n7181), .B(n7180), .ZN(n7192)
         );
  XNOR2_X1 U8919 ( .A(n7182), .B(n7778), .ZN(n7207) );
  XNOR2_X1 U8920 ( .A(n7207), .B(n8127), .ZN(n7190) );
  INV_X1 U8921 ( .A(n7183), .ZN(n7184) );
  NAND2_X1 U8922 ( .A1(n7185), .A2(n7184), .ZN(n7186) );
  INV_X1 U8923 ( .A(n7209), .ZN(n7189) );
  AOI211_X1 U8924 ( .C1(n7190), .C2(n7188), .A(n7887), .B(n7189), .ZN(n7191)
         );
  AOI211_X1 U8925 ( .C1(n10227), .C2(n7883), .A(n7192), .B(n7191), .ZN(n7193)
         );
  INV_X1 U8926 ( .A(n7193), .ZN(P2_U3171) );
  XNOR2_X1 U8927 ( .A(n7194), .B(n8029), .ZN(n7206) );
  INV_X1 U8928 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7197) );
  XOR2_X1 U8929 ( .A(n7195), .B(n8029), .Z(n7196) );
  AOI222_X1 U8930 ( .A1(n8461), .A2(n7196), .B1(n8465), .B2(n8463), .C1(n8125), 
        .C2(n8466), .ZN(n7202) );
  MUX2_X1 U8931 ( .A(n7197), .B(n7202), .S(n10275), .Z(n7199) );
  NAND2_X1 U8932 ( .A1(n8930), .A2(n7679), .ZN(n7198) );
  OAI211_X1 U8933 ( .C1(n7206), .C2(n8919), .A(n7199), .B(n7198), .ZN(P2_U3426) );
  INV_X1 U8934 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7219) );
  MUX2_X1 U8935 ( .A(n7219), .B(n7202), .S(n10289), .Z(n7201) );
  NAND2_X1 U8936 ( .A1(n7679), .A2(n8843), .ZN(n7200) );
  OAI211_X1 U8937 ( .C1(n7206), .C2(n8837), .A(n7201), .B(n7200), .ZN(P2_U3471) );
  INV_X1 U8938 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7203) );
  MUX2_X1 U8939 ( .A(n7203), .B(n7202), .S(n10233), .Z(n7205) );
  AOI22_X1 U8940 ( .A1(n7679), .A2(n10226), .B1(n10228), .B2(n7803), .ZN(n7204) );
  OAI211_X1 U8941 ( .C1(n7206), .C2(n8783), .A(n7205), .B(n7204), .ZN(P2_U3221) );
  NAND2_X1 U8942 ( .A1(n7207), .A2(n8127), .ZN(n7208) );
  XNOR2_X1 U8943 ( .A(n7765), .B(n7778), .ZN(n7760) );
  XNOR2_X1 U8944 ( .A(n7682), .B(n4574), .ZN(n7217) );
  NAND2_X1 U8945 ( .A1(n7895), .A2(n8778), .ZN(n7214) );
  AOI21_X1 U8946 ( .B1(n7891), .B2(n8126), .A(n7212), .ZN(n7213) );
  OAI211_X1 U8947 ( .C1(n8479), .C2(n7893), .A(n7214), .B(n7213), .ZN(n7215)
         );
  AOI21_X1 U8948 ( .B1(n4556), .B2(n7883), .A(n7215), .ZN(n7216) );
  OAI21_X1 U8949 ( .B1(n7217), .B2(n7887), .A(n7216), .ZN(P2_U3176) );
  INV_X1 U8950 ( .A(n7218), .ZN(n8137) );
  XNOR2_X1 U8951 ( .A(n8149), .B(n7219), .ZN(n8138) );
  AOI21_X1 U8952 ( .B1(n8139), .B2(n8137), .A(n8138), .ZN(n8142) );
  AOI21_X1 U8953 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n7233), .A(n8142), .ZN(
        n8173) );
  INV_X1 U8954 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8842) );
  AOI21_X1 U8955 ( .B1(n7220), .B2(n8842), .A(n8175), .ZN(n7241) );
  MUX2_X1 U8956 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8292), .Z(n8165) );
  XNOR2_X1 U8957 ( .A(n8165), .B(n8174), .ZN(n7227) );
  MUX2_X1 U8958 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8292), .Z(n7221) );
  OR2_X1 U8959 ( .A1(n7221), .A2(n7233), .ZN(n7225) );
  XNOR2_X1 U8960 ( .A(n7221), .B(n8149), .ZN(n8152) );
  OR2_X1 U8961 ( .A1(n7222), .A2(n4671), .ZN(n7224) );
  NAND2_X1 U8962 ( .A1(n8152), .A2(n8151), .ZN(n8150) );
  NAND2_X1 U8963 ( .A1(n7225), .A2(n8150), .ZN(n7226) );
  NAND2_X1 U8964 ( .A1(n7227), .A2(n7226), .ZN(n8166) );
  OAI21_X1 U8965 ( .B1(n7227), .B2(n7226), .A(n8166), .ZN(n7239) );
  INV_X1 U8966 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7230) );
  NAND2_X1 U8967 ( .A1(n8297), .A2(n8174), .ZN(n7229) );
  AND2_X1 U8968 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7849) );
  INV_X1 U8969 ( .A(n7849), .ZN(n7228) );
  OAI211_X1 U8970 ( .C1(n8300), .C2(n7230), .A(n7229), .B(n7228), .ZN(n7238)
         );
  INV_X1 U8971 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7235) );
  MUX2_X1 U8972 ( .A(n7203), .B(P2_REG2_REG_12__SCAN_IN), .S(n8149), .Z(n8145)
         );
  NOR2_X1 U8973 ( .A1(n7235), .A2(n7234), .ZN(n8159) );
  AOI21_X1 U8974 ( .B1(n7235), .B2(n7234), .A(n8159), .ZN(n7236) );
  NOR2_X1 U8975 ( .A1(n7236), .A2(n8306), .ZN(n7237) );
  AOI211_X1 U8976 ( .C1(n8309), .C2(n7239), .A(n7238), .B(n7237), .ZN(n7240)
         );
  OAI21_X1 U8977 ( .B1(n7241), .B2(n8310), .A(n7240), .ZN(P2_U3195) );
  INV_X1 U8978 ( .A(SI_29_), .ZN(n7245) );
  INV_X1 U8979 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8766) );
  INV_X1 U8980 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9765) );
  MUX2_X1 U8981 ( .A(n8766), .B(n9765), .S(n4443), .Z(n7247) );
  NAND2_X1 U8982 ( .A1(n7247), .A2(n8598), .ZN(n7250) );
  INV_X1 U8983 ( .A(n7247), .ZN(n7248) );
  NAND2_X1 U8984 ( .A1(n7248), .A2(SI_30_), .ZN(n7249) );
  NAND2_X1 U8985 ( .A1(n7250), .A2(n7249), .ZN(n7256) );
  MUX2_X1 U8986 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4443), .Z(n7251) );
  INV_X1 U8987 ( .A(SI_31_), .ZN(n8706) );
  XNOR2_X1 U8988 ( .A(n7251), .B(n8706), .ZN(n7252) );
  NAND2_X1 U8989 ( .A1(n8937), .A2(n7425), .ZN(n7255) );
  INV_X1 U8990 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9757) );
  OR2_X1 U8991 ( .A1(n7439), .A2(n9757), .ZN(n7254) );
  OR2_X1 U8992 ( .A1(n7439), .A2(n9765), .ZN(n7258) );
  NAND2_X1 U8993 ( .A1(n7589), .A2(n9472), .ZN(n7272) );
  OR2_X1 U8994 ( .A1(n7439), .A2(n9768), .ZN(n7260) );
  INV_X1 U8995 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9221) );
  INV_X1 U8996 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9197) );
  INV_X1 U8997 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9163) );
  INV_X1 U8998 ( .A(n7390), .ZN(n7263) );
  NAND2_X1 U8999 ( .A1(n7263), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7428) );
  INV_X1 U9000 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9087) );
  INV_X1 U9001 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9477) );
  OR2_X1 U9002 ( .A1(n7430), .A2(n9477), .ZN(n7264) );
  OR2_X1 U9003 ( .A1(n9478), .A2(n7264), .ZN(n7271) );
  INV_X1 U9004 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7268) );
  INV_X1 U9005 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8761) );
  OR2_X1 U9006 ( .A1(n7445), .A2(n8761), .ZN(n7267) );
  INV_X1 U9007 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7265) );
  OR2_X1 U9008 ( .A1(n4432), .A2(n7265), .ZN(n7266) );
  OAI211_X1 U9009 ( .C1(n7448), .C2(n7268), .A(n7267), .B(n7266), .ZN(n7269)
         );
  INV_X1 U9010 ( .A(n7269), .ZN(n7270) );
  NAND2_X1 U9011 ( .A1(n7271), .A2(n7270), .ZN(n9270) );
  INV_X1 U9012 ( .A(n9270), .ZN(n7453) );
  NAND2_X1 U9013 ( .A1(n7272), .A2(n7583), .ZN(n7651) );
  NAND2_X1 U9014 ( .A1(n7273), .A2(n7425), .ZN(n7275) );
  AOI22_X1 U9015 ( .A1(n7339), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7338), .B2(
        n9907), .ZN(n7274) );
  INV_X1 U9016 ( .A(n9417), .ZN(n7276) );
  OR2_X1 U9017 ( .A1(n9984), .A2(n7276), .ZN(n7526) );
  NAND2_X1 U9018 ( .A1(n9984), .A2(n7276), .ZN(n7529) );
  INV_X1 U9019 ( .A(n9982), .ZN(n9973) );
  INV_X1 U9020 ( .A(n7519), .ZN(n9974) );
  NOR2_X1 U9021 ( .A1(n9973), .A2(n9974), .ZN(n7277) );
  NAND2_X1 U9022 ( .A1(n7279), .A2(n7425), .ZN(n7281) );
  AOI22_X1 U9023 ( .A1(n7339), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7338), .B2(
        n9911), .ZN(n7280) );
  INV_X1 U9024 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9670) );
  INV_X1 U9025 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9357) );
  OR2_X1 U9026 ( .A1(n7445), .A2(n9357), .ZN(n7282) );
  OAI21_X1 U9027 ( .B1(n7448), .B2(n9670), .A(n7282), .ZN(n7286) );
  INV_X1 U9028 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9097) );
  XNOR2_X1 U9029 ( .A(n7292), .B(n9097), .ZN(n9669) );
  INV_X1 U9030 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7283) );
  OR2_X1 U9031 ( .A1(n4432), .A2(n7283), .ZN(n7284) );
  OAI21_X1 U9032 ( .B1(n7319), .B2(n9669), .A(n7284), .ZN(n7285) );
  NAND2_X1 U9033 ( .A1(n10195), .A2(n9418), .ZN(n7531) );
  NAND2_X1 U9034 ( .A1(n9674), .A2(n9419), .ZN(n7624) );
  NAND2_X1 U9035 ( .A1(n7531), .A2(n7624), .ZN(n9662) );
  INV_X1 U9036 ( .A(n7529), .ZN(n9663) );
  NOR2_X1 U9037 ( .A1(n9662), .A2(n9663), .ZN(n7287) );
  NAND2_X1 U9038 ( .A1(n9976), .A2(n7287), .ZN(n9665) );
  NAND2_X1 U9039 ( .A1(n7288), .A2(n7425), .ZN(n7290) );
  AOI22_X1 U9040 ( .A1(n7339), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7338), .B2(
        n9935), .ZN(n7289) );
  INV_X1 U9041 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7291) );
  OAI21_X1 U9042 ( .B1(n7292), .B2(n9097), .A(n7291), .ZN(n7294) );
  INV_X1 U9043 ( .A(n7293), .ZN(n7308) );
  NAND2_X1 U9044 ( .A1(n7294), .A2(n7308), .ZN(n9838) );
  OR2_X1 U9045 ( .A1(n7430), .A2(n9838), .ZN(n7302) );
  INV_X1 U9046 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7295) );
  OR2_X1 U9047 ( .A1(n7296), .A2(n7295), .ZN(n7301) );
  INV_X1 U9048 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7297) );
  OR2_X1 U9049 ( .A1(n4432), .A2(n7297), .ZN(n7300) );
  INV_X1 U9050 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7298) );
  OR2_X1 U9051 ( .A1(n7445), .A2(n7298), .ZN(n7299) );
  NAND4_X1 U9052 ( .A1(n7302), .A2(n7301), .A3(n7300), .A4(n7299), .ZN(n9421)
         );
  INV_X1 U9053 ( .A(n9421), .ZN(n9422) );
  OR2_X1 U9054 ( .A1(n4438), .A2(n9422), .ZN(n7534) );
  NAND2_X1 U9055 ( .A1(n4437), .A2(n9422), .ZN(n7625) );
  NAND2_X1 U9056 ( .A1(n7534), .A2(n7625), .ZN(n9841) );
  NAND2_X1 U9057 ( .A1(n7303), .A2(n7425), .ZN(n7305) );
  AOI22_X1 U9058 ( .A1(n7339), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7338), .B2(
        n9939), .ZN(n7304) );
  INV_X1 U9059 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9653) );
  INV_X1 U9060 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7306) );
  OR2_X1 U9061 ( .A1(n7445), .A2(n7306), .ZN(n7307) );
  OAI21_X1 U9062 ( .B1(n7448), .B2(n9653), .A(n7307), .ZN(n7313) );
  INV_X1 U9063 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8645) );
  NAND2_X1 U9064 ( .A1(n7308), .A2(n8645), .ZN(n7309) );
  NAND2_X1 U9065 ( .A1(n7329), .A2(n7309), .ZN(n9652) );
  INV_X1 U9066 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7310) );
  OR2_X1 U9067 ( .A1(n4431), .A2(n7310), .ZN(n7311) );
  OAI21_X1 U9068 ( .B1(n7319), .B2(n9652), .A(n7311), .ZN(n7312) );
  NAND2_X1 U9069 ( .A1(n4578), .A2(n9423), .ZN(n7632) );
  NAND2_X1 U9070 ( .A1(n7535), .A2(n7632), .ZN(n9649) );
  INV_X1 U9071 ( .A(n9649), .ZN(n9646) );
  NAND2_X1 U9072 ( .A1(n9644), .A2(n7632), .ZN(n9819) );
  NAND2_X1 U9073 ( .A1(n7314), .A2(n7425), .ZN(n7316) );
  AOI22_X1 U9074 ( .A1(n7339), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7338), .B2(
        n9389), .ZN(n7315) );
  INV_X1 U9075 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9185) );
  XNOR2_X1 U9076 ( .A(n7329), .B(n9185), .ZN(n9823) );
  INV_X1 U9077 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7317) );
  OR2_X1 U9078 ( .A1(n7445), .A2(n7317), .ZN(n7318) );
  OAI21_X1 U9079 ( .B1(n7319), .B2(n9823), .A(n7318), .ZN(n7324) );
  INV_X1 U9080 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7322) );
  INV_X1 U9081 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n7320) );
  OR2_X1 U9082 ( .A1(n4431), .A2(n7320), .ZN(n7321) );
  OAI21_X1 U9083 ( .B1(n7448), .B2(n7322), .A(n7321), .ZN(n7323) );
  NAND2_X1 U9084 ( .A1(n9825), .A2(n9427), .ZN(n7541) );
  NAND2_X1 U9085 ( .A1(n7631), .A2(n7541), .ZN(n9818) );
  NAND2_X1 U9086 ( .A1(n7325), .A2(n7425), .ZN(n7327) );
  AOI22_X1 U9087 ( .A1(n7339), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7338), .B2(
        n9968), .ZN(n7326) );
  INV_X1 U9088 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7328) );
  OAI21_X1 U9089 ( .B1(n7329), .B2(n9185), .A(n7328), .ZN(n7331) );
  NAND2_X1 U9090 ( .A1(n7331), .A2(n7330), .ZN(n9636) );
  OR2_X1 U9091 ( .A1(n7430), .A2(n9636), .ZN(n7336) );
  INV_X1 U9092 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9637) );
  OR2_X1 U9093 ( .A1(n7448), .A2(n9637), .ZN(n7335) );
  INV_X1 U9094 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9385) );
  OR2_X1 U9095 ( .A1(n7445), .A2(n9385), .ZN(n7334) );
  INV_X1 U9096 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n7332) );
  OR2_X1 U9097 ( .A1(n4432), .A2(n7332), .ZN(n7333) );
  NAND4_X1 U9098 ( .A1(n7336), .A2(n7335), .A3(n7334), .A4(n7333), .ZN(n9429)
         );
  INV_X1 U9099 ( .A(n9429), .ZN(n9428) );
  OR2_X1 U9100 ( .A1(n9641), .A2(n9428), .ZN(n7634) );
  NAND2_X1 U9101 ( .A1(n9641), .A2(n9428), .ZN(n7542) );
  NAND2_X1 U9102 ( .A1(n7634), .A2(n7542), .ZN(n9635) );
  NAND2_X1 U9103 ( .A1(n7337), .A2(n7425), .ZN(n7341) );
  AOI22_X1 U9104 ( .A1(n7339), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4434), .B2(
        n7338), .ZN(n7340) );
  INV_X1 U9105 ( .A(n9431), .ZN(n9432) );
  OR2_X1 U9106 ( .A1(n9737), .A2(n9432), .ZN(n7635) );
  NAND2_X1 U9107 ( .A1(n9737), .A2(n9432), .ZN(n7640) );
  INV_X1 U9108 ( .A(n7640), .ZN(n7550) );
  NAND2_X1 U9109 ( .A1(n7342), .A2(n7425), .ZN(n7345) );
  OR2_X1 U9110 ( .A1(n7439), .A2(n7343), .ZN(n7344) );
  XNOR2_X1 U9111 ( .A(n7389), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9553) );
  NAND2_X1 U9112 ( .A1(n9553), .A2(n7450), .ZN(n7353) );
  INV_X1 U9113 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n7350) );
  INV_X1 U9114 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n7346) );
  OR2_X1 U9115 ( .A1(n4432), .A2(n7346), .ZN(n7349) );
  INV_X1 U9116 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7347) );
  OR2_X1 U9117 ( .A1(n7445), .A2(n7347), .ZN(n7348) );
  OAI211_X1 U9118 ( .C1(n7448), .C2(n7350), .A(n7349), .B(n7348), .ZN(n7351)
         );
  INV_X1 U9119 ( .A(n7351), .ZN(n7352) );
  NAND2_X1 U9120 ( .A1(n7353), .A2(n7352), .ZN(n9272) );
  NAND2_X1 U9121 ( .A1(n9713), .A2(n9447), .ZN(n7566) );
  NAND2_X1 U9122 ( .A1(n7354), .A2(n7425), .ZN(n7357) );
  OR2_X1 U9123 ( .A1(n7439), .A2(n7355), .ZN(n7356) );
  INV_X1 U9124 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n7363) );
  INV_X1 U9125 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9107) );
  NAND2_X1 U9126 ( .A1(n7369), .A2(n9107), .ZN(n7358) );
  NAND2_X1 U9127 ( .A1(n7389), .A2(n7358), .ZN(n9561) );
  OR2_X1 U9128 ( .A1(n9561), .A2(n7430), .ZN(n7362) );
  INV_X1 U9129 ( .A(n7445), .ZN(n7359) );
  AOI22_X1 U9130 ( .A1(n7360), .A2(P1_REG0_REG_23__SCAN_IN), .B1(n7359), .B2(
        P1_REG1_REG_23__SCAN_IN), .ZN(n7361) );
  OAI211_X1 U9131 ( .C1(n7448), .C2(n7363), .A(n7362), .B(n7361), .ZN(n9443)
         );
  INV_X1 U9132 ( .A(n9443), .ZN(n9444) );
  OR2_X1 U9133 ( .A1(n9717), .A2(n9444), .ZN(n7459) );
  INV_X1 U9134 ( .A(n7459), .ZN(n7563) );
  NAND2_X1 U9135 ( .A1(n7364), .A2(n7425), .ZN(n7367) );
  OR2_X1 U9136 ( .A1(n7439), .A2(n7365), .ZN(n7366) );
  NAND2_X1 U9137 ( .A1(n7407), .A2(n9221), .ZN(n7368) );
  NAND2_X1 U9138 ( .A1(n7369), .A2(n7368), .ZN(n9576) );
  INV_X1 U9139 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9577) );
  INV_X1 U9140 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7370) );
  OR2_X1 U9141 ( .A1(n7445), .A2(n7370), .ZN(n7371) );
  OAI21_X1 U9142 ( .B1(n7448), .B2(n9577), .A(n7371), .ZN(n7372) );
  INV_X1 U9143 ( .A(n7372), .ZN(n7375) );
  INV_X1 U9144 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n7373) );
  OR2_X1 U9145 ( .A1(n4431), .A2(n7373), .ZN(n7374) );
  OAI211_X1 U9146 ( .C1(n9576), .C2(n7430), .A(n7375), .B(n7374), .ZN(n9442)
         );
  INV_X1 U9147 ( .A(n9442), .ZN(n9441) );
  OR2_X1 U9148 ( .A1(n9723), .A2(n9441), .ZN(n7461) );
  INV_X1 U9149 ( .A(n7461), .ZN(n9463) );
  NOR2_X1 U9150 ( .A1(n7563), .A2(n9463), .ZN(n7562) );
  NAND2_X1 U9151 ( .A1(n9717), .A2(n9444), .ZN(n9464) );
  OAI21_X1 U9152 ( .B1(n7562), .B2(n4845), .A(n9465), .ZN(n7400) );
  NAND2_X1 U9153 ( .A1(n8952), .A2(n7425), .ZN(n7377) );
  OR2_X1 U9154 ( .A1(n7439), .A2(n9778), .ZN(n7376) );
  NAND2_X2 U9155 ( .A1(n7377), .A2(n7376), .ZN(n9703) );
  INV_X1 U9156 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U9157 ( .A1(n7390), .A2(n9254), .ZN(n7378) );
  NAND2_X1 U9158 ( .A1(n7428), .A2(n7378), .ZN(n9521) );
  OR2_X1 U9159 ( .A1(n9521), .A2(n7430), .ZN(n7385) );
  INV_X1 U9160 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9520) );
  INV_X1 U9161 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7379) );
  OR2_X1 U9162 ( .A1(n7445), .A2(n7379), .ZN(n7382) );
  INV_X1 U9163 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n7380) );
  OR2_X1 U9164 ( .A1(n4431), .A2(n7380), .ZN(n7381) );
  OAI211_X1 U9165 ( .C1(n7448), .C2(n9520), .A(n7382), .B(n7381), .ZN(n7383)
         );
  INV_X1 U9166 ( .A(n7383), .ZN(n7384) );
  NAND2_X1 U9167 ( .A1(n7385), .A2(n7384), .ZN(n9271) );
  NAND2_X1 U9168 ( .A1(n7386), .A2(n7425), .ZN(n7388) );
  OR2_X1 U9169 ( .A1(n7439), .A2(n8762), .ZN(n7387) );
  OAI21_X1 U9170 ( .B1(n7389), .B2(n9197), .A(n9163), .ZN(n7391) );
  AND2_X1 U9171 ( .A1(n7391), .A2(n7390), .ZN(n9534) );
  NAND2_X1 U9172 ( .A1(n9534), .A2(n7450), .ZN(n7399) );
  INV_X1 U9173 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n7396) );
  INV_X1 U9174 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7392) );
  OR2_X1 U9175 ( .A1(n7445), .A2(n7392), .ZN(n7395) );
  INV_X1 U9176 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n7393) );
  OR2_X1 U9177 ( .A1(n4432), .A2(n7393), .ZN(n7394) );
  OAI211_X1 U9178 ( .C1(n7448), .C2(n7396), .A(n7395), .B(n7394), .ZN(n7397)
         );
  INV_X1 U9179 ( .A(n7397), .ZN(n7398) );
  NAND2_X1 U9180 ( .A1(n7399), .A2(n7398), .ZN(n9451) );
  INV_X1 U9181 ( .A(n9451), .ZN(n9057) );
  OR2_X1 U9182 ( .A1(n9707), .A2(n9057), .ZN(n9466) );
  NAND2_X1 U9183 ( .A1(n7458), .A2(n9466), .ZN(n7574) );
  NAND2_X1 U9184 ( .A1(n7401), .A2(n7425), .ZN(n7404) );
  OR2_X1 U9185 ( .A1(n7439), .A2(n7402), .ZN(n7403) );
  INV_X1 U9186 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U9187 ( .A1(n7405), .A2(n9145), .ZN(n7406) );
  NAND2_X1 U9188 ( .A1(n7407), .A2(n7406), .ZN(n9144) );
  OR2_X1 U9189 ( .A1(n7430), .A2(n9144), .ZN(n7414) );
  INV_X1 U9190 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n7408) );
  OR2_X1 U9191 ( .A1(n7448), .A2(n7408), .ZN(n7413) );
  INV_X1 U9192 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n7409) );
  OR2_X1 U9193 ( .A1(n7445), .A2(n7409), .ZN(n7412) );
  INV_X1 U9194 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n7410) );
  OR2_X1 U9195 ( .A1(n4431), .A2(n7410), .ZN(n7411) );
  NAND4_X1 U9196 ( .A1(n7414), .A2(n7413), .A3(n7412), .A4(n7411), .ZN(n9438)
         );
  INV_X1 U9197 ( .A(n9438), .ZN(n9437) );
  OR2_X1 U9198 ( .A1(n9728), .A2(n9437), .ZN(n7543) );
  OR2_X1 U9199 ( .A1(n7439), .A2(n7416), .ZN(n7417) );
  INV_X1 U9200 ( .A(n9435), .ZN(n9434) );
  NAND2_X1 U9201 ( .A1(n7543), .A2(n7545), .ZN(n9461) );
  INV_X1 U9202 ( .A(n9461), .ZN(n7419) );
  NAND2_X1 U9203 ( .A1(n7424), .A2(n7419), .ZN(n7638) );
  NAND2_X1 U9204 ( .A1(n9723), .A2(n9441), .ZN(n7460) );
  NAND2_X1 U9205 ( .A1(n9464), .A2(n7460), .ZN(n7560) );
  INV_X1 U9206 ( .A(n7560), .ZN(n7421) );
  NAND2_X1 U9207 ( .A1(n9728), .A2(n9437), .ZN(n7559) );
  NAND2_X1 U9208 ( .A1(n9733), .A2(n9434), .ZN(n7546) );
  NAND2_X1 U9209 ( .A1(n7559), .A2(n7546), .ZN(n7420) );
  NAND2_X1 U9210 ( .A1(n7420), .A2(n7543), .ZN(n9460) );
  NAND3_X1 U9211 ( .A1(n7566), .A2(n7421), .A3(n9460), .ZN(n7423) );
  INV_X1 U9212 ( .A(n7458), .ZN(n7568) );
  NAND2_X1 U9213 ( .A1(n9707), .A2(n9057), .ZN(n7575) );
  NAND2_X1 U9214 ( .A1(n9703), .A2(n9454), .ZN(n7577) );
  OAI21_X1 U9215 ( .B1(n7568), .B2(n7575), .A(n7577), .ZN(n7422) );
  AOI21_X1 U9216 ( .B1(n7424), .B2(n7423), .A(n7422), .ZN(n7641) );
  OAI21_X1 U9217 ( .B1(n9604), .B2(n7638), .A(n7641), .ZN(n7452) );
  NAND2_X1 U9218 ( .A1(n8947), .A2(n7425), .ZN(n7427) );
  OR2_X1 U9219 ( .A1(n7439), .A2(n8764), .ZN(n7426) );
  NAND2_X1 U9220 ( .A1(n7428), .A2(n9087), .ZN(n7429) );
  NAND2_X1 U9221 ( .A1(n9478), .A2(n7429), .ZN(n9504) );
  OR2_X1 U9222 ( .A1(n9504), .A2(n7430), .ZN(n7438) );
  INV_X1 U9223 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n7435) );
  INV_X1 U9224 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n7431) );
  OR2_X1 U9225 ( .A1(n4431), .A2(n7431), .ZN(n7434) );
  INV_X1 U9226 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7432) );
  OR2_X1 U9227 ( .A1(n7445), .A2(n7432), .ZN(n7433) );
  OAI211_X1 U9228 ( .C1(n7448), .C2(n7435), .A(n7434), .B(n7433), .ZN(n7436)
         );
  INV_X1 U9229 ( .A(n7436), .ZN(n7437) );
  INV_X1 U9230 ( .A(n9456), .ZN(n7451) );
  NAND2_X1 U9231 ( .A1(n9770), .A2(n7425), .ZN(n7441) );
  OR2_X1 U9232 ( .A1(n7439), .A2(n9771), .ZN(n7440) );
  NAND2_X2 U9233 ( .A1(n7441), .A2(n7440), .ZN(n9692) );
  XNOR2_X1 U9234 ( .A(n9478), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9497) );
  INV_X1 U9235 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9489) );
  INV_X1 U9236 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7442) );
  OR2_X1 U9237 ( .A1(n4432), .A2(n7442), .ZN(n7447) );
  INV_X1 U9238 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7444) );
  OR2_X1 U9239 ( .A1(n7445), .A2(n7444), .ZN(n7446) );
  OAI211_X1 U9240 ( .C1(n7448), .C2(n9489), .A(n7447), .B(n7446), .ZN(n7449)
         );
  AOI21_X1 U9241 ( .B1(n9497), .B2(n7450), .A(n7449), .ZN(n9474) );
  NAND2_X1 U9242 ( .A1(n9692), .A2(n9474), .ZN(n9469) );
  NAND2_X1 U9243 ( .A1(n9469), .A2(n9468), .ZN(n7645) );
  AOI21_X1 U9244 ( .B1(n7452), .B2(n7642), .A(n7645), .ZN(n7454) );
  NAND2_X1 U9245 ( .A1(n7582), .A2(n7486), .ZN(n7646) );
  NOR2_X1 U9246 ( .A1(n7454), .A2(n7646), .ZN(n7455) );
  AOI211_X1 U9247 ( .C1(n9678), .C2(n7589), .A(n7651), .B(n7455), .ZN(n7457)
         );
  NOR2_X1 U9248 ( .A1(n7589), .A2(n9472), .ZN(n7649) );
  INV_X1 U9249 ( .A(n7588), .ZN(n9407) );
  INV_X1 U9250 ( .A(n7596), .ZN(n7456) );
  OAI21_X1 U9251 ( .B1(n7457), .B2(n7456), .A(n7654), .ZN(n7484) );
  NAND2_X1 U9252 ( .A1(n7458), .A2(n7577), .ZN(n9526) );
  NAND2_X1 U9253 ( .A1(n7461), .A2(n7460), .ZN(n9462) );
  NAND2_X1 U9254 ( .A1(n7545), .A2(n7546), .ZN(n9601) );
  INV_X1 U9255 ( .A(n9623), .ZN(n7478) );
  INV_X1 U9256 ( .A(n9818), .ZN(n9826) );
  INV_X1 U9257 ( .A(n7462), .ZN(n7471) );
  INV_X1 U9258 ( .A(n7463), .ZN(n7470) );
  INV_X1 U9259 ( .A(n10061), .ZN(n7465) );
  INV_X1 U9260 ( .A(n7464), .ZN(n10071) );
  NAND2_X1 U9261 ( .A1(n6285), .A2(n10082), .ZN(n7607) );
  NAND2_X1 U9262 ( .A1(n10071), .A2(n7607), .ZN(n10111) );
  NOR4_X1 U9263 ( .A1(n7465), .A2(n7599), .A3(n10111), .A4(n7490), .ZN(n7467)
         );
  NAND4_X1 U9264 ( .A1(n7467), .A2(n10048), .A3(n10070), .A4(n7466), .ZN(n7468) );
  NOR4_X1 U9265 ( .A1(n7471), .A2(n7470), .A3(n7469), .A4(n7468), .ZN(n7472)
         );
  NAND4_X1 U9266 ( .A1(n7474), .A2(n9995), .A3(n7473), .A4(n7472), .ZN(n7475)
         );
  NOR4_X1 U9267 ( .A1(n9841), .A2(n9973), .A3(n9662), .A4(n7475), .ZN(n7476)
         );
  NAND3_X1 U9268 ( .A1(n9826), .A2(n9646), .A3(n7476), .ZN(n7477) );
  NOR4_X1 U9269 ( .A1(n9601), .A2(n7478), .A3(n9635), .A4(n7477), .ZN(n7479)
         );
  XNOR2_X1 U9270 ( .A(n9728), .B(n9438), .ZN(n9591) );
  NAND4_X1 U9271 ( .A1(n9566), .A2(n9581), .A3(n7479), .A4(n9591), .ZN(n7480)
         );
  NAND2_X1 U9272 ( .A1(n9466), .A2(n7575), .ZN(n9538) );
  NAND2_X1 U9273 ( .A1(n9465), .A2(n7566), .ZN(n9544) );
  NAND2_X1 U9274 ( .A1(n7593), .A2(n9407), .ZN(n7653) );
  XOR2_X1 U9275 ( .A(n9472), .B(n7589), .Z(n7482) );
  NAND4_X1 U9276 ( .A1(n7483), .A2(n7654), .A3(n7653), .A4(n7482), .ZN(n7597)
         );
  NAND2_X1 U9277 ( .A1(n7486), .A2(n7642), .ZN(n7578) );
  OAI211_X1 U9278 ( .C1(n7578), .C2(n9468), .A(n9469), .B(n4734), .ZN(n7572)
         );
  OAI211_X1 U9279 ( .C1(n7645), .C2(n7642), .A(n7600), .B(n7486), .ZN(n7571)
         );
  INV_X1 U9280 ( .A(n7625), .ZN(n7487) );
  NAND2_X1 U9281 ( .A1(n7535), .A2(n7487), .ZN(n7488) );
  OAI211_X1 U9282 ( .C1(n4437), .C2(n4734), .A(n7488), .B(n7632), .ZN(n7540)
         );
  INV_X1 U9283 ( .A(n7632), .ZN(n7489) );
  OAI21_X1 U9284 ( .B1(n7489), .B2(n9422), .A(n7600), .ZN(n7539) );
  NOR2_X1 U9285 ( .A1(n7491), .A2(n7490), .ZN(n7493) );
  OAI211_X1 U9286 ( .C1(n7500), .C2(n7615), .A(n7502), .B(n7497), .ZN(n7495)
         );
  NAND2_X1 U9287 ( .A1(n7495), .A2(n7494), .ZN(n7505) );
  NAND2_X1 U9288 ( .A1(n7497), .A2(n7496), .ZN(n7499) );
  INV_X1 U9289 ( .A(n7615), .ZN(n7498) );
  OAI21_X1 U9290 ( .B1(n7500), .B2(n7499), .A(n7498), .ZN(n7503) );
  AOI21_X1 U9291 ( .B1(n7503), .B2(n7502), .A(n7501), .ZN(n7504) );
  INV_X1 U9292 ( .A(n7507), .ZN(n7521) );
  NAND3_X1 U9293 ( .A1(n7509), .A2(n7508), .A3(n7521), .ZN(n7514) );
  OAI21_X1 U9294 ( .B1(n7512), .B2(n7511), .A(n7510), .ZN(n7513) );
  NAND3_X1 U9295 ( .A1(n7522), .A2(n7617), .A3(n7515), .ZN(n7520) );
  NAND2_X1 U9296 ( .A1(n7517), .A2(n7516), .ZN(n7523) );
  INV_X1 U9297 ( .A(n7523), .ZN(n7620) );
  NAND2_X1 U9298 ( .A1(n7519), .A2(n7518), .ZN(n7619) );
  INV_X1 U9299 ( .A(n7525), .ZN(n7622) );
  NAND2_X1 U9300 ( .A1(n7522), .A2(n7521), .ZN(n7524) );
  AND2_X1 U9301 ( .A1(n7531), .A2(n7526), .ZN(n7532) );
  INV_X1 U9302 ( .A(n7532), .ZN(n7626) );
  AOI21_X1 U9303 ( .B1(n7533), .B2(n7529), .A(n7626), .ZN(n7528) );
  NAND3_X1 U9304 ( .A1(n7632), .A2(n7625), .A3(n7624), .ZN(n7527) );
  OAI21_X1 U9305 ( .B1(n7528), .B2(n7527), .A(n7535), .ZN(n7538) );
  NAND2_X1 U9306 ( .A1(n7624), .A2(n7529), .ZN(n7530) );
  NAND2_X1 U9307 ( .A1(n7535), .A2(n7534), .ZN(n7628) );
  NOR2_X1 U9308 ( .A1(n7536), .A2(n7628), .ZN(n7537) );
  NAND2_X1 U9309 ( .A1(n7542), .A2(n7541), .ZN(n7636) );
  OAI21_X1 U9310 ( .B1(n7631), .B2(n4734), .A(n7634), .ZN(n7544) );
  INV_X1 U9311 ( .A(n7543), .ZN(n7553) );
  AOI211_X1 U9312 ( .C1(n4734), .C2(n7636), .A(n7544), .B(n7553), .ZN(n7549)
         );
  INV_X1 U9313 ( .A(n7546), .ZN(n7548) );
  INV_X1 U9314 ( .A(n7635), .ZN(n7547) );
  INV_X1 U9315 ( .A(n9737), .ZN(n9622) );
  OAI21_X1 U9316 ( .B1(n9429), .B2(n4734), .A(n9641), .ZN(n7552) );
  OAI21_X1 U9317 ( .B1(n9428), .B2(n7600), .A(n9851), .ZN(n7551) );
  AOI21_X1 U9318 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(n7554) );
  AOI21_X1 U9319 ( .B1(n7554), .B2(n7635), .A(n7553), .ZN(n7555) );
  AOI22_X1 U9320 ( .A1(n7556), .A2(n7555), .B1(n9461), .B2(n4734), .ZN(n7557)
         );
  OAI21_X1 U9321 ( .B1(n7600), .B2(n7559), .A(n7558), .ZN(n7561) );
  AOI22_X1 U9322 ( .A1(n7561), .A2(n9581), .B1(n7560), .B2(n4734), .ZN(n7564)
         );
  OAI22_X1 U9323 ( .A1(n7564), .A2(n7563), .B1(n7562), .B2(n4734), .ZN(n7565)
         );
  INV_X1 U9324 ( .A(n9544), .ZN(n9546) );
  MUX2_X1 U9325 ( .A(n9465), .B(n7566), .S(n4734), .Z(n7567) );
  NOR2_X1 U9326 ( .A1(n7573), .A2(n7574), .ZN(n7570) );
  AOI21_X1 U9327 ( .B1(n7577), .B2(n7575), .A(n7568), .ZN(n7569) );
  INV_X1 U9328 ( .A(n7573), .ZN(n7576) );
  AOI21_X1 U9329 ( .B1(n7576), .B2(n7575), .A(n7574), .ZN(n7580) );
  INV_X1 U9330 ( .A(n7577), .ZN(n9467) );
  INV_X1 U9331 ( .A(n7578), .ZN(n7579) );
  OAI211_X1 U9332 ( .C1(n7580), .C2(n9467), .A(n7579), .B(n4734), .ZN(n7586)
         );
  NOR2_X1 U9333 ( .A1(n9472), .A2(n4734), .ZN(n7581) );
  AND2_X1 U9334 ( .A1(n7581), .A2(n7588), .ZN(n7587) );
  NAND3_X1 U9335 ( .A1(n9684), .A2(n7600), .A3(n7583), .ZN(n7584) );
  AOI21_X1 U9336 ( .B1(n7589), .B2(n4734), .A(n7588), .ZN(n7594) );
  INV_X1 U9337 ( .A(n7587), .ZN(n7591) );
  NAND3_X1 U9338 ( .A1(n9472), .A2(n7588), .A3(n4734), .ZN(n7590) );
  MUX2_X1 U9339 ( .A(n7591), .B(n7590), .S(n7589), .Z(n7592) );
  OAI21_X1 U9340 ( .B1(n7594), .B2(n7593), .A(n7592), .ZN(n7595) );
  OAI21_X1 U9341 ( .B1(n7603), .B2(n4922), .A(n7597), .ZN(n7598) );
  NAND2_X1 U9342 ( .A1(n7602), .A2(n7601), .ZN(n7662) );
  OAI21_X1 U9343 ( .B1(n7653), .B2(n4734), .A(n7603), .ZN(n7660) );
  INV_X1 U9344 ( .A(n7654), .ZN(n7605) );
  AOI211_X1 U9345 ( .C1(n7605), .C2(n4434), .A(n4433), .B(n7604), .ZN(n7659)
         );
  INV_X1 U9346 ( .A(n4440), .ZN(n10118) );
  NAND2_X1 U9347 ( .A1(n9283), .A2(n10118), .ZN(n7606) );
  AND2_X1 U9348 ( .A1(n7607), .A2(n7606), .ZN(n7611) );
  AOI21_X1 U9349 ( .B1(n9282), .B2(n10124), .A(n4922), .ZN(n7610) );
  NAND4_X1 U9350 ( .A1(n7611), .A2(n7610), .A3(n7609), .A4(n7608), .ZN(n7614)
         );
  INV_X1 U9351 ( .A(n7612), .ZN(n7613) );
  OAI21_X1 U9352 ( .B1(n7615), .B2(n7614), .A(n7613), .ZN(n7618) );
  NAND3_X1 U9353 ( .A1(n7618), .A2(n7617), .A3(n7616), .ZN(n7621) );
  AOI21_X1 U9354 ( .B1(n7621), .B2(n7620), .A(n7619), .ZN(n7623) );
  NOR3_X1 U9355 ( .A1(n7623), .A2(n9663), .A3(n7622), .ZN(n7627) );
  OAI211_X1 U9356 ( .C1(n7627), .C2(n7626), .A(n7625), .B(n7624), .ZN(n7630)
         );
  INV_X1 U9357 ( .A(n7628), .ZN(n7629) );
  NAND2_X1 U9358 ( .A1(n7630), .A2(n7629), .ZN(n7633) );
  AOI21_X1 U9359 ( .B1(n7633), .B2(n7632), .A(n4838), .ZN(n7637) );
  OAI211_X1 U9360 ( .C1(n7637), .C2(n7636), .A(n7635), .B(n7634), .ZN(n7639)
         );
  INV_X1 U9361 ( .A(n7641), .ZN(n7643) );
  OAI21_X1 U9362 ( .B1(n7644), .B2(n7643), .A(n7642), .ZN(n7648) );
  INV_X1 U9363 ( .A(n7645), .ZN(n7647) );
  INV_X1 U9364 ( .A(n7649), .ZN(n7650) );
  OAI21_X1 U9365 ( .B1(n7652), .B2(n7651), .A(n7650), .ZN(n7656) );
  INV_X1 U9366 ( .A(n7653), .ZN(n7655) );
  NOR3_X1 U9367 ( .A1(n7664), .A2(n9404), .A3(n9475), .ZN(n7666) );
  OAI21_X1 U9368 ( .B1(n7667), .B2(n4433), .A(P1_B_REG_SCAN_IN), .ZN(n7665) );
  INV_X1 U9369 ( .A(n8947), .ZN(n7668) );
  OAI222_X1 U9370 ( .A1(n9769), .A2(n8764), .B1(n9777), .B2(n7668), .C1(n9404), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  NAND2_X1 U9371 ( .A1(n7670), .A2(n10228), .ZN(n8313) );
  NAND2_X1 U9372 ( .A1(n8489), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7671) );
  OAI211_X1 U9373 ( .C1(n7672), .C2(n8431), .A(n8313), .B(n7671), .ZN(n7673)
         );
  AOI21_X1 U9374 ( .B1(n5762), .B2(n7674), .A(n7673), .ZN(n7675) );
  OAI21_X1 U9375 ( .B1(n7669), .B2(n8489), .A(n7675), .ZN(P2_U3204) );
  OAI222_X1 U9376 ( .A1(n8954), .A2(n7677), .B1(P2_U3151), .B2(n5653), .C1(
        n7676), .C2(n8951), .ZN(P2_U3271) );
  INV_X1 U9377 ( .A(n7901), .ZN(n9764) );
  OAI222_X1 U9378 ( .A1(n8951), .A2(n8766), .B1(n8954), .B2(n9764), .C1(
        P2_U3151), .C2(n7678), .ZN(P2_U3265) );
  XNOR2_X1 U9379 ( .A(n8826), .B(n7778), .ZN(n7827) );
  INV_X1 U9380 ( .A(n7827), .ZN(n7696) );
  XNOR2_X1 U9381 ( .A(n8916), .B(n7778), .ZN(n7691) );
  INV_X1 U9382 ( .A(n7691), .ZN(n7692) );
  XNOR2_X1 U9383 ( .A(n8923), .B(n7778), .ZN(n7688) );
  XNOR2_X1 U9384 ( .A(n8929), .B(n7705), .ZN(n7737) );
  INV_X1 U9385 ( .A(n7682), .ZN(n7733) );
  XNOR2_X1 U9386 ( .A(n7679), .B(n7778), .ZN(n7735) );
  OAI211_X1 U9387 ( .C1(n7737), .C2(n8465), .A(n7733), .B(n7736), .ZN(n7690)
         );
  NAND3_X1 U9388 ( .A1(n7736), .A2(n8125), .A3(n7682), .ZN(n7681) );
  INV_X1 U9389 ( .A(n7735), .ZN(n7683) );
  AOI21_X1 U9390 ( .B1(n7683), .B2(n8124), .A(n8465), .ZN(n7680) );
  NAND2_X1 U9391 ( .A1(n7681), .A2(n7680), .ZN(n7687) );
  NAND4_X1 U9392 ( .A1(n7736), .A2(n8465), .A3(n8125), .A4(n7682), .ZN(n7685)
         );
  NAND3_X1 U9393 ( .A1(n7683), .A2(n8465), .A3(n8124), .ZN(n7684) );
  NAND2_X1 U9394 ( .A1(n7685), .A2(n7684), .ZN(n7686) );
  XNOR2_X1 U9395 ( .A(n7688), .B(n8451), .ZN(n7739) );
  XNOR2_X1 U9396 ( .A(n7691), .B(n7743), .ZN(n7889) );
  XNOR2_X1 U9397 ( .A(n8830), .B(n7778), .ZN(n7815) );
  NAND2_X1 U9398 ( .A1(n7817), .A2(n7693), .ZN(n7695) );
  NAND2_X1 U9399 ( .A1(n7695), .A2(n7694), .ZN(n7825) );
  XNOR2_X1 U9400 ( .A(n8903), .B(n7705), .ZN(n7697) );
  NOR2_X1 U9401 ( .A1(n7697), .A2(n8405), .ZN(n7698) );
  AOI21_X1 U9402 ( .B1(n7697), .B2(n8405), .A(n7698), .ZN(n7870) );
  XNOR2_X1 U9403 ( .A(n8819), .B(n7705), .ZN(n7767) );
  NAND2_X1 U9404 ( .A1(n7767), .A2(n8415), .ZN(n7700) );
  INV_X1 U9405 ( .A(n7767), .ZN(n7699) );
  XNOR2_X1 U9406 ( .A(n8896), .B(n7778), .ZN(n7701) );
  XNOR2_X1 U9407 ( .A(n7701), .B(n7791), .ZN(n7843) );
  XNOR2_X1 U9408 ( .A(n8890), .B(n7778), .ZN(n7702) );
  XNOR2_X1 U9409 ( .A(n7702), .B(n8371), .ZN(n7788) );
  XNOR2_X1 U9410 ( .A(n8884), .B(n7778), .ZN(n7703) );
  XNOR2_X1 U9411 ( .A(n7703), .B(n8385), .ZN(n7861) );
  NAND2_X1 U9412 ( .A1(n7862), .A2(n7861), .ZN(n7860) );
  XNOR2_X1 U9413 ( .A(n7706), .B(n7705), .ZN(n7707) );
  NAND2_X1 U9414 ( .A1(n7747), .A2(n8349), .ZN(n7711) );
  INV_X1 U9415 ( .A(n7707), .ZN(n7708) );
  OR2_X1 U9416 ( .A1(n7709), .A2(n7708), .ZN(n7710) );
  NAND2_X1 U9417 ( .A1(n7711), .A2(n7710), .ZN(n7834) );
  XNOR2_X1 U9418 ( .A(n7839), .B(n7778), .ZN(n7712) );
  XNOR2_X1 U9419 ( .A(n7712), .B(n8360), .ZN(n7835) );
  NAND2_X1 U9420 ( .A1(n7834), .A2(n7835), .ZN(n7714) );
  NAND2_X1 U9421 ( .A1(n7712), .A2(n7750), .ZN(n7713) );
  XOR2_X1 U9422 ( .A(n7778), .B(n8867), .Z(n7716) );
  INV_X1 U9423 ( .A(n7716), .ZN(n7715) );
  XNOR2_X1 U9424 ( .A(n7715), .B(n8328), .ZN(n7808) );
  NOR2_X1 U9425 ( .A1(n7716), .A2(n8328), .ZN(n7717) );
  XNOR2_X1 U9426 ( .A(n8861), .B(n7778), .ZN(n7720) );
  XNOR2_X1 U9427 ( .A(n7719), .B(n7720), .ZN(n7878) );
  INV_X1 U9428 ( .A(n7719), .ZN(n7721) );
  NAND2_X1 U9429 ( .A1(n7721), .A2(n7720), .ZN(n7722) );
  XNOR2_X1 U9430 ( .A(n7732), .B(n7778), .ZN(n7723) );
  NAND2_X1 U9431 ( .A1(n7723), .A2(n8329), .ZN(n7776) );
  OAI21_X1 U9432 ( .B1(n7723), .B2(n8329), .A(n7776), .ZN(n7724) );
  NAND2_X1 U9433 ( .A1(n7726), .A2(n7777), .ZN(n7731) );
  INV_X1 U9434 ( .A(n8323), .ZN(n7728) );
  AOI22_X1 U9435 ( .A1(n8338), .A2(n7891), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7727) );
  OAI21_X1 U9436 ( .B1(n7728), .B2(n7821), .A(n7727), .ZN(n7729) );
  AOI21_X1 U9437 ( .B1(n7850), .B2(n8320), .A(n7729), .ZN(n7730) );
  OAI211_X1 U9438 ( .C1(n7732), .C2(n7898), .A(n7731), .B(n7730), .ZN(P2_U3154) );
  MUX2_X1 U9439 ( .A(n7801), .B(n4574), .S(n7733), .Z(n7797) );
  XNOR2_X1 U9440 ( .A(n7735), .B(n8124), .ZN(n7796) );
  NAND2_X1 U9441 ( .A1(n7797), .A2(n7796), .ZN(n7795) );
  NAND2_X1 U9442 ( .A1(n7795), .A2(n7736), .ZN(n7855) );
  XNOR2_X1 U9443 ( .A(n7737), .B(n8465), .ZN(n7856) );
  NOR2_X1 U9444 ( .A1(n7855), .A2(n7856), .ZN(n7854) );
  AOI21_X1 U9445 ( .B1(n7737), .B2(n8465), .A(n7854), .ZN(n7740) );
  OAI21_X1 U9446 ( .B1(n7740), .B2(n7739), .A(n7738), .ZN(n7741) );
  NAND2_X1 U9447 ( .A1(n7741), .A2(n7871), .ZN(n7746) );
  NAND2_X1 U9448 ( .A1(n7891), .A2(n8465), .ZN(n7742) );
  NAND2_X1 U9449 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8170) );
  OAI211_X1 U9450 ( .C1(n7743), .C2(n7893), .A(n7742), .B(n8170), .ZN(n7744)
         );
  AOI21_X1 U9451 ( .B1(n8471), .B2(n7895), .A(n7744), .ZN(n7745) );
  OAI211_X1 U9452 ( .C1(n8459), .C2(n7898), .A(n7746), .B(n7745), .ZN(P2_U3155) );
  XNOR2_X1 U9453 ( .A(n7747), .B(n8372), .ZN(n7753) );
  AOI22_X1 U9454 ( .A1(n8385), .A2(n7891), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7749) );
  NAND2_X1 U9455 ( .A1(n7895), .A2(n8363), .ZN(n7748) );
  OAI211_X1 U9456 ( .C1(n7750), .C2(n7893), .A(n7749), .B(n7748), .ZN(n7751)
         );
  AOI21_X1 U9457 ( .B1(n8878), .B2(n7883), .A(n7751), .ZN(n7752) );
  OAI21_X1 U9458 ( .B1(n7753), .B2(n7887), .A(n7752), .ZN(P2_U3156) );
  INV_X1 U9459 ( .A(n7754), .ZN(n7758) );
  AOI21_X1 U9460 ( .B1(n7850), .B2(n8125), .A(n7755), .ZN(n7757) );
  NAND2_X1 U9461 ( .A1(n7891), .A2(n8127), .ZN(n7756) );
  OAI211_X1 U9462 ( .C1(n7821), .C2(n7758), .A(n7757), .B(n7756), .ZN(n7764)
         );
  NAND2_X1 U9463 ( .A1(n4526), .A2(n7759), .ZN(n7761) );
  XNOR2_X1 U9464 ( .A(n7761), .B(n7760), .ZN(n7762) );
  NOR2_X1 U9465 ( .A1(n7762), .A2(n7887), .ZN(n7763) );
  AOI211_X1 U9466 ( .C1(n7765), .C2(n7883), .A(n7764), .B(n7763), .ZN(n7766)
         );
  INV_X1 U9467 ( .A(n7766), .ZN(P2_U3157) );
  XNOR2_X1 U9468 ( .A(n7767), .B(n8415), .ZN(n7768) );
  XNOR2_X1 U9469 ( .A(n7769), .B(n7768), .ZN(n7775) );
  INV_X1 U9470 ( .A(n7770), .ZN(n8407) );
  NAND2_X1 U9471 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8298) );
  OAI21_X1 U9472 ( .B1(n7893), .B2(n7791), .A(n8298), .ZN(n7771) );
  AOI21_X1 U9473 ( .B1(n7891), .B2(n8405), .A(n7771), .ZN(n7772) );
  OAI21_X1 U9474 ( .B1(n8407), .B2(n7821), .A(n7772), .ZN(n7773) );
  AOI21_X1 U9475 ( .B1(n8819), .B2(n7883), .A(n7773), .ZN(n7774) );
  OAI21_X1 U9476 ( .B1(n7775), .B2(n7887), .A(n7774), .ZN(P2_U3159) );
  XNOR2_X1 U9477 ( .A(n7919), .B(n7778), .ZN(n7779) );
  INV_X1 U9478 ( .A(n7780), .ZN(n7782) );
  INV_X1 U9479 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7781) );
  OAI22_X1 U9480 ( .A1(n7782), .A2(n7821), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7781), .ZN(n7784) );
  OAI22_X1 U9481 ( .A1(n7953), .A2(n7893), .B1(n7881), .B2(n7853), .ZN(n7783)
         );
  AOI211_X1 U9482 ( .C1(n7785), .C2(n7883), .A(n7784), .B(n7783), .ZN(n7786)
         );
  XOR2_X1 U9483 ( .A(n7788), .B(n7787), .Z(n7794) );
  NAND2_X1 U9484 ( .A1(n7895), .A2(n8388), .ZN(n7790) );
  AOI22_X1 U9485 ( .A1(n8385), .A2(n7850), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7789) );
  OAI211_X1 U9486 ( .C1(n7791), .C2(n7853), .A(n7790), .B(n7789), .ZN(n7792)
         );
  AOI21_X1 U9487 ( .B1(n8890), .B2(n7883), .A(n7792), .ZN(n7793) );
  OAI21_X1 U9488 ( .B1(n7794), .B2(n7887), .A(n7793), .ZN(P2_U3163) );
  OAI21_X1 U9489 ( .B1(n7797), .B2(n7796), .A(n7795), .ZN(n7798) );
  NAND2_X1 U9490 ( .A1(n7798), .A2(n7871), .ZN(n7805) );
  NOR2_X1 U9491 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7799), .ZN(n8146) );
  AOI21_X1 U9492 ( .B1(n7850), .B2(n8465), .A(n8146), .ZN(n7800) );
  OAI21_X1 U9493 ( .B1(n7801), .B2(n7853), .A(n7800), .ZN(n7802) );
  AOI21_X1 U9494 ( .B1(n7803), .B2(n7895), .A(n7802), .ZN(n7804) );
  OAI211_X1 U9495 ( .C1(n7806), .C2(n7898), .A(n7805), .B(n7804), .ZN(P2_U3164) );
  XOR2_X1 U9496 ( .A(n7807), .B(n7808), .Z(n7814) );
  INV_X1 U9497 ( .A(n7809), .ZN(n8340) );
  NAND2_X1 U9498 ( .A1(n8338), .A2(n7850), .ZN(n7811) );
  AOI22_X1 U9499 ( .A1(n8360), .A2(n7891), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7810) );
  OAI211_X1 U9500 ( .C1(n8340), .C2(n7821), .A(n7811), .B(n7810), .ZN(n7812)
         );
  AOI21_X1 U9501 ( .B1(n8867), .B2(n7883), .A(n7812), .ZN(n7813) );
  OAI21_X1 U9502 ( .B1(n7814), .B2(n7887), .A(n7813), .ZN(P2_U3165) );
  XNOR2_X1 U9503 ( .A(n7815), .B(n8423), .ZN(n7816) );
  XNOR2_X1 U9504 ( .A(n7817), .B(n7816), .ZN(n7824) );
  INV_X1 U9505 ( .A(n7818), .ZN(n8443) );
  NAND2_X1 U9506 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8214) );
  OAI21_X1 U9507 ( .B1(n7893), .B2(n7826), .A(n8214), .ZN(n7819) );
  AOI21_X1 U9508 ( .B1(n7891), .B2(n8464), .A(n7819), .ZN(n7820) );
  OAI21_X1 U9509 ( .B1(n8443), .B2(n7821), .A(n7820), .ZN(n7822) );
  AOI21_X1 U9510 ( .B1(n8830), .B2(n7883), .A(n7822), .ZN(n7823) );
  OAI21_X1 U9511 ( .B1(n7824), .B2(n7887), .A(n7823), .ZN(P2_U3166) );
  XNOR2_X1 U9512 ( .A(n7827), .B(n7826), .ZN(n7828) );
  XNOR2_X1 U9513 ( .A(n7825), .B(n7828), .ZN(n7833) );
  NAND2_X1 U9514 ( .A1(n7850), .A2(n8405), .ZN(n7829) );
  NAND2_X1 U9515 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8243) );
  OAI211_X1 U9516 ( .C1(n8423), .C2(n7853), .A(n7829), .B(n8243), .ZN(n7831)
         );
  INV_X1 U9517 ( .A(n8826), .ZN(n8432) );
  NOR2_X1 U9518 ( .A1(n8432), .A2(n7898), .ZN(n7830) );
  AOI211_X1 U9519 ( .C1(n8429), .C2(n7895), .A(n7831), .B(n7830), .ZN(n7832)
         );
  OAI21_X1 U9520 ( .B1(n7833), .B2(n7887), .A(n7832), .ZN(P2_U3168) );
  XOR2_X1 U9521 ( .A(n7835), .B(n7834), .Z(n7841) );
  AOI22_X1 U9522 ( .A1(n8372), .A2(n7891), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7837) );
  NAND2_X1 U9523 ( .A1(n7895), .A2(n8351), .ZN(n7836) );
  OAI211_X1 U9524 ( .C1(n8348), .C2(n7893), .A(n7837), .B(n7836), .ZN(n7838)
         );
  AOI21_X1 U9525 ( .B1(n7839), .B2(n7883), .A(n7838), .ZN(n7840) );
  OAI21_X1 U9526 ( .B1(n7841), .B2(n7887), .A(n7840), .ZN(P2_U3169) );
  XOR2_X1 U9527 ( .A(n7843), .B(n7842), .Z(n7848) );
  AOI22_X1 U9528 ( .A1(n8371), .A2(n7850), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7845) );
  NAND2_X1 U9529 ( .A1(n7895), .A2(n8395), .ZN(n7844) );
  OAI211_X1 U9530 ( .C1(n8394), .C2(n7853), .A(n7845), .B(n7844), .ZN(n7846)
         );
  AOI21_X1 U9531 ( .B1(n8896), .B2(n7883), .A(n7846), .ZN(n7847) );
  OAI21_X1 U9532 ( .B1(n7848), .B2(n7887), .A(n7847), .ZN(P2_U3173) );
  NAND2_X1 U9533 ( .A1(n7895), .A2(n8483), .ZN(n7852) );
  AOI21_X1 U9534 ( .B1(n7850), .B2(n8451), .A(n7849), .ZN(n7851) );
  OAI211_X1 U9535 ( .C1(n8479), .C2(n7853), .A(n7852), .B(n7851), .ZN(n7858)
         );
  AOI211_X1 U9536 ( .C1(n7856), .C2(n7855), .A(n7887), .B(n7854), .ZN(n7857)
         );
  AOI211_X1 U9537 ( .C1(n8929), .C2(n7883), .A(n7858), .B(n7857), .ZN(n7859)
         );
  INV_X1 U9538 ( .A(n7859), .ZN(P2_U3174) );
  INV_X1 U9539 ( .A(n8884), .ZN(n7867) );
  OAI211_X1 U9540 ( .C1(n7862), .C2(n7861), .A(n7860), .B(n7871), .ZN(n7866)
         );
  AOI22_X1 U9541 ( .A1(n8371), .A2(n7891), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7863) );
  OAI21_X1 U9542 ( .B1(n8349), .B2(n7893), .A(n7863), .ZN(n7864) );
  AOI21_X1 U9543 ( .B1(n8374), .B2(n7895), .A(n7864), .ZN(n7865) );
  OAI211_X1 U9544 ( .C1(n7867), .C2(n7898), .A(n7866), .B(n7865), .ZN(P2_U3175) );
  OAI21_X1 U9545 ( .B1(n7870), .B2(n7869), .A(n7868), .ZN(n7872) );
  NAND2_X1 U9546 ( .A1(n7872), .A2(n7871), .ZN(n7876) );
  NAND2_X1 U9547 ( .A1(n7891), .A2(n8440), .ZN(n7873) );
  NAND2_X1 U9548 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8270) );
  OAI211_X1 U9549 ( .C1(n8394), .C2(n7893), .A(n7873), .B(n8270), .ZN(n7874)
         );
  AOI21_X1 U9550 ( .B1(n8418), .B2(n7895), .A(n7874), .ZN(n7875) );
  OAI211_X1 U9551 ( .C1(n7877), .C2(n7898), .A(n7876), .B(n7875), .ZN(P2_U3178) );
  XNOR2_X1 U9552 ( .A(n7878), .B(n8338), .ZN(n7885) );
  AOI22_X1 U9553 ( .A1(n8328), .A2(n7891), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7880) );
  NAND2_X1 U9554 ( .A1(n8332), .A2(n7895), .ZN(n7879) );
  OAI211_X1 U9555 ( .C1(n7881), .C2(n7893), .A(n7880), .B(n7879), .ZN(n7882)
         );
  AOI21_X1 U9556 ( .B1(n8861), .B2(n7883), .A(n7882), .ZN(n7884) );
  OAI21_X1 U9557 ( .B1(n7885), .B2(n7887), .A(n7884), .ZN(P2_U3180) );
  INV_X1 U9558 ( .A(n8916), .ZN(n7899) );
  AOI211_X1 U9559 ( .C1(n7889), .C2(n7888), .A(n7887), .B(n7886), .ZN(n7890)
         );
  INV_X1 U9560 ( .A(n7890), .ZN(n7897) );
  NAND2_X1 U9561 ( .A1(n7891), .A2(n8451), .ZN(n7892) );
  NAND2_X1 U9562 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8196) );
  OAI211_X1 U9563 ( .C1(n8423), .C2(n7893), .A(n7892), .B(n8196), .ZN(n7894)
         );
  AOI21_X1 U9564 ( .B1(n8455), .B2(n7895), .A(n7894), .ZN(n7896) );
  OAI211_X1 U9565 ( .C1(n7899), .C2(n7898), .A(n7897), .B(n7896), .ZN(P2_U3181) );
  NAND2_X1 U9566 ( .A1(n7901), .A2(n7900), .ZN(n7903) );
  OR2_X1 U9567 ( .A1(n5746), .A2(n8766), .ZN(n7902) );
  INV_X1 U9568 ( .A(n8123), .ZN(n7907) );
  NAND2_X1 U9569 ( .A1(n8790), .A2(n7907), .ZN(n8099) );
  NAND2_X1 U9570 ( .A1(n8099), .A2(n7908), .ZN(n8094) );
  INV_X1 U9571 ( .A(n8102), .ZN(n7909) );
  NAND2_X1 U9572 ( .A1(n4442), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U9573 ( .A1(n7912), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U9574 ( .A1(n7913), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7914) );
  AND3_X1 U9575 ( .A1(n7916), .A2(n7915), .A3(n7914), .ZN(n7917) );
  NAND2_X1 U9576 ( .A1(n7918), .A2(n7917), .ZN(n8312) );
  AND2_X1 U9577 ( .A1(n8852), .A2(n8123), .ZN(n7947) );
  INV_X1 U9578 ( .A(n8849), .ZN(n8786) );
  NAND2_X1 U9579 ( .A1(n8088), .A2(n8089), .ZN(n8319) );
  INV_X1 U9580 ( .A(n8085), .ZN(n7920) );
  INV_X1 U9581 ( .A(n7921), .ZN(n7923) );
  NAND2_X1 U9582 ( .A1(n8074), .A2(n8071), .ZN(n8354) );
  INV_X1 U9583 ( .A(n8352), .ZN(n7924) );
  NOR2_X1 U9584 ( .A1(n8070), .A2(n7924), .ZN(n8358) );
  INV_X1 U9585 ( .A(n8413), .ZN(n7941) );
  NOR4_X1 U9586 ( .A1(n7927), .A2(n5686), .A3(n7926), .A4(n7925), .ZN(n7931)
         );
  NAND4_X1 U9587 ( .A1(n7931), .A2(n7930), .A3(n7929), .A4(n7928), .ZN(n7934)
         );
  NOR4_X1 U9588 ( .A1(n7934), .A2(n7989), .A3(n7933), .A4(n7932), .ZN(n7937)
         );
  NAND4_X1 U9589 ( .A1(n7937), .A2(n7936), .A3(n8029), .A4(n7935), .ZN(n7939)
         );
  INV_X1 U9590 ( .A(n7938), .ZN(n8031) );
  NAND2_X1 U9591 ( .A1(n8037), .A2(n8034), .ZN(n8473) );
  NOR4_X1 U9592 ( .A1(n8436), .A2(n7939), .A3(n8484), .A4(n8473), .ZN(n7940)
         );
  XNOR2_X1 U9593 ( .A(n8916), .B(n8464), .ZN(n8449) );
  NAND4_X1 U9594 ( .A1(n7941), .A2(n8428), .A3(n7940), .A4(n8449), .ZN(n7942)
         );
  NOR4_X1 U9595 ( .A1(n8381), .A2(n8391), .A3(n8402), .A4(n7942), .ZN(n7943)
         );
  NAND3_X1 U9596 ( .A1(n8358), .A2(n7943), .A3(n8366), .ZN(n7944) );
  NOR4_X1 U9597 ( .A1(n7946), .A2(n5617), .A3(n8319), .A4(n7945), .ZN(n7948)
         );
  INV_X1 U9598 ( .A(n7947), .ZN(n8104) );
  INV_X1 U9599 ( .A(n8312), .ZN(n7949) );
  NAND2_X1 U9600 ( .A1(n7951), .A2(n8103), .ZN(n7952) );
  NAND2_X1 U9601 ( .A1(n8102), .A2(n7952), .ZN(n7955) );
  OR2_X1 U9602 ( .A1(n7953), .A2(n8096), .ZN(n7954) );
  NAND2_X1 U9603 ( .A1(n7955), .A2(n7954), .ZN(n8092) );
  INV_X1 U9604 ( .A(n8092), .ZN(n8093) );
  MUX2_X1 U9605 ( .A(n8095), .B(n8106), .S(n8096), .Z(n8097) );
  AND2_X1 U9606 ( .A1(n7958), .A2(n7956), .ZN(n7996) );
  NAND2_X1 U9607 ( .A1(n8008), .A2(n7957), .ZN(n7960) );
  NAND2_X1 U9608 ( .A1(n7958), .A2(n7992), .ZN(n7959) );
  MUX2_X1 U9609 ( .A(n7960), .B(n7959), .S(n8096), .Z(n8012) );
  INV_X1 U9610 ( .A(n7984), .ZN(n7988) );
  NAND2_X1 U9611 ( .A1(n7968), .A2(n7961), .ZN(n7962) );
  NAND2_X1 U9612 ( .A1(n5884), .A2(n7962), .ZN(n7963) );
  NAND2_X1 U9613 ( .A1(n7963), .A2(n8096), .ZN(n7967) );
  INV_X1 U9614 ( .A(n7964), .ZN(n7965) );
  OAI21_X1 U9615 ( .B1(n7967), .B2(n7965), .A(n5687), .ZN(n7966) );
  MUX2_X1 U9616 ( .A(n5687), .B(n7966), .S(n8096), .Z(n7972) );
  INV_X1 U9617 ( .A(n5686), .ZN(n7969) );
  NAND3_X1 U9618 ( .A1(n7969), .A2(n7968), .A3(n7967), .ZN(n7970) );
  NAND3_X1 U9619 ( .A1(n7972), .A2(n7971), .A3(n7970), .ZN(n7979) );
  OAI21_X1 U9620 ( .B1(n8134), .B2(n7973), .A(n7997), .ZN(n7976) );
  NAND2_X1 U9621 ( .A1(n7982), .A2(n7974), .ZN(n7975) );
  MUX2_X1 U9622 ( .A(n7976), .B(n7975), .S(n8096), .Z(n7977) );
  INV_X1 U9623 ( .A(n7977), .ZN(n7978) );
  NAND2_X1 U9624 ( .A1(n7979), .A2(n7978), .ZN(n7981) );
  NAND2_X1 U9625 ( .A1(n7981), .A2(n7980), .ZN(n8001) );
  INV_X1 U9626 ( .A(n7982), .ZN(n7986) );
  AND2_X1 U9627 ( .A1(n7984), .A2(n7983), .ZN(n8002) );
  OAI211_X1 U9628 ( .C1(n8001), .C2(n7986), .A(n8002), .B(n7985), .ZN(n7987)
         );
  OAI211_X1 U9629 ( .C1(n7988), .C2(n7999), .A(n7987), .B(n8004), .ZN(n7990)
         );
  NAND2_X1 U9630 ( .A1(n7990), .A2(n8005), .ZN(n7995) );
  NAND2_X1 U9631 ( .A1(n7991), .A2(n8103), .ZN(n8015) );
  NAND2_X1 U9632 ( .A1(n8020), .A2(n7992), .ZN(n7993) );
  NOR2_X1 U9633 ( .A1(n8015), .A2(n7993), .ZN(n7994) );
  OAI211_X1 U9634 ( .C1(n7996), .C2(n8012), .A(n7995), .B(n7994), .ZN(n8025)
         );
  INV_X1 U9635 ( .A(n7997), .ZN(n8000) );
  OAI211_X1 U9636 ( .C1(n8001), .C2(n8000), .A(n7999), .B(n7998), .ZN(n8003)
         );
  NAND2_X1 U9637 ( .A1(n8003), .A2(n8002), .ZN(n8006) );
  NAND3_X1 U9638 ( .A1(n8006), .A2(n8005), .A3(n8004), .ZN(n8011) );
  NAND2_X1 U9639 ( .A1(n8007), .A2(n8096), .ZN(n8021) );
  NAND2_X1 U9640 ( .A1(n8014), .A2(n8008), .ZN(n8009) );
  NOR2_X1 U9641 ( .A1(n8021), .A2(n8009), .ZN(n8010) );
  OAI211_X1 U9642 ( .C1(n8013), .C2(n8012), .A(n8011), .B(n8010), .ZN(n8024)
         );
  OR2_X1 U9643 ( .A1(n8015), .A2(n8014), .ZN(n8019) );
  AND2_X1 U9644 ( .A1(n8125), .A2(n8103), .ZN(n8017) );
  OAI21_X1 U9645 ( .B1(n8103), .B2(n8125), .A(n4556), .ZN(n8016) );
  OAI21_X1 U9646 ( .B1(n8017), .B2(n4556), .A(n8016), .ZN(n8018) );
  OAI211_X1 U9647 ( .C1(n8021), .C2(n8020), .A(n8019), .B(n8018), .ZN(n8022)
         );
  INV_X1 U9648 ( .A(n8022), .ZN(n8023) );
  MUX2_X1 U9649 ( .A(n8027), .B(n8026), .S(n8103), .Z(n8028) );
  MUX2_X1 U9650 ( .A(n8032), .B(n8031), .S(n8103), .Z(n8033) );
  NAND3_X1 U9651 ( .A1(n8038), .A2(n8449), .A3(n8034), .ZN(n8036) );
  NAND3_X1 U9652 ( .A1(n8036), .A2(n8044), .A3(n8035), .ZN(n8041) );
  NAND3_X1 U9653 ( .A1(n8050), .A2(n8051), .A3(n8046), .ZN(n8045) );
  NAND3_X1 U9654 ( .A1(n8045), .A2(n8055), .A3(n8047), .ZN(n8054) );
  NAND2_X1 U9655 ( .A1(n8046), .A2(n8411), .ZN(n8049) );
  OAI211_X1 U9656 ( .C1(n8050), .C2(n8049), .A(n8048), .B(n8047), .ZN(n8052)
         );
  NAND2_X1 U9657 ( .A1(n8052), .A2(n8051), .ZN(n8053) );
  INV_X1 U9658 ( .A(n8377), .ZN(n8059) );
  AND2_X1 U9659 ( .A1(n8061), .A2(n8055), .ZN(n8057) );
  MUX2_X1 U9660 ( .A(n8057), .B(n8056), .S(n8096), .Z(n8058) );
  MUX2_X1 U9661 ( .A(n8061), .B(n8060), .S(n8103), .Z(n8062) );
  NAND2_X1 U9662 ( .A1(n8884), .A2(n8063), .ZN(n8064) );
  AND2_X1 U9663 ( .A1(n8352), .A2(n8064), .ZN(n8068) );
  INV_X1 U9664 ( .A(n8065), .ZN(n8066) );
  NOR2_X1 U9665 ( .A1(n8070), .A2(n8066), .ZN(n8067) );
  MUX2_X1 U9666 ( .A(n8068), .B(n8067), .S(n8103), .Z(n8069) );
  AND2_X1 U9667 ( .A1(n4816), .A2(n8074), .ZN(n8073) );
  INV_X1 U9668 ( .A(n8071), .ZN(n8072) );
  AOI21_X1 U9669 ( .B1(n8076), .B2(n8073), .A(n8072), .ZN(n8078) );
  INV_X1 U9670 ( .A(n8074), .ZN(n8075) );
  AOI21_X1 U9671 ( .B1(n8076), .B2(n4508), .A(n8075), .ZN(n8077) );
  INV_X1 U9672 ( .A(n8079), .ZN(n8080) );
  MUX2_X1 U9673 ( .A(n8081), .B(n8080), .S(n8096), .Z(n8082) );
  INV_X1 U9674 ( .A(n8083), .ZN(n8084) );
  MUX2_X1 U9675 ( .A(n8085), .B(n8084), .S(n8103), .Z(n8086) );
  NOR2_X1 U9676 ( .A1(n8319), .A2(n8086), .ZN(n8087) );
  MUX2_X1 U9677 ( .A(n8089), .B(n8088), .S(n8096), .Z(n8090) );
  NAND3_X1 U9678 ( .A1(n8092), .A2(n8091), .A3(n8090), .ZN(n8098) );
  OAI21_X1 U9679 ( .B1(n8093), .B2(n8097), .A(n8098), .ZN(n8105) );
  AOI21_X1 U9680 ( .B1(n8105), .B2(n8095), .A(n8094), .ZN(n8111) );
  INV_X1 U9681 ( .A(n8108), .ZN(n8110) );
  NAND3_X1 U9682 ( .A1(n8101), .A2(n8100), .A3(n8099), .ZN(n8107) );
  XNOR2_X1 U9683 ( .A(n8115), .B(n8291), .ZN(n8122) );
  NOR3_X1 U9684 ( .A1(n8117), .A2(n8116), .A3(n5633), .ZN(n8120) );
  OAI21_X1 U9685 ( .B1(n8121), .B2(n8118), .A(P2_B_REG_SCAN_IN), .ZN(n8119) );
  OAI22_X1 U9686 ( .A1(n8122), .A2(n8121), .B1(n8120), .B2(n8119), .ZN(
        P2_U3296) );
  MUX2_X1 U9687 ( .A(n8312), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8267), .Z(
        P2_U3522) );
  MUX2_X1 U9688 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8123), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9689 ( .A(n8320), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8267), .Z(
        P2_U3519) );
  MUX2_X1 U9690 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8329), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9691 ( .A(n8338), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8267), .Z(
        P2_U3517) );
  MUX2_X1 U9692 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8328), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9693 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8360), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9694 ( .A(n8372), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8267), .Z(
        P2_U3514) );
  MUX2_X1 U9695 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8385), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9696 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8371), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9697 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8404), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9698 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8415), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9699 ( .A(n8405), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8267), .Z(
        P2_U3509) );
  MUX2_X1 U9700 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8440), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9701 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8452), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9702 ( .A(n8464), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8267), .Z(
        P2_U3506) );
  MUX2_X1 U9703 ( .A(n8451), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8267), .Z(
        P2_U3505) );
  MUX2_X1 U9704 ( .A(n8465), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8267), .Z(
        P2_U3504) );
  MUX2_X1 U9705 ( .A(n8124), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8267), .Z(
        P2_U3503) );
  MUX2_X1 U9706 ( .A(n8125), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8267), .Z(
        P2_U3502) );
  MUX2_X1 U9707 ( .A(n8126), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8267), .Z(
        P2_U3501) );
  MUX2_X1 U9708 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8127), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9709 ( .A(n8128), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8267), .Z(
        P2_U3499) );
  MUX2_X1 U9710 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8129), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9711 ( .A(n8130), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8267), .Z(
        P2_U3497) );
  MUX2_X1 U9712 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8131), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9713 ( .A(n8132), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8267), .Z(
        P2_U3495) );
  MUX2_X1 U9714 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8133), .S(P2_U3893), .Z(
        P2_U3494) );
  INV_X1 U9715 ( .A(n8134), .ZN(n8135) );
  MUX2_X1 U9716 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8135), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9717 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n5248), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U9718 ( .A(n8136), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8267), .Z(
        P2_U3491) );
  AND3_X1 U9719 ( .A1(n8139), .A2(n8138), .A3(n8137), .ZN(n8141) );
  OAI21_X1 U9720 ( .B1(n8142), .B2(n8141), .A(n8140), .ZN(n8157) );
  OAI21_X1 U9721 ( .B1(n8145), .B2(n8144), .A(n8143), .ZN(n8147) );
  AOI21_X1 U9722 ( .B1(n8148), .B2(n8147), .A(n8146), .ZN(n8156) );
  AOI22_X1 U9723 ( .A1(n8195), .A2(P2_ADDR_REG_12__SCAN_IN), .B1(n8297), .B2(
        n8149), .ZN(n8155) );
  OAI21_X1 U9724 ( .B1(n8152), .B2(n8151), .A(n8150), .ZN(n8153) );
  NAND2_X1 U9725 ( .A1(n8153), .A2(n8309), .ZN(n8154) );
  NAND4_X1 U9726 ( .A1(n8157), .A2(n8156), .A3(n8155), .A4(n8154), .ZN(
        P2_U3194) );
  NOR2_X1 U9727 ( .A1(n8174), .A2(n8158), .ZN(n8160) );
  NOR2_X1 U9728 ( .A1(n8160), .A2(n8159), .ZN(n8163) );
  INV_X1 U9729 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8161) );
  AOI22_X1 U9730 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8177), .B1(n8193), .B2(
        n8161), .ZN(n8162) );
  NOR2_X1 U9731 ( .A1(n8163), .A2(n8162), .ZN(n8185) );
  AOI21_X1 U9732 ( .B1(n8163), .B2(n8162), .A(n8185), .ZN(n8184) );
  MUX2_X1 U9733 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8292), .Z(n8187) );
  XNOR2_X1 U9734 ( .A(n8187), .B(n8177), .ZN(n8169) );
  OR2_X1 U9735 ( .A1(n8165), .A2(n8164), .ZN(n8167) );
  NAND2_X1 U9736 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  NAND2_X1 U9737 ( .A1(n8169), .A2(n8168), .ZN(n8188) );
  OAI21_X1 U9738 ( .B1(n8169), .B2(n8168), .A(n8188), .ZN(n8182) );
  INV_X1 U9739 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U9740 ( .A1(n8297), .A2(n8177), .ZN(n8171) );
  OAI211_X1 U9741 ( .C1(n8300), .C2(n8172), .A(n8171), .B(n8170), .ZN(n8181)
         );
  NOR2_X1 U9742 ( .A1(n8174), .A2(n8173), .ZN(n8176) );
  INV_X1 U9743 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8838) );
  XNOR2_X1 U9744 ( .A(n8177), .B(n8838), .ZN(n8178) );
  AOI21_X1 U9745 ( .B1(n4521), .B2(n8178), .A(n8192), .ZN(n8179) );
  NOR2_X1 U9746 ( .A1(n8179), .A2(n8310), .ZN(n8180) );
  AOI211_X1 U9747 ( .C1(n8309), .C2(n8182), .A(n8181), .B(n8180), .ZN(n8183)
         );
  OAI21_X1 U9748 ( .B1(n8184), .B2(n8306), .A(n8183), .ZN(P2_U3196) );
  INV_X1 U9749 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8454) );
  AOI21_X1 U9750 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8193), .A(n8185), .ZN(
        n8217) );
  XNOR2_X1 U9751 ( .A(n8217), .B(n8218), .ZN(n8186) );
  AOI21_X1 U9752 ( .B1(n8454), .B2(n8186), .A(n8219), .ZN(n8202) );
  INV_X1 U9753 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8834) );
  MUX2_X1 U9754 ( .A(n8454), .B(n8834), .S(n8292), .Z(n8209) );
  XOR2_X1 U9755 ( .A(n8218), .B(n8209), .Z(n8191) );
  OR2_X1 U9756 ( .A1(n8187), .A2(n8193), .ZN(n8189) );
  NAND2_X1 U9757 ( .A1(n8189), .A2(n8188), .ZN(n8190) );
  NAND2_X1 U9758 ( .A1(n8191), .A2(n8190), .ZN(n8210) );
  OAI21_X1 U9759 ( .B1(n8191), .B2(n8190), .A(n8210), .ZN(n8200) );
  AOI21_X1 U9760 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8193), .A(n8192), .ZN(
        n8203) );
  AOI21_X1 U9761 ( .B1(n8194), .B2(n8834), .A(n8204), .ZN(n8198) );
  AOI22_X1 U9762 ( .A1(n8195), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(n8297), .B2(
        n8218), .ZN(n8197) );
  OAI211_X1 U9763 ( .C1(n8198), .C2(n8310), .A(n8197), .B(n8196), .ZN(n8199)
         );
  AOI21_X1 U9764 ( .B1(n8309), .B2(n8200), .A(n8199), .ZN(n8201) );
  OAI21_X1 U9765 ( .B1(n8202), .B2(n8306), .A(n8201), .ZN(P2_U3197) );
  NAND2_X1 U9766 ( .A1(n8237), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8232) );
  INV_X1 U9767 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U9768 ( .A1(n8222), .A2(n8575), .ZN(n8205) );
  NAND2_X1 U9769 ( .A1(n8232), .A2(n8205), .ZN(n8207) );
  INV_X1 U9770 ( .A(n8233), .ZN(n8206) );
  AOI21_X1 U9771 ( .B1(n8208), .B2(n8207), .A(n8206), .ZN(n8231) );
  MUX2_X1 U9772 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8292), .Z(n8238) );
  XNOR2_X1 U9773 ( .A(n8238), .B(n8222), .ZN(n8213) );
  NAND2_X1 U9774 ( .A1(n8209), .A2(n8218), .ZN(n8211) );
  NAND2_X1 U9775 ( .A1(n8211), .A2(n8210), .ZN(n8212) );
  NAND2_X1 U9776 ( .A1(n8213), .A2(n8212), .ZN(n8239) );
  OAI21_X1 U9777 ( .B1(n8213), .B2(n8212), .A(n8239), .ZN(n8229) );
  INV_X1 U9778 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U9779 ( .A1(n8297), .A2(n8222), .ZN(n8215) );
  OAI211_X1 U9780 ( .C1(n8300), .C2(n8216), .A(n8215), .B(n8214), .ZN(n8228)
         );
  NOR2_X1 U9781 ( .A1(n8218), .A2(n8217), .ZN(n8220) );
  NAND2_X1 U9782 ( .A1(n8237), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8246) );
  INV_X1 U9783 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8221) );
  NAND2_X1 U9784 ( .A1(n8222), .A2(n8221), .ZN(n8223) );
  NAND2_X1 U9785 ( .A1(n8246), .A2(n8223), .ZN(n8224) );
  NAND2_X1 U9786 ( .A1(n8225), .A2(n8224), .ZN(n8226) );
  AOI21_X1 U9787 ( .B1(n8247), .B2(n8226), .A(n8306), .ZN(n8227) );
  AOI211_X1 U9788 ( .C1(n8309), .C2(n8229), .A(n8228), .B(n8227), .ZN(n8230)
         );
  OAI21_X1 U9789 ( .B1(n8231), .B2(n8310), .A(n8230), .ZN(P2_U3198) );
  XNOR2_X1 U9790 ( .A(n8256), .B(n8273), .ZN(n8234) );
  INV_X1 U9791 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8235) );
  NOR2_X1 U9792 ( .A1(n8235), .A2(n8234), .ZN(n8257) );
  AOI21_X1 U9793 ( .B1(n8234), .B2(n8235), .A(n8257), .ZN(n8255) );
  MUX2_X1 U9794 ( .A(n8249), .B(n8235), .S(n8292), .Z(n8261) );
  XNOR2_X1 U9795 ( .A(n8261), .B(n8236), .ZN(n8242) );
  OR2_X1 U9796 ( .A1(n8238), .A2(n8237), .ZN(n8240) );
  NAND2_X1 U9797 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  NAND2_X1 U9798 ( .A1(n8242), .A2(n8241), .ZN(n8262) );
  OAI21_X1 U9799 ( .B1(n8242), .B2(n8241), .A(n8262), .ZN(n8253) );
  INV_X1 U9800 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U9801 ( .A1(n8297), .A2(n8273), .ZN(n8244) );
  OAI211_X1 U9802 ( .C1(n8300), .C2(n8245), .A(n8244), .B(n8243), .ZN(n8252)
         );
  AOI21_X1 U9803 ( .B1(n8249), .B2(n8248), .A(n8274), .ZN(n8250) );
  NOR2_X1 U9804 ( .A1(n8250), .A2(n8306), .ZN(n8251) );
  AOI211_X1 U9805 ( .C1(n8309), .C2(n8253), .A(n8252), .B(n8251), .ZN(n8254)
         );
  OAI21_X1 U9806 ( .B1(n8255), .B2(n8310), .A(n8254), .ZN(P2_U3199) );
  NOR2_X1 U9807 ( .A1(n8273), .A2(n8256), .ZN(n8258) );
  NAND2_X1 U9808 ( .A1(n8276), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8283) );
  OAI21_X1 U9809 ( .B1(n8276), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8283), .ZN(
        n8259) );
  NOR2_X1 U9810 ( .A1(n8260), .A2(n8259), .ZN(n8285) );
  AOI21_X1 U9811 ( .B1(n8260), .B2(n8259), .A(n8285), .ZN(n8281) );
  NAND2_X1 U9812 ( .A1(n8261), .A2(n8273), .ZN(n8263) );
  NAND2_X1 U9813 ( .A1(n8263), .A2(n8262), .ZN(n8265) );
  INV_X1 U9814 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8417) );
  INV_X1 U9815 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8823) );
  MUX2_X1 U9816 ( .A(n8417), .B(n8823), .S(n8292), .Z(n8264) );
  NAND2_X1 U9817 ( .A1(n8265), .A2(n8264), .ZN(n8289) );
  NAND2_X1 U9818 ( .A1(n8288), .A2(n8289), .ZN(n8268) );
  OAI21_X1 U9819 ( .B1(n8267), .B2(n8268), .A(n8266), .ZN(n8280) );
  INV_X1 U9820 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8271) );
  NAND3_X1 U9821 ( .A1(n8309), .A2(n8276), .A3(n8268), .ZN(n8269) );
  OAI211_X1 U9822 ( .C1(n8300), .C2(n8271), .A(n8270), .B(n8269), .ZN(n8279)
         );
  NOR2_X1 U9823 ( .A1(n8273), .A2(n8272), .ZN(n8275) );
  NAND2_X1 U9824 ( .A1(n8276), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8301) );
  OAI21_X1 U9825 ( .B1(n8276), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8301), .ZN(
        n8277) );
  NOR2_X1 U9826 ( .A1(n8278), .A2(n8277), .ZN(n8303) );
  INV_X1 U9827 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8282) );
  XNOR2_X1 U9828 ( .A(n8291), .B(n8282), .ZN(n8293) );
  INV_X1 U9829 ( .A(n8293), .ZN(n8286) );
  INV_X1 U9830 ( .A(n8283), .ZN(n8284) );
  NAND2_X1 U9831 ( .A1(n8288), .A2(n8287), .ZN(n8290) );
  NAND2_X1 U9832 ( .A1(n8290), .A2(n8289), .ZN(n8295) );
  INV_X1 U9833 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8696) );
  MUX2_X1 U9834 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8696), .S(n8291), .Z(n8304)
         );
  MUX2_X1 U9835 ( .A(n8304), .B(n8293), .S(n8292), .Z(n8294) );
  XNOR2_X1 U9836 ( .A(n8295), .B(n8294), .ZN(n8308) );
  INV_X1 U9837 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U9838 ( .A1(n8297), .A2(n8296), .ZN(n8299) );
  OAI211_X1 U9839 ( .C1(n8678), .C2(n8300), .A(n8299), .B(n8298), .ZN(n8307)
         );
  INV_X1 U9840 ( .A(n8301), .ZN(n8302) );
  NOR2_X1 U9841 ( .A1(n8303), .A2(n8302), .ZN(n8305) );
  NAND2_X1 U9842 ( .A1(n8312), .A2(n8311), .ZN(n8847) );
  AOI21_X1 U9843 ( .B1(n8313), .B2(n8847), .A(n8489), .ZN(n8315) );
  AOI21_X1 U9844 ( .B1(n8489), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8315), .ZN(
        n8314) );
  OAI21_X1 U9845 ( .B1(n8849), .B2(n8431), .A(n8314), .ZN(P2_U3202) );
  AOI21_X1 U9846 ( .B1(n8489), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8315), .ZN(
        n8316) );
  OAI21_X1 U9847 ( .B1(n8852), .B2(n8431), .A(n8316), .ZN(P2_U3203) );
  XOR2_X1 U9848 ( .A(n8319), .B(n8317), .Z(n8858) );
  INV_X1 U9849 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8322) );
  XOR2_X1 U9850 ( .A(n8319), .B(n8318), .Z(n8321) );
  AOI222_X2 U9851 ( .A1(n8321), .A2(n8461), .B1(n8338), .B2(n8466), .C1(n8320), 
        .C2(n8463), .ZN(n8853) );
  MUX2_X1 U9852 ( .A(n8322), .B(n8853), .S(n10233), .Z(n8325) );
  AOI22_X1 U9853 ( .A1(n8855), .A2(n10226), .B1(n10228), .B2(n8323), .ZN(n8324) );
  OAI211_X1 U9854 ( .C1(n8858), .C2(n8783), .A(n8325), .B(n8324), .ZN(P2_U3206) );
  XNOR2_X1 U9855 ( .A(n8326), .B(n4463), .ZN(n8864) );
  INV_X1 U9856 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8331) );
  XNOR2_X1 U9857 ( .A(n8327), .B(n4463), .ZN(n8330) );
  AOI222_X1 U9858 ( .A1(n8461), .A2(n8330), .B1(n8329), .B2(n8463), .C1(n8328), 
        .C2(n8466), .ZN(n8859) );
  MUX2_X1 U9859 ( .A(n8331), .B(n8859), .S(n10233), .Z(n8334) );
  AOI22_X1 U9860 ( .A1(n8861), .A2(n10226), .B1(n10228), .B2(n8332), .ZN(n8333) );
  OAI211_X1 U9861 ( .C1(n8864), .C2(n8783), .A(n8334), .B(n8333), .ZN(P2_U3207) );
  XOR2_X1 U9862 ( .A(n8337), .B(n8335), .Z(n8870) );
  XOR2_X1 U9863 ( .A(n8336), .B(n8337), .Z(n8339) );
  AOI222_X1 U9864 ( .A1(n8461), .A2(n8339), .B1(n8338), .B2(n8463), .C1(n8360), 
        .C2(n8466), .ZN(n8865) );
  INV_X1 U9865 ( .A(n8865), .ZN(n8343) );
  INV_X1 U9866 ( .A(n8867), .ZN(n8341) );
  OAI22_X1 U9867 ( .A1(n8341), .A2(n8458), .B1(n8340), .B2(n8444), .ZN(n8342)
         );
  OAI21_X1 U9868 ( .B1(n8343), .B2(n8342), .A(n10233), .ZN(n8345) );
  NAND2_X1 U9869 ( .A1(n8489), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8344) );
  OAI211_X1 U9870 ( .C1(n8870), .C2(n8783), .A(n8345), .B(n8344), .ZN(P2_U3208) );
  NOR2_X1 U9871 ( .A1(n8872), .A2(n8458), .ZN(n8350) );
  XOR2_X1 U9872 ( .A(n8346), .B(n8354), .Z(n8347) );
  OAI222_X1 U9873 ( .A1(n8480), .A2(n8349), .B1(n8481), .B2(n8348), .C1(n8477), 
        .C2(n8347), .ZN(n8871) );
  AOI211_X1 U9874 ( .C1(n10228), .C2(n8351), .A(n8350), .B(n8871), .ZN(n8356)
         );
  NAND2_X1 U9875 ( .A1(n5054), .A2(n8352), .ZN(n8353) );
  XOR2_X1 U9876 ( .A(n8354), .B(n8353), .Z(n8803) );
  AOI22_X1 U9877 ( .A1(n8803), .A2(n8486), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8489), .ZN(n8355) );
  OAI21_X1 U9878 ( .B1(n8356), .B2(n8489), .A(n8355), .ZN(P2_U3209) );
  XNOR2_X1 U9879 ( .A(n8357), .B(n8358), .ZN(n8881) );
  INV_X1 U9880 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8362) );
  XOR2_X1 U9881 ( .A(n8359), .B(n8358), .Z(n8361) );
  AOI222_X1 U9882 ( .A1(n8461), .A2(n8361), .B1(n8385), .B2(n8466), .C1(n8360), 
        .C2(n8463), .ZN(n8876) );
  MUX2_X1 U9883 ( .A(n8362), .B(n8876), .S(n10233), .Z(n8365) );
  AOI22_X1 U9884 ( .A1(n8878), .A2(n10226), .B1(n10228), .B2(n8363), .ZN(n8364) );
  OAI211_X1 U9885 ( .C1(n8881), .C2(n8783), .A(n8365), .B(n8364), .ZN(P2_U3210) );
  XNOR2_X1 U9886 ( .A(n8367), .B(n8366), .ZN(n8887) );
  OAI21_X1 U9887 ( .B1(n8370), .B2(n8369), .A(n8368), .ZN(n8373) );
  AOI222_X1 U9888 ( .A1(n8461), .A2(n8373), .B1(n8372), .B2(n8463), .C1(n8371), 
        .C2(n8466), .ZN(n8882) );
  MUX2_X1 U9889 ( .A(n8591), .B(n8882), .S(n10233), .Z(n8376) );
  AOI22_X1 U9890 ( .A1(n8884), .A2(n10226), .B1(n10228), .B2(n8374), .ZN(n8375) );
  OAI211_X1 U9891 ( .C1(n8887), .C2(n8783), .A(n8376), .B(n8375), .ZN(P2_U3211) );
  NAND2_X1 U9892 ( .A1(n8378), .A2(n8377), .ZN(n8379) );
  XNOR2_X1 U9893 ( .A(n8379), .B(n8381), .ZN(n8893) );
  INV_X1 U9894 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8387) );
  OR3_X1 U9895 ( .A1(n8380), .A2(n8382), .A3(n8381), .ZN(n8383) );
  NAND2_X1 U9896 ( .A1(n8384), .A2(n8383), .ZN(n8386) );
  AOI222_X1 U9897 ( .A1(n8461), .A2(n8386), .B1(n8385), .B2(n8463), .C1(n8404), 
        .C2(n8466), .ZN(n8888) );
  MUX2_X1 U9898 ( .A(n8387), .B(n8888), .S(n10233), .Z(n8390) );
  AOI22_X1 U9899 ( .A1(n8890), .A2(n10226), .B1(n10228), .B2(n8388), .ZN(n8389) );
  OAI211_X1 U9900 ( .C1(n8893), .C2(n8783), .A(n8390), .B(n8389), .ZN(P2_U3212) );
  INV_X1 U9901 ( .A(n8391), .ZN(n8397) );
  AOI21_X1 U9902 ( .B1(n8397), .B2(n4520), .A(n8380), .ZN(n8392) );
  OAI222_X1 U9903 ( .A1(n8480), .A2(n8394), .B1(n8481), .B2(n8393), .C1(n8477), 
        .C2(n8392), .ZN(n8815) );
  AOI21_X1 U9904 ( .B1(n10228), .B2(n8395), .A(n8815), .ZN(n8400) );
  AOI22_X1 U9905 ( .A1(n8896), .A2(n10226), .B1(P2_REG2_REG_20__SCAN_IN), .B2(
        n8489), .ZN(n8399) );
  XNOR2_X1 U9906 ( .A(n8396), .B(n8397), .ZN(n8897) );
  NAND2_X1 U9907 ( .A1(n8897), .A2(n8486), .ZN(n8398) );
  OAI211_X1 U9908 ( .C1(n8400), .C2(n8489), .A(n8399), .B(n8398), .ZN(P2_U3213) );
  XNOR2_X1 U9909 ( .A(n8401), .B(n8402), .ZN(n8822) );
  XOR2_X1 U9910 ( .A(n8403), .B(n8402), .Z(n8406) );
  AOI222_X1 U9911 ( .A1(n8461), .A2(n8406), .B1(n8405), .B2(n8466), .C1(n8404), 
        .C2(n8463), .ZN(n8821) );
  OR2_X1 U9912 ( .A1(n8821), .A2(n8489), .ZN(n8410) );
  OAI22_X1 U9913 ( .A1(n10233), .A2(n8696), .B1(n8407), .B2(n8444), .ZN(n8408)
         );
  AOI21_X1 U9914 ( .B1(n8819), .B2(n10226), .A(n8408), .ZN(n8409) );
  OAI211_X1 U9915 ( .C1(n8822), .C2(n8783), .A(n8410), .B(n8409), .ZN(P2_U3214) );
  NAND2_X1 U9916 ( .A1(n8427), .A2(n8411), .ZN(n8412) );
  XNOR2_X1 U9917 ( .A(n8412), .B(n8413), .ZN(n8906) );
  XNOR2_X1 U9918 ( .A(n8414), .B(n8413), .ZN(n8416) );
  AOI222_X1 U9919 ( .A1(n8461), .A2(n8416), .B1(n8440), .B2(n8466), .C1(n8415), 
        .C2(n8463), .ZN(n8901) );
  MUX2_X1 U9920 ( .A(n8417), .B(n8901), .S(n10233), .Z(n8420) );
  AOI22_X1 U9921 ( .A1(n8903), .A2(n10226), .B1(n10228), .B2(n8418), .ZN(n8419) );
  OAI211_X1 U9922 ( .C1(n8906), .C2(n8783), .A(n8420), .B(n8419), .ZN(P2_U3215) );
  AOI211_X1 U9923 ( .C1(n8428), .C2(n8421), .A(n8477), .B(n8422), .ZN(n8426)
         );
  OAI22_X1 U9924 ( .A1(n8424), .A2(n8481), .B1(n8423), .B2(n8480), .ZN(n8425)
         );
  NOR2_X1 U9925 ( .A1(n8426), .A2(n8425), .ZN(n8829) );
  OAI21_X1 U9926 ( .B1(n4525), .B2(n8428), .A(n8427), .ZN(n8827) );
  AOI22_X1 U9927 ( .A1(n8489), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n10228), .B2(
        n8429), .ZN(n8430) );
  OAI21_X1 U9928 ( .B1(n8432), .B2(n8431), .A(n8430), .ZN(n8433) );
  AOI21_X1 U9929 ( .B1(n8827), .B2(n8486), .A(n8433), .ZN(n8434) );
  OAI21_X1 U9930 ( .B1(n8829), .B2(n8489), .A(n8434), .ZN(P2_U3216) );
  XNOR2_X1 U9931 ( .A(n8435), .B(n8436), .ZN(n8911) );
  OAI21_X1 U9932 ( .B1(n8437), .B2(n8436), .A(n8461), .ZN(n8438) );
  OR2_X1 U9933 ( .A1(n8439), .A2(n8438), .ZN(n8442) );
  AOI22_X1 U9934 ( .A1(n8440), .A2(n8463), .B1(n8466), .B2(n8464), .ZN(n8441)
         );
  NAND2_X1 U9935 ( .A1(n8442), .A2(n8441), .ZN(n8908) );
  NOR2_X1 U9936 ( .A1(n8444), .A2(n8443), .ZN(n8445) );
  OAI21_X1 U9937 ( .B1(n8908), .B2(n8445), .A(n10233), .ZN(n8447) );
  AOI22_X1 U9938 ( .A1(n8830), .A2(n10226), .B1(P2_REG2_REG_16__SCAN_IN), .B2(
        n8489), .ZN(n8446) );
  OAI211_X1 U9939 ( .C1(n8911), .C2(n8783), .A(n8447), .B(n8446), .ZN(P2_U3217) );
  XOR2_X1 U9940 ( .A(n8449), .B(n8448), .Z(n8920) );
  XOR2_X1 U9941 ( .A(n8450), .B(n8449), .Z(n8453) );
  AOI222_X1 U9942 ( .A1(n8461), .A2(n8453), .B1(n8452), .B2(n8463), .C1(n8451), 
        .C2(n8466), .ZN(n8914) );
  MUX2_X1 U9943 ( .A(n8454), .B(n8914), .S(n10233), .Z(n8457) );
  AOI22_X1 U9944 ( .A1(n8916), .A2(n10226), .B1(n10228), .B2(n8455), .ZN(n8456) );
  OAI211_X1 U9945 ( .C1(n8920), .C2(n8783), .A(n8457), .B(n8456), .ZN(P2_U3218) );
  NOR2_X1 U9946 ( .A1(n8459), .A2(n8458), .ZN(n8470) );
  XNOR2_X1 U9947 ( .A(n8460), .B(n8473), .ZN(n8462) );
  NAND2_X1 U9948 ( .A1(n8462), .A2(n8461), .ZN(n8468) );
  AOI22_X1 U9949 ( .A1(n8466), .A2(n8465), .B1(n8464), .B2(n8463), .ZN(n8467)
         );
  AND2_X1 U9950 ( .A1(n8468), .A2(n8467), .ZN(n8921) );
  INV_X1 U9951 ( .A(n8921), .ZN(n8469) );
  AOI211_X1 U9952 ( .C1(n10228), .C2(n8471), .A(n8470), .B(n8469), .ZN(n8475)
         );
  XOR2_X1 U9953 ( .A(n8473), .B(n8472), .Z(n8924) );
  AOI22_X1 U9954 ( .A1(n8924), .A2(n8486), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8489), .ZN(n8474) );
  OAI21_X1 U9955 ( .B1(n8475), .B2(n8489), .A(n8474), .ZN(P2_U3219) );
  XNOR2_X1 U9956 ( .A(n8476), .B(n8484), .ZN(n8478) );
  OAI222_X1 U9957 ( .A1(n8481), .A2(n4972), .B1(n8480), .B2(n8479), .C1(n8478), 
        .C2(n8477), .ZN(n8841) );
  AOI21_X1 U9958 ( .B1(n8482), .B2(n8929), .A(n8841), .ZN(n8490) );
  AOI22_X1 U9959 ( .A1(n8489), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10228), .B2(
        n8483), .ZN(n8488) );
  XNOR2_X1 U9960 ( .A(n8485), .B(n8484), .ZN(n8932) );
  NAND2_X1 U9961 ( .A1(n8932), .A2(n8486), .ZN(n8487) );
  OAI211_X1 U9962 ( .C1(n8490), .C2(n8489), .A(n8488), .B(n8487), .ZN(P2_U3220) );
  NOR2_X1 U9963 ( .A1(keyinput114), .A2(keyinput36), .ZN(n8491) );
  NAND3_X1 U9964 ( .A1(keyinput39), .A2(keyinput51), .A3(n8491), .ZN(n8492) );
  NOR4_X1 U9965 ( .A1(keyinput109), .A2(keyinput115), .A3(keyinput78), .A4(
        n8492), .ZN(n8503) );
  INV_X1 U9966 ( .A(keyinput106), .ZN(n8493) );
  NOR4_X1 U9967 ( .A1(keyinput77), .A2(keyinput81), .A3(keyinput94), .A4(n8493), .ZN(n8502) );
  NAND2_X1 U9968 ( .A1(keyinput57), .A2(keyinput61), .ZN(n8494) );
  NOR3_X1 U9969 ( .A1(keyinput4), .A2(keyinput24), .A3(n8494), .ZN(n8501) );
  NOR2_X1 U9970 ( .A1(keyinput9), .A2(keyinput127), .ZN(n8495) );
  NAND3_X1 U9971 ( .A1(keyinput105), .A2(keyinput74), .A3(n8495), .ZN(n8499)
         );
  NAND4_X1 U9972 ( .A1(keyinput40), .A2(keyinput99), .A3(keyinput26), .A4(
        keyinput20), .ZN(n8498) );
  OR4_X1 U9973 ( .A1(keyinput97), .A2(keyinput117), .A3(keyinput112), .A4(
        keyinput121), .ZN(n8497) );
  INV_X1 U9974 ( .A(keyinput54), .ZN(n8559) );
  NAND4_X1 U9975 ( .A1(keyinput21), .A2(keyinput101), .A3(keyinput73), .A4(
        n8559), .ZN(n8496) );
  NOR4_X1 U9976 ( .A1(n8499), .A2(n8498), .A3(n8497), .A4(n8496), .ZN(n8500)
         );
  NAND4_X1 U9977 ( .A1(n8503), .A2(n8502), .A3(n8501), .A4(n8500), .ZN(n8553)
         );
  NOR4_X1 U9978 ( .A1(keyinput10), .A2(keyinput7), .A3(keyinput30), .A4(
        keyinput42), .ZN(n8504) );
  NAND3_X1 U9979 ( .A1(keyinput84), .A2(keyinput64), .A3(n8504), .ZN(n8517) );
  NOR2_X1 U9980 ( .A1(keyinput58), .A2(keyinput65), .ZN(n8505) );
  NAND3_X1 U9981 ( .A1(keyinput33), .A2(keyinput56), .A3(n8505), .ZN(n8506) );
  NOR3_X1 U9982 ( .A1(keyinput43), .A2(keyinput38), .A3(n8506), .ZN(n8515) );
  INV_X1 U9983 ( .A(keyinput25), .ZN(n8507) );
  NAND4_X1 U9984 ( .A1(keyinput89), .A2(keyinput71), .A3(keyinput100), .A4(
        n8507), .ZN(n8513) );
  OR4_X1 U9985 ( .A1(keyinput76), .A2(keyinput126), .A3(keyinput17), .A4(
        keyinput62), .ZN(n8512) );
  NOR3_X1 U9986 ( .A1(keyinput107), .A2(keyinput113), .A3(keyinput87), .ZN(
        n8508) );
  NAND2_X1 U9987 ( .A1(keyinput83), .A2(n8508), .ZN(n8511) );
  INV_X1 U9988 ( .A(keyinput90), .ZN(n8509) );
  NAND4_X1 U9989 ( .A1(keyinput119), .A2(keyinput80), .A3(keyinput88), .A4(
        n8509), .ZN(n8510) );
  NOR4_X1 U9990 ( .A1(n8513), .A2(n8512), .A3(n8511), .A4(n8510), .ZN(n8514)
         );
  NAND4_X1 U9991 ( .A1(keyinput22), .A2(keyinput35), .A3(n8515), .A4(n8514), 
        .ZN(n8516) );
  NOR4_X1 U9992 ( .A1(keyinput104), .A2(keyinput3), .A3(n8517), .A4(n8516), 
        .ZN(n8551) );
  NAND2_X1 U9993 ( .A1(keyinput91), .A2(keyinput60), .ZN(n8518) );
  NOR3_X1 U9994 ( .A1(keyinput70), .A2(keyinput52), .A3(n8518), .ZN(n8519) );
  NAND3_X1 U9995 ( .A1(keyinput15), .A2(keyinput92), .A3(n8519), .ZN(n8532) );
  NOR2_X1 U9996 ( .A1(keyinput108), .A2(keyinput13), .ZN(n8520) );
  NAND3_X1 U9997 ( .A1(keyinput41), .A2(keyinput5), .A3(n8520), .ZN(n8521) );
  NOR3_X1 U9998 ( .A1(keyinput67), .A2(keyinput6), .A3(n8521), .ZN(n8530) );
  NOR2_X1 U9999 ( .A1(keyinput27), .A2(keyinput103), .ZN(n8522) );
  NAND3_X1 U10000 ( .A1(keyinput124), .A2(keyinput8), .A3(n8522), .ZN(n8528)
         );
  NOR2_X1 U10001 ( .A1(keyinput53), .A2(keyinput12), .ZN(n8523) );
  NAND3_X1 U10002 ( .A1(keyinput11), .A2(keyinput44), .A3(n8523), .ZN(n8527)
         );
  OR4_X1 U10003 ( .A1(keyinput1), .A2(keyinput48), .A3(keyinput37), .A4(
        keyinput86), .ZN(n8526) );
  INV_X1 U10004 ( .A(keyinput72), .ZN(n8524) );
  NAND4_X1 U10005 ( .A1(keyinput47), .A2(keyinput75), .A3(keyinput120), .A4(
        n8524), .ZN(n8525) );
  NOR4_X1 U10006 ( .A1(n8528), .A2(n8527), .A3(n8526), .A4(n8525), .ZN(n8529)
         );
  NAND4_X1 U10007 ( .A1(keyinput116), .A2(keyinput125), .A3(n8530), .A4(n8529), 
        .ZN(n8531) );
  NOR4_X1 U10008 ( .A1(keyinput122), .A2(keyinput66), .A3(n8532), .A4(n8531), 
        .ZN(n8550) );
  INV_X1 U10009 ( .A(keyinput32), .ZN(n8533) );
  NAND4_X1 U10010 ( .A1(keyinput93), .A2(keyinput2), .A3(keyinput95), .A4(
        n8533), .ZN(n8540) );
  NOR2_X1 U10011 ( .A1(keyinput68), .A2(keyinput29), .ZN(n8534) );
  NAND3_X1 U10012 ( .A1(keyinput31), .A2(keyinput50), .A3(n8534), .ZN(n8539)
         );
  NOR2_X1 U10013 ( .A1(keyinput14), .A2(keyinput46), .ZN(n8535) );
  NAND3_X1 U10014 ( .A1(keyinput98), .A2(keyinput34), .A3(n8535), .ZN(n8538)
         );
  INV_X1 U10015 ( .A(keyinput123), .ZN(n8536) );
  NAND4_X1 U10016 ( .A1(keyinput23), .A2(keyinput96), .A3(keyinput118), .A4(
        n8536), .ZN(n8537) );
  NOR4_X1 U10017 ( .A1(n8540), .A2(n8539), .A3(n8538), .A4(n8537), .ZN(n8549)
         );
  NOR3_X1 U10018 ( .A1(keyinput110), .A2(keyinput19), .A3(keyinput59), .ZN(
        n8541) );
  NAND2_X1 U10019 ( .A1(keyinput85), .A2(n8541), .ZN(n8547) );
  INV_X1 U10020 ( .A(keyinput49), .ZN(n8542) );
  NAND4_X1 U10021 ( .A1(keyinput16), .A2(keyinput102), .A3(keyinput55), .A4(
        n8542), .ZN(n8546) );
  NAND4_X1 U10022 ( .A1(keyinput111), .A2(keyinput82), .A3(keyinput69), .A4(
        keyinput18), .ZN(n8545) );
  NOR3_X1 U10023 ( .A1(keyinput0), .A2(keyinput45), .A3(keyinput79), .ZN(n8543) );
  NAND2_X1 U10024 ( .A1(keyinput63), .A2(n8543), .ZN(n8544) );
  NOR4_X1 U10025 ( .A1(n8547), .A2(n8546), .A3(n8545), .A4(n8544), .ZN(n8548)
         );
  NAND4_X1 U10026 ( .A1(n8551), .A2(n8550), .A3(n8549), .A4(n8548), .ZN(n8552)
         );
  OAI21_X1 U10027 ( .B1(n8553), .B2(n8552), .A(keyinput28), .ZN(n8775) );
  INV_X1 U10028 ( .A(keyinput117), .ZN(n8555) );
  OAI22_X1 U10029 ( .A1(n7435), .A2(keyinput112), .B1(n8555), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n8554) );
  AOI221_X1 U10030 ( .B1(n7435), .B2(keyinput112), .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n8555), .A(n8554), .ZN(n8566) );
  OAI22_X1 U10031 ( .A1(n8557), .A2(keyinput21), .B1(n7332), .B2(keyinput97), 
        .ZN(n8556) );
  AOI221_X1 U10032 ( .B1(n8557), .B2(keyinput21), .C1(keyinput97), .C2(n7332), 
        .A(n8556), .ZN(n8565) );
  OAI22_X1 U10033 ( .A1(keyinput73), .A2(n5939), .B1(n8559), .B2(
        P2_ADDR_REG_5__SCAN_IN), .ZN(n8558) );
  AOI221_X1 U10034 ( .B1(n5939), .B2(keyinput73), .C1(n8559), .C2(
        P2_ADDR_REG_5__SCAN_IN), .A(n8558), .ZN(n8564) );
  OAI22_X1 U10035 ( .A1(n8562), .A2(keyinput121), .B1(n8561), .B2(keyinput61), 
        .ZN(n8560) );
  AOI221_X1 U10036 ( .B1(n8562), .B2(keyinput121), .C1(keyinput61), .C2(n8561), 
        .A(n8560), .ZN(n8563) );
  AND4_X1 U10037 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(n8586)
         );
  AOI22_X1 U10038 ( .A1(n9116), .A2(keyinput38), .B1(keyinput33), .B2(n8568), 
        .ZN(n8567) );
  OAI221_X1 U10039 ( .B1(n9116), .B2(keyinput38), .C1(n8568), .C2(keyinput33), 
        .A(n8567), .ZN(n8571) );
  XNOR2_X1 U10040 ( .A(n8569), .B(keyinput51), .ZN(n8570) );
  NOR2_X1 U10041 ( .A1(n8571), .A2(n8570), .ZN(n8585) );
  AOI22_X1 U10042 ( .A1(n5175), .A2(keyinput85), .B1(n8573), .B2(keyinput68), 
        .ZN(n8572) );
  OAI221_X1 U10043 ( .B1(n5175), .B2(keyinput85), .C1(n8573), .C2(keyinput68), 
        .A(n8572), .ZN(n8578) );
  INV_X1 U10044 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8576) );
  AOI22_X1 U10045 ( .A1(n8576), .A2(keyinput47), .B1(keyinput120), .B2(n8575), 
        .ZN(n8574) );
  OAI221_X1 U10046 ( .B1(n8576), .B2(keyinput47), .C1(n8575), .C2(keyinput120), 
        .A(n8574), .ZN(n8577) );
  NOR2_X1 U10047 ( .A1(n8578), .A2(n8577), .ZN(n8584) );
  INV_X1 U10048 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U10049 ( .A1(n10103), .A2(keyinput99), .B1(keyinput26), .B2(n9477), 
        .ZN(n8579) );
  OAI221_X1 U10050 ( .B1(n10103), .B2(keyinput99), .C1(n9477), .C2(keyinput26), 
        .A(n8579), .ZN(n8582) );
  AOI22_X1 U10051 ( .A1(n9185), .A2(keyinput18), .B1(keyinput79), .B2(n8777), 
        .ZN(n8580) );
  OAI221_X1 U10052 ( .B1(n9185), .B2(keyinput18), .C1(n8777), .C2(keyinput79), 
        .A(n8580), .ZN(n8581) );
  NOR2_X1 U10053 ( .A1(n8582), .A2(n8581), .ZN(n8583) );
  NAND4_X1 U10054 ( .A1(n8586), .A2(n8585), .A3(n8584), .A4(n8583), .ZN(n8624)
         );
  AOI22_X1 U10055 ( .A1(n8589), .A2(keyinput114), .B1(keyinput39), .B2(n8588), 
        .ZN(n8587) );
  OAI221_X1 U10056 ( .B1(n8589), .B2(keyinput114), .C1(n8588), .C2(keyinput39), 
        .A(n8587), .ZN(n8596) );
  AOI22_X1 U10057 ( .A1(n9768), .A2(keyinput55), .B1(keyinput110), .B2(n8591), 
        .ZN(n8590) );
  OAI221_X1 U10058 ( .B1(n9768), .B2(keyinput55), .C1(n8591), .C2(keyinput110), 
        .A(n8590), .ZN(n8595) );
  AOI22_X1 U10059 ( .A1(n9254), .A2(keyinput6), .B1(n8593), .B2(keyinput49), 
        .ZN(n8592) );
  OAI221_X1 U10060 ( .B1(n9254), .B2(keyinput6), .C1(n8593), .C2(keyinput49), 
        .A(n8592), .ZN(n8594) );
  NOR3_X1 U10061 ( .A1(n8596), .A2(n8595), .A3(n8594), .ZN(n8622) );
  INV_X1 U10062 ( .A(SI_30_), .ZN(n8598) );
  AOI22_X1 U10063 ( .A1(n7297), .A2(keyinput119), .B1(keyinput107), .B2(n8598), 
        .ZN(n8597) );
  OAI221_X1 U10064 ( .B1(n7297), .B2(keyinput119), .C1(n8598), .C2(keyinput107), .A(n8597), .ZN(n8601) );
  INV_X1 U10065 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U10066 ( .A1(n10102), .A2(keyinput20), .B1(keyinput105), .B2(n9520), 
        .ZN(n8599) );
  OAI221_X1 U10067 ( .B1(n10102), .B2(keyinput20), .C1(n9520), .C2(keyinput105), .A(n8599), .ZN(n8600) );
  NOR2_X1 U10068 ( .A1(n8601), .A2(n8600), .ZN(n8621) );
  AOI22_X1 U10069 ( .A1(n8604), .A2(keyinput52), .B1(n8603), .B2(keyinput122), 
        .ZN(n8602) );
  OAI221_X1 U10070 ( .B1(n8604), .B2(keyinput52), .C1(n8603), .C2(keyinput122), 
        .A(n8602), .ZN(n8612) );
  AOI22_X1 U10071 ( .A1(n8607), .A2(keyinput31), .B1(n8606), .B2(keyinput50), 
        .ZN(n8605) );
  OAI221_X1 U10072 ( .B1(n8607), .B2(keyinput31), .C1(n8606), .C2(keyinput50), 
        .A(n8605), .ZN(n8611) );
  XNOR2_X1 U10073 ( .A(keyinput35), .B(P1_REG0_REG_5__SCAN_IN), .ZN(n8609) );
  XNOR2_X1 U10074 ( .A(keyinput7), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10075 ( .A1(n8609), .A2(n8608), .ZN(n8610) );
  NOR3_X1 U10076 ( .A1(n8612), .A2(n8611), .A3(n8610), .ZN(n8620) );
  AOI22_X1 U10077 ( .A1(n9778), .A2(keyinput113), .B1(keyinput60), .B2(n8614), 
        .ZN(n8613) );
  OAI221_X1 U10078 ( .B1(n9778), .B2(keyinput113), .C1(n8614), .C2(keyinput60), 
        .A(n8613), .ZN(n8618) );
  AOI22_X1 U10079 ( .A1(n8616), .A2(keyinput92), .B1(n6855), .B2(keyinput70), 
        .ZN(n8615) );
  OAI221_X1 U10080 ( .B1(n8616), .B2(keyinput92), .C1(n6855), .C2(keyinput70), 
        .A(n8615), .ZN(n8617) );
  NOR2_X1 U10081 ( .A1(n8618), .A2(n8617), .ZN(n8619) );
  NAND4_X1 U10082 ( .A1(n8622), .A2(n8621), .A3(n8620), .A4(n8619), .ZN(n8623)
         );
  NOR2_X1 U10083 ( .A1(n8624), .A2(n8623), .ZN(n8744) );
  AOI22_X1 U10084 ( .A1(n6701), .A2(keyinput23), .B1(n8626), .B2(keyinput96), 
        .ZN(n8625) );
  OAI221_X1 U10085 ( .B1(n6701), .B2(keyinput23), .C1(n8626), .C2(keyinput96), 
        .A(n8625), .ZN(n8634) );
  INV_X1 U10086 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8812) );
  AOI22_X1 U10087 ( .A1(n8877), .A2(keyinput118), .B1(keyinput14), .B2(n8812), 
        .ZN(n8627) );
  OAI221_X1 U10088 ( .B1(n8877), .B2(keyinput118), .C1(n8812), .C2(keyinput14), 
        .A(n8627), .ZN(n8633) );
  AOI22_X1 U10089 ( .A1(n7350), .A2(keyinput98), .B1(n8629), .B2(keyinput46), 
        .ZN(n8628) );
  OAI221_X1 U10090 ( .B1(n7350), .B2(keyinput98), .C1(n8629), .C2(keyinput46), 
        .A(n8628), .ZN(n8632) );
  INV_X1 U10091 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U10092 ( .A1(n6071), .A2(keyinput34), .B1(n10101), .B2(keyinput0), 
        .ZN(n8630) );
  OAI221_X1 U10093 ( .B1(n6071), .B2(keyinput34), .C1(n10101), .C2(keyinput0), 
        .A(n8630), .ZN(n8631) );
  NOR4_X1 U10094 ( .A1(n8634), .A2(n8633), .A3(n8632), .A4(n8631), .ZN(n8743)
         );
  AOI22_X1 U10095 ( .A1(n5825), .A2(keyinput13), .B1(n8636), .B2(keyinput67), 
        .ZN(n8635) );
  OAI221_X1 U10096 ( .B1(n5825), .B2(keyinput13), .C1(n8636), .C2(keyinput67), 
        .A(n8635), .ZN(n8641) );
  AOI22_X1 U10097 ( .A1(n8639), .A2(keyinput9), .B1(keyinput74), .B2(n8638), 
        .ZN(n8637) );
  OAI221_X1 U10098 ( .B1(n8639), .B2(keyinput9), .C1(n8638), .C2(keyinput74), 
        .A(n8637), .ZN(n8640) );
  NOR2_X1 U10099 ( .A1(n8641), .A2(n8640), .ZN(n8671) );
  AOI22_X1 U10100 ( .A1(n5177), .A2(keyinput78), .B1(n8643), .B2(keyinput36), 
        .ZN(n8642) );
  OAI221_X1 U10101 ( .B1(n5177), .B2(keyinput78), .C1(n8643), .C2(keyinput36), 
        .A(n8642), .ZN(n8648) );
  AOI22_X1 U10102 ( .A1(n8646), .A2(keyinput59), .B1(n8645), .B2(keyinput19), 
        .ZN(n8644) );
  OAI221_X1 U10103 ( .B1(n8646), .B2(keyinput59), .C1(n8645), .C2(keyinput19), 
        .A(n8644), .ZN(n8647) );
  NOR2_X1 U10104 ( .A1(n8648), .A2(n8647), .ZN(n8670) );
  XNOR2_X1 U10105 ( .A(SI_5_), .B(keyinput30), .ZN(n8652) );
  XNOR2_X1 U10106 ( .A(SI_7_), .B(keyinput37), .ZN(n8651) );
  XNOR2_X1 U10107 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput125), .ZN(n8650) );
  XNOR2_X1 U10108 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput127), .ZN(n8649)
         );
  NAND4_X1 U10109 ( .A1(n8652), .A2(n8651), .A3(n8650), .A4(n8649), .ZN(n8657)
         );
  XNOR2_X1 U10110 ( .A(SI_8_), .B(keyinput10), .ZN(n8655) );
  XNOR2_X1 U10111 ( .A(keyinput16), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n8654)
         );
  NAND2_X1 U10112 ( .A1(keyinput28), .A2(n9329), .ZN(n8653) );
  NAND3_X1 U10113 ( .A1(n8655), .A2(n8654), .A3(n8653), .ZN(n8656) );
  NOR2_X1 U10114 ( .A1(n8657), .A2(n8656), .ZN(n8669) );
  XNOR2_X1 U10115 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput64), .ZN(n8661) );
  XNOR2_X1 U10116 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput56), .ZN(n8660) );
  XNOR2_X1 U10117 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput123), .ZN(n8659) );
  XNOR2_X1 U10118 ( .A(P1_REG0_REG_23__SCAN_IN), .B(keyinput65), .ZN(n8658) );
  NAND4_X1 U10119 ( .A1(n8661), .A2(n8660), .A3(n8659), .A4(n8658), .ZN(n8667)
         );
  XNOR2_X1 U10120 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput102), .ZN(n8665) );
  XNOR2_X1 U10121 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput69), .ZN(n8664) );
  XNOR2_X1 U10122 ( .A(P1_REG1_REG_20__SCAN_IN), .B(keyinput76), .ZN(n8663) );
  XNOR2_X1 U10123 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput83), .ZN(n8662) );
  NAND4_X1 U10124 ( .A1(n8665), .A2(n8664), .A3(n8663), .A4(n8662), .ZN(n8666)
         );
  NOR2_X1 U10125 ( .A1(n8667), .A2(n8666), .ZN(n8668) );
  NAND4_X1 U10126 ( .A1(n8671), .A2(n8670), .A3(n8669), .A4(n8668), .ZN(n8686)
         );
  INV_X1 U10127 ( .A(keyinput77), .ZN(n8673) );
  OAI22_X1 U10128 ( .A1(keyinput24), .A2(n8674), .B1(n8673), .B2(
        P1_ADDR_REG_2__SCAN_IN), .ZN(n8672) );
  AOI221_X1 U10129 ( .B1(n8674), .B2(keyinput24), .C1(n8673), .C2(
        P1_ADDR_REG_2__SCAN_IN), .A(n8672), .ZN(n8684) );
  INV_X1 U10130 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10107) );
  OAI22_X1 U10131 ( .A1(n10107), .A2(keyinput4), .B1(n8834), .B2(keyinput57), 
        .ZN(n8675) );
  AOI221_X1 U10132 ( .B1(n10107), .B2(keyinput4), .C1(keyinput57), .C2(n8834), 
        .A(n8675), .ZN(n8683) );
  INV_X1 U10133 ( .A(keyinput81), .ZN(n8677) );
  OAI22_X1 U10134 ( .A1(n8678), .A2(keyinput104), .B1(n8677), .B2(
        P2_D_REG_13__SCAN_IN), .ZN(n8676) );
  AOI221_X1 U10135 ( .B1(n8678), .B2(keyinput104), .C1(P2_D_REG_13__SCAN_IN), 
        .C2(n8677), .A(n8676), .ZN(n8682) );
  OAI22_X1 U10136 ( .A1(n8680), .A2(keyinput106), .B1(n6636), .B2(keyinput94), 
        .ZN(n8679) );
  AOI221_X1 U10137 ( .B1(n8680), .B2(keyinput106), .C1(keyinput94), .C2(n6636), 
        .A(n8679), .ZN(n8681) );
  NAND4_X1 U10138 ( .A1(n8684), .A2(n8683), .A3(n8682), .A4(n8681), .ZN(n8685)
         );
  NOR2_X1 U10139 ( .A1(n8686), .A2(n8685), .ZN(n8742) );
  INV_X1 U10140 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U10141 ( .A1(n6179), .A2(keyinput86), .B1(n10105), .B2(keyinput116), 
        .ZN(n8687) );
  OAI221_X1 U10142 ( .B1(n6179), .B2(keyinput86), .C1(n10105), .C2(keyinput116), .A(n8687), .ZN(n8690) );
  INV_X1 U10143 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8889) );
  AOI22_X1 U10144 ( .A1(n8889), .A2(keyinput66), .B1(n6707), .B2(keyinput15), 
        .ZN(n8688) );
  OAI221_X1 U10145 ( .B1(n8889), .B2(keyinput66), .C1(n6707), .C2(keyinput15), 
        .A(n8688), .ZN(n8689) );
  NOR2_X1 U10146 ( .A1(n8690), .A2(n8689), .ZN(n8712) );
  INV_X1 U10147 ( .A(keyinput108), .ZN(n8692) );
  AOI22_X1 U10148 ( .A1(n8693), .A2(keyinput5), .B1(P2_ADDR_REG_6__SCAN_IN), 
        .B2(n8692), .ZN(n8691) );
  OAI221_X1 U10149 ( .B1(n8693), .B2(keyinput5), .C1(n8692), .C2(
        P2_ADDR_REG_6__SCAN_IN), .A(n8691), .ZN(n8698) );
  AOI22_X1 U10150 ( .A1(n8696), .A2(keyinput42), .B1(n8695), .B2(keyinput43), 
        .ZN(n8694) );
  OAI221_X1 U10151 ( .B1(n8696), .B2(keyinput42), .C1(n8695), .C2(keyinput43), 
        .A(n8694), .ZN(n8697) );
  NOR2_X1 U10152 ( .A1(n8698), .A2(n8697), .ZN(n8711) );
  AOI22_X1 U10153 ( .A1(n5828), .A2(keyinput109), .B1(n6873), .B2(keyinput45), 
        .ZN(n8699) );
  OAI221_X1 U10154 ( .B1(n5828), .B2(keyinput109), .C1(n6873), .C2(keyinput45), 
        .A(n8699), .ZN(n8702) );
  AOI22_X1 U10155 ( .A1(n8842), .A2(keyinput87), .B1(n6852), .B2(keyinput90), 
        .ZN(n8700) );
  OAI221_X1 U10156 ( .B1(n8842), .B2(keyinput87), .C1(n6852), .C2(keyinput90), 
        .A(n8700), .ZN(n8701) );
  NOR2_X1 U10157 ( .A1(n8702), .A2(n8701), .ZN(n8710) );
  AOI22_X1 U10158 ( .A1(n8704), .A2(keyinput93), .B1(n7781), .B2(keyinput32), 
        .ZN(n8703) );
  OAI221_X1 U10159 ( .B1(n8704), .B2(keyinput93), .C1(n7781), .C2(keyinput32), 
        .A(n8703), .ZN(n8708) );
  AOI22_X1 U10160 ( .A1(n5352), .A2(keyinput72), .B1(keyinput1), .B2(n8706), 
        .ZN(n8705) );
  OAI221_X1 U10161 ( .B1(n5352), .B2(keyinput72), .C1(n8706), .C2(keyinput1), 
        .A(n8705), .ZN(n8707) );
  NOR2_X1 U10162 ( .A1(n8708), .A2(n8707), .ZN(n8709) );
  NAND4_X1 U10163 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), .ZN(n8740)
         );
  XNOR2_X1 U10164 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(keyinput53), .ZN(n8716)
         );
  XNOR2_X1 U10165 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput84), .ZN(n8715) );
  XNOR2_X1 U10166 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput22), .ZN(n8714) );
  XNOR2_X1 U10167 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput3), .ZN(n8713) );
  NAND4_X1 U10168 ( .A1(n8716), .A2(n8715), .A3(n8714), .A4(n8713), .ZN(n8722)
         );
  XNOR2_X1 U10169 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput115), .ZN(n8720) );
  XNOR2_X1 U10170 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput111), .ZN(n8719) );
  XNOR2_X1 U10171 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput2), .ZN(n8718) );
  XNOR2_X1 U10172 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput91), .ZN(n8717) );
  NAND4_X1 U10173 ( .A1(n8720), .A2(n8719), .A3(n8718), .A4(n8717), .ZN(n8721)
         );
  NOR2_X1 U10174 ( .A1(n8722), .A2(n8721), .ZN(n8738) );
  INV_X1 U10175 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10104) );
  INV_X1 U10176 ( .A(keyinput88), .ZN(n8723) );
  XNOR2_X1 U10177 ( .A(n10104), .B(n8723), .ZN(n8737) );
  INV_X1 U10178 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10108) );
  INV_X1 U10179 ( .A(keyinput41), .ZN(n8724) );
  XNOR2_X1 U10180 ( .A(n10108), .B(n8724), .ZN(n8736) );
  XNOR2_X1 U10181 ( .A(P2_REG0_REG_18__SCAN_IN), .B(keyinput82), .ZN(n8728) );
  XNOR2_X1 U10182 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput63), .ZN(n8727) );
  XNOR2_X1 U10183 ( .A(P2_REG1_REG_23__SCAN_IN), .B(keyinput48), .ZN(n8726) );
  XNOR2_X1 U10184 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput58), .ZN(n8725) );
  NAND4_X1 U10185 ( .A1(n8728), .A2(n8727), .A3(n8726), .A4(n8725), .ZN(n8734)
         );
  XNOR2_X1 U10186 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput101), .ZN(n8732)
         );
  XNOR2_X1 U10187 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput40), .ZN(n8731) );
  XNOR2_X1 U10188 ( .A(keyinput95), .B(P1_REG0_REG_17__SCAN_IN), .ZN(n8730) );
  XNOR2_X1 U10189 ( .A(keyinput29), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n8729) );
  NAND4_X1 U10190 ( .A1(n8732), .A2(n8731), .A3(n8730), .A4(n8729), .ZN(n8733)
         );
  NOR2_X1 U10191 ( .A1(n8734), .A2(n8733), .ZN(n8735) );
  NAND4_X1 U10192 ( .A1(n8738), .A2(n8737), .A3(n8736), .A4(n8735), .ZN(n8739)
         );
  NOR2_X1 U10193 ( .A1(n8740), .A2(n8739), .ZN(n8741) );
  NAND4_X1 U10194 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(n8774)
         );
  AOI22_X1 U10195 ( .A1(n8854), .A2(keyinput89), .B1(n8746), .B2(keyinput17), 
        .ZN(n8745) );
  OAI221_X1 U10196 ( .B1(n8854), .B2(keyinput89), .C1(n8746), .C2(keyinput17), 
        .A(n8745), .ZN(n8757) );
  AOI22_X1 U10197 ( .A1(n8748), .A2(keyinput126), .B1(keyinput71), .B2(n7363), 
        .ZN(n8747) );
  OAI221_X1 U10198 ( .B1(n8748), .B2(keyinput126), .C1(n7363), .C2(keyinput71), 
        .A(n8747), .ZN(n8756) );
  INV_X1 U10199 ( .A(keyinput80), .ZN(n8750) );
  AOI22_X1 U10200 ( .A1(n7298), .A2(keyinput100), .B1(P2_ADDR_REG_1__SCAN_IN), 
        .B2(n8750), .ZN(n8749) );
  OAI221_X1 U10201 ( .B1(n7298), .B2(keyinput100), .C1(n8750), .C2(
        P2_ADDR_REG_1__SCAN_IN), .A(n8749), .ZN(n8755) );
  INV_X1 U10202 ( .A(keyinput62), .ZN(n8752) );
  AOI22_X1 U10203 ( .A1(n8753), .A2(keyinput25), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n8752), .ZN(n8751) );
  OAI221_X1 U10204 ( .B1(n8753), .B2(keyinput25), .C1(n8752), .C2(
        P1_ADDR_REG_16__SCAN_IN), .A(n8751), .ZN(n8754) );
  NOR4_X1 U10205 ( .A1(n8757), .A2(n8756), .A3(n8755), .A4(n8754), .ZN(n8772)
         );
  INV_X1 U10206 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U10207 ( .A1(n10276), .A2(keyinput11), .B1(n8759), .B2(keyinput12), 
        .ZN(n8758) );
  OAI221_X1 U10208 ( .B1(n10276), .B2(keyinput11), .C1(n8759), .C2(keyinput12), 
        .A(n8758), .ZN(n8770) );
  AOI22_X1 U10209 ( .A1(n8762), .A2(keyinput44), .B1(keyinput27), .B2(n8761), 
        .ZN(n8760) );
  OAI221_X1 U10210 ( .B1(n8762), .B2(keyinput44), .C1(n8761), .C2(keyinput27), 
        .A(n8760), .ZN(n8769) );
  AOI22_X1 U10211 ( .A1(n7396), .A2(keyinput124), .B1(n8764), .B2(keyinput8), 
        .ZN(n8763) );
  OAI221_X1 U10212 ( .B1(n7396), .B2(keyinput124), .C1(n8764), .C2(keyinput8), 
        .A(n8763), .ZN(n8768) );
  INV_X1 U10213 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U10214 ( .A1(n8766), .A2(keyinput103), .B1(n10106), .B2(keyinput75), 
        .ZN(n8765) );
  OAI221_X1 U10215 ( .B1(n8766), .B2(keyinput103), .C1(n10106), .C2(keyinput75), .A(n8765), .ZN(n8767) );
  NOR4_X1 U10216 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n8771)
         );
  NAND2_X1 U10217 ( .A1(n8772), .A2(n8771), .ZN(n8773) );
  AOI211_X1 U10218 ( .C1(n8775), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n8774), .B(
        n8773), .ZN(n8785) );
  MUX2_X1 U10219 ( .A(n8777), .B(n8776), .S(n10233), .Z(n8781) );
  AOI22_X1 U10220 ( .A1(n4556), .A2(n10226), .B1(n10228), .B2(n8778), .ZN(
        n8780) );
  OAI211_X1 U10221 ( .C1(n8783), .C2(n8782), .A(n8781), .B(n8780), .ZN(n8784)
         );
  XOR2_X1 U10222 ( .A(n8785), .B(n8784), .Z(P2_U3222) );
  INV_X1 U10223 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U10224 ( .A1(n8786), .A2(n8843), .ZN(n8788) );
  INV_X1 U10225 ( .A(n8847), .ZN(n8787) );
  NAND2_X1 U10226 ( .A1(n8787), .A2(n10289), .ZN(n8791) );
  OAI211_X1 U10227 ( .C1(n10289), .C2(n8789), .A(n8788), .B(n8791), .ZN(
        P2_U3490) );
  INV_X1 U10228 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U10229 ( .A1(n8790), .A2(n8843), .ZN(n8792) );
  OAI211_X1 U10230 ( .C1(n10289), .C2(n8793), .A(n8792), .B(n8791), .ZN(
        P2_U3489) );
  INV_X1 U10231 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8794) );
  MUX2_X1 U10232 ( .A(n8794), .B(n8853), .S(n10289), .Z(n8796) );
  NAND2_X1 U10233 ( .A1(n8855), .A2(n8843), .ZN(n8795) );
  OAI211_X1 U10234 ( .C1(n8858), .C2(n8837), .A(n8796), .B(n8795), .ZN(
        P2_U3486) );
  MUX2_X1 U10235 ( .A(n8797), .B(n8859), .S(n10289), .Z(n8799) );
  NAND2_X1 U10236 ( .A1(n8861), .A2(n8843), .ZN(n8798) );
  OAI211_X1 U10237 ( .C1(n8837), .C2(n8864), .A(n8799), .B(n8798), .ZN(
        P2_U3485) );
  MUX2_X1 U10238 ( .A(n8800), .B(n8865), .S(n10289), .Z(n8802) );
  NAND2_X1 U10239 ( .A1(n8867), .A2(n8843), .ZN(n8801) );
  OAI211_X1 U10240 ( .C1(n8837), .C2(n8870), .A(n8802), .B(n8801), .ZN(
        P2_U3484) );
  MUX2_X1 U10241 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8871), .S(n10289), .Z(
        n8805) );
  INV_X1 U10242 ( .A(n8803), .ZN(n8873) );
  OAI22_X1 U10243 ( .A1(n8873), .A2(n8837), .B1(n8872), .B2(n8831), .ZN(n8804)
         );
  OR2_X1 U10244 ( .A1(n8805), .A2(n8804), .ZN(P2_U3483) );
  INV_X1 U10245 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8806) );
  MUX2_X1 U10246 ( .A(n8806), .B(n8876), .S(n10289), .Z(n8808) );
  NAND2_X1 U10247 ( .A1(n8878), .A2(n8843), .ZN(n8807) );
  OAI211_X1 U10248 ( .C1(n8881), .C2(n8837), .A(n8808), .B(n8807), .ZN(
        P2_U3482) );
  INV_X1 U10249 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8809) );
  MUX2_X1 U10250 ( .A(n8809), .B(n8882), .S(n10289), .Z(n8811) );
  NAND2_X1 U10251 ( .A1(n8884), .A2(n8843), .ZN(n8810) );
  OAI211_X1 U10252 ( .C1(n8837), .C2(n8887), .A(n8811), .B(n8810), .ZN(
        P2_U3481) );
  MUX2_X1 U10253 ( .A(n8812), .B(n8888), .S(n10289), .Z(n8814) );
  NAND2_X1 U10254 ( .A1(n8890), .A2(n8843), .ZN(n8813) );
  OAI211_X1 U10255 ( .C1(n8837), .C2(n8893), .A(n8814), .B(n8813), .ZN(
        P2_U3480) );
  INV_X1 U10256 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8816) );
  INV_X1 U10257 ( .A(n8815), .ZN(n8894) );
  MUX2_X1 U10258 ( .A(n8816), .B(n8894), .S(n10289), .Z(n8818) );
  INV_X1 U10259 ( .A(n8837), .ZN(n8844) );
  AOI22_X1 U10260 ( .A1(n8897), .A2(n8844), .B1(n8843), .B2(n8896), .ZN(n8817)
         );
  NAND2_X1 U10261 ( .A1(n8818), .A2(n8817), .ZN(P2_U3479) );
  NAND2_X1 U10262 ( .A1(n8819), .A2(n10244), .ZN(n8820) );
  OAI211_X1 U10263 ( .C1(n10263), .C2(n8822), .A(n8821), .B(n8820), .ZN(n8900)
         );
  MUX2_X1 U10264 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8900), .S(n10289), .Z(
        P2_U3478) );
  MUX2_X1 U10265 ( .A(n8823), .B(n8901), .S(n10289), .Z(n8825) );
  NAND2_X1 U10266 ( .A1(n8903), .A2(n8843), .ZN(n8824) );
  OAI211_X1 U10267 ( .C1(n8837), .C2(n8906), .A(n8825), .B(n8824), .ZN(
        P2_U3477) );
  AOI22_X1 U10268 ( .A1(n8827), .A2(n10274), .B1(n10244), .B2(n8826), .ZN(
        n8828) );
  NAND2_X1 U10269 ( .A1(n8829), .A2(n8828), .ZN(n8907) );
  MUX2_X1 U10270 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8907), .S(n10289), .Z(
        P2_U3476) );
  MUX2_X1 U10271 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8908), .S(n10289), .Z(
        n8833) );
  INV_X1 U10272 ( .A(n8830), .ZN(n8910) );
  OAI22_X1 U10273 ( .A1(n8911), .A2(n8837), .B1(n8910), .B2(n8831), .ZN(n8832)
         );
  OR2_X1 U10274 ( .A1(n8833), .A2(n8832), .ZN(P2_U3475) );
  MUX2_X1 U10275 ( .A(n8834), .B(n8914), .S(n10289), .Z(n8836) );
  NAND2_X1 U10276 ( .A1(n8916), .A2(n8843), .ZN(n8835) );
  OAI211_X1 U10277 ( .C1(n8920), .C2(n8837), .A(n8836), .B(n8835), .ZN(
        P2_U3474) );
  MUX2_X1 U10278 ( .A(n8838), .B(n8921), .S(n10289), .Z(n8840) );
  AOI22_X1 U10279 ( .A1(n8924), .A2(n8844), .B1(n8843), .B2(n8923), .ZN(n8839)
         );
  NAND2_X1 U10280 ( .A1(n8840), .A2(n8839), .ZN(P2_U3473) );
  INV_X1 U10281 ( .A(n8841), .ZN(n8927) );
  MUX2_X1 U10282 ( .A(n8842), .B(n8927), .S(n10289), .Z(n8846) );
  AOI22_X1 U10283 ( .A1(n8932), .A2(n8844), .B1(n8843), .B2(n8929), .ZN(n8845)
         );
  NAND2_X1 U10284 ( .A1(n8846), .A2(n8845), .ZN(P2_U3472) );
  NOR2_X1 U10285 ( .A1(n8847), .A2(n10277), .ZN(n8850) );
  AOI21_X1 U10286 ( .B1(n10277), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8850), .ZN(
        n8848) );
  OAI21_X1 U10287 ( .B1(n8849), .B2(n8909), .A(n8848), .ZN(P2_U3458) );
  AOI21_X1 U10288 ( .B1(n10277), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8850), .ZN(
        n8851) );
  OAI21_X1 U10289 ( .B1(n8852), .B2(n8909), .A(n8851), .ZN(P2_U3457) );
  MUX2_X1 U10290 ( .A(n8854), .B(n8853), .S(n10275), .Z(n8857) );
  NAND2_X1 U10291 ( .A1(n8855), .A2(n8930), .ZN(n8856) );
  OAI211_X1 U10292 ( .C1(n8858), .C2(n8919), .A(n8857), .B(n8856), .ZN(
        P2_U3454) );
  INV_X1 U10293 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8860) );
  MUX2_X1 U10294 ( .A(n8860), .B(n8859), .S(n10275), .Z(n8863) );
  NAND2_X1 U10295 ( .A1(n8861), .A2(n8930), .ZN(n8862) );
  OAI211_X1 U10296 ( .C1(n8864), .C2(n8919), .A(n8863), .B(n8862), .ZN(
        P2_U3453) );
  INV_X1 U10297 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8866) );
  MUX2_X1 U10298 ( .A(n8866), .B(n8865), .S(n10275), .Z(n8869) );
  NAND2_X1 U10299 ( .A1(n8867), .A2(n8930), .ZN(n8868) );
  OAI211_X1 U10300 ( .C1(n8870), .C2(n8919), .A(n8869), .B(n8868), .ZN(
        P2_U3452) );
  MUX2_X1 U10301 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8871), .S(n10275), .Z(
        n8875) );
  OAI22_X1 U10302 ( .A1(n8873), .A2(n8919), .B1(n8872), .B2(n8909), .ZN(n8874)
         );
  OR2_X1 U10303 ( .A1(n8875), .A2(n8874), .ZN(P2_U3451) );
  MUX2_X1 U10304 ( .A(n8877), .B(n8876), .S(n10275), .Z(n8880) );
  NAND2_X1 U10305 ( .A1(n8878), .A2(n8930), .ZN(n8879) );
  OAI211_X1 U10306 ( .C1(n8881), .C2(n8919), .A(n8880), .B(n8879), .ZN(
        P2_U3450) );
  INV_X1 U10307 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8883) );
  MUX2_X1 U10308 ( .A(n8883), .B(n8882), .S(n10275), .Z(n8886) );
  NAND2_X1 U10309 ( .A1(n8884), .A2(n8930), .ZN(n8885) );
  OAI211_X1 U10310 ( .C1(n8887), .C2(n8919), .A(n8886), .B(n8885), .ZN(
        P2_U3449) );
  MUX2_X1 U10311 ( .A(n8889), .B(n8888), .S(n10275), .Z(n8892) );
  NAND2_X1 U10312 ( .A1(n8890), .A2(n8930), .ZN(n8891) );
  OAI211_X1 U10313 ( .C1(n8893), .C2(n8919), .A(n8892), .B(n8891), .ZN(
        P2_U3448) );
  INV_X1 U10314 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U10315 ( .A(n8895), .B(n8894), .S(n10275), .Z(n8899) );
  INV_X1 U10316 ( .A(n8919), .ZN(n8931) );
  AOI22_X1 U10317 ( .A1(n8897), .A2(n8931), .B1(n8930), .B2(n8896), .ZN(n8898)
         );
  NAND2_X1 U10318 ( .A1(n8899), .A2(n8898), .ZN(P2_U3447) );
  MUX2_X1 U10319 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8900), .S(n10275), .Z(
        P2_U3446) );
  INV_X1 U10320 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8902) );
  MUX2_X1 U10321 ( .A(n8902), .B(n8901), .S(n10275), .Z(n8905) );
  NAND2_X1 U10322 ( .A1(n8903), .A2(n8930), .ZN(n8904) );
  OAI211_X1 U10323 ( .C1(n8906), .C2(n8919), .A(n8905), .B(n8904), .ZN(
        P2_U3444) );
  MUX2_X1 U10324 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8907), .S(n10275), .Z(
        P2_U3441) );
  MUX2_X1 U10325 ( .A(n8908), .B(P2_REG0_REG_16__SCAN_IN), .S(n10277), .Z(
        n8913) );
  OAI22_X1 U10326 ( .A1(n8911), .A2(n8919), .B1(n8910), .B2(n8909), .ZN(n8912)
         );
  OR2_X1 U10327 ( .A1(n8913), .A2(n8912), .ZN(P2_U3438) );
  INV_X1 U10328 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8915) );
  MUX2_X1 U10329 ( .A(n8915), .B(n8914), .S(n10275), .Z(n8918) );
  NAND2_X1 U10330 ( .A1(n8916), .A2(n8930), .ZN(n8917) );
  OAI211_X1 U10331 ( .C1(n8920), .C2(n8919), .A(n8918), .B(n8917), .ZN(
        P2_U3435) );
  INV_X1 U10332 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8922) );
  MUX2_X1 U10333 ( .A(n8922), .B(n8921), .S(n10275), .Z(n8926) );
  AOI22_X1 U10334 ( .A1(n8924), .A2(n8931), .B1(n8930), .B2(n8923), .ZN(n8925)
         );
  NAND2_X1 U10335 ( .A1(n8926), .A2(n8925), .ZN(P2_U3432) );
  INV_X1 U10336 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8928) );
  MUX2_X1 U10337 ( .A(n8928), .B(n8927), .S(n10275), .Z(n8934) );
  AOI22_X1 U10338 ( .A1(n8932), .A2(n8931), .B1(n8930), .B2(n8929), .ZN(n8933)
         );
  NAND2_X1 U10339 ( .A1(n8934), .A2(n8933), .ZN(P2_U3429) );
  MUX2_X1 U10340 ( .A(P2_D_REG_1__SCAN_IN), .B(n8936), .S(n8935), .Z(P2_U3377)
         );
  INV_X1 U10341 ( .A(n8937), .ZN(n9762) );
  NOR4_X1 U10342 ( .A1(n5199), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5405), .ZN(n8938) );
  AOI21_X1 U10343 ( .B1(n8939), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8938), .ZN(
        n8940) );
  OAI21_X1 U10344 ( .B1(n9762), .B2(n8954), .A(n8940), .ZN(P2_U3264) );
  INV_X1 U10345 ( .A(n7259), .ZN(n9766) );
  OAI222_X1 U10346 ( .A1(n8954), .A2(n9766), .B1(n8942), .B2(P2_U3151), .C1(
        n8941), .C2(n8951), .ZN(P2_U3266) );
  NAND2_X1 U10347 ( .A1(n9770), .A2(n8946), .ZN(n8944) );
  OAI211_X1 U10348 ( .C1(n8951), .C2(n8945), .A(n8944), .B(n8943), .ZN(
        P2_U3267) );
  NAND2_X1 U10349 ( .A1(n8947), .A2(n8946), .ZN(n8949) );
  OAI211_X1 U10350 ( .C1(n8951), .C2(n8950), .A(n8949), .B(n8948), .ZN(
        P2_U3268) );
  INV_X1 U10351 ( .A(n8952), .ZN(n9776) );
  OAI222_X1 U10352 ( .A1(n8954), .A2(n9776), .B1(P2_U3151), .B2(n4575), .C1(
        n8953), .C2(n8951), .ZN(P2_U3269) );
  MUX2_X1 U10353 ( .A(n8955), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10354 ( .A(n9697), .ZN(n9507) );
  NAND2_X1 U10355 ( .A1(n10002), .A2(n9127), .ZN(n8961) );
  NAND2_X1 U10356 ( .A1(n8963), .A2(n9121), .ZN(n8960) );
  NAND2_X1 U10357 ( .A1(n8961), .A2(n8960), .ZN(n8962) );
  XNOR2_X1 U10358 ( .A(n8962), .B(n9075), .ZN(n8964) );
  AOI22_X1 U10359 ( .A1(n10002), .A2(n9121), .B1(n6421), .B2(n8963), .ZN(n8965) );
  XNOR2_X1 U10360 ( .A(n8964), .B(n8965), .ZN(n9227) );
  INV_X1 U10361 ( .A(n8964), .ZN(n8966) );
  AOI22_X1 U10362 ( .A1(n9156), .A2(n9121), .B1(n6421), .B2(n9274), .ZN(n8970)
         );
  NAND2_X1 U10363 ( .A1(n9156), .A2(n9127), .ZN(n8968) );
  NAND2_X1 U10364 ( .A1(n9274), .A2(n9121), .ZN(n8967) );
  NAND2_X1 U10365 ( .A1(n8968), .A2(n8967), .ZN(n8969) );
  XNOR2_X1 U10366 ( .A(n8969), .B(n9075), .ZN(n8972) );
  XOR2_X1 U10367 ( .A(n8970), .B(n8972), .Z(n9149) );
  INV_X1 U10368 ( .A(n8970), .ZN(n8971) );
  NAND2_X1 U10369 ( .A1(n9984), .A2(n9127), .ZN(n8974) );
  NAND2_X1 U10370 ( .A1(n9417), .A2(n9121), .ZN(n8973) );
  NAND2_X1 U10371 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  XNOR2_X1 U10372 ( .A(n8975), .B(n9075), .ZN(n8976) );
  AOI22_X1 U10373 ( .A1(n9984), .A2(n9121), .B1(n6421), .B2(n9417), .ZN(n8977)
         );
  XNOR2_X1 U10374 ( .A(n8976), .B(n8977), .ZN(n9213) );
  INV_X1 U10375 ( .A(n8976), .ZN(n8978) );
  NAND2_X1 U10376 ( .A1(n9674), .A2(n9127), .ZN(n8980) );
  NAND2_X1 U10377 ( .A1(n9418), .A2(n9121), .ZN(n8979) );
  NAND2_X1 U10378 ( .A1(n8980), .A2(n8979), .ZN(n8981) );
  XNOR2_X1 U10379 ( .A(n8981), .B(n9075), .ZN(n8983) );
  INV_X1 U10380 ( .A(n8983), .ZN(n8982) );
  AOI22_X1 U10381 ( .A1(n9674), .A2(n9121), .B1(n6421), .B2(n9418), .ZN(n9092)
         );
  OR2_X1 U10382 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  NAND2_X1 U10383 ( .A1(n9656), .A2(n9127), .ZN(n8987) );
  NAND2_X1 U10384 ( .A1(n9273), .A2(n9121), .ZN(n8986) );
  NAND2_X1 U10385 ( .A1(n8987), .A2(n8986), .ZN(n8988) );
  XNOR2_X1 U10386 ( .A(n8988), .B(n9075), .ZN(n9171) );
  AOI22_X1 U10387 ( .A1(n9656), .A2(n9121), .B1(n6421), .B2(n9273), .ZN(n9170)
         );
  INV_X1 U10388 ( .A(n9170), .ZN(n8997) );
  NAND2_X1 U10389 ( .A1(n4437), .A2(n9121), .ZN(n8990) );
  NAND2_X1 U10390 ( .A1(n9421), .A2(n6421), .ZN(n8989) );
  NAND2_X1 U10391 ( .A1(n4436), .A2(n9127), .ZN(n8992) );
  NAND2_X1 U10392 ( .A1(n9421), .A2(n9121), .ZN(n8991) );
  NAND2_X1 U10393 ( .A1(n8992), .A2(n8991), .ZN(n8993) );
  INV_X1 U10394 ( .A(n9169), .ZN(n8996) );
  AOI22_X1 U10395 ( .A1(n9171), .A2(n8997), .B1(n9260), .B2(n8996), .ZN(n9000)
         );
  AOI21_X1 U10396 ( .B1(n9169), .B2(n8994), .A(n9170), .ZN(n8995) );
  NOR2_X1 U10397 ( .A1(n8995), .A2(n9171), .ZN(n8999) );
  NAND2_X1 U10398 ( .A1(n9825), .A2(n9127), .ZN(n9002) );
  NAND2_X1 U10399 ( .A1(n9424), .A2(n9121), .ZN(n9001) );
  NAND2_X1 U10400 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  XNOR2_X1 U10401 ( .A(n9003), .B(n9125), .ZN(n9006) );
  AND2_X1 U10402 ( .A1(n9424), .A2(n6421), .ZN(n9004) );
  AOI21_X1 U10403 ( .B1(n9825), .B2(n9121), .A(n9004), .ZN(n9005) );
  NOR2_X1 U10404 ( .A1(n9006), .A2(n9005), .ZN(n9180) );
  NAND2_X1 U10405 ( .A1(n9641), .A2(n9127), .ZN(n9008) );
  NAND2_X1 U10406 ( .A1(n9429), .A2(n9121), .ZN(n9007) );
  NAND2_X1 U10407 ( .A1(n9008), .A2(n9007), .ZN(n9009) );
  XNOR2_X1 U10408 ( .A(n9009), .B(n9125), .ZN(n9011) );
  AOI22_X1 U10409 ( .A1(n9641), .A2(n9121), .B1(n6421), .B2(n9429), .ZN(n9010)
         );
  AND2_X1 U10410 ( .A1(n9011), .A2(n9010), .ZN(n9236) );
  OR2_X1 U10411 ( .A1(n9011), .A2(n9010), .ZN(n9237) );
  NAND2_X1 U10412 ( .A1(n9737), .A2(n9127), .ZN(n9013) );
  NAND2_X1 U10413 ( .A1(n9431), .A2(n9121), .ZN(n9012) );
  NAND2_X1 U10414 ( .A1(n9013), .A2(n9012), .ZN(n9014) );
  XNOR2_X1 U10415 ( .A(n9014), .B(n9125), .ZN(n9016) );
  AOI22_X1 U10416 ( .A1(n9737), .A2(n9121), .B1(n6421), .B2(n9431), .ZN(n9015)
         );
  NOR2_X1 U10417 ( .A1(n9016), .A2(n9015), .ZN(n9111) );
  NAND2_X1 U10418 ( .A1(n9733), .A2(n9127), .ZN(n9018) );
  NAND2_X1 U10419 ( .A1(n9435), .A2(n9121), .ZN(n9017) );
  NAND2_X1 U10420 ( .A1(n9018), .A2(n9017), .ZN(n9019) );
  XNOR2_X1 U10421 ( .A(n9019), .B(n9075), .ZN(n9023) );
  NAND2_X1 U10422 ( .A1(n9733), .A2(n9121), .ZN(n9021) );
  NAND2_X1 U10423 ( .A1(n9435), .A2(n6421), .ZN(n9020) );
  NAND2_X1 U10424 ( .A1(n9021), .A2(n9020), .ZN(n9022) );
  NOR2_X1 U10425 ( .A1(n9023), .A2(n9022), .ZN(n9024) );
  AOI21_X1 U10426 ( .B1(n9023), .B2(n9022), .A(n9024), .ZN(n9203) );
  INV_X1 U10427 ( .A(n9024), .ZN(n9025) );
  NAND2_X1 U10428 ( .A1(n9728), .A2(n9127), .ZN(n9027) );
  NAND2_X1 U10429 ( .A1(n9438), .A2(n9121), .ZN(n9026) );
  NAND2_X1 U10430 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  XNOR2_X1 U10431 ( .A(n9028), .B(n9075), .ZN(n9031) );
  AOI22_X1 U10432 ( .A1(n9728), .A2(n9121), .B1(n6421), .B2(n9438), .ZN(n9029)
         );
  XNOR2_X1 U10433 ( .A(n9031), .B(n9029), .ZN(n9142) );
  INV_X1 U10434 ( .A(n9029), .ZN(n9030) );
  AOI22_X1 U10435 ( .A1(n9723), .A2(n9127), .B1(n9121), .B2(n9442), .ZN(n9033)
         );
  XNOR2_X1 U10436 ( .A(n9033), .B(n9075), .ZN(n9034) );
  INV_X1 U10437 ( .A(n9034), .ZN(n9035) );
  OAI22_X1 U10438 ( .A1(n9575), .A2(n5045), .B1(n9441), .B2(n4435), .ZN(n9220)
         );
  INV_X1 U10439 ( .A(n9036), .ZN(n9105) );
  NAND2_X1 U10440 ( .A1(n9717), .A2(n9127), .ZN(n9038) );
  NAND2_X1 U10441 ( .A1(n9443), .A2(n9121), .ZN(n9037) );
  NAND2_X1 U10442 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  XNOR2_X1 U10443 ( .A(n9039), .B(n9125), .ZN(n9041) );
  AND2_X1 U10444 ( .A1(n9443), .A2(n6421), .ZN(n9040) );
  AOI21_X1 U10445 ( .B1(n9717), .B2(n9121), .A(n9040), .ZN(n9042) );
  NAND2_X1 U10446 ( .A1(n9041), .A2(n9042), .ZN(n9190) );
  INV_X1 U10447 ( .A(n9041), .ZN(n9044) );
  INV_X1 U10448 ( .A(n9042), .ZN(n9043) );
  NAND2_X1 U10449 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  AND2_X1 U10450 ( .A1(n9190), .A2(n9045), .ZN(n9104) );
  NAND2_X1 U10451 ( .A1(n9102), .A2(n9190), .ZN(n9055) );
  NAND2_X1 U10452 ( .A1(n9713), .A2(n9127), .ZN(n9047) );
  NAND2_X1 U10453 ( .A1(n9272), .A2(n9121), .ZN(n9046) );
  NAND2_X1 U10454 ( .A1(n9047), .A2(n9046), .ZN(n9048) );
  XNOR2_X1 U10455 ( .A(n9048), .B(n9125), .ZN(n9050) );
  AND2_X1 U10456 ( .A1(n9272), .A2(n6421), .ZN(n9049) );
  AOI21_X1 U10457 ( .B1(n9713), .B2(n9121), .A(n9049), .ZN(n9051) );
  NAND2_X1 U10458 ( .A1(n9050), .A2(n9051), .ZN(n9056) );
  INV_X1 U10459 ( .A(n9050), .ZN(n9053) );
  INV_X1 U10460 ( .A(n9051), .ZN(n9052) );
  NAND2_X1 U10461 ( .A1(n9053), .A2(n9052), .ZN(n9054) );
  INV_X1 U10462 ( .A(n9707), .ZN(n9536) );
  OAI22_X1 U10463 ( .A1(n9536), .A2(n5045), .B1(n9057), .B2(n4435), .ZN(n9066)
         );
  NAND2_X1 U10464 ( .A1(n9707), .A2(n9127), .ZN(n9059) );
  NAND2_X1 U10465 ( .A1(n9451), .A2(n9121), .ZN(n9058) );
  NAND2_X1 U10466 ( .A1(n9059), .A2(n9058), .ZN(n9060) );
  XNOR2_X1 U10467 ( .A(n9060), .B(n9075), .ZN(n9065) );
  XOR2_X1 U10468 ( .A(n9066), .B(n9065), .Z(n9161) );
  NAND2_X1 U10469 ( .A1(n9703), .A2(n9127), .ZN(n9062) );
  NAND2_X1 U10470 ( .A1(n9271), .A2(n9121), .ZN(n9061) );
  NAND2_X1 U10471 ( .A1(n9062), .A2(n9061), .ZN(n9063) );
  XNOR2_X1 U10472 ( .A(n9063), .B(n9075), .ZN(n9072) );
  AND2_X1 U10473 ( .A1(n9271), .A2(n6421), .ZN(n9064) );
  AOI21_X1 U10474 ( .B1(n9703), .B2(n9121), .A(n9064), .ZN(n9070) );
  XNOR2_X1 U10475 ( .A(n9072), .B(n9070), .ZN(n9248) );
  INV_X1 U10476 ( .A(n9065), .ZN(n9068) );
  INV_X1 U10477 ( .A(n9066), .ZN(n9067) );
  NAND2_X1 U10478 ( .A1(n9068), .A2(n9067), .ZN(n9245) );
  INV_X1 U10479 ( .A(n9070), .ZN(n9071) );
  NAND2_X1 U10480 ( .A1(n9072), .A2(n9071), .ZN(n9082) );
  NAND2_X1 U10481 ( .A1(n9697), .A2(n9127), .ZN(n9074) );
  NAND2_X1 U10482 ( .A1(n9456), .A2(n9121), .ZN(n9073) );
  NAND2_X1 U10483 ( .A1(n9074), .A2(n9073), .ZN(n9076) );
  XNOR2_X1 U10484 ( .A(n9076), .B(n9075), .ZN(n9080) );
  NAND2_X1 U10485 ( .A1(n9697), .A2(n9121), .ZN(n9078) );
  NAND2_X1 U10486 ( .A1(n9456), .A2(n6421), .ZN(n9077) );
  NAND2_X1 U10487 ( .A1(n9078), .A2(n9077), .ZN(n9079) );
  NOR2_X1 U10488 ( .A1(n9080), .A2(n9079), .ZN(n9134) );
  AOI21_X1 U10489 ( .B1(n9080), .B2(n9079), .A(n9134), .ZN(n9081) );
  AOI21_X1 U10490 ( .B1(n9246), .B2(n9082), .A(n9081), .ZN(n9086) );
  INV_X1 U10491 ( .A(n9081), .ZN(n9084) );
  INV_X1 U10492 ( .A(n9082), .ZN(n9083) );
  NOR2_X1 U10493 ( .A1(n9084), .A2(n9083), .ZN(n9085) );
  OAI22_X1 U10494 ( .A1(n9474), .A2(n9406), .B1(n9454), .B2(n9475), .ZN(n9510)
         );
  OAI22_X1 U10495 ( .A1(n9504), .A2(n9264), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9087), .ZN(n9088) );
  AOI21_X1 U10496 ( .B1(n9510), .B2(n9262), .A(n9088), .ZN(n9089) );
  OAI211_X1 U10497 ( .C1(n9507), .C2(n9258), .A(n9090), .B(n9089), .ZN(
        P1_U3214) );
  OAI21_X1 U10498 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9094) );
  NAND2_X1 U10499 ( .A1(n9094), .A2(n9247), .ZN(n9101) );
  INV_X1 U10500 ( .A(n9669), .ZN(n9099) );
  NAND2_X1 U10501 ( .A1(n9421), .A2(n9250), .ZN(n9096) );
  NAND2_X1 U10502 ( .A1(n9417), .A2(n9251), .ZN(n9095) );
  AND2_X1 U10503 ( .A1(n9096), .A2(n9095), .ZN(n9668) );
  OAI22_X1 U10504 ( .A1(n9668), .A2(n9222), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9097), .ZN(n9098) );
  AOI21_X1 U10505 ( .B1(n9099), .B2(n9210), .A(n9098), .ZN(n9100) );
  OAI211_X1 U10506 ( .C1(n10195), .C2(n9258), .A(n9101), .B(n9100), .ZN(
        P1_U3215) );
  INV_X1 U10507 ( .A(n9102), .ZN(n9193) );
  NOR3_X1 U10508 ( .A1(n4580), .A2(n9105), .A3(n9104), .ZN(n9106) );
  OAI21_X1 U10509 ( .B1(n9193), .B2(n9106), .A(n9247), .ZN(n9110) );
  OAI22_X1 U10510 ( .A1(n9447), .A2(n9406), .B1(n9441), .B2(n9475), .ZN(n9567)
         );
  OAI22_X1 U10511 ( .A1(n9264), .A2(n9561), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9107), .ZN(n9108) );
  AOI21_X1 U10512 ( .B1(n9567), .B2(n9262), .A(n9108), .ZN(n9109) );
  OAI211_X1 U10513 ( .C1(n4581), .C2(n9258), .A(n9110), .B(n9109), .ZN(
        P1_U3216) );
  NOR2_X1 U10514 ( .A1(n9111), .A2(n4518), .ZN(n9112) );
  XNOR2_X1 U10515 ( .A(n9113), .B(n9112), .ZN(n9120) );
  NAND2_X1 U10516 ( .A1(n9435), .A2(n9250), .ZN(n9115) );
  NAND2_X1 U10517 ( .A1(n9429), .A2(n9251), .ZN(n9114) );
  NAND2_X1 U10518 ( .A1(n9115), .A2(n9114), .ZN(n9625) );
  NOR2_X1 U10519 ( .A1(n9116), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9400) );
  AOI21_X1 U10520 ( .B1(n9625), .B2(n9262), .A(n9400), .ZN(n9117) );
  OAI21_X1 U10521 ( .B1(n9264), .B2(n9618), .A(n9117), .ZN(n9118) );
  AOI21_X1 U10522 ( .B1(n9737), .B2(n9266), .A(n9118), .ZN(n9119) );
  OAI21_X1 U10523 ( .B1(n9120), .B2(n9268), .A(n9119), .ZN(P1_U3219) );
  NAND2_X1 U10524 ( .A1(n9692), .A2(n9121), .ZN(n9124) );
  OR2_X1 U10525 ( .A1(n9474), .A2(n4435), .ZN(n9123) );
  NAND2_X1 U10526 ( .A1(n9124), .A2(n9123), .ZN(n9126) );
  XNOR2_X1 U10527 ( .A(n9126), .B(n9125), .ZN(n9130) );
  NAND2_X1 U10528 ( .A1(n9692), .A2(n9127), .ZN(n9128) );
  OAI21_X1 U10529 ( .B1(n9474), .B2(n5045), .A(n9128), .ZN(n9129) );
  XNOR2_X1 U10530 ( .A(n9130), .B(n9129), .ZN(n9135) );
  OR4_X2 U10531 ( .A1(n9131), .A2(n9134), .A3(n9135), .A4(n9268), .ZN(n9139)
         );
  AOI22_X1 U10532 ( .A1(n9456), .A2(n9251), .B1(n9250), .B2(n9270), .ZN(n9494)
         );
  AOI22_X1 U10533 ( .A1(n9497), .A2(n9210), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9132) );
  OAI21_X1 U10534 ( .B1(n9494), .B2(n9222), .A(n9132), .ZN(n9133) );
  AOI21_X1 U10535 ( .B1(n9692), .B2(n9266), .A(n9133), .ZN(n9137) );
  NAND3_X1 U10536 ( .A1(n9135), .A2(n9134), .A3(n9247), .ZN(n9136) );
  NAND4_X1 U10537 ( .A1(n9139), .A2(n9138), .A3(n9137), .A4(n9136), .ZN(
        P1_U3220) );
  INV_X1 U10538 ( .A(n9728), .ZN(n9598) );
  OAI21_X1 U10539 ( .B1(n9142), .B2(n9141), .A(n9140), .ZN(n9143) );
  NAND2_X1 U10540 ( .A1(n9143), .A2(n9247), .ZN(n9148) );
  INV_X1 U10541 ( .A(n9144), .ZN(n9595) );
  AOI22_X1 U10542 ( .A1(n9442), .A2(n9250), .B1(n9251), .B2(n9435), .ZN(n9592)
         );
  OAI22_X1 U10543 ( .A1(n9592), .A2(n9222), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9145), .ZN(n9146) );
  AOI21_X1 U10544 ( .B1(n9595), .B2(n9210), .A(n9146), .ZN(n9147) );
  OAI211_X1 U10545 ( .C1(n9598), .C2(n9258), .A(n9148), .B(n9147), .ZN(
        P1_U3223) );
  XOR2_X1 U10546 ( .A(n9150), .B(n9149), .Z(n9158) );
  NAND2_X1 U10547 ( .A1(n9151), .A2(n9262), .ZN(n9153) );
  OAI211_X1 U10548 ( .C1(n9264), .C2(n9154), .A(n9153), .B(n9152), .ZN(n9155)
         );
  AOI21_X1 U10549 ( .B1(n9156), .B2(n9266), .A(n9155), .ZN(n9157) );
  OAI21_X1 U10550 ( .B1(n9158), .B2(n9268), .A(n9157), .ZN(P1_U3224) );
  OAI21_X1 U10551 ( .B1(n9161), .B2(n9160), .A(n9159), .ZN(n9162) );
  NAND2_X1 U10552 ( .A1(n9162), .A2(n9247), .ZN(n9167) );
  OAI22_X1 U10553 ( .A1(n9454), .A2(n9406), .B1(n9447), .B2(n9475), .ZN(n9539)
         );
  INV_X1 U10554 ( .A(n9534), .ZN(n9164) );
  OAI22_X1 U10555 ( .A1(n9164), .A2(n9264), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9163), .ZN(n9165) );
  AOI21_X1 U10556 ( .B1(n9539), .B2(n9262), .A(n9165), .ZN(n9166) );
  OAI211_X1 U10557 ( .C1(n9536), .C2(n9258), .A(n9167), .B(n9166), .ZN(
        P1_U3225) );
  XNOR2_X1 U10558 ( .A(n9169), .B(n9168), .ZN(n9261) );
  NOR2_X1 U10559 ( .A1(n9261), .A2(n9260), .ZN(n9259) );
  AOI21_X1 U10560 ( .B1(n9169), .B2(n9168), .A(n9259), .ZN(n9173) );
  XNOR2_X1 U10561 ( .A(n9171), .B(n9170), .ZN(n9172) );
  XNOR2_X1 U10562 ( .A(n9173), .B(n9172), .ZN(n9179) );
  NAND2_X1 U10563 ( .A1(n9424), .A2(n9250), .ZN(n9175) );
  NAND2_X1 U10564 ( .A1(n9421), .A2(n9251), .ZN(n9174) );
  NAND2_X1 U10565 ( .A1(n9175), .A2(n9174), .ZN(n9647) );
  AOI22_X1 U10566 ( .A1(n9647), .A2(n9262), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n9176) );
  OAI21_X1 U10567 ( .B1(n9264), .B2(n9652), .A(n9176), .ZN(n9177) );
  AOI21_X1 U10568 ( .B1(n4578), .B2(n9266), .A(n9177), .ZN(n9178) );
  OAI21_X1 U10569 ( .B1(n9179), .B2(n9268), .A(n9178), .ZN(P1_U3226) );
  NOR2_X1 U10570 ( .A1(n9180), .A2(n4527), .ZN(n9181) );
  XNOR2_X1 U10571 ( .A(n9182), .B(n9181), .ZN(n9189) );
  NAND2_X1 U10572 ( .A1(n9273), .A2(n9251), .ZN(n9184) );
  NAND2_X1 U10573 ( .A1(n9429), .A2(n9250), .ZN(n9183) );
  NAND2_X1 U10574 ( .A1(n9184), .A2(n9183), .ZN(n9820) );
  NOR2_X1 U10575 ( .A1(n9185), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9380) );
  AOI21_X1 U10576 ( .B1(n9820), .B2(n9262), .A(n9380), .ZN(n9186) );
  OAI21_X1 U10577 ( .B1(n9264), .B2(n9823), .A(n9186), .ZN(n9187) );
  AOI21_X1 U10578 ( .B1(n9825), .B2(n9266), .A(n9187), .ZN(n9188) );
  OAI21_X1 U10579 ( .B1(n9189), .B2(n9268), .A(n9188), .ZN(P1_U3228) );
  INV_X1 U10580 ( .A(n9190), .ZN(n9192) );
  NOR3_X1 U10581 ( .A1(n9193), .A2(n9192), .A3(n9191), .ZN(n9196) );
  INV_X1 U10582 ( .A(n9194), .ZN(n9195) );
  OAI21_X1 U10583 ( .B1(n9196), .B2(n9195), .A(n9247), .ZN(n9200) );
  AOI22_X1 U10584 ( .A1(n9451), .A2(n9250), .B1(n9251), .B2(n9443), .ZN(n9547)
         );
  OAI22_X1 U10585 ( .A1(n9547), .A2(n9222), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9197), .ZN(n9198) );
  AOI21_X1 U10586 ( .B1(n9553), .B2(n9210), .A(n9198), .ZN(n9199) );
  OAI211_X1 U10587 ( .C1(n9556), .C2(n9258), .A(n9200), .B(n9199), .ZN(
        P1_U3229) );
  OAI21_X1 U10588 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n9204) );
  NAND2_X1 U10589 ( .A1(n9204), .A2(n9247), .ZN(n9212) );
  INV_X1 U10590 ( .A(n9205), .ZN(n9610) );
  NAND2_X1 U10591 ( .A1(n9438), .A2(n9250), .ZN(n9207) );
  NAND2_X1 U10592 ( .A1(n9431), .A2(n9251), .ZN(n9206) );
  AND2_X1 U10593 ( .A1(n9207), .A2(n9206), .ZN(n9605) );
  OAI22_X1 U10594 ( .A1(n9605), .A2(n9222), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9208), .ZN(n9209) );
  AOI21_X1 U10595 ( .B1(n9610), .B2(n9210), .A(n9209), .ZN(n9211) );
  OAI211_X1 U10596 ( .C1(n9613), .C2(n9258), .A(n9212), .B(n9211), .ZN(
        P1_U3233) );
  XOR2_X1 U10597 ( .A(n9214), .B(n9213), .Z(n9218) );
  OAI22_X1 U10598 ( .A1(n9419), .A2(n9406), .B1(n9414), .B2(n9475), .ZN(n9978)
         );
  AOI22_X1 U10599 ( .A1(n9978), .A2(n9262), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n9215) );
  OAI21_X1 U10600 ( .B1(n9264), .B2(n9980), .A(n9215), .ZN(n9216) );
  AOI21_X1 U10601 ( .B1(n9984), .B2(n9266), .A(n9216), .ZN(n9217) );
  OAI21_X1 U10602 ( .B1(n9218), .B2(n9268), .A(n9217), .ZN(P1_U3234) );
  AOI21_X1 U10603 ( .B1(n9220), .B2(n9219), .A(n4580), .ZN(n9226) );
  NOR2_X1 U10604 ( .A1(n9264), .A2(n9576), .ZN(n9224) );
  AOI22_X1 U10605 ( .A1(n9443), .A2(n9250), .B1(n9251), .B2(n9438), .ZN(n9583)
         );
  OAI22_X1 U10606 ( .A1(n9583), .A2(n9222), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9221), .ZN(n9223) );
  AOI211_X1 U10607 ( .C1(n9723), .C2(n9266), .A(n9224), .B(n9223), .ZN(n9225)
         );
  OAI21_X1 U10608 ( .B1(n9226), .B2(n9268), .A(n9225), .ZN(P1_U3235) );
  XOR2_X1 U10609 ( .A(n9228), .B(n9227), .Z(n9234) );
  NAND2_X1 U10610 ( .A1(n9274), .A2(n9250), .ZN(n9230) );
  NAND2_X1 U10611 ( .A1(n9275), .A2(n9251), .ZN(n9229) );
  NAND2_X1 U10612 ( .A1(n9230), .A2(n9229), .ZN(n9997) );
  AOI22_X1 U10613 ( .A1(n9997), .A2(n9262), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n9231) );
  OAI21_X1 U10614 ( .B1(n9264), .B2(n9999), .A(n9231), .ZN(n9232) );
  AOI21_X1 U10615 ( .B1(n10002), .B2(n9266), .A(n9232), .ZN(n9233) );
  OAI21_X1 U10616 ( .B1(n9234), .B2(n9268), .A(n9233), .ZN(P1_U3236) );
  NAND2_X1 U10617 ( .A1(n4899), .A2(n9237), .ZN(n9238) );
  XNOR2_X1 U10618 ( .A(n9235), .B(n9238), .ZN(n9244) );
  NAND2_X1 U10619 ( .A1(n9424), .A2(n9251), .ZN(n9240) );
  NAND2_X1 U10620 ( .A1(n9431), .A2(n9250), .ZN(n9239) );
  NAND2_X1 U10621 ( .A1(n9240), .A2(n9239), .ZN(n9632) );
  AOI22_X1 U10622 ( .A1(n9632), .A2(n9262), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9241) );
  OAI21_X1 U10623 ( .B1(n9264), .B2(n9636), .A(n9241), .ZN(n9242) );
  AOI21_X1 U10624 ( .B1(n9641), .B2(n9266), .A(n9242), .ZN(n9243) );
  OAI21_X1 U10625 ( .B1(n9244), .B2(n9268), .A(n9243), .ZN(P1_U3238) );
  AND2_X1 U10626 ( .A1(n9159), .A2(n9245), .ZN(n9249) );
  OAI211_X1 U10627 ( .C1(n9249), .C2(n9248), .A(n9247), .B(n9246), .ZN(n9257)
         );
  NAND2_X1 U10628 ( .A1(n9456), .A2(n9250), .ZN(n9253) );
  NAND2_X1 U10629 ( .A1(n9451), .A2(n9251), .ZN(n9252) );
  NAND2_X1 U10630 ( .A1(n9253), .A2(n9252), .ZN(n9527) );
  OAI22_X1 U10631 ( .A1(n9521), .A2(n9264), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9254), .ZN(n9255) );
  AOI21_X1 U10632 ( .B1(n9527), .B2(n9262), .A(n9255), .ZN(n9256) );
  OAI211_X1 U10633 ( .C1(n9519), .C2(n9258), .A(n9257), .B(n9256), .ZN(
        P1_U3240) );
  AOI21_X1 U10634 ( .B1(n9261), .B2(n9260), .A(n9259), .ZN(n9269) );
  OAI22_X1 U10635 ( .A1(n9423), .A2(n9406), .B1(n9419), .B2(n9475), .ZN(n9836)
         );
  AOI22_X1 U10636 ( .A1(n9836), .A2(n9262), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9263) );
  OAI21_X1 U10637 ( .B1(n9264), .B2(n9838), .A(n9263), .ZN(n9265) );
  AOI21_X1 U10638 ( .B1(n4437), .B2(n9266), .A(n9265), .ZN(n9267) );
  OAI21_X1 U10639 ( .B1(n9269), .B2(n9268), .A(n9267), .ZN(P1_U3241) );
  MUX2_X1 U10640 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9270), .S(P1_U3973), .Z(
        P1_U3583) );
  INV_X1 U10641 ( .A(n9474), .ZN(n9457) );
  MUX2_X1 U10642 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9457), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10643 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9456), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10644 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9271), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10645 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9451), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10646 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9272), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10647 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9443), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10648 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9442), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10649 ( .A(n9438), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9284), .Z(
        P1_U3575) );
  MUX2_X1 U10650 ( .A(n9429), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9284), .Z(
        P1_U3572) );
  MUX2_X1 U10651 ( .A(n9424), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9284), .Z(
        P1_U3571) );
  MUX2_X1 U10652 ( .A(n9273), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9284), .Z(
        P1_U3570) );
  MUX2_X1 U10653 ( .A(n9421), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9284), .Z(
        P1_U3569) );
  MUX2_X1 U10654 ( .A(n9418), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9284), .Z(
        P1_U3568) );
  MUX2_X1 U10655 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9274), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10656 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9275), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10657 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9276), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10658 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9277), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10659 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9278), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10660 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9279), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10661 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9280), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10662 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9281), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10663 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9282), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10664 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9283), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10665 ( .A(n6285), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9284), .Z(
        P1_U3554) );
  OAI211_X1 U10666 ( .C1(n9287), .C2(n9286), .A(n9961), .B(n9285), .ZN(n9295)
         );
  OAI211_X1 U10667 ( .C1(n9290), .C2(n9289), .A(n9948), .B(n9288), .ZN(n9294)
         );
  AOI22_X1 U10668 ( .A1(n9883), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9293) );
  NAND2_X1 U10669 ( .A1(n9969), .A2(n9291), .ZN(n9292) );
  NAND4_X1 U10670 ( .A1(n9295), .A2(n9294), .A3(n9293), .A4(n9292), .ZN(
        P1_U3244) );
  INV_X1 U10671 ( .A(n9296), .ZN(n9300) );
  INV_X1 U10672 ( .A(n9883), .ZN(n9972) );
  INV_X1 U10673 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U10674 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9297) );
  OAI21_X1 U10675 ( .B1(n9972), .B2(n9298), .A(n9297), .ZN(n9299) );
  AOI21_X1 U10676 ( .B1(n9300), .B2(n9969), .A(n9299), .ZN(n9309) );
  OAI211_X1 U10677 ( .C1(n9303), .C2(n9302), .A(n9948), .B(n9301), .ZN(n9308)
         );
  OAI211_X1 U10678 ( .C1(n9306), .C2(n9305), .A(n9961), .B(n9304), .ZN(n9307)
         );
  NAND3_X1 U10679 ( .A1(n9309), .A2(n9308), .A3(n9307), .ZN(P1_U3246) );
  NAND2_X1 U10680 ( .A1(n9883), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9310) );
  OAI211_X1 U10681 ( .C1(n9952), .C2(n9312), .A(n9311), .B(n9310), .ZN(n9313)
         );
  INV_X1 U10682 ( .A(n9313), .ZN(n9322) );
  OAI211_X1 U10683 ( .C1(n9316), .C2(n9315), .A(n9961), .B(n9314), .ZN(n9321)
         );
  OAI211_X1 U10684 ( .C1(n9319), .C2(n9318), .A(n9948), .B(n9317), .ZN(n9320)
         );
  NAND4_X1 U10685 ( .A1(n9323), .A2(n9322), .A3(n9321), .A4(n9320), .ZN(
        P1_U3247) );
  AOI211_X1 U10686 ( .C1(n9326), .C2(n9325), .A(n9324), .B(n9958), .ZN(n9327)
         );
  INV_X1 U10687 ( .A(n9327), .ZN(n9337) );
  NAND2_X1 U10688 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9328) );
  OAI21_X1 U10689 ( .B1(n9972), .B2(n9329), .A(n9328), .ZN(n9330) );
  AOI21_X1 U10690 ( .B1(n9331), .B2(n9969), .A(n9330), .ZN(n9336) );
  OAI211_X1 U10691 ( .C1(n9334), .C2(n9333), .A(n9961), .B(n9332), .ZN(n9335)
         );
  NAND3_X1 U10692 ( .A1(n9337), .A2(n9336), .A3(n9335), .ZN(P1_U3248) );
  AOI211_X1 U10693 ( .C1(n9340), .C2(n9339), .A(n9958), .B(n9338), .ZN(n9341)
         );
  INV_X1 U10694 ( .A(n9341), .ZN(n9351) );
  INV_X1 U10695 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9343) );
  NAND2_X1 U10696 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9342) );
  OAI21_X1 U10697 ( .B1(n9972), .B2(n9343), .A(n9342), .ZN(n9344) );
  AOI21_X1 U10698 ( .B1(n9345), .B2(n9969), .A(n9344), .ZN(n9350) );
  OAI211_X1 U10699 ( .C1(n9348), .C2(n9347), .A(n9961), .B(n9346), .ZN(n9349)
         );
  NAND3_X1 U10700 ( .A1(n9351), .A2(n9350), .A3(n9349), .ZN(P1_U3249) );
  AOI22_X1 U10701 ( .A1(n9389), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n7317), .B2(
        n9378), .ZN(n9363) );
  OR2_X1 U10702 ( .A1(n9939), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U10703 ( .A1(n9939), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9352) );
  AND2_X1 U10704 ( .A1(n9353), .A2(n9352), .ZN(n9945) );
  INV_X1 U10705 ( .A(n9935), .ZN(n9370) );
  NAND2_X1 U10706 ( .A1(n9911), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9359) );
  NOR2_X1 U10707 ( .A1(n9355), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9354) );
  AOI21_X1 U10708 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n9355), .A(n9354), .ZN(
        n9900) );
  OAI21_X1 U10709 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9368), .A(n9356), .ZN(
        n9901) );
  NOR2_X1 U10710 ( .A1(n9900), .A2(n9901), .ZN(n9899) );
  MUX2_X1 U10711 ( .A(n9357), .B(P1_REG1_REG_14__SCAN_IN), .S(n9911), .Z(n9913) );
  NOR2_X1 U10712 ( .A1(n9914), .A2(n9913), .ZN(n9912) );
  INV_X1 U10713 ( .A(n9912), .ZN(n9358) );
  NAND2_X1 U10714 ( .A1(n9359), .A2(n9358), .ZN(n9360) );
  XNOR2_X1 U10715 ( .A(n9370), .B(n9360), .ZN(n9927) );
  AND2_X1 U10716 ( .A1(n9360), .A2(n9935), .ZN(n9361) );
  NAND2_X1 U10717 ( .A1(n9945), .A2(n9946), .ZN(n9944) );
  OAI21_X1 U10718 ( .B1(n9939), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9944), .ZN(
        n9362) );
  NAND2_X1 U10719 ( .A1(n9363), .A2(n9362), .ZN(n9384) );
  OAI21_X1 U10720 ( .B1(n9363), .B2(n9362), .A(n9384), .ZN(n9364) );
  INV_X1 U10721 ( .A(n9364), .ZN(n9383) );
  NOR2_X1 U10722 ( .A1(n9389), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9365) );
  AOI21_X1 U10723 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9389), .A(n9365), .ZN(
        n9376) );
  NAND2_X1 U10724 ( .A1(n9907), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9366) );
  OAI21_X1 U10725 ( .B1(n9907), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9366), .ZN(
        n9903) );
  OAI21_X1 U10726 ( .B1(n9368), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9367), .ZN(
        n9904) );
  NOR2_X1 U10727 ( .A1(n9903), .A2(n9904), .ZN(n9902) );
  NAND2_X1 U10728 ( .A1(n9911), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9369) );
  OAI21_X1 U10729 ( .B1(n9911), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9369), .ZN(
        n9918) );
  NOR2_X1 U10730 ( .A1(n9917), .A2(n9918), .ZN(n9916) );
  NOR2_X1 U10731 ( .A1(n9371), .A2(n9370), .ZN(n9373) );
  AOI21_X1 U10732 ( .B1(n9371), .B2(n9370), .A(n9373), .ZN(n9372) );
  INV_X1 U10733 ( .A(n9372), .ZN(n9932) );
  NOR2_X1 U10734 ( .A1(n9373), .A2(n9931), .ZN(n9941) );
  NAND2_X1 U10735 ( .A1(n9939), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9374) );
  OAI21_X1 U10736 ( .B1(n9939), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9374), .ZN(
        n9942) );
  NOR2_X1 U10737 ( .A1(n9941), .A2(n9942), .ZN(n9940) );
  AOI21_X1 U10738 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9939), .A(n9940), .ZN(
        n9375) );
  NAND2_X1 U10739 ( .A1(n9376), .A2(n9375), .ZN(n9388) );
  OAI21_X1 U10740 ( .B1(n9376), .B2(n9375), .A(n9388), .ZN(n9377) );
  NAND2_X1 U10741 ( .A1(n9377), .A2(n9961), .ZN(n9382) );
  NOR2_X1 U10742 ( .A1(n9952), .A2(n9378), .ZN(n9379) );
  AOI211_X1 U10743 ( .C1(n9883), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9380), .B(
        n9379), .ZN(n9381) );
  OAI211_X1 U10744 ( .C1(n9958), .C2(n9383), .A(n9382), .B(n9381), .ZN(
        P1_U3260) );
  OAI21_X1 U10745 ( .B1(n9389), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9384), .ZN(
        n9959) );
  NOR2_X1 U10746 ( .A1(n9968), .A2(n9385), .ZN(n9386) );
  AOI21_X1 U10747 ( .B1(n9968), .B2(n9385), .A(n9386), .ZN(n9960) );
  NOR2_X1 U10748 ( .A1(n9959), .A2(n9960), .ZN(n9957) );
  XNOR2_X1 U10749 ( .A(n9387), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9394) );
  OR2_X1 U10750 ( .A1(n9968), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U10751 ( .A1(n9968), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9391) );
  AND2_X1 U10752 ( .A1(n9390), .A2(n9391), .ZN(n9963) );
  NAND2_X1 U10753 ( .A1(n9964), .A2(n9963), .ZN(n9962) );
  NAND2_X1 U10754 ( .A1(n9962), .A2(n9391), .ZN(n9392) );
  XNOR2_X1 U10755 ( .A(n9392), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U10756 ( .A1(n9396), .A2(n9961), .ZN(n9393) );
  OAI211_X1 U10757 ( .C1(n9958), .C2(n9394), .A(n9393), .B(n9952), .ZN(n9398)
         );
  INV_X1 U10758 ( .A(n9394), .ZN(n9395) );
  OAI22_X1 U10759 ( .A1(n9396), .A2(n9930), .B1(n9395), .B2(n9958), .ZN(n9397)
         );
  INV_X1 U10760 ( .A(n9401), .ZN(P1_U3262) );
  NAND2_X1 U10761 ( .A1(n9843), .A2(n9862), .ZN(n9828) );
  NAND2_X1 U10762 ( .A1(n9829), .A2(n9851), .ZN(n9638) );
  NAND2_X1 U10763 ( .A1(n9560), .A2(n9556), .ZN(n9550) );
  INV_X1 U10764 ( .A(n9692), .ZN(n9490) );
  NAND2_X1 U10765 ( .A1(n9476), .A2(n9684), .ZN(n9410) );
  XNOR2_X1 U10766 ( .A(n9678), .B(n9410), .ZN(n9402) );
  NAND2_X1 U10767 ( .A1(n9402), .A2(n10081), .ZN(n9677) );
  INV_X1 U10768 ( .A(P1_B_REG_SCAN_IN), .ZN(n9403) );
  NOR2_X1 U10769 ( .A1(n9404), .A2(n9403), .ZN(n9405) );
  OR2_X1 U10770 ( .A1(n9406), .A2(n9405), .ZN(n9473) );
  OR2_X1 U10771 ( .A1(n9407), .A2(n9473), .ZN(n9682) );
  NOR2_X1 U10772 ( .A1(n9682), .A2(n10100), .ZN(n9412) );
  NOR2_X1 U10773 ( .A1(n9678), .A2(n9621), .ZN(n9408) );
  AOI211_X1 U10774 ( .C1(n10100), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9412), .B(
        n9408), .ZN(n9409) );
  OAI21_X1 U10775 ( .B1(n9677), .B2(n9671), .A(n9409), .ZN(P1_U3263) );
  OAI211_X1 U10776 ( .C1(n9684), .C2(n9476), .A(n10081), .B(n9410), .ZN(n9683)
         );
  NOR2_X1 U10777 ( .A1(n9684), .A2(n9621), .ZN(n9411) );
  AOI211_X1 U10778 ( .C1(n10100), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9412), .B(
        n9411), .ZN(n9413) );
  OAI21_X1 U10779 ( .B1(n9671), .B2(n9683), .A(n9413), .ZN(P1_U3264) );
  INV_X1 U10780 ( .A(n9825), .ZN(n9856) );
  INV_X1 U10781 ( .A(n4438), .ZN(n9868) );
  NOR2_X1 U10782 ( .A1(n9674), .A2(n9418), .ZN(n9420) );
  NAND2_X1 U10783 ( .A1(n9650), .A2(n9649), .ZN(n9864) );
  NAND2_X1 U10784 ( .A1(n9864), .A2(n5046), .ZN(n9827) );
  NAND2_X1 U10785 ( .A1(n9827), .A2(n9425), .ZN(n9426) );
  OAI21_X1 U10786 ( .B1(n9856), .B2(n9427), .A(n9426), .ZN(n9634) );
  NAND2_X1 U10787 ( .A1(n9851), .A2(n9428), .ZN(n9430) );
  NAND2_X1 U10788 ( .A1(n9737), .A2(n9431), .ZN(n9433) );
  AOI22_X2 U10789 ( .A1(n9616), .A2(n9433), .B1(n9622), .B2(n9432), .ZN(n9602)
         );
  NAND2_X1 U10790 ( .A1(n9613), .A2(n9434), .ZN(n9436) );
  NAND2_X1 U10791 ( .A1(n9588), .A2(n5047), .ZN(n9440) );
  NOR2_X1 U10792 ( .A1(n9717), .A2(n9443), .ZN(n9445) );
  NOR2_X1 U10793 ( .A1(n9556), .A2(n9447), .ZN(n9446) );
  NAND2_X1 U10794 ( .A1(n9556), .A2(n9447), .ZN(n9448) );
  NAND2_X1 U10795 ( .A1(n9449), .A2(n9448), .ZN(n9532) );
  INV_X1 U10796 ( .A(n9532), .ZN(n9450) );
  NAND2_X1 U10797 ( .A1(n9707), .A2(n9451), .ZN(n9452) );
  NAND2_X1 U10798 ( .A1(n9519), .A2(n9454), .ZN(n9455) );
  NAND2_X1 U10799 ( .A1(n9490), .A2(n9474), .ZN(n9458) );
  XNOR2_X1 U10800 ( .A(n9459), .B(n9470), .ZN(n9686) );
  INV_X1 U10801 ( .A(n9686), .ZN(n9483) );
  NOR2_X1 U10802 ( .A1(n9580), .A2(n9462), .ZN(n9584) );
  NAND2_X1 U10803 ( .A1(n9492), .A2(n9493), .ZN(n9491) );
  NAND2_X1 U10804 ( .A1(n9491), .A2(n9469), .ZN(n9471) );
  AOI211_X1 U10805 ( .C1(n9689), .C2(n9486), .A(n10012), .B(n9476), .ZN(n9688)
         );
  NAND2_X1 U10806 ( .A1(n9688), .A2(n10097), .ZN(n9481) );
  NOR3_X1 U10807 ( .A1(n9478), .A2(n10090), .A3(n9477), .ZN(n9479) );
  AOI21_X1 U10808 ( .B1(n10100), .B2(P1_REG2_REG_29__SCAN_IN), .A(n9479), .ZN(
        n9480) );
  OAI211_X1 U10809 ( .C1(n4591), .C2(n9621), .A(n9481), .B(n9480), .ZN(n9482)
         );
  XNOR2_X1 U10810 ( .A(n9485), .B(n9484), .ZN(n9695) );
  INV_X1 U10811 ( .A(n9503), .ZN(n9488) );
  INV_X1 U10812 ( .A(n9486), .ZN(n9487) );
  AOI211_X1 U10813 ( .C1(n9692), .C2(n9488), .A(n10012), .B(n9487), .ZN(n9691)
         );
  OAI22_X1 U10814 ( .A1(n9490), .A2(n9621), .B1(n9489), .B2(n10058), .ZN(n9500) );
  OAI21_X1 U10815 ( .B1(n9493), .B2(n9492), .A(n9491), .ZN(n9496) );
  INV_X1 U10816 ( .A(n9494), .ZN(n9495) );
  INV_X1 U10817 ( .A(n10090), .ZN(n10079) );
  NAND2_X1 U10818 ( .A1(n9497), .A2(n10079), .ZN(n9498) );
  AOI21_X1 U10819 ( .B1(n9694), .B2(n9498), .A(n10100), .ZN(n9499) );
  OAI21_X1 U10820 ( .B1(n9695), .B2(n9630), .A(n9501), .ZN(P1_U3265) );
  XOR2_X1 U10821 ( .A(n9508), .B(n9502), .Z(n9700) );
  AOI211_X1 U10822 ( .C1(n9697), .C2(n9516), .A(n10012), .B(n9503), .ZN(n9696)
         );
  INV_X1 U10823 ( .A(n9504), .ZN(n9505) );
  AOI22_X1 U10824 ( .A1(n9505), .A2(n10079), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10100), .ZN(n9506) );
  OAI21_X1 U10825 ( .B1(n9507), .B2(n9621), .A(n9506), .ZN(n9513) );
  XNOR2_X1 U10826 ( .A(n9509), .B(n9508), .ZN(n9511) );
  AOI21_X1 U10827 ( .B1(n9511), .B2(n10112), .A(n9510), .ZN(n9699) );
  NOR2_X1 U10828 ( .A1(n9699), .A2(n10100), .ZN(n9512) );
  AOI211_X1 U10829 ( .C1(n10097), .C2(n9696), .A(n9513), .B(n9512), .ZN(n9514)
         );
  OAI21_X1 U10830 ( .B1(n9700), .B2(n9630), .A(n9514), .ZN(P1_U3266) );
  XNOR2_X1 U10831 ( .A(n9515), .B(n9526), .ZN(n9705) );
  INV_X1 U10832 ( .A(n9533), .ZN(n9518) );
  INV_X1 U10833 ( .A(n9516), .ZN(n9517) );
  AOI211_X1 U10834 ( .C1(n9703), .C2(n9518), .A(n10012), .B(n9517), .ZN(n9702)
         );
  NOR2_X1 U10835 ( .A1(n9519), .A2(n9621), .ZN(n9523) );
  OAI22_X1 U10836 ( .A1(n9521), .A2(n10090), .B1(n9520), .B2(n10058), .ZN(
        n9522) );
  AOI211_X1 U10837 ( .C1(n9702), .C2(n10097), .A(n9523), .B(n9522), .ZN(n9531)
         );
  AOI21_X1 U10838 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9529) );
  INV_X1 U10839 ( .A(n9527), .ZN(n9528) );
  OAI21_X1 U10840 ( .B1(n9529), .B2(n10072), .A(n9528), .ZN(n9701) );
  NAND2_X1 U10841 ( .A1(n9701), .A2(n10058), .ZN(n9530) );
  OAI211_X1 U10842 ( .C1(n9705), .C2(n9630), .A(n9531), .B(n9530), .ZN(
        P1_U3267) );
  XOR2_X1 U10843 ( .A(n9532), .B(n9538), .Z(n9710) );
  AOI211_X1 U10844 ( .C1(n9707), .C2(n9550), .A(n10012), .B(n9533), .ZN(n9706)
         );
  AOI22_X1 U10845 ( .A1(n9534), .A2(n10079), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10100), .ZN(n9535) );
  OAI21_X1 U10846 ( .B1(n9536), .B2(n9621), .A(n9535), .ZN(n9542) );
  XOR2_X1 U10847 ( .A(n9538), .B(n9537), .Z(n9540) );
  AOI21_X1 U10848 ( .B1(n9540), .B2(n10112), .A(n9539), .ZN(n9709) );
  NOR2_X1 U10849 ( .A1(n9709), .A2(n10100), .ZN(n9541) );
  AOI211_X1 U10850 ( .C1(n9706), .C2(n10097), .A(n9542), .B(n9541), .ZN(n9543)
         );
  OAI21_X1 U10851 ( .B1(n9710), .B2(n9630), .A(n9543), .ZN(P1_U3268) );
  XNOR2_X1 U10852 ( .A(n9545), .B(n9544), .ZN(n9715) );
  OAI21_X1 U10853 ( .B1(n4477), .B2(n9546), .A(n10112), .ZN(n9549) );
  OAI21_X1 U10854 ( .B1(n9549), .B2(n9548), .A(n9547), .ZN(n9711) );
  INV_X1 U10855 ( .A(n9560), .ZN(n9552) );
  INV_X1 U10856 ( .A(n9550), .ZN(n9551) );
  AOI211_X1 U10857 ( .C1(n9713), .C2(n9552), .A(n10012), .B(n9551), .ZN(n9712)
         );
  NAND2_X1 U10858 ( .A1(n9712), .A2(n10097), .ZN(n9555) );
  AOI22_X1 U10859 ( .A1(n9553), .A2(n10079), .B1(n10100), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9554) );
  OAI211_X1 U10860 ( .C1(n9556), .C2(n9621), .A(n9555), .B(n9554), .ZN(n9557)
         );
  AOI21_X1 U10861 ( .B1(n9711), .B2(n10058), .A(n9557), .ZN(n9558) );
  OAI21_X1 U10862 ( .B1(n9715), .B2(n9630), .A(n9558), .ZN(P1_U3269) );
  XNOR2_X1 U10863 ( .A(n9559), .B(n9566), .ZN(n9720) );
  AOI211_X1 U10864 ( .C1(n9717), .C2(n9573), .A(n10012), .B(n9560), .ZN(n9716)
         );
  INV_X1 U10865 ( .A(n9561), .ZN(n9562) );
  AOI22_X1 U10866 ( .A1(n9562), .A2(n10079), .B1(n10100), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9563) );
  OAI21_X1 U10867 ( .B1(n4581), .B2(n9621), .A(n9563), .ZN(n9570) );
  OAI21_X1 U10868 ( .B1(n9566), .B2(n9565), .A(n9564), .ZN(n9568) );
  AOI21_X1 U10869 ( .B1(n9568), .B2(n10112), .A(n9567), .ZN(n9719) );
  NOR2_X1 U10870 ( .A1(n9719), .A2(n10100), .ZN(n9569) );
  AOI211_X1 U10871 ( .C1(n9716), .C2(n10097), .A(n9570), .B(n9569), .ZN(n9571)
         );
  OAI21_X1 U10872 ( .B1(n9720), .B2(n9630), .A(n9571), .ZN(P1_U3270) );
  XNOR2_X1 U10873 ( .A(n9572), .B(n9581), .ZN(n9725) );
  INV_X1 U10874 ( .A(n9573), .ZN(n9574) );
  AOI211_X1 U10875 ( .C1(n9723), .C2(n4585), .A(n10012), .B(n9574), .ZN(n9722)
         );
  NOR2_X1 U10876 ( .A1(n9575), .A2(n9621), .ZN(n9579) );
  OAI22_X1 U10877 ( .A1(n10058), .A2(n9577), .B1(n9576), .B2(n10090), .ZN(
        n9578) );
  AOI211_X1 U10878 ( .C1(n9722), .C2(n10097), .A(n9579), .B(n9578), .ZN(n9587)
         );
  INV_X1 U10879 ( .A(n9580), .ZN(n9582) );
  OAI21_X1 U10880 ( .B1(n9582), .B2(n9581), .A(n10112), .ZN(n9585) );
  OAI21_X1 U10881 ( .B1(n9585), .B2(n9584), .A(n9583), .ZN(n9721) );
  NAND2_X1 U10882 ( .A1(n9721), .A2(n10058), .ZN(n9586) );
  OAI211_X1 U10883 ( .C1(n9725), .C2(n9630), .A(n9587), .B(n9586), .ZN(
        P1_U3271) );
  XNOR2_X1 U10884 ( .A(n9588), .B(n9591), .ZN(n9730) );
  INV_X1 U10885 ( .A(n9601), .ZN(n9603) );
  AOI21_X1 U10886 ( .B1(n9604), .B2(n9603), .A(n9589), .ZN(n9590) );
  XOR2_X1 U10887 ( .A(n9591), .B(n9590), .Z(n9593) );
  OAI21_X1 U10888 ( .B1(n9593), .B2(n10072), .A(n9592), .ZN(n9726) );
  AOI211_X1 U10889 ( .C1(n9728), .C2(n9607), .A(n10012), .B(n9594), .ZN(n9727)
         );
  NAND2_X1 U10890 ( .A1(n9727), .A2(n10097), .ZN(n9597) );
  AOI22_X1 U10891 ( .A1(n10100), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9595), 
        .B2(n10079), .ZN(n9596) );
  OAI211_X1 U10892 ( .C1(n9598), .C2(n9621), .A(n9597), .B(n9596), .ZN(n9599)
         );
  AOI21_X1 U10893 ( .B1(n9726), .B2(n10058), .A(n9599), .ZN(n9600) );
  OAI21_X1 U10894 ( .B1(n9730), .B2(n9630), .A(n9600), .ZN(P1_U3272) );
  XNOR2_X1 U10895 ( .A(n9602), .B(n9601), .ZN(n9735) );
  XNOR2_X1 U10896 ( .A(n9604), .B(n9603), .ZN(n9606) );
  OAI21_X1 U10897 ( .B1(n9606), .B2(n10072), .A(n9605), .ZN(n9731) );
  INV_X1 U10898 ( .A(n9617), .ZN(n9609) );
  INV_X1 U10899 ( .A(n9607), .ZN(n9608) );
  AOI211_X1 U10900 ( .C1(n9733), .C2(n9609), .A(n10012), .B(n9608), .ZN(n9732)
         );
  NAND2_X1 U10901 ( .A1(n9732), .A2(n10097), .ZN(n9612) );
  AOI22_X1 U10902 ( .A1(n10100), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9610), 
        .B2(n10079), .ZN(n9611) );
  OAI211_X1 U10903 ( .C1(n9613), .C2(n9621), .A(n9612), .B(n9611), .ZN(n9614)
         );
  AOI21_X1 U10904 ( .B1(n10058), .B2(n9731), .A(n9614), .ZN(n9615) );
  OAI21_X1 U10905 ( .B1(n9735), .B2(n9630), .A(n9615), .ZN(P1_U3273) );
  XNOR2_X1 U10906 ( .A(n9616), .B(n9623), .ZN(n9740) );
  AOI211_X1 U10907 ( .C1(n9737), .C2(n9638), .A(n10012), .B(n9617), .ZN(n9736)
         );
  INV_X1 U10908 ( .A(n9618), .ZN(n9619) );
  AOI22_X1 U10909 ( .A1(n10100), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9619), 
        .B2(n10079), .ZN(n9620) );
  OAI21_X1 U10910 ( .B1(n9622), .B2(n9621), .A(n9620), .ZN(n9628) );
  XNOR2_X1 U10911 ( .A(n9624), .B(n9623), .ZN(n9626) );
  AOI21_X1 U10912 ( .B1(n9626), .B2(n10112), .A(n9625), .ZN(n9739) );
  NOR2_X1 U10913 ( .A1(n9739), .A2(n10100), .ZN(n9627) );
  AOI211_X1 U10914 ( .C1(n9736), .C2(n10097), .A(n9628), .B(n9627), .ZN(n9629)
         );
  OAI21_X1 U10915 ( .B1(n9740), .B2(n9630), .A(n9629), .ZN(P1_U3274) );
  XNOR2_X1 U10916 ( .A(n9631), .B(n9635), .ZN(n9633) );
  AOI21_X1 U10917 ( .B1(n9633), .B2(n10112), .A(n9632), .ZN(n9850) );
  XOR2_X1 U10918 ( .A(n9635), .B(n9634), .Z(n9853) );
  NAND2_X1 U10919 ( .A1(n9853), .A2(n10066), .ZN(n9643) );
  OAI22_X1 U10920 ( .A1(n10058), .A2(n9637), .B1(n9636), .B2(n10090), .ZN(
        n9640) );
  OAI211_X1 U10921 ( .C1(n9829), .C2(n9851), .A(n9638), .B(n10081), .ZN(n9849)
         );
  NOR2_X1 U10922 ( .A1(n9849), .A2(n9671), .ZN(n9639) );
  AOI211_X1 U10923 ( .C1(n10077), .C2(n9641), .A(n9640), .B(n9639), .ZN(n9642)
         );
  OAI211_X1 U10924 ( .C1(n10100), .C2(n9850), .A(n9643), .B(n9642), .ZN(
        P1_U3275) );
  OAI21_X1 U10925 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9648) );
  AOI21_X1 U10926 ( .B1(n9648), .B2(n10112), .A(n9647), .ZN(n9861) );
  NOR2_X1 U10927 ( .A1(n9650), .A2(n9649), .ZN(n9859) );
  INV_X1 U10928 ( .A(n9859), .ZN(n9651) );
  NAND3_X1 U10929 ( .A1(n9651), .A2(n10066), .A3(n9864), .ZN(n9658) );
  OAI22_X1 U10930 ( .A1(n10058), .A2(n9653), .B1(n9652), .B2(n10090), .ZN(
        n9655) );
  OAI211_X1 U10931 ( .C1(n9843), .C2(n9862), .A(n9828), .B(n10081), .ZN(n9860)
         );
  NOR2_X1 U10932 ( .A1(n9860), .A2(n9671), .ZN(n9654) );
  AOI211_X1 U10933 ( .C1(n10077), .C2(n4578), .A(n9655), .B(n9654), .ZN(n9657)
         );
  OAI211_X1 U10934 ( .C1(n10100), .C2(n9861), .A(n9658), .B(n9657), .ZN(
        P1_U3277) );
  XOR2_X1 U10935 ( .A(n9659), .B(n9662), .Z(n10192) );
  INV_X1 U10936 ( .A(n9660), .ZN(n9661) );
  NAND2_X1 U10937 ( .A1(n10058), .A2(n9661), .ZN(n10001) );
  INV_X1 U10938 ( .A(n9976), .ZN(n9664) );
  OAI21_X1 U10939 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9666) );
  NAND3_X1 U10940 ( .A1(n9666), .A2(n9665), .A3(n10112), .ZN(n9667) );
  OAI211_X1 U10941 ( .C1(n10192), .C2(n9992), .A(n9668), .B(n9667), .ZN(n10196) );
  NAND2_X1 U10942 ( .A1(n10196), .A2(n10058), .ZN(n9676) );
  OAI22_X1 U10943 ( .A1(n10058), .A2(n9670), .B1(n9669), .B2(n10090), .ZN(
        n9673) );
  OAI211_X1 U10944 ( .C1(n9986), .C2(n10195), .A(n9842), .B(n10081), .ZN(
        n10193) );
  NOR2_X1 U10945 ( .A1(n10193), .A2(n9671), .ZN(n9672) );
  AOI211_X1 U10946 ( .C1(n10077), .C2(n9674), .A(n9673), .B(n9672), .ZN(n9675)
         );
  OAI211_X1 U10947 ( .C1(n10192), .C2(n10001), .A(n9676), .B(n9675), .ZN(
        P1_U3279) );
  OAI211_X1 U10948 ( .C1(n9678), .C2(n10194), .A(n9677), .B(n9682), .ZN(n9744)
         );
  NOR2_X1 U10949 ( .A1(n9680), .A2(n9679), .ZN(n9743) );
  MUX2_X1 U10950 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9744), .S(n10221), .Z(
        P1_U3553) );
  OAI211_X1 U10951 ( .C1(n9684), .C2(n10194), .A(n9683), .B(n9682), .ZN(n9745)
         );
  MUX2_X1 U10952 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9745), .S(n10221), .Z(
        P1_U3552) );
  NAND2_X1 U10953 ( .A1(n4555), .A2(n9685), .ZN(n10116) );
  NAND2_X1 U10954 ( .A1(n9686), .A2(n10190), .ZN(n9690) );
  MUX2_X1 U10955 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9746), .S(n10221), .Z(
        P1_U3551) );
  AOI21_X1 U10956 ( .B1(n10148), .B2(n9692), .A(n9691), .ZN(n9693) );
  OAI211_X1 U10957 ( .C1(n9695), .C2(n10150), .A(n9694), .B(n9693), .ZN(n9747)
         );
  MUX2_X1 U10958 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9747), .S(n10221), .Z(
        P1_U3550) );
  AOI21_X1 U10959 ( .B1(n10148), .B2(n9697), .A(n9696), .ZN(n9698) );
  OAI211_X1 U10960 ( .C1(n9700), .C2(n10150), .A(n9699), .B(n9698), .ZN(n9748)
         );
  MUX2_X1 U10961 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9748), .S(n10221), .Z(
        P1_U3549) );
  AOI211_X1 U10962 ( .C1(n10148), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9704)
         );
  OAI21_X1 U10963 ( .B1(n9705), .B2(n10150), .A(n9704), .ZN(n9749) );
  MUX2_X1 U10964 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9749), .S(n10221), .Z(
        P1_U3548) );
  AOI21_X1 U10965 ( .B1(n10148), .B2(n9707), .A(n9706), .ZN(n9708) );
  OAI211_X1 U10966 ( .C1(n9710), .C2(n10150), .A(n9709), .B(n9708), .ZN(n9750)
         );
  MUX2_X1 U10967 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9750), .S(n10221), .Z(
        P1_U3547) );
  AOI211_X1 U10968 ( .C1(n10148), .C2(n9713), .A(n9712), .B(n9711), .ZN(n9714)
         );
  OAI21_X1 U10969 ( .B1(n9715), .B2(n10150), .A(n9714), .ZN(n9751) );
  MUX2_X1 U10970 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9751), .S(n10221), .Z(
        P1_U3546) );
  AOI21_X1 U10971 ( .B1(n10148), .B2(n9717), .A(n9716), .ZN(n9718) );
  OAI211_X1 U10972 ( .C1(n9720), .C2(n10150), .A(n9719), .B(n9718), .ZN(n9752)
         );
  MUX2_X1 U10973 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9752), .S(n10221), .Z(
        P1_U3545) );
  AOI211_X1 U10974 ( .C1(n10148), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9724)
         );
  OAI21_X1 U10975 ( .B1(n9725), .B2(n10150), .A(n9724), .ZN(n9753) );
  MUX2_X1 U10976 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9753), .S(n10221), .Z(
        P1_U3544) );
  AOI211_X1 U10977 ( .C1(n10148), .C2(n9728), .A(n9727), .B(n9726), .ZN(n9729)
         );
  OAI21_X1 U10978 ( .B1(n9730), .B2(n10150), .A(n9729), .ZN(n9754) );
  MUX2_X1 U10979 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9754), .S(n10221), .Z(
        P1_U3543) );
  AOI211_X1 U10980 ( .C1(n10148), .C2(n9733), .A(n9732), .B(n9731), .ZN(n9734)
         );
  OAI21_X1 U10981 ( .B1(n9735), .B2(n10150), .A(n9734), .ZN(n9755) );
  MUX2_X1 U10982 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9755), .S(n10221), .Z(
        P1_U3542) );
  AOI21_X1 U10983 ( .B1(n10148), .B2(n9737), .A(n9736), .ZN(n9738) );
  OAI211_X1 U10984 ( .C1(n9740), .C2(n10150), .A(n9739), .B(n9738), .ZN(n9756)
         );
  MUX2_X1 U10985 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9756), .S(n10221), .Z(
        P1_U3541) );
  MUX2_X1 U10986 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9744), .S(n10201), .Z(
        P1_U3521) );
  MUX2_X1 U10987 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9745), .S(n10201), .Z(
        P1_U3520) );
  MUX2_X1 U10988 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9746), .S(n10201), .Z(
        P1_U3519) );
  MUX2_X1 U10989 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9747), .S(n10201), .Z(
        P1_U3518) );
  MUX2_X1 U10990 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9748), .S(n10201), .Z(
        P1_U3517) );
  MUX2_X1 U10991 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9749), .S(n10201), .Z(
        P1_U3516) );
  MUX2_X1 U10992 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9750), .S(n10201), .Z(
        P1_U3515) );
  MUX2_X1 U10993 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9751), .S(n10201), .Z(
        P1_U3514) );
  MUX2_X1 U10994 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9752), .S(n10201), .Z(
        P1_U3513) );
  MUX2_X1 U10995 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9753), .S(n10201), .Z(
        P1_U3512) );
  MUX2_X1 U10996 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9754), .S(n10201), .Z(
        P1_U3511) );
  MUX2_X1 U10997 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9755), .S(n10201), .Z(
        P1_U3510) );
  MUX2_X1 U10998 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9756), .S(n10201), .Z(
        P1_U3509) );
  NAND2_X1 U10999 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .ZN(n9758) );
  OAI22_X1 U11000 ( .A1(n9759), .A2(n9758), .B1(n9757), .B2(n9769), .ZN(n9760)
         );
  INV_X1 U11001 ( .A(n9760), .ZN(n9761) );
  OAI21_X1 U11002 ( .B1(n9762), .B2(n9773), .A(n9761), .ZN(P1_U3324) );
  OAI222_X1 U11003 ( .A1(n9769), .A2(n9765), .B1(n9773), .B2(n9764), .C1(n9763), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U11004 ( .A1(n9769), .A2(n9768), .B1(P1_U3086), .B2(n9767), .C1(
        n9773), .C2(n9766), .ZN(P1_U3326) );
  INV_X1 U11005 ( .A(n9770), .ZN(n9772) );
  OAI222_X1 U11006 ( .A1(n9774), .A2(P1_U3086), .B1(n9773), .B2(n9772), .C1(
        n9771), .C2(n9769), .ZN(P1_U3327) );
  OAI222_X1 U11007 ( .A1(n9769), .A2(n9778), .B1(n9777), .B2(n9776), .C1(n9775), .C2(P1_U3086), .ZN(P1_U3329) );
  MUX2_X1 U11008 ( .A(n9780), .B(n9779), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11009 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9792) );
  AOI211_X1 U11010 ( .C1(n9783), .C2(n9782), .A(n9781), .B(n9958), .ZN(n9788)
         );
  AOI211_X1 U11011 ( .C1(n9786), .C2(n9785), .A(n9784), .B(n9930), .ZN(n9787)
         );
  AOI211_X1 U11012 ( .C1(n9969), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9791)
         );
  NAND2_X1 U11013 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9790) );
  OAI211_X1 U11014 ( .C1(n9972), .C2(n9792), .A(n9791), .B(n9790), .ZN(
        P1_U3253) );
  INV_X1 U11015 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9805) );
  INV_X1 U11016 ( .A(n9793), .ZN(n9796) );
  AOI211_X1 U11017 ( .C1(n9796), .C2(n9795), .A(n9794), .B(n9930), .ZN(n9801)
         );
  AOI211_X1 U11018 ( .C1(n9799), .C2(n9798), .A(n9958), .B(n9797), .ZN(n9800)
         );
  AOI211_X1 U11019 ( .C1(n9969), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9804)
         );
  NAND2_X1 U11020 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9803) );
  OAI211_X1 U11021 ( .C1(n9972), .C2(n9805), .A(n9804), .B(n9803), .ZN(
        P1_U3250) );
  INV_X1 U11022 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9817) );
  AOI211_X1 U11023 ( .C1(n9808), .C2(n9807), .A(n9806), .B(n9930), .ZN(n9813)
         );
  AOI211_X1 U11024 ( .C1(n9811), .C2(n9810), .A(n9809), .B(n9958), .ZN(n9812)
         );
  AOI211_X1 U11025 ( .C1(n9969), .C2(n9814), .A(n9813), .B(n9812), .ZN(n9816)
         );
  OAI211_X1 U11026 ( .C1(n9972), .C2(n9817), .A(n9816), .B(n9815), .ZN(
        P1_U3251) );
  AOI21_X1 U11027 ( .B1(n9819), .B2(n9818), .A(n10072), .ZN(n9822) );
  AOI21_X1 U11028 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9855) );
  INV_X1 U11029 ( .A(n9823), .ZN(n9824) );
  AOI222_X1 U11030 ( .A1(n9825), .A2(n10077), .B1(P1_REG2_REG_17__SCAN_IN), 
        .B2(n10100), .C1(n10079), .C2(n9824), .ZN(n9834) );
  XNOR2_X1 U11031 ( .A(n9827), .B(n9826), .ZN(n9858) );
  INV_X1 U11032 ( .A(n9828), .ZN(n9831) );
  INV_X1 U11033 ( .A(n9829), .ZN(n9830) );
  OAI211_X1 U11034 ( .C1(n9856), .C2(n9831), .A(n9830), .B(n10081), .ZN(n9854)
         );
  INV_X1 U11035 ( .A(n9854), .ZN(n9832) );
  AOI22_X1 U11036 ( .A1(n9858), .A2(n10066), .B1(n10097), .B2(n9832), .ZN(
        n9833) );
  OAI211_X1 U11037 ( .C1(n10100), .C2(n9855), .A(n9834), .B(n9833), .ZN(
        P1_U3276) );
  XNOR2_X1 U11038 ( .A(n9835), .B(n9841), .ZN(n9837) );
  AOI21_X1 U11039 ( .B1(n9837), .B2(n10112), .A(n9836), .ZN(n9867) );
  INV_X1 U11040 ( .A(n9838), .ZN(n9839) );
  AOI222_X1 U11041 ( .A1(n4438), .A2(n10077), .B1(P1_REG2_REG_15__SCAN_IN), 
        .B2(n10100), .C1(n9839), .C2(n10079), .ZN(n9848) );
  XOR2_X1 U11042 ( .A(n9841), .B(n9840), .Z(n9870) );
  INV_X1 U11043 ( .A(n9842), .ZN(n9845) );
  INV_X1 U11044 ( .A(n9843), .ZN(n9844) );
  OAI211_X1 U11045 ( .C1(n9868), .C2(n9845), .A(n9844), .B(n10081), .ZN(n9866)
         );
  INV_X1 U11046 ( .A(n9866), .ZN(n9846) );
  AOI22_X1 U11047 ( .A1(n9870), .A2(n10066), .B1(n10097), .B2(n9846), .ZN(
        n9847) );
  OAI211_X1 U11048 ( .C1(n10100), .C2(n9867), .A(n9848), .B(n9847), .ZN(
        P1_U3278) );
  OAI211_X1 U11049 ( .C1(n9851), .C2(n10194), .A(n9850), .B(n9849), .ZN(n9852)
         );
  AOI21_X1 U11050 ( .B1(n9853), .B2(n10190), .A(n9852), .ZN(n9871) );
  AOI22_X1 U11051 ( .A1(n10221), .A2(n9871), .B1(n9385), .B2(n10219), .ZN(
        P1_U3540) );
  OAI211_X1 U11052 ( .C1(n9856), .C2(n10194), .A(n9855), .B(n9854), .ZN(n9857)
         );
  AOI21_X1 U11053 ( .B1(n9858), .B2(n10190), .A(n9857), .ZN(n9872) );
  AOI22_X1 U11054 ( .A1(n10221), .A2(n9872), .B1(n7317), .B2(n10219), .ZN(
        P1_U3539) );
  NOR2_X1 U11055 ( .A1(n9859), .A2(n10150), .ZN(n9865) );
  OAI211_X1 U11056 ( .C1(n9862), .C2(n10194), .A(n9861), .B(n9860), .ZN(n9863)
         );
  AOI21_X1 U11057 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n9873) );
  AOI22_X1 U11058 ( .A1(n10221), .A2(n9873), .B1(n7306), .B2(n10219), .ZN(
        P1_U3538) );
  OAI211_X1 U11059 ( .C1(n9868), .C2(n10194), .A(n9867), .B(n9866), .ZN(n9869)
         );
  AOI21_X1 U11060 ( .B1(n9870), .B2(n10190), .A(n9869), .ZN(n9874) );
  AOI22_X1 U11061 ( .A1(n10221), .A2(n9874), .B1(n7298), .B2(n10219), .ZN(
        P1_U3537) );
  AOI22_X1 U11062 ( .A1(n10201), .A2(n9871), .B1(n7332), .B2(n10200), .ZN(
        P1_U3507) );
  AOI22_X1 U11063 ( .A1(n10201), .A2(n9872), .B1(n7320), .B2(n10200), .ZN(
        P1_U3504) );
  AOI22_X1 U11064 ( .A1(n10201), .A2(n9873), .B1(n7310), .B2(n10200), .ZN(
        P1_U3501) );
  AOI22_X1 U11065 ( .A1(n10201), .A2(n9874), .B1(n7297), .B2(n10200), .ZN(
        P1_U3498) );
  XNOR2_X1 U11066 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  NOR2_X1 U11067 ( .A1(n9875), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9877) );
  OR2_X1 U11068 ( .A1(n9876), .A2(n9877), .ZN(n9880) );
  INV_X1 U11069 ( .A(n9877), .ZN(n9879) );
  MUX2_X1 U11070 ( .A(n9880), .B(n9879), .S(n9878), .Z(n9882) );
  NAND2_X1 U11071 ( .A1(n9882), .A2(n9881), .ZN(n9886) );
  AOI22_X1 U11072 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9883), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9884) );
  OAI21_X1 U11073 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(P1_U3243) );
  INV_X1 U11074 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9898) );
  AOI211_X1 U11075 ( .C1(n9889), .C2(n9888), .A(n9887), .B(n9930), .ZN(n9894)
         );
  AOI211_X1 U11076 ( .C1(n9892), .C2(n9891), .A(n9890), .B(n9958), .ZN(n9893)
         );
  AOI211_X1 U11077 ( .C1(n9969), .C2(n9895), .A(n9894), .B(n9893), .ZN(n9897)
         );
  NAND2_X1 U11078 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9896) );
  OAI211_X1 U11079 ( .C1(n9972), .C2(n9898), .A(n9897), .B(n9896), .ZN(
        P1_U3254) );
  INV_X1 U11080 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9910) );
  AOI211_X1 U11081 ( .C1(n9901), .C2(n9900), .A(n9899), .B(n9958), .ZN(n9906)
         );
  AOI211_X1 U11082 ( .C1(n9904), .C2(n9903), .A(n9902), .B(n9930), .ZN(n9905)
         );
  AOI211_X1 U11083 ( .C1(n9969), .C2(n9907), .A(n9906), .B(n9905), .ZN(n9909)
         );
  NAND2_X1 U11084 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9908) );
  OAI211_X1 U11085 ( .C1(n9972), .C2(n9910), .A(n9909), .B(n9908), .ZN(
        P1_U3256) );
  INV_X1 U11086 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9926) );
  INV_X1 U11087 ( .A(n9911), .ZN(n9922) );
  AOI21_X1 U11088 ( .B1(n9914), .B2(n9913), .A(n9912), .ZN(n9915) );
  NAND2_X1 U11089 ( .A1(n9948), .A2(n9915), .ZN(n9921) );
  AOI21_X1 U11090 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n9919) );
  NAND2_X1 U11091 ( .A1(n9961), .A2(n9919), .ZN(n9920) );
  OAI211_X1 U11092 ( .C1(n9952), .C2(n9922), .A(n9921), .B(n9920), .ZN(n9923)
         );
  INV_X1 U11093 ( .A(n9923), .ZN(n9925) );
  NAND2_X1 U11094 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9924) );
  OAI211_X1 U11095 ( .C1(n9972), .C2(n9926), .A(n9925), .B(n9924), .ZN(
        P1_U3257) );
  INV_X1 U11096 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9938) );
  INV_X1 U11097 ( .A(n9927), .ZN(n9929) );
  AOI211_X1 U11098 ( .C1(n7298), .C2(n9929), .A(n9928), .B(n9958), .ZN(n9934)
         );
  AOI211_X1 U11099 ( .C1(n7295), .C2(n9932), .A(n9931), .B(n9930), .ZN(n9933)
         );
  AOI211_X1 U11100 ( .C1(n9969), .C2(n9935), .A(n9934), .B(n9933), .ZN(n9937)
         );
  NAND2_X1 U11101 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9936) );
  OAI211_X1 U11102 ( .C1(n9972), .C2(n9938), .A(n9937), .B(n9936), .ZN(
        P1_U3258) );
  INV_X1 U11103 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9956) );
  INV_X1 U11104 ( .A(n9939), .ZN(n9951) );
  AOI21_X1 U11105 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(n9943) );
  NAND2_X1 U11106 ( .A1(n9961), .A2(n9943), .ZN(n9950) );
  OAI21_X1 U11107 ( .B1(n9946), .B2(n9945), .A(n9944), .ZN(n9947) );
  NAND2_X1 U11108 ( .A1(n9948), .A2(n9947), .ZN(n9949) );
  OAI211_X1 U11109 ( .C1(n9952), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9953)
         );
  INV_X1 U11110 ( .A(n9953), .ZN(n9955) );
  NAND2_X1 U11111 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n9954) );
  OAI211_X1 U11112 ( .C1(n9956), .C2(n9972), .A(n9955), .B(n9954), .ZN(
        P1_U3259) );
  AOI211_X1 U11113 ( .C1(n9960), .C2(n9959), .A(n9958), .B(n9957), .ZN(n9967)
         );
  OAI211_X1 U11114 ( .C1(n9964), .C2(n9963), .A(n9962), .B(n9961), .ZN(n9965)
         );
  INV_X1 U11115 ( .A(n9965), .ZN(n9966) );
  AOI211_X1 U11116 ( .C1(n9969), .C2(n9968), .A(n9967), .B(n9966), .ZN(n9971)
         );
  NAND2_X1 U11117 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9970) );
  OAI211_X1 U11118 ( .C1(n9972), .C2(n10295), .A(n9971), .B(n9970), .ZN(
        P1_U3261) );
  OAI21_X1 U11119 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(n9977) );
  AOI21_X1 U11120 ( .B1(n9977), .B2(n9976), .A(n10072), .ZN(n9979) );
  NOR2_X1 U11121 ( .A1(n9979), .A2(n9978), .ZN(n10187) );
  INV_X1 U11122 ( .A(n9980), .ZN(n9981) );
  AOI222_X1 U11123 ( .A1(n9984), .A2(n10077), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n10100), .C1(n9981), .C2(n10079), .ZN(n9990) );
  XNOR2_X1 U11124 ( .A(n9983), .B(n9982), .ZN(n10191) );
  INV_X1 U11125 ( .A(n9984), .ZN(n10188) );
  INV_X1 U11126 ( .A(n9985), .ZN(n9987) );
  OAI211_X1 U11127 ( .C1(n10188), .C2(n9987), .A(n4590), .B(n10081), .ZN(
        n10186) );
  INV_X1 U11128 ( .A(n10186), .ZN(n9988) );
  AOI22_X1 U11129 ( .A1(n10191), .A2(n10066), .B1(n10097), .B2(n9988), .ZN(
        n9989) );
  OAI211_X1 U11130 ( .C1(n10100), .C2(n10187), .A(n9990), .B(n9989), .ZN(
        P1_U3280) );
  XNOR2_X1 U11131 ( .A(n9991), .B(n9995), .ZN(n10180) );
  INV_X1 U11132 ( .A(n9992), .ZN(n10076) );
  OAI211_X1 U11133 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n10112), .ZN(n9996)
         );
  INV_X1 U11134 ( .A(n9996), .ZN(n9998) );
  AOI211_X1 U11135 ( .C1(n10180), .C2(n10076), .A(n9998), .B(n9997), .ZN(
        n10177) );
  INV_X1 U11136 ( .A(n9999), .ZN(n10000) );
  AOI222_X1 U11137 ( .A1(n10002), .A2(n10077), .B1(n10000), .B2(n10079), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(n10100), .ZN(n10009) );
  INV_X1 U11138 ( .A(n10001), .ZN(n10084) );
  INV_X1 U11139 ( .A(n10002), .ZN(n10176) );
  INV_X1 U11140 ( .A(n10003), .ZN(n10006) );
  INV_X1 U11141 ( .A(n10004), .ZN(n10005) );
  OAI211_X1 U11142 ( .C1(n10176), .C2(n10006), .A(n10005), .B(n10081), .ZN(
        n10175) );
  INV_X1 U11143 ( .A(n10175), .ZN(n10007) );
  AOI22_X1 U11144 ( .A1(n10180), .A2(n10084), .B1(n10097), .B2(n10007), .ZN(
        n10008) );
  OAI211_X1 U11145 ( .C1(n10100), .C2(n10177), .A(n10009), .B(n10008), .ZN(
        P1_U3282) );
  XNOR2_X1 U11146 ( .A(n10010), .B(n10019), .ZN(n10169) );
  AOI211_X1 U11147 ( .C1(n10024), .C2(n10013), .A(n10012), .B(n10011), .ZN(
        n10015) );
  NOR2_X1 U11148 ( .A1(n10015), .A2(n10014), .ZN(n10165) );
  NAND2_X1 U11149 ( .A1(n10017), .A2(n10016), .ZN(n10018) );
  XOR2_X1 U11150 ( .A(n10019), .B(n10018), .Z(n10020) );
  NAND2_X1 U11151 ( .A1(n10020), .A2(n10112), .ZN(n10166) );
  INV_X1 U11152 ( .A(n10021), .ZN(n10022) );
  AOI22_X1 U11153 ( .A1(n10024), .A2(n10023), .B1(n10022), .B2(n10079), .ZN(
        n10025) );
  OAI211_X1 U11154 ( .C1(n4434), .C2(n10165), .A(n10166), .B(n10025), .ZN(
        n10027) );
  AOI21_X1 U11155 ( .B1(n10169), .B2(n10028), .A(n10027), .ZN(n10029) );
  AOI22_X1 U11156 ( .A1(n10100), .A2(n6855), .B1(n10029), .B2(n10058), .ZN(
        P1_U3284) );
  XNOR2_X1 U11157 ( .A(n10030), .B(n10032), .ZN(n10159) );
  XOR2_X1 U11158 ( .A(n10032), .B(n10031), .Z(n10033) );
  NOR2_X1 U11159 ( .A1(n10033), .A2(n10072), .ZN(n10034) );
  AOI211_X1 U11160 ( .C1(n10159), .C2(n10076), .A(n10035), .B(n10034), .ZN(
        n10156) );
  INV_X1 U11161 ( .A(n10036), .ZN(n10037) );
  AOI222_X1 U11162 ( .A1(n10038), .A2(n10077), .B1(P1_REG2_REG_7__SCAN_IN), 
        .B2(n10100), .C1(n10079), .C2(n10037), .ZN(n10042) );
  OAI211_X1 U11163 ( .C1(n10155), .C2(n4462), .A(n4597), .B(n10081), .ZN(
        n10154) );
  INV_X1 U11164 ( .A(n10154), .ZN(n10040) );
  AOI22_X1 U11165 ( .A1(n10159), .A2(n10084), .B1(n10097), .B2(n10040), .ZN(
        n10041) );
  OAI211_X1 U11166 ( .C1(n10100), .C2(n10156), .A(n10042), .B(n10041), .ZN(
        P1_U3286) );
  XOR2_X1 U11167 ( .A(n10043), .B(n10048), .Z(n10045) );
  AOI21_X1 U11168 ( .B1(n10045), .B2(n10112), .A(n10044), .ZN(n10142) );
  AOI222_X1 U11169 ( .A1(n10047), .A2(n10077), .B1(P1_REG2_REG_5__SCAN_IN), 
        .B2(n10100), .C1(n10079), .C2(n10046), .ZN(n10054) );
  XNOR2_X1 U11170 ( .A(n10049), .B(n10048), .ZN(n10145) );
  OAI211_X1 U11171 ( .C1(n10051), .C2(n10141), .A(n10081), .B(n10050), .ZN(
        n10140) );
  INV_X1 U11172 ( .A(n10140), .ZN(n10052) );
  AOI22_X1 U11173 ( .A1(n10145), .A2(n10066), .B1(n10097), .B2(n10052), .ZN(
        n10053) );
  OAI211_X1 U11174 ( .C1(n10100), .C2(n10142), .A(n10054), .B(n10053), .ZN(
        P1_U3288) );
  XNOR2_X1 U11175 ( .A(n10055), .B(n10061), .ZN(n10057) );
  AOI21_X1 U11176 ( .B1(n10057), .B2(n10112), .A(n10056), .ZN(n10130) );
  OAI22_X1 U11177 ( .A1(n10058), .A2(n8639), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10090), .ZN(n10059) );
  AOI21_X1 U11178 ( .B1(n10077), .B2(n10060), .A(n10059), .ZN(n10068) );
  XNOR2_X1 U11179 ( .A(n10062), .B(n10061), .ZN(n10133) );
  OAI211_X1 U11180 ( .C1(n10129), .C2(n10064), .A(n10063), .B(n10081), .ZN(
        n10128) );
  INV_X1 U11181 ( .A(n10128), .ZN(n10065) );
  AOI22_X1 U11182 ( .A1(n10133), .A2(n10066), .B1(n10097), .B2(n10065), .ZN(
        n10067) );
  OAI211_X1 U11183 ( .C1(n10100), .C2(n10130), .A(n10068), .B(n10067), .ZN(
        P1_U3290) );
  XNOR2_X1 U11184 ( .A(n10069), .B(n10070), .ZN(n10122) );
  XNOR2_X1 U11185 ( .A(n10071), .B(n10070), .ZN(n10073) );
  NOR2_X1 U11186 ( .A1(n10073), .A2(n10072), .ZN(n10074) );
  AOI211_X1 U11187 ( .C1(n10076), .C2(n10122), .A(n10075), .B(n10074), .ZN(
        n10119) );
  AOI222_X1 U11188 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(n10100), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10079), .C1(n4440), .C2(n10077), .ZN(
        n10086) );
  OAI211_X1 U11189 ( .C1(n10118), .C2(n10082), .A(n10081), .B(n10080), .ZN(
        n10117) );
  INV_X1 U11190 ( .A(n10117), .ZN(n10083) );
  AOI22_X1 U11191 ( .A1(n10122), .A2(n10084), .B1(n10097), .B2(n10083), .ZN(
        n10085) );
  OAI211_X1 U11192 ( .C1(n10100), .C2(n10119), .A(n10086), .B(n10085), .ZN(
        P1_U3292) );
  INV_X1 U11193 ( .A(n10087), .ZN(n10095) );
  INV_X1 U11194 ( .A(n10114), .ZN(n10094) );
  NAND2_X1 U11195 ( .A1(n10089), .A2(n10088), .ZN(n10113) );
  OAI22_X1 U11196 ( .A1(n10113), .A2(n10092), .B1(n10091), .B2(n10090), .ZN(
        n10093) );
  AOI211_X1 U11197 ( .C1(n10111), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10099) );
  INV_X1 U11198 ( .A(n10113), .ZN(n10096) );
  AOI22_X1 U11199 ( .A1(n10097), .A2(n10096), .B1(n10100), .B2(
        P1_REG2_REG_0__SCAN_IN), .ZN(n10098) );
  OAI21_X1 U11200 ( .B1(n10100), .B2(n10099), .A(n10098), .ZN(P1_U3293) );
  NOR2_X1 U11201 ( .A1(n10109), .A2(n10101), .ZN(P1_U3294) );
  AND2_X1 U11202 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10110), .ZN(P1_U3295) );
  AND2_X1 U11203 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10110), .ZN(P1_U3296) );
  AND2_X1 U11204 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10110), .ZN(P1_U3297) );
  AND2_X1 U11205 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10110), .ZN(P1_U3298) );
  AND2_X1 U11206 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10110), .ZN(P1_U3299) );
  AND2_X1 U11207 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10110), .ZN(P1_U3300) );
  AND2_X1 U11208 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10110), .ZN(P1_U3301) );
  NOR2_X1 U11209 ( .A1(n10109), .A2(n10102), .ZN(P1_U3302) );
  AND2_X1 U11210 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10110), .ZN(P1_U3303) );
  NOR2_X1 U11211 ( .A1(n10109), .A2(n10103), .ZN(P1_U3304) );
  AND2_X1 U11212 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10110), .ZN(P1_U3305) );
  AND2_X1 U11213 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10110), .ZN(P1_U3306) );
  AND2_X1 U11214 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10110), .ZN(P1_U3307) );
  NOR2_X1 U11215 ( .A1(n10109), .A2(n10104), .ZN(P1_U3308) );
  AND2_X1 U11216 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10110), .ZN(P1_U3309) );
  AND2_X1 U11217 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10110), .ZN(P1_U3310) );
  AND2_X1 U11218 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10110), .ZN(P1_U3311) );
  AND2_X1 U11219 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10110), .ZN(P1_U3312) );
  NOR2_X1 U11220 ( .A1(n10109), .A2(n10105), .ZN(P1_U3313) );
  NOR2_X1 U11221 ( .A1(n10109), .A2(n10106), .ZN(P1_U3314) );
  NOR2_X1 U11222 ( .A1(n10109), .A2(n10107), .ZN(P1_U3315) );
  AND2_X1 U11223 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10110), .ZN(P1_U3316) );
  NOR2_X1 U11224 ( .A1(n10109), .A2(n10108), .ZN(P1_U3317) );
  AND2_X1 U11225 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10110), .ZN(P1_U3318) );
  AND2_X1 U11226 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10110), .ZN(P1_U3319) );
  AND2_X1 U11227 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10110), .ZN(P1_U3320) );
  AND2_X1 U11228 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10110), .ZN(P1_U3321) );
  AND2_X1 U11229 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10110), .ZN(P1_U3322) );
  AND2_X1 U11230 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10110), .ZN(P1_U3323) );
  OAI21_X1 U11231 ( .B1(n10190), .B2(n10112), .A(n10111), .ZN(n10115) );
  AND3_X1 U11232 ( .A1(n10115), .A2(n10114), .A3(n10113), .ZN(n10202) );
  AOI22_X1 U11233 ( .A1(n10201), .A2(n10202), .B1(n6127), .B2(n10200), .ZN(
        P1_U3453) );
  INV_X1 U11234 ( .A(n10116), .ZN(n10199) );
  OAI21_X1 U11235 ( .B1(n10118), .B2(n10194), .A(n10117), .ZN(n10121) );
  INV_X1 U11236 ( .A(n10119), .ZN(n10120) );
  AOI211_X1 U11237 ( .C1(n10199), .C2(n10122), .A(n10121), .B(n10120), .ZN(
        n10203) );
  AOI22_X1 U11238 ( .A1(n10201), .A2(n10203), .B1(n6177), .B2(n10200), .ZN(
        P1_U3456) );
  OAI21_X1 U11239 ( .B1(n10124), .B2(n10194), .A(n10123), .ZN(n10126) );
  AOI211_X1 U11240 ( .C1(n10127), .C2(n10190), .A(n10126), .B(n10125), .ZN(
        n10205) );
  AOI22_X1 U11241 ( .A1(n10201), .A2(n10205), .B1(n6280), .B2(n10200), .ZN(
        P1_U3459) );
  OAI21_X1 U11242 ( .B1(n10129), .B2(n10194), .A(n10128), .ZN(n10132) );
  INV_X1 U11243 ( .A(n10130), .ZN(n10131) );
  AOI211_X1 U11244 ( .C1(n10190), .C2(n10133), .A(n10132), .B(n10131), .ZN(
        n10206) );
  AOI22_X1 U11245 ( .A1(n10201), .A2(n10206), .B1(n6317), .B2(n10200), .ZN(
        P1_U3462) );
  AOI21_X1 U11246 ( .B1(n10148), .B2(n10135), .A(n10134), .ZN(n10136) );
  OAI211_X1 U11247 ( .C1(n10138), .C2(n10150), .A(n10137), .B(n10136), .ZN(
        n10139) );
  INV_X1 U11248 ( .A(n10139), .ZN(n10208) );
  AOI22_X1 U11249 ( .A1(n10201), .A2(n10208), .B1(n6430), .B2(n10200), .ZN(
        P1_U3465) );
  OAI21_X1 U11250 ( .B1(n10141), .B2(n10194), .A(n10140), .ZN(n10144) );
  INV_X1 U11251 ( .A(n10142), .ZN(n10143) );
  AOI211_X1 U11252 ( .C1(n10190), .C2(n10145), .A(n10144), .B(n10143), .ZN(
        n10209) );
  AOI22_X1 U11253 ( .A1(n10201), .A2(n10209), .B1(n6485), .B2(n10200), .ZN(
        P1_U3468) );
  AOI21_X1 U11254 ( .B1(n10148), .B2(n10147), .A(n10146), .ZN(n10149) );
  OAI21_X1 U11255 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(n10153) );
  NOR2_X1 U11256 ( .A1(n10153), .A2(n10152), .ZN(n10210) );
  AOI22_X1 U11257 ( .A1(n10201), .A2(n10210), .B1(n6635), .B2(n10200), .ZN(
        P1_U3471) );
  OAI21_X1 U11258 ( .B1(n10155), .B2(n10194), .A(n10154), .ZN(n10158) );
  INV_X1 U11259 ( .A(n10156), .ZN(n10157) );
  AOI211_X1 U11260 ( .C1(n10199), .C2(n10159), .A(n10158), .B(n10157), .ZN(
        n10211) );
  AOI22_X1 U11261 ( .A1(n10201), .A2(n10211), .B1(n6707), .B2(n10200), .ZN(
        P1_U3474) );
  OAI211_X1 U11262 ( .C1(n10162), .C2(n10194), .A(n10161), .B(n10160), .ZN(
        n10163) );
  AOI21_X1 U11263 ( .B1(n10190), .B2(n10164), .A(n10163), .ZN(n10212) );
  AOI22_X1 U11264 ( .A1(n10201), .A2(n10212), .B1(n6063), .B2(n10200), .ZN(
        P1_U3477) );
  OAI211_X1 U11265 ( .C1(n10167), .C2(n10194), .A(n10166), .B(n10165), .ZN(
        n10168) );
  AOI21_X1 U11266 ( .B1(n10169), .B2(n10190), .A(n10168), .ZN(n10213) );
  AOI22_X1 U11267 ( .A1(n10201), .A2(n10213), .B1(n6856), .B2(n10200), .ZN(
        P1_U3480) );
  OAI211_X1 U11268 ( .C1(n10172), .C2(n10194), .A(n10171), .B(n10170), .ZN(
        n10173) );
  AOI21_X1 U11269 ( .B1(n10174), .B2(n10190), .A(n10173), .ZN(n10214) );
  AOI22_X1 U11270 ( .A1(n10201), .A2(n10214), .B1(n6873), .B2(n10200), .ZN(
        P1_U3483) );
  OAI21_X1 U11271 ( .B1(n10176), .B2(n10194), .A(n10175), .ZN(n10179) );
  INV_X1 U11272 ( .A(n10177), .ZN(n10178) );
  AOI211_X1 U11273 ( .C1(n10199), .C2(n10180), .A(n10179), .B(n10178), .ZN(
        n10215) );
  AOI22_X1 U11274 ( .A1(n10201), .A2(n10215), .B1(n6071), .B2(n10200), .ZN(
        P1_U3486) );
  OAI211_X1 U11275 ( .C1(n10183), .C2(n10194), .A(n10182), .B(n10181), .ZN(
        n10184) );
  AOI21_X1 U11276 ( .B1(n10185), .B2(n10190), .A(n10184), .ZN(n10217) );
  AOI22_X1 U11277 ( .A1(n10201), .A2(n10217), .B1(n7000), .B2(n10200), .ZN(
        P1_U3489) );
  OAI211_X1 U11278 ( .C1(n10188), .C2(n10194), .A(n10187), .B(n10186), .ZN(
        n10189) );
  AOI21_X1 U11279 ( .B1(n10191), .B2(n10190), .A(n10189), .ZN(n10218) );
  AOI22_X1 U11280 ( .A1(n10201), .A2(n10218), .B1(n6109), .B2(n10200), .ZN(
        P1_U3492) );
  INV_X1 U11281 ( .A(n10192), .ZN(n10198) );
  OAI21_X1 U11282 ( .B1(n10195), .B2(n10194), .A(n10193), .ZN(n10197) );
  AOI211_X1 U11283 ( .C1(n10199), .C2(n10198), .A(n10197), .B(n10196), .ZN(
        n10220) );
  AOI22_X1 U11284 ( .A1(n10201), .A2(n10220), .B1(n7283), .B2(n10200), .ZN(
        P1_U3495) );
  AOI22_X1 U11285 ( .A1(n10221), .A2(n10202), .B1(n6128), .B2(n10219), .ZN(
        P1_U3522) );
  AOI22_X1 U11286 ( .A1(n10221), .A2(n10203), .B1(n6182), .B2(n10219), .ZN(
        P1_U3523) );
  AOI22_X1 U11287 ( .A1(n10221), .A2(n10205), .B1(n10204), .B2(n10219), .ZN(
        P1_U3524) );
  AOI22_X1 U11288 ( .A1(n10221), .A2(n10206), .B1(n6315), .B2(n10219), .ZN(
        P1_U3525) );
  AOI22_X1 U11289 ( .A1(n10221), .A2(n10208), .B1(n10207), .B2(n10219), .ZN(
        P1_U3526) );
  AOI22_X1 U11290 ( .A1(n10221), .A2(n10209), .B1(n6480), .B2(n10219), .ZN(
        P1_U3527) );
  AOI22_X1 U11291 ( .A1(n10221), .A2(n10210), .B1(n6636), .B2(n10219), .ZN(
        P1_U3528) );
  AOI22_X1 U11292 ( .A1(n10221), .A2(n10211), .B1(n6706), .B2(n10219), .ZN(
        P1_U3529) );
  AOI22_X1 U11293 ( .A1(n10221), .A2(n10212), .B1(n6057), .B2(n10219), .ZN(
        P1_U3530) );
  AOI22_X1 U11294 ( .A1(n10221), .A2(n10213), .B1(n6857), .B2(n10219), .ZN(
        P1_U3531) );
  AOI22_X1 U11295 ( .A1(n10221), .A2(n10214), .B1(n6874), .B2(n10219), .ZN(
        P1_U3532) );
  AOI22_X1 U11296 ( .A1(n10221), .A2(n10215), .B1(n6673), .B2(n10219), .ZN(
        P1_U3533) );
  AOI22_X1 U11297 ( .A1(n10221), .A2(n10217), .B1(n10216), .B2(n10219), .ZN(
        P1_U3534) );
  AOI22_X1 U11298 ( .A1(n10221), .A2(n10218), .B1(n6110), .B2(n10219), .ZN(
        P1_U3535) );
  AOI22_X1 U11299 ( .A1(n10221), .A2(n10220), .B1(n9357), .B2(n10219), .ZN(
        P1_U3536) );
  INV_X1 U11300 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10232) );
  INV_X1 U11301 ( .A(n10222), .ZN(n10225) );
  OAI21_X1 U11302 ( .B1(n10225), .B2(n10224), .A(n10223), .ZN(n10230) );
  AOI222_X1 U11303 ( .A1(n10233), .A2(n10230), .B1(n10229), .B2(n10228), .C1(
        n10227), .C2(n10226), .ZN(n10231) );
  OAI21_X1 U11304 ( .B1(n10233), .B2(n10232), .A(n10231), .ZN(P2_U3224) );
  INV_X1 U11305 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10240) );
  INV_X1 U11306 ( .A(n10234), .ZN(n10239) );
  OAI22_X1 U11307 ( .A1(n10237), .A2(n10236), .B1(n10270), .B2(n10235), .ZN(
        n10238) );
  NOR2_X1 U11308 ( .A1(n10239), .A2(n10238), .ZN(n10279) );
  AOI22_X1 U11309 ( .A1(n10277), .A2(n10240), .B1(n10279), .B2(n10275), .ZN(
        P2_U3393) );
  INV_X1 U11310 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U11311 ( .A1(n10277), .A2(n10242), .B1(n10241), .B2(n10275), .ZN(
        P2_U3396) );
  INV_X1 U11312 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10249) );
  NAND2_X1 U11313 ( .A1(n10243), .A2(n10274), .ZN(n10247) );
  NAND2_X1 U11314 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  AND3_X1 U11315 ( .A1(n10248), .A2(n10247), .A3(n10246), .ZN(n10281) );
  AOI22_X1 U11316 ( .A1(n10277), .A2(n10249), .B1(n10281), .B2(n10275), .ZN(
        P2_U3399) );
  INV_X1 U11317 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10255) );
  INV_X1 U11318 ( .A(n10250), .ZN(n10254) );
  OAI22_X1 U11319 ( .A1(n10252), .A2(n10263), .B1(n10251), .B2(n10270), .ZN(
        n10253) );
  NOR2_X1 U11320 ( .A1(n10254), .A2(n10253), .ZN(n10283) );
  AOI22_X1 U11321 ( .A1(n10277), .A2(n10255), .B1(n10283), .B2(n10275), .ZN(
        P2_U3402) );
  INV_X1 U11322 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10260) );
  NOR2_X1 U11323 ( .A1(n10256), .A2(n10270), .ZN(n10258) );
  AOI211_X1 U11324 ( .C1(n5763), .C2(n10259), .A(n10258), .B(n10257), .ZN(
        n10285) );
  AOI22_X1 U11325 ( .A1(n10277), .A2(n10260), .B1(n10285), .B2(n10275), .ZN(
        P2_U3405) );
  INV_X1 U11326 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10267) );
  INV_X1 U11327 ( .A(n10261), .ZN(n10266) );
  OAI22_X1 U11328 ( .A1(n10264), .A2(n10263), .B1(n10262), .B2(n10270), .ZN(
        n10265) );
  NOR2_X1 U11329 ( .A1(n10266), .A2(n10265), .ZN(n10287) );
  AOI22_X1 U11330 ( .A1(n10277), .A2(n10267), .B1(n10287), .B2(n10275), .ZN(
        P2_U3408) );
  INV_X1 U11331 ( .A(n10268), .ZN(n10273) );
  OAI21_X1 U11332 ( .B1(n10271), .B2(n10270), .A(n10269), .ZN(n10272) );
  AOI21_X1 U11333 ( .B1(n10274), .B2(n10273), .A(n10272), .ZN(n10288) );
  AOI22_X1 U11334 ( .A1(n10277), .A2(n10276), .B1(n10288), .B2(n10275), .ZN(
        P2_U3414) );
  AOI22_X1 U11335 ( .A1(n10289), .A2(n10279), .B1(n10278), .B2(n5770), .ZN(
        P2_U3460) );
  INV_X1 U11336 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U11337 ( .A1(n10289), .A2(n10281), .B1(n10280), .B2(n5770), .ZN(
        P2_U3462) );
  AOI22_X1 U11338 ( .A1(n10289), .A2(n10283), .B1(n10282), .B2(n5770), .ZN(
        P2_U3463) );
  INV_X1 U11339 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U11340 ( .A1(n10289), .A2(n10285), .B1(n10284), .B2(n5770), .ZN(
        P2_U3464) );
  AOI22_X1 U11341 ( .A1(n10289), .A2(n10287), .B1(n10286), .B2(n5770), .ZN(
        P2_U3465) );
  AOI22_X1 U11342 ( .A1(n10289), .A2(n10288), .B1(n5825), .B2(n5770), .ZN(
        P2_U3467) );
  INV_X1 U11343 ( .A(n10292), .ZN(n10291) );
  OAI222_X1 U11344 ( .A1(n5951), .A2(n10293), .B1(n5951), .B2(n10292), .C1(
        n10291), .C2(n10290), .ZN(ADD_1068_U5) );
  XOR2_X1 U11345 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11346 ( .B1(n10296), .B2(n10295), .A(n10294), .ZN(n10297) );
  XOR2_X1 U11347 ( .A(n10297), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55)
         );
  OAI21_X1 U11348 ( .B1(n10300), .B2(n10299), .A(n10298), .ZN(ADD_1068_U56) );
  OAI21_X1 U11349 ( .B1(n10303), .B2(n10302), .A(n10301), .ZN(ADD_1068_U57) );
  OAI21_X1 U11350 ( .B1(n10306), .B2(n10305), .A(n10304), .ZN(ADD_1068_U58) );
  OAI21_X1 U11351 ( .B1(n10309), .B2(n10308), .A(n10307), .ZN(ADD_1068_U59) );
  OAI21_X1 U11352 ( .B1(n10312), .B2(n10311), .A(n10310), .ZN(ADD_1068_U60) );
  OAI21_X1 U11353 ( .B1(n10315), .B2(n10314), .A(n10313), .ZN(ADD_1068_U61) );
  OAI21_X1 U11354 ( .B1(n10318), .B2(n10317), .A(n10316), .ZN(ADD_1068_U62) );
  OAI21_X1 U11355 ( .B1(n10321), .B2(n10320), .A(n10319), .ZN(ADD_1068_U63) );
  OAI21_X1 U11356 ( .B1(n10324), .B2(n10323), .A(n10322), .ZN(ADD_1068_U50) );
  OAI21_X1 U11357 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(ADD_1068_U51) );
  OAI21_X1 U11358 ( .B1(n10330), .B2(n10329), .A(n10328), .ZN(ADD_1068_U47) );
  OAI21_X1 U11359 ( .B1(n10333), .B2(n10332), .A(n10331), .ZN(ADD_1068_U49) );
  OAI21_X1 U11360 ( .B1(n10336), .B2(n10335), .A(n10334), .ZN(ADD_1068_U48) );
  AOI21_X1 U11361 ( .B1(n10339), .B2(n10338), .A(n10337), .ZN(ADD_1068_U54) );
  AOI21_X1 U11362 ( .B1(n10342), .B2(n10341), .A(n10340), .ZN(ADD_1068_U53) );
  OAI21_X1 U11363 ( .B1(n10345), .B2(n10344), .A(n10343), .ZN(ADD_1068_U52) );
  XNOR2_X1 U5011 ( .A(n5985), .B(n5984), .ZN(n9312) );
  NAND2_X1 U6398 ( .A1(n4854), .A2(n6520), .ZN(n10055) );
  INV_X1 U4942 ( .A(n7778), .ZN(n7705) );
  NOR2_X2 U4951 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5978) );
  CLKBUF_X1 U4991 ( .A(n9103), .Z(n4580) );
  CLKBUF_X2 U5049 ( .A(n5963), .Z(n4443) );
endmodule

