

module b20_C_gen_AntiSAT_k_256_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4511, n4512, n4513, n4515, n4516, n4517, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571;

  INV_X1 U5017 ( .A(n5706), .ZN(n5726) );
  INV_X2 U5018 ( .A(n6792), .ZN(n6741) );
  INV_X1 U5019 ( .A(n5728), .ZN(n5587) );
  INV_X1 U5020 ( .A(n7578), .ZN(n7584) );
  CLKBUF_X2 U5021 ( .A(n6337), .Z(n4513) );
  BUF_X2 U5022 ( .A(n6338), .Z(n4517) );
  CLKBUF_X1 U5023 ( .A(n7131), .Z(n4512) );
  NAND2_X2 U5024 ( .A1(n6795), .A2(n6318), .ZN(n6346) );
  XNOR2_X1 U5025 ( .A(n4833), .B(n7131), .ZN(n7024) );
  INV_X1 U5026 ( .A(n6056), .ZN(n5855) );
  NAND3_X1 U5027 ( .A1(n5552), .A2(n5556), .A3(n4918), .ZN(n5106) );
  NOR2_X1 U5028 ( .A1(n6074), .A2(n6073), .ZN(n6075) );
  INV_X1 U5029 ( .A(n8233), .ZN(n8293) );
  NOR3_X2 U5030 ( .A1(n5106), .A2(P1_IR_REG_14__SCAN_IN), .A3(
        P1_IR_REG_20__SCAN_IN), .ZN(n5105) );
  CLKBUF_X2 U5031 ( .A(n7133), .Z(n8277) );
  INV_X1 U5032 ( .A(n5708), .ZN(n5614) );
  NAND2_X1 U5033 ( .A1(n7923), .A2(n6001), .ZN(n6056) );
  INV_X2 U5034 ( .A(n6337), .ZN(n6393) );
  INV_X1 U5035 ( .A(n8310), .ZN(n9149) );
  AND3_X1 U5036 ( .A1(n5404), .A2(n5403), .A3(n5402), .ZN(n7674) );
  NAND2_X1 U5037 ( .A1(n4830), .A2(n4831), .ZN(n7306) );
  INV_X1 U5038 ( .A(n6346), .ZN(n6431) );
  INV_X2 U5039 ( .A(n6678), .ZN(n8565) );
  XNOR2_X1 U5040 ( .A(n6333), .B(n6332), .ZN(n7178) );
  AND2_X1 U5041 ( .A1(n7043), .A2(n7042), .ZN(n4511) );
  OAI21_X2 U5042 ( .B1(n8656), .B2(n8658), .A(n8655), .ZN(n8674) );
  NAND2_X2 U5043 ( .A1(n9104), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6095) );
  OAI21_X2 U5044 ( .B1(n7671), .B2(n4902), .A(n4643), .ZN(n8104) );
  OAI21_X2 U5045 ( .B1(n7577), .B2(n7618), .A(n4642), .ZN(n7671) );
  NAND3_X1 U5046 ( .A1(n5308), .A2(n5307), .A3(n4832), .ZN(n7131) );
  AOI21_X2 U5047 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n8072), .A(n8051), .ZN(
        n8052) );
  XOR2_X2 U5048 ( .A(n7975), .B(n7974), .Z(n7623) );
  NAND2_X1 U5049 ( .A1(n8345), .A2(n8330), .ZN(n6337) );
  XNOR2_X2 U5050 ( .A(n4680), .B(n6084), .ZN(n6673) );
  NAND2_X2 U5051 ( .A1(n6083), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4680) );
  BUF_X4 U5052 ( .A(n6344), .Z(n4515) );
  NAND2_X1 U5053 ( .A1(n6795), .A2(n6847), .ZN(n6344) );
  AND2_X1 U5054 ( .A1(n6745), .A2(n6744), .ZN(n4809) );
  AND2_X1 U5055 ( .A1(n8042), .A2(n6557), .ZN(n8172) );
  NAND2_X2 U5056 ( .A1(n6466), .A2(n6465), .ZN(n7440) );
  NAND2_X1 U5057 ( .A1(n9302), .A2(n7584), .ZN(n5897) );
  OR2_X1 U5058 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  NAND2_X1 U5059 ( .A1(n5399), .A2(n5220), .ZN(n5440) );
  NAND2_X1 U5060 ( .A1(n5339), .A2(n5338), .ZN(n7256) );
  NAND4_X1 U5061 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n9305)
         );
  INV_X2 U5063 ( .A(n8284), .ZN(n9148) );
  AND2_X1 U5064 ( .A1(n7240), .A2(n7034), .ZN(n8231) );
  AND2_X1 U5065 ( .A1(n7033), .A2(n5937), .ZN(n7146) );
  XNOR2_X1 U5066 ( .A(n5179), .B(n5178), .ZN(n9877) );
  CLKBUF_X1 U5067 ( .A(n5967), .Z(n9927) );
  AOI21_X1 U5068 ( .B1(n4639), .B2(n4641), .A(n4641), .ZN(n4636) );
  OAI21_X1 U5069 ( .B1(n4534), .B2(n4641), .A(n5582), .ZN(n4640) );
  CLKBUF_X2 U5070 ( .A(n6823), .Z(n6998) );
  INV_X1 U5071 ( .A(n5203), .ZN(n6318) );
  NOR2_X1 U5072 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5315) );
  AND2_X1 U5073 ( .A1(n9484), .A2(n9979), .ZN(n4854) );
  OAI21_X1 U5074 ( .B1(n4809), .B2(n8920), .A(n4807), .ZN(n4805) );
  INV_X1 U5075 ( .A(n4808), .ZN(n4807) );
  OR2_X1 U5076 ( .A1(n8328), .A2(n8927), .ZN(n6745) );
  NAND2_X1 U5077 ( .A1(n5117), .A2(n5116), .ZN(n5114) );
  NAND2_X1 U5078 ( .A1(n5596), .A2(n5837), .ZN(n9637) );
  NAND2_X1 U5079 ( .A1(n6031), .A2(n6030), .ZN(n9667) );
  AOI21_X1 U5080 ( .B1(n8344), .B2(n6431), .A(n6106), .ZN(n8949) );
  NAND2_X1 U5081 ( .A1(n4629), .A2(n4628), .ZN(n9127) );
  XNOR2_X1 U5082 ( .A(n5721), .B(n5720), .ZN(n8344) );
  NAND2_X1 U5083 ( .A1(n8043), .A2(n8199), .ZN(n8042) );
  NOR2_X1 U5084 ( .A1(n8107), .A2(n8106), .ZN(n8110) );
  AND2_X1 U5085 ( .A1(n8107), .A2(n8106), .ZN(n8108) );
  NAND2_X1 U5086 ( .A1(n4795), .A2(n4794), .ZN(n5146) );
  OR2_X1 U5087 ( .A1(n4531), .A2(n4903), .ZN(n4902) );
  NOR2_X1 U5088 ( .A1(n7821), .A2(n4728), .ZN(n7872) );
  NAND2_X1 U5089 ( .A1(n4702), .A2(n4701), .ZN(n7969) );
  NAND2_X1 U5090 ( .A1(n5442), .A2(n5441), .ZN(n6860) );
  INV_X1 U5091 ( .A(n7256), .ZN(n8338) );
  INV_X1 U5092 ( .A(n7572), .ZN(n9302) );
  INV_X1 U5093 ( .A(n7448), .ZN(n10038) );
  NAND2_X2 U5094 ( .A1(n7089), .A2(n7088), .ZN(n8198) );
  AND4_X2 U5095 ( .A1(n6294), .A2(n6293), .A3(n6292), .A4(n6291), .ZN(n8929)
         );
  NAND2_X1 U5096 ( .A1(n6308), .A2(n6307), .ZN(n10032) );
  AND2_X1 U5097 ( .A1(n9990), .A2(n9989), .ZN(n10002) );
  NAND2_X1 U5098 ( .A1(n7040), .A2(n4657), .ZN(n7133) );
  AND2_X2 U5099 ( .A1(n5306), .A2(n5305), .ZN(n5354) );
  INV_X4 U5100 ( .A(n6340), .ZN(n6372) );
  OAI21_X1 U5101 ( .B1(n5332), .B2(n4989), .A(n4988), .ZN(n5361) );
  AOI21_X1 U5102 ( .B1(n4750), .B2(n4752), .A(n4563), .ZN(n4749) );
  NAND2_X2 U5103 ( .A1(n7919), .A2(n7300), .ZN(n6792) );
  NAND2_X1 U5104 ( .A1(n6871), .A2(n6847), .ZN(n5706) );
  BUF_X4 U5105 ( .A(n6673), .Z(n8699) );
  CLKBUF_X2 U5106 ( .A(n6672), .Z(n4516) );
  XNOR2_X1 U5107 ( .A(n6491), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7300) );
  OR2_X1 U5108 ( .A1(n9868), .A2(n4641), .ZN(n5177) );
  XNOR2_X1 U5109 ( .A(n6499), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7919) );
  XNOR2_X1 U5110 ( .A(n5950), .B(n5949), .ZN(n7923) );
  NAND2_X1 U5111 ( .A1(n4637), .A2(n4636), .ZN(n5585) );
  NAND2_X1 U5112 ( .A1(n5301), .A2(n5300), .ZN(n5966) );
  NAND2_X1 U5113 ( .A1(n5300), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5179) );
  OR2_X1 U5114 ( .A1(n6097), .A2(n6096), .ZN(n6098) );
  NAND2_X1 U5115 ( .A1(n5298), .A2(n5175), .ZN(n5300) );
  INV_X4 U5116 ( .A(n6318), .ZN(n6847) );
  NOR2_X1 U5117 ( .A1(n5140), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5137) );
  AND2_X1 U5118 ( .A1(n4985), .A2(n6079), .ZN(n4695) );
  AND2_X1 U5119 ( .A1(n5085), .A2(n4987), .ZN(n4986) );
  NAND2_X1 U5120 ( .A1(n4674), .A2(n4678), .ZN(n9998) );
  AND2_X1 U5121 ( .A1(n6077), .A2(n6076), .ZN(n5085) );
  AND2_X1 U5122 ( .A1(n4920), .A2(n4919), .ZN(n5552) );
  NAND4_X1 U5123 ( .A1(n5364), .A2(n5092), .A3(n5163), .A4(n5315), .ZN(n5408)
         );
  INV_X1 U5124 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5949) );
  NOR2_X1 U5125 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6077) );
  INV_X1 U5126 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6416) );
  INV_X1 U5127 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6242) );
  INV_X1 U5128 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n10551) );
  INV_X1 U5129 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5037) );
  NOR2_X1 U5130 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6067) );
  INV_X1 U5131 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9473) );
  NOR2_X1 U5132 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n6068) );
  NOR2_X1 U5133 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6069) );
  INV_X1 U5134 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5736) );
  INV_X1 U5135 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5178) );
  NOR2_X2 U5136 ( .A1(n7134), .A2(n5152), .ZN(n7249) );
  AND2_X1 U5137 ( .A1(n7044), .A2(n7046), .ZN(n7134) );
  OR2_X1 U5138 ( .A1(n7033), .A2(n7039), .ZN(n9946) );
  NAND2_X1 U5139 ( .A1(n6678), .A2(n7306), .ZN(n6507) );
  AND4_X2 U5140 ( .A1(n6343), .A2(n5143), .A3(n6342), .A4(n6341), .ZN(n6678)
         );
  OAI21_X2 U5141 ( .B1(n7789), .B2(n7790), .A(n6544), .ZN(n7895) );
  NAND2_X1 U5142 ( .A1(n6099), .A2(n6100), .ZN(n6338) );
  NAND2_X4 U5143 ( .A1(n6100), .A2(n8345), .ZN(n6340) );
  INV_X1 U5145 ( .A(n9137), .ZN(n4917) );
  NAND2_X1 U5146 ( .A1(n6645), .A2(n6641), .ZN(n4700) );
  AND2_X1 U5147 ( .A1(n7822), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4728) );
  OR2_X1 U5148 ( .A1(n6772), .A2(n8555), .ZN(n6487) );
  OR2_X1 U5149 ( .A1(n9056), .A2(n8808), .ZN(n6610) );
  NAND2_X1 U5150 ( .A1(n5013), .A2(n5017), .ZN(n5286) );
  INV_X1 U5151 ( .A(n5018), .ZN(n5017) );
  AND2_X1 U5152 ( .A1(n5285), .A2(n5284), .ZN(n5689) );
  AND3_X1 U5153 ( .A1(n5736), .A2(n5952), .A3(n5949), .ZN(n5170) );
  INV_X1 U5154 ( .A(SI_9_), .ZN(n10290) );
  INV_X1 U5155 ( .A(n4517), .ZN(n6202) );
  OR2_X1 U5156 ( .A1(n6356), .A2(n6096), .ZN(n6400) );
  NAND2_X1 U5157 ( .A1(n8274), .A2(n8273), .ZN(n4654) );
  AOI21_X1 U5158 ( .B1(n4913), .B2(n4910), .A(n4909), .ZN(n4908) );
  INV_X1 U5159 ( .A(n4537), .ZN(n4910) );
  NAND2_X1 U5160 ( .A1(n5114), .A2(n5113), .ZN(n6035) );
  AND2_X1 U5161 ( .A1(n4566), .A2(n6033), .ZN(n5113) );
  NOR2_X1 U5162 ( .A1(n5154), .A2(n4550), .ZN(n5093) );
  XNOR2_X1 U5163 ( .A(n5957), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U5164 ( .A1(n5964), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U5165 ( .A1(n4688), .A2(n4687), .ZN(n6548) );
  NAND2_X1 U5166 ( .A1(n6537), .A2(n6792), .ZN(n4688) );
  NAND2_X1 U5167 ( .A1(n6538), .A2(n6741), .ZN(n4687) );
  NAND2_X1 U5168 ( .A1(n4613), .A2(n6741), .ZN(n4612) );
  INV_X1 U5169 ( .A(n6535), .ZN(n4613) );
  NAND2_X1 U5170 ( .A1(n4692), .A2(n4690), .ZN(n4689) );
  NOR2_X1 U5171 ( .A1(n4691), .A2(n6741), .ZN(n4690) );
  OAI22_X1 U5172 ( .A1(n4540), .A2(n6056), .B1(n4789), .B2(n4786), .ZN(n5840)
         );
  AND2_X1 U5173 ( .A1(n6694), .A2(n6693), .ZN(n4800) );
  NAND2_X1 U5174 ( .A1(n5249), .A2(n10229), .ZN(n5252) );
  NOR2_X1 U5175 ( .A1(n5466), .A2(n4774), .ZN(n4773) );
  INV_X1 U5176 ( .A(n5234), .ZN(n4774) );
  NOR2_X1 U5177 ( .A1(n5422), .A2(n4753), .ZN(n4752) );
  INV_X1 U5178 ( .A(n5225), .ZN(n4753) );
  NOR2_X1 U5179 ( .A1(n4980), .A2(n8720), .ZN(n4977) );
  INV_X1 U5180 ( .A(n4983), .ZN(n4980) );
  INV_X1 U5181 ( .A(n8345), .ZN(n6099) );
  OR2_X1 U5182 ( .A1(n9998), .A2(n6812), .ZN(n4677) );
  NAND2_X1 U5183 ( .A1(n7184), .A2(n7185), .ZN(n7183) );
  INV_X1 U5184 ( .A(n6541), .ZN(n4966) );
  OR2_X1 U5185 ( .A1(n10071), .A2(n8196), .ZN(n6551) );
  OR2_X1 U5186 ( .A1(n10067), .A2(n8133), .ZN(n6546) );
  OR2_X1 U5187 ( .A1(n9023), .A2(n8389), .ZN(n6632) );
  AOI21_X1 U5188 ( .B1(n4821), .B2(n6721), .A(n4820), .ZN(n4819) );
  NOR2_X1 U5189 ( .A1(n9035), .A2(n8789), .ZN(n4820) );
  OR2_X1 U5190 ( .A1(n9072), .A2(n8855), .ZN(n6577) );
  XNOR2_X1 U5191 ( .A(n6749), .B(n6748), .ZN(n5080) );
  INV_X1 U5192 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4694) );
  INV_X1 U5193 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5090) );
  AND2_X1 U5194 ( .A1(n8286), .A2(n8285), .ZN(n8288) );
  NOR2_X1 U5195 ( .A1(n7607), .A2(n7608), .ZN(n7618) );
  NOR4_X1 U5196 ( .A1(n5934), .A2(n5945), .A3(n5756), .A4(n5755), .ZN(n5759)
         );
  OR2_X1 U5197 ( .A1(n5732), .A2(n5731), .ZN(n5933) );
  INV_X1 U5198 ( .A(n5131), .ZN(n5128) );
  OR2_X1 U5199 ( .A1(n9798), .A2(n9292), .ZN(n5837) );
  OR2_X1 U5200 ( .A1(n7811), .A2(n7140), .ZN(n7039) );
  NAND2_X1 U5201 ( .A1(n4994), .A2(n5294), .ZN(n4993) );
  NAND2_X1 U5202 ( .A1(n4996), .A2(n4998), .ZN(n4994) );
  INV_X1 U5203 ( .A(n4997), .ZN(n4996) );
  AND2_X1 U5204 ( .A1(n5294), .A2(n5293), .ZN(n5598) );
  NAND2_X1 U5205 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  AND2_X1 U5206 ( .A1(n5281), .A2(n5280), .ZN(n5649) );
  NOR2_X1 U5207 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4918) );
  NAND2_X1 U5208 ( .A1(n5024), .A2(n4579), .ZN(n5023) );
  AOI21_X1 U5209 ( .B1(n4526), .B2(n5024), .A(n5022), .ZN(n5021) );
  NOR2_X1 U5210 ( .A1(n5254), .A2(n5255), .ZN(n5022) );
  OAI21_X1 U5211 ( .B1(n5509), .B2(n4757), .A(n4754), .ZN(n5539) );
  NOR2_X1 U5212 ( .A1(n4759), .A2(n4758), .ZN(n4757) );
  INV_X1 U5213 ( .A(n4755), .ZN(n4754) );
  NOR2_X1 U5214 ( .A1(n4763), .A2(n5523), .ZN(n4758) );
  NAND2_X1 U5215 ( .A1(n5497), .A2(n5245), .ZN(n5509) );
  AND2_X1 U5216 ( .A1(n4775), .A2(n5238), .ZN(n4771) );
  INV_X1 U5217 ( .A(n5479), .ZN(n4775) );
  INV_X1 U5218 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5163) );
  INV_X1 U5219 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5039) );
  INV_X1 U5220 ( .A(n6526), .ZN(n7727) );
  XNOR2_X1 U5221 ( .A(n8195), .B(n8196), .ZN(n8184) );
  AND2_X1 U5222 ( .A1(n4538), .A2(n6653), .ZN(n5033) );
  AOI21_X1 U5223 ( .B1(n6652), .B2(n6792), .A(n6651), .ZN(n6653) );
  AOI21_X1 U5224 ( .B1(n4700), .B2(n8393), .A(n6642), .ZN(n6655) );
  AND2_X1 U5225 ( .A1(n6162), .A2(n6161), .ZN(n8529) );
  NAND2_X1 U5226 ( .A1(n4723), .A2(n4724), .ZN(n7821) );
  OR2_X1 U5227 ( .A1(n10025), .A2(n4726), .ZN(n4723) );
  OR2_X1 U5228 ( .A1(n7715), .A2(n7796), .ZN(n4726) );
  XNOR2_X1 U5229 ( .A(n7693), .B(n7711), .ZN(n10021) );
  NOR2_X1 U5230 ( .A1(n7812), .A2(n4664), .ZN(n7866) );
  AND2_X1 U5231 ( .A1(n7822), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4664) );
  NOR2_X1 U5232 ( .A1(n8653), .A2(n5148), .ZN(n8684) );
  AND2_X1 U5233 ( .A1(n6124), .A2(n6091), .ZN(n8323) );
  AOI21_X1 U5234 ( .B1(n4827), .B2(n4826), .A(n4556), .ZN(n4825) );
  INV_X1 U5235 ( .A(n6717), .ZN(n4826) );
  OR2_X1 U5236 ( .A1(n8817), .A2(n8798), .ZN(n6612) );
  AND2_X1 U5237 ( .A1(n6610), .A2(n6603), .ZN(n4974) );
  AND3_X1 U5238 ( .A1(n6186), .A2(n6185), .A3(n6184), .ZN(n8809) );
  OR2_X1 U5239 ( .A1(n7214), .A2(n7213), .ZN(n7216) );
  OAI21_X1 U5240 ( .B1(n9876), .B2(n6346), .A(n6113), .ZN(n6772) );
  XNOR2_X1 U5241 ( .A(n6737), .B(n6733), .ZN(n8328) );
  AND2_X1 U5242 ( .A1(n6632), .A2(n6633), .ZN(n8749) );
  NAND2_X1 U5243 ( .A1(n9041), .A2(n8799), .ZN(n8771) );
  AND2_X1 U5244 ( .A1(n6179), .A2(n8776), .ZN(n8770) );
  OR2_X1 U5245 ( .A1(n9062), .A2(n8854), .ZN(n6603) );
  NAND2_X1 U5246 ( .A1(n8848), .A2(n6578), .ZN(n8838) );
  AOI21_X1 U5247 ( .B1(n4972), .B2(n4521), .A(n4970), .ZN(n4969) );
  INV_X1 U5248 ( .A(n4515), .ZN(n6446) );
  NAND2_X2 U5249 ( .A1(n6779), .A2(n6735), .ZN(n8914) );
  INV_X1 U5250 ( .A(n9120), .ZN(n6753) );
  NAND2_X1 U5251 ( .A1(n6092), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4679) );
  INV_X1 U5252 ( .A(n9944), .ZN(n4833) );
  AOI21_X1 U5253 ( .B1(n4652), .B2(n4551), .A(n4650), .ZN(n4649) );
  INV_X1 U5254 ( .A(n9216), .ZN(n4650) );
  NAND2_X1 U5255 ( .A1(n7248), .A2(n7247), .ZN(n4619) );
  NOR2_X1 U5256 ( .A1(n6007), .A2(n9487), .ZN(n9478) );
  AND2_X1 U5257 ( .A1(n5868), .A2(n5998), .ZN(n9505) );
  INV_X1 U5258 ( .A(n9288), .ZN(n9524) );
  AOI21_X1 U5259 ( .B1(n5118), .B2(n6032), .A(n4555), .ZN(n5116) );
  NOR2_X1 U5260 ( .A1(n4544), .A2(n5096), .ZN(n5095) );
  INV_X1 U5261 ( .A(n6026), .ZN(n5096) );
  NAND2_X1 U5262 ( .A1(n5691), .A2(n5690), .ZN(n9763) );
  OR2_X1 U5263 ( .A1(n7175), .A2(n7140), .ZN(n9969) );
  INV_X1 U5264 ( .A(n4907), .ZN(n4906) );
  OR2_X1 U5265 ( .A1(n5733), .A2(n4641), .ZN(n4904) );
  OAI21_X1 U5266 ( .B1(n4535), .B2(n4641), .A(n5171), .ZN(n4907) );
  AND2_X1 U5267 ( .A1(n5272), .A2(n5271), .ZN(n5630) );
  AND2_X1 U5268 ( .A1(n5233), .A2(n5231), .ZN(n5029) );
  AND2_X1 U5269 ( .A1(n6369), .A2(n6368), .ZN(n10013) );
  NAND2_X1 U5270 ( .A1(n6123), .A2(n6122), .ZN(n8743) );
  NAND2_X1 U5271 ( .A1(n9014), .A2(n10099), .ZN(n8952) );
  NOR2_X1 U5272 ( .A1(n4686), .A2(n4685), .ZN(n4684) );
  NAND2_X1 U5273 ( .A1(n6542), .A2(n6741), .ZN(n4685) );
  INV_X1 U5274 ( .A(n6553), .ZN(n4686) );
  NAND2_X1 U5275 ( .A1(n4615), .A2(n6792), .ZN(n4614) );
  INV_X1 U5276 ( .A(n6536), .ZN(n4615) );
  OAI21_X1 U5277 ( .B1(n6548), .B2(n6547), .A(n4682), .ZN(n4681) );
  AND2_X1 U5278 ( .A1(n6551), .A2(n4568), .ZN(n4682) );
  INV_X1 U5279 ( .A(n6703), .ZN(n4611) );
  INV_X1 U5280 ( .A(n5818), .ZN(n4791) );
  AOI21_X1 U5281 ( .B1(n5849), .B2(n5848), .A(n4744), .ZN(n4743) );
  NOR2_X1 U5282 ( .A1(n5991), .A2(n6056), .ZN(n4742) );
  NAND2_X1 U5283 ( .A1(n4565), .A2(n4817), .ZN(n4816) );
  NAND2_X1 U5284 ( .A1(n6727), .A2(n4818), .ZN(n4817) );
  INV_X1 U5285 ( .A(n4819), .ZN(n4818) );
  INV_X1 U5286 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6071) );
  NOR2_X1 U5287 ( .A1(n8014), .A2(n4873), .ZN(n4872) );
  INV_X1 U5288 ( .A(n5910), .ZN(n4873) );
  NOR2_X1 U5289 ( .A1(n5103), .A2(n5100), .ZN(n5099) );
  INV_X1 U5290 ( .A(n7465), .ZN(n5103) );
  NAND2_X1 U5291 ( .A1(n5059), .A2(n5058), .ZN(n5057) );
  INV_X1 U5292 ( .A(n8419), .ZN(n5058) );
  NAND2_X1 U5293 ( .A1(n4677), .A2(n4527), .ZN(n9993) );
  OR2_X1 U5294 ( .A1(n7004), .A2(n6831), .ZN(n7180) );
  NAND2_X1 U5295 ( .A1(n7180), .A2(n7181), .ZN(n7179) );
  NAND2_X1 U5296 ( .A1(n7183), .A2(n6816), .ZN(n7358) );
  NOR2_X1 U5297 ( .A1(n6381), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6356) );
  NOR2_X1 U5298 ( .A1(n4816), .A2(n4814), .ZN(n4813) );
  INV_X1 U5299 ( .A(n6718), .ZN(n4814) );
  INV_X1 U5300 ( .A(n4816), .ZN(n4811) );
  AOI21_X1 U5301 ( .B1(n4799), .B2(n4798), .A(n4557), .ZN(n4797) );
  INV_X1 U5302 ( .A(n6693), .ZN(n4798) );
  NAND2_X1 U5303 ( .A1(n4796), .A2(n4799), .ZN(n4795) );
  INV_X1 U5304 ( .A(n6519), .ZN(n4950) );
  NAND2_X1 U5305 ( .A1(n7727), .A2(n10044), .ZN(n6686) );
  NAND2_X1 U5306 ( .A1(n6526), .A2(n7506), .ZN(n6687) );
  NOR2_X1 U5307 ( .A1(n6722), .A2(n4822), .ZN(n4821) );
  INV_X1 U5308 ( .A(n6720), .ZN(n4822) );
  OR2_X1 U5309 ( .A1(n9035), .A2(n8475), .ZN(n6626) );
  OR2_X1 U5310 ( .A1(n8988), .A2(n8466), .ZN(n6578) );
  NOR2_X1 U5311 ( .A1(n6777), .A2(n9103), .ZN(n7105) );
  CLKBUF_X1 U5312 ( .A(n6229), .Z(n6259) );
  INV_X1 U5313 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U5314 ( .A1(n9232), .A2(n4631), .ZN(n4630) );
  OR2_X1 U5315 ( .A1(n8228), .A2(n8229), .ZN(n4631) );
  OAI21_X1 U5316 ( .B1(n5872), .B2(n4782), .A(n4780), .ZN(n5942) );
  NAND2_X1 U5317 ( .A1(n4784), .A2(n6050), .ZN(n4782) );
  AOI21_X1 U5318 ( .B1(n4784), .B2(n4781), .A(n4777), .ZN(n4780) );
  INV_X1 U5319 ( .A(n9877), .ZN(n5305) );
  NAND2_X1 U5320 ( .A1(n4708), .A2(n4707), .ZN(n6007) );
  NOR2_X1 U5321 ( .A1(n9538), .A2(n9529), .ZN(n4708) );
  OR2_X1 U5322 ( .A1(n9529), .A2(n9537), .ZN(n5764) );
  AND2_X1 U5323 ( .A1(n5134), .A2(n6039), .ZN(n5127) );
  NOR2_X1 U5324 ( .A1(n9734), .A2(n9812), .ZN(n4718) );
  AND2_X1 U5325 ( .A1(n8155), .A2(n9976), .ZN(n8154) );
  NAND2_X1 U5326 ( .A1(n7907), .A2(n4872), .ZN(n4871) );
  AND2_X1 U5327 ( .A1(n4523), .A2(n6024), .ZN(n4714) );
  NOR2_X1 U5328 ( .A1(n7776), .A2(n4840), .ZN(n4839) );
  INV_X1 U5329 ( .A(n5903), .ZN(n4840) );
  NOR2_X1 U5330 ( .A1(n5112), .A2(n5109), .ZN(n5108) );
  INV_X1 U5331 ( .A(n7656), .ZN(n5109) );
  INV_X1 U5332 ( .A(n7642), .ZN(n5112) );
  INV_X1 U5333 ( .A(n6020), .ZN(n5111) );
  AND2_X1 U5334 ( .A1(n7546), .A2(n7630), .ZN(n7545) );
  NAND2_X1 U5335 ( .A1(n7404), .A2(n5891), .ZN(n5896) );
  OR2_X1 U5336 ( .A1(n9305), .A2(n8338), .ZN(n5091) );
  AND2_X1 U5337 ( .A1(n9571), .A2(n9838), .ZN(n9555) );
  AND2_X1 U5338 ( .A1(n9589), .A2(n9576), .ZN(n9571) );
  INV_X1 U5339 ( .A(n5173), .ZN(n5141) );
  INV_X1 U5340 ( .A(n5168), .ZN(n4875) );
  INV_X1 U5341 ( .A(n5290), .ZN(n4998) );
  AND2_X1 U5342 ( .A1(n5290), .A2(n5289), .ZN(n5611) );
  NAND2_X1 U5343 ( .A1(n5001), .A2(n4999), .ZN(n5619) );
  AOI21_X1 U5344 ( .B1(n5003), .B2(n5006), .A(n5000), .ZN(n4999) );
  INV_X1 U5345 ( .A(n5272), .ZN(n5000) );
  AND2_X1 U5346 ( .A1(n5276), .A2(n5275), .ZN(n5620) );
  INV_X1 U5347 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5952) );
  INV_X1 U5348 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U5349 ( .A1(n5453), .A2(n4773), .ZN(n4772) );
  INV_X1 U5350 ( .A(n5197), .ZN(n4991) );
  OAI21_X1 U5351 ( .B1(n6847), .B2(n5206), .A(n5205), .ZN(n5209) );
  OR2_X1 U5352 ( .A1(n6318), .A2(n5204), .ZN(n5205) );
  AND2_X1 U5353 ( .A1(n7852), .A2(n7851), .ZN(n7858) );
  INV_X1 U5354 ( .A(n5055), .ZN(n5054) );
  OAI21_X1 U5355 ( .B1(n5057), .B2(n5062), .A(n5056), .ZN(n5055) );
  OR2_X1 U5356 ( .A1(n8418), .A2(n8530), .ZN(n5056) );
  NAND2_X1 U5357 ( .A1(n8454), .A2(n4584), .ZN(n8462) );
  AOI21_X1 U5358 ( .B1(n8502), .B2(n8503), .A(n8382), .ZN(n8473) );
  NOR2_X1 U5359 ( .A1(n5046), .A2(n5042), .ZN(n5041) );
  INV_X1 U5360 ( .A(n8511), .ZN(n5042) );
  INV_X1 U5361 ( .A(n8411), .ZN(n5046) );
  NAND2_X1 U5362 ( .A1(n8411), .A2(n5045), .ZN(n5044) );
  INV_X1 U5363 ( .A(n8371), .ZN(n5045) );
  NAND2_X1 U5364 ( .A1(n7522), .A2(n7521), .ZN(n7593) );
  NOR2_X1 U5365 ( .A1(n8398), .A2(n5084), .ZN(n5083) );
  AOI21_X1 U5366 ( .B1(n4983), .B2(n4548), .A(n4979), .ZN(n4978) );
  AND2_X1 U5367 ( .A1(n6118), .A2(n6105), .ZN(n8553) );
  AND4_X1 U5368 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n7590)
         );
  NAND2_X1 U5369 ( .A1(n6300), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6312) );
  OR2_X1 U5370 ( .A1(n4517), .A2(n6302), .ZN(n6309) );
  OR2_X1 U5371 ( .A1(n4513), .A2(n6303), .ZN(n6310) );
  OR2_X1 U5372 ( .A1(n6340), .A2(n6301), .ZN(n6311) );
  NAND2_X1 U5373 ( .A1(n6984), .A2(n6814), .ZN(n4665) );
  NAND2_X1 U5374 ( .A1(n4666), .A2(n6984), .ZN(n4669) );
  NOR2_X1 U5375 ( .A1(n7015), .A2(n4667), .ZN(n4666) );
  INV_X1 U5376 ( .A(n6814), .ZN(n4667) );
  XNOR2_X1 U5377 ( .A(n7358), .B(n7342), .ZN(n6817) );
  NOR2_X1 U5378 ( .A1(n6817), .A2(n6280), .ZN(n7361) );
  NOR2_X1 U5379 ( .A1(n8071), .A2(n4671), .ZN(n8073) );
  NOR2_X1 U5380 ( .A1(n7888), .A2(n6420), .ZN(n4671) );
  NAND2_X1 U5381 ( .A1(n4922), .A2(n4921), .ZN(n8567) );
  NAND2_X1 U5382 ( .A1(n8074), .A2(n4926), .ZN(n4921) );
  OR2_X1 U5383 ( .A1(n8085), .A2(n4923), .ZN(n4922) );
  NAND2_X1 U5384 ( .A1(n4926), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4923) );
  AOI21_X1 U5385 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8570), .A(n8569), .ZN(
        n8586) );
  OR2_X1 U5386 ( .A1(n8568), .A2(n9003), .ZN(n4932) );
  INV_X1 U5387 ( .A(n8601), .ZN(n4931) );
  OR2_X1 U5388 ( .A1(n8568), .A2(n4930), .ZN(n4927) );
  OR2_X1 U5389 ( .A1(n8603), .A2(n9003), .ZN(n4930) );
  NAND2_X1 U5390 ( .A1(n8601), .A2(n4929), .ZN(n4928) );
  INV_X1 U5391 ( .A(n8603), .ZN(n4929) );
  AOI21_X1 U5392 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8619), .A(n8610), .ZN(
        n8628) );
  XNOR2_X1 U5393 ( .A(n8667), .B(n8685), .ZN(n8659) );
  NAND2_X1 U5394 ( .A1(n4670), .A2(n4536), .ZN(n4941) );
  NAND2_X1 U5395 ( .A1(n4941), .A2(n4942), .ZN(n4940) );
  NOR2_X1 U5396 ( .A1(n4961), .A2(n4959), .ZN(n4958) );
  INV_X1 U5397 ( .A(n6628), .ZN(n4959) );
  AND3_X1 U5398 ( .A1(n6196), .A2(n6195), .A3(n6194), .ZN(n8798) );
  AND2_X1 U5399 ( .A1(n6481), .A2(n6616), .ZN(n8795) );
  INV_X1 U5400 ( .A(n8795), .ZN(n8801) );
  AND4_X1 U5401 ( .A1(n6206), .A2(n6205), .A3(n6204), .A4(n6203), .ZN(n8808)
         );
  OR2_X1 U5402 ( .A1(n6424), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6437) );
  AOI21_X1 U5403 ( .B1(n4965), .B2(n6471), .A(n4964), .ZN(n4963) );
  INV_X1 U5404 ( .A(n6546), .ZN(n4964) );
  NAND2_X1 U5405 ( .A1(n8135), .A2(n7969), .ZN(n6541) );
  OR2_X1 U5406 ( .A1(n7854), .A2(n10053), .ZN(n6693) );
  NAND2_X1 U5407 ( .A1(n6686), .A2(n6687), .ZN(n7501) );
  INV_X1 U5408 ( .A(n8911), .ZN(n8930) );
  NAND2_X1 U5409 ( .A1(n8757), .A2(n6629), .ZN(n4960) );
  OR2_X1 U5410 ( .A1(n9029), .A2(n8529), .ZN(n6628) );
  AND2_X1 U5411 ( .A1(n6626), .A2(n6622), .ZN(n8775) );
  INV_X1 U5412 ( .A(n6616), .ZN(n4947) );
  AND2_X1 U5413 ( .A1(n6481), .A2(n4945), .ZN(n4944) );
  NAND2_X1 U5414 ( .A1(n6616), .A2(n4946), .ZN(n4945) );
  OR2_X1 U5415 ( .A1(n8825), .A2(n8826), .ZN(n8827) );
  AND2_X1 U5416 ( .A1(n6610), .A2(n8813), .ZN(n8826) );
  NOR2_X1 U5417 ( .A1(n4586), .A2(n4802), .ZN(n4801) );
  NAND2_X1 U5418 ( .A1(n8838), .A2(n8839), .ZN(n8837) );
  AND2_X1 U5419 ( .A1(n6603), .A2(n6601), .ZN(n8839) );
  NAND2_X1 U5420 ( .A1(n6583), .A2(n6582), .ZN(n4951) );
  INV_X1 U5421 ( .A(n4954), .ZN(n4953) );
  NOR2_X1 U5422 ( .A1(n6579), .A2(n4957), .ZN(n4956) );
  INV_X1 U5423 ( .A(n6574), .ZN(n4957) );
  OR2_X1 U5424 ( .A1(n9084), .A2(n8399), .ZN(n6574) );
  INV_X1 U5425 ( .A(n4973), .ZN(n4972) );
  OAI21_X1 U5426 ( .B1(n4521), .B2(n8171), .A(n4542), .ZN(n4973) );
  AND2_X1 U5427 ( .A1(n6570), .A2(n6569), .ZN(n8895) );
  NAND2_X1 U5428 ( .A1(n8172), .A2(n8171), .ZN(n8170) );
  INV_X1 U5429 ( .A(n7969), .ZN(n10059) );
  INV_X1 U5430 ( .A(n7735), .ZN(n10048) );
  OR2_X1 U5431 ( .A1(n7919), .A2(n7300), .ZN(n10073) );
  NAND2_X1 U5432 ( .A1(n5077), .A2(n6753), .ZN(n6752) );
  INV_X1 U5433 ( .A(n5080), .ZN(n5079) );
  NOR3_X1 U5434 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U5435 ( .A1(n6662), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6668) );
  INV_X1 U5436 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U5437 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4676) );
  AND2_X1 U5438 ( .A1(n8313), .A2(n8312), .ZN(n9161) );
  INV_X1 U5439 ( .A(n8110), .ZN(n4635) );
  NAND2_X1 U5440 ( .A1(n8216), .A2(n8121), .ZN(n4887) );
  INV_X1 U5441 ( .A(n9896), .ZN(n4883) );
  INV_X1 U5442 ( .A(n9294), .ZN(n9179) );
  NOR2_X1 U5443 ( .A1(n4901), .A2(n4531), .ZN(n4644) );
  NOR2_X1 U5444 ( .A1(n9165), .A2(n9166), .ZN(n8274) );
  NOR2_X1 U5445 ( .A1(n8255), .A2(n4899), .ZN(n4898) );
  INV_X1 U5446 ( .A(n9206), .ZN(n4899) );
  AND2_X1 U5447 ( .A1(n7617), .A2(n4571), .ZN(n4642) );
  INV_X1 U5448 ( .A(n7616), .ZN(n7617) );
  AOI211_X1 U5449 ( .C1(n5738), .C2(n5933), .A(n5739), .B(n6004), .ZN(n5757)
         );
  AND4_X1 U5450 ( .A1(n5421), .A2(n5420), .A3(n5419), .A4(n5418), .ZN(n7985)
         );
  AND4_X1 U5451 ( .A1(n5378), .A2(n5377), .A3(n5376), .A4(n5375), .ZN(n7572)
         );
  NAND2_X1 U5452 ( .A1(n4857), .A2(n4856), .ZN(n9519) );
  AOI21_X1 U5453 ( .B1(n4859), .B2(n4862), .A(n5753), .ZN(n4856) );
  AOI21_X1 U5454 ( .B1(n4861), .B2(n4860), .A(n9520), .ZN(n4859) );
  INV_X1 U5455 ( .A(n4708), .ZN(n9516) );
  NOR2_X1 U5456 ( .A1(n6046), .A2(n5122), .ZN(n5121) );
  INV_X1 U5457 ( .A(n6044), .ZN(n5122) );
  AND2_X1 U5458 ( .A1(n5653), .A2(n5693), .ZN(n9558) );
  AOI21_X1 U5459 ( .B1(n9580), .B2(n5994), .A(n5993), .ZN(n9550) );
  INV_X1 U5460 ( .A(n9609), .ZN(n9569) );
  NOR2_X1 U5461 ( .A1(n5132), .A2(n4554), .ZN(n5131) );
  NOR2_X1 U5462 ( .A1(n6037), .A2(n5133), .ZN(n5132) );
  NAND2_X1 U5463 ( .A1(n5136), .A2(n6036), .ZN(n5133) );
  NOR2_X1 U5464 ( .A1(n6037), .A2(n5135), .ZN(n5134) );
  INV_X1 U5465 ( .A(n5136), .ZN(n5135) );
  AND2_X1 U5466 ( .A1(n5851), .A2(n9565), .ZN(n9582) );
  NAND2_X1 U5467 ( .A1(n4844), .A2(n4846), .ZN(n9606) );
  INV_X1 U5468 ( .A(n4847), .ZN(n4846) );
  OAI21_X1 U5469 ( .B1(n5988), .B2(n4848), .A(n9607), .ZN(n4847) );
  NAND2_X1 U5470 ( .A1(n9848), .A2(n9246), .ZN(n5136) );
  NAND2_X1 U5471 ( .A1(n9637), .A2(n9635), .ZN(n9618) );
  NAND2_X1 U5472 ( .A1(n9618), .A2(n5988), .ZN(n9619) );
  NAND2_X1 U5473 ( .A1(n5966), .A2(n7136), .ZN(n9664) );
  AND2_X1 U5474 ( .A1(n5589), .A2(n5588), .ZN(n9652) );
  NAND2_X1 U5475 ( .A1(n9674), .A2(n9661), .ZN(n5118) );
  NOR2_X1 U5476 ( .A1(n9674), .A2(n9661), .ZN(n6032) );
  NAND2_X1 U5477 ( .A1(n9685), .A2(n4547), .ZN(n9675) );
  NAND2_X1 U5478 ( .A1(n9690), .A2(n9702), .ZN(n6030) );
  NAND2_X1 U5479 ( .A1(n7903), .A2(n6025), .ZN(n6027) );
  OR2_X1 U5480 ( .A1(n9299), .A2(n9921), .ZN(n6020) );
  NAND2_X1 U5481 ( .A1(n7655), .A2(n7656), .ZN(n7654) );
  NAND2_X1 U5482 ( .A1(n7408), .A2(n6018), .ZN(n7377) );
  NAND2_X1 U5483 ( .A1(n7377), .A2(n7379), .ZN(n7376) );
  NAND2_X1 U5484 ( .A1(n7226), .A2(n5091), .ZN(n7154) );
  NAND2_X1 U5485 ( .A1(n9944), .A2(n9888), .ZN(n7153) );
  OAI21_X1 U5486 ( .B1(n9876), .B2(n5706), .A(n5705), .ZN(n9487) );
  INV_X1 U5487 ( .A(n9576), .ZN(n9773) );
  INV_X1 U5488 ( .A(n9134), .ZN(n9976) );
  NAND2_X1 U5489 ( .A1(n5504), .A2(n5503), .ZN(n8212) );
  NAND2_X1 U5490 ( .A1(n5704), .A2(n5297), .ZN(n5721) );
  NAND2_X1 U5491 ( .A1(n5703), .A2(SI_29_), .ZN(n5704) );
  XNOR2_X1 U5492 ( .A(n5302), .B(n5174), .ZN(n5967) );
  NAND2_X1 U5493 ( .A1(n4713), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5302) );
  NOR2_X1 U5494 ( .A1(n5173), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5138) );
  INV_X1 U5495 ( .A(n5016), .ZN(n5688) );
  AOI21_X1 U5496 ( .B1(n5648), .B2(n5649), .A(n5019), .ZN(n5016) );
  INV_X1 U5497 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5171) );
  AND2_X1 U5498 ( .A1(n5105), .A2(n5512), .ZN(n5733) );
  XNOR2_X1 U5499 ( .A(n5648), .B(n5649), .ZN(n9121) );
  NOR2_X1 U5500 ( .A1(n5638), .A2(n5012), .ZN(n5011) );
  INV_X1 U5501 ( .A(n5263), .ZN(n5012) );
  AOI21_X1 U5502 ( .B1(n5010), .B2(n5009), .A(n5008), .ZN(n5007) );
  AND2_X1 U5503 ( .A1(n5264), .A2(n5263), .ZN(n5010) );
  INV_X1 U5504 ( .A(n5268), .ZN(n5008) );
  INV_X1 U5505 ( .A(n5638), .ZN(n5009) );
  NAND2_X1 U5506 ( .A1(n5735), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U5507 ( .A(n5886), .B(P1_IR_REG_20__SCAN_IN), .ZN(n7140) );
  NOR2_X1 U5508 ( .A1(n5106), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U5509 ( .A1(n5020), .A2(n5024), .ZN(n5568) );
  NAND2_X1 U5510 ( .A1(n5539), .A2(n5027), .ZN(n5020) );
  NAND2_X1 U5511 ( .A1(n5512), .A2(n5169), .ZN(n5526) );
  OAI21_X1 U5512 ( .B1(n5539), .B2(n5246), .A(n5247), .ZN(n5551) );
  NAND2_X1 U5513 ( .A1(n4761), .A2(n4764), .ZN(n5525) );
  NAND2_X1 U5514 ( .A1(n5509), .A2(n4765), .ZN(n4761) );
  AOI21_X1 U5515 ( .B1(n4769), .B2(n4771), .A(n4768), .ZN(n4767) );
  INV_X1 U5516 ( .A(n4771), .ZN(n4770) );
  INV_X1 U5517 ( .A(n5240), .ZN(n4768) );
  NAND2_X1 U5518 ( .A1(n4748), .A2(n4746), .ZN(n5030) );
  AOI21_X1 U5519 ( .B1(n4749), .B2(n4751), .A(n4747), .ZN(n4746) );
  INV_X1 U5520 ( .A(n5406), .ZN(n4747) );
  NAND2_X1 U5521 ( .A1(n5442), .A2(n5225), .ZN(n5423) );
  NAND2_X1 U5522 ( .A1(n5440), .A2(n5439), .ZN(n5442) );
  AND2_X1 U5523 ( .A1(n5201), .A2(n5202), .ZN(n5344) );
  INV_X1 U5524 ( .A(n8559), .ZN(n8135) );
  NAND2_X1 U5525 ( .A1(n7290), .A2(n5089), .ZN(n7427) );
  AND2_X1 U5526 ( .A1(n7291), .A2(n7289), .ZN(n5089) );
  NAND2_X1 U5527 ( .A1(n7092), .A2(n8565), .ZN(n5081) );
  NAND2_X1 U5528 ( .A1(n6188), .A2(n6187), .ZN(n8817) );
  AND4_X1 U5529 ( .A1(n6428), .A2(n6427), .A3(n6426), .A4(n6425), .ZN(n8196)
         );
  AND3_X1 U5530 ( .A1(n6178), .A2(n6177), .A3(n6176), .ZN(n8799) );
  AND4_X1 U5531 ( .A1(n6216), .A2(n6215), .A3(n6214), .A4(n6213), .ZN(n8854)
         );
  AND2_X1 U5532 ( .A1(n7083), .A2(n7082), .ZN(n8538) );
  AND2_X1 U5533 ( .A1(n7114), .A2(n7113), .ZN(n8548) );
  XNOR2_X1 U5534 ( .A(n6208), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8705) );
  INV_X1 U5535 ( .A(n8799), .ZN(n8776) );
  INV_X1 U5536 ( .A(n7590), .ZN(n8562) );
  OAI21_X1 U5537 ( .B1(n9998), .B2(n6826), .A(n6827), .ZN(n10007) );
  AOI21_X1 U5538 ( .B1(n6801), .B2(n9998), .A(n10002), .ZN(n6981) );
  AND2_X1 U5539 ( .A1(n4725), .A2(n4729), .ZN(n7716) );
  INV_X1 U5540 ( .A(n7713), .ZN(n4725) );
  NAND2_X1 U5541 ( .A1(n4661), .A2(n4660), .ZN(n7812) );
  OR2_X1 U5542 ( .A1(n10021), .A2(n4662), .ZN(n4660) );
  OR2_X1 U5543 ( .A1(n7696), .A2(n6360), .ZN(n4662) );
  AND2_X1 U5544 ( .A1(n6404), .A2(n6415), .ZN(n7873) );
  OR2_X1 U5545 ( .A1(n8085), .A2(n8057), .ZN(n4925) );
  XNOR2_X1 U5546 ( .A(n8073), .B(n8097), .ZN(n8085) );
  OR2_X1 U5547 ( .A1(n8611), .A2(n8887), .ZN(n4733) );
  OR2_X1 U5548 ( .A1(n8654), .A2(n8991), .ZN(n4670) );
  OAI21_X1 U5549 ( .B1(n8668), .B2(n8661), .A(n8660), .ZN(n8663) );
  AND2_X1 U5550 ( .A1(n8659), .A2(n8866), .ZN(n8661) );
  AOI21_X1 U5551 ( .B1(n8665), .B2(n10020), .A(n4739), .ZN(n4738) );
  OAI21_X1 U5552 ( .B1(n8679), .B2(n8664), .A(n4740), .ZN(n4739) );
  AOI21_X1 U5553 ( .B1(n10018), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n4598), .ZN(
        n4740) );
  XNOR2_X1 U5554 ( .A(n8684), .B(n8685), .ZN(n8654) );
  OAI21_X1 U5555 ( .B1(n4942), .B2(n4941), .A(n4940), .ZN(n4939) );
  NAND2_X1 U5556 ( .A1(n8689), .A2(n8697), .ZN(n4938) );
  NOR2_X1 U5557 ( .A1(n4606), .A2(n4605), .ZN(n4604) );
  XNOR2_X1 U5558 ( .A(n4659), .B(n4593), .ZN(n4658) );
  NAND2_X1 U5559 ( .A1(n4940), .A2(n8695), .ZN(n4659) );
  OAI21_X1 U5560 ( .B1(n8328), .B2(n8327), .A(n8326), .ZN(n4808) );
  NAND2_X1 U5561 ( .A1(n6435), .A2(n6434), .ZN(n10084) );
  NAND2_X1 U5562 ( .A1(n6419), .A2(n6418), .ZN(n10071) );
  OR2_X1 U5563 ( .A1(n6346), .A2(n6853), .ZN(n4830) );
  NAND2_X1 U5564 ( .A1(n6086), .A2(n6085), .ZN(n9008) );
  INV_X1 U5565 ( .A(n6772), .ZN(n8324) );
  NAND2_X1 U5566 ( .A1(n6135), .A2(n6134), .ZN(n9016) );
  AOI21_X1 U5567 ( .B1(n8726), .B2(n8914), .A(n8725), .ZN(n9014) );
  NAND2_X1 U5568 ( .A1(n8724), .A2(n8723), .ZN(n8725) );
  XNOR2_X1 U5569 ( .A(n4601), .B(n4600), .ZN(n8751) );
  INV_X1 U5570 ( .A(n8749), .ZN(n4600) );
  NAND2_X1 U5571 ( .A1(n8748), .A2(n8747), .ZN(n4601) );
  NAND2_X1 U5572 ( .A1(n6173), .A2(n6172), .ZN(n9041) );
  NAND2_X1 U5573 ( .A1(n6448), .A2(n6447), .ZN(n9097) );
  XNOR2_X1 U5574 ( .A(n6359), .B(n6358), .ZN(n7822) );
  NOR2_X1 U5575 ( .A1(n8050), .A2(n9885), .ZN(n4879) );
  INV_X1 U5576 ( .A(n4622), .ZN(n4621) );
  AOI21_X1 U5577 ( .B1(n8318), .B2(n4623), .A(n4587), .ZN(n4622) );
  NOR2_X1 U5578 ( .A1(n8301), .A2(n9916), .ZN(n4623) );
  INV_X1 U5579 ( .A(n4915), .ZN(n4911) );
  AOI22_X1 U5580 ( .A1(n9148), .A2(n4512), .B1(n4833), .B2(n8233), .ZN(n7132)
         );
  NAND2_X1 U5581 ( .A1(n4648), .A2(n4646), .ZN(n9187) );
  AOI21_X1 U5582 ( .B1(n4649), .B2(n4653), .A(n4647), .ZN(n4646) );
  INV_X1 U5583 ( .A(n8292), .ZN(n4647) );
  NAND2_X1 U5584 ( .A1(n5677), .A2(n5676), .ZN(n9643) );
  NAND2_X1 U5585 ( .A1(n5641), .A2(n5640), .ZN(n9782) );
  INV_X1 U5586 ( .A(n7999), .ZN(n9299) );
  AND2_X1 U5587 ( .A1(n9476), .A2(n9746), .ZN(n9743) );
  NAND2_X1 U5588 ( .A1(n4522), .A2(n9724), .ZN(n4855) );
  AND2_X1 U5589 ( .A1(n5633), .A2(n5632), .ZN(n9843) );
  AND3_X1 U5590 ( .A1(n5352), .A2(n5351), .A3(n5350), .ZN(n7421) );
  NAND2_X1 U5591 ( .A1(n6510), .A2(n6741), .ZN(n6513) );
  NAND2_X1 U5592 ( .A1(n4683), .A2(n4681), .ZN(n6549) );
  OAI21_X1 U5593 ( .B1(n6548), .B2(n6543), .A(n4684), .ZN(n4683) );
  NAND2_X1 U5594 ( .A1(n6567), .A2(n4610), .ZN(n6568) );
  NAND2_X1 U5595 ( .A1(n6566), .A2(n4611), .ZN(n4610) );
  OR2_X1 U5596 ( .A1(n5810), .A2(n4790), .ZN(n5816) );
  AOI21_X1 U5597 ( .B1(n5835), .B2(n5921), .A(n5927), .ZN(n4789) );
  NAND2_X1 U5598 ( .A1(n5836), .A2(n4787), .ZN(n4786) );
  NOR2_X1 U5599 ( .A1(n4788), .A2(n5855), .ZN(n4787) );
  INV_X1 U5600 ( .A(n5925), .ZN(n4788) );
  INV_X1 U5601 ( .A(n6619), .ZN(n4616) );
  NAND2_X1 U5602 ( .A1(n4745), .A2(n4741), .ZN(n5854) );
  NAND2_X1 U5603 ( .A1(n5850), .A2(n6056), .ZN(n4745) );
  OAI21_X1 U5604 ( .B1(n4743), .B2(n5844), .A(n4742), .ZN(n4741) );
  AOI22_X1 U5605 ( .A1(n8675), .A2(n8674), .B1(n8685), .B2(n8673), .ZN(n8677)
         );
  AND2_X1 U5606 ( .A1(n6753), .A2(n5076), .ZN(n5075) );
  AND2_X1 U5607 ( .A1(n9048), .A2(n8788), .ZN(n6618) );
  OAI21_X1 U5608 ( .B1(n4778), .B2(n5882), .A(n4783), .ZN(n4777) );
  OR2_X1 U5609 ( .A1(n4785), .A2(n9828), .ZN(n4778) );
  AOI21_X1 U5610 ( .B1(n5881), .B2(n9828), .A(n5739), .ZN(n4783) );
  INV_X1 U5611 ( .A(n5876), .ZN(n4781) );
  NAND2_X1 U5612 ( .A1(n4779), .A2(n5880), .ZN(n4784) );
  NAND2_X1 U5613 ( .A1(n4776), .A2(n5877), .ZN(n4779) );
  NOR2_X1 U5614 ( .A1(n5766), .A2(n5765), .ZN(n5871) );
  AND2_X1 U5615 ( .A1(n5859), .A2(n6056), .ZN(n5765) );
  OAI21_X1 U5616 ( .B1(n5611), .B2(n4998), .A(n5598), .ZN(n4997) );
  NOR2_X1 U5617 ( .A1(n5015), .A2(n5019), .ZN(n5014) );
  INV_X1 U5618 ( .A(n5276), .ZN(n5015) );
  OAI21_X1 U5619 ( .B1(n5649), .B2(n5019), .A(n5689), .ZN(n5018) );
  AOI21_X1 U5620 ( .B1(n5007), .B2(n5005), .A(n5004), .ZN(n5003) );
  INV_X1 U5621 ( .A(n5630), .ZN(n5004) );
  INV_X1 U5622 ( .A(n5011), .ZN(n5005) );
  INV_X1 U5623 ( .A(n5007), .ZN(n5006) );
  INV_X1 U5624 ( .A(SI_18_), .ZN(n5255) );
  INV_X1 U5625 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5248) );
  INV_X1 U5626 ( .A(n4764), .ZN(n4763) );
  OAI21_X1 U5627 ( .B1(n4762), .B2(n5523), .A(n4756), .ZN(n4755) );
  NAND2_X1 U5628 ( .A1(n4759), .A2(n4766), .ZN(n4756) );
  AOI21_X1 U5629 ( .B1(n4766), .B2(n4764), .A(n4760), .ZN(n4762) );
  AND2_X1 U5630 ( .A1(n4764), .A2(n4760), .ZN(n4759) );
  AND2_X1 U5631 ( .A1(n8349), .A2(n8183), .ZN(n5068) );
  INV_X1 U5632 ( .A(n5066), .ZN(n5065) );
  OAI21_X1 U5633 ( .B1(n5069), .B2(n8347), .A(n8437), .ZN(n5066) );
  NAND2_X1 U5634 ( .A1(n5080), .A2(n5075), .ZN(n5073) );
  NAND2_X1 U5635 ( .A1(n6750), .A2(n5075), .ZN(n5072) );
  INV_X1 U5636 ( .A(n7084), .ZN(n5071) );
  INV_X1 U5637 ( .A(n8493), .ZN(n5084) );
  INV_X1 U5638 ( .A(n6485), .ZN(n4981) );
  NOR2_X1 U5639 ( .A1(n9008), .A2(n8949), .ZN(n4984) );
  INV_X1 U5640 ( .A(n6488), .ZN(n4979) );
  OR2_X1 U5641 ( .A1(n6648), .A2(n6647), .ZN(n6649) );
  INV_X1 U5642 ( .A(n4700), .ZN(n6646) );
  NAND2_X1 U5643 ( .A1(n6829), .A2(n7015), .ZN(n6830) );
  NAND2_X1 U5644 ( .A1(n7179), .A2(n6833), .ZN(n7346) );
  INV_X1 U5645 ( .A(n7715), .ZN(n4727) );
  NAND2_X1 U5646 ( .A1(n7709), .A2(n7708), .ZN(n7712) );
  INV_X1 U5647 ( .A(n8075), .ZN(n4926) );
  NOR2_X1 U5648 ( .A1(n6147), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U5649 ( .A1(n8826), .A2(n6717), .ZN(n4829) );
  NOR2_X1 U5650 ( .A1(n6224), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6199) );
  AND2_X1 U5651 ( .A1(n6251), .A2(n6089), .ZN(n6233) );
  NOR2_X1 U5652 ( .A1(n6275), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6251) );
  INV_X1 U5653 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10480) );
  NOR2_X1 U5654 ( .A1(n6437), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6436) );
  AND2_X1 U5655 ( .A1(n6350), .A2(n6088), .ZN(n6349) );
  NOR2_X1 U5656 ( .A1(n6376), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6350) );
  AND4_X1 U5657 ( .A1(n6312), .A2(n6311), .A3(n6309), .A4(n6310), .ZN(n6682)
         );
  NAND2_X1 U5658 ( .A1(n5074), .A2(n6881), .ZN(n7085) );
  OAI21_X1 U5659 ( .B1(n5080), .B2(n6750), .A(n5075), .ZN(n5074) );
  INV_X1 U5660 ( .A(n6626), .ZN(n6621) );
  INV_X1 U5661 ( .A(n6612), .ZN(n4946) );
  INV_X1 U5662 ( .A(n6713), .ZN(n4802) );
  OAI21_X1 U5663 ( .B1(n4956), .B2(n4955), .A(n6577), .ZN(n4954) );
  INV_X1 U5664 ( .A(n6570), .ZN(n4970) );
  NOR2_X1 U5665 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4975) );
  NAND2_X1 U5666 ( .A1(n5086), .A2(n4985), .ZN(n6659) );
  INV_X1 U5667 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4987) );
  INV_X1 U5668 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6217) );
  INV_X1 U5669 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6072) );
  INV_X1 U5670 ( .A(n8273), .ZN(n4655) );
  OAI21_X1 U5671 ( .B1(n7615), .B2(n7614), .A(n7669), .ZN(n7616) );
  NAND2_X1 U5672 ( .A1(n9126), .A2(n9129), .ZN(n8238) );
  NAND2_X1 U5673 ( .A1(n5768), .A2(n5829), .ZN(n5920) );
  INV_X1 U5674 ( .A(n4863), .ZN(n4860) );
  AOI21_X1 U5675 ( .B1(n5686), .B2(n5862), .A(n9534), .ZN(n4865) );
  NOR2_X1 U5676 ( .A1(n5995), .A2(n4864), .ZN(n4863) );
  INV_X1 U5677 ( .A(n5994), .ZN(n4864) );
  NOR2_X1 U5678 ( .A1(n4848), .A2(n9636), .ZN(n4845) );
  NAND2_X1 U5679 ( .A1(n5543), .A2(n4792), .ZN(n5829) );
  AND2_X1 U5680 ( .A1(n4793), .A2(n5542), .ZN(n4792) );
  INV_X1 U5681 ( .A(n4872), .ZN(n4868) );
  AND2_X1 U5682 ( .A1(n4874), .A2(n5913), .ZN(n4870) );
  NAND2_X1 U5683 ( .A1(n5405), .A2(n4842), .ZN(n4841) );
  NOR2_X1 U5684 ( .A1(n5449), .A2(n5772), .ZN(n4842) );
  NOR2_X1 U5685 ( .A1(n8109), .A2(n7987), .ZN(n4716) );
  NOR2_X1 U5686 ( .A1(n6009), .A2(n9499), .ZN(n5873) );
  AOI21_X1 U5687 ( .B1(n7465), .B2(n5102), .A(n4553), .ZN(n5101) );
  INV_X1 U5688 ( .A(n6019), .ZN(n5102) );
  NAND2_X1 U5689 ( .A1(n5405), .A2(n5900), .ZN(n7540) );
  INV_X1 U5690 ( .A(n5281), .ZN(n5019) );
  NAND2_X1 U5691 ( .A1(n5257), .A2(n5256), .ZN(n5260) );
  INV_X1 U5692 ( .A(SI_19_), .ZN(n5256) );
  INV_X1 U5693 ( .A(n5247), .ZN(n5028) );
  AOI21_X1 U5694 ( .B1(n5027), .B2(n5246), .A(n5025), .ZN(n5024) );
  INV_X1 U5695 ( .A(n5252), .ZN(n5025) );
  INV_X1 U5696 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U5697 ( .A1(n5510), .A2(SI_14_), .ZN(n4764) );
  INV_X1 U5698 ( .A(SI_13_), .ZN(n10481) );
  INV_X1 U5699 ( .A(n4773), .ZN(n4769) );
  OR2_X1 U5700 ( .A1(n5468), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5483) );
  INV_X1 U5701 ( .A(n4752), .ZN(n4751) );
  INV_X1 U5702 ( .A(n5439), .ZN(n4750) );
  NOR2_X2 U5703 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5092) );
  NOR2_X2 U5704 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5364) );
  INV_X1 U5705 ( .A(n5060), .ZN(n5059) );
  OAI21_X1 U5706 ( .B1(n8525), .B2(n5061), .A(n8523), .ZN(n5060) );
  INV_X1 U5707 ( .A(n5064), .ZN(n5061) );
  NOR2_X1 U5708 ( .A1(n8525), .A2(n5063), .ZN(n5062) );
  INV_X1 U5709 ( .A(n8448), .ZN(n5063) );
  NAND2_X1 U5710 ( .A1(n7858), .A2(n7857), .ZN(n7961) );
  NAND2_X1 U5711 ( .A1(n7427), .A2(n5088), .ZN(n7520) );
  AND2_X1 U5712 ( .A1(n7431), .A2(n7426), .ZN(n5088) );
  NAND2_X1 U5713 ( .A1(n8182), .A2(n8181), .ZN(n8195) );
  NAND2_X1 U5714 ( .A1(n8369), .A2(n8511), .ZN(n8514) );
  AND2_X1 U5715 ( .A1(n8388), .A2(n8529), .ZN(n5064) );
  AND4_X1 U5716 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n8466)
         );
  AND4_X1 U5717 ( .A1(n6279), .A2(n6278), .A3(n6277), .A4(n6276), .ZN(n8496)
         );
  OR2_X1 U5718 ( .A1(n10007), .A2(n7305), .ZN(n10005) );
  NAND2_X1 U5719 ( .A1(n4677), .A2(n6813), .ZN(n9991) );
  OAI21_X1 U5720 ( .B1(n6829), .B2(n7015), .A(n6830), .ZN(n7005) );
  NOR2_X1 U5721 ( .A1(n7446), .A2(n7005), .ZN(n7004) );
  AOI21_X1 U5722 ( .B1(n6805), .B2(n7178), .A(n7190), .ZN(n6807) );
  NOR2_X1 U5723 ( .A1(n6807), .A2(n6808), .ZN(n7341) );
  NOR2_X1 U5724 ( .A1(n7361), .A2(n7362), .ZN(n7366) );
  INV_X1 U5725 ( .A(n7358), .ZN(n7359) );
  OR2_X1 U5726 ( .A1(n7366), .A2(n7365), .ZN(n7691) );
  OR2_X1 U5727 ( .A1(n7353), .A2(n7352), .ZN(n7709) );
  AOI21_X1 U5728 ( .B1(n7343), .B2(n7342), .A(n7341), .ZN(n7345) );
  NAND2_X1 U5729 ( .A1(n7345), .A2(n7344), .ZN(n7702) );
  XNOR2_X1 U5730 ( .A(n7712), .B(n7711), .ZN(n10025) );
  NAND2_X1 U5731 ( .A1(n7691), .A2(n7690), .ZN(n7693) );
  OR2_X1 U5732 ( .A1(n10025), .A2(n7796), .ZN(n4729) );
  INV_X1 U5733 ( .A(n7696), .ZN(n4663) );
  AND2_X1 U5734 ( .A1(n6400), .A2(n6399), .ZN(n6403) );
  AOI21_X1 U5735 ( .B1(n7885), .B2(n7884), .A(n7883), .ZN(n7890) );
  NOR2_X1 U5736 ( .A1(n7890), .A2(n7889), .ZN(n8059) );
  NOR2_X1 U5737 ( .A1(n7875), .A2(n7874), .ZN(n7878) );
  NOR2_X1 U5738 ( .A1(n8060), .A2(n8059), .ZN(n8087) );
  NOR2_X1 U5739 ( .A1(n8087), .A2(n8088), .ZN(n8086) );
  NOR2_X1 U5740 ( .A1(n8065), .A2(n8086), .ZN(n8579) );
  NOR2_X1 U5741 ( .A1(n8093), .A2(n8058), .ZN(n8092) );
  AND2_X1 U5742 ( .A1(n4673), .A2(n4672), .ZN(n8598) );
  NAND2_X1 U5743 ( .A1(n8570), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4672) );
  INV_X1 U5744 ( .A(n8567), .ZN(n4673) );
  INV_X1 U5745 ( .A(n8688), .ZN(n4942) );
  NOR2_X1 U5746 ( .A1(n8657), .A2(n4595), .ZN(n8667) );
  NOR2_X1 U5747 ( .A1(n10011), .A2(n8683), .ZN(n4606) );
  INV_X1 U5748 ( .A(n8682), .ZN(n4605) );
  NAND2_X1 U5749 ( .A1(n8681), .A2(n4608), .ZN(n4607) );
  AND2_X1 U5750 ( .A1(n10020), .A2(n8687), .ZN(n4608) );
  NAND2_X1 U5751 ( .A1(n4811), .A2(n4559), .ZN(n4810) );
  OR2_X1 U5752 ( .A1(n6183), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U5753 ( .A1(n6191), .A2(n8431), .ZN(n6193) );
  OR2_X1 U5754 ( .A1(n6235), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U5755 ( .A1(n6233), .A2(n8465), .ZN(n6235) );
  OR2_X1 U5756 ( .A1(n6451), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U5757 ( .A1(n6698), .A2(n6697), .ZN(n8037) );
  AND4_X1 U5758 ( .A1(n6414), .A2(n6413), .A3(n6412), .A4(n6411), .ZN(n8133)
         );
  NAND2_X1 U5759 ( .A1(n6349), .A2(n10394), .ZN(n6422) );
  AND2_X1 U5760 ( .A1(n4797), .A2(n7932), .ZN(n4794) );
  OR2_X1 U5761 ( .A1(n6374), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6376) );
  NOR2_X1 U5762 ( .A1(n6470), .A2(n4950), .ZN(n4949) );
  NAND2_X1 U5763 ( .A1(n7725), .A2(n6689), .ZN(n4824) );
  NAND2_X1 U5764 ( .A1(n6682), .A2(n10032), .ZN(n7441) );
  NAND2_X1 U5765 ( .A1(n6739), .A2(n7217), .ZN(n8927) );
  OR2_X1 U5766 ( .A1(n6792), .A2(n7086), .ZN(n7217) );
  NAND2_X1 U5767 ( .A1(n6628), .A2(n6629), .ZN(n8758) );
  NAND2_X1 U5768 ( .A1(n4815), .A2(n4819), .ZN(n8759) );
  NAND2_X1 U5769 ( .A1(n8787), .A2(n4821), .ZN(n4815) );
  INV_X1 U5770 ( .A(n8758), .ZN(n8756) );
  NAND2_X1 U5771 ( .A1(n8850), .A2(n8849), .ZN(n8848) );
  AND2_X1 U5772 ( .A1(n6574), .A2(n6580), .ZN(n8883) );
  INV_X1 U5773 ( .A(n8883), .ZN(n8881) );
  AND2_X1 U5774 ( .A1(n7113), .A2(n6741), .ZN(n8911) );
  AND3_X1 U5775 ( .A1(n6336), .A2(n6335), .A3(n6334), .ZN(n10044) );
  AND2_X1 U5776 ( .A1(n7105), .A2(n6880), .ZN(n7111) );
  NAND2_X1 U5777 ( .A1(n8927), .A2(n6746), .ZN(n10078) );
  XNOR2_X1 U5778 ( .A(n6661), .B(n6660), .ZN(n6793) );
  INV_X1 U5779 ( .A(n9102), .ZN(n6880) );
  INV_X1 U5780 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6078) );
  OR2_X1 U5781 ( .A1(n6432), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6243) );
  INV_X1 U5782 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6358) );
  OR2_X1 U5783 ( .A1(n6287), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6381) );
  INV_X1 U5784 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6332) );
  INV_X1 U5785 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6296) );
  XNOR2_X1 U5786 ( .A(n6305), .B(n6304), .ZN(n6823) );
  NAND2_X1 U5787 ( .A1(n4943), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U5788 ( .A1(n7671), .A2(n7621), .ZN(n7622) );
  NAND2_X1 U5789 ( .A1(n7622), .A2(n7623), .ZN(n7995) );
  NAND2_X1 U5790 ( .A1(n9529), .A2(n9920), .ZN(n4627) );
  NAND2_X1 U5791 ( .A1(n4630), .A2(n8232), .ZN(n9126) );
  INV_X1 U5792 ( .A(n8232), .ZN(n4628) );
  INV_X1 U5793 ( .A(n4630), .ZN(n4629) );
  NAND2_X1 U5794 ( .A1(n9241), .A2(n9242), .ZN(n4915) );
  AND2_X1 U5795 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  NAND2_X1 U5796 ( .A1(n5678), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5680) );
  AND2_X1 U5797 ( .A1(n7577), .A2(n7576), .ZN(n7619) );
  NOR2_X1 U5798 ( .A1(n5643), .A2(n9138), .ZN(n5634) );
  AND2_X1 U5799 ( .A1(n8292), .A2(n8291), .ZN(n9216) );
  AND2_X1 U5800 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5373) );
  OAI21_X1 U5801 ( .B1(n9896), .B2(n4886), .A(n4880), .ZN(n9233) );
  INV_X1 U5802 ( .A(n4881), .ZN(n4880) );
  AOI21_X1 U5803 ( .B1(n4635), .B2(n4882), .A(n4528), .ZN(n4881) );
  NOR2_X1 U5804 ( .A1(n4884), .A2(n9175), .ZN(n4882) );
  NAND2_X1 U5805 ( .A1(n9233), .A2(n9234), .ZN(n9232) );
  OR2_X1 U5806 ( .A1(n5680), .A2(n9168), .ZN(n5666) );
  NAND2_X1 U5807 ( .A1(n9896), .A2(n4635), .ZN(n4634) );
  INV_X1 U5808 ( .A(n8121), .ZN(n4633) );
  NAND2_X1 U5809 ( .A1(n7251), .A2(n7252), .ZN(n4618) );
  OR2_X1 U5810 ( .A1(n5560), .A2(n5559), .ZN(n5573) );
  AND2_X1 U5811 ( .A1(n7126), .A2(n9866), .ZN(n7147) );
  OR3_X1 U5812 ( .A1(n5517), .A2(n5516), .A3(n9130), .ZN(n5529) );
  AOI21_X1 U5813 ( .B1(n9127), .B2(n8238), .A(n8237), .ZN(n9273) );
  AND4_X1 U5814 ( .A1(n5565), .A2(n5564), .A3(n5563), .A4(n5562), .ZN(n9256)
         );
  AND4_X1 U5815 ( .A1(n5431), .A2(n5430), .A3(n5429), .A4(n5428), .ZN(n7999)
         );
  NAND2_X1 U5816 ( .A1(n9478), .A2(n9828), .ZN(n9477) );
  AND2_X1 U5817 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5692), .ZN(n5602) );
  NOR2_X1 U5818 ( .A1(n9527), .A2(n5124), .ZN(n5119) );
  NOR2_X1 U5819 ( .A1(n5693), .A2(n9266), .ZN(n5692) );
  OR2_X1 U5820 ( .A1(n5862), .A2(n5995), .ZN(n9548) );
  NAND2_X1 U5821 ( .A1(n5126), .A2(n5125), .ZN(n9564) );
  NAND2_X1 U5822 ( .A1(n4564), .A2(n6039), .ZN(n5125) );
  AND2_X1 U5823 ( .A1(n5629), .A2(n5628), .ZN(n9585) );
  NAND2_X1 U5824 ( .A1(n9599), .A2(n9605), .ZN(n9600) );
  NAND2_X1 U5825 ( .A1(n9675), .A2(n4546), .ZN(n5596) );
  INV_X1 U5826 ( .A(n9657), .ZN(n4843) );
  NOR2_X1 U5827 ( .A1(n5573), .A2(n9255), .ZN(n5590) );
  AND2_X1 U5828 ( .A1(n4519), .A2(n9674), .ZN(n4717) );
  AND2_X1 U5829 ( .A1(n5832), .A2(n5834), .ZN(n9676) );
  NAND2_X1 U5830 ( .A1(n9706), .A2(n5149), .ZN(n9688) );
  OR2_X1 U5831 ( .A1(n9710), .A2(n9278), .ZN(n5149) );
  INV_X1 U5832 ( .A(n9682), .ZN(n5566) );
  NOR2_X1 U5833 ( .A1(n5529), .A2(n9277), .ZN(n5544) );
  NAND2_X1 U5834 ( .A1(n8154), .A2(n9865), .ZN(n9731) );
  NAND2_X1 U5835 ( .A1(n8154), .A2(n4718), .ZN(n9708) );
  OAI21_X1 U5836 ( .B1(n7907), .B2(n4869), .A(n4866), .ZN(n9722) );
  INV_X1 U5837 ( .A(n4870), .ZN(n4869) );
  AOI21_X1 U5838 ( .B1(n4870), .B2(n4868), .A(n4867), .ZN(n4866) );
  INV_X1 U5839 ( .A(n5817), .ZN(n4867) );
  AND2_X1 U5840 ( .A1(n5768), .A2(n5821), .ZN(n9723) );
  AND2_X1 U5841 ( .A1(n7777), .A2(n4575), .ZN(n8155) );
  NAND2_X1 U5842 ( .A1(n4871), .A2(n5913), .ZN(n8148) );
  NAND2_X1 U5843 ( .A1(n4871), .A2(n4870), .ZN(n8150) );
  NAND2_X1 U5844 ( .A1(n7907), .A2(n5910), .ZN(n8016) );
  NAND2_X1 U5845 ( .A1(n7777), .A2(n4523), .ZN(n7941) );
  NAND2_X1 U5846 ( .A1(n4841), .A2(n5903), .ZN(n7769) );
  AOI21_X1 U5847 ( .B1(n7642), .B2(n5111), .A(n4560), .ZN(n5110) );
  NAND2_X1 U5848 ( .A1(n7774), .A2(n7776), .ZN(n7775) );
  NAND2_X1 U5849 ( .A1(n7777), .A2(n4716), .ZN(n7943) );
  OR2_X1 U5850 ( .A1(n5434), .A2(n5416), .ZN(n5459) );
  AND2_X1 U5851 ( .A1(n7545), .A2(n7764), .ZN(n7777) );
  NOR2_X1 U5852 ( .A1(n7470), .A2(n7469), .ZN(n7546) );
  NAND2_X1 U5853 ( .A1(n4705), .A2(n7584), .ZN(n7470) );
  INV_X1 U5854 ( .A(n7412), .ZN(n4705) );
  NAND2_X1 U5855 ( .A1(n4706), .A2(n9957), .ZN(n7412) );
  NAND2_X1 U5856 ( .A1(n7410), .A2(n7409), .ZN(n7408) );
  NAND2_X1 U5857 ( .A1(n4836), .A2(n4835), .ZN(n7404) );
  AOI21_X1 U5858 ( .B1(n5893), .B2(n4837), .A(n4561), .ZN(n4835) );
  INV_X1 U5859 ( .A(n5091), .ZN(n4837) );
  NAND2_X1 U5860 ( .A1(n4838), .A2(n5091), .ZN(n7227) );
  INV_X1 U5861 ( .A(n7155), .ZN(n4838) );
  NAND2_X1 U5862 ( .A1(n7152), .A2(n7154), .ZN(n7151) );
  CLKBUF_X1 U5863 ( .A(n6013), .Z(n7022) );
  NOR2_X1 U5864 ( .A1(n7038), .A2(n9888), .ZN(n7023) );
  INV_X1 U5865 ( .A(n6006), .ZN(n4850) );
  INV_X1 U5866 ( .A(n9969), .ZN(n9813) );
  OR2_X1 U5867 ( .A1(n6056), .A2(n7140), .ZN(n7758) );
  NOR2_X1 U5868 ( .A1(n5160), .A2(n4539), .ZN(n5339) );
  NAND2_X1 U5869 ( .A1(n7923), .A2(n7811), .ZN(n7175) );
  XNOR2_X1 U5870 ( .A(n5295), .B(n5296), .ZN(n5703) );
  NAND2_X1 U5871 ( .A1(n5141), .A2(n5174), .ZN(n5140) );
  INV_X1 U5872 ( .A(n4995), .ZN(n5597) );
  AOI21_X1 U5873 ( .B1(n5610), .B2(n5611), .A(n4998), .ZN(n4995) );
  XNOR2_X1 U5874 ( .A(n5610), .B(n5611), .ZN(n9113) );
  NAND2_X1 U5875 ( .A1(n5734), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5737) );
  INV_X1 U5876 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5584) );
  INV_X1 U5877 ( .A(n4640), .ZN(n4639) );
  NAND2_X1 U5878 ( .A1(n4638), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U5879 ( .A1(n5555), .A2(n4534), .ZN(n4638) );
  NAND2_X1 U5880 ( .A1(n5494), .A2(n5244), .ZN(n5497) );
  NAND2_X1 U5881 ( .A1(n4772), .A2(n4771), .ZN(n5482) );
  NAND2_X1 U5882 ( .A1(n4772), .A2(n5238), .ZN(n5480) );
  NAND2_X1 U5883 ( .A1(n5453), .A2(n5234), .ZN(n5467) );
  CLKBUF_X1 U5884 ( .A(n5408), .Z(n5409) );
  INV_X1 U5885 ( .A(n5344), .ZN(n4989) );
  INV_X1 U5886 ( .A(n5202), .ZN(n4990) );
  AND2_X1 U5887 ( .A1(n5210), .A2(n5211), .ZN(n5360) );
  CLKBUF_X1 U5888 ( .A(n5315), .Z(n5334) );
  NAND2_X1 U5889 ( .A1(n5053), .A2(n5059), .ZN(n8420) );
  NAND2_X1 U5890 ( .A1(n8447), .A2(n5062), .ZN(n5053) );
  NAND2_X1 U5891 ( .A1(n8357), .A2(n8493), .ZN(n8397) );
  AND4_X1 U5892 ( .A1(n6398), .A2(n6397), .A3(n6396), .A4(n6395), .ZN(n8191)
         );
  NAND2_X1 U5893 ( .A1(n8514), .A2(n8371), .ZN(n8410) );
  AND2_X1 U5894 ( .A1(n6118), .A2(n6117), .ZN(n8555) );
  AOI21_X1 U5895 ( .B1(n8473), .B2(n5051), .A(n5048), .ZN(n5047) );
  OAI21_X1 U5896 ( .B1(n5050), .B2(n5049), .A(n5054), .ZN(n5048) );
  INV_X1 U5897 ( .A(n8387), .ZN(n5049) );
  AND2_X1 U5898 ( .A1(n6171), .A2(n6170), .ZN(n8475) );
  AND2_X1 U5899 ( .A1(n6262), .A2(n6261), .ZN(n8461) );
  AND4_X1 U5900 ( .A1(n6239), .A2(n6238), .A3(n6237), .A4(n6236), .ZN(n8855)
         );
  NAND2_X1 U5901 ( .A1(n8456), .A2(n8455), .ZN(n8454) );
  NAND2_X1 U5902 ( .A1(n8454), .A2(n8366), .ZN(n8463) );
  AND2_X1 U5903 ( .A1(n7427), .A2(n7426), .ZN(n7432) );
  NAND2_X1 U5904 ( .A1(n8138), .A2(n8137), .ZN(n8141) );
  NAND2_X1 U5905 ( .A1(n5040), .A2(n5043), .ZN(n8485) );
  AND2_X1 U5906 ( .A1(n5044), .A2(n8374), .ZN(n5043) );
  NAND2_X1 U5907 ( .A1(n8369), .A2(n5041), .ZN(n5040) );
  NAND2_X1 U5908 ( .A1(n6181), .A2(n6180), .ZN(n8507) );
  AND2_X1 U5909 ( .A1(n8201), .A2(n8347), .ZN(n5070) );
  NAND2_X1 U5910 ( .A1(n8184), .A2(n8183), .ZN(n8200) );
  AND4_X1 U5911 ( .A1(n6366), .A2(n6365), .A3(n6364), .A4(n6363), .ZN(n7854)
         );
  AND2_X1 U5912 ( .A1(n7596), .A2(n7592), .ZN(n5087) );
  NAND2_X1 U5913 ( .A1(n7593), .A2(n7592), .ZN(n7594) );
  AOI21_X1 U5914 ( .B1(n8447), .B2(n8448), .A(n5064), .ZN(n8527) );
  NAND2_X1 U5915 ( .A1(n7285), .A2(n7928), .ZN(n8533) );
  AND2_X1 U5916 ( .A1(n6657), .A2(n6778), .ZN(n4703) );
  NAND2_X1 U5917 ( .A1(n6143), .A2(n6142), .ZN(n8736) );
  INV_X1 U5918 ( .A(n8389), .ZN(n8760) );
  INV_X1 U5919 ( .A(n8529), .ZN(n8777) );
  INV_X1 U5920 ( .A(n8475), .ZN(n8789) );
  INV_X1 U5921 ( .A(n8809), .ZN(n8788) );
  INV_X1 U5922 ( .A(n8798), .ZN(n8831) );
  INV_X1 U5923 ( .A(n8855), .ZN(n8874) );
  INV_X1 U5924 ( .A(n8399), .ZN(n8897) );
  INV_X1 U5925 ( .A(n8496), .ZN(n8910) );
  INV_X1 U5926 ( .A(n7854), .ZN(n8560) );
  AND2_X1 U5927 ( .A1(n6329), .A2(n5161), .ZN(n6330) );
  OR2_X1 U5928 ( .A1(n6821), .A2(n6797), .ZN(n8680) );
  NOR2_X1 U5929 ( .A1(n6981), .A2(n6982), .ZN(n6980) );
  NAND2_X1 U5930 ( .A1(n4669), .A2(n6815), .ZN(n7009) );
  INV_X1 U5931 ( .A(n4668), .ZN(n7008) );
  NOR2_X1 U5932 ( .A1(n7191), .A2(n7192), .ZN(n7190) );
  INV_X1 U5933 ( .A(n10014), .ZN(n8679) );
  XNOR2_X1 U5934 ( .A(n4933), .B(n7814), .ZN(n7813) );
  NOR2_X1 U5935 ( .A1(n7813), .A2(n6407), .ZN(n7867) );
  OAI21_X1 U5936 ( .B1(n7813), .B2(n4935), .A(n4934), .ZN(n8071) );
  NAND2_X1 U5937 ( .A1(n4936), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U5938 ( .A1(n7868), .A2(n4936), .ZN(n4934) );
  INV_X1 U5939 ( .A(n7870), .ZN(n4936) );
  INV_X1 U5940 ( .A(n8074), .ZN(n4924) );
  OAI21_X1 U5941 ( .B1(n8093), .B2(n4722), .A(n4721), .ZN(n8569) );
  NAND2_X1 U5942 ( .A1(n8055), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U5943 ( .A1(n8053), .A2(n8055), .ZN(n4721) );
  NOR2_X1 U5944 ( .A1(n8572), .A2(n8571), .ZN(n8587) );
  NAND2_X1 U5945 ( .A1(n4928), .A2(n4927), .ZN(n8620) );
  NAND2_X1 U5946 ( .A1(n4737), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4736) );
  NAND2_X1 U5947 ( .A1(n8588), .A2(n4737), .ZN(n4735) );
  INV_X1 U5948 ( .A(n8589), .ZN(n4737) );
  INV_X1 U5949 ( .A(n8630), .ZN(n4732) );
  OAI21_X1 U5950 ( .B1(n8611), .B2(n4731), .A(n4730), .ZN(n8657) );
  NAND2_X1 U5951 ( .A1(n4734), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U5952 ( .A1(n8630), .A2(n4734), .ZN(n4730) );
  INV_X1 U5953 ( .A(n8632), .ZN(n4734) );
  NAND2_X1 U5954 ( .A1(n6480), .A2(n6612), .ZN(n8800) );
  NAND2_X1 U5955 ( .A1(n8827), .A2(n6717), .ZN(n8807) );
  NAND2_X1 U5956 ( .A1(n6222), .A2(n6221), .ZN(n8988) );
  NAND2_X1 U5957 ( .A1(n7215), .A2(n8938), .ZN(n8820) );
  NAND2_X1 U5958 ( .A1(n4962), .A2(n4963), .ZN(n8028) );
  NAND2_X1 U5959 ( .A1(n4967), .A2(n6541), .ZN(n7931) );
  NAND2_X1 U5960 ( .A1(n4968), .A2(n6545), .ZN(n4967) );
  AOI22_X1 U5961 ( .A1(n6446), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7698), .B2(
        n6445), .ZN(n4701) );
  NAND2_X1 U5962 ( .A1(n6862), .A2(n6431), .ZN(n4702) );
  OR2_X1 U5963 ( .A1(n6860), .A2(n6346), .ZN(n6371) );
  NAND2_X1 U5964 ( .A1(n7498), .A2(n6519), .ZN(n7723) );
  INV_X1 U5965 ( .A(n8820), .ZN(n8890) );
  OR2_X1 U5966 ( .A1(n8958), .A2(n8957), .ZN(n9020) );
  NAND2_X1 U5967 ( .A1(n6145), .A2(n6144), .ZN(n9023) );
  NAND2_X1 U5968 ( .A1(n4960), .A2(n6628), .ZN(n8746) );
  NAND2_X1 U5969 ( .A1(n6154), .A2(n6153), .ZN(n9029) );
  NAND2_X1 U5970 ( .A1(n6164), .A2(n6163), .ZN(n9035) );
  XOR2_X1 U5971 ( .A(n8775), .B(n8773), .Z(n9038) );
  INV_X1 U5972 ( .A(n8507), .ZN(n9048) );
  NAND2_X1 U5973 ( .A1(n6198), .A2(n6197), .ZN(n9056) );
  NAND2_X1 U5974 ( .A1(n8837), .A2(n6603), .ZN(n8824) );
  NAND2_X1 U5975 ( .A1(n6210), .A2(n6209), .ZN(n9062) );
  NAND2_X1 U5976 ( .A1(n6232), .A2(n6231), .ZN(n9072) );
  NAND2_X1 U5977 ( .A1(n4952), .A2(n6582), .ZN(n8861) );
  NAND2_X1 U5978 ( .A1(n6477), .A2(n4956), .ZN(n4952) );
  INV_X1 U5979 ( .A(n8461), .ZN(n9078) );
  NAND2_X1 U5980 ( .A1(n6477), .A2(n6574), .ZN(n8871) );
  NAND2_X1 U5981 ( .A1(n6250), .A2(n6249), .ZN(n9084) );
  NAND2_X1 U5982 ( .A1(n6272), .A2(n6271), .ZN(n9090) );
  OAI21_X1 U5983 ( .B1(n8172), .B2(n4521), .A(n4972), .ZN(n8893) );
  INV_X1 U5984 ( .A(n9052), .ZN(n9096) );
  NAND2_X1 U5985 ( .A1(n8170), .A2(n6473), .ZN(n8906) );
  AND3_X1 U5986 ( .A1(n6386), .A2(n6385), .A3(n6384), .ZN(n7754) );
  OR2_X1 U5987 ( .A1(n10087), .A2(n10073), .ZN(n9052) );
  AND2_X1 U5988 ( .A1(n6755), .A2(n6754), .ZN(n9103) );
  AND2_X1 U5989 ( .A1(n6793), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7109) );
  XNOR2_X1 U5990 ( .A(n6666), .B(n6080), .ZN(n9120) );
  CLKBUF_X1 U5991 ( .A(n6664), .Z(n6665) );
  OR2_X1 U5992 ( .A1(n6668), .A2(n6667), .ZN(n6670) );
  INV_X1 U5993 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7921) );
  INV_X1 U5994 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7532) );
  INV_X1 U5995 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7299) );
  INV_X1 U5996 ( .A(n8644), .ZN(n8658) );
  INV_X1 U5997 ( .A(n10013), .ZN(n7711) );
  INV_X1 U5998 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U5999 ( .A1(n4676), .A2(n4675), .ZN(n4674) );
  INV_X1 U6000 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4675) );
  AND2_X1 U6001 ( .A1(n7239), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6790) );
  INV_X1 U6002 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U6003 ( .A1(n5515), .A2(n5514), .ZN(n9134) );
  INV_X1 U6004 ( .A(n9843), .ZN(n9590) );
  INV_X1 U6005 ( .A(n9652), .ZN(n9798) );
  OR2_X1 U6006 ( .A1(n9162), .A2(n4897), .ZN(n4896) );
  OR2_X1 U6007 ( .A1(n9161), .A2(n9916), .ZN(n4897) );
  AND2_X1 U6008 ( .A1(n8318), .A2(n4893), .ZN(n4891) );
  AND2_X1 U6009 ( .A1(n9162), .A2(n9906), .ZN(n4893) );
  OR2_X1 U6010 ( .A1(n8318), .A2(n4896), .ZN(n4889) );
  NOR2_X1 U6011 ( .A1(n4580), .A2(n4895), .ZN(n4894) );
  INV_X1 U6012 ( .A(n9163), .ZN(n4895) );
  OAI21_X1 U6013 ( .B1(n4883), .B2(n4888), .A(n4885), .ZN(n9173) );
  NAND2_X1 U6014 ( .A1(n4635), .A2(n8216), .ZN(n4888) );
  NAND2_X1 U6015 ( .A1(n5543), .A2(n5542), .ZN(n9812) );
  NOR3_X1 U6016 ( .A1(n4520), .A2(n4909), .A3(n9216), .ZN(n9217) );
  OR2_X1 U6017 ( .A1(n8275), .A2(n4653), .ZN(n4645) );
  NOR2_X1 U6018 ( .A1(n4533), .A2(n4644), .ZN(n4643) );
  INV_X1 U6019 ( .A(n7041), .ZN(n9888) );
  INV_X1 U6020 ( .A(n9143), .ZN(n4877) );
  OR2_X1 U6021 ( .A1(n8275), .A2(n8274), .ZN(n4651) );
  AND4_X1 U6022 ( .A1(n5464), .A2(n5463), .A3(n5462), .A4(n5461), .ZN(n8123)
         );
  NOR2_X1 U6023 ( .A1(n4634), .A2(n4633), .ZN(n8122) );
  INV_X1 U6024 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9255) );
  AND2_X1 U6025 ( .A1(n7147), .A2(n7146), .ZN(n9900) );
  INV_X1 U6026 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U6027 ( .A1(n7243), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9923) );
  NAND2_X1 U6028 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  NOR2_X1 U6029 ( .A1(n5948), .A2(n5947), .ZN(n5955) );
  INV_X1 U6030 ( .A(n5944), .ZN(n5948) );
  INV_X1 U6031 ( .A(n7923), .ZN(n6053) );
  INV_X1 U6032 ( .A(n9585), .ZN(n9289) );
  INV_X1 U6033 ( .A(n9256), .ZN(n9702) );
  AOI22_X1 U6034 ( .A1(n5708), .A2(P1_REG1_REG_1__SCAN_IN), .B1(n5707), .B2(
        P1_REG0_REG_1__SCAN_IN), .ZN(n4832) );
  INV_X1 U6035 ( .A(P1_U3973), .ZN(n9306) );
  AND2_X1 U6036 ( .A1(n9441), .A2(n9440), .ZN(n9447) );
  OR2_X1 U6037 ( .A1(n9437), .A2(n9436), .ZN(n9456) );
  INV_X1 U6038 ( .A(n9478), .ZN(n6008) );
  NAND2_X1 U6039 ( .A1(n4855), .A2(n6006), .ZN(n9493) );
  AOI21_X1 U6040 ( .B1(n9502), .B2(n9724), .A(n9501), .ZN(n9754) );
  OAI21_X1 U6041 ( .B1(n9537), .B2(n9662), .A(n9500), .ZN(n9501) );
  NAND2_X1 U6042 ( .A1(n9497), .A2(n5157), .ZN(n9502) );
  NOR2_X1 U6043 ( .A1(n9522), .A2(n9521), .ZN(n9523) );
  AND2_X1 U6044 ( .A1(n9517), .A2(n9516), .ZN(n9757) );
  NAND2_X1 U6045 ( .A1(n5120), .A2(n5123), .ZN(n9528) );
  INV_X1 U6046 ( .A(n9763), .ZN(n9544) );
  AOI21_X1 U6047 ( .B1(n9550), .B2(n5996), .A(n5995), .ZN(n9535) );
  NAND2_X1 U6048 ( .A1(n6045), .A2(n6044), .ZN(n9533) );
  AND2_X1 U6049 ( .A1(n5622), .A2(n5621), .ZN(n9576) );
  NAND2_X1 U6050 ( .A1(n5129), .A2(n5131), .ZN(n9579) );
  NAND2_X1 U6051 ( .A1(n9616), .A2(n5134), .ZN(n5129) );
  NAND2_X1 U6052 ( .A1(n9619), .A2(n5989), .ZN(n9608) );
  NAND2_X1 U6053 ( .A1(n5130), .A2(n5136), .ZN(n9598) );
  OR2_X1 U6054 ( .A1(n9616), .A2(n6036), .ZN(n5130) );
  NAND2_X1 U6055 ( .A1(n5114), .A2(n6033), .ZN(n9634) );
  NAND2_X1 U6056 ( .A1(n9675), .A2(n5834), .ZN(n9658) );
  NAND2_X1 U6057 ( .A1(n5115), .A2(n5118), .ZN(n9650) );
  OR2_X1 U6058 ( .A1(n9667), .A2(n6032), .ZN(n5115) );
  AND2_X1 U6059 ( .A1(n5094), .A2(n5097), .ZN(n8146) );
  NAND2_X1 U6060 ( .A1(n6027), .A2(n6026), .ZN(n8013) );
  INV_X1 U6061 ( .A(n9642), .ZN(n9945) );
  NAND2_X1 U6062 ( .A1(n7643), .A2(n7642), .ZN(n7641) );
  NAND2_X1 U6063 ( .A1(n7654), .A2(n6020), .ZN(n7643) );
  NOR2_X1 U6064 ( .A1(n9612), .A2(n7394), .ZN(n9642) );
  NAND2_X1 U6065 ( .A1(n7463), .A2(n7465), .ZN(n7462) );
  NAND2_X1 U6066 ( .A1(n7376), .A2(n6019), .ZN(n7463) );
  INV_X1 U6067 ( .A(n9741), .ZN(n9707) );
  NAND2_X1 U6068 ( .A1(n9866), .A2(n7129), .ZN(n9711) );
  AND2_X1 U6069 ( .A1(n5651), .A2(n5650), .ZN(n9838) );
  INV_X1 U6070 ( .A(n9643), .ZN(n9852) );
  NAND2_X1 U6071 ( .A1(n6871), .A2(n4710), .ZN(n4709) );
  NAND2_X1 U6072 ( .A1(n5586), .A2(n9309), .ZN(n4834) );
  OAI22_X1 U6073 ( .A1(n6853), .A2(n6318), .B1(n6842), .B2(n6847), .ZN(n4710)
         );
  NAND2_X1 U6074 ( .A1(n9860), .A2(n9956), .ZN(n9864) );
  AND2_X1 U6075 ( .A1(n7240), .A2(n6790), .ZN(n9866) );
  XNOR2_X1 U6076 ( .A(n5725), .B(n5724), .ZN(n6066) );
  OAI22_X1 U6077 ( .A1(n5721), .A2(n5720), .B1(SI_30_), .B2(n5719), .ZN(n5725)
         );
  OAI21_X1 U6078 ( .B1(n5703), .B2(SI_29_), .A(n5704), .ZN(n9876) );
  INV_X1 U6079 ( .A(n5973), .ZN(n9881) );
  NAND2_X1 U6080 ( .A1(n4905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U6081 ( .A1(n5733), .A2(n4535), .ZN(n4905) );
  INV_X1 U6082 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U6083 ( .A1(n5002), .A2(n5007), .ZN(n5631) );
  NAND2_X1 U6084 ( .A1(n5662), .A2(n5011), .ZN(n5002) );
  INV_X1 U6085 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10278) );
  INV_X1 U6086 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7633) );
  NAND2_X1 U6087 ( .A1(n5555), .A2(n5554), .ZN(n5569) );
  NAND2_X1 U6088 ( .A1(n5030), .A2(n5231), .ZN(n5451) );
  NAND2_X1 U6089 ( .A1(n5345), .A2(n5344), .ZN(n5347) );
  NAND2_X1 U6090 ( .A1(n5332), .A2(n5197), .ZN(n5345) );
  AND2_X1 U6091 ( .A1(n7290), .A2(n7289), .ZN(n7292) );
  NAND2_X1 U6092 ( .A1(n5081), .A2(n7201), .ZN(n7096) );
  NOR2_X1 U6093 ( .A1(n4594), .A2(n7694), .ZN(n7697) );
  INV_X1 U6094 ( .A(n4925), .ZN(n8084) );
  INV_X1 U6095 ( .A(n4733), .ZN(n8629) );
  INV_X1 U6096 ( .A(n4670), .ZN(n8686) );
  OAI21_X1 U6097 ( .B1(n8690), .B2(n10026), .A(n4602), .ZN(P2_U3200) );
  NOR2_X1 U6098 ( .A1(n4937), .A2(n4603), .ZN(n4602) );
  AND2_X1 U6099 ( .A1(n4939), .A2(n9997), .ZN(n4603) );
  AOI21_X1 U6100 ( .B1(n4658), .B2(n9997), .A(n8709), .ZN(n8710) );
  OAI21_X1 U6101 ( .B1(n4806), .B2(n8920), .A(n4804), .ZN(P2_U3204) );
  INV_X1 U6102 ( .A(n4805), .ZN(n4804) );
  NOR2_X1 U6103 ( .A1(n6773), .A2(n6775), .ZN(n6776) );
  NOR2_X1 U6104 ( .A1(n8324), .A2(n8980), .ZN(n6773) );
  NAND2_X1 U6105 ( .A1(n8952), .A2(n8951), .ZN(n8954) );
  OAI21_X1 U6106 ( .B1(n9186), .B2(n4530), .A(n4624), .ZN(n4625) );
  AOI21_X1 U6107 ( .B1(n9263), .B2(n4524), .A(n4621), .ZN(n4620) );
  NOR2_X1 U6108 ( .A1(n4626), .A2(n9916), .ZN(n4624) );
  OAI21_X1 U6109 ( .B1(n9743), .B2(n9985), .A(n4711), .ZN(P1_U3553) );
  AOI21_X1 U6110 ( .B1(n5732), .B2(n7806), .A(n4712), .ZN(n4711) );
  NOR2_X1 U6111 ( .A1(n9988), .A2(n9744), .ZN(n4712) );
  OR2_X1 U6112 ( .A1(n4852), .A2(n9985), .ZN(n4851) );
  INV_X1 U6113 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n4853) );
  AND2_X1 U6114 ( .A1(n4718), .A2(n9858), .ZN(n4519) );
  OAI21_X1 U6115 ( .B1(n8301), .B2(n4530), .A(n8317), .ZN(n4626) );
  INV_X2 U6116 ( .A(n6339), .ZN(n6300) );
  AND2_X1 U6117 ( .A1(n4916), .A2(n4913), .ZN(n4520) );
  OR2_X1 U6118 ( .A1(n6474), .A2(n6559), .ZN(n4521) );
  OR2_X1 U6119 ( .A1(n9773), .A2(n9585), .ZN(n5992) );
  XOR2_X1 U6120 ( .A(n6000), .B(n5999), .Z(n4522) );
  INV_X1 U6121 ( .A(n4653), .ZN(n4652) );
  OAI21_X1 U6122 ( .B1(n4914), .B2(n4654), .A(n4908), .ZN(n4653) );
  AND2_X1 U6123 ( .A1(n4716), .A2(n4715), .ZN(n4523) );
  INV_X1 U6124 ( .A(n7379), .ZN(n5100) );
  AND2_X1 U6125 ( .A1(n8318), .A2(n9906), .ZN(n4524) );
  AND3_X1 U6126 ( .A1(n4927), .A2(n4928), .A3(n4590), .ZN(n4525) );
  AND2_X1 U6127 ( .A1(n5026), .A2(n4579), .ZN(n4526) );
  AND4_X1 U6128 ( .A1(n5670), .A2(n5669), .A3(n5668), .A4(n5667), .ZN(n9246)
         );
  AND2_X1 U6129 ( .A1(n6813), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4527) );
  INV_X1 U6130 ( .A(n4862), .ZN(n4861) );
  OAI21_X1 U6131 ( .B1(n5995), .B2(n5992), .A(n4865), .ZN(n4862) );
  INV_X1 U6132 ( .A(n9957), .ZN(n7414) );
  AND3_X1 U6133 ( .A1(n5370), .A2(n5369), .A3(n5368), .ZN(n9957) );
  INV_X1 U6134 ( .A(n8227), .ZN(n4884) );
  AND2_X1 U6135 ( .A1(n4886), .A2(n8227), .ZN(n4528) );
  OR2_X1 U6136 ( .A1(n9734), .A2(n9701), .ZN(n4529) );
  AND2_X1 U6137 ( .A1(n5571), .A2(n5570), .ZN(n9674) );
  INV_X1 U6138 ( .A(n9674), .ZN(n4719) );
  AND2_X1 U6139 ( .A1(n8305), .A2(n8304), .ZN(n4530) );
  AND2_X1 U6140 ( .A1(n5730), .A2(n5729), .ZN(n9745) );
  INV_X1 U6141 ( .A(n9745), .ZN(n5732) );
  INV_X1 U6142 ( .A(n9529), .ZN(n9833) );
  NAND2_X1 U6143 ( .A1(n5613), .A2(n5612), .ZN(n9529) );
  XNOR2_X1 U6144 ( .A(n6663), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6750) );
  NAND3_X1 U6145 ( .A1(n8332), .A2(n4618), .A3(n4619), .ZN(n8331) );
  INV_X1 U6146 ( .A(n9607), .ZN(n4744) );
  AND2_X1 U6147 ( .A1(n7988), .A2(n9914), .ZN(n4531) );
  AND2_X1 U6148 ( .A1(n5086), .A2(n4986), .ZN(n6490) );
  OR2_X1 U6149 ( .A1(n7260), .A2(n7259), .ZN(n4532) );
  NAND3_X1 U6150 ( .A1(n7994), .A2(n7996), .A3(n7993), .ZN(n4533) );
  AND2_X1 U6151 ( .A1(n6541), .A2(n6545), .ZN(n7897) );
  AND2_X1 U6152 ( .A1(n5554), .A2(n5556), .ZN(n4534) );
  AND2_X1 U6153 ( .A1(n5170), .A2(n5960), .ZN(n4535) );
  INV_X1 U6154 ( .A(n4914), .ZN(n4913) );
  NAND2_X1 U6155 ( .A1(n4917), .A2(n4915), .ZN(n4914) );
  NAND2_X1 U6156 ( .A1(n6331), .A2(n6330), .ZN(n6526) );
  OR2_X1 U6157 ( .A1(n8685), .A2(n8684), .ZN(n4536) );
  XNOR2_X1 U6158 ( .A(n9016), .B(n8736), .ZN(n8718) );
  OR2_X1 U6159 ( .A1(n9241), .A2(n9242), .ZN(n4537) );
  OAI21_X1 U6160 ( .B1(n8787), .B2(n6721), .A(n6720), .ZN(n8774) );
  INV_X1 U6161 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4641) );
  NAND2_X1 U6162 ( .A1(n4812), .A2(n4810), .ZN(n8733) );
  NAND2_X1 U6163 ( .A1(n4803), .A2(n6713), .ZN(n8851) );
  AND2_X1 U6164 ( .A1(n5304), .A2(n5303), .ZN(n9828) );
  NAND2_X1 U6165 ( .A1(n6487), .A2(n6486), .ZN(n6732) );
  INV_X1 U6166 ( .A(n5989), .ZN(n4848) );
  NAND2_X1 U6167 ( .A1(n5528), .A2(n5527), .ZN(n9734) );
  INV_X1 U6168 ( .A(n6557), .ZN(n4691) );
  OR2_X1 U6169 ( .A1(n9008), .A2(n8553), .ZN(n4538) );
  NAND2_X1 U6170 ( .A1(n5471), .A2(n5470), .ZN(n8115) );
  INV_X1 U6171 ( .A(n8115), .ZN(n4715) );
  NAND2_X1 U6172 ( .A1(n6670), .A2(n6669), .ZN(n6749) );
  AND3_X1 U6173 ( .A1(n5966), .A2(n7070), .A3(n9927), .ZN(n4539) );
  AND3_X1 U6174 ( .A1(n5831), .A2(n5834), .A3(n5925), .ZN(n4540) );
  AND3_X1 U6175 ( .A1(n5512), .A2(n5105), .A3(n5170), .ZN(n5958) );
  AND2_X1 U6176 ( .A1(n4858), .A2(n4861), .ZN(n4541) );
  OR2_X1 U6177 ( .A1(n8916), .A2(n8896), .ZN(n4542) );
  NAND2_X1 U6178 ( .A1(n8561), .A2(n7687), .ZN(n4543) );
  AND2_X1 U6179 ( .A1(n8212), .A2(n9294), .ZN(n4544) );
  AND2_X1 U6180 ( .A1(n6555), .A2(n6557), .ZN(n8199) );
  INV_X1 U6181 ( .A(n6582), .ZN(n4955) );
  NAND2_X1 U6182 ( .A1(n5485), .A2(n5484), .ZN(n8221) );
  NAND2_X1 U6183 ( .A1(n5085), .A2(n5086), .ZN(n6494) );
  NAND2_X1 U6184 ( .A1(n5512), .A2(n5104), .ZN(n5885) );
  NAND2_X1 U6185 ( .A1(n5086), .A2(n6076), .ZN(n6207) );
  NAND2_X1 U6186 ( .A1(n6490), .A2(n6078), .ZN(n6498) );
  INV_X1 U6187 ( .A(n9858), .ZN(n9690) );
  AND2_X1 U6188 ( .A1(n5558), .A2(n5557), .ZN(n9858) );
  INV_X1 U6189 ( .A(n6050), .ZN(n5999) );
  NOR2_X1 U6190 ( .A1(n5873), .A2(n5741), .ZN(n6050) );
  AND3_X1 U6191 ( .A1(n4876), .A2(n5170), .A3(n4875), .ZN(n4545) );
  AND2_X1 U6192 ( .A1(n4843), .A2(n5834), .ZN(n4546) );
  INV_X1 U6193 ( .A(n5051), .ZN(n5050) );
  NOR2_X1 U6194 ( .A1(n5057), .A2(n5052), .ZN(n5051) );
  INV_X1 U6195 ( .A(n5880), .ZN(n5881) );
  OAI211_X1 U6196 ( .C1(n5879), .C2(n6056), .A(n5732), .B(n9286), .ZN(n5880)
         );
  AND2_X1 U6197 ( .A1(n9676), .A2(n5767), .ZN(n4547) );
  NOR2_X1 U6198 ( .A1(n7897), .A2(n4800), .ZN(n4799) );
  OR2_X1 U6199 ( .A1(n6732), .A2(n4981), .ZN(n4548) );
  OR2_X1 U6200 ( .A1(n4912), .A2(n4911), .ZN(n4549) );
  NOR2_X1 U6201 ( .A1(n9134), .A2(n9726), .ZN(n4550) );
  OR2_X1 U6202 ( .A1(n4914), .A2(n4655), .ZN(n4551) );
  INV_X1 U6203 ( .A(n8212), .ZN(n9240) );
  AND2_X1 U6204 ( .A1(n4733), .A2(n4732), .ZN(n4552) );
  INV_X1 U6205 ( .A(n5124), .ZN(n5123) );
  INV_X1 U6206 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5556) );
  INV_X1 U6207 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6082) );
  NOR2_X1 U6208 ( .A1(n9301), .A2(n7469), .ZN(n4553) );
  INV_X1 U6209 ( .A(n5877), .ZN(n4785) );
  NAND2_X1 U6210 ( .A1(n5879), .A2(n6056), .ZN(n5877) );
  NOR2_X1 U6211 ( .A1(n9605), .A2(n9584), .ZN(n4554) );
  NOR2_X1 U6212 ( .A1(n9292), .A2(n9652), .ZN(n4555) );
  NOR2_X1 U6213 ( .A1(n8817), .A2(n8831), .ZN(n4556) );
  AND2_X1 U6214 ( .A1(n7969), .A2(n8559), .ZN(n4557) );
  INV_X1 U6215 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5174) );
  AND2_X1 U6216 ( .A1(n4645), .A2(n4649), .ZN(n4558) );
  NAND2_X1 U6217 ( .A1(n6727), .A2(n4821), .ZN(n4559) );
  XNOR2_X1 U6218 ( .A(n5597), .B(n5598), .ZN(n6132) );
  NOR2_X1 U6219 ( .A1(n9298), .A2(n7987), .ZN(n4560) );
  INV_X1 U6220 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5960) );
  AND2_X1 U6221 ( .A1(n6016), .A2(n7395), .ZN(n4561) );
  AOI21_X1 U6222 ( .B1(n5610), .B2(n4996), .A(n4993), .ZN(n4992) );
  INV_X1 U6223 ( .A(n8147), .ZN(n4874) );
  AND2_X1 U6224 ( .A1(n4607), .A2(n4604), .ZN(n4562) );
  INV_X1 U6225 ( .A(n4766), .ZN(n4765) );
  NOR2_X1 U6226 ( .A1(n5510), .A2(SI_14_), .ZN(n4766) );
  INV_X1 U6227 ( .A(n9848), .ZN(n9626) );
  AND2_X1 U6228 ( .A1(n5664), .A2(n5663), .ZN(n9848) );
  AND2_X1 U6229 ( .A1(n5764), .A2(n5997), .ZN(n9527) );
  AND2_X1 U6230 ( .A1(n5228), .A2(n5227), .ZN(n4563) );
  OR2_X1 U6231 ( .A1(n5128), .A2(n6038), .ZN(n4564) );
  OR2_X1 U6232 ( .A1(n6726), .A2(n6725), .ZN(n4565) );
  INV_X1 U6233 ( .A(n4886), .ZN(n4885) );
  NAND2_X1 U6234 ( .A1(n9174), .A2(n4887), .ZN(n4886) );
  OR2_X1 U6235 ( .A1(n9643), .A2(n9291), .ZN(n4566) );
  AND2_X1 U6236 ( .A1(n9734), .A2(n9701), .ZN(n4567) );
  AND2_X1 U6237 ( .A1(n6546), .A2(n6792), .ZN(n4568) );
  AND2_X1 U6238 ( .A1(n4963), .A2(n6551), .ZN(n4569) );
  AND2_X1 U6239 ( .A1(n4975), .A2(n6082), .ZN(n4570) );
  OR2_X1 U6240 ( .A1(n7576), .A2(n7618), .ZN(n4571) );
  AND2_X1 U6241 ( .A1(n9685), .A2(n5767), .ZN(n4572) );
  AND2_X1 U6242 ( .A1(n8663), .A2(n4738), .ZN(n4573) );
  AND2_X1 U6243 ( .A1(n4894), .A2(n4889), .ZN(n4574) );
  AND2_X1 U6244 ( .A1(n4714), .A2(n9240), .ZN(n4575) );
  AND2_X1 U6245 ( .A1(n8139), .A2(n8137), .ZN(n4576) );
  AND2_X1 U6246 ( .A1(n6078), .A2(n5090), .ZN(n4577) );
  AND2_X1 U6247 ( .A1(n6429), .A2(n6697), .ZN(n4578) );
  INV_X1 U6248 ( .A(n4828), .ZN(n4827) );
  NAND2_X1 U6249 ( .A1(n8814), .A2(n4829), .ZN(n4828) );
  NOR2_X1 U6250 ( .A1(n7932), .A2(n4966), .ZN(n4965) );
  XNOR2_X1 U6251 ( .A(n5737), .B(n5736), .ZN(n7811) );
  INV_X1 U6252 ( .A(n9215), .ZN(n4909) );
  AND4_X1 U6253 ( .A1(n5579), .A2(n5578), .A3(n5577), .A4(n5576), .ZN(n9661)
         );
  INV_X1 U6254 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5206) );
  XOR2_X1 U6255 ( .A(n5253), .B(SI_18_), .Z(n4579) );
  AND3_X1 U6256 ( .A1(n9162), .A2(n9906), .A3(n9161), .ZN(n4580) );
  NAND2_X1 U6257 ( .A1(n5600), .A2(n5599), .ZN(n9752) );
  INV_X1 U6258 ( .A(n9752), .ZN(n4707) );
  INV_X1 U6259 ( .A(n9295), .ZN(n6023) );
  AND2_X1 U6260 ( .A1(n4634), .A2(n4633), .ZN(n4581) );
  NAND2_X1 U6261 ( .A1(n6240), .A2(n6075), .ZN(n6257) );
  NOR2_X1 U6262 ( .A1(n8092), .A2(n8053), .ZN(n4582) );
  NOR2_X1 U6263 ( .A1(n8587), .A2(n8588), .ZN(n4583) );
  NOR2_X1 U6264 ( .A1(n9640), .A2(n9626), .ZN(n9599) );
  INV_X1 U6265 ( .A(n5027), .ZN(n5026) );
  NOR2_X1 U6266 ( .A1(n5550), .A2(n5028), .ZN(n5027) );
  NAND2_X1 U6267 ( .A1(n8154), .A2(n4519), .ZN(n4720) );
  AND2_X1 U6268 ( .A1(n8367), .A2(n8366), .ZN(n4584) );
  AND2_X1 U6269 ( .A1(n4925), .A2(n4924), .ZN(n4585) );
  AND2_X1 U6270 ( .A1(n8988), .A2(n8864), .ZN(n4586) );
  NAND2_X1 U6271 ( .A1(n8321), .A2(n4627), .ZN(n4587) );
  INV_X1 U6272 ( .A(n8386), .ZN(n5052) );
  AND4_X1 U6273 ( .A1(n5549), .A2(n5548), .A3(n5547), .A4(n5546), .ZN(n9278)
         );
  INV_X1 U6274 ( .A(n9278), .ZN(n4793) );
  AND2_X1 U6275 ( .A1(n4932), .A2(n4931), .ZN(n4588) );
  INV_X1 U6276 ( .A(n9903), .ZN(n9920) );
  NAND2_X1 U6277 ( .A1(n6659), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U6278 ( .A1(n7777), .A2(n4714), .ZN(n4589) );
  NAND2_X1 U6279 ( .A1(n4824), .A2(n6690), .ZN(n7681) );
  OR2_X1 U6280 ( .A1(n8602), .A2(n9000), .ZN(n4590) );
  NOR2_X1 U6281 ( .A1(n7867), .A2(n7868), .ZN(n4591) );
  AND2_X1 U6282 ( .A1(n4797), .A2(n4795), .ZN(n4592) );
  INV_X1 U6283 ( .A(SI_15_), .ZN(n4760) );
  INV_X1 U6284 ( .A(n5154), .ZN(n5097) );
  AND2_X1 U6285 ( .A1(n6835), .A2(n8699), .ZN(n9997) );
  INV_X2 U6286 ( .A(n9985), .ZN(n9988) );
  XNOR2_X1 U6287 ( .A(n4679), .B(n6082), .ZN(n6672) );
  INV_X1 U6288 ( .A(n7411), .ZN(n4706) );
  XOR2_X1 U6289 ( .A(n8705), .B(n8984), .Z(n4593) );
  AND2_X1 U6290 ( .A1(n6003), .A2(n6002), .ZN(n9659) );
  AND2_X1 U6291 ( .A1(n7147), .A2(n7137), .ZN(n9906) );
  NOR2_X1 U6292 ( .A1(n10021), .A2(n6360), .ZN(n4594) );
  AND2_X1 U6293 ( .A1(n8658), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4595) );
  OR2_X1 U6294 ( .A1(n9988), .A2(n4853), .ZN(n4596) );
  AND2_X1 U6295 ( .A1(n4619), .A2(n4618), .ZN(n4597) );
  AND2_X1 U6296 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n4598) );
  INV_X1 U6297 ( .A(n8705), .ZN(n7531) );
  INV_X1 U6298 ( .A(n6750), .ZN(n5078) );
  INV_X1 U6299 ( .A(n7652), .ZN(n6778) );
  NAND2_X1 U6300 ( .A1(n6497), .A2(n6496), .ZN(n7652) );
  INV_X1 U6301 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5076) );
  XNOR2_X1 U6302 ( .A(n8586), .B(n8599), .ZN(n8572) );
  XNOR2_X1 U6303 ( .A(n8598), .B(n8599), .ZN(n8568) );
  NAND2_X1 U6304 ( .A1(n7020), .A2(n6014), .ZN(n7152) );
  NAND2_X1 U6305 ( .A1(n4599), .A2(n9860), .ZN(n6059) );
  NAND2_X1 U6306 ( .A1(n4852), .A2(n4855), .ZN(n4599) );
  NAND2_X1 U6307 ( .A1(n7537), .A2(n5153), .ZN(n7655) );
  NAND2_X1 U6308 ( .A1(n6045), .A2(n5121), .ZN(n5120) );
  NAND2_X1 U6309 ( .A1(n5958), .A2(n5138), .ZN(n4713) );
  OAI21_X1 U6310 ( .B1(n9720), .B2(n4567), .A(n4529), .ZN(n4609) );
  NAND2_X1 U6311 ( .A1(n9244), .A2(n4537), .ZN(n4916) );
  OR2_X1 U6312 ( .A1(n6860), .A2(n5706), .ZN(n5445) );
  INV_X1 U6313 ( .A(n7623), .ZN(n4903) );
  NAND2_X2 U6314 ( .A1(n9897), .A2(n9898), .ZN(n9896) );
  NAND2_X1 U6315 ( .A1(n4651), .A2(n8273), .ZN(n9244) );
  INV_X1 U6316 ( .A(n4916), .ZN(n4912) );
  NAND2_X1 U6317 ( .A1(n8104), .A2(n8103), .ZN(n8107) );
  NAND2_X1 U6318 ( .A1(n9204), .A2(n9205), .ZN(n4900) );
  NAND3_X4 U6319 ( .A1(n9946), .A2(n7240), .A3(n4656), .ZN(n8310) );
  INV_X2 U6320 ( .A(n6664), .ZN(n6081) );
  NAND2_X1 U6321 ( .A1(n4695), .A2(n4693), .ZN(n6664) );
  OAI22_X2 U6322 ( .A1(n8840), .A2(n8839), .B1(n8854), .B2(n6716), .ZN(n8825)
         );
  OR2_X1 U6323 ( .A1(n5187), .A2(SI_1_), .ZN(n5188) );
  NAND2_X1 U6324 ( .A1(n4971), .A2(n4969), .ZN(n6475) );
  NAND2_X1 U6325 ( .A1(n8862), .A2(n8863), .ZN(n4803) );
  NAND2_X1 U6326 ( .A1(n6698), .A2(n4578), .ZN(n8039) );
  INV_X1 U6327 ( .A(n8769), .ZN(n6482) );
  NAND2_X1 U6328 ( .A1(n4806), .A2(n4809), .ZN(n8322) );
  INV_X1 U6329 ( .A(n7306), .ZN(n6679) );
  OAI21_X1 U6330 ( .B1(n7680), .B2(n6532), .A(n6531), .ZN(n7789) );
  NAND2_X1 U6331 ( .A1(n6028), .A2(n5155), .ZN(n9720) );
  INV_X1 U6332 ( .A(n4609), .ZN(n9705) );
  NOR2_X2 U6333 ( .A1(n8677), .A2(n8676), .ZN(n8698) );
  AOI21_X2 U6334 ( .B1(n6802), .B2(n6998), .A(n6980), .ZN(n7002) );
  NAND2_X1 U6335 ( .A1(n5107), .A2(n5110), .ZN(n7774) );
  NAND2_X1 U6336 ( .A1(n5098), .A2(n5101), .ZN(n7535) );
  NAND2_X1 U6337 ( .A1(n4562), .A2(n4938), .ZN(n4937) );
  XNOR2_X2 U6338 ( .A(n5177), .B(n5176), .ZN(n9874) );
  OAI211_X1 U6339 ( .C1(n4855), .C2(n9985), .A(n4851), .B(n4596), .ZN(P1_U3551) );
  NOR2_X2 U6340 ( .A1(n5147), .A2(n4849), .ZN(n4852) );
  MUX2_X1 U6341 ( .A(n6504), .B(n6503), .S(n6792), .Z(n6516) );
  NAND3_X1 U6342 ( .A1(n6539), .A2(n4614), .A3(n4612), .ZN(n6550) );
  NAND2_X1 U6343 ( .A1(n6556), .A2(n6555), .ZN(n4692) );
  OAI211_X1 U6344 ( .C1(n6558), .C2(n6792), .A(n8171), .B(n4689), .ZN(n6563)
         );
  NAND2_X1 U6345 ( .A1(n5034), .A2(n5033), .ZN(n5031) );
  OAI21_X1 U6346 ( .B1(n6614), .B2(n6615), .A(n4616), .ZN(n6625) );
  AOI21_X1 U6347 ( .B1(n4704), .B2(n7652), .A(n4703), .ZN(n6658) );
  NAND2_X1 U6348 ( .A1(n6640), .A2(n6733), .ZN(n6645) );
  NOR2_X1 U6349 ( .A1(n6650), .A2(n6649), .ZN(n5035) );
  AND2_X1 U6350 ( .A1(n4532), .A2(n4617), .ZN(n8332) );
  NAND2_X1 U6351 ( .A1(n7260), .A2(n7259), .ZN(n4617) );
  NAND2_X1 U6352 ( .A1(n8331), .A2(n4532), .ZN(n7261) );
  NAND2_X1 U6353 ( .A1(n9186), .A2(n8301), .ZN(n9264) );
  NAND2_X1 U6354 ( .A1(n4625), .A2(n4620), .ZN(P1_U3214) );
  NAND2_X1 U6355 ( .A1(n9225), .A2(n9223), .ZN(n8269) );
  NAND2_X1 U6356 ( .A1(n4632), .A2(n8260), .ZN(n9225) );
  NAND3_X1 U6357 ( .A1(n8256), .A2(n9252), .A3(n4877), .ZN(n4632) );
  NAND2_X1 U6358 ( .A1(n8254), .A2(n8255), .ZN(n9252) );
  NAND2_X1 U6359 ( .A1(n9251), .A2(n9253), .ZN(n8256) );
  NAND2_X1 U6360 ( .A1(n5555), .A2(n4639), .ZN(n4637) );
  NAND2_X1 U6361 ( .A1(n8275), .A2(n4649), .ZN(n4648) );
  NAND2_X1 U6362 ( .A1(n7146), .A2(n7923), .ZN(n4656) );
  NAND2_X4 U6363 ( .A1(n7133), .A2(n8310), .ZN(n8233) );
  AND2_X1 U6364 ( .A1(n7240), .A2(n7039), .ZN(n4657) );
  NOR2_X2 U6365 ( .A1(n5408), .A2(n5168), .ZN(n5512) );
  NAND4_X1 U6366 ( .A1(n5165), .A2(n5166), .A3(n5167), .A4(n5164), .ZN(n5168)
         );
  NAND2_X1 U6367 ( .A1(n7694), .A2(n4663), .ZN(n4661) );
  NAND2_X1 U6368 ( .A1(n4665), .A2(n7015), .ZN(n6815) );
  NAND2_X1 U6369 ( .A1(n6815), .A2(n4668), .ZN(n7184) );
  NAND3_X1 U6370 ( .A1(n4669), .A2(n6815), .A3(P2_REG1_REG_3__SCAN_IN), .ZN(
        n4668) );
  NAND3_X1 U6371 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4678) );
  NAND2_X2 U6372 ( .A1(n6673), .A2(n4516), .ZN(n6795) );
  INV_X1 U6373 ( .A(n6229), .ZN(n4693) );
  NAND3_X1 U6374 ( .A1(n6240), .A2(n4694), .A3(n6075), .ZN(n6229) );
  AND2_X2 U6375 ( .A1(n4986), .A2(n4577), .ZN(n4985) );
  NAND2_X1 U6376 ( .A1(n4699), .A2(n4696), .ZN(n6631) );
  NAND2_X1 U6377 ( .A1(n4697), .A2(n6741), .ZN(n4696) );
  NAND2_X1 U6378 ( .A1(n4698), .A2(n6626), .ZN(n4697) );
  OAI21_X1 U6379 ( .B1(n6625), .B2(n8770), .A(n6624), .ZN(n4698) );
  NAND2_X1 U6380 ( .A1(n6627), .A2(n6792), .ZN(n4699) );
  NAND3_X1 U6381 ( .A1(n5032), .A2(n5031), .A3(n6656), .ZN(n4704) );
  NAND2_X2 U6382 ( .A1(n6871), .A2(n6318), .ZN(n5728) );
  AND2_X2 U6383 ( .A1(n4834), .A2(n4709), .ZN(n9944) );
  NAND2_X1 U6384 ( .A1(n6060), .A2(n9813), .ZN(n9476) );
  NAND2_X1 U6385 ( .A1(n8154), .A2(n4717), .ZN(n9669) );
  INV_X1 U6386 ( .A(n4720), .ZN(n9689) );
  XNOR2_X1 U6387 ( .A(n8052), .B(n8097), .ZN(n8093) );
  NAND2_X1 U6388 ( .A1(n7713), .A2(n4727), .ZN(n4724) );
  INV_X1 U6389 ( .A(n4729), .ZN(n10024) );
  XNOR2_X1 U6390 ( .A(n8628), .B(n8641), .ZN(n8611) );
  OAI21_X1 U6391 ( .B1(n8572), .B2(n4736), .A(n4735), .ZN(n8610) );
  NAND2_X1 U6392 ( .A1(n5440), .A2(n4749), .ZN(n4748) );
  OAI21_X1 U6393 ( .B1(n5440), .B2(n4751), .A(n4749), .ZN(n5407) );
  OAI21_X1 U6394 ( .B1(n5453), .B2(n4770), .A(n4767), .ZN(n5494) );
  INV_X1 U6395 ( .A(n5882), .ZN(n4776) );
  NAND3_X1 U6396 ( .A1(n5829), .A2(n5768), .A3(n4791), .ZN(n4790) );
  INV_X1 U6397 ( .A(n7791), .ZN(n4796) );
  OAI21_X1 U6398 ( .B1(n7791), .B2(n6694), .A(n6693), .ZN(n7896) );
  NAND2_X1 U6399 ( .A1(n4803), .A2(n4801), .ZN(n6715) );
  NAND2_X1 U6400 ( .A1(n6736), .A2(n8914), .ZN(n4806) );
  NAND2_X1 U6401 ( .A1(n6719), .A2(n6718), .ZN(n8787) );
  NAND2_X1 U6402 ( .A1(n6719), .A2(n4813), .ZN(n4812) );
  NAND2_X1 U6403 ( .A1(n4824), .A2(n4823), .ZN(n6692) );
  AND2_X1 U6404 ( .A1(n6690), .A2(n4543), .ZN(n4823) );
  OAI21_X1 U6405 ( .B1(n8825), .B2(n4828), .A(n4825), .ZN(n8796) );
  NAND2_X1 U6406 ( .A1(n8039), .A2(n6699), .ZN(n8173) );
  INV_X1 U6407 ( .A(n6345), .ZN(n4831) );
  INV_X1 U6409 ( .A(n6259), .ZN(n5086) );
  INV_X1 U6410 ( .A(n7024), .ZN(n6013) );
  NAND2_X1 U6411 ( .A1(n7155), .A2(n5893), .ZN(n4836) );
  NAND2_X1 U6412 ( .A1(n4841), .A2(n4839), .ZN(n7947) );
  NAND2_X1 U6413 ( .A1(n9637), .A2(n4845), .ZN(n4844) );
  OR2_X2 U6414 ( .A1(n4854), .A2(n4850), .ZN(n4849) );
  NAND2_X1 U6415 ( .A1(n9580), .A2(n4859), .ZN(n4857) );
  NAND2_X1 U6416 ( .A1(n9580), .A2(n4863), .ZN(n4858) );
  INV_X1 U6417 ( .A(n5408), .ZN(n4876) );
  NAND3_X1 U6418 ( .A1(n5105), .A2(n5137), .A3(n4545), .ZN(n5139) );
  XNOR2_X2 U6419 ( .A(n6297), .B(n6296), .ZN(n7015) );
  NAND2_X1 U6420 ( .A1(n8256), .A2(n9252), .ZN(n4878) );
  XNOR2_X1 U6421 ( .A(n4878), .B(n9143), .ZN(n9147) );
  NAND2_X2 U6422 ( .A1(n5973), .A2(n4879), .ZN(n7240) );
  NAND3_X1 U6423 ( .A1(n4892), .A2(n4890), .A3(n4574), .ZN(P1_U3220) );
  NAND2_X1 U6424 ( .A1(n9264), .A2(n4891), .ZN(n4890) );
  OR2_X1 U6425 ( .A1(n9264), .A2(n4896), .ZN(n4892) );
  NAND2_X1 U6426 ( .A1(n4900), .A2(n9206), .ZN(n8254) );
  NAND2_X1 U6427 ( .A1(n4900), .A2(n4898), .ZN(n9251) );
  NAND2_X1 U6428 ( .A1(n7623), .A2(n7620), .ZN(n4901) );
  NAND2_X1 U6429 ( .A1(n4904), .A2(n4906), .ZN(n5964) );
  INV_X2 U6430 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4919) );
  INV_X1 U6431 ( .A(n4932), .ZN(n8600) );
  INV_X1 U6432 ( .A(n7866), .ZN(n4933) );
  NOR2_X4 U6433 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6811) );
  INV_X1 U6434 ( .A(n6811), .ZN(n4943) );
  OAI21_X2 U6435 ( .B1(n6480), .B2(n4947), .A(n4944), .ZN(n8769) );
  NAND2_X1 U6436 ( .A1(n6469), .A2(n7501), .ZN(n7498) );
  NAND2_X1 U6437 ( .A1(n7498), .A2(n4949), .ZN(n4948) );
  NAND2_X1 U6438 ( .A1(n4948), .A2(n6527), .ZN(n7680) );
  OAI22_X2 U6439 ( .A1(n6477), .A2(n4951), .B1(n4953), .B2(n6478), .ZN(n8850)
         );
  NAND2_X1 U6440 ( .A1(n4960), .A2(n4958), .ZN(n6483) );
  INV_X1 U6441 ( .A(n6632), .ZN(n4961) );
  NAND2_X1 U6442 ( .A1(n7895), .A2(n4965), .ZN(n4962) );
  NAND2_X1 U6443 ( .A1(n4962), .A2(n4569), .ZN(n6472) );
  INV_X1 U6444 ( .A(n7895), .ZN(n4968) );
  NAND2_X1 U6445 ( .A1(n8172), .A2(n4972), .ZN(n4971) );
  NAND2_X1 U6446 ( .A1(n8837), .A2(n4974), .ZN(n8812) );
  NAND2_X1 U6447 ( .A1(n6081), .A2(n4975), .ZN(n6092) );
  AND2_X2 U6448 ( .A1(n6081), .A2(n4570), .ZN(n6097) );
  NAND2_X1 U6449 ( .A1(n6081), .A2(n6080), .ZN(n6083) );
  NAND2_X1 U6450 ( .A1(n8719), .A2(n4977), .ZN(n4976) );
  NAND2_X1 U6451 ( .A1(n8719), .A2(n8718), .ZN(n4982) );
  NAND2_X1 U6452 ( .A1(n4976), .A2(n4978), .ZN(n6492) );
  NAND2_X1 U6453 ( .A1(n4982), .A2(n6485), .ZN(n6737) );
  NOR2_X1 U6454 ( .A1(n6489), .A2(n4984), .ZN(n4983) );
  AOI21_X1 U6455 ( .B1(n5344), .B2(n4991), .A(n4990), .ZN(n4988) );
  NAND2_X1 U6456 ( .A1(n5361), .A2(n5360), .ZN(n5363) );
  INV_X1 U6457 ( .A(n4992), .ZN(n5295) );
  NAND2_X1 U6458 ( .A1(n5662), .A2(n5003), .ZN(n5001) );
  OAI21_X1 U6459 ( .B1(n5662), .B2(n5264), .A(n5263), .ZN(n5639) );
  NAND2_X1 U6460 ( .A1(n5277), .A2(n5276), .ZN(n5648) );
  NAND2_X1 U6461 ( .A1(n5277), .A2(n5014), .ZN(n5013) );
  OAI21_X1 U6462 ( .B1(n5539), .B2(n5023), .A(n5021), .ZN(n5580) );
  NAND2_X1 U6463 ( .A1(n5030), .A2(n5029), .ZN(n5453) );
  NAND3_X1 U6464 ( .A1(n6655), .A2(n6654), .A3(n4538), .ZN(n5032) );
  OAI21_X1 U6465 ( .B1(n6646), .B2(n9016), .A(n5035), .ZN(n5034) );
  NAND2_X2 U6466 ( .A1(n5038), .A2(n5036), .ZN(n5203) );
  NAND3_X1 U6467 ( .A1(n5037), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5036) );
  NAND3_X1 U6468 ( .A1(n10551), .A2(n9473), .A3(n5039), .ZN(n5038) );
  OAI21_X1 U6469 ( .B1(n8473), .B2(n8387), .A(n8386), .ZN(n8447) );
  INV_X1 U6470 ( .A(n5047), .ZN(n8423) );
  NAND2_X1 U6471 ( .A1(n8184), .A2(n5068), .ZN(n5067) );
  OAI211_X1 U6472 ( .C1(n8201), .C2(n5069), .A(n5067), .B(n5065), .ZN(n8354)
         );
  NAND2_X1 U6473 ( .A1(n8350), .A2(n8349), .ZN(n8438) );
  NAND2_X1 U6474 ( .A1(n5070), .A2(n8200), .ZN(n8350) );
  INV_X1 U6475 ( .A(n8349), .ZN(n5069) );
  NAND4_X1 U6476 ( .A1(n6881), .A2(n5073), .A3(n5072), .A4(n5071), .ZN(n7089)
         );
  NAND2_X1 U6477 ( .A1(n5078), .A2(n5079), .ZN(n5077) );
  NAND3_X1 U6478 ( .A1(n5081), .A2(n7094), .A3(n7201), .ZN(n7202) );
  NAND2_X1 U6479 ( .A1(n7093), .A2(n6678), .ZN(n7201) );
  NAND2_X1 U6480 ( .A1(n8357), .A2(n5083), .ZN(n5082) );
  NAND2_X1 U6481 ( .A1(n5082), .A2(n8359), .ZN(n8540) );
  INV_X1 U6482 ( .A(n8540), .ZN(n8361) );
  NAND2_X1 U6483 ( .A1(n8138), .A2(n4576), .ZN(n8182) );
  NAND2_X1 U6484 ( .A1(n7593), .A2(n5087), .ZN(n7852) );
  NAND3_X1 U6485 ( .A1(n5092), .A2(n5334), .A3(n5364), .ZN(n5400) );
  NAND2_X1 U6486 ( .A1(n5094), .A2(n5093), .ZN(n6028) );
  NAND2_X1 U6487 ( .A1(n6027), .A2(n5095), .ZN(n5094) );
  NAND2_X1 U6488 ( .A1(n7377), .A2(n5099), .ZN(n5098) );
  NAND2_X1 U6489 ( .A1(n7655), .A2(n5108), .ZN(n5107) );
  NAND2_X1 U6490 ( .A1(n9667), .A2(n5118), .ZN(n5117) );
  NAND2_X1 U6491 ( .A1(n5120), .A2(n5119), .ZN(n9504) );
  NOR2_X1 U6492 ( .A1(n9544), .A2(n9524), .ZN(n5124) );
  NAND2_X1 U6493 ( .A1(n9616), .A2(n5127), .ZN(n5126) );
  INV_X1 U6494 ( .A(n5139), .ZN(n5298) );
  NAND2_X1 U6495 ( .A1(n5139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5299) );
  INV_X2 U6496 ( .A(n6871), .ZN(n5586) );
  NAND2_X2 U6497 ( .A1(n5966), .A2(n5967), .ZN(n6871) );
  OAI21_X2 U6498 ( .B1(n8732), .B2(n8731), .A(n6484), .ZN(n8719) );
  OR2_X1 U6499 ( .A1(n6339), .A2(n7305), .ZN(n6342) );
  INV_X1 U6500 ( .A(n6465), .ZN(n8925) );
  INV_X1 U6501 ( .A(n5709), .ZN(n5605) );
  OAI21_X2 U6502 ( .B1(n8894), .B2(n6708), .A(n6707), .ZN(n8884) );
  OAI21_X1 U6503 ( .B1(n5941), .B2(n5940), .A(n5939), .ZN(n5956) );
  INV_X1 U6504 ( .A(n9487), .ZN(n6009) );
  XNOR2_X1 U6505 ( .A(n5688), .B(n5689), .ZN(n9118) );
  AOI21_X2 U6506 ( .B1(n6482), .B2(n5151), .A(n5150), .ZN(n8757) );
  OAI21_X1 U6507 ( .B1(n5203), .B2(n5186), .A(n5185), .ZN(n5187) );
  NAND2_X1 U6508 ( .A1(n5203), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6509 ( .A1(n7254), .A2(n7253), .ZN(n7255) );
  OAI22_X1 U6510 ( .A1(n8733), .A2(n6728), .B1(n8750), .B2(n8743), .ZN(n8721)
         );
  AOI211_X1 U6511 ( .C1(n5926), .C2(n5714), .A(n5870), .B(n5741), .ZN(n5932)
         );
  OAI22_X2 U6512 ( .A1(n7444), .A2(n6685), .B1(n10038), .B2(n8929), .ZN(n7502)
         );
  NAND2_X1 U6513 ( .A1(n6880), .A2(n6752), .ZN(n6883) );
  OR2_X1 U6514 ( .A1(n6752), .A2(n6770), .ZN(n7210) );
  OR2_X1 U6515 ( .A1(n6752), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6755) );
  NAND2_X1 U6516 ( .A1(n6669), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6663) );
  AND2_X1 U6517 ( .A1(n9508), .A2(n9507), .ZN(n9750) );
  OAI21_X1 U6518 ( .B1(n7085), .B2(n6757), .A(n6756), .ZN(n7214) );
  AND2_X1 U6519 ( .A1(n7537), .A2(n7536), .ZN(n7738) );
  NAND2_X1 U6520 ( .A1(n9508), .A2(n6049), .ZN(n6051) );
  INV_X1 U6521 ( .A(n9874), .ZN(n5306) );
  OR2_X1 U6522 ( .A1(n6795), .A2(n6998), .ZN(n5142) );
  OR2_X1 U6523 ( .A1(n6338), .A2(n9994), .ZN(n5143) );
  OR2_X1 U6524 ( .A1(n7240), .A2(n9926), .ZN(n5144) );
  INV_X1 U6525 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8465) );
  AND2_X1 U6526 ( .A1(n4715), .A2(n9180), .ZN(n5145) );
  NAND2_X1 U6527 ( .A1(n5162), .A2(n6012), .ZN(n5147) );
  AND2_X1 U6528 ( .A1(n8658), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5148) );
  NOR2_X1 U6529 ( .A1(n6621), .A2(n6624), .ZN(n5150) );
  NOR2_X1 U6530 ( .A1(n8770), .A2(n6621), .ZN(n5151) );
  AND2_X1 U6531 ( .A1(n4511), .A2(n9152), .ZN(n5152) );
  OR2_X1 U6532 ( .A1(n7745), .A2(n9300), .ZN(n5153) );
  AND2_X1 U6533 ( .A1(n9240), .A2(n9179), .ZN(n5154) );
  OR2_X1 U6534 ( .A1(n9976), .A2(n9280), .ZN(n5155) );
  NAND2_X1 U6535 ( .A1(n7178), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U6536 ( .A1(n7178), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6833) );
  INV_X1 U6537 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6088) );
  AND2_X1 U6538 ( .A1(n7049), .A2(n7136), .ZN(n9727) );
  NOR2_X1 U6539 ( .A1(n8324), .A2(n9052), .ZN(n6785) );
  INV_X1 U6540 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5169) );
  INV_X1 U6541 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8431) );
  AND4_X1 U6542 ( .A1(n5618), .A2(n5617), .A3(n5616), .A4(n5615), .ZN(n9537)
         );
  INV_X1 U6543 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5175) );
  INV_X1 U6544 ( .A(n9646), .ZN(n9950) );
  INV_X1 U6545 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6094) );
  AND4_X1 U6546 ( .A1(n5869), .A2(n5868), .A3(n5867), .A4(n5866), .ZN(n5156)
         );
  OR2_X1 U6547 ( .A1(n9496), .A2(n9505), .ZN(n5157) );
  AND2_X1 U6548 ( .A1(n5870), .A2(n6056), .ZN(n5158) );
  OR2_X1 U6549 ( .A1(n9838), .A2(n9570), .ZN(n5159) );
  NOR2_X1 U6550 ( .A1(n5706), .A2(n6856), .ZN(n5160) );
  AND3_X2 U6551 ( .A1(n7214), .A2(n6771), .A3(n7101), .ZN(n10099) );
  NOR2_X1 U6552 ( .A1(n7919), .A2(n6781), .ZN(n10033) );
  INV_X1 U6553 ( .A(n8602), .ZN(n8619) );
  AND2_X1 U6554 ( .A1(n6328), .A2(n6327), .ZN(n5161) );
  INV_X1 U6555 ( .A(n8221), .ZN(n6024) );
  OR2_X1 U6556 ( .A1(n9491), .A2(n9969), .ZN(n5162) );
  INV_X1 U6557 ( .A(n7140), .ZN(n5937) );
  INV_X2 U6558 ( .A(n9612), .ZN(n9714) );
  AND4_X1 U6559 ( .A1(n5609), .A2(n5608), .A3(n5607), .A4(n5606), .ZN(n9525)
         );
  INV_X1 U6560 ( .A(n8123), .ZN(n9297) );
  NAND2_X1 U6561 ( .A1(n6511), .A2(n6792), .ZN(n6512) );
  AND2_X1 U6562 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  AOI21_X1 U6563 ( .B1(n6639), .B2(n6638), .A(n6637), .ZN(n6640) );
  NAND2_X1 U6564 ( .A1(n6733), .A2(n6643), .ZN(n6641) );
  AOI21_X1 U6565 ( .B1(n5871), .B2(n5156), .A(n5158), .ZN(n5872) );
  INV_X1 U6566 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6076) );
  INV_X1 U6567 ( .A(n8101), .ZN(n8102) );
  INV_X1 U6568 ( .A(n7776), .ZN(n5465) );
  INV_X1 U6569 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5172) );
  INV_X1 U6570 ( .A(n10026), .ZN(n8660) );
  AND2_X1 U6571 ( .A1(n9016), .A2(n8736), .ZN(n6730) );
  NAND2_X1 U6572 ( .A1(n8100), .A2(n8102), .ZN(n8103) );
  INV_X1 U6573 ( .A(n7904), .ZN(n5492) );
  INV_X1 U6574 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5164) );
  INV_X1 U6575 ( .A(n8142), .ZN(n8139) );
  NOR2_X1 U6576 ( .A1(n6175), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6155) );
  INV_X1 U6577 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10394) );
  INV_X1 U6578 ( .A(n6618), .ZN(n6481) );
  INV_X1 U6579 ( .A(P2_B_REG_SCAN_IN), .ZN(n6748) );
  INV_X1 U6580 ( .A(n7574), .ZN(n7575) );
  INV_X1 U6581 ( .A(n7811), .ZN(n5883) );
  NAND2_X1 U6582 ( .A1(n9487), .A2(n9956), .ZN(n6012) );
  NAND2_X1 U6583 ( .A1(n5896), .A2(n5770), .ZN(n5769) );
  INV_X1 U6584 ( .A(SI_24_), .ZN(n10388) );
  INV_X1 U6585 ( .A(SI_17_), .ZN(n10229) );
  INV_X1 U6586 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6084) );
  INV_X1 U6587 ( .A(n8464), .ZN(n8367) );
  OR2_X1 U6588 ( .A1(n6193), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6183) );
  AND2_X1 U6589 ( .A1(n6199), .A2(n10380), .ZN(n6191) );
  OR2_X1 U6590 ( .A1(n6422), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U6591 ( .A1(n7573), .A2(n7575), .ZN(n7576) );
  INV_X1 U6592 ( .A(n8284), .ZN(n8306) );
  AND2_X1 U6593 ( .A1(n5634), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5652) );
  AND2_X1 U6594 ( .A1(n5472), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5486) );
  AND2_X1 U6595 ( .A1(n9557), .A2(n9570), .ZN(n5995) );
  AND2_X1 U6596 ( .A1(n5590), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U6597 ( .A1(n6053), .A2(n5883), .ZN(n6004) );
  OR2_X1 U6598 ( .A1(n4512), .A2(n4833), .ZN(n6014) );
  INV_X1 U6599 ( .A(SI_20_), .ZN(n5672) );
  NAND2_X1 U6600 ( .A1(n5241), .A2(SI_13_), .ZN(n5245) );
  INV_X1 U6601 ( .A(n7199), .ZN(n8421) );
  INV_X1 U6602 ( .A(n6795), .ZN(n6445) );
  INV_X1 U6603 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6087) );
  INV_X1 U6604 ( .A(n8750), .ZN(n8530) );
  AND2_X1 U6605 ( .A1(n6810), .A2(n9111), .ZN(n6835) );
  OR2_X1 U6606 ( .A1(n6157), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6147) );
  OR2_X1 U6607 ( .A1(n10073), .A2(n7301), .ZN(n8915) );
  INV_X1 U6608 ( .A(n7085), .ZN(n7212) );
  INV_X1 U6609 ( .A(n8928), .ZN(n8909) );
  NAND2_X1 U6610 ( .A1(n6742), .A2(n6741), .ZN(n8928) );
  NOR2_X1 U6611 ( .A1(n7101), .A2(n6782), .ZN(n7115) );
  INV_X1 U6612 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U6613 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  NAND2_X1 U6614 ( .A1(n5486), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5517) );
  INV_X1 U6615 ( .A(n9726), .ZN(n9280) );
  INV_X1 U6616 ( .A(n5946), .ZN(n5947) );
  NAND2_X1 U6617 ( .A1(n5652), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5693) );
  OR2_X1 U6618 ( .A1(n5666), .A2(n9245), .ZN(n5643) );
  INV_X1 U6619 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9378) );
  OR2_X1 U6620 ( .A1(n7835), .A2(n7834), .ZN(n9441) );
  NAND2_X1 U6621 ( .A1(n9504), .A2(n6048), .ZN(n9508) );
  INV_X1 U6622 ( .A(n9599), .ZN(n9625) );
  INV_X1 U6623 ( .A(n9727), .ZN(n9662) );
  INV_X1 U6624 ( .A(n6004), .ZN(n7136) );
  INV_X1 U6625 ( .A(n7128), .ZN(n7129) );
  NAND2_X1 U6626 ( .A1(n9866), .A2(n7238), .ZN(n7028) );
  INV_X1 U6627 ( .A(n7146), .ZN(n6054) );
  OR2_X1 U6628 ( .A1(n9969), .A2(n7033), .ZN(n7128) );
  OAI21_X1 U6629 ( .B1(n5580), .B2(n5581), .A(n5260), .ZN(n5675) );
  INV_X1 U6630 ( .A(n5450), .ZN(n5233) );
  AND2_X1 U6631 ( .A1(n5225), .A2(n5224), .ZN(n5439) );
  INV_X1 U6632 ( .A(n8538), .ZN(n8515) );
  AND2_X1 U6633 ( .A1(n6152), .A2(n6151), .ZN(n8389) );
  AND4_X1 U6634 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n8399)
         );
  INV_X1 U6635 ( .A(n10011), .ZN(n10018) );
  OR2_X1 U6636 ( .A1(n8680), .A2(n6806), .ZN(n8707) );
  INV_X1 U6637 ( .A(n8707), .ZN(n10020) );
  OR2_X1 U6638 ( .A1(n9102), .A2(n7116), .ZN(n8899) );
  INV_X1 U6639 ( .A(n10044), .ZN(n7506) );
  INV_X1 U6640 ( .A(n8899), .ZN(n8937) );
  INV_X1 U6641 ( .A(n8980), .ZN(n9004) );
  NAND2_X1 U6642 ( .A1(n9103), .A2(n7212), .ZN(n7101) );
  INV_X1 U6643 ( .A(n10078), .ZN(n10080) );
  NAND2_X1 U6644 ( .A1(n6750), .A2(n6671), .ZN(n6821) );
  NOR2_X1 U6645 ( .A1(n5459), .A2(n9378), .ZN(n5472) );
  OR2_X1 U6646 ( .A1(n7127), .A2(n7394), .ZN(n7130) );
  INV_X1 U6647 ( .A(n5707), .ZN(n5656) );
  AND4_X1 U6648 ( .A1(n5595), .A2(n5594), .A3(n5593), .A4(n5592), .ZN(n9292)
         );
  NAND2_X1 U6649 ( .A1(n5708), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5325) );
  INV_X1 U6650 ( .A(n9936), .ZN(n6926) );
  XNOR2_X1 U6651 ( .A(n9745), .B(n9477), .ZN(n6060) );
  INV_X1 U6652 ( .A(n9664), .ZN(n9728) );
  NAND2_X1 U6653 ( .A1(n7775), .A2(n6021), .ZN(n7940) );
  INV_X1 U6654 ( .A(n9659), .ZN(n9724) );
  NOR2_X1 U6655 ( .A1(n7028), .A2(n7125), .ZN(n7029) );
  INV_X1 U6656 ( .A(n9979), .ZN(n9804) );
  AND2_X1 U6657 ( .A1(n6010), .A2(n6054), .ZN(n9956) );
  NAND2_X1 U6658 ( .A1(n7658), .A2(n7758), .ZN(n9979) );
  AND3_X1 U6659 ( .A1(n7123), .A2(n7122), .A3(n7128), .ZN(n7030) );
  XNOR2_X1 U6660 ( .A(n5953), .B(n5952), .ZN(n7239) );
  NAND2_X1 U6661 ( .A1(n5191), .A2(n5309), .ZN(n5313) );
  INV_X1 U6662 ( .A(n8533), .ZN(n8545) );
  AND2_X1 U6663 ( .A1(n7117), .A2(n8899), .ZN(n8551) );
  NAND2_X1 U6664 ( .A1(n6131), .A2(n6130), .ZN(n8750) );
  INV_X1 U6665 ( .A(n8466), .ZN(n8864) );
  OR2_X1 U6666 ( .A1(P2_U3150), .A2(n6822), .ZN(n10011) );
  INV_X1 U6667 ( .A(n9997), .ZN(n10022) );
  OR2_X1 U6668 ( .A1(n6970), .A2(n8699), .ZN(n10026) );
  AND2_X1 U6669 ( .A1(n7216), .A2(n8899), .ZN(n8920) );
  INV_X2 U6670 ( .A(n8920), .ZN(n8942) );
  NAND2_X1 U6671 ( .A1(n8942), .A2(n7302), .ZN(n8923) );
  NAND2_X1 U6672 ( .A1(n10099), .A2(n10085), .ZN(n8980) );
  NAND2_X1 U6673 ( .A1(n10099), .A2(n10078), .ZN(n9007) );
  INV_X1 U6674 ( .A(n10099), .ZN(n10097) );
  NOR2_X1 U6675 ( .A1(n6785), .A2(n6787), .ZN(n6788) );
  XNOR2_X1 U6676 ( .A(n8757), .B(n8756), .ZN(n9032) );
  OR2_X1 U6677 ( .A1(n10087), .A2(n10080), .ZN(n9100) );
  AND2_X1 U6678 ( .A1(n6784), .A2(n6783), .ZN(n10087) );
  INV_X2 U6679 ( .A(n10087), .ZN(n10086) );
  NAND2_X1 U6680 ( .A1(n6821), .A2(n7109), .ZN(n9102) );
  INV_X1 U6681 ( .A(n6100), .ZN(n8330) );
  INV_X1 U6682 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7651) );
  INV_X1 U6683 ( .A(n7360), .ZN(n7342) );
  INV_X1 U6684 ( .A(n9115), .ZN(n9105) );
  AND2_X1 U6685 ( .A1(n7130), .A2(n9711), .ZN(n9903) );
  AOI21_X1 U6686 ( .B1(n9558), .B2(n5354), .A(n5657), .ZN(n9570) );
  INV_X1 U6687 ( .A(n9661), .ZN(n9293) );
  OR2_X1 U6688 ( .A1(n6908), .A2(n6907), .ZN(n9936) );
  NAND2_X1 U6689 ( .A1(n6926), .A2(n5966), .ZN(n9459) );
  OR2_X1 U6690 ( .A1(n9612), .A2(n7391), .ZN(n9741) );
  NAND2_X1 U6691 ( .A1(n9988), .A2(n9956), .ZN(n9823) );
  NAND2_X1 U6692 ( .A1(n7030), .A2(n7029), .ZN(n9985) );
  INV_X1 U6693 ( .A(n9734), .ZN(n9865) );
  AND2_X2 U6694 ( .A1(n7390), .A2(n7030), .ZN(n9860) );
  INV_X1 U6695 ( .A(n9955), .ZN(n9954) );
  AND2_X1 U6696 ( .A1(n9866), .A2(n6864), .ZN(n9955) );
  INV_X1 U6697 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10495) );
  INV_X1 U6698 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10508) );
  INV_X2 U6699 ( .A(n8680), .ZN(P2_U3893) );
  NOR2_X2 U6700 ( .A1(n6791), .A2(n7240), .ZN(P1_U3973) );
  INV_X2 U6701 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U6702 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5167) );
  NOR2_X1 U6703 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5166) );
  NOR2_X1 U6704 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5165) );
  NOR2_X2 U6705 ( .A1(n5300), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n9868) );
  INV_X1 U6706 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5176) );
  AND2_X4 U6707 ( .A1(n5305), .A2(n9874), .ZN(n5708) );
  NAND2_X1 U6708 ( .A1(n5708), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5182) );
  AND2_X4 U6709 ( .A1(n5306), .A2(n9877), .ZN(n5709) );
  NAND2_X1 U6710 ( .A1(n5709), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5181) );
  AND2_X4 U6711 ( .A1(n9874), .A2(n9877), .ZN(n5707) );
  NAND2_X1 U6712 ( .A1(n5707), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5180) );
  NAND3_X1 U6713 ( .A1(n5182), .A2(n5181), .A3(n5180), .ZN(n9285) );
  INV_X1 U6714 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U6715 ( .A1(n5709), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6716 ( .A1(n5708), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5183) );
  OAI211_X1 U6717 ( .C1(n5656), .C2(n9825), .A(n5184), .B(n5183), .ZN(n9286)
         );
  NAND2_X1 U6718 ( .A1(n9285), .A2(n9286), .ZN(n5878) );
  NAND2_X1 U6719 ( .A1(n5187), .A2(SI_1_), .ZN(n5192) );
  INV_X1 U6720 ( .A(SI_1_), .ZN(n10222) );
  NAND2_X1 U6721 ( .A1(n5192), .A2(n5188), .ZN(n5311) );
  INV_X1 U6722 ( .A(n5311), .ZN(n5191) );
  INV_X1 U6723 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6319) );
  INV_X1 U6724 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5189) );
  MUX2_X1 U6725 ( .A(n6319), .B(n5189), .S(n5203), .Z(n5190) );
  NOR2_X1 U6726 ( .A1(n5190), .A2(n10280), .ZN(n5309) );
  NAND2_X1 U6727 ( .A1(n5313), .A2(n5192), .ZN(n5329) );
  MUX2_X1 U6728 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5203), .Z(n5193) );
  NAND2_X1 U6729 ( .A1(n5193), .A2(SI_2_), .ZN(n5197) );
  INV_X1 U6730 ( .A(n5193), .ZN(n5194) );
  INV_X1 U6731 ( .A(SI_2_), .ZN(n10395) );
  NAND2_X1 U6732 ( .A1(n5194), .A2(n10395), .ZN(n5195) );
  NAND2_X1 U6733 ( .A1(n5197), .A2(n5195), .ZN(n5330) );
  INV_X1 U6734 ( .A(n5330), .ZN(n5196) );
  NAND2_X1 U6735 ( .A1(n5329), .A2(n5196), .ZN(n5332) );
  MUX2_X1 U6736 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5203), .Z(n5200) );
  INV_X1 U6737 ( .A(n5200), .ZN(n5199) );
  INV_X1 U6738 ( .A(SI_3_), .ZN(n5198) );
  NAND2_X1 U6739 ( .A1(n5199), .A2(n5198), .ZN(n5201) );
  NAND2_X1 U6740 ( .A1(n5200), .A2(SI_3_), .ZN(n5202) );
  INV_X1 U6741 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5204) );
  INV_X1 U6742 ( .A(n5209), .ZN(n5208) );
  INV_X1 U6743 ( .A(SI_4_), .ZN(n5207) );
  NAND2_X1 U6744 ( .A1(n5208), .A2(n5207), .ZN(n5210) );
  NAND2_X1 U6745 ( .A1(n5209), .A2(SI_4_), .ZN(n5211) );
  NAND2_X1 U6746 ( .A1(n5363), .A2(n5211), .ZN(n5383) );
  MUX2_X1 U6747 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6847), .Z(n5212) );
  NAND2_X1 U6748 ( .A1(n5212), .A2(SI_5_), .ZN(n5215) );
  INV_X1 U6749 ( .A(n5212), .ZN(n5213) );
  INV_X1 U6750 ( .A(SI_5_), .ZN(n10483) );
  NAND2_X1 U6751 ( .A1(n5213), .A2(n10483), .ZN(n5214) );
  AND2_X1 U6752 ( .A1(n5215), .A2(n5214), .ZN(n5382) );
  NAND2_X1 U6753 ( .A1(n5383), .A2(n5382), .ZN(n5385) );
  NAND2_X1 U6754 ( .A1(n5385), .A2(n5215), .ZN(n5397) );
  MUX2_X1 U6755 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6847), .Z(n5216) );
  NAND2_X1 U6756 ( .A1(n5216), .A2(SI_6_), .ZN(n5220) );
  INV_X1 U6757 ( .A(n5216), .ZN(n5218) );
  INV_X1 U6758 ( .A(SI_6_), .ZN(n5217) );
  NAND2_X1 U6759 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  AND2_X1 U6760 ( .A1(n5220), .A2(n5219), .ZN(n5396) );
  NAND2_X1 U6761 ( .A1(n5397), .A2(n5396), .ZN(n5399) );
  MUX2_X1 U6762 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6847), .Z(n5221) );
  NAND2_X1 U6763 ( .A1(n5221), .A2(SI_7_), .ZN(n5225) );
  INV_X1 U6764 ( .A(n5221), .ZN(n5223) );
  INV_X1 U6765 ( .A(SI_7_), .ZN(n5222) );
  NAND2_X1 U6766 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  MUX2_X1 U6767 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6847), .Z(n5226) );
  XNOR2_X1 U6768 ( .A(n5226), .B(SI_8_), .ZN(n5422) );
  INV_X1 U6769 ( .A(n5226), .ZN(n5228) );
  INV_X1 U6770 ( .A(SI_8_), .ZN(n5227) );
  MUX2_X1 U6771 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n6847), .Z(n5229) );
  XNOR2_X1 U6772 ( .A(n5229), .B(n10290), .ZN(n5406) );
  INV_X1 U6773 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6774 ( .A1(n5230), .A2(n10290), .ZN(n5231) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6847), .Z(n5232) );
  NAND2_X1 U6776 ( .A1(n5232), .A2(SI_10_), .ZN(n5234) );
  OAI21_X1 U6777 ( .B1(n5232), .B2(SI_10_), .A(n5234), .ZN(n5450) );
  MUX2_X1 U6778 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6847), .Z(n5235) );
  XNOR2_X1 U6779 ( .A(n5235), .B(SI_11_), .ZN(n5466) );
  INV_X1 U6780 ( .A(n5235), .ZN(n5237) );
  INV_X1 U6781 ( .A(SI_11_), .ZN(n5236) );
  NAND2_X1 U6782 ( .A1(n5237), .A2(n5236), .ZN(n5238) );
  MUX2_X1 U6783 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6847), .Z(n5239) );
  NAND2_X1 U6784 ( .A1(n5239), .A2(SI_12_), .ZN(n5240) );
  OAI21_X1 U6785 ( .B1(n5239), .B2(SI_12_), .A(n5240), .ZN(n5479) );
  MUX2_X1 U6786 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6847), .Z(n5241) );
  INV_X1 U6787 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U6788 ( .A1(n5242), .A2(n10481), .ZN(n5243) );
  NAND2_X1 U6789 ( .A1(n5245), .A2(n5243), .ZN(n5495) );
  INV_X1 U6790 ( .A(n5495), .ZN(n5244) );
  MUX2_X1 U6791 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6847), .Z(n5510) );
  MUX2_X1 U6792 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6847), .Z(n5523) );
  MUX2_X1 U6793 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6847), .Z(n5536) );
  NOR2_X1 U6794 ( .A1(n5536), .A2(SI_16_), .ZN(n5246) );
  NAND2_X1 U6795 ( .A1(n5536), .A2(SI_16_), .ZN(n5247) );
  MUX2_X1 U6796 ( .A(n7299), .B(n5248), .S(n6847), .Z(n5249) );
  INV_X1 U6797 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6798 ( .A1(n5250), .A2(SI_17_), .ZN(n5251) );
  NAND2_X1 U6799 ( .A1(n5252), .A2(n5251), .ZN(n5550) );
  MUX2_X1 U6800 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6847), .Z(n5253) );
  INV_X1 U6801 ( .A(n5253), .ZN(n5254) );
  MUX2_X1 U6802 ( .A(n7532), .B(n10508), .S(n6847), .Z(n5257) );
  INV_X1 U6803 ( .A(n5257), .ZN(n5258) );
  NAND2_X1 U6804 ( .A1(n5258), .A2(SI_19_), .ZN(n5259) );
  NAND2_X1 U6805 ( .A1(n5260), .A2(n5259), .ZN(n5581) );
  MUX2_X1 U6806 ( .A(n7651), .B(n7633), .S(n6847), .Z(n5671) );
  OAI21_X1 U6807 ( .B1(n5675), .B2(n5672), .A(n5671), .ZN(n5262) );
  NAND2_X1 U6808 ( .A1(n5675), .A2(n5672), .ZN(n5261) );
  NAND2_X1 U6809 ( .A1(n5262), .A2(n5261), .ZN(n5662) );
  MUX2_X1 U6810 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6847), .Z(n5660) );
  NOR2_X1 U6811 ( .A1(n5660), .A2(SI_21_), .ZN(n5264) );
  NAND2_X1 U6812 ( .A1(n5660), .A2(SI_21_), .ZN(n5263) );
  MUX2_X1 U6813 ( .A(n7921), .B(n10278), .S(n6847), .Z(n5265) );
  INV_X1 U6814 ( .A(SI_22_), .ZN(n10484) );
  NAND2_X1 U6815 ( .A1(n5265), .A2(n10484), .ZN(n5268) );
  INV_X1 U6816 ( .A(n5265), .ZN(n5266) );
  NAND2_X1 U6817 ( .A1(n5266), .A2(SI_22_), .ZN(n5267) );
  NAND2_X1 U6818 ( .A1(n5268), .A2(n5267), .ZN(n5638) );
  INV_X1 U6819 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7930) );
  MUX2_X1 U6820 ( .A(n7930), .B(n10300), .S(n6847), .Z(n5269) );
  INV_X1 U6821 ( .A(SI_23_), .ZN(n10227) );
  NAND2_X1 U6822 ( .A1(n5269), .A2(n10227), .ZN(n5272) );
  INV_X1 U6823 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6824 ( .A1(n5270), .A2(SI_23_), .ZN(n5271) );
  INV_X1 U6825 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8026) );
  MUX2_X1 U6826 ( .A(n8026), .B(n10495), .S(n6847), .Z(n5273) );
  NAND2_X1 U6827 ( .A1(n5273), .A2(n10388), .ZN(n5276) );
  INV_X1 U6828 ( .A(n5273), .ZN(n5274) );
  NAND2_X1 U6829 ( .A1(n5274), .A2(SI_24_), .ZN(n5275) );
  NAND2_X1 U6830 ( .A1(n5619), .A2(n5620), .ZN(n5277) );
  INV_X1 U6831 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9123) );
  INV_X1 U6832 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10221) );
  MUX2_X1 U6833 ( .A(n9123), .B(n10221), .S(n6847), .Z(n5278) );
  INV_X1 U6834 ( .A(SI_25_), .ZN(n10365) );
  NAND2_X1 U6835 ( .A1(n5278), .A2(n10365), .ZN(n5281) );
  INV_X1 U6836 ( .A(n5278), .ZN(n5279) );
  NAND2_X1 U6837 ( .A1(n5279), .A2(SI_25_), .ZN(n5280) );
  INV_X1 U6838 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9119) );
  INV_X1 U6839 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10246) );
  MUX2_X1 U6840 ( .A(n9119), .B(n10246), .S(n6847), .Z(n5282) );
  INV_X1 U6841 ( .A(SI_26_), .ZN(n10404) );
  NAND2_X1 U6842 ( .A1(n5282), .A2(n10404), .ZN(n5285) );
  INV_X1 U6843 ( .A(n5282), .ZN(n5283) );
  NAND2_X1 U6844 ( .A1(n5283), .A2(SI_26_), .ZN(n5284) );
  NAND2_X1 U6845 ( .A1(n5286), .A2(n5285), .ZN(n5610) );
  INV_X1 U6846 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6121) );
  INV_X1 U6847 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10265) );
  MUX2_X1 U6848 ( .A(n6121), .B(n10265), .S(n6847), .Z(n5287) );
  INV_X1 U6849 ( .A(SI_27_), .ZN(n10379) );
  NAND2_X1 U6850 ( .A1(n5287), .A2(n10379), .ZN(n5290) );
  INV_X1 U6851 ( .A(n5287), .ZN(n5288) );
  NAND2_X1 U6852 ( .A1(n5288), .A2(SI_27_), .ZN(n5289) );
  INV_X1 U6853 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6133) );
  INV_X1 U6854 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10244) );
  MUX2_X1 U6855 ( .A(n6133), .B(n10244), .S(n6847), .Z(n5291) );
  INV_X1 U6856 ( .A(SI_28_), .ZN(n10520) );
  NAND2_X1 U6857 ( .A1(n5291), .A2(n10520), .ZN(n5294) );
  INV_X1 U6858 ( .A(n5291), .ZN(n5292) );
  NAND2_X1 U6859 ( .A1(n5292), .A2(SI_28_), .ZN(n5293) );
  MUX2_X1 U6860 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6847), .Z(n5296) );
  NAND2_X1 U6861 ( .A1(n4992), .A2(n5296), .ZN(n5297) );
  MUX2_X1 U6862 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6847), .Z(n5719) );
  XNOR2_X1 U6863 ( .A(n5719), .B(SI_30_), .ZN(n5720) );
  MUX2_X1 U6864 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5299), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5301) );
  NAND2_X1 U6865 ( .A1(n8344), .A2(n5726), .ZN(n5304) );
  INV_X1 U6866 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10522) );
  OR2_X1 U6867 ( .A1(n5728), .A2(n10522), .ZN(n5303) );
  INV_X1 U6868 ( .A(n9828), .ZN(n5879) );
  NAND2_X1 U6869 ( .A1(n5709), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6870 ( .A1(n5354), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5307) );
  INV_X1 U6871 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6842) );
  INV_X1 U6872 ( .A(n5309), .ZN(n5310) );
  NAND2_X1 U6873 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  NAND2_X1 U6874 ( .A1(n5313), .A2(n5312), .ZN(n6853) );
  NAND2_X1 U6875 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5314) );
  MUX2_X1 U6876 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5314), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5317) );
  INV_X1 U6877 ( .A(n5334), .ZN(n5316) );
  NAND2_X1 U6878 ( .A1(n5317), .A2(n5316), .ZN(n6911) );
  INV_X1 U6879 ( .A(n6911), .ZN(n9309) );
  NAND2_X1 U6880 ( .A1(n5708), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6881 ( .A1(n5707), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6882 ( .A1(n5709), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6883 ( .A1(n5354), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5318) );
  NAND4_X1 U6884 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), .ZN(n7038)
         );
  NAND2_X1 U6885 ( .A1(n6847), .A2(SI_0_), .ZN(n5322) );
  XNOR2_X1 U6886 ( .A(n5322), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9886) );
  MUX2_X1 U6887 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9886), .S(n6871), .Z(n7041) );
  NAND2_X1 U6888 ( .A1(n7024), .A2(n7023), .ZN(n5324) );
  INV_X1 U6889 ( .A(n4512), .ZN(n9889) );
  NAND2_X1 U6890 ( .A1(n9889), .A2(n4833), .ZN(n5323) );
  NAND2_X1 U6891 ( .A1(n5324), .A2(n5323), .ZN(n7155) );
  NAND2_X1 U6892 ( .A1(n5709), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6893 ( .A1(n5707), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6894 ( .A1(n5354), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5326) );
  INV_X1 U6895 ( .A(n5329), .ZN(n5331) );
  NAND2_X1 U6896 ( .A1(n5331), .A2(n5330), .ZN(n5333) );
  NAND2_X1 U6897 ( .A1(n5333), .A2(n5332), .ZN(n6856) );
  OR2_X1 U6898 ( .A1(n5334), .A2(n4641), .ZN(n5366) );
  INV_X1 U6899 ( .A(n5366), .ZN(n5335) );
  NAND2_X1 U6900 ( .A1(n5335), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5337) );
  INV_X1 U6901 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6902 ( .A1(n5366), .A2(n5336), .ZN(n5348) );
  AND2_X1 U6903 ( .A1(n5337), .A2(n5348), .ZN(n7070) );
  INV_X1 U6904 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6845) );
  OR2_X1 U6905 ( .A1(n5728), .A2(n6845), .ZN(n5338) );
  NAND2_X1 U6906 ( .A1(n9305), .A2(n8338), .ZN(n7226) );
  INV_X4 U6907 ( .A(n5354), .ZN(n5372) );
  OR2_X1 U6908 ( .A1(n5372), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6909 ( .A1(n5707), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6910 ( .A1(n5708), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6911 ( .A1(n5709), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5340) );
  NAND4_X2 U6912 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n9304)
         );
  INV_X1 U6913 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6844) );
  OR2_X1 U6914 ( .A1(n5728), .A2(n6844), .ZN(n5352) );
  OR2_X1 U6915 ( .A1(n5345), .A2(n5344), .ZN(n5346) );
  NAND2_X1 U6916 ( .A1(n5347), .A2(n5346), .ZN(n6854) );
  OR2_X1 U6917 ( .A1(n5706), .A2(n6854), .ZN(n5351) );
  NAND2_X1 U6918 ( .A1(n5348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5349) );
  XNOR2_X1 U6919 ( .A(n5349), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9327) );
  NAND2_X1 U6920 ( .A1(n5586), .A2(n9327), .ZN(n5350) );
  NAND2_X1 U6921 ( .A1(n9304), .A2(n7421), .ZN(n5353) );
  AND2_X1 U6922 ( .A1(n7226), .A2(n5353), .ZN(n5893) );
  INV_X1 U6923 ( .A(n9304), .ZN(n6016) );
  INV_X1 U6924 ( .A(n7421), .ZN(n7395) );
  NAND2_X1 U6925 ( .A1(n5709), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6926 ( .A1(n5707), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5358) );
  NOR2_X1 U6927 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5355) );
  NOR2_X1 U6928 ( .A1(n5373), .A2(n5355), .ZN(n7413) );
  NAND2_X1 U6929 ( .A1(n5354), .A2(n7413), .ZN(n5357) );
  NAND2_X1 U6930 ( .A1(n5708), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5356) );
  NAND4_X1 U6931 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .ZN(n9303)
         );
  OR2_X1 U6932 ( .A1(n5728), .A2(n5204), .ZN(n5370) );
  OR2_X1 U6933 ( .A1(n5361), .A2(n5360), .ZN(n5362) );
  NAND2_X1 U6934 ( .A1(n5363), .A2(n5362), .ZN(n6858) );
  OR2_X1 U6935 ( .A1(n5706), .A2(n6858), .ZN(n5369) );
  OR2_X1 U6936 ( .A1(n5364), .A2(n4641), .ZN(n5365) );
  NAND2_X1 U6937 ( .A1(n5366), .A2(n5365), .ZN(n5379) );
  INV_X1 U6938 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5367) );
  XNOR2_X1 U6939 ( .A(n5379), .B(n5367), .ZN(n7051) );
  NAND2_X1 U6940 ( .A1(n5586), .A2(n7051), .ZN(n5368) );
  NAND2_X1 U6941 ( .A1(n9303), .A2(n9957), .ZN(n5891) );
  OR2_X1 U6942 ( .A1(n9303), .A2(n9957), .ZN(n5770) );
  NAND2_X1 U6943 ( .A1(n5709), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5378) );
  INV_X1 U6944 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5371) );
  OR2_X1 U6945 ( .A1(n5656), .A2(n5371), .ZN(n5377) );
  NAND2_X1 U6946 ( .A1(n5373), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5390) );
  OAI21_X1 U6947 ( .B1(n5373), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5390), .ZN(
        n7581) );
  OR2_X1 U6948 ( .A1(n5372), .A2(n7581), .ZN(n5376) );
  INV_X1 U6949 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5374) );
  OR2_X1 U6950 ( .A1(n5614), .A2(n5374), .ZN(n5375) );
  OAI21_X1 U6951 ( .B1(n5379), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5381) );
  INV_X1 U6952 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5380) );
  XNOR2_X1 U6953 ( .A(n5381), .B(n5380), .ZN(n9335) );
  OR2_X1 U6954 ( .A1(n5383), .A2(n5382), .ZN(n5384) );
  NAND2_X1 U6955 ( .A1(n5385), .A2(n5384), .ZN(n6849) );
  OR2_X1 U6956 ( .A1(n5706), .A2(n6849), .ZN(n5387) );
  INV_X1 U6957 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6846) );
  OR2_X1 U6958 ( .A1(n5728), .A2(n6846), .ZN(n5386) );
  OAI211_X1 U6959 ( .C1(n6871), .C2(n9335), .A(n5387), .B(n5386), .ZN(n7578)
         );
  NAND2_X1 U6960 ( .A1(n7572), .A2(n7578), .ZN(n5771) );
  NAND2_X1 U6961 ( .A1(n5771), .A2(n5897), .ZN(n7379) );
  NAND2_X1 U6962 ( .A1(n5769), .A2(n5100), .ZN(n5388) );
  NAND2_X1 U6963 ( .A1(n5388), .A2(n5771), .ZN(n7466) );
  INV_X1 U6964 ( .A(n7466), .ZN(n5405) );
  NAND2_X1 U6965 ( .A1(n5709), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6966 ( .A1(n5707), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5394) );
  INV_X1 U6967 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5389) );
  NOR2_X1 U6968 ( .A1(n5390), .A2(n5389), .ZN(n5432) );
  AND2_X1 U6969 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  NOR2_X1 U6970 ( .A1(n5432), .A2(n5391), .ZN(n7473) );
  NAND2_X1 U6971 ( .A1(n5354), .A2(n7473), .ZN(n5393) );
  NAND2_X1 U6972 ( .A1(n5708), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5392) );
  NAND4_X1 U6973 ( .A1(n5395), .A2(n5394), .A3(n5393), .A4(n5392), .ZN(n9301)
         );
  OR2_X1 U6974 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  NAND2_X1 U6975 ( .A1(n5399), .A2(n5398), .ZN(n6852) );
  OR2_X1 U6976 ( .A1(n6852), .A2(n5706), .ZN(n5404) );
  NAND2_X1 U6977 ( .A1(n5400), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5401) );
  XNOR2_X1 U6978 ( .A(n5401), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U6979 ( .A1(n5586), .A2(n6920), .ZN(n5403) );
  INV_X1 U6980 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6851) );
  OR2_X1 U6981 ( .A1(n5728), .A2(n6851), .ZN(n5402) );
  OR2_X1 U6982 ( .A1(n9301), .A2(n7674), .ZN(n5900) );
  INV_X1 U6983 ( .A(n5900), .ZN(n5772) );
  XNOR2_X1 U6984 ( .A(n5407), .B(n5406), .ZN(n6873) );
  NAND2_X1 U6985 ( .A1(n6873), .A2(n5726), .ZN(n5414) );
  NOR2_X1 U6986 ( .A1(n5409), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5455) );
  OR2_X1 U6987 ( .A1(n5455), .A2(n4641), .ZN(n5424) );
  INV_X1 U6988 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U6989 ( .A1(n5424), .A2(n5410), .ZN(n5411) );
  NAND2_X1 U6990 ( .A1(n5411), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5412) );
  XNOR2_X1 U6991 ( .A(n5412), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U6992 ( .A1(n5587), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5586), .B2(
        n6950), .ZN(n5413) );
  NAND2_X1 U6993 ( .A1(n5414), .A2(n5413), .ZN(n7987) );
  NAND2_X1 U6994 ( .A1(n5707), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5421) );
  INV_X1 U6995 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7644) );
  OR2_X1 U6996 ( .A1(n5605), .A2(n7644), .ZN(n5420) );
  NAND2_X1 U6997 ( .A1(n5432), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5434) );
  INV_X1 U6998 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5427) );
  INV_X1 U6999 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5415) );
  OAI21_X1 U7000 ( .B1(n5434), .B2(n5427), .A(n5415), .ZN(n5417) );
  NAND2_X1 U7001 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n5416) );
  NAND2_X1 U7002 ( .A1(n5417), .A2(n5459), .ZN(n7998) );
  OR2_X1 U7003 ( .A1(n5372), .A2(n7998), .ZN(n5419) );
  INV_X1 U7004 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6904) );
  OR2_X1 U7005 ( .A1(n5614), .A2(n6904), .ZN(n5418) );
  NAND2_X1 U7006 ( .A1(n7987), .A2(n7985), .ZN(n5799) );
  XNOR2_X1 U7007 ( .A(n5423), .B(n5422), .ZN(n6862) );
  NAND2_X1 U7008 ( .A1(n6862), .A2(n5726), .ZN(n5426) );
  XNOR2_X1 U7009 ( .A(n5424), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6944) );
  AOI22_X1 U7010 ( .A1(n5587), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5586), .B2(
        n6944), .ZN(n5425) );
  NAND2_X1 U7011 ( .A1(n5426), .A2(n5425), .ZN(n9921) );
  NAND2_X1 U7012 ( .A1(n5707), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5431) );
  INV_X1 U7013 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7662) );
  OR2_X1 U7014 ( .A1(n5605), .A2(n7662), .ZN(n5430) );
  XNOR2_X1 U7015 ( .A(n5434), .B(n5427), .ZN(n9924) );
  OR2_X1 U7016 ( .A1(n5372), .A2(n9924), .ZN(n5429) );
  INV_X1 U7017 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6936) );
  OR2_X1 U7018 ( .A1(n5614), .A2(n6936), .ZN(n5428) );
  NAND2_X1 U7019 ( .A1(n9921), .A2(n7999), .ZN(n7636) );
  OR2_X1 U7020 ( .A1(n5432), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U7021 ( .A1(n5434), .A2(n5433), .ZN(n7743) );
  OR2_X1 U7022 ( .A1(n5372), .A2(n7743), .ZN(n5438) );
  NAND2_X1 U7023 ( .A1(n5709), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U7024 ( .A1(n5707), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U7025 ( .A1(n5708), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5435) );
  NAND4_X1 U7026 ( .A1(n5438), .A2(n5437), .A3(n5436), .A4(n5435), .ZN(n9300)
         );
  INV_X1 U7027 ( .A(n9300), .ZN(n7467) );
  NAND2_X1 U7028 ( .A1(n5409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5443) );
  XNOR2_X1 U7029 ( .A(n5443), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9372) );
  AOI22_X1 U7030 ( .A1(n5587), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5586), .B2(
        n9372), .ZN(n5444) );
  AND2_X2 U7031 ( .A1(n5445), .A2(n5444), .ZN(n7630) );
  INV_X1 U7032 ( .A(n7630), .ZN(n7745) );
  NAND2_X1 U7033 ( .A1(n7467), .A2(n7745), .ZN(n7634) );
  NAND2_X1 U7034 ( .A1(n7636), .A2(n7634), .ZN(n5446) );
  INV_X1 U7035 ( .A(n5446), .ZN(n5787) );
  NAND2_X1 U7036 ( .A1(n5799), .A2(n5787), .ZN(n5449) );
  OR2_X1 U7037 ( .A1(n7987), .A2(n7985), .ZN(n5798) );
  OR2_X1 U7038 ( .A1(n9921), .A2(n7999), .ZN(n7637) );
  NAND2_X1 U7039 ( .A1(n7630), .A2(n9300), .ZN(n5777) );
  AND2_X1 U7040 ( .A1(n7637), .A2(n5777), .ZN(n5788) );
  NAND2_X1 U7041 ( .A1(n9301), .A2(n7674), .ZN(n7539) );
  AND3_X1 U7042 ( .A1(n5798), .A2(n5788), .A3(n7539), .ZN(n5448) );
  NAND3_X1 U7043 ( .A1(n5798), .A2(n5446), .A3(n7637), .ZN(n5447) );
  NAND2_X1 U7044 ( .A1(n5447), .A2(n5799), .ZN(n5899) );
  OR2_X1 U7045 ( .A1(n5448), .A2(n5899), .ZN(n5903) );
  NAND2_X1 U7046 ( .A1(n5451), .A2(n5450), .ZN(n5452) );
  NAND2_X1 U7047 ( .A1(n5453), .A2(n5452), .ZN(n6879) );
  OR2_X1 U7048 ( .A1(n6879), .A2(n5706), .ZN(n5458) );
  NOR2_X1 U7049 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5454) );
  NAND2_X1 U7050 ( .A1(n5455), .A2(n5454), .ZN(n5468) );
  NAND2_X1 U7051 ( .A1(n5468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5456) );
  XNOR2_X1 U7052 ( .A(n5456), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6957) );
  AOI22_X1 U7053 ( .A1(n5587), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5586), .B2(
        n6957), .ZN(n5457) );
  NAND2_X1 U7054 ( .A1(n5458), .A2(n5457), .ZN(n8109) );
  NAND2_X1 U7055 ( .A1(n5707), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5464) );
  INV_X1 U7056 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7780) );
  OR2_X1 U7057 ( .A1(n5605), .A2(n7780), .ZN(n5463) );
  AND2_X1 U7058 ( .A1(n5459), .A2(n9378), .ZN(n5460) );
  OR2_X1 U7059 ( .A1(n5460), .A2(n5472), .ZN(n9909) );
  OR2_X1 U7060 ( .A1(n5372), .A2(n9909), .ZN(n5462) );
  INV_X1 U7061 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6958) );
  OR2_X1 U7062 ( .A1(n5614), .A2(n6958), .ZN(n5461) );
  OR2_X1 U7063 ( .A1(n8109), .A2(n8123), .ZN(n5904) );
  NAND2_X1 U7064 ( .A1(n8109), .A2(n8123), .ZN(n7946) );
  NAND2_X1 U7065 ( .A1(n5904), .A2(n7946), .ZN(n7776) );
  XNOR2_X1 U7066 ( .A(n5467), .B(n5466), .ZN(n6884) );
  NAND2_X1 U7067 ( .A1(n6884), .A2(n5726), .ZN(n5471) );
  NAND2_X1 U7068 ( .A1(n5483), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5469) );
  XNOR2_X1 U7069 ( .A(n5469), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6955) );
  AOI22_X1 U7070 ( .A1(n5587), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5586), .B2(
        n6955), .ZN(n5470) );
  NOR2_X1 U7071 ( .A1(n5472), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5473) );
  OR2_X1 U7072 ( .A1(n5486), .A2(n5473), .ZN(n7944) );
  OR2_X1 U7073 ( .A1(n5372), .A2(n7944), .ZN(n5477) );
  NAND2_X1 U7074 ( .A1(n5707), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U7075 ( .A1(n5708), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7076 ( .A1(n5709), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5474) );
  NAND4_X1 U7077 ( .A1(n5477), .A2(n5476), .A3(n5475), .A4(n5474), .ZN(n9296)
         );
  INV_X1 U7078 ( .A(n9296), .ZN(n9180) );
  OR2_X1 U7079 ( .A1(n8115), .A2(n9180), .ZN(n5804) );
  NAND2_X1 U7080 ( .A1(n8115), .A2(n9180), .ZN(n5802) );
  NAND2_X1 U7081 ( .A1(n5804), .A2(n5802), .ZN(n7951) );
  INV_X1 U7082 ( .A(n7946), .ZN(n5794) );
  NOR2_X1 U7083 ( .A1(n7951), .A2(n5794), .ZN(n5478) );
  NAND2_X1 U7084 ( .A1(n7947), .A2(n5478), .ZN(n7948) );
  NAND2_X1 U7085 ( .A1(n7948), .A2(n5804), .ZN(n7905) );
  INV_X1 U7086 ( .A(n7905), .ZN(n5493) );
  NAND2_X1 U7087 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  AND2_X1 U7088 ( .A1(n5482), .A2(n5481), .ZN(n6968) );
  NAND2_X1 U7089 ( .A1(n6968), .A2(n5726), .ZN(n5485) );
  OAI21_X1 U7090 ( .B1(n5483), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5500) );
  XNOR2_X1 U7091 ( .A(n5500), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7323) );
  AOI22_X1 U7092 ( .A1(n5587), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5586), .B2(
        n7323), .ZN(n5484) );
  OR2_X1 U7093 ( .A1(n5486), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7094 ( .A1(n5517), .A2(n5487), .ZN(n9178) );
  OR2_X1 U7095 ( .A1(n5372), .A2(n9178), .ZN(n5491) );
  NAND2_X1 U7096 ( .A1(n5707), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U7097 ( .A1(n5708), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7098 ( .A1(n5709), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5488) );
  NAND4_X1 U7099 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n9295)
         );
  XNOR2_X1 U7100 ( .A(n8221), .B(n6023), .ZN(n7904) );
  NAND2_X1 U7101 ( .A1(n5493), .A2(n5492), .ZN(n7907) );
  NAND2_X1 U7102 ( .A1(n8221), .A2(n6023), .ZN(n5910) );
  INV_X1 U7103 ( .A(n5494), .ZN(n5496) );
  NAND2_X1 U7104 ( .A1(n5496), .A2(n5495), .ZN(n5498) );
  NAND2_X1 U7105 ( .A1(n5498), .A2(n5497), .ZN(n6979) );
  OR2_X1 U7106 ( .A1(n6979), .A2(n5706), .ZN(n5504) );
  INV_X1 U7107 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U7108 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  NAND2_X1 U7109 ( .A1(n5501), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5502) );
  XNOR2_X1 U7110 ( .A(n5502), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7330) );
  AOI22_X1 U7111 ( .A1(n5587), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5586), .B2(
        n7330), .ZN(n5503) );
  NAND2_X1 U7112 ( .A1(n5709), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7113 ( .A1(n5707), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5507) );
  XNOR2_X1 U7114 ( .A(n5517), .B(P1_REG3_REG_13__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U7115 ( .A1(n5354), .A2(n9237), .ZN(n5506) );
  NAND2_X1 U7116 ( .A1(n5708), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5505) );
  NAND4_X1 U7117 ( .A1(n5508), .A2(n5507), .A3(n5506), .A4(n5505), .ZN(n9294)
         );
  XNOR2_X1 U7118 ( .A(n8212), .B(n9179), .ZN(n8014) );
  NAND2_X1 U7119 ( .A1(n9240), .A2(n9294), .ZN(n5913) );
  XNOR2_X1 U7120 ( .A(n5510), .B(SI_14_), .ZN(n5511) );
  XNOR2_X1 U7121 ( .A(n5509), .B(n5511), .ZN(n7016) );
  NAND2_X1 U7122 ( .A1(n7016), .A2(n5726), .ZN(n5515) );
  OR2_X1 U7123 ( .A1(n5512), .A2(n4641), .ZN(n5513) );
  XNOR2_X1 U7124 ( .A(n5513), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7327) );
  AOI22_X1 U7125 ( .A1(n5587), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5586), .B2(
        n7327), .ZN(n5514) );
  INV_X1 U7126 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5516) );
  OAI21_X1 U7127 ( .B1(n5517), .B2(n5516), .A(n9130), .ZN(n5518) );
  NAND2_X1 U7128 ( .A1(n5518), .A2(n5529), .ZN(n9131) );
  OR2_X1 U7129 ( .A1(n5372), .A2(n9131), .ZN(n5522) );
  NAND2_X1 U7130 ( .A1(n5707), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7131 ( .A1(n5709), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7132 ( .A1(n5708), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5519) );
  NAND4_X1 U7133 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), .ZN(n9726)
         );
  OR2_X1 U7134 ( .A1(n9134), .A2(n9280), .ZN(n5916) );
  NAND2_X1 U7135 ( .A1(n9134), .A2(n9280), .ZN(n5817) );
  NAND2_X1 U7136 ( .A1(n5916), .A2(n5817), .ZN(n8147) );
  XNOR2_X1 U7137 ( .A(n5523), .B(SI_15_), .ZN(n5524) );
  XNOR2_X1 U7138 ( .A(n5525), .B(n5524), .ZN(n7162) );
  NAND2_X1 U7139 ( .A1(n7162), .A2(n5726), .ZN(n5528) );
  NAND2_X1 U7140 ( .A1(n5526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5555) );
  XNOR2_X1 U7141 ( .A(n5555), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7555) );
  AOI22_X1 U7142 ( .A1(n5587), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5586), .B2(
        n7555), .ZN(n5527) );
  INV_X1 U7143 ( .A(n5544), .ZN(n5531) );
  NAND2_X1 U7144 ( .A1(n5529), .A2(n9277), .ZN(n5530) );
  NAND2_X1 U7145 ( .A1(n5531), .A2(n5530), .ZN(n9735) );
  OR2_X1 U7146 ( .A1(n5372), .A2(n9735), .ZN(n5535) );
  NAND2_X1 U7147 ( .A1(n5709), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7148 ( .A1(n5707), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7149 ( .A1(n5708), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5532) );
  NAND4_X1 U7150 ( .A1(n5535), .A2(n5534), .A3(n5533), .A4(n5532), .ZN(n9701)
         );
  INV_X1 U7151 ( .A(n9701), .ZN(n9199) );
  OR2_X1 U7152 ( .A1(n9734), .A2(n9199), .ZN(n5768) );
  NAND2_X1 U7153 ( .A1(n9734), .A2(n9199), .ZN(n5821) );
  NAND2_X1 U7154 ( .A1(n9722), .A2(n9723), .ZN(n9721) );
  NAND2_X1 U7155 ( .A1(n9721), .A2(n5821), .ZN(n9699) );
  INV_X1 U7156 ( .A(n5536), .ZN(n5537) );
  XNOR2_X1 U7157 ( .A(n5537), .B(SI_16_), .ZN(n5538) );
  XNOR2_X1 U7158 ( .A(n5539), .B(n5538), .ZN(n7197) );
  NAND2_X1 U7159 ( .A1(n7197), .A2(n5726), .ZN(n5543) );
  NAND2_X1 U7160 ( .A1(n5555), .A2(n4919), .ZN(n5540) );
  NAND2_X1 U7161 ( .A1(n5540), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5541) );
  XNOR2_X1 U7162 ( .A(n5541), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7833) );
  AOI22_X1 U7163 ( .A1(n5587), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5586), .B2(
        n7833), .ZN(n5542) );
  NAND2_X1 U7164 ( .A1(n5707), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5549) );
  INV_X1 U7165 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9713) );
  OR2_X1 U7166 ( .A1(n5605), .A2(n9713), .ZN(n5548) );
  NAND2_X1 U7167 ( .A1(n5544), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5560) );
  OR2_X1 U7168 ( .A1(n5544), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U7169 ( .A1(n5560), .A2(n5545), .ZN(n9712) );
  OR2_X1 U7170 ( .A1(n5372), .A2(n9712), .ZN(n5547) );
  INV_X1 U7171 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7839) );
  OR2_X1 U7172 ( .A1(n5614), .A2(n7839), .ZN(n5546) );
  NAND2_X1 U7173 ( .A1(n9812), .A2(n9278), .ZN(n5918) );
  NAND2_X1 U7174 ( .A1(n5829), .A2(n5918), .ZN(n9704) );
  INV_X1 U7175 ( .A(n9704), .ZN(n9700) );
  NAND2_X1 U7176 ( .A1(n9699), .A2(n9700), .ZN(n9698) );
  NAND2_X1 U7177 ( .A1(n9698), .A2(n5918), .ZN(n9683) );
  INV_X1 U7178 ( .A(n9683), .ZN(n5567) );
  XNOR2_X1 U7179 ( .A(n5551), .B(n5550), .ZN(n7236) );
  NAND2_X1 U7180 ( .A1(n7236), .A2(n5726), .ZN(n5558) );
  INV_X1 U7181 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U7182 ( .A1(n5553), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5554) );
  XNOR2_X1 U7183 ( .A(n5569), .B(n5556), .ZN(n9433) );
  AOI22_X1 U7184 ( .A1(n5587), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5586), .B2(
        n9433), .ZN(n5557) );
  NAND2_X1 U7185 ( .A1(n5707), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5565) );
  INV_X1 U7186 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9692) );
  OR2_X1 U7187 ( .A1(n5605), .A2(n9692), .ZN(n5564) );
  INV_X1 U7188 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7189 ( .A1(n5560), .A2(n5559), .ZN(n5561) );
  NAND2_X1 U7190 ( .A1(n5573), .A2(n5561), .ZN(n9691) );
  OR2_X1 U7191 ( .A1(n5372), .A2(n9691), .ZN(n5563) );
  INV_X1 U7192 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9809) );
  OR2_X1 U7193 ( .A1(n5614), .A2(n9809), .ZN(n5562) );
  OR2_X1 U7194 ( .A1(n9690), .A2(n9256), .ZN(n5767) );
  NAND2_X1 U7195 ( .A1(n9690), .A2(n9256), .ZN(n5833) );
  NAND2_X1 U7196 ( .A1(n5767), .A2(n5833), .ZN(n9682) );
  NAND2_X1 U7197 ( .A1(n5567), .A2(n5566), .ZN(n9685) );
  XNOR2_X1 U7198 ( .A(n5568), .B(n4579), .ZN(n7451) );
  NAND2_X1 U7199 ( .A1(n7451), .A2(n5726), .ZN(n5571) );
  XNOR2_X1 U7200 ( .A(n5583), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9454) );
  AOI22_X1 U7201 ( .A1(n5587), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5586), .B2(
        n9454), .ZN(n5570) );
  NAND2_X1 U7202 ( .A1(n5709), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5579) );
  INV_X1 U7203 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n5572) );
  OR2_X1 U7204 ( .A1(n5656), .A2(n5572), .ZN(n5578) );
  AND2_X1 U7205 ( .A1(n5573), .A2(n9255), .ZN(n5574) );
  OR2_X1 U7206 ( .A1(n5574), .A2(n5590), .ZN(n9671) );
  OR2_X1 U7207 ( .A1(n5372), .A2(n9671), .ZN(n5577) );
  INV_X1 U7208 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n5575) );
  OR2_X1 U7209 ( .A1(n5614), .A2(n5575), .ZN(n5576) );
  OR2_X1 U7210 ( .A1(n4719), .A2(n9661), .ZN(n5832) );
  NAND2_X1 U7211 ( .A1(n4719), .A2(n9661), .ZN(n5834) );
  XNOR2_X1 U7212 ( .A(n5580), .B(n5581), .ZN(n7530) );
  NAND2_X1 U7213 ( .A1(n7530), .A2(n5726), .ZN(n5589) );
  XNOR2_X2 U7214 ( .A(n5585), .B(n5584), .ZN(n7033) );
  INV_X1 U7215 ( .A(n7033), .ZN(n6001) );
  AOI22_X1 U7216 ( .A1(n5587), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6001), .B2(
        n5586), .ZN(n5588) );
  NAND2_X1 U7217 ( .A1(n5707), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5595) );
  INV_X1 U7218 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9654) );
  OR2_X1 U7219 ( .A1(n5605), .A2(n9654), .ZN(n5594) );
  NOR2_X1 U7220 ( .A1(n5590), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5591) );
  OR2_X1 U7221 ( .A1(n5678), .A2(n5591), .ZN(n9653) );
  OR2_X1 U7222 ( .A1(n5372), .A2(n9653), .ZN(n5593) );
  INV_X1 U7223 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9457) );
  OR2_X1 U7224 ( .A1(n5614), .A2(n9457), .ZN(n5592) );
  NAND2_X1 U7225 ( .A1(n9798), .A2(n9292), .ZN(n5925) );
  NAND2_X1 U7226 ( .A1(n5837), .A2(n5925), .ZN(n9657) );
  INV_X1 U7227 ( .A(n9637), .ZN(n5716) );
  NAND2_X1 U7228 ( .A1(n6132), .A2(n5726), .ZN(n5600) );
  OR2_X1 U7229 ( .A1(n5728), .A2(n10244), .ZN(n5599) );
  NAND2_X1 U7230 ( .A1(n5707), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5609) );
  INV_X1 U7231 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5601) );
  OR2_X1 U7232 ( .A1(n5614), .A2(n5601), .ZN(n5608) );
  INV_X1 U7233 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9168) );
  INV_X1 U7234 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9245) );
  INV_X1 U7235 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9138) );
  INV_X1 U7236 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U7237 ( .A1(n5602), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9485) );
  INV_X1 U7238 ( .A(n5602), .ZN(n5603) );
  INV_X1 U7239 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U7240 ( .A1(n5603), .A2(n9157), .ZN(n5604) );
  NAND2_X1 U7241 ( .A1(n9485), .A2(n5604), .ZN(n9510) );
  OR2_X1 U7242 ( .A1(n5372), .A2(n9510), .ZN(n5607) );
  INV_X1 U7243 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9511) );
  OR2_X1 U7244 ( .A1(n5605), .A2(n9511), .ZN(n5606) );
  NAND2_X1 U7245 ( .A1(n9752), .A2(n9525), .ZN(n5998) );
  NAND2_X1 U7246 ( .A1(n9113), .A2(n5726), .ZN(n5613) );
  OR2_X1 U7247 ( .A1(n5728), .A2(n10265), .ZN(n5612) );
  NAND2_X1 U7248 ( .A1(n5709), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5618) );
  INV_X1 U7249 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9831) );
  OR2_X1 U7250 ( .A1(n5656), .A2(n9831), .ZN(n5617) );
  XNOR2_X1 U7251 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n5692), .ZN(n9518) );
  OR2_X1 U7252 ( .A1(n5372), .A2(n9518), .ZN(n5616) );
  INV_X1 U7253 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9759) );
  OR2_X1 U7254 ( .A1(n5614), .A2(n9759), .ZN(n5615) );
  NAND2_X1 U7255 ( .A1(n9529), .A2(n9537), .ZN(n5997) );
  NAND2_X1 U7256 ( .A1(n5998), .A2(n5997), .ZN(n5859) );
  XNOR2_X1 U7257 ( .A(n5619), .B(n5620), .ZN(n8025) );
  NAND2_X1 U7258 ( .A1(n8025), .A2(n5726), .ZN(n5622) );
  OR2_X1 U7259 ( .A1(n5728), .A2(n10495), .ZN(n5621) );
  NOR2_X1 U7260 ( .A1(n5634), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5623) );
  OR2_X1 U7261 ( .A1(n5652), .A2(n5623), .ZN(n9218) );
  INV_X1 U7262 ( .A(n9218), .ZN(n9573) );
  NAND2_X1 U7263 ( .A1(n9573), .A2(n5354), .ZN(n5629) );
  INV_X1 U7264 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7265 ( .A1(n5709), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7266 ( .A1(n5708), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5624) );
  OAI211_X1 U7267 ( .C1(n5656), .C2(n5626), .A(n5625), .B(n5624), .ZN(n5627)
         );
  INV_X1 U7268 ( .A(n5627), .ZN(n5628) );
  NAND2_X1 U7269 ( .A1(n9773), .A2(n9585), .ZN(n5856) );
  XNOR2_X1 U7270 ( .A(n5631), .B(n5630), .ZN(n7927) );
  NAND2_X1 U7271 ( .A1(n7927), .A2(n5726), .ZN(n5633) );
  OR2_X1 U7272 ( .A1(n5728), .A2(n10300), .ZN(n5632) );
  AND2_X1 U7273 ( .A1(n5643), .A2(n9138), .ZN(n5635) );
  OR2_X1 U7274 ( .A1(n5635), .A2(n5634), .ZN(n9591) );
  AOI22_X1 U7275 ( .A1(n5707), .A2(P1_REG0_REG_23__SCAN_IN), .B1(n5709), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7276 ( .A1(n5708), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5636) );
  OAI211_X1 U7277 ( .C1(n9591), .C2(n5372), .A(n5637), .B(n5636), .ZN(n9609)
         );
  NAND2_X1 U7278 ( .A1(n9590), .A2(n9569), .ZN(n9565) );
  OR2_X1 U7279 ( .A1(n9590), .A2(n9569), .ZN(n5851) );
  XNOR2_X1 U7280 ( .A(n5639), .B(n5638), .ZN(n7918) );
  NAND2_X1 U7281 ( .A1(n7918), .A2(n5726), .ZN(n5641) );
  OR2_X1 U7282 ( .A1(n5728), .A2(n10278), .ZN(n5640) );
  NAND2_X1 U7283 ( .A1(n5666), .A2(n9245), .ZN(n5642) );
  NAND2_X1 U7284 ( .A1(n5643), .A2(n5642), .ZN(n9602) );
  AOI22_X1 U7285 ( .A1(n5707), .A2(P1_REG0_REG_22__SCAN_IN), .B1(n5708), .B2(
        P1_REG1_REG_22__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7286 ( .A1(n5709), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5644) );
  OAI211_X1 U7287 ( .C1(n9602), .C2(n5372), .A(n5645), .B(n5644), .ZN(n9290)
         );
  INV_X1 U7288 ( .A(n9290), .ZN(n9584) );
  OR2_X1 U7289 ( .A1(n9782), .A2(n9584), .ZN(n5646) );
  NAND2_X1 U7290 ( .A1(n5851), .A2(n5646), .ZN(n5844) );
  NAND3_X1 U7291 ( .A1(n5856), .A2(n9565), .A3(n5844), .ZN(n5647) );
  AND2_X1 U7292 ( .A1(n5647), .A2(n5992), .ZN(n5658) );
  NAND2_X1 U7293 ( .A1(n9121), .A2(n5726), .ZN(n5651) );
  OR2_X1 U7294 ( .A1(n5728), .A2(n10221), .ZN(n5650) );
  INV_X1 U7295 ( .A(n9838), .ZN(n9557) );
  OR2_X1 U7296 ( .A1(n5652), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5653) );
  INV_X1 U7297 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U7298 ( .A1(n5709), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7299 ( .A1(n5708), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5654) );
  OAI211_X1 U7300 ( .C1(n5656), .C2(n9836), .A(n5655), .B(n5654), .ZN(n5657)
         );
  OR2_X1 U7301 ( .A1(n9557), .A2(n9570), .ZN(n5996) );
  NAND2_X1 U7302 ( .A1(n5658), .A2(n5996), .ZN(n5701) );
  NAND2_X1 U7303 ( .A1(n9782), .A2(n9584), .ZN(n5990) );
  AND2_X1 U7304 ( .A1(n9565), .A2(n5990), .ZN(n5842) );
  INV_X1 U7305 ( .A(SI_21_), .ZN(n5659) );
  XNOR2_X1 U7306 ( .A(n5660), .B(n5659), .ZN(n5661) );
  XNOR2_X1 U7307 ( .A(n5662), .B(n5661), .ZN(n7786) );
  NAND2_X1 U7308 ( .A1(n7786), .A2(n5726), .ZN(n5664) );
  INV_X1 U7309 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7809) );
  OR2_X1 U7310 ( .A1(n5728), .A2(n7809), .ZN(n5663) );
  NAND2_X1 U7311 ( .A1(n5680), .A2(n9168), .ZN(n5665) );
  NAND2_X1 U7312 ( .A1(n5666), .A2(n5665), .ZN(n9627) );
  OR2_X1 U7313 ( .A1(n9627), .A2(n5372), .ZN(n5670) );
  NAND2_X1 U7314 ( .A1(n5709), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7315 ( .A1(n5707), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7316 ( .A1(n5708), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7317 ( .A1(n9626), .A2(n9246), .ZN(n5989) );
  INV_X1 U7318 ( .A(n5671), .ZN(n5673) );
  XNOR2_X1 U7319 ( .A(n5673), .B(n5672), .ZN(n5674) );
  XNOR2_X1 U7320 ( .A(n5675), .B(n5674), .ZN(n7650) );
  NAND2_X1 U7321 ( .A1(n7650), .A2(n5726), .ZN(n5677) );
  OR2_X1 U7322 ( .A1(n5728), .A2(n7633), .ZN(n5676) );
  NAND2_X1 U7323 ( .A1(n5709), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7324 ( .A1(n5707), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5683) );
  OR2_X1 U7325 ( .A1(n5678), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5679) );
  AND2_X1 U7326 ( .A1(n5680), .A2(n5679), .ZN(n9641) );
  NAND2_X1 U7327 ( .A1(n5354), .A2(n9641), .ZN(n5682) );
  NAND2_X1 U7328 ( .A1(n5708), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5681) );
  NAND4_X1 U7329 ( .A1(n5684), .A2(n5683), .A3(n5682), .A4(n5681), .ZN(n9291)
         );
  INV_X1 U7330 ( .A(n9291), .ZN(n9663) );
  NAND2_X1 U7331 ( .A1(n9643), .A2(n9663), .ZN(n5836) );
  NAND2_X1 U7332 ( .A1(n5989), .A2(n5836), .ZN(n5845) );
  OR2_X1 U7333 ( .A1(n9626), .A2(n9246), .ZN(n5848) );
  NAND2_X1 U7334 ( .A1(n5845), .A2(n5848), .ZN(n5685) );
  AND3_X1 U7335 ( .A1(n5856), .A2(n5842), .A3(n5685), .ZN(n5687) );
  INV_X1 U7336 ( .A(n5995), .ZN(n5686) );
  OAI21_X1 U7337 ( .B1(n5701), .B2(n5687), .A(n5686), .ZN(n5698) );
  NAND2_X1 U7338 ( .A1(n9118), .A2(n5726), .ZN(n5691) );
  OR2_X1 U7339 ( .A1(n5728), .A2(n10246), .ZN(n5690) );
  NAND2_X1 U7340 ( .A1(n5707), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7341 ( .A1(n5708), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5696) );
  AOI21_X1 U7342 ( .B1(n9266), .B2(n5693), .A(n5692), .ZN(n9541) );
  NAND2_X1 U7343 ( .A1(n5354), .A2(n9541), .ZN(n5695) );
  NAND2_X1 U7344 ( .A1(n5709), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5694) );
  NAND4_X1 U7345 ( .A1(n5697), .A2(n5696), .A3(n5695), .A4(n5694), .ZN(n9288)
         );
  OR2_X1 U7346 ( .A1(n9763), .A2(n9524), .ZN(n5863) );
  AND2_X1 U7347 ( .A1(n5698), .A2(n5863), .ZN(n5699) );
  OR2_X1 U7348 ( .A1(n5859), .A2(n5699), .ZN(n5700) );
  AND2_X1 U7349 ( .A1(n9763), .A2(n9524), .ZN(n9520) );
  NOR2_X1 U7350 ( .A1(n5700), .A2(n9520), .ZN(n5926) );
  INV_X1 U7351 ( .A(n5926), .ZN(n5715) );
  INV_X1 U7352 ( .A(n5701), .ZN(n5702) );
  NOR2_X1 U7353 ( .A1(n9643), .A2(n9663), .ZN(n5987) );
  INV_X1 U7354 ( .A(n5987), .ZN(n9617) );
  AND2_X1 U7355 ( .A1(n5848), .A2(n9617), .ZN(n5841) );
  NAND3_X1 U7356 ( .A1(n5702), .A2(n5863), .A3(n5841), .ZN(n5714) );
  OR2_X1 U7357 ( .A1(n9752), .A2(n9525), .ZN(n5868) );
  OAI21_X1 U7358 ( .B1(n5859), .B2(n5764), .A(n5868), .ZN(n5870) );
  INV_X1 U7359 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10247) );
  OR2_X1 U7360 ( .A1(n5728), .A2(n10247), .ZN(n5705) );
  OR2_X1 U7361 ( .A1(n5372), .A2(n9485), .ZN(n5713) );
  NAND2_X1 U7362 ( .A1(n5707), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7363 ( .A1(n5708), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7364 ( .A1(n5709), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5710) );
  NAND4_X1 U7365 ( .A1(n5713), .A2(n5712), .A3(n5711), .A4(n5710), .ZN(n9499)
         );
  INV_X1 U7366 ( .A(n9499), .ZN(n9158) );
  NOR2_X1 U7367 ( .A1(n9487), .A2(n9158), .ZN(n5741) );
  OAI21_X1 U7368 ( .B1(n5716), .B2(n5715), .A(n5932), .ZN(n5717) );
  NOR2_X1 U7369 ( .A1(n9828), .A2(n9286), .ZN(n5755) );
  NOR2_X1 U7370 ( .A1(n5755), .A2(n5873), .ZN(n5929) );
  OAI211_X1 U7371 ( .C1(n9828), .C2(n9285), .A(n5717), .B(n5929), .ZN(n5718)
         );
  OAI21_X1 U7372 ( .B1(n5878), .B2(n5879), .A(n5718), .ZN(n5738) );
  MUX2_X1 U7373 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6847), .Z(n5723) );
  INV_X1 U7374 ( .A(SI_31_), .ZN(n5722) );
  XNOR2_X1 U7375 ( .A(n5723), .B(n5722), .ZN(n5724) );
  NAND2_X1 U7376 ( .A1(n6066), .A2(n5726), .ZN(n5730) );
  INV_X1 U7377 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5727) );
  OR2_X1 U7378 ( .A1(n5728), .A2(n5727), .ZN(n5729) );
  INV_X1 U7379 ( .A(n9285), .ZN(n5731) );
  NOR2_X1 U7380 ( .A1(n9745), .A2(n9285), .ZN(n5739) );
  INV_X1 U7381 ( .A(n5733), .ZN(n5734) );
  NAND2_X1 U7382 ( .A1(n5737), .A2(n5736), .ZN(n5735) );
  INV_X1 U7383 ( .A(n9286), .ZN(n5740) );
  INV_X1 U7384 ( .A(n5739), .ZN(n5943) );
  OAI21_X1 U7385 ( .B1(n5740), .B2(n5879), .A(n5943), .ZN(n5934) );
  INV_X1 U7386 ( .A(n5933), .ZN(n5945) );
  INV_X1 U7387 ( .A(n9527), .ZN(n5753) );
  XNOR2_X1 U7388 ( .A(n9763), .B(n9524), .ZN(n9534) );
  INV_X1 U7389 ( .A(n5996), .ZN(n5862) );
  NAND2_X1 U7390 ( .A1(n5992), .A2(n5856), .ZN(n9566) );
  INV_X1 U7391 ( .A(n9566), .ZN(n5751) );
  NAND2_X1 U7392 ( .A1(n5848), .A2(n5989), .ZN(n9622) );
  XNOR2_X1 U7393 ( .A(n9643), .B(n9291), .ZN(n9635) );
  INV_X1 U7394 ( .A(n9635), .ZN(n9636) );
  INV_X1 U7395 ( .A(n9723), .ZN(n5747) );
  NAND2_X1 U7396 ( .A1(n5798), .A2(n5799), .ZN(n7642) );
  XNOR2_X1 U7397 ( .A(n9304), .B(n7421), .ZN(n7228) );
  AND2_X1 U7398 ( .A1(n7038), .A2(n9888), .ZN(n5889) );
  NOR2_X1 U7399 ( .A1(n7023), .A2(n5889), .ZN(n7454) );
  NAND2_X1 U7400 ( .A1(n5770), .A2(n5891), .ZN(n7409) );
  NOR2_X1 U7401 ( .A1(n7409), .A2(n7154), .ZN(n5742) );
  NAND4_X1 U7402 ( .A1(n7454), .A2(n5742), .A3(n5100), .A4(n7811), .ZN(n5743)
         );
  NAND2_X1 U7403 ( .A1(n5900), .A2(n7539), .ZN(n7465) );
  NOR4_X1 U7404 ( .A1(n7022), .A2(n7228), .A3(n5743), .A4(n7465), .ZN(n5744)
         );
  NAND4_X1 U7405 ( .A1(n5465), .A2(n5787), .A3(n5788), .A4(n5744), .ZN(n5745)
         );
  OR4_X1 U7406 ( .A1(n7904), .A2(n7951), .A3(n7642), .A4(n5745), .ZN(n5746) );
  NOR4_X1 U7407 ( .A1(n5747), .A2(n8014), .A3(n8147), .A4(n5746), .ZN(n5748)
         );
  NAND4_X1 U7408 ( .A1(n9676), .A2(n5566), .A3(n9700), .A4(n5748), .ZN(n5749)
         );
  NOR4_X1 U7409 ( .A1(n9622), .A2(n9636), .A3(n9657), .A4(n5749), .ZN(n5750)
         );
  XNOR2_X1 U7410 ( .A(n9782), .B(n9290), .ZN(n9607) );
  NAND4_X1 U7411 ( .A1(n5751), .A2(n9582), .A3(n5750), .A4(n9607), .ZN(n5752)
         );
  NOR4_X1 U7412 ( .A1(n5753), .A2(n9534), .A3(n9548), .A4(n5752), .ZN(n5754)
         );
  NAND3_X1 U7413 ( .A1(n6050), .A2(n9505), .A3(n5754), .ZN(n5756) );
  NOR2_X1 U7414 ( .A1(n5757), .A2(n5759), .ZN(n5758) );
  NAND2_X1 U7415 ( .A1(n5758), .A2(n7033), .ZN(n5761) );
  NAND2_X1 U7416 ( .A1(n5759), .A2(n6001), .ZN(n5760) );
  NAND2_X1 U7417 ( .A1(n5761), .A2(n5760), .ZN(n5941) );
  INV_X1 U7418 ( .A(n5863), .ZN(n5762) );
  NAND2_X1 U7419 ( .A1(n5762), .A2(n5855), .ZN(n5763) );
  AOI21_X1 U7420 ( .B1(n5764), .B2(n5763), .A(n5859), .ZN(n5766) );
  AND2_X1 U7421 ( .A1(n5832), .A2(n5767), .ZN(n5924) );
  NAND4_X1 U7422 ( .A1(n5769), .A2(n5855), .A3(n7539), .A4(n5897), .ZN(n5786)
         );
  NAND2_X1 U7423 ( .A1(n5771), .A2(n5770), .ZN(n5888) );
  NOR3_X1 U7424 ( .A1(n5888), .A2(n5772), .A3(n5855), .ZN(n5784) );
  NAND2_X1 U7425 ( .A1(n9302), .A2(n6056), .ZN(n5774) );
  INV_X1 U7426 ( .A(n9301), .ZN(n7625) );
  OAI22_X1 U7427 ( .A1(n5774), .A2(n7578), .B1(n5855), .B2(n7625), .ZN(n5773)
         );
  NAND2_X1 U7428 ( .A1(n5773), .A2(n7674), .ZN(n5782) );
  OAI21_X1 U7429 ( .B1(n5774), .B2(n7625), .A(n7584), .ZN(n5776) );
  NAND2_X1 U7430 ( .A1(n7572), .A2(n5855), .ZN(n5778) );
  OAI21_X1 U7431 ( .B1(n5778), .B2(n9301), .A(n7578), .ZN(n5775) );
  NAND2_X1 U7432 ( .A1(n5776), .A2(n5775), .ZN(n5781) );
  NAND2_X1 U7433 ( .A1(n5777), .A2(n7634), .ZN(n7534) );
  INV_X1 U7434 ( .A(n7534), .ZN(n7538) );
  OAI22_X1 U7435 ( .A1(n5778), .A2(n7584), .B1(n6056), .B2(n9301), .ZN(n5779)
         );
  INV_X1 U7436 ( .A(n7674), .ZN(n7469) );
  NAND2_X1 U7437 ( .A1(n5779), .A2(n7469), .ZN(n5780) );
  NAND4_X1 U7438 ( .A1(n5782), .A2(n5781), .A3(n7538), .A4(n5780), .ZN(n5783)
         );
  AOI21_X1 U7439 ( .B1(n5896), .B2(n5784), .A(n5783), .ZN(n5785) );
  NAND2_X1 U7440 ( .A1(n5786), .A2(n5785), .ZN(n5790) );
  MUX2_X1 U7441 ( .A(n5788), .B(n5787), .S(n6056), .Z(n5789) );
  NAND2_X1 U7442 ( .A1(n5790), .A2(n5789), .ZN(n5793) );
  AND2_X1 U7443 ( .A1(n5799), .A2(n7636), .ZN(n5791) );
  MUX2_X1 U7444 ( .A(n7637), .B(n5791), .S(n5855), .Z(n5792) );
  NAND2_X1 U7445 ( .A1(n5793), .A2(n5792), .ZN(n5801) );
  AOI21_X1 U7446 ( .B1(n5801), .B2(n5798), .A(n5794), .ZN(n5796) );
  NAND2_X1 U7447 ( .A1(n5804), .A2(n5904), .ZN(n5795) );
  OAI211_X1 U7448 ( .C1(n5796), .C2(n5795), .A(n5910), .B(n5802), .ZN(n5797)
         );
  OR2_X1 U7449 ( .A1(n8221), .A2(n6023), .ZN(n5805) );
  NAND2_X1 U7450 ( .A1(n5797), .A2(n5805), .ZN(n5808) );
  INV_X1 U7451 ( .A(n5798), .ZN(n5800) );
  OAI21_X1 U7452 ( .B1(n5801), .B2(n5800), .A(n5799), .ZN(n5803) );
  NAND2_X1 U7453 ( .A1(n5802), .A2(n7946), .ZN(n5906) );
  AOI21_X1 U7454 ( .B1(n5803), .B2(n5904), .A(n5906), .ZN(n5806) );
  NAND2_X1 U7455 ( .A1(n5805), .A2(n5804), .ZN(n5911) );
  OAI21_X1 U7456 ( .B1(n5806), .B2(n5911), .A(n5910), .ZN(n5807) );
  MUX2_X1 U7457 ( .A(n5808), .B(n5807), .S(n6056), .Z(n5812) );
  AND2_X1 U7458 ( .A1(n8212), .A2(n9179), .ZN(n5811) );
  OR2_X1 U7459 ( .A1(n8147), .A2(n5811), .ZN(n5809) );
  AOI21_X1 U7460 ( .B1(n5812), .B2(n5913), .A(n5809), .ZN(n5810) );
  NAND2_X1 U7461 ( .A1(n5916), .A2(n6056), .ZN(n5818) );
  INV_X1 U7462 ( .A(n5811), .ZN(n5909) );
  NAND2_X1 U7463 ( .A1(n5812), .A2(n5909), .ZN(n5813) );
  NAND3_X1 U7464 ( .A1(n5813), .A2(n4874), .A3(n5913), .ZN(n5814) );
  NAND3_X1 U7465 ( .A1(n5814), .A2(n5855), .A3(n5918), .ZN(n5815) );
  NAND2_X1 U7466 ( .A1(n5816), .A2(n5815), .ZN(n5820) );
  NAND2_X1 U7467 ( .A1(n5821), .A2(n5817), .ZN(n5915) );
  NAND2_X1 U7468 ( .A1(n5915), .A2(n5818), .ZN(n5819) );
  NAND2_X1 U7469 ( .A1(n5820), .A2(n5819), .ZN(n5828) );
  INV_X1 U7470 ( .A(n5821), .ZN(n5822) );
  NAND2_X1 U7471 ( .A1(n5829), .A2(n5822), .ZN(n5823) );
  OAI211_X1 U7472 ( .C1(n9734), .C2(n6056), .A(n5823), .B(n5918), .ZN(n5826)
         );
  NAND2_X1 U7473 ( .A1(n5918), .A2(n9701), .ZN(n5824) );
  NAND2_X1 U7474 ( .A1(n5824), .A2(n5855), .ZN(n5825) );
  NAND2_X1 U7475 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  OAI211_X1 U7476 ( .C1(n5829), .C2(n6056), .A(n5828), .B(n5827), .ZN(n5830)
         );
  NAND2_X1 U7477 ( .A1(n5830), .A2(n5566), .ZN(n5835) );
  NAND2_X1 U7478 ( .A1(n5924), .A2(n5835), .ZN(n5831) );
  NAND2_X1 U7479 ( .A1(n5837), .A2(n5832), .ZN(n5927) );
  AND2_X1 U7480 ( .A1(n5834), .A2(n5833), .ZN(n5921) );
  INV_X1 U7481 ( .A(n5837), .ZN(n5838) );
  OAI21_X1 U7482 ( .B1(n5987), .B2(n5838), .A(n5855), .ZN(n5839) );
  NAND2_X1 U7483 ( .A1(n5840), .A2(n5839), .ZN(n5847) );
  AOI21_X1 U7484 ( .B1(n5847), .B2(n5841), .A(n4848), .ZN(n5843) );
  OAI21_X1 U7485 ( .B1(n4744), .B2(n5843), .A(n5842), .ZN(n5850) );
  INV_X1 U7486 ( .A(n5845), .ZN(n5846) );
  NAND2_X1 U7487 ( .A1(n5847), .A2(n5846), .ZN(n5849) );
  INV_X1 U7488 ( .A(n9565), .ZN(n5991) );
  NOR2_X1 U7489 ( .A1(n5851), .A2(n5855), .ZN(n5852) );
  NOR2_X1 U7490 ( .A1(n9566), .A2(n5852), .ZN(n5853) );
  NAND2_X1 U7491 ( .A1(n5854), .A2(n5853), .ZN(n5858) );
  MUX2_X1 U7492 ( .A(n5856), .B(n5992), .S(n5855), .Z(n5857) );
  NAND2_X1 U7493 ( .A1(n5858), .A2(n5857), .ZN(n5865) );
  INV_X1 U7494 ( .A(n5859), .ZN(n5861) );
  NOR3_X1 U7495 ( .A1(n9520), .A2(n5995), .A3(n6056), .ZN(n5860) );
  OAI211_X1 U7496 ( .C1(n5862), .C2(n5865), .A(n5861), .B(n5860), .ZN(n5869)
         );
  AND3_X1 U7497 ( .A1(n5863), .A2(n6056), .A3(n5996), .ZN(n5864) );
  OAI21_X1 U7498 ( .B1(n5865), .B2(n5995), .A(n5864), .ZN(n5867) );
  NAND3_X1 U7499 ( .A1(n9763), .A2(n9524), .A3(n6056), .ZN(n5866) );
  INV_X1 U7500 ( .A(n5873), .ZN(n5875) );
  INV_X1 U7501 ( .A(n5741), .ZN(n5874) );
  MUX2_X1 U7502 ( .A(n5875), .B(n5874), .S(n6056), .Z(n5876) );
  NAND2_X1 U7503 ( .A1(n5933), .A2(n5878), .ZN(n5882) );
  OAI21_X1 U7504 ( .B1(n5942), .B2(n7033), .A(n6056), .ZN(n5884) );
  NAND2_X1 U7505 ( .A1(n5884), .A2(n5883), .ZN(n5887) );
  NAND2_X1 U7506 ( .A1(n5885), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7507 ( .A1(n5887), .A2(n7140), .ZN(n5940) );
  INV_X1 U7508 ( .A(n5888), .ZN(n5895) );
  AOI21_X1 U7509 ( .B1(n4512), .B2(n9944), .A(n7811), .ZN(n5892) );
  INV_X1 U7510 ( .A(n5889), .ZN(n5890) );
  NAND4_X1 U7511 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n5894)
         );
  NAND3_X1 U7512 ( .A1(n5896), .A2(n5895), .A3(n5894), .ZN(n5898) );
  NAND2_X1 U7513 ( .A1(n5898), .A2(n5897), .ZN(n5902) );
  INV_X1 U7514 ( .A(n5899), .ZN(n5901) );
  NAND3_X1 U7515 ( .A1(n5902), .A2(n5901), .A3(n5900), .ZN(n5905) );
  NAND3_X1 U7516 ( .A1(n5905), .A2(n5904), .A3(n5903), .ZN(n5908) );
  INV_X1 U7517 ( .A(n5906), .ZN(n5907) );
  AND2_X1 U7518 ( .A1(n5908), .A2(n5907), .ZN(n5912) );
  OAI211_X1 U7519 ( .C1(n5912), .C2(n5911), .A(n5910), .B(n5909), .ZN(n5914)
         );
  AND2_X1 U7520 ( .A1(n5914), .A2(n5913), .ZN(n5917) );
  AOI21_X1 U7521 ( .B1(n5917), .B2(n5916), .A(n5915), .ZN(n5919) );
  OAI21_X1 U7522 ( .B1(n5920), .B2(n5919), .A(n5918), .ZN(n5923) );
  INV_X1 U7523 ( .A(n5921), .ZN(n5922) );
  AOI21_X1 U7524 ( .B1(n5924), .B2(n5923), .A(n5922), .ZN(n5928) );
  OAI211_X1 U7525 ( .C1(n5928), .C2(n5927), .A(n5926), .B(n5925), .ZN(n5931)
         );
  INV_X1 U7526 ( .A(n5929), .ZN(n5930) );
  AOI21_X1 U7527 ( .B1(n5932), .B2(n5931), .A(n5930), .ZN(n5935) );
  OAI21_X1 U7528 ( .B1(n5935), .B2(n5934), .A(n5933), .ZN(n5936) );
  XNOR2_X1 U7529 ( .A(n5936), .B(n7033), .ZN(n5938) );
  OAI21_X1 U7530 ( .B1(n5943), .B2(n6056), .A(n5942), .ZN(n5944) );
  NAND2_X1 U7531 ( .A1(n5883), .A2(n7140), .ZN(n6002) );
  AOI211_X1 U7532 ( .C1(n5945), .C2(n6001), .A(n6053), .B(n6002), .ZN(n5946)
         );
  NAND2_X1 U7533 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  NAND2_X1 U7534 ( .A1(n5951), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5953) );
  OR2_X1 U7535 ( .A1(n7239), .A2(P1_U3086), .ZN(n7925) );
  INV_X1 U7536 ( .A(n7925), .ZN(n5954) );
  OAI21_X1 U7537 ( .B1(n5956), .B2(n5955), .A(n5954), .ZN(n5970) );
  INV_X1 U7538 ( .A(n5958), .ZN(n5959) );
  NAND2_X1 U7539 ( .A1(n5959), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5961) );
  XNOR2_X1 U7540 ( .A(n5961), .B(n5960), .ZN(n8050) );
  OR2_X1 U7541 ( .A1(n5962), .A2(n5171), .ZN(n5963) );
  NAND2_X1 U7542 ( .A1(n5964), .A2(n5963), .ZN(n9885) );
  OR2_X1 U7543 ( .A1(n6004), .A2(n6054), .ZN(n6052) );
  INV_X1 U7544 ( .A(n6052), .ZN(n5965) );
  AND2_X1 U7545 ( .A1(n9866), .A2(n5965), .ZN(n7139) );
  NOR2_X1 U7546 ( .A1(n5966), .A2(n9927), .ZN(n6909) );
  NAND2_X1 U7547 ( .A1(n7139), .A2(n6909), .ZN(n5968) );
  OAI211_X1 U7548 ( .C1(n6053), .C2(n7925), .A(n5968), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5969) );
  NAND2_X1 U7549 ( .A1(n5970), .A2(n5969), .ZN(P1_U3242) );
  OR2_X1 U7550 ( .A1(n6004), .A2(n7146), .ZN(n7238) );
  INV_X1 U7551 ( .A(n7028), .ZN(n7145) );
  NAND2_X1 U7552 ( .A1(n9885), .A2(P1_B_REG_SCAN_IN), .ZN(n5971) );
  MUX2_X1 U7553 ( .A(P1_B_REG_SCAN_IN), .B(n5971), .S(n8050), .Z(n5972) );
  NAND2_X1 U7554 ( .A1(n5973), .A2(n5972), .ZN(n6864) );
  INV_X1 U7555 ( .A(n6864), .ZN(n5986) );
  INV_X1 U7556 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10387) );
  NAND2_X1 U7557 ( .A1(n5986), .A2(n10387), .ZN(n5975) );
  NAND2_X1 U7558 ( .A1(n9881), .A2(n8050), .ZN(n5974) );
  NAND2_X1 U7559 ( .A1(n5975), .A2(n5974), .ZN(n7125) );
  AND2_X1 U7560 ( .A1(n7145), .A2(n7125), .ZN(n7390) );
  NAND2_X1 U7561 ( .A1(n9881), .A2(n9885), .ZN(n6865) );
  OAI21_X1 U7562 ( .B1(n6864), .B2(P1_D_REG_1__SCAN_IN), .A(n6865), .ZN(n7123)
         );
  NOR4_X1 U7563 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5984) );
  NOR4_X1 U7564 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5983) );
  INV_X1 U7565 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10211) );
  INV_X1 U7566 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10498) );
  INV_X1 U7567 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10524) );
  INV_X1 U7568 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10368) );
  NAND4_X1 U7569 ( .A1(n10211), .A2(n10498), .A3(n10524), .A4(n10368), .ZN(
        n5981) );
  NOR4_X1 U7570 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5979) );
  NOR4_X1 U7571 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5978) );
  NOR4_X1 U7572 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5977) );
  NOR4_X1 U7573 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5976) );
  NAND4_X1 U7574 ( .A1(n5979), .A2(n5978), .A3(n5977), .A4(n5976), .ZN(n5980)
         );
  NOR4_X1 U7575 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5981), .A4(n5980), .ZN(n5982) );
  NAND3_X1 U7576 ( .A1(n5984), .A2(n5983), .A3(n5982), .ZN(n5985) );
  NAND2_X1 U7577 ( .A1(n5986), .A2(n5985), .ZN(n7122) );
  NOR2_X1 U7578 ( .A1(n9622), .A2(n5987), .ZN(n5988) );
  NAND2_X1 U7579 ( .A1(n9606), .A2(n5990), .ZN(n9581) );
  NAND2_X1 U7580 ( .A1(n9581), .A2(n9582), .ZN(n9580) );
  NOR2_X1 U7581 ( .A1(n9566), .A2(n5991), .ZN(n5994) );
  INV_X1 U7582 ( .A(n5992), .ZN(n5993) );
  NAND2_X1 U7583 ( .A1(n9519), .A2(n5997), .ZN(n9496) );
  NAND2_X1 U7584 ( .A1(n9496), .A2(n9505), .ZN(n9497) );
  NAND2_X1 U7585 ( .A1(n9497), .A2(n5998), .ZN(n6000) );
  NAND2_X1 U7586 ( .A1(n6053), .A2(n6001), .ZN(n6003) );
  INV_X1 U7587 ( .A(n9525), .ZN(n9287) );
  INV_X1 U7588 ( .A(n5966), .ZN(n7049) );
  INV_X1 U7589 ( .A(n9927), .ZN(n7047) );
  AND2_X1 U7590 ( .A1(n7047), .A2(P1_B_REG_SCAN_IN), .ZN(n6005) );
  NOR2_X1 U7591 ( .A1(n9664), .A2(n6005), .ZN(n6061) );
  AOI22_X1 U7592 ( .A1(n9287), .A2(n9727), .B1(n9286), .B2(n6061), .ZN(n6006)
         );
  NOR2_X1 U7593 ( .A1(n7153), .A2(n7256), .ZN(n7232) );
  NAND2_X1 U7594 ( .A1(n7232), .A2(n7421), .ZN(n7411) );
  INV_X1 U7595 ( .A(n9921), .ZN(n7764) );
  INV_X1 U7596 ( .A(n8109), .ZN(n9904) );
  INV_X1 U7597 ( .A(n7987), .ZN(n9965) );
  NOR2_X1 U7598 ( .A1(n9798), .A2(n9669), .ZN(n9651) );
  NAND2_X1 U7599 ( .A1(n9852), .A2(n9651), .ZN(n9640) );
  NOR2_X1 U7600 ( .A1(n9590), .A2(n9600), .ZN(n9589) );
  NAND2_X1 U7601 ( .A1(n9544), .A2(n9555), .ZN(n9538) );
  INV_X1 U7602 ( .A(n6007), .ZN(n9509) );
  OAI21_X1 U7603 ( .B1(n6009), .B2(n9509), .A(n6008), .ZN(n9491) );
  INV_X1 U7604 ( .A(n7175), .ZN(n6010) );
  INV_X1 U7605 ( .A(n9956), .ZN(n6011) );
  NAND2_X1 U7606 ( .A1(n7038), .A2(n7041), .ZN(n7021) );
  NAND2_X1 U7607 ( .A1(n6013), .A2(n7021), .ZN(n7020) );
  OR2_X1 U7608 ( .A1(n9305), .A2(n7256), .ZN(n6015) );
  NAND2_X1 U7609 ( .A1(n7151), .A2(n6015), .ZN(n7225) );
  NAND2_X1 U7610 ( .A1(n7225), .A2(n7228), .ZN(n7224) );
  NAND2_X1 U7611 ( .A1(n6016), .A2(n7421), .ZN(n6017) );
  NAND2_X1 U7612 ( .A1(n7224), .A2(n6017), .ZN(n7410) );
  OR2_X1 U7613 ( .A1(n9303), .A2(n7414), .ZN(n6018) );
  NAND2_X1 U7614 ( .A1(n7572), .A2(n7584), .ZN(n6019) );
  NAND2_X1 U7615 ( .A1(n7535), .A2(n7534), .ZN(n7537) );
  NAND2_X1 U7616 ( .A1(n7637), .A2(n7636), .ZN(n7656) );
  INV_X1 U7617 ( .A(n7985), .ZN(n9298) );
  NAND2_X1 U7618 ( .A1(n9904), .A2(n8123), .ZN(n6021) );
  NAND2_X1 U7619 ( .A1(n8115), .A2(n9296), .ZN(n6022) );
  AOI21_X2 U7620 ( .B1(n7940), .B2(n6022), .A(n5145), .ZN(n7903) );
  NAND2_X1 U7621 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  NAND2_X1 U7622 ( .A1(n8221), .A2(n9295), .ZN(n6026) );
  NAND2_X1 U7623 ( .A1(n9705), .A2(n9704), .ZN(n9706) );
  INV_X1 U7624 ( .A(n9812), .ZN(n9710) );
  NAND2_X1 U7625 ( .A1(n9858), .A2(n9256), .ZN(n6029) );
  NAND2_X1 U7626 ( .A1(n9688), .A2(n6029), .ZN(n6031) );
  NAND2_X1 U7627 ( .A1(n9652), .A2(n9292), .ZN(n6033) );
  NAND2_X1 U7628 ( .A1(n9643), .A2(n9291), .ZN(n6034) );
  NAND2_X2 U7629 ( .A1(n6035), .A2(n6034), .ZN(n9616) );
  NOR2_X1 U7630 ( .A1(n9848), .A2(n9246), .ZN(n6036) );
  INV_X1 U7631 ( .A(n9246), .ZN(n9610) );
  NOR2_X1 U7632 ( .A1(n9782), .A2(n9290), .ZN(n6037) );
  INV_X1 U7633 ( .A(n9782), .ZN(n9605) );
  NOR2_X1 U7634 ( .A1(n9843), .A2(n9569), .ZN(n6038) );
  NAND2_X1 U7635 ( .A1(n9843), .A2(n9569), .ZN(n6039) );
  NAND2_X1 U7636 ( .A1(n9576), .A2(n9585), .ZN(n6040) );
  NAND2_X1 U7637 ( .A1(n9564), .A2(n6040), .ZN(n6042) );
  NAND2_X1 U7638 ( .A1(n9773), .A2(n9289), .ZN(n6041) );
  NAND2_X1 U7639 ( .A1(n6042), .A2(n6041), .ZN(n9547) );
  INV_X1 U7640 ( .A(n9547), .ZN(n6043) );
  NAND2_X1 U7641 ( .A1(n6043), .A2(n5159), .ZN(n6045) );
  NAND2_X1 U7642 ( .A1(n9838), .A2(n9570), .ZN(n6044) );
  NOR2_X1 U7643 ( .A1(n9763), .A2(n9288), .ZN(n6046) );
  NAND2_X1 U7644 ( .A1(n9833), .A2(n9537), .ZN(n9503) );
  INV_X1 U7645 ( .A(n9505), .ZN(n6047) );
  AND2_X1 U7646 ( .A1(n9503), .A2(n6047), .ZN(n6048) );
  NAND2_X1 U7647 ( .A1(n9752), .A2(n9287), .ZN(n6049) );
  XNOR2_X1 U7648 ( .A(n6051), .B(n6050), .ZN(n9484) );
  NAND2_X1 U7649 ( .A1(n6052), .A2(n7175), .ZN(n7453) );
  NAND2_X1 U7650 ( .A1(n6053), .A2(n7033), .ZN(n7040) );
  AND2_X1 U7651 ( .A1(n7040), .A2(n6054), .ZN(n6055) );
  OR2_X1 U7652 ( .A1(n7453), .A2(n6055), .ZN(n7658) );
  INV_X1 U7653 ( .A(n9860), .ZN(n6057) );
  NAND2_X1 U7654 ( .A1(n6057), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7655 ( .A1(n6059), .A2(n6058), .ZN(P1_U3519) );
  INV_X1 U7656 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7657 ( .A1(n9285), .A2(n6061), .ZN(n9746) );
  MUX2_X1 U7658 ( .A(n6062), .B(n9743), .S(n9860), .Z(n6065) );
  INV_X1 U7659 ( .A(n9864), .ZN(n6063) );
  NAND2_X1 U7660 ( .A1(n5732), .A2(n6063), .ZN(n6064) );
  NAND2_X1 U7661 ( .A1(n6065), .A2(n6064), .ZN(P1_U3521) );
  AND2_X2 U7662 ( .A1(n6811), .A2(n6304), .ZN(n6295) );
  AND2_X2 U7663 ( .A1(n6295), .A2(n6296), .ZN(n6240) );
  NOR2_X1 U7664 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n6070) );
  NAND4_X1 U7665 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(n6074)
         );
  NAND4_X1 U7666 ( .A1(n6416), .A2(n6072), .A3(n6242), .A4(n6071), .ZN(n6073)
         );
  INV_X1 U7667 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7668 ( .A1(n6066), .A2(n6431), .ZN(n6086) );
  INV_X1 U7669 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9106) );
  OR2_X1 U7670 ( .A1(n4515), .A2(n9106), .ZN(n6085) );
  NOR2_X1 U7671 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6281) );
  NAND2_X1 U7672 ( .A1(n6281), .A2(n6087), .ZN(n6374) );
  NAND2_X1 U7673 ( .A1(n6436), .A2(n10480), .ZN(n6451) );
  INV_X1 U7674 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6089) );
  INV_X1 U7675 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10380) );
  INV_X1 U7676 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7677 ( .A1(n6155), .A2(n6090), .ZN(n6157) );
  INV_X1 U7678 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6091) );
  INV_X1 U7679 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7680 ( .A1(n6097), .A2(n6093), .ZN(n9104) );
  XNOR2_X2 U7681 ( .A(n6095), .B(n6094), .ZN(n8345) );
  INV_X1 U7682 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6096) );
  XNOR2_X2 U7683 ( .A(n6098), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7684 ( .A1(n8323), .A2(n6202), .ZN(n6118) );
  INV_X1 U7685 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6103) );
  NAND2_X2 U7686 ( .A1(n6099), .A2(n8330), .ZN(n6339) );
  NAND2_X1 U7687 ( .A1(n6300), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7688 ( .A1(n6372), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6101) );
  OAI211_X1 U7689 ( .C1(n6103), .C2(n4513), .A(n6102), .B(n6101), .ZN(n6104)
         );
  INV_X1 U7690 ( .A(n6104), .ZN(n6105) );
  INV_X1 U7691 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8346) );
  NOR2_X1 U7692 ( .A1(n4515), .A2(n8346), .ZN(n6106) );
  INV_X1 U7693 ( .A(n8949), .ZN(n9011) );
  INV_X1 U7694 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7695 ( .A1(n6300), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7696 ( .A1(n6372), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6107) );
  OAI211_X1 U7697 ( .C1(n6109), .C2(n4513), .A(n6108), .B(n6107), .ZN(n6110)
         );
  INV_X1 U7698 ( .A(n6110), .ZN(n6111) );
  NAND2_X1 U7699 ( .A1(n6118), .A2(n6111), .ZN(n8554) );
  INV_X1 U7700 ( .A(n8554), .ZN(n6112) );
  AND2_X1 U7701 ( .A1(n9011), .A2(n6112), .ZN(n6651) );
  INV_X1 U7702 ( .A(n6651), .ZN(n6119) );
  INV_X1 U7703 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8329) );
  OR2_X1 U7704 ( .A1(n4515), .A2(n8329), .ZN(n6113) );
  INV_X1 U7705 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U7706 ( .A1(n6300), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7707 ( .A1(n6372), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6114) );
  OAI211_X1 U7708 ( .C1(n6786), .C2(n4513), .A(n6115), .B(n6114), .ZN(n6116)
         );
  INV_X1 U7709 ( .A(n6116), .ZN(n6117) );
  NAND2_X1 U7710 ( .A1(n6772), .A2(n8555), .ZN(n6486) );
  NAND2_X1 U7711 ( .A1(n6119), .A2(n6486), .ZN(n6642) );
  INV_X1 U7712 ( .A(n6642), .ZN(n6120) );
  NAND2_X1 U7713 ( .A1(n4538), .A2(n6120), .ZN(n6489) );
  INV_X1 U7714 ( .A(n6489), .ZN(n6463) );
  INV_X1 U7715 ( .A(n6487), .ZN(n6647) );
  NAND2_X1 U7716 ( .A1(n9113), .A2(n6431), .ZN(n6123) );
  OR2_X1 U7717 ( .A1(n4515), .A2(n6121), .ZN(n6122) );
  INV_X1 U7718 ( .A(n6124), .ZN(n6136) );
  NAND2_X1 U7719 ( .A1(n6147), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7720 ( .A1(n6136), .A2(n6125), .ZN(n8739) );
  NAND2_X1 U7721 ( .A1(n8739), .A2(n6202), .ZN(n6131) );
  INV_X1 U7722 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7723 ( .A1(n6300), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7724 ( .A1(n6372), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6126) );
  OAI211_X1 U7725 ( .C1(n6128), .C2(n4513), .A(n6127), .B(n6126), .ZN(n6129)
         );
  INV_X1 U7726 ( .A(n6129), .ZN(n6130) );
  XNOR2_X1 U7727 ( .A(n8743), .B(n8750), .ZN(n8734) );
  INV_X1 U7728 ( .A(n8734), .ZN(n8731) );
  NAND2_X1 U7729 ( .A1(n6132), .A2(n6431), .ZN(n6135) );
  OR2_X1 U7730 ( .A1(n4515), .A2(n6133), .ZN(n6134) );
  INV_X1 U7731 ( .A(n8323), .ZN(n6138) );
  NAND2_X1 U7732 ( .A1(n6136), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7733 ( .A1(n6138), .A2(n6137), .ZN(n8728) );
  NAND2_X1 U7734 ( .A1(n8728), .A2(n6202), .ZN(n6143) );
  INV_X1 U7735 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U7736 ( .A1(n6300), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7737 ( .A1(n6372), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6139) );
  OAI211_X1 U7738 ( .C1(n9015), .C2(n4513), .A(n6140), .B(n6139), .ZN(n6141)
         );
  INV_X1 U7739 ( .A(n6141), .ZN(n6142) );
  INV_X1 U7740 ( .A(n8718), .ZN(n8720) );
  NAND2_X1 U7741 ( .A1(n9118), .A2(n6431), .ZN(n6145) );
  OR2_X1 U7742 ( .A1(n4515), .A2(n9119), .ZN(n6144) );
  NAND2_X1 U7743 ( .A1(n6157), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7744 ( .A1(n6147), .A2(n6146), .ZN(n8753) );
  NAND2_X1 U7745 ( .A1(n8753), .A2(n6202), .ZN(n6152) );
  INV_X1 U7746 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U7747 ( .A1(n6300), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7748 ( .A1(n6372), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6148) );
  OAI211_X1 U7749 ( .C1(n9022), .C2(n4513), .A(n6149), .B(n6148), .ZN(n6150)
         );
  INV_X1 U7750 ( .A(n6150), .ZN(n6151) );
  NAND2_X1 U7751 ( .A1(n9023), .A2(n8389), .ZN(n6633) );
  NAND2_X1 U7752 ( .A1(n9121), .A2(n6431), .ZN(n6154) );
  OR2_X1 U7753 ( .A1(n4515), .A2(n9123), .ZN(n6153) );
  INV_X1 U7754 ( .A(n6155), .ZN(n6166) );
  NAND2_X1 U7755 ( .A1(n6166), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7756 ( .A1(n6157), .A2(n6156), .ZN(n8762) );
  NAND2_X1 U7757 ( .A1(n8762), .A2(n6202), .ZN(n6162) );
  INV_X1 U7758 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U7759 ( .A1(n6300), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7760 ( .A1(n6372), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6158) );
  OAI211_X1 U7761 ( .C1(n9028), .C2(n4513), .A(n6159), .B(n6158), .ZN(n6160)
         );
  INV_X1 U7762 ( .A(n6160), .ZN(n6161) );
  NAND2_X1 U7763 ( .A1(n9029), .A2(n8529), .ZN(n6629) );
  NAND2_X1 U7764 ( .A1(n8025), .A2(n6431), .ZN(n6164) );
  OR2_X1 U7765 ( .A1(n4515), .A2(n8026), .ZN(n6163) );
  NAND2_X1 U7766 ( .A1(n6175), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7767 ( .A1(n6166), .A2(n6165), .ZN(n8779) );
  NAND2_X1 U7768 ( .A1(n8779), .A2(n6202), .ZN(n6171) );
  INV_X1 U7769 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U7770 ( .A1(n6300), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7771 ( .A1(n6372), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6167) );
  OAI211_X1 U7772 ( .C1(n9034), .C2(n4513), .A(n6168), .B(n6167), .ZN(n6169)
         );
  INV_X1 U7773 ( .A(n6169), .ZN(n6170) );
  NAND2_X1 U7774 ( .A1(n9035), .A2(n8475), .ZN(n6622) );
  NAND2_X1 U7775 ( .A1(n7927), .A2(n6431), .ZN(n6173) );
  OR2_X1 U7776 ( .A1(n4515), .A2(n7930), .ZN(n6172) );
  INV_X1 U7777 ( .A(n9041), .ZN(n6179) );
  NAND2_X1 U7778 ( .A1(n6183), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7779 ( .A1(n6175), .A2(n6174), .ZN(n8792) );
  NAND2_X1 U7780 ( .A1(n8792), .A2(n6202), .ZN(n6178) );
  AOI22_X1 U7781 ( .A1(n6300), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n6372), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7782 ( .A1(n6393), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6176) );
  INV_X1 U7783 ( .A(n8770), .ZN(n6620) );
  NAND2_X1 U7784 ( .A1(n6620), .A2(n8771), .ZN(n8786) );
  NAND2_X1 U7785 ( .A1(n7918), .A2(n6431), .ZN(n6181) );
  OR2_X1 U7786 ( .A1(n4515), .A2(n7921), .ZN(n6180) );
  NAND2_X1 U7787 ( .A1(n6193), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7788 ( .A1(n6183), .A2(n6182), .ZN(n8802) );
  NAND2_X1 U7789 ( .A1(n8802), .A2(n6202), .ZN(n6186) );
  AOI22_X1 U7790 ( .A1(n6300), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n6372), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7791 ( .A1(n6393), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7792 ( .A1(n8507), .A2(n8809), .ZN(n6616) );
  NAND2_X1 U7793 ( .A1(n7786), .A2(n6431), .ZN(n6188) );
  INV_X1 U7794 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7787) );
  OR2_X1 U7795 ( .A1(n4515), .A2(n7787), .ZN(n6187) );
  NAND2_X1 U7796 ( .A1(n6300), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7797 ( .A1(n6372), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6189) );
  AND2_X1 U7798 ( .A1(n6190), .A2(n6189), .ZN(n6196) );
  INV_X1 U7799 ( .A(n6191), .ZN(n6201) );
  NAND2_X1 U7800 ( .A1(n6201), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7801 ( .A1(n6193), .A2(n6192), .ZN(n8818) );
  NAND2_X1 U7802 ( .A1(n8818), .A2(n6202), .ZN(n6195) );
  NAND2_X1 U7803 ( .A1(n6393), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7804 ( .A1(n8817), .A2(n8798), .ZN(n6500) );
  NAND2_X1 U7805 ( .A1(n6612), .A2(n6500), .ZN(n8814) );
  NAND2_X1 U7806 ( .A1(n7650), .A2(n6431), .ZN(n6198) );
  OR2_X1 U7807 ( .A1(n4515), .A2(n7651), .ZN(n6197) );
  INV_X1 U7808 ( .A(n6199), .ZN(n6212) );
  NAND2_X1 U7809 ( .A1(n6212), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7810 ( .A1(n6201), .A2(n6200), .ZN(n8834) );
  NAND2_X1 U7811 ( .A1(n6202), .A2(n8834), .ZN(n6206) );
  INV_X1 U7812 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8833) );
  OR2_X1 U7813 ( .A1(n6339), .A2(n8833), .ZN(n6205) );
  INV_X1 U7814 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8981) );
  OR2_X1 U7815 ( .A1(n6340), .A2(n8981), .ZN(n6204) );
  INV_X1 U7816 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9055) );
  OR2_X1 U7817 ( .A1(n4513), .A2(n9055), .ZN(n6203) );
  NAND2_X1 U7818 ( .A1(n9056), .A2(n8808), .ZN(n8813) );
  NAND2_X1 U7819 ( .A1(n7530), .A2(n6431), .ZN(n6210) );
  NAND2_X1 U7820 ( .A1(n6207), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7821 ( .A1(n6218), .A2(n6217), .ZN(n6220) );
  NAND2_X1 U7822 ( .A1(n6220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6208) );
  AOI22_X1 U7823 ( .A1(n6446), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8705), .B2(
        n6445), .ZN(n6209) );
  NAND2_X1 U7824 ( .A1(n6393), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6216) );
  INV_X1 U7825 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8843) );
  OR2_X1 U7826 ( .A1(n6339), .A2(n8843), .ZN(n6215) );
  INV_X1 U7827 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8984) );
  OR2_X1 U7828 ( .A1(n6340), .A2(n8984), .ZN(n6214) );
  NAND2_X1 U7829 ( .A1(n6224), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6211) );
  AND2_X1 U7830 ( .A1(n6212), .A2(n6211), .ZN(n8844) );
  OR2_X1 U7831 ( .A1(n4517), .A2(n8844), .ZN(n6213) );
  NAND2_X1 U7832 ( .A1(n9062), .A2(n8854), .ZN(n6601) );
  NAND2_X1 U7833 ( .A1(n7451), .A2(n6431), .ZN(n6222) );
  OR2_X1 U7834 ( .A1(n6218), .A2(n6217), .ZN(n6219) );
  AND2_X1 U7835 ( .A1(n6220), .A2(n6219), .ZN(n8697) );
  AOI22_X1 U7836 ( .A1(n6446), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6445), .B2(
        n8697), .ZN(n6221) );
  NAND2_X1 U7837 ( .A1(n6300), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6228) );
  INV_X1 U7838 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8989) );
  OR2_X1 U7839 ( .A1(n6340), .A2(n8989), .ZN(n6227) );
  NAND2_X1 U7840 ( .A1(n6235), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6223) );
  AND2_X1 U7841 ( .A1(n6224), .A2(n6223), .ZN(n8856) );
  OR2_X1 U7842 ( .A1(n4517), .A2(n8856), .ZN(n6226) );
  INV_X1 U7843 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9067) );
  OR2_X1 U7844 ( .A1(n4513), .A2(n9067), .ZN(n6225) );
  NAND2_X1 U7845 ( .A1(n8988), .A2(n8466), .ZN(n6584) );
  NAND2_X1 U7846 ( .A1(n6578), .A2(n6584), .ZN(n8852) );
  INV_X1 U7847 ( .A(n8852), .ZN(n8849) );
  NAND2_X1 U7848 ( .A1(n7236), .A2(n6431), .ZN(n6232) );
  NAND2_X1 U7849 ( .A1(n6259), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6230) );
  XNOR2_X1 U7850 ( .A(n6230), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8685) );
  AOI22_X1 U7851 ( .A1(n6446), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6445), .B2(
        n8685), .ZN(n6231) );
  NAND2_X1 U7852 ( .A1(n6393), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6239) );
  INV_X1 U7853 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8866) );
  OR2_X1 U7854 ( .A1(n6339), .A2(n8866), .ZN(n6238) );
  INV_X1 U7855 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8991) );
  OR2_X1 U7856 ( .A1(n6340), .A2(n8991), .ZN(n6237) );
  INV_X1 U7857 ( .A(n6233), .ZN(n6265) );
  NAND2_X1 U7858 ( .A1(n6265), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6234) );
  AND2_X1 U7859 ( .A1(n6235), .A2(n6234), .ZN(n8867) );
  OR2_X1 U7860 ( .A1(n4517), .A2(n8867), .ZN(n6236) );
  NAND2_X1 U7861 ( .A1(n9072), .A2(n8855), .ZN(n6583) );
  NAND2_X1 U7862 ( .A1(n6577), .A2(n6583), .ZN(n8863) );
  NAND2_X1 U7863 ( .A1(n7162), .A2(n6431), .ZN(n6250) );
  NAND2_X1 U7864 ( .A1(n6240), .A2(n6332), .ZN(n6287) );
  INV_X1 U7865 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6402) );
  INV_X1 U7866 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6357) );
  AND4_X1 U7867 ( .A1(n6358), .A2(n6402), .A3(n6357), .A4(n6416), .ZN(n6241)
         );
  AND2_X1 U7868 ( .A1(n6356), .A2(n6241), .ZN(n6389) );
  NAND2_X1 U7869 ( .A1(n6389), .A2(n6242), .ZN(n6432) );
  NAND2_X1 U7870 ( .A1(n6243), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6444) );
  INV_X1 U7871 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7872 ( .A1(n6444), .A2(n6244), .ZN(n6245) );
  NAND2_X1 U7873 ( .A1(n6245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6270) );
  INV_X1 U7874 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7875 ( .A1(n6270), .A2(n6246), .ZN(n6247) );
  NAND2_X1 U7876 ( .A1(n6247), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6248) );
  XNOR2_X1 U7877 ( .A(n6248), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8641) );
  AOI22_X1 U7878 ( .A1(n6446), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6445), .B2(
        n8641), .ZN(n6249) );
  NAND2_X1 U7879 ( .A1(n6393), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6256) );
  INV_X1 U7880 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8997) );
  OR2_X1 U7881 ( .A1(n6340), .A2(n8997), .ZN(n6255) );
  INV_X1 U7882 ( .A(n6251), .ZN(n6263) );
  NAND2_X1 U7883 ( .A1(n6275), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6252) );
  AND2_X1 U7884 ( .A1(n6263), .A2(n6252), .ZN(n8888) );
  OR2_X1 U7885 ( .A1(n4517), .A2(n8888), .ZN(n6254) );
  INV_X1 U7886 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8887) );
  OR2_X1 U7887 ( .A1(n6339), .A2(n8887), .ZN(n6253) );
  NAND2_X1 U7888 ( .A1(n9084), .A2(n8399), .ZN(n6580) );
  NAND2_X1 U7889 ( .A1(n7197), .A2(n6431), .ZN(n6262) );
  NAND2_X1 U7890 ( .A1(n6257), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6258) );
  MUX2_X1 U7891 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6258), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6260) );
  AND2_X1 U7892 ( .A1(n6260), .A2(n6259), .ZN(n8644) );
  AOI22_X1 U7893 ( .A1(n6446), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6445), .B2(
        n8644), .ZN(n6261) );
  NAND2_X1 U7894 ( .A1(n6393), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6269) );
  INV_X1 U7895 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8994) );
  OR2_X1 U7896 ( .A1(n6340), .A2(n8994), .ZN(n6268) );
  NAND2_X1 U7897 ( .A1(n6263), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6264) );
  AND2_X1 U7898 ( .A1(n6265), .A2(n6264), .ZN(n8877) );
  OR2_X1 U7899 ( .A1(n4517), .A2(n8877), .ZN(n6267) );
  INV_X1 U7900 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8876) );
  OR2_X1 U7901 ( .A1(n6339), .A2(n8876), .ZN(n6266) );
  NAND4_X1 U7902 ( .A1(n6269), .A2(n6268), .A3(n6267), .A4(n6266), .ZN(n8885)
         );
  AND2_X1 U7903 ( .A1(n8461), .A2(n8885), .ZN(n6579) );
  INV_X1 U7904 ( .A(n6579), .ZN(n6575) );
  INV_X1 U7905 ( .A(n8885), .ZN(n8543) );
  NAND2_X1 U7906 ( .A1(n9078), .A2(n8543), .ZN(n6582) );
  NAND2_X1 U7907 ( .A1(n6575), .A2(n6582), .ZN(n8873) );
  NAND2_X1 U7908 ( .A1(n7016), .A2(n6431), .ZN(n6272) );
  XNOR2_X1 U7909 ( .A(n6270), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8602) );
  AOI22_X1 U7910 ( .A1(n6446), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6445), .B2(
        n8602), .ZN(n6271) );
  NAND2_X1 U7911 ( .A1(n6393), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6279) );
  INV_X1 U7912 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6273) );
  OR2_X1 U7913 ( .A1(n6339), .A2(n6273), .ZN(n6278) );
  INV_X1 U7914 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9000) );
  OR2_X1 U7915 ( .A1(n6340), .A2(n9000), .ZN(n6277) );
  NAND2_X1 U7916 ( .A1(n6451), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6274) );
  AND2_X1 U7917 ( .A1(n6275), .A2(n6274), .ZN(n8900) );
  OR2_X1 U7918 ( .A1(n4517), .A2(n8900), .ZN(n6276) );
  OR2_X1 U7919 ( .A1(n9090), .A2(n8496), .ZN(n6570) );
  NAND2_X1 U7920 ( .A1(n9090), .A2(n8496), .ZN(n6569) );
  NAND2_X1 U7921 ( .A1(n6393), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6286) );
  INV_X1 U7922 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7732) );
  OR2_X1 U7923 ( .A1(n6339), .A2(n7732), .ZN(n6285) );
  INV_X1 U7924 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6280) );
  OR2_X1 U7925 ( .A1(n6340), .A2(n6280), .ZN(n6284) );
  INV_X1 U7926 ( .A(n6281), .ZN(n6324) );
  NAND2_X1 U7927 ( .A1(n6324), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6282) );
  AND2_X1 U7928 ( .A1(n6374), .A2(n6282), .ZN(n7733) );
  OR2_X1 U7929 ( .A1(n4517), .A2(n7733), .ZN(n6283) );
  NAND2_X1 U7930 ( .A1(n6287), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6288) );
  XNOR2_X1 U7931 ( .A(n6288), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7360) );
  OR2_X1 U7932 ( .A1(n6346), .A2(n6849), .ZN(n6290) );
  INV_X1 U7933 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6848) );
  OR2_X1 U7934 ( .A1(n4515), .A2(n6848), .ZN(n6289) );
  OAI211_X1 U7935 ( .C1(n6795), .C2(n7342), .A(n6290), .B(n6289), .ZN(n7735)
         );
  XNOR2_X1 U7936 ( .A(n8562), .B(n10048), .ZN(n7726) );
  NAND2_X1 U7937 ( .A1(n6393), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6294) );
  INV_X1 U7938 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7446) );
  OR2_X1 U7939 ( .A1(n6339), .A2(n7446), .ZN(n6293) );
  INV_X1 U7940 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6798) );
  OR2_X1 U7941 ( .A1(n6340), .A2(n6798), .ZN(n6292) );
  OR2_X1 U7942 ( .A1(n4517), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6291) );
  OR2_X1 U7943 ( .A1(n6295), .A2(n6096), .ZN(n6297) );
  INV_X1 U7944 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6855) );
  OR2_X1 U7945 ( .A1(n4515), .A2(n6855), .ZN(n6299) );
  OR2_X1 U7946 ( .A1(n6346), .A2(n6854), .ZN(n6298) );
  OAI211_X1 U7947 ( .C1(n6795), .C2(n7015), .A(n6299), .B(n6298), .ZN(n7448)
         );
  NAND2_X1 U7948 ( .A1(n8929), .A2(n7448), .ZN(n6525) );
  INV_X1 U7949 ( .A(n8929), .ZN(n8563) );
  NAND2_X1 U7950 ( .A1(n8563), .A2(n10038), .ZN(n6518) );
  AND2_X1 U7951 ( .A1(n6525), .A2(n6518), .ZN(n6467) );
  INV_X1 U7952 ( .A(n6467), .ZN(n7443) );
  INV_X1 U7953 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6301) );
  INV_X1 U7954 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6302) );
  INV_X1 U7955 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6303) );
  INV_X1 U7956 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6857) );
  OR2_X1 U7957 ( .A1(n4515), .A2(n6857), .ZN(n6308) );
  OR2_X1 U7958 ( .A1(n6346), .A2(n6856), .ZN(n6306) );
  AND2_X1 U7959 ( .A1(n6306), .A2(n5142), .ZN(n6307) );
  INV_X1 U7960 ( .A(n10032), .ZN(n7200) );
  NAND4_X1 U7961 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n8564)
         );
  NAND2_X1 U7962 ( .A1(n7200), .A2(n8564), .ZN(n6509) );
  AND2_X2 U7963 ( .A1(n7441), .A2(n6509), .ZN(n6465) );
  NAND2_X1 U7964 ( .A1(n6393), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6317) );
  INV_X1 U7965 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10384) );
  OR2_X1 U7966 ( .A1(n4517), .A2(n10384), .ZN(n6316) );
  INV_X1 U7967 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6313) );
  OR2_X1 U7968 ( .A1(n6339), .A2(n6313), .ZN(n6315) );
  NAND2_X1 U7969 ( .A1(n6372), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6314) );
  NAND4_X1 U7970 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n6322)
         );
  INV_X1 U7971 ( .A(n6322), .ZN(n6321) );
  INV_X1 U7972 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U7973 ( .A1(n6318), .A2(SI_0_), .ZN(n6320) );
  XNOR2_X1 U7974 ( .A(n6320), .B(n6319), .ZN(n9124) );
  MUX2_X1 U7975 ( .A(n6825), .B(n9124), .S(n6795), .Z(n7167) );
  INV_X1 U7976 ( .A(n7167), .ZN(n8339) );
  NAND2_X1 U7977 ( .A1(n6321), .A2(n8339), .ZN(n7091) );
  CLKBUF_X1 U7978 ( .A(n6322), .Z(n8566) );
  NAND2_X1 U7979 ( .A1(n6322), .A2(n7167), .ZN(n6505) );
  AND2_X1 U7980 ( .A1(n7091), .A2(n6505), .ZN(n7165) );
  NAND2_X1 U7981 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6323) );
  AND2_X1 U7982 ( .A1(n6324), .A2(n6323), .ZN(n7504) );
  OR2_X1 U7983 ( .A1(n4517), .A2(n7504), .ZN(n6331) );
  NAND2_X1 U7984 ( .A1(n6300), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6329) );
  INV_X1 U7985 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6325) );
  OR2_X1 U7986 ( .A1(n4513), .A2(n6325), .ZN(n6328) );
  INV_X1 U7987 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6326) );
  OR2_X1 U7988 ( .A1(n6340), .A2(n6326), .ZN(n6327) );
  OR2_X1 U7989 ( .A1(n4515), .A2(n5206), .ZN(n6336) );
  OR2_X1 U7990 ( .A1(n6346), .A2(n6858), .ZN(n6335) );
  OR2_X1 U7991 ( .A1(n6240), .A2(n6096), .ZN(n6333) );
  OR2_X1 U7992 ( .A1(n6795), .A2(n7178), .ZN(n6334) );
  NAND3_X1 U7993 ( .A1(n6465), .A2(n7165), .A3(n7501), .ZN(n6347) );
  NAND2_X1 U7994 ( .A1(n6393), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6343) );
  INV_X1 U7995 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9994) );
  INV_X1 U7996 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7305) );
  NAND2_X1 U7997 ( .A1(n6372), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6341) );
  OAI22_X1 U7998 ( .A1(n6344), .A2(n5186), .B1(n6795), .B2(n9998), .ZN(n6345)
         );
  NAND2_X1 U7999 ( .A1(n6507), .A2(n6502), .ZN(n6677) );
  NOR4_X1 U8000 ( .A1(n7726), .A2(n7443), .A3(n6347), .A4(n6677), .ZN(n6388)
         );
  NAND2_X1 U8001 ( .A1(n6393), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6355) );
  INV_X1 U8002 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6348) );
  OR2_X1 U8003 ( .A1(n6340), .A2(n6348), .ZN(n6354) );
  INV_X1 U8004 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7899) );
  OR2_X1 U8005 ( .A1(n6339), .A2(n7899), .ZN(n6353) );
  INV_X1 U8006 ( .A(n6349), .ZN(n6408) );
  INV_X1 U8007 ( .A(n6350), .ZN(n6362) );
  NAND2_X1 U8008 ( .A1(n6362), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6351) );
  AND2_X1 U8009 ( .A1(n6408), .A2(n6351), .ZN(n7960) );
  OR2_X1 U8010 ( .A1(n4517), .A2(n7960), .ZN(n6352) );
  NAND4_X1 U8011 ( .A1(n6355), .A2(n6354), .A3(n6353), .A4(n6352), .ZN(n8559)
         );
  NAND2_X1 U8012 ( .A1(n6400), .A2(n6357), .ZN(n6368) );
  NAND2_X1 U8013 ( .A1(n6368), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6359) );
  INV_X1 U8014 ( .A(n7822), .ZN(n7698) );
  NAND2_X1 U8015 ( .A1(n10059), .A2(n8559), .ZN(n6545) );
  NAND2_X1 U8016 ( .A1(n6393), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6366) );
  INV_X1 U8017 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7796) );
  OR2_X1 U8018 ( .A1(n6339), .A2(n7796), .ZN(n6365) );
  INV_X1 U8019 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6360) );
  OR2_X1 U8020 ( .A1(n6340), .A2(n6360), .ZN(n6364) );
  NAND2_X1 U8021 ( .A1(n6376), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6361) );
  AND2_X1 U8022 ( .A1(n6362), .A2(n6361), .ZN(n7865) );
  OR2_X1 U8023 ( .A1(n4517), .A2(n7865), .ZN(n6363) );
  INV_X1 U8024 ( .A(n6400), .ZN(n6367) );
  NAND2_X1 U8025 ( .A1(n6367), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6369) );
  INV_X1 U8026 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6859) );
  OR2_X1 U8027 ( .A1(n4515), .A2(n6859), .ZN(n6370) );
  OAI211_X1 U8028 ( .C1(n6795), .C2(n7711), .A(n6371), .B(n6370), .ZN(n7860)
         );
  NAND2_X1 U8029 ( .A1(n7854), .A2(n7860), .ZN(n6540) );
  INV_X1 U8030 ( .A(n7860), .ZN(n10053) );
  NAND2_X1 U8031 ( .A1(n8560), .A2(n10053), .ZN(n6544) );
  NAND2_X1 U8032 ( .A1(n6540), .A2(n6544), .ZN(n7790) );
  INV_X1 U8033 ( .A(n7790), .ZN(n6387) );
  NAND2_X1 U8034 ( .A1(n6372), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6380) );
  INV_X1 U8035 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6373) );
  OR2_X1 U8036 ( .A1(n4513), .A2(n6373), .ZN(n6379) );
  NAND2_X1 U8037 ( .A1(n6374), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6375) );
  AND2_X1 U8038 ( .A1(n6376), .A2(n6375), .ZN(n7685) );
  OR2_X1 U8039 ( .A1(n4517), .A2(n7685), .ZN(n6378) );
  INV_X1 U8040 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7684) );
  OR2_X1 U8041 ( .A1(n6339), .A2(n7684), .ZN(n6377) );
  NAND4_X1 U8042 ( .A1(n6380), .A2(n6379), .A3(n6378), .A4(n6377), .ZN(n8561)
         );
  OR2_X1 U8043 ( .A1(n6346), .A2(n6852), .ZN(n6386) );
  INV_X1 U8044 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6850) );
  OR2_X1 U8045 ( .A1(n4515), .A2(n6850), .ZN(n6385) );
  NAND2_X1 U8046 ( .A1(n6381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6383) );
  INV_X1 U8047 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U8048 ( .A(n6383), .B(n6382), .ZN(n7700) );
  OR2_X1 U8049 ( .A1(n6795), .A2(n7700), .ZN(n6384) );
  INV_X1 U8050 ( .A(n7754), .ZN(n7687) );
  XNOR2_X1 U8051 ( .A(n8561), .B(n7687), .ZN(n7682) );
  NAND4_X1 U8052 ( .A1(n6388), .A2(n7897), .A3(n6387), .A4(n7682), .ZN(n6430)
         );
  NAND2_X1 U8053 ( .A1(n6884), .A2(n6431), .ZN(n6392) );
  OR2_X1 U8054 ( .A1(n6389), .A2(n6096), .ZN(n6390) );
  XNOR2_X1 U8055 ( .A(n6390), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8097) );
  AOI22_X1 U8056 ( .A1(n6446), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6445), .B2(
        n8097), .ZN(n6391) );
  NAND2_X1 U8057 ( .A1(n6392), .A2(n6391), .ZN(n8208) );
  NAND2_X1 U8058 ( .A1(n6393), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6398) );
  INV_X1 U8059 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8058) );
  OR2_X1 U8060 ( .A1(n6339), .A2(n8058), .ZN(n6397) );
  INV_X1 U8061 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8057) );
  OR2_X1 U8062 ( .A1(n6340), .A2(n8057), .ZN(n6396) );
  NAND2_X1 U8063 ( .A1(n6424), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6394) );
  AND2_X1 U8064 ( .A1(n6437), .A2(n6394), .ZN(n8044) );
  OR2_X1 U8065 ( .A1(n4517), .A2(n8044), .ZN(n6395) );
  OR2_X1 U8066 ( .A1(n8208), .A2(n8191), .ZN(n6555) );
  NAND2_X1 U8067 ( .A1(n8208), .A2(n8191), .ZN(n6557) );
  INV_X1 U8068 ( .A(n8199), .ZN(n6429) );
  NAND2_X1 U8069 ( .A1(n6873), .A2(n6431), .ZN(n6406) );
  OAI21_X1 U8070 ( .B1(P2_IR_REG_8__SCAN_IN), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6399) );
  INV_X1 U8071 ( .A(n6403), .ZN(n6401) );
  NAND2_X1 U8072 ( .A1(n6401), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U8073 ( .A1(n6403), .A2(n6402), .ZN(n6415) );
  AOI22_X1 U8074 ( .A1(n6446), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6445), .B2(
        n7873), .ZN(n6405) );
  NAND2_X1 U8075 ( .A1(n6406), .A2(n6405), .ZN(n10067) );
  NAND2_X1 U8076 ( .A1(n6300), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6414) );
  INV_X1 U8077 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6407) );
  OR2_X1 U8078 ( .A1(n6340), .A2(n6407), .ZN(n6413) );
  NAND2_X1 U8079 ( .A1(n6408), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6409) );
  AND2_X1 U8080 ( .A1(n6422), .A2(n6409), .ZN(n8129) );
  OR2_X1 U8081 ( .A1(n4517), .A2(n8129), .ZN(n6412) );
  INV_X1 U8082 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6410) );
  OR2_X1 U8083 ( .A1(n4513), .A2(n6410), .ZN(n6411) );
  NAND2_X1 U8084 ( .A1(n10067), .A2(n8133), .ZN(n6542) );
  NAND2_X1 U8085 ( .A1(n6546), .A2(n6542), .ZN(n7932) );
  OR2_X1 U8086 ( .A1(n6879), .A2(n6346), .ZN(n6419) );
  NAND2_X1 U8087 ( .A1(n6415), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6417) );
  XNOR2_X1 U8088 ( .A(n6417), .B(n6416), .ZN(n8072) );
  INV_X1 U8089 ( .A(n8072), .ZN(n7888) );
  AOI22_X1 U8090 ( .A1(n6446), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6445), .B2(
        n7888), .ZN(n6418) );
  NAND2_X1 U8091 ( .A1(n6393), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6428) );
  INV_X1 U8092 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6420) );
  OR2_X1 U8093 ( .A1(n6340), .A2(n6420), .ZN(n6427) );
  INV_X1 U8094 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6421) );
  OR2_X1 U8095 ( .A1(n6339), .A2(n6421), .ZN(n6426) );
  NAND2_X1 U8096 ( .A1(n6422), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6423) );
  AND2_X1 U8097 ( .A1(n6424), .A2(n6423), .ZN(n8187) );
  OR2_X1 U8098 ( .A1(n4517), .A2(n8187), .ZN(n6425) );
  NAND2_X1 U8099 ( .A1(n10071), .A2(n8196), .ZN(n6553) );
  NAND2_X1 U8100 ( .A1(n6551), .A2(n6553), .ZN(n8029) );
  NOR4_X1 U8101 ( .A1(n6430), .A2(n6429), .A3(n7932), .A4(n8029), .ZN(n6456)
         );
  NAND2_X1 U8102 ( .A1(n6968), .A2(n6431), .ZN(n6435) );
  NAND2_X1 U8103 ( .A1(n6432), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6433) );
  XNOR2_X1 U8104 ( .A(n6433), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8080) );
  AOI22_X1 U8105 ( .A1(n6446), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6445), .B2(
        n8080), .ZN(n6434) );
  NAND2_X1 U8106 ( .A1(n6300), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6443) );
  INV_X1 U8107 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8067) );
  OR2_X1 U8108 ( .A1(n6340), .A2(n8067), .ZN(n6442) );
  INV_X1 U8109 ( .A(n6436), .ZN(n6449) );
  NAND2_X1 U8110 ( .A1(n6437), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6438) );
  AND2_X1 U8111 ( .A1(n6449), .A2(n6438), .ZN(n8443) );
  OR2_X1 U8112 ( .A1(n4517), .A2(n8443), .ZN(n6441) );
  INV_X1 U8113 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6439) );
  OR2_X1 U8114 ( .A1(n4513), .A2(n6439), .ZN(n6440) );
  NAND4_X1 U8115 ( .A1(n6443), .A2(n6442), .A3(n6441), .A4(n6440), .ZN(n8912)
         );
  XNOR2_X1 U8116 ( .A(n10084), .B(n8912), .ZN(n8171) );
  OR2_X1 U8117 ( .A1(n6979), .A2(n6346), .ZN(n6448) );
  XNOR2_X1 U8118 ( .A(n6444), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8599) );
  AOI22_X1 U8119 ( .A1(n6446), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6445), .B2(
        n8599), .ZN(n6447) );
  NAND2_X1 U8120 ( .A1(n6393), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6455) );
  INV_X1 U8121 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8571) );
  OR2_X1 U8122 ( .A1(n6339), .A2(n8571), .ZN(n6454) );
  INV_X1 U8123 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9003) );
  OR2_X1 U8124 ( .A1(n6340), .A2(n9003), .ZN(n6453) );
  NAND2_X1 U8125 ( .A1(n6449), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6450) );
  AND2_X1 U8126 ( .A1(n6451), .A2(n6450), .ZN(n8918) );
  OR2_X1 U8127 ( .A1(n4517), .A2(n8918), .ZN(n6452) );
  NAND4_X1 U8128 ( .A1(n6455), .A2(n6454), .A3(n6453), .A4(n6452), .ZN(n8896)
         );
  XNOR2_X1 U8129 ( .A(n9097), .B(n8896), .ZN(n8908) );
  NAND4_X1 U8130 ( .A1(n8895), .A2(n6456), .A3(n8171), .A4(n8908), .ZN(n6457)
         );
  NOR4_X1 U8131 ( .A1(n8863), .A2(n8881), .A3(n8873), .A4(n6457), .ZN(n6458)
         );
  NAND4_X1 U8132 ( .A1(n8826), .A2(n8839), .A3(n8849), .A4(n6458), .ZN(n6459)
         );
  NOR4_X1 U8133 ( .A1(n8786), .A2(n8801), .A3(n8814), .A4(n6459), .ZN(n6460)
         );
  NAND4_X1 U8134 ( .A1(n8749), .A2(n8756), .A3(n8775), .A4(n6460), .ZN(n6461)
         );
  NOR4_X1 U8135 ( .A1(n6647), .A2(n8731), .A3(n8720), .A4(n6461), .ZN(n6462)
         );
  NAND2_X1 U8136 ( .A1(n9008), .A2(n8553), .ZN(n6656) );
  AND2_X1 U8137 ( .A1(n8949), .A2(n8554), .ZN(n6648) );
  INV_X1 U8138 ( .A(n6648), .ZN(n6652) );
  NAND4_X1 U8139 ( .A1(n6463), .A2(n6462), .A3(n6656), .A4(n6652), .ZN(n6493)
         );
  NAND2_X1 U8140 ( .A1(n6507), .A2(n7091), .ZN(n6464) );
  NAND2_X1 U8141 ( .A1(n6464), .A2(n6502), .ZN(n8924) );
  INV_X1 U8142 ( .A(n8924), .ZN(n6466) );
  NAND2_X1 U8143 ( .A1(n7440), .A2(n7441), .ZN(n6468) );
  NAND2_X1 U8144 ( .A1(n6468), .A2(n6467), .ZN(n7439) );
  NAND2_X1 U8145 ( .A1(n7439), .A2(n6525), .ZN(n6469) );
  NAND2_X1 U8146 ( .A1(n7727), .A2(n7506), .ZN(n6519) );
  NAND2_X1 U8147 ( .A1(n7590), .A2(n7735), .ZN(n6530) );
  INV_X1 U8148 ( .A(n6530), .ZN(n6470) );
  NAND2_X1 U8149 ( .A1(n8562), .A2(n10048), .ZN(n6527) );
  NAND2_X1 U8150 ( .A1(n8561), .A2(n7754), .ZN(n6521) );
  INV_X1 U8151 ( .A(n6521), .ZN(n6532) );
  NOR2_X1 U8152 ( .A1(n8561), .A2(n7754), .ZN(n6522) );
  INV_X1 U8153 ( .A(n6522), .ZN(n6531) );
  INV_X1 U8154 ( .A(n6545), .ZN(n6471) );
  NAND2_X1 U8155 ( .A1(n6472), .A2(n6553), .ZN(n8043) );
  INV_X1 U8156 ( .A(n8171), .ZN(n8174) );
  INV_X1 U8157 ( .A(n8912), .ZN(n8206) );
  NOR2_X1 U8158 ( .A1(n10084), .A2(n8206), .ZN(n6559) );
  INV_X1 U8159 ( .A(n6559), .ZN(n6473) );
  INV_X1 U8160 ( .A(n8896), .ZN(n8439) );
  NOR2_X1 U8161 ( .A1(n9097), .A2(n8439), .ZN(n6474) );
  INV_X1 U8162 ( .A(n9097), .ZN(n8916) );
  NAND2_X1 U8163 ( .A1(n6475), .A2(n6569), .ZN(n8882) );
  INV_X1 U8164 ( .A(n8882), .ZN(n6476) );
  NAND2_X1 U8165 ( .A1(n6476), .A2(n6580), .ZN(n6477) );
  INV_X1 U8166 ( .A(n6583), .ZN(n6478) );
  NAND2_X1 U8167 ( .A1(n6500), .A2(n8813), .ZN(n6606) );
  INV_X1 U8168 ( .A(n6606), .ZN(n6479) );
  NAND2_X1 U8169 ( .A1(n8812), .A2(n6479), .ZN(n6480) );
  AND2_X1 U8170 ( .A1(n6622), .A2(n8771), .ZN(n6624) );
  NAND2_X1 U8171 ( .A1(n6483), .A2(n6633), .ZN(n8732) );
  NOR2_X1 U8172 ( .A1(n8743), .A2(n8530), .ZN(n6635) );
  INV_X1 U8173 ( .A(n6635), .ZN(n6484) );
  INV_X1 U8174 ( .A(n8736), .ZN(n8393) );
  OR2_X1 U8175 ( .A1(n9016), .A2(n8393), .ZN(n6485) );
  OAI21_X1 U8176 ( .B1(n6648), .B2(n8553), .A(n9008), .ZN(n6488) );
  INV_X1 U8177 ( .A(n6490), .ZN(n6496) );
  NAND2_X1 U8178 ( .A1(n6496), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6491) );
  MUX2_X1 U8179 ( .A(n6493), .B(n6492), .S(n7300), .Z(n6657) );
  NAND2_X1 U8180 ( .A1(n6494), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6495) );
  MUX2_X1 U8181 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6495), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6497) );
  NAND2_X1 U8182 ( .A1(n6498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6499) );
  MUX2_X1 U8183 ( .A(n8736), .B(n9016), .S(n6792), .Z(n6643) );
  OAI21_X1 U8184 ( .B1(n6792), .B2(n6500), .A(n8795), .ZN(n6615) );
  NAND2_X1 U8185 ( .A1(n6502), .A2(n6505), .ZN(n6501) );
  NAND2_X1 U8186 ( .A1(n6507), .A2(n6501), .ZN(n6504) );
  INV_X1 U8187 ( .A(n6502), .ZN(n6503) );
  NAND2_X1 U8188 ( .A1(n6505), .A2(n7300), .ZN(n6506) );
  NAND4_X1 U8189 ( .A1(n6507), .A2(n7091), .A3(n6792), .A4(n6506), .ZN(n6508)
         );
  NAND2_X1 U8190 ( .A1(n6465), .A2(n6508), .ZN(n6515) );
  NAND2_X1 U8191 ( .A1(n6518), .A2(n6509), .ZN(n6510) );
  NAND2_X1 U8192 ( .A1(n6525), .A2(n7441), .ZN(n6511) );
  OAI21_X2 U8193 ( .B1(n6516), .B2(n6515), .A(n6514), .ZN(n6517) );
  NAND2_X1 U8194 ( .A1(n6517), .A2(n7501), .ZN(n6529) );
  INV_X1 U8195 ( .A(n6518), .ZN(n6520) );
  OAI211_X1 U8196 ( .C1(n6529), .C2(n6520), .A(n6519), .B(n6530), .ZN(n6524)
         );
  AND2_X1 U8197 ( .A1(n6521), .A2(n6527), .ZN(n6523) );
  AOI21_X1 U8198 ( .B1(n6524), .B2(n6523), .A(n6522), .ZN(n6536) );
  INV_X1 U8199 ( .A(n6525), .ZN(n7497) );
  NAND2_X1 U8200 ( .A1(n6526), .A2(n10044), .ZN(n6528) );
  OAI211_X1 U8201 ( .C1(n6529), .C2(n7497), .A(n6528), .B(n6527), .ZN(n6534)
         );
  AND2_X1 U8202 ( .A1(n6531), .A2(n6530), .ZN(n6533) );
  AOI21_X1 U8203 ( .B1(n6534), .B2(n6533), .A(n6532), .ZN(n6535) );
  NAND2_X1 U8204 ( .A1(n6546), .A2(n6545), .ZN(n6538) );
  NAND2_X1 U8205 ( .A1(n6542), .A2(n6541), .ZN(n6537) );
  NOR2_X1 U8206 ( .A1(n6548), .A2(n7790), .ZN(n6539) );
  AND2_X1 U8207 ( .A1(n6541), .A2(n6540), .ZN(n6543) );
  AND2_X1 U8208 ( .A1(n6545), .A2(n6544), .ZN(n6547) );
  NAND2_X1 U8209 ( .A1(n6550), .A2(n6549), .ZN(n6554) );
  AND2_X1 U8210 ( .A1(n6555), .A2(n6551), .ZN(n6552) );
  AOI21_X1 U8211 ( .B1(n6554), .B2(n6552), .A(n4691), .ZN(n6558) );
  NAND2_X1 U8212 ( .A1(n6554), .A2(n6553), .ZN(n6556) );
  AND2_X1 U8213 ( .A1(n10084), .A2(n8206), .ZN(n6560) );
  MUX2_X1 U8214 ( .A(n6560), .B(n6559), .S(n6741), .Z(n6561) );
  INV_X1 U8215 ( .A(n6561), .ZN(n6562) );
  NAND2_X1 U8216 ( .A1(n6563), .A2(n6562), .ZN(n6566) );
  NAND2_X1 U8217 ( .A1(n8916), .A2(n8439), .ZN(n6705) );
  MUX2_X1 U8218 ( .A(n9097), .B(n8896), .S(n6792), .Z(n6564) );
  INV_X1 U8219 ( .A(n6564), .ZN(n6565) );
  OAI21_X1 U8220 ( .B1(n6566), .B2(n6705), .A(n6565), .ZN(n6567) );
  NAND2_X1 U8221 ( .A1(n9097), .A2(n8896), .ZN(n6703) );
  NAND2_X1 U8222 ( .A1(n6568), .A2(n8895), .ZN(n6572) );
  MUX2_X1 U8223 ( .A(n6570), .B(n6569), .S(n6792), .Z(n6571) );
  NAND2_X1 U8224 ( .A1(n6572), .A2(n6571), .ZN(n6573) );
  NAND2_X1 U8225 ( .A1(n6573), .A2(n8883), .ZN(n6581) );
  AND2_X1 U8226 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  AOI21_X1 U8227 ( .B1(n6581), .B2(n6576), .A(n4955), .ZN(n6600) );
  NAND4_X1 U8228 ( .A1(n6603), .A2(n6741), .A3(n6578), .A4(n6577), .ZN(n6599)
         );
  AOI21_X1 U8229 ( .B1(n6581), .B2(n6580), .A(n6579), .ZN(n6586) );
  NAND4_X1 U8230 ( .A1(n6584), .A2(n6792), .A3(n6583), .A4(n6582), .ZN(n6585)
         );
  OR2_X1 U8231 ( .A1(n6586), .A2(n6585), .ZN(n6598) );
  NOR2_X1 U8232 ( .A1(n8874), .A2(n6792), .ZN(n6587) );
  NAND2_X1 U8233 ( .A1(n9072), .A2(n6587), .ZN(n6590) );
  OAI21_X1 U8234 ( .B1(n8864), .B2(n6792), .A(n6590), .ZN(n6588) );
  NAND2_X1 U8235 ( .A1(n6588), .A2(n8988), .ZN(n6589) );
  OAI21_X1 U8236 ( .B1(n6590), .B2(n8864), .A(n6589), .ZN(n6596) );
  INV_X1 U8237 ( .A(n8988), .ZN(n8522) );
  NAND2_X1 U8238 ( .A1(n8874), .A2(n6792), .ZN(n6592) );
  OAI22_X1 U8239 ( .A1(n9072), .A2(n6592), .B1(n6741), .B2(n8466), .ZN(n6591)
         );
  NAND2_X1 U8240 ( .A1(n8522), .A2(n6591), .ZN(n6594) );
  OR3_X1 U8241 ( .A1(n9072), .A2(n8466), .A3(n6592), .ZN(n6593) );
  NAND2_X1 U8242 ( .A1(n6594), .A2(n6593), .ZN(n6595) );
  AOI21_X1 U8243 ( .B1(n6603), .B2(n6596), .A(n6595), .ZN(n6597) );
  OAI211_X1 U8244 ( .C1(n6600), .C2(n6599), .A(n6598), .B(n6597), .ZN(n6602)
         );
  MUX2_X1 U8245 ( .A(n6741), .B(n6602), .S(n6601), .Z(n6609) );
  NAND2_X1 U8246 ( .A1(n6610), .A2(n6603), .ZN(n6604) );
  NAND2_X1 U8247 ( .A1(n6604), .A2(n6792), .ZN(n6605) );
  NAND2_X1 U8248 ( .A1(n6605), .A2(n8813), .ZN(n6608) );
  NAND2_X1 U8249 ( .A1(n6606), .A2(n6792), .ZN(n6607) );
  OAI21_X1 U8250 ( .B1(n6609), .B2(n6608), .A(n6607), .ZN(n6613) );
  AOI21_X1 U8251 ( .B1(n6612), .B2(n6610), .A(n6792), .ZN(n6611) );
  AOI21_X1 U8252 ( .B1(n6613), .B2(n6612), .A(n6611), .ZN(n6614) );
  NAND2_X1 U8253 ( .A1(n8771), .A2(n6616), .ZN(n6617) );
  MUX2_X1 U8254 ( .A(n6618), .B(n6617), .S(n6792), .Z(n6619) );
  NAND2_X1 U8255 ( .A1(n6625), .A2(n6620), .ZN(n6623) );
  AOI21_X1 U8256 ( .B1(n6623), .B2(n6622), .A(n6621), .ZN(n6627) );
  MUX2_X1 U8257 ( .A(n6629), .B(n6628), .S(n6792), .Z(n6630) );
  OAI211_X1 U8258 ( .C1(n6631), .C2(n8758), .A(n8749), .B(n6630), .ZN(n6639)
         );
  MUX2_X1 U8259 ( .A(n6633), .B(n6632), .S(n6741), .Z(n6634) );
  AND2_X1 U8260 ( .A1(n8734), .A2(n6634), .ZN(n6638) );
  AND2_X1 U8261 ( .A1(n8743), .A2(n8530), .ZN(n6636) );
  MUX2_X1 U8262 ( .A(n6636), .B(n6635), .S(n6792), .Z(n6637) );
  INV_X1 U8263 ( .A(n6643), .ZN(n6644) );
  NOR2_X1 U8264 ( .A1(n6645), .A2(n6644), .ZN(n6650) );
  NOR2_X1 U8265 ( .A1(n6650), .A2(n6741), .ZN(n6654) );
  XNOR2_X1 U8266 ( .A(n6658), .B(n8705), .ZN(n6676) );
  INV_X1 U8267 ( .A(n6793), .ZN(n6820) );
  NAND2_X1 U8268 ( .A1(n6820), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7928) );
  NAND2_X1 U8269 ( .A1(n6661), .A2(n6660), .ZN(n6662) );
  NAND2_X1 U8270 ( .A1(n6665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6666) );
  NOR2_X1 U8271 ( .A1(n9120), .A2(n6749), .ZN(n6671) );
  NAND2_X1 U8272 ( .A1(n7652), .A2(n7531), .ZN(n7086) );
  NOR2_X1 U8273 ( .A1(n9102), .A2(n7217), .ZN(n7106) );
  INV_X1 U8274 ( .A(n4516), .ZN(n6806) );
  NAND3_X1 U8275 ( .A1(n7106), .A2(n6806), .A3(n8699), .ZN(n6674) );
  OAI211_X1 U8276 ( .C1(n7919), .C2(n7928), .A(n6674), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6675) );
  OAI21_X1 U8277 ( .B1(n6676), .B2(n7928), .A(n6675), .ZN(P2_U3296) );
  INV_X1 U8278 ( .A(n9016), .ZN(n6729) );
  NAND2_X1 U8279 ( .A1(n8566), .A2(n8339), .ZN(n7303) );
  NAND2_X1 U8280 ( .A1(n6677), .A2(n7303), .ZN(n6681) );
  NAND2_X1 U8281 ( .A1(n6678), .A2(n6679), .ZN(n6680) );
  NAND2_X1 U8282 ( .A1(n6681), .A2(n6680), .ZN(n8931) );
  NAND2_X1 U8283 ( .A1(n8931), .A2(n8925), .ZN(n6684) );
  NAND2_X1 U8284 ( .A1(n6682), .A2(n7200), .ZN(n6683) );
  NAND2_X1 U8285 ( .A1(n6684), .A2(n6683), .ZN(n7444) );
  AND2_X1 U8286 ( .A1(n8929), .A2(n10038), .ZN(n6685) );
  NAND2_X1 U8287 ( .A1(n7502), .A2(n6686), .ZN(n6688) );
  NAND2_X1 U8288 ( .A1(n6688), .A2(n6687), .ZN(n7725) );
  NAND2_X1 U8289 ( .A1(n7590), .A2(n10048), .ZN(n6689) );
  OR2_X1 U8290 ( .A1(n7590), .A2(n10048), .ZN(n6690) );
  INV_X1 U8291 ( .A(n8561), .ZN(n7792) );
  NAND2_X1 U8292 ( .A1(n7792), .A2(n7754), .ZN(n6691) );
  NAND2_X1 U8293 ( .A1(n6692), .A2(n6691), .ZN(n7791) );
  AND2_X1 U8294 ( .A1(n7854), .A2(n10053), .ZN(n6694) );
  INV_X1 U8295 ( .A(n8133), .ZN(n8558) );
  OR2_X1 U8296 ( .A1(n8558), .A2(n10067), .ZN(n6695) );
  NAND2_X1 U8297 ( .A1(n5146), .A2(n6695), .ZN(n8030) );
  INV_X1 U8298 ( .A(n8196), .ZN(n8557) );
  NAND2_X1 U8299 ( .A1(n10071), .A2(n8557), .ZN(n6696) );
  NAND2_X1 U8300 ( .A1(n8030), .A2(n6696), .ZN(n6698) );
  OR2_X1 U8301 ( .A1(n10071), .A2(n8557), .ZN(n6697) );
  INV_X1 U8302 ( .A(n8191), .ZN(n8556) );
  NAND2_X1 U8303 ( .A1(n8208), .A2(n8556), .ZN(n6699) );
  OR2_X1 U8304 ( .A1(n10084), .A2(n8912), .ZN(n6700) );
  NAND2_X1 U8305 ( .A1(n8173), .A2(n6700), .ZN(n6702) );
  NAND2_X1 U8306 ( .A1(n10084), .A2(n8912), .ZN(n6701) );
  NAND2_X1 U8307 ( .A1(n6702), .A2(n6701), .ZN(n8907) );
  INV_X1 U8308 ( .A(n8907), .ZN(n6704) );
  NAND2_X1 U8309 ( .A1(n6704), .A2(n6703), .ZN(n6706) );
  NAND2_X1 U8310 ( .A1(n6706), .A2(n6705), .ZN(n8894) );
  NOR2_X1 U8311 ( .A1(n9090), .A2(n8910), .ZN(n6708) );
  NAND2_X1 U8312 ( .A1(n9090), .A2(n8910), .ZN(n6707) );
  NAND2_X1 U8313 ( .A1(n8884), .A2(n8881), .ZN(n6710) );
  NAND2_X1 U8314 ( .A1(n9084), .A2(n8897), .ZN(n6709) );
  NAND2_X1 U8315 ( .A1(n6710), .A2(n6709), .ZN(n8872) );
  NAND2_X1 U8316 ( .A1(n8872), .A2(n8873), .ZN(n6712) );
  OR2_X1 U8317 ( .A1(n8461), .A2(n8543), .ZN(n6711) );
  NAND2_X1 U8318 ( .A1(n6712), .A2(n6711), .ZN(n8862) );
  NAND2_X1 U8319 ( .A1(n9072), .A2(n8874), .ZN(n6713) );
  OR2_X1 U8320 ( .A1(n8988), .A2(n8864), .ZN(n6714) );
  NAND2_X1 U8321 ( .A1(n6715), .A2(n6714), .ZN(n8840) );
  INV_X1 U8322 ( .A(n9062), .ZN(n6716) );
  INV_X1 U8323 ( .A(n8808), .ZN(n8841) );
  OR2_X1 U8324 ( .A1(n9056), .A2(n8841), .ZN(n6717) );
  NAND2_X1 U8325 ( .A1(n8796), .A2(n8801), .ZN(n6719) );
  OR2_X1 U8326 ( .A1(n8507), .A2(n8788), .ZN(n6718) );
  NOR2_X1 U8327 ( .A1(n9041), .A2(n8776), .ZN(n6721) );
  NAND2_X1 U8328 ( .A1(n9041), .A2(n8776), .ZN(n6720) );
  AND2_X1 U8329 ( .A1(n9035), .A2(n8789), .ZN(n6722) );
  NAND2_X1 U8330 ( .A1(n9023), .A2(n8760), .ZN(n6723) );
  AND2_X1 U8331 ( .A1(n8758), .A2(n6723), .ZN(n6727) );
  INV_X1 U8332 ( .A(n6723), .ZN(n6726) );
  OR2_X1 U8333 ( .A1(n9029), .A2(n8777), .ZN(n8747) );
  OR2_X1 U8334 ( .A1(n9023), .A2(n8760), .ZN(n6724) );
  AND2_X1 U8335 ( .A1(n8747), .A2(n6724), .ZN(n6725) );
  INV_X1 U8336 ( .A(n8743), .ZN(n8955) );
  NOR2_X1 U8337 ( .A1(n8955), .A2(n8530), .ZN(n6728) );
  AOI21_X1 U8338 ( .B1(n6729), .B2(n8393), .A(n8721), .ZN(n6731) );
  NOR2_X1 U8339 ( .A1(n6731), .A2(n6730), .ZN(n6734) );
  INV_X1 U8340 ( .A(n6732), .ZN(n6733) );
  XNOR2_X1 U8341 ( .A(n6734), .B(n6732), .ZN(n6736) );
  NAND2_X1 U8342 ( .A1(n7919), .A2(n8705), .ZN(n6779) );
  NAND2_X1 U8343 ( .A1(n7300), .A2(n6778), .ZN(n6735) );
  OAI211_X1 U8344 ( .C1(n7919), .C2(n7652), .A(n10073), .B(n7531), .ZN(n6738)
         );
  INV_X1 U8345 ( .A(n6738), .ZN(n6739) );
  OR2_X1 U8346 ( .A1(n4516), .A2(n8699), .ZN(n6740) );
  NAND2_X1 U8347 ( .A1(n6795), .A2(n6740), .ZN(n6742) );
  INV_X1 U8348 ( .A(n6742), .ZN(n7113) );
  AND2_X1 U8349 ( .A1(n6795), .A2(P2_B_REG_SCAN_IN), .ZN(n6743) );
  NOR2_X1 U8350 ( .A1(n8928), .A2(n6743), .ZN(n8712) );
  AOI22_X1 U8351 ( .A1(n8911), .A2(n8736), .B1(n8554), .B2(n8712), .ZN(n6744)
         );
  NAND2_X1 U8352 ( .A1(n7652), .A2(n8705), .ZN(n6781) );
  INV_X1 U8353 ( .A(n10033), .ZN(n6746) );
  NOR2_X1 U8354 ( .A1(n8328), .A2(n6746), .ZN(n6747) );
  NOR2_X2 U8355 ( .A1(n8322), .A2(n6747), .ZN(n6789) );
  NAND2_X1 U8356 ( .A1(n9120), .A2(n6749), .ZN(n6881) );
  NAND3_X1 U8357 ( .A1(n7919), .A2(n6778), .A3(n7531), .ZN(n6751) );
  NAND2_X1 U8358 ( .A1(n6792), .A2(n6751), .ZN(n6757) );
  OR2_X1 U8359 ( .A1(n6750), .A2(n6753), .ZN(n6754) );
  NAND2_X1 U8360 ( .A1(n9103), .A2(n6757), .ZN(n6756) );
  INV_X1 U8361 ( .A(n7086), .ZN(n6758) );
  OR2_X1 U8362 ( .A1(n6758), .A2(n6792), .ZN(n6759) );
  NAND2_X1 U8363 ( .A1(n6821), .A2(n6759), .ZN(n7098) );
  INV_X1 U8364 ( .A(n7109), .ZN(n6797) );
  NOR2_X1 U8365 ( .A1(n7098), .A2(n6797), .ZN(n7211) );
  NOR2_X1 U8366 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6763) );
  NOR4_X1 U8367 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6762) );
  NOR4_X1 U8368 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6761) );
  NOR4_X1 U8369 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6760) );
  NAND4_X1 U8370 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n6769)
         );
  NOR4_X1 U8371 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6767) );
  NOR4_X1 U8372 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6766) );
  NOR4_X1 U8373 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6765) );
  NOR4_X1 U8374 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6764) );
  NAND4_X1 U8375 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6768)
         );
  NOR2_X1 U8376 ( .A1(n6769), .A2(n6768), .ZN(n6770) );
  INV_X1 U8377 ( .A(n7300), .ZN(n7788) );
  NAND2_X1 U8378 ( .A1(n10033), .A2(n7788), .ZN(n7116) );
  AND3_X1 U8379 ( .A1(n7211), .A2(n7210), .A3(n7116), .ZN(n6771) );
  INV_X1 U8380 ( .A(n10073), .ZN(n10085) );
  INV_X1 U8381 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6774) );
  NOR2_X1 U8382 ( .A1(n10099), .A2(n6774), .ZN(n6775) );
  OAI21_X1 U8383 ( .B1(n6789), .B2(n10097), .A(n6776), .ZN(P2_U3488) );
  NAND2_X1 U8384 ( .A1(n7085), .A2(n7210), .ZN(n6777) );
  AND2_X1 U8385 ( .A1(n10073), .A2(n6792), .ZN(n6780) );
  NAND2_X1 U8386 ( .A1(n7788), .A2(n6778), .ZN(n7084) );
  OR2_X1 U8387 ( .A1(n7084), .A2(n6779), .ZN(n7104) );
  NAND2_X1 U8388 ( .A1(n6780), .A2(n7104), .ZN(n7080) );
  INV_X1 U8389 ( .A(n6781), .ZN(n7301) );
  NAND2_X1 U8390 ( .A1(n7080), .A2(n8915), .ZN(n7100) );
  NAND2_X1 U8391 ( .A1(n7111), .A2(n7100), .ZN(n6784) );
  INV_X1 U8392 ( .A(n7217), .ZN(n7110) );
  INV_X1 U8393 ( .A(n7104), .ZN(n7079) );
  NAND2_X1 U8394 ( .A1(n7210), .A2(n6880), .ZN(n6782) );
  OAI21_X1 U8395 ( .B1(n7110), .B2(n7079), .A(n7115), .ZN(n6783) );
  NOR2_X1 U8396 ( .A1(n10086), .A2(n6786), .ZN(n6787) );
  OAI21_X1 U8397 ( .B1(n6789), .B2(n10087), .A(n6788), .ZN(P2_U3456) );
  INV_X1 U8398 ( .A(n6790), .ZN(n6791) );
  NAND2_X1 U8399 ( .A1(n6821), .A2(n6792), .ZN(n6794) );
  NAND2_X1 U8400 ( .A1(n6794), .A2(n6793), .ZN(n6810) );
  NAND2_X1 U8401 ( .A1(n6810), .A2(n6795), .ZN(n6796) );
  NAND2_X1 U8402 ( .A1(n6796), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  MUX2_X1 U8403 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8699), .Z(n7343) );
  XNOR2_X1 U8404 ( .A(n7343), .B(n7342), .ZN(n6808) );
  MUX2_X1 U8405 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8699), .Z(n6805) );
  MUX2_X1 U8406 ( .A(n7446), .B(n6798), .S(n8699), .Z(n6803) );
  INV_X1 U8407 ( .A(n6803), .ZN(n6804) );
  MUX2_X1 U8408 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8699), .Z(n6802) );
  INV_X1 U8409 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6799) );
  MUX2_X1 U8410 ( .A(n7305), .B(n6799), .S(n8699), .Z(n6800) );
  INV_X1 U8411 ( .A(n6800), .ZN(n6801) );
  XNOR2_X1 U8412 ( .A(n6800), .B(n9998), .ZN(n9990) );
  INV_X1 U8413 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7172) );
  MUX2_X1 U8414 ( .A(n6313), .B(n7172), .S(n8699), .Z(n6971) );
  NAND2_X1 U8415 ( .A1(n6971), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9989) );
  XNOR2_X1 U8416 ( .A(n6802), .B(n6998), .ZN(n6982) );
  XNOR2_X1 U8417 ( .A(n6803), .B(n7015), .ZN(n7001) );
  NAND2_X1 U8418 ( .A1(n7002), .A2(n7001), .ZN(n7000) );
  OAI21_X1 U8419 ( .B1(n6804), .B2(n7015), .A(n7000), .ZN(n7191) );
  XNOR2_X1 U8420 ( .A(n6805), .B(n7178), .ZN(n7192) );
  AOI211_X1 U8421 ( .C1(n6808), .C2(n6807), .A(n8707), .B(n7341), .ZN(n6841)
         );
  NOR2_X1 U8422 ( .A1(n8699), .A2(P2_U3151), .ZN(n9114) );
  AND2_X1 U8423 ( .A1(n6810), .A2(n9114), .ZN(n6809) );
  MUX2_X1 U8424 ( .A(P2_U3893), .B(n6809), .S(n4516), .Z(n10014) );
  NOR2_X1 U8425 ( .A1(n8679), .A2(n7342), .ZN(n6840) );
  NOR2_X1 U8426 ( .A1(n4516), .A2(P2_U3151), .ZN(n9111) );
  MUX2_X1 U8427 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6301), .S(n6998), .Z(n6986)
         );
  AND2_X1 U8428 ( .A1(n6825), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6812) );
  NAND2_X1 U8429 ( .A1(n6811), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6813) );
  NAND2_X1 U8430 ( .A1(n9993), .A2(n6813), .ZN(n6985) );
  NAND2_X1 U8431 ( .A1(n6986), .A2(n6985), .ZN(n6984) );
  NAND2_X1 U8432 ( .A1(n6998), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6814) );
  MUX2_X1 U8433 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6326), .S(n7178), .Z(n7185)
         );
  AOI21_X1 U8434 ( .B1(n6280), .B2(n6817), .A(n7361), .ZN(n6819) );
  NOR2_X1 U8435 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6087), .ZN(n7525) );
  INV_X1 U8436 ( .A(n7525), .ZN(n6818) );
  OAI21_X1 U8437 ( .B1(n10022), .B2(n6819), .A(n6818), .ZN(n6839) );
  NOR2_X1 U8438 ( .A1(n6821), .A2(n6820), .ZN(n6822) );
  INV_X1 U8439 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6837) );
  INV_X1 U8440 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6824) );
  MUX2_X1 U8441 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6824), .S(n6823), .Z(n6989)
         );
  AND2_X1 U8442 ( .A1(n6825), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6826) );
  NAND2_X1 U8443 ( .A1(n6811), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U8444 ( .A1(n10005), .A2(n6827), .ZN(n6988) );
  NAND2_X1 U8445 ( .A1(n6989), .A2(n6988), .ZN(n6987) );
  NAND2_X1 U8446 ( .A1(n6998), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U8447 ( .A1(n6987), .A2(n6828), .ZN(n6829) );
  INV_X1 U8448 ( .A(n6830), .ZN(n6831) );
  INV_X1 U8449 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6832) );
  MUX2_X1 U8450 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6832), .S(n7178), .Z(n7181)
         );
  XNOR2_X1 U8451 ( .A(n7346), .B(n7342), .ZN(n6834) );
  NOR2_X1 U8452 ( .A1(n7732), .A2(n6834), .ZN(n7349) );
  AOI21_X1 U8453 ( .B1(n7732), .B2(n6834), .A(n7349), .ZN(n6836) );
  INV_X1 U8454 ( .A(n6835), .ZN(n6970) );
  OAI22_X1 U8455 ( .A1(n10011), .A2(n6837), .B1(n6836), .B2(n10026), .ZN(n6838) );
  OR4_X1 U8456 ( .A1(n6841), .A2(n6840), .A3(n6839), .A4(n6838), .ZN(P2_U3187)
         );
  NOR2_X1 U8457 ( .A1(n6847), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9871) );
  INV_X2 U8458 ( .A(n9871), .ZN(n9882) );
  AND2_X1 U8459 ( .A1(n6847), .A2(P1_U3086), .ZN(n7924) );
  INV_X2 U8460 ( .A(n7924), .ZN(n9884) );
  OAI222_X1 U8461 ( .A1(n9882), .A2(n6842), .B1(n9884), .B2(n6853), .C1(
        P1_U3086), .C2(n6911), .ZN(P1_U3354) );
  INV_X1 U8462 ( .A(n9327), .ZN(n6843) );
  OAI222_X1 U8463 ( .A1(n9882), .A2(n6844), .B1(n9884), .B2(n6854), .C1(
        P1_U3086), .C2(n6843), .ZN(P1_U3352) );
  INV_X1 U8464 ( .A(n7070), .ZN(n7066) );
  OAI222_X1 U8465 ( .A1(n9882), .A2(n6845), .B1(n9884), .B2(n6856), .C1(
        P1_U3086), .C2(n7066), .ZN(P1_U3353) );
  INV_X1 U8466 ( .A(n7051), .ZN(n7061) );
  OAI222_X1 U8467 ( .A1(n9882), .A2(n5204), .B1(P1_U3086), .B2(n7061), .C1(
        n6858), .C2(n9884), .ZN(P1_U3351) );
  OAI222_X1 U8468 ( .A1(P1_U3086), .A2(n9335), .B1(n9884), .B2(n6849), .C1(
        n6846), .C2(n9882), .ZN(P1_U3350) );
  NOR2_X1 U8469 ( .A1(n6847), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9109) );
  INV_X2 U8470 ( .A(n9109), .ZN(n9117) );
  NAND2_X1 U8471 ( .A1(n6847), .A2(P2_U3151), .ZN(n9122) );
  INV_X1 U8472 ( .A(n9122), .ZN(n9115) );
  OAI222_X1 U8473 ( .A1(n9117), .A2(n6849), .B1(n7342), .B2(P2_U3151), .C1(
        n6848), .C2(n9105), .ZN(P2_U3290) );
  OAI222_X1 U8474 ( .A1(n9117), .A2(n6852), .B1(n7700), .B2(P2_U3151), .C1(
        n6850), .C2(n9105), .ZN(P2_U3289) );
  INV_X1 U8475 ( .A(n6920), .ZN(n9348) );
  OAI222_X1 U8476 ( .A1(P1_U3086), .A2(n9348), .B1(n9884), .B2(n6852), .C1(
        n6851), .C2(n9882), .ZN(P1_U3349) );
  OAI222_X1 U8477 ( .A1(n9105), .A2(n5186), .B1(n9998), .B2(P2_U3151), .C1(
        n9117), .C2(n6853), .ZN(P2_U3294) );
  OAI222_X1 U8478 ( .A1(n9105), .A2(n6855), .B1(n7015), .B2(P2_U3151), .C1(
        n9117), .C2(n6854), .ZN(P2_U3292) );
  OAI222_X1 U8479 ( .A1(n9105), .A2(n6857), .B1(n6998), .B2(P2_U3151), .C1(
        n9117), .C2(n6856), .ZN(P2_U3293) );
  OAI222_X1 U8480 ( .A1(n9122), .A2(n5206), .B1(n7178), .B2(P2_U3151), .C1(
        n9117), .C2(n6858), .ZN(P2_U3291) );
  OAI222_X1 U8481 ( .A1(n9117), .A2(n6860), .B1(n7711), .B2(P2_U3151), .C1(
        n6859), .C2(n9105), .ZN(P2_U3288) );
  INV_X1 U8482 ( .A(n9372), .ZN(n6861) );
  INV_X1 U8483 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10382) );
  OAI222_X1 U8484 ( .A1(P1_U3086), .A2(n6861), .B1(n9884), .B2(n6860), .C1(
        n10382), .C2(n9882), .ZN(P1_U3348) );
  INV_X1 U8485 ( .A(n6862), .ZN(n6867) );
  AOI22_X1 U8486 ( .A1(n6944), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9871), .ZN(n6863) );
  OAI21_X1 U8487 ( .B1(n6867), .B2(n9884), .A(n6863), .ZN(P1_U3347) );
  INV_X1 U8488 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10512) );
  NAND2_X1 U8489 ( .A1(n9955), .A2(n6865), .ZN(n6866) );
  OAI21_X1 U8490 ( .B1(n9955), .B2(n10512), .A(n6866), .ZN(P1_U3440) );
  INV_X1 U8491 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6868) );
  OAI222_X1 U8492 ( .A1(n9105), .A2(n6868), .B1(n9117), .B2(n6867), .C1(
        P2_U3151), .C2(n7822), .ZN(P2_U3287) );
  INV_X1 U8493 ( .A(n7239), .ZN(n6869) );
  OAI21_X1 U8494 ( .B1(n7240), .B2(n6869), .A(P1_STATE_REG_SCAN_IN), .ZN(n6907) );
  INV_X1 U8495 ( .A(n6907), .ZN(n6872) );
  NAND2_X1 U8496 ( .A1(n7136), .A2(n7239), .ZN(n6870) );
  NAND2_X1 U8497 ( .A1(n6871), .A2(n6870), .ZN(n6908) );
  AND2_X1 U8498 ( .A1(n6872), .A2(n6908), .ZN(n9933) );
  NOR2_X1 U8499 ( .A1(n9933), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8500 ( .A(n6873), .ZN(n6876) );
  INV_X1 U8501 ( .A(n7873), .ZN(n7814) );
  INV_X1 U8502 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6874) );
  OAI222_X1 U8503 ( .A1(n9117), .A2(n6876), .B1(n7814), .B2(P2_U3151), .C1(
        n6874), .C2(n9122), .ZN(P2_U3286) );
  INV_X1 U8504 ( .A(n6950), .ZN(n6960) );
  INV_X1 U8505 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6875) );
  OAI222_X1 U8506 ( .A1(P1_U3086), .A2(n6960), .B1(n9884), .B2(n6876), .C1(
        n6875), .C2(n9882), .ZN(P1_U3346) );
  INV_X1 U8507 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6877) );
  OAI222_X1 U8508 ( .A1(n9117), .A2(n6879), .B1(n8072), .B2(P2_U3151), .C1(
        n6877), .C2(n9105), .ZN(P2_U3285) );
  INV_X1 U8509 ( .A(n6957), .ZN(n9379) );
  INV_X1 U8510 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6878) );
  OAI222_X1 U8511 ( .A1(P1_U3086), .A2(n9379), .B1(n9884), .B2(n6879), .C1(
        n6878), .C2(n9882), .ZN(P1_U3345) );
  INV_X1 U8512 ( .A(n6881), .ZN(n6882) );
  AOI22_X1 U8513 ( .A1(n6883), .A2(n5076), .B1(n7109), .B2(n6882), .ZN(
        P2_U3376) );
  AND2_X1 U8514 ( .A1(n6883), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8515 ( .A1(n6883), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8516 ( .A1(n6883), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8517 ( .A1(n6883), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8518 ( .A1(n6883), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8519 ( .A1(n6883), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8520 ( .A1(n6883), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8521 ( .A1(n6883), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8522 ( .A1(n6883), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8523 ( .A1(n6883), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8524 ( .A1(n6883), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8525 ( .A1(n6883), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8526 ( .A1(n6883), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8527 ( .A1(n6883), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8528 ( .A1(n6883), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8529 ( .A1(n6883), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8530 ( .A1(n6883), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8531 ( .A1(n6883), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8532 ( .A1(n6883), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8533 ( .A1(n6883), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8534 ( .A1(n6883), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8535 ( .A1(n6883), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8536 ( .A1(n6883), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8537 ( .A1(n6883), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8538 ( .A1(n6883), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8539 ( .A1(n6883), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8540 ( .A1(n6883), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8541 ( .A1(n6883), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8542 ( .A1(n6883), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8543 ( .A1(n6883), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8544 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6885) );
  INV_X1 U8545 ( .A(n6884), .ZN(n6886) );
  INV_X1 U8546 ( .A(n8097), .ZN(n8062) );
  OAI222_X1 U8547 ( .A1(n9105), .A2(n6885), .B1(n9117), .B2(n6886), .C1(
        P2_U3151), .C2(n8062), .ZN(P2_U3284) );
  INV_X1 U8548 ( .A(n6955), .ZN(n9391) );
  INV_X1 U8549 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10367) );
  OAI222_X1 U8550 ( .A1(n9391), .A2(P1_U3086), .B1(n9884), .B2(n6886), .C1(
        n10367), .C2(n9882), .ZN(P1_U3344) );
  INV_X1 U8551 ( .A(n6944), .ZN(n6903) );
  INV_X1 U8552 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6887) );
  MUX2_X1 U8553 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6887), .S(n7070), .Z(n6890)
         );
  INV_X1 U8554 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6888) );
  MUX2_X1 U8555 ( .A(n6888), .B(P1_REG1_REG_1__SCAN_IN), .S(n6911), .Z(n9311)
         );
  AND2_X1 U8556 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9312) );
  NAND2_X1 U8557 ( .A1(n9311), .A2(n9312), .ZN(n9310) );
  NAND2_X1 U8558 ( .A1(n9309), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7071) );
  NAND2_X1 U8559 ( .A1(n9310), .A2(n7071), .ZN(n6889) );
  NAND2_X1 U8560 ( .A1(n6890), .A2(n6889), .ZN(n9324) );
  NAND2_X1 U8561 ( .A1(n7070), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U8562 ( .A1(n9324), .A2(n9322), .ZN(n6893) );
  INV_X1 U8563 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6891) );
  MUX2_X1 U8564 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6891), .S(n9327), .Z(n6892)
         );
  NAND2_X1 U8565 ( .A1(n6893), .A2(n6892), .ZN(n9326) );
  NAND2_X1 U8566 ( .A1(n9327), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7053) );
  NAND2_X1 U8567 ( .A1(n9326), .A2(n7053), .ZN(n6896) );
  INV_X1 U8568 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6894) );
  MUX2_X1 U8569 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6894), .S(n7051), .Z(n6895)
         );
  NAND2_X1 U8570 ( .A1(n6896), .A2(n6895), .ZN(n9343) );
  NAND2_X1 U8571 ( .A1(n7051), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9342) );
  MUX2_X1 U8572 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5374), .S(n9335), .Z(n9341)
         );
  AOI21_X1 U8573 ( .B1(n9343), .B2(n9342), .A(n9341), .ZN(n6897) );
  INV_X1 U8574 ( .A(n6897), .ZN(n9356) );
  INV_X1 U8575 ( .A(n9335), .ZN(n6898) );
  NAND2_X1 U8576 ( .A1(n6898), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9355) );
  INV_X1 U8577 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7493) );
  MUX2_X1 U8578 ( .A(n7493), .B(P1_REG1_REG_6__SCAN_IN), .S(n6920), .Z(n9354)
         );
  AOI21_X1 U8579 ( .B1(n9356), .B2(n9355), .A(n9354), .ZN(n9370) );
  NOR2_X1 U8580 ( .A1(n9348), .A2(n7493), .ZN(n9365) );
  INV_X1 U8581 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6899) );
  MUX2_X1 U8582 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6899), .S(n9372), .Z(n6900)
         );
  OAI21_X1 U8583 ( .B1(n9370), .B2(n9365), .A(n6900), .ZN(n9368) );
  NAND2_X1 U8584 ( .A1(n9372), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6935) );
  MUX2_X1 U8585 ( .A(n6936), .B(P1_REG1_REG_8__SCAN_IN), .S(n6944), .Z(n6901)
         );
  AOI21_X1 U8586 ( .B1(n9368), .B2(n6935), .A(n6901), .ZN(n6941) );
  INV_X1 U8587 ( .A(n6941), .ZN(n6902) );
  OAI21_X1 U8588 ( .B1(n6936), .B2(n6903), .A(n6902), .ZN(n6906) );
  MUX2_X1 U8589 ( .A(n6904), .B(P1_REG1_REG_9__SCAN_IN), .S(n6950), .Z(n6905)
         );
  NOR2_X1 U8590 ( .A1(n6905), .A2(n6906), .ZN(n6959) );
  AOI21_X1 U8591 ( .B1(n6906), .B2(n6905), .A(n6959), .ZN(n6931) );
  NAND2_X1 U8592 ( .A1(n6926), .A2(n9927), .ZN(n9464) );
  NAND2_X1 U8593 ( .A1(n6926), .A2(n6909), .ZN(n9465) );
  INV_X1 U8594 ( .A(n9465), .ZN(n9445) );
  AOI22_X1 U8595 ( .A1(n6950), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7644), .B2(
        n6960), .ZN(n6925) );
  INV_X1 U8596 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6910) );
  XNOR2_X1 U8597 ( .A(n7070), .B(n6910), .ZN(n7069) );
  XNOR2_X1 U8598 ( .A(n6911), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9315) );
  AND2_X1 U8599 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9314) );
  NAND2_X1 U8600 ( .A1(n9315), .A2(n9314), .ZN(n9313) );
  NAND2_X1 U8601 ( .A1(n9309), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8602 ( .A1(n9313), .A2(n6912), .ZN(n7068) );
  NAND2_X1 U8603 ( .A1(n7069), .A2(n7068), .ZN(n7067) );
  NAND2_X1 U8604 ( .A1(n7070), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6913) );
  NAND2_X1 U8605 ( .A1(n7067), .A2(n6913), .ZN(n9320) );
  INV_X1 U8606 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6914) );
  XNOR2_X1 U8607 ( .A(n9327), .B(n6914), .ZN(n9321) );
  NAND2_X1 U8608 ( .A1(n9320), .A2(n9321), .ZN(n9319) );
  NAND2_X1 U8609 ( .A1(n9327), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U8610 ( .A1(n9319), .A2(n6915), .ZN(n7059) );
  INV_X1 U8611 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6916) );
  XNOR2_X1 U8612 ( .A(n7051), .B(n6916), .ZN(n7058) );
  NAND2_X1 U8613 ( .A1(n7059), .A2(n7058), .ZN(n7057) );
  NAND2_X1 U8614 ( .A1(n7051), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U8615 ( .A1(n7057), .A2(n6917), .ZN(n9339) );
  INV_X1 U8616 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7479) );
  MUX2_X1 U8617 ( .A(n7479), .B(P1_REG2_REG_5__SCAN_IN), .S(n9335), .Z(n9340)
         );
  NAND2_X1 U8618 ( .A1(n9339), .A2(n9340), .ZN(n9338) );
  OR2_X1 U8619 ( .A1(n9335), .A2(n7479), .ZN(n6918) );
  NAND2_X1 U8620 ( .A1(n9338), .A2(n6918), .ZN(n9352) );
  INV_X1 U8621 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6919) );
  MUX2_X1 U8622 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6919), .S(n6920), .Z(n9353)
         );
  NAND2_X1 U8623 ( .A1(n9352), .A2(n9353), .ZN(n9351) );
  NAND2_X1 U8624 ( .A1(n6920), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U8625 ( .A1(n9351), .A2(n6921), .ZN(n9363) );
  INV_X1 U8626 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6922) );
  MUX2_X1 U8627 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6922), .S(n9372), .Z(n9364)
         );
  NAND2_X1 U8628 ( .A1(n9363), .A2(n9364), .ZN(n9362) );
  NAND2_X1 U8629 ( .A1(n9372), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8630 ( .A1(n9362), .A2(n6923), .ZN(n6932) );
  MUX2_X1 U8631 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7662), .S(n6944), .Z(n6933)
         );
  AND2_X1 U8632 ( .A1(n6932), .A2(n6933), .ZN(n6947) );
  AOI21_X1 U8633 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6944), .A(n6947), .ZN(
        n6924) );
  NAND2_X1 U8634 ( .A1(n6925), .A2(n6924), .ZN(n6949) );
  OAI21_X1 U8635 ( .B1(n6925), .B2(n6924), .A(n6949), .ZN(n6929) );
  AND2_X1 U8636 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8001) );
  AOI21_X1 U8637 ( .B1(n9933), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n8001), .ZN(
        n6927) );
  OAI21_X1 U8638 ( .B1(n9459), .B2(n6960), .A(n6927), .ZN(n6928) );
  AOI21_X1 U8639 ( .B1(n9445), .B2(n6929), .A(n6928), .ZN(n6930) );
  OAI21_X1 U8640 ( .B1(n6931), .B2(n9464), .A(n6930), .ZN(P1_U3252) );
  OAI21_X1 U8641 ( .B1(n6933), .B2(n6932), .A(n9445), .ZN(n6946) );
  INV_X1 U8642 ( .A(n9459), .ZN(n9373) );
  INV_X1 U8643 ( .A(n9933), .ZN(n9472) );
  INV_X1 U8644 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U8645 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9910) );
  OAI21_X1 U8646 ( .B1(n9472), .B2(n6934), .A(n9910), .ZN(n6943) );
  INV_X1 U8647 ( .A(n9368), .ZN(n6939) );
  INV_X1 U8648 ( .A(n6935), .ZN(n6938) );
  MUX2_X1 U8649 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6936), .S(n6944), .Z(n6937)
         );
  NOR3_X1 U8650 ( .A1(n6939), .A2(n6938), .A3(n6937), .ZN(n6940) );
  NOR3_X1 U8651 ( .A1(n9464), .A2(n6941), .A3(n6940), .ZN(n6942) );
  AOI211_X1 U8652 ( .C1(n9373), .C2(n6944), .A(n6943), .B(n6942), .ZN(n6945)
         );
  OAI21_X1 U8653 ( .B1(n6947), .B2(n6946), .A(n6945), .ZN(P1_U3251) );
  INV_X1 U8654 ( .A(n7323), .ZN(n7332) );
  NOR2_X1 U8655 ( .A1(n7323), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6948) );
  AOI21_X1 U8656 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7323), .A(n6948), .ZN(
        n6953) );
  AOI22_X1 U8657 ( .A1(n6957), .A2(n7780), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n9379), .ZN(n9382) );
  OAI21_X1 U8658 ( .B1(n6950), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6949), .ZN(
        n9383) );
  NOR2_X1 U8659 ( .A1(n9382), .A2(n9383), .ZN(n9381) );
  AOI21_X1 U8660 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6957), .A(n9381), .ZN(
        n9399) );
  NAND2_X1 U8661 ( .A1(n6955), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6951) );
  OAI21_X1 U8662 ( .B1(n6955), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6951), .ZN(
        n9398) );
  NOR2_X1 U8663 ( .A1(n9399), .A2(n9398), .ZN(n9397) );
  AOI21_X1 U8664 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6955), .A(n9397), .ZN(
        n6952) );
  NAND2_X1 U8665 ( .A1(n6953), .A2(n6952), .ZN(n7322) );
  OAI21_X1 U8666 ( .B1(n6953), .B2(n6952), .A(n7322), .ZN(n6965) );
  INV_X1 U8667 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6954) );
  MUX2_X1 U8668 ( .A(n6954), .B(P1_REG1_REG_12__SCAN_IN), .S(n7323), .Z(n6962)
         );
  INV_X1 U8669 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6956) );
  MUX2_X1 U8670 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6956), .S(n6955), .Z(n9395)
         );
  MUX2_X1 U8671 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6958), .S(n6957), .Z(n9386)
         );
  AOI21_X1 U8672 ( .B1(n6960), .B2(n6904), .A(n6959), .ZN(n9387) );
  NAND2_X1 U8673 ( .A1(n9386), .A2(n9387), .ZN(n9385) );
  OAI21_X1 U8674 ( .B1(n9379), .B2(n6958), .A(n9385), .ZN(n9396) );
  NAND2_X1 U8675 ( .A1(n9395), .A2(n9396), .ZN(n9394) );
  OAI21_X1 U8676 ( .B1(n9391), .B2(n6956), .A(n9394), .ZN(n6961) );
  NOR2_X1 U8677 ( .A1(n6961), .A2(n6962), .ZN(n7331) );
  AOI21_X1 U8678 ( .B1(n6962), .B2(n6961), .A(n7331), .ZN(n6963) );
  NOR2_X1 U8679 ( .A1(n9464), .A2(n6963), .ZN(n6964) );
  AOI21_X1 U8680 ( .B1(n9445), .B2(n6965), .A(n6964), .ZN(n6967) );
  AND2_X1 U8681 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9182) );
  AOI21_X1 U8682 ( .B1(n9933), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9182), .ZN(
        n6966) );
  OAI211_X1 U8683 ( .C1(n7332), .C2(n9459), .A(n6967), .B(n6966), .ZN(P1_U3255) );
  INV_X1 U8684 ( .A(n6968), .ZN(n6978) );
  INV_X1 U8685 ( .A(n8080), .ZN(n8570) );
  INV_X1 U8686 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6969) );
  OAI222_X1 U8687 ( .A1(n9117), .A2(n6978), .B1(n8570), .B2(P2_U3151), .C1(
        n6969), .C2(n9105), .ZN(P2_U3283) );
  INV_X1 U8688 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6976) );
  NAND2_X1 U8689 ( .A1(n6970), .A2(n8707), .ZN(n6973) );
  OAI21_X1 U8690 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6971), .A(n9989), .ZN(n6972) );
  AOI22_X1 U8691 ( .A1(n6973), .A2(n6972), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6975) );
  NAND2_X1 U8692 ( .A1(n10014), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6974) );
  OAI211_X1 U8693 ( .C1(n10011), .C2(n6976), .A(n6975), .B(n6974), .ZN(
        P2_U3182) );
  AOI22_X1 U8694 ( .A1(n8599), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n9115), .ZN(n6977) );
  OAI21_X1 U8695 ( .B1(n6979), .B2(n9117), .A(n6977), .ZN(P2_U3282) );
  INV_X1 U8696 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10511) );
  OAI222_X1 U8697 ( .A1(P1_U3086), .A2(n7332), .B1(n9884), .B2(n6978), .C1(
        n10511), .C2(n9882), .ZN(P1_U3343) );
  INV_X1 U8698 ( .A(n7330), .ZN(n9404) );
  INV_X1 U8699 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10385) );
  OAI222_X1 U8700 ( .A1(P1_U3086), .A2(n9404), .B1(n9884), .B2(n6979), .C1(
        n10385), .C2(n9882), .ZN(P1_U3342) );
  AOI211_X1 U8701 ( .C1(n6982), .C2(n6981), .A(n8707), .B(n6980), .ZN(n6983)
         );
  INV_X1 U8702 ( .A(n6983), .ZN(n6997) );
  OAI21_X1 U8703 ( .B1(n6986), .B2(n6985), .A(n6984), .ZN(n6995) );
  OAI21_X1 U8704 ( .B1(n6989), .B2(n6988), .A(n6987), .ZN(n6990) );
  INV_X1 U8705 ( .A(n6990), .ZN(n6991) );
  OAI22_X1 U8706 ( .A1(n10026), .A2(n6991), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6302), .ZN(n6994) );
  INV_X1 U8707 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6992) );
  NOR2_X1 U8708 ( .A1(n10011), .A2(n6992), .ZN(n6993) );
  AOI211_X1 U8709 ( .C1(n9997), .C2(n6995), .A(n6994), .B(n6993), .ZN(n6996)
         );
  OAI211_X1 U8710 ( .C1(n8679), .C2(n6998), .A(n6997), .B(n6996), .ZN(P2_U3184) );
  NAND2_X1 U8711 ( .A1(n9306), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6999) );
  OAI21_X1 U8712 ( .B1(n9570), .B2(n9306), .A(n6999), .ZN(P1_U3579) );
  OAI21_X1 U8713 ( .B1(n7002), .B2(n7001), .A(n7000), .ZN(n7003) );
  NAND2_X1 U8714 ( .A1(n7003), .A2(n10020), .ZN(n7014) );
  AOI21_X1 U8715 ( .B1(n7005), .B2(n7446), .A(n7004), .ZN(n7007) );
  INV_X1 U8716 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7447) );
  NOR2_X1 U8717 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7447), .ZN(n7293) );
  INV_X1 U8718 ( .A(n7293), .ZN(n7006) );
  OAI21_X1 U8719 ( .B1(n10026), .B2(n7007), .A(n7006), .ZN(n7012) );
  AOI21_X1 U8720 ( .B1(n7009), .B2(n6798), .A(n7008), .ZN(n7010) );
  NOR2_X1 U8721 ( .A1(n10022), .A2(n7010), .ZN(n7011) );
  AOI211_X1 U8722 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n10018), .A(n7012), .B(
        n7011), .ZN(n7013) );
  OAI211_X1 U8723 ( .C1(n8679), .C2(n7015), .A(n7014), .B(n7013), .ZN(P2_U3185) );
  INV_X1 U8724 ( .A(n7327), .ZN(n9417) );
  INV_X1 U8725 ( .A(n7016), .ZN(n7018) );
  INV_X1 U8726 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7017) );
  OAI222_X1 U8727 ( .A1(n9417), .A2(P1_U3086), .B1(n9884), .B2(n7018), .C1(
        n7017), .C2(n9882), .ZN(P1_U3341) );
  INV_X1 U8728 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7019) );
  OAI222_X1 U8729 ( .A1(n9105), .A2(n7019), .B1(n9117), .B2(n7018), .C1(
        P2_U3151), .C2(n8619), .ZN(P2_U3281) );
  OAI21_X1 U8730 ( .B1(n7022), .B2(n7021), .A(n7020), .ZN(n9939) );
  INV_X1 U8731 ( .A(n9939), .ZN(n9947) );
  XNOR2_X1 U8732 ( .A(n7024), .B(n7023), .ZN(n7027) );
  NAND2_X1 U8733 ( .A1(n9305), .A2(n9728), .ZN(n7026) );
  NAND2_X1 U8734 ( .A1(n7038), .A2(n9727), .ZN(n7025) );
  NAND2_X1 U8735 ( .A1(n7026), .A2(n7025), .ZN(n7148) );
  AOI21_X1 U8736 ( .B1(n7027), .B2(n9724), .A(n7148), .ZN(n9937) );
  OAI211_X1 U8737 ( .C1(n9888), .C2(n9944), .A(n9813), .B(n7153), .ZN(n9941)
         );
  OAI211_X1 U8738 ( .C1(n9804), .C2(n9947), .A(n9937), .B(n9941), .ZN(n7374)
         );
  OAI22_X1 U8739 ( .A1(n9823), .A2(n9944), .B1(n9988), .B2(n6888), .ZN(n7031)
         );
  AOI21_X1 U8740 ( .B1(n7374), .B2(n9988), .A(n7031), .ZN(n7032) );
  INV_X1 U8741 ( .A(n7032), .ZN(P1_U3523) );
  NAND2_X1 U8742 ( .A1(n7038), .A2(n9149), .ZN(n7037) );
  INV_X1 U8743 ( .A(n7039), .ZN(n7034) );
  INV_X1 U8744 ( .A(n7240), .ZN(n7035) );
  AOI22_X1 U8745 ( .A1(n7041), .A2(n8231), .B1(n7035), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n7036) );
  NAND2_X1 U8746 ( .A1(n7037), .A2(n7036), .ZN(n7046) );
  NAND2_X1 U8747 ( .A1(n7038), .A2(n8231), .ZN(n7043) );
  NAND2_X1 U8748 ( .A1(n7041), .A2(n8233), .ZN(n7042) );
  INV_X1 U8749 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U8750 ( .A1(n4511), .A2(n5144), .ZN(n7044) );
  INV_X1 U8751 ( .A(n7134), .ZN(n7045) );
  OAI21_X1 U8752 ( .B1(n7046), .B2(n7044), .A(n7045), .ZN(n9887) );
  MUX2_X1 U8753 ( .A(n9887), .B(n9314), .S(n7047), .Z(n7050) );
  NOR2_X1 U8754 ( .A1(n9927), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7048) );
  NOR2_X1 U8755 ( .A1(n5966), .A2(n7048), .ZN(n9928) );
  NOR2_X1 U8756 ( .A1(n9928), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9925) );
  AOI211_X1 U8757 ( .C1(n7050), .C2(n7049), .A(n9925), .B(n9306), .ZN(n7078)
         );
  MUX2_X1 U8758 ( .A(n6894), .B(P1_REG1_REG_4__SCAN_IN), .S(n7051), .Z(n7052)
         );
  NAND3_X1 U8759 ( .A1(n9326), .A2(n7053), .A3(n7052), .ZN(n7054) );
  NAND2_X1 U8760 ( .A1(n9343), .A2(n7054), .ZN(n7056) );
  NAND2_X1 U8761 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n7278) );
  NAND2_X1 U8762 ( .A1(n9933), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n7055) );
  OAI211_X1 U8763 ( .C1(n9464), .C2(n7056), .A(n7278), .B(n7055), .ZN(n7063)
         );
  OAI21_X1 U8764 ( .B1(n7059), .B2(n7058), .A(n7057), .ZN(n7060) );
  OAI22_X1 U8765 ( .A1(n7061), .A2(n9459), .B1(n9465), .B2(n7060), .ZN(n7062)
         );
  OR3_X1 U8766 ( .A1(n7078), .A2(n7063), .A3(n7062), .ZN(P1_U3247) );
  INV_X1 U8767 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7509) );
  NOR2_X1 U8768 ( .A1(n7509), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7064) );
  AOI21_X1 U8769 ( .B1(n9933), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n7064), .ZN(
        n7065) );
  OAI21_X1 U8770 ( .B1(n9459), .B2(n7066), .A(n7065), .ZN(n7077) );
  OAI21_X1 U8771 ( .B1(n7069), .B2(n7068), .A(n7067), .ZN(n7075) );
  MUX2_X1 U8772 ( .A(n6887), .B(P1_REG1_REG_2__SCAN_IN), .S(n7070), .Z(n7072)
         );
  NAND3_X1 U8773 ( .A1(n7072), .A2(n9310), .A3(n7071), .ZN(n7073) );
  NAND2_X1 U8774 ( .A1(n9324), .A2(n7073), .ZN(n7074) );
  OAI22_X1 U8775 ( .A1(n9465), .A2(n7075), .B1(n9464), .B2(n7074), .ZN(n7076)
         );
  OR3_X1 U8776 ( .A1(n7078), .A2(n7077), .A3(n7076), .ZN(P1_U3245) );
  NAND2_X1 U8777 ( .A1(n7111), .A2(n7079), .ZN(n7083) );
  INV_X1 U8778 ( .A(n7080), .ZN(n7081) );
  NAND2_X1 U8779 ( .A1(n7115), .A2(n7081), .ZN(n7082) );
  NAND2_X1 U8780 ( .A1(n7300), .A2(n7652), .ZN(n7087) );
  AND2_X1 U8781 ( .A1(n7087), .A2(n7086), .ZN(n7088) );
  INV_X1 U8782 ( .A(n8198), .ZN(n7199) );
  NAND2_X1 U8783 ( .A1(n7199), .A2(n7167), .ZN(n7090) );
  AND2_X1 U8784 ( .A1(n7091), .A2(n7090), .ZN(n7097) );
  XNOR2_X1 U8785 ( .A(n7306), .B(n8198), .ZN(n7093) );
  INV_X1 U8786 ( .A(n7093), .ZN(n7092) );
  INV_X1 U8787 ( .A(n7097), .ZN(n7094) );
  INV_X1 U8788 ( .A(n7202), .ZN(n7095) );
  AOI21_X1 U8789 ( .B1(n7097), .B2(n7096), .A(n7095), .ZN(n7121) );
  INV_X1 U8790 ( .A(n7210), .ZN(n7099) );
  AOI21_X1 U8791 ( .B1(n7099), .B2(n7100), .A(n7098), .ZN(n7103) );
  NAND2_X1 U8792 ( .A1(n7101), .A2(n7100), .ZN(n7102) );
  OAI211_X1 U8793 ( .C1(n7105), .C2(n7104), .A(n7103), .B(n7102), .ZN(n7108)
         );
  INV_X1 U8794 ( .A(n7105), .ZN(n7107) );
  AOI22_X1 U8795 ( .A1(n7108), .A2(P2_STATE_REG_SCAN_IN), .B1(n7107), .B2(
        n7106), .ZN(n7285) );
  NAND2_X1 U8796 ( .A1(n7285), .A2(n7109), .ZN(n8341) );
  INV_X1 U8797 ( .A(n8564), .ZN(n7287) );
  AND2_X1 U8798 ( .A1(n7111), .A2(n7110), .ZN(n7114) );
  INV_X1 U8799 ( .A(n7114), .ZN(n7112) );
  OR2_X2 U8800 ( .A1(n7112), .A2(n7113), .ZN(n8544) );
  NAND2_X1 U8801 ( .A1(n7115), .A2(n10085), .ZN(n7117) );
  INV_X2 U8802 ( .A(n8551), .ZN(n8534) );
  AOI22_X1 U8803 ( .A1(n8548), .A2(n8566), .B1(n7306), .B2(n8534), .ZN(n7118)
         );
  OAI21_X1 U8804 ( .B1(n7287), .B2(n8544), .A(n7118), .ZN(n7119) );
  AOI21_X1 U8805 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8341), .A(n7119), .ZN(
        n7120) );
  OAI21_X1 U8806 ( .B1(n8538), .B2(n7121), .A(n7120), .ZN(P2_U3162) );
  INV_X1 U8807 ( .A(n7122), .ZN(n7124) );
  NOR2_X1 U8808 ( .A1(n7124), .A2(n7123), .ZN(n7389) );
  INV_X1 U8809 ( .A(n7125), .ZN(n9867) );
  NAND2_X1 U8810 ( .A1(n7389), .A2(n9867), .ZN(n7144) );
  INV_X1 U8811 ( .A(n7144), .ZN(n7126) );
  INV_X1 U8812 ( .A(n7147), .ZN(n7127) );
  OR2_X1 U8813 ( .A1(n7175), .A2(n5937), .ZN(n7394) );
  XNOR2_X1 U8814 ( .A(n7132), .B(n8277), .ZN(n7250) );
  INV_X2 U8815 ( .A(n8231), .ZN(n8284) );
  OAI22_X1 U8816 ( .A1(n9889), .A2(n8310), .B1(n9944), .B2(n8284), .ZN(n7247)
         );
  XNOR2_X1 U8817 ( .A(n7249), .B(n7247), .ZN(n7135) );
  XNOR2_X1 U8818 ( .A(n7250), .B(n7135), .ZN(n7138) );
  OR2_X1 U8819 ( .A1(n9956), .A2(n7136), .ZN(n7141) );
  INV_X1 U8820 ( .A(n7141), .ZN(n7137) );
  NAND2_X1 U8821 ( .A1(n7138), .A2(n9906), .ZN(n7150) );
  INV_X1 U8822 ( .A(n7139), .ZN(n7142) );
  NAND2_X1 U8823 ( .A1(n7140), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7631) );
  NAND3_X1 U8824 ( .A1(n7142), .A2(n7141), .A3(n7631), .ZN(n7143) );
  NAND2_X1 U8825 ( .A1(n7144), .A2(n7143), .ZN(n7242) );
  AND2_X1 U8826 ( .A1(n7242), .A2(n7145), .ZN(n9895) );
  INV_X1 U8827 ( .A(n9895), .ZN(n8335) );
  AOI22_X1 U8828 ( .A1(n8335), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9900), .B2(
        n7148), .ZN(n7149) );
  OAI211_X1 U8829 ( .C1(n9944), .C2(n9903), .A(n7150), .B(n7149), .ZN(P1_U3222) );
  OAI21_X1 U8830 ( .B1(n7152), .B2(n7154), .A(n7151), .ZN(n7514) );
  AOI211_X1 U8831 ( .C1(n7256), .C2(n7153), .A(n9969), .B(n7232), .ZN(n7512)
         );
  XNOR2_X1 U8832 ( .A(n7155), .B(n7154), .ZN(n7159) );
  NAND2_X1 U8833 ( .A1(n9304), .A2(n9728), .ZN(n7157) );
  NAND2_X1 U8834 ( .A1(n4512), .A2(n9727), .ZN(n7156) );
  NAND2_X1 U8835 ( .A1(n7157), .A2(n7156), .ZN(n8334) );
  INV_X1 U8836 ( .A(n8334), .ZN(n7158) );
  OAI21_X1 U8837 ( .B1(n7159), .B2(n9659), .A(n7158), .ZN(n7510) );
  AOI211_X1 U8838 ( .C1(n9979), .C2(n7514), .A(n7512), .B(n7510), .ZN(n7320)
         );
  OAI22_X1 U8839 ( .A1(n9823), .A2(n8338), .B1(n9988), .B2(n6887), .ZN(n7160)
         );
  INV_X1 U8840 ( .A(n7160), .ZN(n7161) );
  OAI21_X1 U8841 ( .B1(n7320), .B2(n9985), .A(n7161), .ZN(P1_U3524) );
  INV_X1 U8842 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7163) );
  INV_X1 U8843 ( .A(n7162), .ZN(n7164) );
  INV_X1 U8844 ( .A(n8641), .ZN(n8633) );
  OAI222_X1 U8845 ( .A1(n9122), .A2(n7163), .B1(n9117), .B2(n7164), .C1(
        P2_U3151), .C2(n8633), .ZN(P2_U3280) );
  INV_X1 U8846 ( .A(n7555), .ZN(n7560) );
  INV_X1 U8847 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10403) );
  OAI222_X1 U8848 ( .A1(n7560), .A2(P1_U3086), .B1(n9884), .B2(n7164), .C1(
        n10403), .C2(n9882), .ZN(P1_U3340) );
  INV_X1 U8849 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7169) );
  INV_X1 U8850 ( .A(n7165), .ZN(n8340) );
  OAI21_X1 U8851 ( .B1(n8914), .B2(n10078), .A(n8340), .ZN(n7166) );
  OR2_X1 U8852 ( .A1(n6678), .A2(n8928), .ZN(n7218) );
  OAI211_X1 U8853 ( .C1(n10073), .C2(n7167), .A(n7166), .B(n7218), .ZN(n7170)
         );
  NAND2_X1 U8854 ( .A1(n7170), .A2(n10086), .ZN(n7168) );
  OAI21_X1 U8855 ( .B1(n7169), .B2(n10086), .A(n7168), .ZN(P2_U3390) );
  NAND2_X1 U8856 ( .A1(n7170), .A2(n10099), .ZN(n7171) );
  OAI21_X1 U8857 ( .B1(n10099), .B2(n7172), .A(n7171), .ZN(P2_U3459) );
  INV_X1 U8858 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7177) );
  INV_X1 U8859 ( .A(n7454), .ZN(n7173) );
  OAI21_X1 U8860 ( .B1(n9979), .B2(n9724), .A(n7173), .ZN(n7174) );
  NAND2_X1 U8861 ( .A1(n4512), .A2(n9728), .ZN(n7452) );
  OAI211_X1 U8862 ( .C1(n7175), .C2(n9888), .A(n7174), .B(n7452), .ZN(n9824)
         );
  NAND2_X1 U8863 ( .A1(n9824), .A2(n9860), .ZN(n7176) );
  OAI21_X1 U8864 ( .B1(n9860), .B2(n7177), .A(n7176), .ZN(P1_U3453) );
  INV_X1 U8865 ( .A(n7178), .ZN(n7195) );
  INV_X1 U8866 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7189) );
  OAI21_X1 U8867 ( .B1(n7181), .B2(n7180), .A(n7179), .ZN(n7182) );
  INV_X1 U8868 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10486) );
  NOR2_X1 U8869 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10486), .ZN(n7434) );
  AOI21_X1 U8870 ( .B1(n8660), .B2(n7182), .A(n7434), .ZN(n7188) );
  OAI21_X1 U8871 ( .B1(n7185), .B2(n7184), .A(n7183), .ZN(n7186) );
  NAND2_X1 U8872 ( .A1(n9997), .A2(n7186), .ZN(n7187) );
  OAI211_X1 U8873 ( .C1(n7189), .C2(n10011), .A(n7188), .B(n7187), .ZN(n7194)
         );
  AOI211_X1 U8874 ( .C1(n7192), .C2(n7191), .A(n8707), .B(n7190), .ZN(n7193)
         );
  AOI211_X1 U8875 ( .C1(n10014), .C2(n7195), .A(n7194), .B(n7193), .ZN(n7196)
         );
  INV_X1 U8876 ( .A(n7196), .ZN(P2_U3186) );
  INV_X1 U8877 ( .A(n7197), .ZN(n7223) );
  INV_X1 U8878 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7198) );
  OAI222_X1 U8879 ( .A1(n9117), .A2(n7223), .B1(n8658), .B2(P2_U3151), .C1(
        n7198), .C2(n9122), .ZN(P2_U3279) );
  XNOR2_X1 U8880 ( .A(n8198), .B(n7200), .ZN(n7286) );
  XNOR2_X1 U8881 ( .A(n7286), .B(n7287), .ZN(n7204) );
  NAND2_X1 U8882 ( .A1(n7202), .A2(n7201), .ZN(n7203) );
  NAND2_X1 U8883 ( .A1(n7203), .A2(n7204), .ZN(n7290) );
  OAI21_X1 U8884 ( .B1(n7204), .B2(n7203), .A(n7290), .ZN(n7208) );
  AOI22_X1 U8885 ( .A1(n8548), .A2(n8565), .B1(n10032), .B2(n8534), .ZN(n7206)
         );
  NAND2_X1 U8886 ( .A1(n8341), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7205) );
  OAI211_X1 U8887 ( .C1(n8929), .C2(n8544), .A(n7206), .B(n7205), .ZN(n7207)
         );
  AOI21_X1 U8888 ( .B1(n8515), .B2(n7208), .A(n7207), .ZN(n7209) );
  INV_X1 U8889 ( .A(n7209), .ZN(P2_U3177) );
  OAI211_X1 U8890 ( .C1(n7212), .C2(n9103), .A(n7211), .B(n7210), .ZN(n7213)
         );
  INV_X1 U8891 ( .A(n7216), .ZN(n7215) );
  INV_X1 U8892 ( .A(n8915), .ZN(n8938) );
  OAI22_X1 U8893 ( .A1(n8942), .A2(n6313), .B1(n10384), .B2(n8899), .ZN(n7221)
         );
  NAND3_X1 U8894 ( .A1(n8340), .A2(n7217), .A3(n10073), .ZN(n7219) );
  AOI21_X1 U8895 ( .B1(n7219), .B2(n7218), .A(n8920), .ZN(n7220) );
  AOI211_X1 U8896 ( .C1(n8890), .C2(n8339), .A(n7221), .B(n7220), .ZN(n7222)
         );
  INV_X1 U8897 ( .A(n7222), .ZN(P2_U3233) );
  INV_X1 U8898 ( .A(n7833), .ZN(n7840) );
  INV_X1 U8899 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10401) );
  OAI222_X1 U8900 ( .A1(P1_U3086), .A2(n7840), .B1(n9884), .B2(n7223), .C1(
        n10401), .C2(n9882), .ZN(P1_U3339) );
  OAI21_X1 U8901 ( .B1(n7225), .B2(n7228), .A(n7224), .ZN(n7400) );
  INV_X1 U8902 ( .A(n7400), .ZN(n7233) );
  NAND2_X1 U8903 ( .A1(n7227), .A2(n7226), .ZN(n7229) );
  XNOR2_X1 U8904 ( .A(n7229), .B(n7228), .ZN(n7231) );
  AOI22_X1 U8905 ( .A1(n9727), .A2(n9305), .B1(n9303), .B2(n9728), .ZN(n7264)
         );
  INV_X1 U8906 ( .A(n7264), .ZN(n7230) );
  AOI21_X1 U8907 ( .B1(n7231), .B2(n9724), .A(n7230), .ZN(n7402) );
  OAI211_X1 U8908 ( .C1(n7232), .C2(n7421), .A(n9813), .B(n7411), .ZN(n7398)
         );
  OAI211_X1 U8909 ( .C1(n7233), .C2(n9804), .A(n7402), .B(n7398), .ZN(n7423)
         );
  OAI22_X1 U8910 ( .A1(n9823), .A2(n7421), .B1(n9988), .B2(n6891), .ZN(n7234)
         );
  AOI21_X1 U8911 ( .B1(n7423), .B2(n9988), .A(n7234), .ZN(n7235) );
  INV_X1 U8912 ( .A(n7235), .ZN(P1_U3525) );
  INV_X1 U8913 ( .A(n7236), .ZN(n7298) );
  AOI22_X1 U8914 ( .A1(n9433), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9871), .ZN(n7237) );
  OAI21_X1 U8915 ( .B1(n7298), .B2(n9884), .A(n7237), .ZN(P1_U3338) );
  INV_X1 U8916 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9328) );
  AND3_X1 U8917 ( .A1(n7240), .A2(n7239), .A3(n7238), .ZN(n7241) );
  NAND2_X1 U8918 ( .A1(n7242), .A2(n7241), .ZN(n7243) );
  AOI22_X1 U8919 ( .A1(n9148), .A2(n9304), .B1(n7395), .B2(n8233), .ZN(n7244)
         );
  XNOR2_X1 U8920 ( .A(n7244), .B(n8277), .ZN(n7273) );
  NAND2_X1 U8921 ( .A1(n9304), .A2(n9149), .ZN(n7246) );
  NAND2_X1 U8922 ( .A1(n7395), .A2(n9148), .ZN(n7245) );
  NAND2_X1 U8923 ( .A1(n7246), .A2(n7245), .ZN(n7271) );
  XNOR2_X1 U8924 ( .A(n7273), .B(n7271), .ZN(n7262) );
  NAND2_X1 U8925 ( .A1(n7249), .A2(n7250), .ZN(n7248) );
  INV_X1 U8926 ( .A(n7249), .ZN(n7252) );
  INV_X1 U8927 ( .A(n7250), .ZN(n7251) );
  NAND2_X1 U8928 ( .A1(n7256), .A2(n8233), .ZN(n7254) );
  NAND2_X1 U8929 ( .A1(n9305), .A2(n9148), .ZN(n7253) );
  XNOR2_X1 U8930 ( .A(n7255), .B(n8277), .ZN(n7260) );
  NAND2_X1 U8931 ( .A1(n9305), .A2(n9149), .ZN(n7258) );
  NAND2_X1 U8932 ( .A1(n7256), .A2(n9148), .ZN(n7257) );
  NAND2_X1 U8933 ( .A1(n7258), .A2(n7257), .ZN(n7259) );
  NAND2_X1 U8934 ( .A1(n7261), .A2(n7262), .ZN(n7276) );
  OAI21_X1 U8935 ( .B1(n7262), .B2(n7261), .A(n7276), .ZN(n7263) );
  NAND2_X1 U8936 ( .A1(n7263), .A2(n9906), .ZN(n7267) );
  INV_X1 U8937 ( .A(n9900), .ZN(n9911) );
  OAI22_X1 U8938 ( .A1(n9911), .A2(n7264), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9328), .ZN(n7265) );
  AOI21_X1 U8939 ( .B1(n7395), .B2(n9920), .A(n7265), .ZN(n7266) );
  OAI211_X1 U8940 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9923), .A(n7267), .B(
        n7266), .ZN(P1_U3218) );
  NAND2_X1 U8941 ( .A1(n9303), .A2(n9148), .ZN(n7269) );
  NAND2_X1 U8942 ( .A1(n7414), .A2(n8233), .ZN(n7268) );
  NAND2_X1 U8943 ( .A1(n7269), .A2(n7268), .ZN(n7270) );
  XNOR2_X1 U8944 ( .A(n7270), .B(n8277), .ZN(n7573) );
  AOI22_X1 U8945 ( .A1(n9149), .A2(n9303), .B1(n7414), .B2(n8306), .ZN(n7574)
         );
  XNOR2_X1 U8946 ( .A(n7573), .B(n7574), .ZN(n7274) );
  INV_X1 U8947 ( .A(n7271), .ZN(n7272) );
  NAND2_X1 U8948 ( .A1(n7273), .A2(n7272), .ZN(n7275) );
  NAND3_X1 U8949 ( .A1(n7276), .A2(n7274), .A3(n7275), .ZN(n7577) );
  NAND2_X1 U8950 ( .A1(n7577), .A2(n9906), .ZN(n7284) );
  AOI21_X1 U8951 ( .B1(n7276), .B2(n7275), .A(n7274), .ZN(n7283) );
  NAND2_X1 U8952 ( .A1(n9900), .A2(n9728), .ZN(n9890) );
  INV_X1 U8953 ( .A(n9890), .ZN(n7277) );
  INV_X1 U8954 ( .A(n9923), .ZN(n9269) );
  AOI22_X1 U8955 ( .A1(n7277), .A2(n9302), .B1(n7413), .B2(n9269), .ZN(n7282)
         );
  NAND2_X1 U8956 ( .A1(n9900), .A2(n9727), .ZN(n9279) );
  INV_X1 U8957 ( .A(n9279), .ZN(n7280) );
  OAI21_X1 U8958 ( .B1(n9903), .B2(n9957), .A(n7278), .ZN(n7279) );
  AOI21_X1 U8959 ( .B1(n7280), .B2(n9304), .A(n7279), .ZN(n7281) );
  OAI211_X1 U8960 ( .C1(n7284), .C2(n7283), .A(n7282), .B(n7281), .ZN(P1_U3230) );
  INV_X1 U8961 ( .A(n7286), .ZN(n7288) );
  NAND2_X1 U8962 ( .A1(n7288), .A2(n7287), .ZN(n7289) );
  XNOR2_X1 U8963 ( .A(n8198), .B(n10038), .ZN(n7425) );
  XNOR2_X1 U8964 ( .A(n7425), .B(n8929), .ZN(n7291) );
  OAI211_X1 U8965 ( .C1(n7292), .C2(n7291), .A(n7427), .B(n8515), .ZN(n7297)
         );
  AOI21_X1 U8966 ( .B1(n8534), .B2(n7448), .A(n7293), .ZN(n7294) );
  OAI21_X1 U8967 ( .B1(n8544), .B2(n7727), .A(n7294), .ZN(n7295) );
  AOI21_X1 U8968 ( .B1(n8548), .B2(n8564), .A(n7295), .ZN(n7296) );
  OAI211_X1 U8969 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8545), .A(n7297), .B(
        n7296), .ZN(P2_U3158) );
  INV_X1 U8970 ( .A(n8685), .ZN(n8664) );
  OAI222_X1 U8971 ( .A1(n9122), .A2(n7299), .B1(n9117), .B2(n7298), .C1(
        P2_U3151), .C2(n8664), .ZN(P2_U3278) );
  XOR2_X1 U8972 ( .A(n6677), .B(n7091), .Z(n7310) );
  AND2_X1 U8973 ( .A1(n7301), .A2(n7300), .ZN(n7724) );
  INV_X1 U8974 ( .A(n7724), .ZN(n8940) );
  NAND2_X1 U8975 ( .A1(n8927), .A2(n8940), .ZN(n7302) );
  XNOR2_X1 U8976 ( .A(n6677), .B(n7303), .ZN(n7304) );
  AOI222_X1 U8977 ( .A1(n8914), .A2(n7304), .B1(n8564), .B2(n8909), .C1(n8566), 
        .C2(n8911), .ZN(n7309) );
  MUX2_X1 U8978 ( .A(n7305), .B(n7309), .S(n8942), .Z(n7308) );
  AOI22_X1 U8979 ( .A1(n8890), .A2(n7306), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8937), .ZN(n7307) );
  OAI211_X1 U8980 ( .C1(n7310), .C2(n8923), .A(n7308), .B(n7307), .ZN(P2_U3232) );
  OAI21_X1 U8981 ( .B1(n10080), .B2(n7310), .A(n7309), .ZN(n7315) );
  INV_X1 U8982 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7311) );
  OAI22_X1 U8983 ( .A1(n6679), .A2(n9052), .B1(n10086), .B2(n7311), .ZN(n7312)
         );
  AOI21_X1 U8984 ( .B1(n7315), .B2(n10086), .A(n7312), .ZN(n7313) );
  INV_X1 U8985 ( .A(n7313), .ZN(P2_U3393) );
  OAI22_X1 U8986 ( .A1(n8980), .A2(n6679), .B1(n10099), .B2(n6799), .ZN(n7314)
         );
  AOI21_X1 U8987 ( .B1(n7315), .B2(n10099), .A(n7314), .ZN(n7316) );
  INV_X1 U8988 ( .A(n7316), .ZN(P2_U3460) );
  INV_X1 U8989 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7317) );
  OAI22_X1 U8990 ( .A1(n9864), .A2(n8338), .B1(n9860), .B2(n7317), .ZN(n7318)
         );
  INV_X1 U8991 ( .A(n7318), .ZN(n7319) );
  OAI21_X1 U8992 ( .B1(n7320), .B2(n6057), .A(n7319), .ZN(P1_U3459) );
  NAND2_X1 U8993 ( .A1(n7330), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7321) );
  OAI21_X1 U8994 ( .B1(n7330), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7321), .ZN(
        n9411) );
  OAI21_X1 U8995 ( .B1(n7323), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7322), .ZN(
        n9412) );
  NOR2_X1 U8996 ( .A1(n9411), .A2(n9412), .ZN(n9410) );
  AOI21_X1 U8997 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7330), .A(n9410), .ZN(
        n9425) );
  NAND2_X1 U8998 ( .A1(n7327), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7324) );
  OAI21_X1 U8999 ( .B1(n7327), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7324), .ZN(
        n9424) );
  NOR2_X1 U9000 ( .A1(n9425), .A2(n9424), .ZN(n9423) );
  AOI21_X1 U9001 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7327), .A(n9423), .ZN(
        n7561) );
  XNOR2_X1 U9002 ( .A(n7561), .B(n7560), .ZN(n7326) );
  INV_X1 U9003 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7325) );
  NOR2_X1 U9004 ( .A1(n7325), .A2(n7326), .ZN(n7562) );
  AOI211_X1 U9005 ( .C1(n7326), .C2(n7325), .A(n7562), .B(n9465), .ZN(n7340)
         );
  INV_X1 U9006 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9986) );
  OR2_X1 U9007 ( .A1(n7327), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7329) );
  NAND2_X1 U9008 ( .A1(n7327), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7328) );
  AND2_X1 U9009 ( .A1(n7329), .A2(n7328), .ZN(n9422) );
  INV_X1 U9010 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n8165) );
  MUX2_X1 U9011 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n8165), .S(n7330), .Z(n9408)
         );
  AOI21_X1 U9012 ( .B1(n7332), .B2(n6954), .A(n7331), .ZN(n9409) );
  NAND2_X1 U9013 ( .A1(n9408), .A2(n9409), .ZN(n9407) );
  OAI21_X1 U9014 ( .B1(n9404), .B2(n8165), .A(n9407), .ZN(n9421) );
  NAND2_X1 U9015 ( .A1(n9422), .A2(n9421), .ZN(n9420) );
  OAI21_X1 U9016 ( .B1(n9986), .B2(n9417), .A(n9420), .ZN(n7554) );
  INV_X1 U9017 ( .A(n7554), .ZN(n7333) );
  XNOR2_X1 U9018 ( .A(n7555), .B(n7333), .ZN(n7334) );
  NAND2_X1 U9019 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7334), .ZN(n7556) );
  OAI21_X1 U9020 ( .B1(n7334), .B2(P1_REG1_REG_15__SCAN_IN), .A(n7556), .ZN(
        n7335) );
  NOR2_X1 U9021 ( .A1(n9464), .A2(n7335), .ZN(n7339) );
  NOR2_X1 U9022 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9277), .ZN(n7336) );
  AOI21_X1 U9023 ( .B1(n9933), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n7336), .ZN(
        n7337) );
  OAI21_X1 U9024 ( .B1(n9459), .B2(n7560), .A(n7337), .ZN(n7338) );
  OR3_X1 U9025 ( .A1(n7340), .A2(n7339), .A3(n7338), .ZN(P1_U3258) );
  MUX2_X1 U9026 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8699), .Z(n7701) );
  XOR2_X1 U9027 ( .A(n7700), .B(n7701), .Z(n7344) );
  OAI21_X1 U9028 ( .B1(n7345), .B2(n7344), .A(n7702), .ZN(n7370) );
  INV_X1 U9029 ( .A(n7346), .ZN(n7347) );
  NOR2_X1 U9030 ( .A1(n7360), .A2(n7347), .ZN(n7348) );
  NOR2_X1 U9031 ( .A1(n7349), .A2(n7348), .ZN(n7353) );
  NAND2_X1 U9032 ( .A1(n7700), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7708) );
  OR2_X1 U9033 ( .A1(n7700), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7350) );
  NAND2_X1 U9034 ( .A1(n7708), .A2(n7350), .ZN(n7352) );
  INV_X1 U9035 ( .A(n7709), .ZN(n7351) );
  AOI21_X1 U9036 ( .B1(n7353), .B2(n7352), .A(n7351), .ZN(n7357) );
  INV_X1 U9037 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7354) );
  NOR2_X1 U9038 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7354), .ZN(n7598) );
  INV_X1 U9039 ( .A(n7598), .ZN(n7356) );
  NAND2_X1 U9040 ( .A1(n10018), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7355) );
  OAI211_X1 U9041 ( .C1(n7357), .C2(n10026), .A(n7356), .B(n7355), .ZN(n7369)
         );
  NOR2_X1 U9042 ( .A1(n7360), .A2(n7359), .ZN(n7362) );
  NAND2_X1 U9043 ( .A1(n7700), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7690) );
  OR2_X1 U9044 ( .A1(n7700), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U9045 ( .A1(n7690), .A2(n7363), .ZN(n7365) );
  INV_X1 U9046 ( .A(n7691), .ZN(n7364) );
  AOI21_X1 U9047 ( .B1(n7366), .B2(n7365), .A(n7364), .ZN(n7367) );
  OAI22_X1 U9048 ( .A1(n7367), .A2(n10022), .B1(n7700), .B2(n8679), .ZN(n7368)
         );
  AOI211_X1 U9049 ( .C1(n7370), .C2(n10020), .A(n7369), .B(n7368), .ZN(n7371)
         );
  INV_X1 U9050 ( .A(n7371), .ZN(P2_U3188) );
  INV_X1 U9051 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7372) );
  OAI22_X1 U9052 ( .A1(n9864), .A2(n9944), .B1(n9860), .B2(n7372), .ZN(n7373)
         );
  AOI21_X1 U9053 ( .B1(n7374), .B2(n9860), .A(n7373), .ZN(n7375) );
  INV_X1 U9054 ( .A(n7375), .ZN(P1_U3456) );
  OAI21_X1 U9055 ( .B1(n7377), .B2(n7379), .A(n7376), .ZN(n7478) );
  INV_X1 U9056 ( .A(n7470), .ZN(n7378) );
  AOI211_X1 U9057 ( .C1(n7578), .C2(n7412), .A(n9969), .B(n7378), .ZN(n7482)
         );
  XNOR2_X1 U9058 ( .A(n5769), .B(n7379), .ZN(n7383) );
  NAND2_X1 U9059 ( .A1(n9303), .A2(n9727), .ZN(n7381) );
  NAND2_X1 U9060 ( .A1(n9301), .A2(n9728), .ZN(n7380) );
  NAND2_X1 U9061 ( .A1(n7381), .A2(n7380), .ZN(n7582) );
  INV_X1 U9062 ( .A(n7582), .ZN(n7382) );
  OAI21_X1 U9063 ( .B1(n7383), .B2(n9659), .A(n7382), .ZN(n7483) );
  AOI211_X1 U9064 ( .C1(n9979), .C2(n7478), .A(n7482), .B(n7483), .ZN(n7388)
         );
  OAI22_X1 U9065 ( .A1(n9864), .A2(n7584), .B1(n9860), .B2(n5371), .ZN(n7384)
         );
  INV_X1 U9066 ( .A(n7384), .ZN(n7385) );
  OAI21_X1 U9067 ( .B1(n7388), .B2(n6057), .A(n7385), .ZN(P1_U3468) );
  OAI22_X1 U9068 ( .A1(n9823), .A2(n7584), .B1(n9988), .B2(n5374), .ZN(n7386)
         );
  INV_X1 U9069 ( .A(n7386), .ZN(n7387) );
  OAI21_X1 U9070 ( .B1(n7388), .B2(n9985), .A(n7387), .ZN(P1_U3527) );
  NAND2_X1 U9071 ( .A1(n7390), .A2(n7389), .ZN(n7392) );
  AND2_X2 U9072 ( .A1(n7392), .A2(n9711), .ZN(n9612) );
  AND2_X1 U9073 ( .A1(n7658), .A2(n9946), .ZN(n7391) );
  INV_X1 U9074 ( .A(n7392), .ZN(n7393) );
  NAND2_X1 U9075 ( .A1(n7393), .A2(n7033), .ZN(n9646) );
  INV_X1 U9076 ( .A(n9711), .ZN(n9942) );
  AOI22_X1 U9077 ( .A1(n9612), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9942), .B2(
        n9328), .ZN(n7397) );
  NAND2_X1 U9078 ( .A1(n9642), .A2(n7395), .ZN(n7396) );
  OAI211_X1 U9079 ( .C1(n7398), .C2(n9646), .A(n7397), .B(n7396), .ZN(n7399)
         );
  AOI21_X1 U9080 ( .B1(n7400), .B2(n9707), .A(n7399), .ZN(n7401) );
  OAI21_X1 U9081 ( .B1(n7402), .B2(n9612), .A(n7401), .ZN(P1_U3290) );
  INV_X1 U9082 ( .A(n7409), .ZN(n7403) );
  XNOR2_X1 U9083 ( .A(n7404), .B(n7403), .ZN(n7405) );
  NAND2_X1 U9084 ( .A1(n7405), .A2(n9724), .ZN(n7407) );
  AOI22_X1 U9085 ( .A1(n9302), .A2(n9728), .B1(n9727), .B2(n9304), .ZN(n7406)
         );
  NAND2_X1 U9086 ( .A1(n7407), .A2(n7406), .ZN(n9959) );
  INV_X1 U9087 ( .A(n9959), .ZN(n7419) );
  OAI21_X1 U9088 ( .B1(n7410), .B2(n7409), .A(n7408), .ZN(n9961) );
  OAI21_X1 U9089 ( .B1(n4706), .B2(n9957), .A(n7412), .ZN(n9958) );
  OR2_X1 U9090 ( .A1(n9646), .A2(n9969), .ZN(n9490) );
  AOI22_X1 U9091 ( .A1(n9612), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7413), .B2(
        n9942), .ZN(n7416) );
  NAND2_X1 U9092 ( .A1(n9642), .A2(n7414), .ZN(n7415) );
  OAI211_X1 U9093 ( .C1(n9958), .C2(n9490), .A(n7416), .B(n7415), .ZN(n7417)
         );
  AOI21_X1 U9094 ( .B1(n9961), .B2(n9707), .A(n7417), .ZN(n7418) );
  OAI21_X1 U9095 ( .B1(n7419), .B2(n9612), .A(n7418), .ZN(P1_U3289) );
  INV_X1 U9096 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7420) );
  OAI22_X1 U9097 ( .A1(n9864), .A2(n7421), .B1(n9860), .B2(n7420), .ZN(n7422)
         );
  AOI21_X1 U9098 ( .B1(n7423), .B2(n9860), .A(n7422), .ZN(n7424) );
  INV_X1 U9099 ( .A(n7424), .ZN(P1_U3462) );
  NAND2_X1 U9100 ( .A1(n8563), .A2(n7425), .ZN(n7426) );
  XNOR2_X1 U9101 ( .A(n8198), .B(n10044), .ZN(n7428) );
  NAND2_X1 U9102 ( .A1(n6526), .A2(n7428), .ZN(n7430) );
  INV_X1 U9103 ( .A(n7428), .ZN(n7429) );
  NAND2_X1 U9104 ( .A1(n7429), .A2(n7727), .ZN(n7519) );
  AND2_X1 U9105 ( .A1(n7430), .A2(n7519), .ZN(n7431) );
  OAI21_X1 U9106 ( .B1(n7432), .B2(n7431), .A(n7520), .ZN(n7433) );
  NAND2_X1 U9107 ( .A1(n7433), .A2(n8515), .ZN(n7438) );
  AOI21_X1 U9108 ( .B1(n8534), .B2(n7506), .A(n7434), .ZN(n7435) );
  OAI21_X1 U9109 ( .B1(n8544), .B2(n7590), .A(n7435), .ZN(n7436) );
  AOI21_X1 U9110 ( .B1(n8548), .B2(n8563), .A(n7436), .ZN(n7437) );
  OAI211_X1 U9111 ( .C1(n7504), .C2(n8545), .A(n7438), .B(n7437), .ZN(P2_U3170) );
  NAND3_X1 U9112 ( .A1(n7440), .A2(n7441), .A3(n7443), .ZN(n7442) );
  AND2_X1 U9113 ( .A1(n7439), .A2(n7442), .ZN(n10039) );
  XNOR2_X1 U9114 ( .A(n7444), .B(n7443), .ZN(n7445) );
  AOI222_X1 U9115 ( .A1(n8914), .A2(n7445), .B1(n6526), .B2(n8909), .C1(n8564), 
        .C2(n8911), .ZN(n10037) );
  MUX2_X1 U9116 ( .A(n7446), .B(n10037), .S(n8942), .Z(n7450) );
  AOI22_X1 U9117 ( .A1(n8890), .A2(n7448), .B1(n8937), .B2(n7447), .ZN(n7449)
         );
  OAI211_X1 U9118 ( .C1(n10039), .C2(n8923), .A(n7450), .B(n7449), .ZN(
        P2_U3230) );
  INV_X1 U9119 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10371) );
  INV_X1 U9120 ( .A(n7451), .ZN(n7460) );
  INV_X1 U9121 ( .A(n9454), .ZN(n9430) );
  OAI222_X1 U9122 ( .A1(n9882), .A2(n10371), .B1(n9884), .B2(n7460), .C1(
        P1_U3086), .C2(n9430), .ZN(P1_U3337) );
  OAI21_X1 U9123 ( .B1(n7454), .B2(n7453), .A(n7452), .ZN(n7458) );
  INV_X1 U9124 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7455) );
  INV_X1 U9125 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9894) );
  OAI22_X1 U9126 ( .A1(n9714), .A2(n7455), .B1(n9894), .B2(n9711), .ZN(n7457)
         );
  AOI21_X1 U9127 ( .B1(n9945), .B2(n9490), .A(n9888), .ZN(n7456) );
  AOI211_X1 U9128 ( .C1(n9714), .C2(n7458), .A(n7457), .B(n7456), .ZN(n7459)
         );
  INV_X1 U9129 ( .A(n7459), .ZN(P1_U3293) );
  INV_X1 U9130 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7461) );
  INV_X1 U9131 ( .A(n8697), .ZN(n8687) );
  OAI222_X1 U9132 ( .A1(n9122), .A2(n7461), .B1(n8687), .B2(P2_U3151), .C1(
        n9117), .C2(n7460), .ZN(P2_U3277) );
  OAI21_X1 U9133 ( .B1(n7463), .B2(n7465), .A(n7462), .ZN(n7464) );
  INV_X1 U9134 ( .A(n7464), .ZN(n7489) );
  XOR2_X1 U9135 ( .A(n7466), .B(n7465), .Z(n7468) );
  OAI22_X1 U9136 ( .A1(n7467), .A2(n9664), .B1(n7572), .B2(n9662), .ZN(n7676)
         );
  AOI21_X1 U9137 ( .B1(n7468), .B2(n9724), .A(n7676), .ZN(n7488) );
  MUX2_X1 U9138 ( .A(n6919), .B(n7488), .S(n9714), .Z(n7477) );
  INV_X1 U9139 ( .A(n7546), .ZN(n7472) );
  AOI21_X1 U9140 ( .B1(n7470), .B2(n7469), .A(n9969), .ZN(n7471) );
  NAND2_X1 U9141 ( .A1(n7472), .A2(n7471), .ZN(n7487) );
  INV_X1 U9142 ( .A(n7487), .ZN(n7475) );
  INV_X1 U9143 ( .A(n7473), .ZN(n7679) );
  OAI22_X1 U9144 ( .A1(n9945), .A2(n7674), .B1(n9711), .B2(n7679), .ZN(n7474)
         );
  AOI21_X1 U9145 ( .B1(n7475), .B2(n9950), .A(n7474), .ZN(n7476) );
  OAI211_X1 U9146 ( .C1(n7489), .C2(n9741), .A(n7477), .B(n7476), .ZN(P1_U3287) );
  INV_X1 U9147 ( .A(n7478), .ZN(n7486) );
  NOR2_X1 U9148 ( .A1(n9945), .A2(n7584), .ZN(n7481) );
  OAI22_X1 U9149 ( .A1(n9714), .A2(n7479), .B1(n7581), .B2(n9711), .ZN(n7480)
         );
  AOI211_X1 U9150 ( .C1(n7482), .C2(n9950), .A(n7481), .B(n7480), .ZN(n7485)
         );
  NAND2_X1 U9151 ( .A1(n7483), .A2(n9714), .ZN(n7484) );
  OAI211_X1 U9152 ( .C1(n7486), .C2(n9741), .A(n7485), .B(n7484), .ZN(P1_U3288) );
  OAI211_X1 U9153 ( .C1(n7489), .C2(n9804), .A(n7488), .B(n7487), .ZN(n7495)
         );
  INV_X1 U9154 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7490) );
  OAI22_X1 U9155 ( .A1(n9864), .A2(n7674), .B1(n9860), .B2(n7490), .ZN(n7491)
         );
  AOI21_X1 U9156 ( .B1(n7495), .B2(n9860), .A(n7491), .ZN(n7492) );
  INV_X1 U9157 ( .A(n7492), .ZN(P1_U3471) );
  OAI22_X1 U9158 ( .A1(n9823), .A2(n7674), .B1(n9988), .B2(n7493), .ZN(n7494)
         );
  AOI21_X1 U9159 ( .B1(n7495), .B2(n9988), .A(n7494), .ZN(n7496) );
  INV_X1 U9160 ( .A(n7496), .ZN(P1_U3528) );
  NOR2_X1 U9161 ( .A1(n7501), .A2(n7497), .ZN(n7500) );
  INV_X1 U9162 ( .A(n7498), .ZN(n7499) );
  AOI21_X1 U9163 ( .B1(n7500), .B2(n7439), .A(n7499), .ZN(n10045) );
  XNOR2_X1 U9164 ( .A(n7502), .B(n7501), .ZN(n7503) );
  AOI222_X1 U9165 ( .A1(n8914), .A2(n7503), .B1(n8563), .B2(n8911), .C1(n8562), 
        .C2(n8909), .ZN(n10043) );
  MUX2_X1 U9166 ( .A(n6832), .B(n10043), .S(n8942), .Z(n7508) );
  INV_X1 U9167 ( .A(n7504), .ZN(n7505) );
  AOI22_X1 U9168 ( .A1(n8890), .A2(n7506), .B1(n8937), .B2(n7505), .ZN(n7507)
         );
  OAI211_X1 U9169 ( .C1(n10045), .C2(n8923), .A(n7508), .B(n7507), .ZN(
        P2_U3229) );
  NOR2_X1 U9170 ( .A1(n9711), .A2(n7509), .ZN(n7511) );
  AOI211_X1 U9171 ( .C1(n7512), .C2(n7033), .A(n7511), .B(n7510), .ZN(n7516)
         );
  OAI22_X1 U9172 ( .A1(n9945), .A2(n8338), .B1(n6910), .B2(n9714), .ZN(n7513)
         );
  AOI21_X1 U9173 ( .B1(n7514), .B2(n9707), .A(n7513), .ZN(n7515) );
  OAI21_X1 U9174 ( .B1(n7516), .B2(n9612), .A(n7515), .ZN(P1_U3291) );
  INV_X1 U9175 ( .A(n7520), .ZN(n7518) );
  INV_X1 U9176 ( .A(n7519), .ZN(n7517) );
  XNOR2_X1 U9177 ( .A(n8198), .B(n10048), .ZN(n7589) );
  XNOR2_X1 U9178 ( .A(n7589), .B(n7590), .ZN(n7521) );
  NOR3_X1 U9179 ( .A1(n7518), .A2(n7517), .A3(n7521), .ZN(n7524) );
  NAND2_X1 U9180 ( .A1(n7520), .A2(n7519), .ZN(n7522) );
  INV_X1 U9181 ( .A(n7593), .ZN(n7523) );
  OAI21_X1 U9182 ( .B1(n7524), .B2(n7523), .A(n8515), .ZN(n7529) );
  AOI21_X1 U9183 ( .B1(n8534), .B2(n7735), .A(n7525), .ZN(n7526) );
  OAI21_X1 U9184 ( .B1(n8544), .B2(n7792), .A(n7526), .ZN(n7527) );
  AOI21_X1 U9185 ( .B1(n8548), .B2(n6526), .A(n7527), .ZN(n7528) );
  OAI211_X1 U9186 ( .C1(n7733), .C2(n8545), .A(n7529), .B(n7528), .ZN(P2_U3167) );
  INV_X1 U9187 ( .A(n7530), .ZN(n7533) );
  OAI222_X1 U9188 ( .A1(n9122), .A2(n7532), .B1(n9117), .B2(n7533), .C1(n7531), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U9189 ( .A1(n7033), .A2(P1_U3086), .B1(n9884), .B2(n7533), .C1(
        n10508), .C2(n9882), .ZN(P1_U3336) );
  OR2_X1 U9190 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  AOI22_X1 U9191 ( .A1(n9299), .A2(n9728), .B1(n9727), .B2(n9301), .ZN(n7544)
         );
  NAND3_X1 U9192 ( .A1(n7540), .A2(n7538), .A3(n7539), .ZN(n7635) );
  INV_X1 U9193 ( .A(n7635), .ZN(n7542) );
  AOI21_X1 U9194 ( .B1(n7540), .B2(n7539), .A(n7538), .ZN(n7541) );
  OAI21_X1 U9195 ( .B1(n7542), .B2(n7541), .A(n9724), .ZN(n7543) );
  OAI211_X1 U9196 ( .C1(n7738), .C2(n7658), .A(n7544), .B(n7543), .ZN(n7739)
         );
  INV_X1 U9197 ( .A(n7545), .ZN(n7661) );
  OAI21_X1 U9198 ( .B1(n7630), .B2(n7546), .A(n7661), .ZN(n7748) );
  OAI22_X1 U9199 ( .A1(n7738), .A2(n7758), .B1(n9969), .B2(n7748), .ZN(n7547)
         );
  NOR2_X1 U9200 ( .A1(n7739), .A2(n7547), .ZN(n7553) );
  OAI22_X1 U9201 ( .A1(n7630), .A2(n9823), .B1(n9988), .B2(n6899), .ZN(n7548)
         );
  INV_X1 U9202 ( .A(n7548), .ZN(n7549) );
  OAI21_X1 U9203 ( .B1(n7553), .B2(n9985), .A(n7549), .ZN(P1_U3529) );
  INV_X1 U9204 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7550) );
  OAI22_X1 U9205 ( .A1(n9864), .A2(n7630), .B1(n9860), .B2(n7550), .ZN(n7551)
         );
  INV_X1 U9206 ( .A(n7551), .ZN(n7552) );
  OAI21_X1 U9207 ( .B1(n7553), .B2(n6057), .A(n7552), .ZN(P1_U3474) );
  NAND2_X1 U9208 ( .A1(n7555), .A2(n7554), .ZN(n7557) );
  NAND2_X1 U9209 ( .A1(n7557), .A2(n7556), .ZN(n7559) );
  XNOR2_X1 U9210 ( .A(n7833), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7558) );
  NOR2_X1 U9211 ( .A1(n7558), .A2(n7559), .ZN(n7838) );
  AOI21_X1 U9212 ( .B1(n7559), .B2(n7558), .A(n7838), .ZN(n7571) );
  NOR2_X1 U9213 ( .A1(n7561), .A2(n7560), .ZN(n7563) );
  NOR2_X1 U9214 ( .A1(n7563), .A2(n7562), .ZN(n7565) );
  AOI22_X1 U9215 ( .A1(n7833), .A2(n9713), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n7840), .ZN(n7564) );
  NOR2_X1 U9216 ( .A1(n7565), .A2(n7564), .ZN(n7832) );
  AOI211_X1 U9217 ( .C1(n7565), .C2(n7564), .A(n7832), .B(n9465), .ZN(n7566)
         );
  INV_X1 U9218 ( .A(n7566), .ZN(n7570) );
  AND2_X1 U9219 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7568) );
  NOR2_X1 U9220 ( .A1(n9459), .A2(n7840), .ZN(n7567) );
  AOI211_X1 U9221 ( .C1(n9933), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n7568), .B(
        n7567), .ZN(n7569) );
  OAI211_X1 U9222 ( .C1(n7571), .C2(n9464), .A(n7570), .B(n7569), .ZN(P1_U3259) );
  OAI22_X1 U9223 ( .A1(n7572), .A2(n8310), .B1(n7584), .B2(n8284), .ZN(n7608)
         );
  AOI22_X1 U9224 ( .A1(n9302), .A2(n8306), .B1(n7578), .B2(n8233), .ZN(n7579)
         );
  XOR2_X1 U9225 ( .A(n8277), .B(n7579), .Z(n7607) );
  INV_X1 U9226 ( .A(n7607), .ZN(n7615) );
  NAND2_X1 U9227 ( .A1(n7619), .A2(n7615), .ZN(n7667) );
  OAI21_X1 U9228 ( .B1(n7619), .B2(n7615), .A(n7667), .ZN(n7580) );
  NOR2_X1 U9229 ( .A1(n7580), .A2(n7608), .ZN(n7670) );
  AOI21_X1 U9230 ( .B1(n7608), .B2(n7580), .A(n7670), .ZN(n7588) );
  INV_X1 U9231 ( .A(n9906), .ZN(n9916) );
  INV_X1 U9232 ( .A(n7581), .ZN(n7586) );
  NAND2_X1 U9233 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9334) );
  NAND2_X1 U9234 ( .A1(n9900), .A2(n7582), .ZN(n7583) );
  OAI211_X1 U9235 ( .C1(n9903), .C2(n7584), .A(n9334), .B(n7583), .ZN(n7585)
         );
  AOI21_X1 U9236 ( .B1(n7586), .B2(n9269), .A(n7585), .ZN(n7587) );
  OAI21_X1 U9237 ( .B1(n7588), .B2(n9916), .A(n7587), .ZN(P1_U3227) );
  INV_X1 U9238 ( .A(n7589), .ZN(n7591) );
  NAND2_X1 U9239 ( .A1(n7591), .A2(n7590), .ZN(n7592) );
  XNOR2_X1 U9240 ( .A(n8198), .B(n7754), .ZN(n7850) );
  XNOR2_X1 U9241 ( .A(n7850), .B(n8561), .ZN(n7595) );
  AOI21_X1 U9242 ( .B1(n7594), .B2(n7595), .A(n8538), .ZN(n7597) );
  INV_X1 U9243 ( .A(n7595), .ZN(n7596) );
  NAND2_X1 U9244 ( .A1(n7597), .A2(n7852), .ZN(n7602) );
  AOI21_X1 U9245 ( .B1(n8534), .B2(n7687), .A(n7598), .ZN(n7599) );
  OAI21_X1 U9246 ( .B1(n8544), .B2(n7854), .A(n7599), .ZN(n7600) );
  AOI21_X1 U9247 ( .B1(n8548), .B2(n8562), .A(n7600), .ZN(n7601) );
  OAI211_X1 U9248 ( .C1(n7685), .C2(n8545), .A(n7602), .B(n7601), .ZN(P2_U3179) );
  OR2_X1 U9249 ( .A1(n7630), .A2(n8284), .ZN(n7604) );
  NAND2_X1 U9250 ( .A1(n9300), .A2(n9149), .ZN(n7603) );
  NAND2_X1 U9251 ( .A1(n7604), .A2(n7603), .ZN(n7975) );
  NAND2_X1 U9252 ( .A1(n9300), .A2(n9148), .ZN(n7605) );
  OAI21_X1 U9253 ( .B1(n7630), .B2(n8293), .A(n7605), .ZN(n7606) );
  XNOR2_X1 U9254 ( .A(n7606), .B(n8277), .ZN(n7974) );
  INV_X1 U9255 ( .A(n7608), .ZN(n7614) );
  NAND2_X1 U9256 ( .A1(n9301), .A2(n9148), .ZN(n7609) );
  OAI21_X1 U9257 ( .B1(n7674), .B2(n8293), .A(n7609), .ZN(n7610) );
  XNOR2_X1 U9258 ( .A(n7610), .B(n8277), .ZN(n7613) );
  NAND2_X1 U9259 ( .A1(n9301), .A2(n9149), .ZN(n7611) );
  OAI21_X1 U9260 ( .B1(n7674), .B2(n8284), .A(n7611), .ZN(n7612) );
  NOR2_X1 U9261 ( .A1(n7613), .A2(n7612), .ZN(n7620) );
  AOI21_X1 U9262 ( .B1(n7613), .B2(n7612), .A(n7620), .ZN(n7669) );
  INV_X1 U9263 ( .A(n7620), .ZN(n7621) );
  OAI21_X1 U9264 ( .B1(n7623), .B2(n7622), .A(n7995), .ZN(n7624) );
  NAND2_X1 U9265 ( .A1(n7624), .A2(n9906), .ZN(n7629) );
  INV_X1 U9266 ( .A(n7743), .ZN(n7627) );
  AND2_X1 U9267 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9371) );
  OAI22_X1 U9268 ( .A1(n7625), .A2(n9279), .B1(n9890), .B2(n7999), .ZN(n7626)
         );
  AOI211_X1 U9269 ( .C1(n7627), .C2(n9269), .A(n9371), .B(n7626), .ZN(n7628)
         );
  OAI211_X1 U9270 ( .C1(n7630), .C2(n9903), .A(n7629), .B(n7628), .ZN(P1_U3213) );
  NAND2_X1 U9271 ( .A1(n7650), .A2(n7924), .ZN(n7632) );
  OAI211_X1 U9272 ( .C1(n7633), .C2(n9882), .A(n7632), .B(n7631), .ZN(P1_U3335) );
  NAND2_X1 U9273 ( .A1(n7635), .A2(n7634), .ZN(n7657) );
  INV_X1 U9274 ( .A(n7636), .ZN(n7638) );
  OAI21_X1 U9275 ( .B1(n7657), .B2(n7638), .A(n7637), .ZN(n7639) );
  XNOR2_X1 U9276 ( .A(n7639), .B(n7642), .ZN(n7640) );
  AOI22_X1 U9277 ( .A1(n7640), .A2(n9724), .B1(n9727), .B2(n9299), .ZN(n9964)
         );
  OAI21_X1 U9278 ( .B1(n7643), .B2(n7642), .A(n7641), .ZN(n9967) );
  NAND2_X1 U9279 ( .A1(n9967), .A2(n9707), .ZN(n7649) );
  OAI22_X1 U9280 ( .A1(n9714), .A2(n7644), .B1(n7998), .B2(n9711), .ZN(n7647)
         );
  XNOR2_X1 U9281 ( .A(n7777), .B(n7987), .ZN(n7645) );
  AOI22_X1 U9282 ( .A1(n7645), .A2(n9813), .B1(n9728), .B2(n9297), .ZN(n9963)
         );
  NOR2_X1 U9283 ( .A1(n9963), .A2(n9646), .ZN(n7646) );
  AOI211_X1 U9284 ( .C1(n9642), .C2(n7987), .A(n7647), .B(n7646), .ZN(n7648)
         );
  OAI211_X1 U9285 ( .C1(n9612), .C2(n9964), .A(n7649), .B(n7648), .ZN(P1_U3284) );
  INV_X1 U9286 ( .A(n7650), .ZN(n7653) );
  OAI222_X1 U9287 ( .A1(n9117), .A2(n7653), .B1(P2_U3151), .B2(n7652), .C1(
        n7651), .C2(n9105), .ZN(P2_U3275) );
  INV_X1 U9288 ( .A(n9946), .ZN(n7741) );
  OAI21_X1 U9289 ( .B1(n7655), .B2(n7656), .A(n7654), .ZN(n7761) );
  XNOR2_X1 U9290 ( .A(n7657), .B(n7656), .ZN(n7660) );
  INV_X1 U9291 ( .A(n7658), .ZN(n9940) );
  NAND2_X1 U9292 ( .A1(n7761), .A2(n9940), .ZN(n7659) );
  AOI22_X1 U9293 ( .A1(n9298), .A2(n9728), .B1(n9727), .B2(n9300), .ZN(n9912)
         );
  OAI211_X1 U9294 ( .C1(n9659), .C2(n7660), .A(n7659), .B(n9912), .ZN(n7759)
         );
  AOI21_X1 U9295 ( .B1(n7741), .B2(n7761), .A(n7759), .ZN(n7666) );
  AOI211_X1 U9296 ( .C1(n9921), .C2(n7661), .A(n9969), .B(n7777), .ZN(n7760)
         );
  NOR2_X1 U9297 ( .A1(n9945), .A2(n7764), .ZN(n7664) );
  OAI22_X1 U9298 ( .A1(n9714), .A2(n7662), .B1(n9924), .B2(n9711), .ZN(n7663)
         );
  AOI211_X1 U9299 ( .C1(n7760), .C2(n9950), .A(n7664), .B(n7663), .ZN(n7665)
         );
  OAI21_X1 U9300 ( .B1(n7666), .B2(n9612), .A(n7665), .ZN(P1_U3285) );
  INV_X1 U9301 ( .A(n7667), .ZN(n7668) );
  NOR3_X1 U9302 ( .A1(n7670), .A2(n7669), .A3(n7668), .ZN(n7673) );
  INV_X1 U9303 ( .A(n7671), .ZN(n7672) );
  OAI21_X1 U9304 ( .B1(n7673), .B2(n7672), .A(n9906), .ZN(n7678) );
  AND2_X1 U9305 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9350) );
  NOR2_X1 U9306 ( .A1(n9903), .A2(n7674), .ZN(n7675) );
  AOI211_X1 U9307 ( .C1(n9900), .C2(n7676), .A(n9350), .B(n7675), .ZN(n7677)
         );
  OAI211_X1 U9308 ( .C1(n9923), .C2(n7679), .A(n7678), .B(n7677), .ZN(P1_U3239) );
  XNOR2_X1 U9309 ( .A(n7680), .B(n7682), .ZN(n7750) );
  XNOR2_X1 U9310 ( .A(n7681), .B(n7682), .ZN(n7683) );
  AOI222_X1 U9311 ( .A1(n8914), .A2(n7683), .B1(n8560), .B2(n8909), .C1(n8562), 
        .C2(n8911), .ZN(n7749) );
  MUX2_X1 U9312 ( .A(n7684), .B(n7749), .S(n8942), .Z(n7689) );
  INV_X1 U9313 ( .A(n7685), .ZN(n7686) );
  AOI22_X1 U9314 ( .A1(n8890), .A2(n7687), .B1(n8937), .B2(n7686), .ZN(n7688)
         );
  OAI211_X1 U9315 ( .C1(n8923), .C2(n7750), .A(n7689), .B(n7688), .ZN(P2_U3227) );
  INV_X1 U9316 ( .A(n7693), .ZN(n7692) );
  NOR2_X1 U9317 ( .A1(n10013), .A2(n7692), .ZN(n7694) );
  NAND2_X1 U9318 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7822), .ZN(n7695) );
  OAI21_X1 U9319 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7822), .A(n7695), .ZN(
        n7696) );
  AOI21_X1 U9320 ( .B1(n7697), .B2(n7696), .A(n7812), .ZN(n7722) );
  MUX2_X1 U9321 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8699), .Z(n7816) );
  XNOR2_X1 U9322 ( .A(n7816), .B(n7698), .ZN(n7706) );
  MUX2_X1 U9323 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8699), .Z(n7699) );
  OR2_X1 U9324 ( .A1(n7699), .A2(n7711), .ZN(n7704) );
  XNOR2_X1 U9325 ( .A(n7699), .B(n10013), .ZN(n10017) );
  OR2_X1 U9326 ( .A1(n7701), .A2(n7700), .ZN(n7703) );
  NAND2_X1 U9327 ( .A1(n7703), .A2(n7702), .ZN(n10016) );
  NAND2_X1 U9328 ( .A1(n10017), .A2(n10016), .ZN(n10015) );
  NAND2_X1 U9329 ( .A1(n7704), .A2(n10015), .ZN(n7705) );
  NAND2_X1 U9330 ( .A1(n7706), .A2(n7705), .ZN(n7817) );
  OAI21_X1 U9331 ( .B1(n7706), .B2(n7705), .A(n7817), .ZN(n7720) );
  NOR2_X1 U9332 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6088), .ZN(n7958) );
  AOI21_X1 U9333 ( .B1(n10018), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7958), .ZN(
        n7707) );
  OAI21_X1 U9334 ( .B1(n7822), .B2(n8679), .A(n7707), .ZN(n7719) );
  INV_X1 U9335 ( .A(n7712), .ZN(n7710) );
  NOR2_X1 U9336 ( .A1(n10013), .A2(n7710), .ZN(n7713) );
  NAND2_X1 U9337 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7822), .ZN(n7714) );
  OAI21_X1 U9338 ( .B1(n7822), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7714), .ZN(
        n7715) );
  AOI21_X1 U9339 ( .B1(n7716), .B2(n7715), .A(n7821), .ZN(n7717) );
  NOR2_X1 U9340 ( .A1(n7717), .A2(n10026), .ZN(n7718) );
  AOI211_X1 U9341 ( .C1(n10020), .C2(n7720), .A(n7719), .B(n7718), .ZN(n7721)
         );
  OAI21_X1 U9342 ( .B1(n7722), .B2(n10022), .A(n7721), .ZN(P2_U3190) );
  XNOR2_X1 U9343 ( .A(n7723), .B(n7726), .ZN(n10049) );
  NAND2_X1 U9344 ( .A1(n8942), .A2(n7724), .ZN(n8327) );
  XOR2_X1 U9345 ( .A(n7725), .B(n7726), .Z(n7729) );
  OAI22_X1 U9346 ( .A1(n7792), .A2(n8928), .B1(n7727), .B2(n8930), .ZN(n7728)
         );
  AOI21_X1 U9347 ( .B1(n7729), .B2(n8914), .A(n7728), .ZN(n7730) );
  OAI21_X1 U9348 ( .B1(n10049), .B2(n8927), .A(n7730), .ZN(n10051) );
  INV_X1 U9349 ( .A(n10051), .ZN(n7731) );
  MUX2_X1 U9350 ( .A(n7732), .B(n7731), .S(n8942), .Z(n7737) );
  INV_X1 U9351 ( .A(n7733), .ZN(n7734) );
  AOI22_X1 U9352 ( .A1(n8890), .A2(n7735), .B1(n8937), .B2(n7734), .ZN(n7736)
         );
  OAI211_X1 U9353 ( .C1(n10049), .C2(n8327), .A(n7737), .B(n7736), .ZN(
        P2_U3228) );
  INV_X1 U9354 ( .A(n7738), .ZN(n7740) );
  AOI21_X1 U9355 ( .B1(n7741), .B2(n7740), .A(n7739), .ZN(n7742) );
  MUX2_X1 U9356 ( .A(n6922), .B(n7742), .S(n9714), .Z(n7747) );
  NOR2_X1 U9357 ( .A1(n9711), .A2(n7743), .ZN(n7744) );
  AOI21_X1 U9358 ( .B1(n9642), .B2(n7745), .A(n7744), .ZN(n7746) );
  OAI211_X1 U9359 ( .C1(n9490), .C2(n7748), .A(n7747), .B(n7746), .ZN(P1_U3286) );
  OAI21_X1 U9360 ( .B1(n10080), .B2(n7750), .A(n7749), .ZN(n7756) );
  OAI22_X1 U9361 ( .A1(n7754), .A2(n9052), .B1(n10086), .B2(n6373), .ZN(n7751)
         );
  AOI21_X1 U9362 ( .B1(n7756), .B2(n10086), .A(n7751), .ZN(n7752) );
  INV_X1 U9363 ( .A(n7752), .ZN(P2_U3408) );
  INV_X1 U9364 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7753) );
  OAI22_X1 U9365 ( .A1(n8980), .A2(n7754), .B1(n10099), .B2(n7753), .ZN(n7755)
         );
  AOI21_X1 U9366 ( .B1(n7756), .B2(n10099), .A(n7755), .ZN(n7757) );
  INV_X1 U9367 ( .A(n7757), .ZN(P2_U3465) );
  INV_X1 U9368 ( .A(n7758), .ZN(n7762) );
  AOI211_X1 U9369 ( .C1(n7762), .C2(n7761), .A(n7760), .B(n7759), .ZN(n7768)
         );
  INV_X1 U9370 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7763) );
  OAI22_X1 U9371 ( .A1(n7764), .A2(n9864), .B1(n9860), .B2(n7763), .ZN(n7765)
         );
  INV_X1 U9372 ( .A(n7765), .ZN(n7766) );
  OAI21_X1 U9373 ( .B1(n7768), .B2(n6057), .A(n7766), .ZN(P1_U3477) );
  INV_X1 U9374 ( .A(n9823), .ZN(n7806) );
  AOI22_X1 U9375 ( .A1(n9921), .A2(n7806), .B1(n9985), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7767) );
  OAI21_X1 U9376 ( .B1(n7768), .B2(n9985), .A(n7767), .ZN(P1_U3530) );
  XNOR2_X1 U9377 ( .A(n7769), .B(n7776), .ZN(n7770) );
  NAND2_X1 U9378 ( .A1(n7770), .A2(n9724), .ZN(n7773) );
  NAND2_X1 U9379 ( .A1(n9296), .A2(n9728), .ZN(n7771) );
  OAI21_X1 U9380 ( .B1(n7985), .B2(n9662), .A(n7771), .ZN(n9901) );
  INV_X1 U9381 ( .A(n9901), .ZN(n7772) );
  NAND2_X1 U9382 ( .A1(n7773), .A2(n7772), .ZN(n7800) );
  INV_X1 U9383 ( .A(n7800), .ZN(n7785) );
  OAI21_X1 U9384 ( .B1(n7774), .B2(n7776), .A(n7775), .ZN(n7802) );
  NAND2_X1 U9385 ( .A1(n7802), .A2(n9707), .ZN(n7784) );
  INV_X1 U9386 ( .A(n7943), .ZN(n7779) );
  AOI21_X1 U9387 ( .B1(n7777), .B2(n9965), .A(n9904), .ZN(n7778) );
  NOR3_X1 U9388 ( .A1(n7779), .A2(n7778), .A3(n9969), .ZN(n7801) );
  NOR2_X1 U9389 ( .A1(n9904), .A2(n9945), .ZN(n7782) );
  OAI22_X1 U9390 ( .A1(n9714), .A2(n7780), .B1(n9909), .B2(n9711), .ZN(n7781)
         );
  AOI211_X1 U9391 ( .C1(n7801), .C2(n9950), .A(n7782), .B(n7781), .ZN(n7783)
         );
  OAI211_X1 U9392 ( .C1(n9612), .C2(n7785), .A(n7784), .B(n7783), .ZN(P1_U3283) );
  INV_X1 U9393 ( .A(n7786), .ZN(n7810) );
  OAI222_X1 U9394 ( .A1(n9117), .A2(n7810), .B1(P2_U3151), .B2(n7788), .C1(
        n7787), .C2(n9105), .ZN(P2_U3274) );
  XNOR2_X1 U9395 ( .A(n7789), .B(n7790), .ZN(n10054) );
  XNOR2_X1 U9396 ( .A(n7791), .B(n7790), .ZN(n7794) );
  OAI22_X1 U9397 ( .A1(n7792), .A2(n8930), .B1(n8135), .B2(n8928), .ZN(n7793)
         );
  AOI21_X1 U9398 ( .B1(n7794), .B2(n8914), .A(n7793), .ZN(n7795) );
  OAI21_X1 U9399 ( .B1(n8927), .B2(n10054), .A(n7795), .ZN(n10056) );
  NAND2_X1 U9400 ( .A1(n10056), .A2(n8942), .ZN(n7799) );
  OAI22_X1 U9401 ( .A1(n8942), .A2(n7796), .B1(n7865), .B2(n8899), .ZN(n7797)
         );
  AOI21_X1 U9402 ( .B1(n8890), .B2(n7860), .A(n7797), .ZN(n7798) );
  OAI211_X1 U9403 ( .C1(n10054), .C2(n8327), .A(n7799), .B(n7798), .ZN(
        P2_U3226) );
  AOI211_X1 U9404 ( .C1(n7802), .C2(n9979), .A(n7801), .B(n7800), .ZN(n7808)
         );
  INV_X1 U9405 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7803) );
  OAI22_X1 U9406 ( .A1(n9904), .A2(n9864), .B1(n9860), .B2(n7803), .ZN(n7804)
         );
  INV_X1 U9407 ( .A(n7804), .ZN(n7805) );
  OAI21_X1 U9408 ( .B1(n7808), .B2(n6057), .A(n7805), .ZN(P1_U3483) );
  AOI22_X1 U9409 ( .A1(n8109), .A2(n7806), .B1(n9985), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7807) );
  OAI21_X1 U9410 ( .B1(n7808), .B2(n9985), .A(n7807), .ZN(P1_U3532) );
  OAI222_X1 U9411 ( .A1(P1_U3086), .A2(n7811), .B1(n9884), .B2(n7810), .C1(
        n7809), .C2(n9882), .ZN(P1_U3334) );
  AOI21_X1 U9412 ( .B1(n6407), .B2(n7813), .A(n7867), .ZN(n7830) );
  MUX2_X1 U9413 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8699), .Z(n7815) );
  NOR2_X1 U9414 ( .A1(n7815), .A2(n7814), .ZN(n7883) );
  AND2_X1 U9415 ( .A1(n7815), .A2(n7814), .ZN(n7882) );
  NOR2_X1 U9416 ( .A1(n7883), .A2(n7882), .ZN(n7819) );
  OR2_X1 U9417 ( .A1(n7816), .A2(n7822), .ZN(n7818) );
  NAND2_X1 U9418 ( .A1(n7818), .A2(n7817), .ZN(n7884) );
  XNOR2_X1 U9419 ( .A(n7819), .B(n7884), .ZN(n7820) );
  NAND2_X1 U9420 ( .A1(n7820), .A2(n10020), .ZN(n7829) );
  XNOR2_X1 U9421 ( .A(n7873), .B(n7872), .ZN(n7823) );
  INV_X1 U9422 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7936) );
  NOR2_X1 U9423 ( .A1(n7936), .A2(n7823), .ZN(n7874) );
  AOI21_X1 U9424 ( .B1(n7823), .B2(n7936), .A(n7874), .ZN(n7825) );
  NOR2_X1 U9425 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10394), .ZN(n8128) );
  INV_X1 U9426 ( .A(n8128), .ZN(n7824) );
  OAI21_X1 U9427 ( .B1(n10026), .B2(n7825), .A(n7824), .ZN(n7827) );
  INV_X1 U9428 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10122) );
  NOR2_X1 U9429 ( .A1(n10011), .A2(n10122), .ZN(n7826) );
  AOI211_X1 U9430 ( .C1(n10014), .C2(n7873), .A(n7827), .B(n7826), .ZN(n7828)
         );
  OAI211_X1 U9431 ( .C1(n7830), .C2(n10022), .A(n7829), .B(n7828), .ZN(
        P2_U3191) );
  INV_X1 U9432 ( .A(n9433), .ZN(n7849) );
  OR2_X1 U9433 ( .A1(n9433), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U9434 ( .A1(n9433), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U9435 ( .A1(n9440), .A2(n7831), .ZN(n7835) );
  INV_X1 U9436 ( .A(n7835), .ZN(n7837) );
  AOI21_X1 U9437 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n7833), .A(n7832), .ZN(
        n7836) );
  INV_X1 U9438 ( .A(n7836), .ZN(n7834) );
  OAI21_X1 U9439 ( .B1(n7837), .B2(n7836), .A(n9441), .ZN(n7845) );
  INV_X1 U9440 ( .A(n9464), .ZN(n9439) );
  XNOR2_X1 U9441 ( .A(n9433), .B(n9809), .ZN(n7843) );
  AOI21_X1 U9442 ( .B1(n7840), .B2(n7839), .A(n7838), .ZN(n7841) );
  INV_X1 U9443 ( .A(n7841), .ZN(n7842) );
  NAND2_X1 U9444 ( .A1(n7843), .A2(n7842), .ZN(n9435) );
  OAI21_X1 U9445 ( .B1(n7843), .B2(n7842), .A(n9435), .ZN(n7844) );
  AOI22_X1 U9446 ( .A1(n9445), .A2(n7845), .B1(n9439), .B2(n7844), .ZN(n7848)
         );
  NAND2_X1 U9447 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9210) );
  INV_X1 U9448 ( .A(n9210), .ZN(n7846) );
  AOI21_X1 U9449 ( .B1(n9933), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n7846), .ZN(
        n7847) );
  OAI211_X1 U9450 ( .C1(n7849), .C2(n9459), .A(n7848), .B(n7847), .ZN(P1_U3260) );
  NAND2_X1 U9451 ( .A1(n7850), .A2(n8561), .ZN(n7851) );
  XNOR2_X1 U9452 ( .A(n10053), .B(n8198), .ZN(n7853) );
  NAND2_X1 U9453 ( .A1(n8560), .A2(n7853), .ZN(n7856) );
  INV_X1 U9454 ( .A(n7853), .ZN(n7855) );
  NAND2_X1 U9455 ( .A1(n7855), .A2(n7854), .ZN(n7964) );
  AND2_X1 U9456 ( .A1(n7856), .A2(n7964), .ZN(n7857) );
  OAI21_X1 U9457 ( .B1(n7858), .B2(n7857), .A(n7961), .ZN(n7859) );
  NAND2_X1 U9458 ( .A1(n7859), .A2(n8515), .ZN(n7864) );
  INV_X1 U9459 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10400) );
  NOR2_X1 U9460 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10400), .ZN(n10012) );
  AOI21_X1 U9461 ( .B1(n8534), .B2(n7860), .A(n10012), .ZN(n7861) );
  OAI21_X1 U9462 ( .B1(n8544), .B2(n8135), .A(n7861), .ZN(n7862) );
  AOI21_X1 U9463 ( .B1(n8548), .B2(n8561), .A(n7862), .ZN(n7863) );
  OAI211_X1 U9464 ( .C1(n7865), .C2(n8545), .A(n7864), .B(n7863), .ZN(P2_U3153) );
  NOR2_X1 U9465 ( .A1(n7873), .A2(n7866), .ZN(n7868) );
  NAND2_X1 U9466 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n8072), .ZN(n7869) );
  OAI21_X1 U9467 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n8072), .A(n7869), .ZN(
        n7870) );
  AOI21_X1 U9468 ( .B1(n4591), .B2(n7870), .A(n8071), .ZN(n7894) );
  INV_X1 U9469 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10126) );
  INV_X1 U9470 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10494) );
  NOR2_X1 U9471 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10494), .ZN(n8186) );
  INV_X1 U9472 ( .A(n8186), .ZN(n7871) );
  OAI21_X1 U9473 ( .B1(n10011), .B2(n10126), .A(n7871), .ZN(n7881) );
  NOR2_X1 U9474 ( .A1(n7873), .A2(n7872), .ZN(n7875) );
  NAND2_X1 U9475 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n8072), .ZN(n7876) );
  OAI21_X1 U9476 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n8072), .A(n7876), .ZN(
        n7877) );
  NOR2_X1 U9477 ( .A1(n7878), .A2(n7877), .ZN(n8051) );
  AOI21_X1 U9478 ( .B1(n7878), .B2(n7877), .A(n8051), .ZN(n7879) );
  NOR2_X1 U9479 ( .A1(n7879), .A2(n10026), .ZN(n7880) );
  AOI211_X1 U9480 ( .C1(n10014), .C2(n7888), .A(n7881), .B(n7880), .ZN(n7893)
         );
  INV_X1 U9481 ( .A(n7882), .ZN(n7885) );
  MUX2_X1 U9482 ( .A(n6421), .B(n6420), .S(n8699), .Z(n7887) );
  AND2_X1 U9483 ( .A1(n7887), .A2(n7888), .ZN(n8060) );
  INV_X1 U9484 ( .A(n8060), .ZN(n7886) );
  OAI21_X1 U9485 ( .B1(n7888), .B2(n7887), .A(n7886), .ZN(n7889) );
  AOI21_X1 U9486 ( .B1(n7890), .B2(n7889), .A(n8059), .ZN(n7891) );
  OR2_X1 U9487 ( .A1(n7891), .A2(n8707), .ZN(n7892) );
  OAI211_X1 U9488 ( .C1(n7894), .C2(n10022), .A(n7893), .B(n7892), .ZN(
        P2_U3192) );
  XNOR2_X1 U9489 ( .A(n7895), .B(n7897), .ZN(n10060) );
  XNOR2_X1 U9490 ( .A(n7896), .B(n7897), .ZN(n7898) );
  AOI222_X1 U9491 ( .A1(n8914), .A2(n7898), .B1(n8558), .B2(n8909), .C1(n8560), 
        .C2(n8911), .ZN(n10058) );
  MUX2_X1 U9492 ( .A(n7899), .B(n10058), .S(n8942), .Z(n7902) );
  INV_X1 U9493 ( .A(n7960), .ZN(n7900) );
  AOI22_X1 U9494 ( .A1(n8890), .A2(n7969), .B1(n8937), .B2(n7900), .ZN(n7901)
         );
  OAI211_X1 U9495 ( .C1(n10060), .C2(n8923), .A(n7902), .B(n7901), .ZN(
        P2_U3225) );
  XOR2_X1 U9496 ( .A(n7903), .B(n7904), .Z(n9973) );
  INV_X1 U9497 ( .A(n9973), .ZN(n7917) );
  NAND2_X1 U9498 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  NAND2_X1 U9499 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  NAND2_X1 U9500 ( .A1(n7908), .A2(n9724), .ZN(n7910) );
  AOI22_X1 U9501 ( .A1(n9727), .A2(n9296), .B1(n9294), .B2(n9728), .ZN(n7909)
         );
  NAND2_X1 U9502 ( .A1(n7910), .A2(n7909), .ZN(n9972) );
  NAND2_X1 U9503 ( .A1(n7941), .A2(n8221), .ZN(n7911) );
  NAND2_X1 U9504 ( .A1(n4589), .A2(n7911), .ZN(n9970) );
  NAND2_X1 U9505 ( .A1(n9612), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7912) );
  OAI21_X1 U9506 ( .B1(n9711), .B2(n9178), .A(n7912), .ZN(n7913) );
  AOI21_X1 U9507 ( .B1(n8221), .B2(n9642), .A(n7913), .ZN(n7914) );
  OAI21_X1 U9508 ( .B1(n9970), .B2(n9490), .A(n7914), .ZN(n7915) );
  AOI21_X1 U9509 ( .B1(n9972), .B2(n9714), .A(n7915), .ZN(n7916) );
  OAI21_X1 U9510 ( .B1(n7917), .B2(n9741), .A(n7916), .ZN(P1_U3281) );
  INV_X1 U9511 ( .A(n7918), .ZN(n7922) );
  INV_X1 U9512 ( .A(n7919), .ZN(n7920) );
  OAI222_X1 U9513 ( .A1(n9122), .A2(n7921), .B1(n9117), .B2(n7922), .C1(n7920), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9514 ( .A1(n7923), .A2(P1_U3086), .B1(n9884), .B2(n7922), .C1(
        n10278), .C2(n9882), .ZN(P1_U3333) );
  NAND2_X1 U9515 ( .A1(n7927), .A2(n7924), .ZN(n7926) );
  OAI211_X1 U9516 ( .C1(n10300), .C2(n9882), .A(n7926), .B(n7925), .ZN(
        P1_U3332) );
  NAND2_X1 U9517 ( .A1(n7927), .A2(n9109), .ZN(n7929) );
  OAI211_X1 U9518 ( .C1(n7930), .C2(n9105), .A(n7929), .B(n7928), .ZN(P2_U3272) );
  XNOR2_X1 U9519 ( .A(n7931), .B(n7932), .ZN(n10064) );
  OAI21_X1 U9520 ( .B1(n4592), .B2(n7932), .A(n5146), .ZN(n7934) );
  OAI22_X1 U9521 ( .A1(n8135), .A2(n8930), .B1(n8196), .B2(n8928), .ZN(n7933)
         );
  AOI21_X1 U9522 ( .B1(n7934), .B2(n8914), .A(n7933), .ZN(n7935) );
  OAI21_X1 U9523 ( .B1(n8927), .B2(n10064), .A(n7935), .ZN(n10065) );
  NAND2_X1 U9524 ( .A1(n10065), .A2(n8942), .ZN(n7939) );
  OAI22_X1 U9525 ( .A1(n8942), .A2(n7936), .B1(n8129), .B2(n8899), .ZN(n7937)
         );
  AOI21_X1 U9526 ( .B1(n8890), .B2(n10067), .A(n7937), .ZN(n7938) );
  OAI211_X1 U9527 ( .C1(n10064), .C2(n8327), .A(n7939), .B(n7938), .ZN(
        P2_U3224) );
  XOR2_X1 U9528 ( .A(n7940), .B(n7951), .Z(n8008) );
  INV_X1 U9529 ( .A(n7941), .ZN(n7942) );
  AOI21_X1 U9530 ( .B1(n8115), .B2(n7943), .A(n7942), .ZN(n8005) );
  INV_X1 U9531 ( .A(n9490), .ZN(n9717) );
  INV_X1 U9532 ( .A(n7944), .ZN(n8125) );
  AOI22_X1 U9533 ( .A1(n9612), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8125), .B2(
        n9942), .ZN(n7945) );
  OAI21_X1 U9534 ( .B1(n4715), .B2(n9945), .A(n7945), .ZN(n7955) );
  NOR2_X1 U9535 ( .A1(n8123), .A2(n9662), .ZN(n7953) );
  NAND2_X1 U9536 ( .A1(n7947), .A2(n7946), .ZN(n7950) );
  INV_X1 U9537 ( .A(n7948), .ZN(n7949) );
  AOI211_X1 U9538 ( .C1(n7951), .C2(n7950), .A(n9659), .B(n7949), .ZN(n7952)
         );
  AOI211_X1 U9539 ( .C1(n9728), .C2(n9295), .A(n7953), .B(n7952), .ZN(n8007)
         );
  NOR2_X1 U9540 ( .A1(n8007), .A2(n9612), .ZN(n7954) );
  AOI211_X1 U9541 ( .C1(n8005), .C2(n9717), .A(n7955), .B(n7954), .ZN(n7956)
         );
  OAI21_X1 U9542 ( .B1(n8008), .B2(n9741), .A(n7956), .ZN(P1_U3282) );
  NOR2_X1 U9543 ( .A1(n8544), .A2(n8133), .ZN(n7957) );
  AOI211_X1 U9544 ( .C1(n8548), .C2(n8560), .A(n7958), .B(n7957), .ZN(n7959)
         );
  OAI21_X1 U9545 ( .B1(n7960), .B2(n8545), .A(n7959), .ZN(n7968) );
  NAND2_X1 U9546 ( .A1(n7961), .A2(n7964), .ZN(n7962) );
  XNOR2_X1 U9547 ( .A(n10059), .B(n8198), .ZN(n8134) );
  XNOR2_X1 U9548 ( .A(n8134), .B(n8135), .ZN(n7963) );
  NAND2_X1 U9549 ( .A1(n7962), .A2(n7963), .ZN(n8138) );
  INV_X1 U9550 ( .A(n7963), .ZN(n7965) );
  NAND3_X1 U9551 ( .A1(n7961), .A2(n7965), .A3(n7964), .ZN(n7966) );
  AOI21_X1 U9552 ( .B1(n8138), .B2(n7966), .A(n8538), .ZN(n7967) );
  AOI211_X1 U9553 ( .C1(n7969), .C2(n8534), .A(n7968), .B(n7967), .ZN(n7970)
         );
  INV_X1 U9554 ( .A(n7970), .ZN(P2_U3161) );
  NAND2_X1 U9555 ( .A1(n9921), .A2(n8233), .ZN(n7972) );
  NAND2_X1 U9556 ( .A1(n9299), .A2(n9148), .ZN(n7971) );
  NAND2_X1 U9557 ( .A1(n7972), .A2(n7971), .ZN(n7973) );
  XNOR2_X1 U9558 ( .A(n7973), .B(n8277), .ZN(n7988) );
  INV_X1 U9559 ( .A(n7988), .ZN(n7981) );
  INV_X1 U9560 ( .A(n7974), .ZN(n7977) );
  INV_X1 U9561 ( .A(n7975), .ZN(n7976) );
  NAND2_X1 U9562 ( .A1(n7977), .A2(n7976), .ZN(n7990) );
  NAND2_X1 U9563 ( .A1(n7995), .A2(n7990), .ZN(n7980) );
  XOR2_X1 U9564 ( .A(n7988), .B(n7980), .Z(n9915) );
  NAND2_X1 U9565 ( .A1(n9921), .A2(n8306), .ZN(n7979) );
  NAND2_X1 U9566 ( .A1(n9299), .A2(n9149), .ZN(n7978) );
  NAND2_X1 U9567 ( .A1(n7979), .A2(n7978), .ZN(n9914) );
  NOR2_X1 U9568 ( .A1(n9915), .A2(n9914), .ZN(n9913) );
  AOI21_X1 U9569 ( .B1(n7981), .B2(n7980), .A(n9913), .ZN(n7997) );
  NAND2_X1 U9570 ( .A1(n7987), .A2(n8233), .ZN(n7983) );
  NAND2_X1 U9571 ( .A1(n9298), .A2(n9148), .ZN(n7982) );
  NAND2_X1 U9572 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  XNOR2_X1 U9573 ( .A(n7984), .B(n8277), .ZN(n8100) );
  NOR2_X1 U9574 ( .A1(n7985), .A2(n8310), .ZN(n7986) );
  AOI21_X1 U9575 ( .B1(n7987), .B2(n8306), .A(n7986), .ZN(n8101) );
  XNOR2_X1 U9576 ( .A(n8100), .B(n8101), .ZN(n7996) );
  AOI21_X1 U9577 ( .B1(n9914), .B2(n7990), .A(n7988), .ZN(n7989) );
  INV_X1 U9578 ( .A(n7989), .ZN(n7994) );
  INV_X1 U9579 ( .A(n7990), .ZN(n7992) );
  INV_X1 U9580 ( .A(n9914), .ZN(n7991) );
  NAND2_X1 U9581 ( .A1(n7992), .A2(n7991), .ZN(n7993) );
  OAI211_X1 U9582 ( .C1(n7997), .C2(n7996), .A(n9906), .B(n8104), .ZN(n8004)
         );
  INV_X1 U9583 ( .A(n7998), .ZN(n8002) );
  OAI22_X1 U9584 ( .A1(n7999), .A2(n9279), .B1(n9890), .B2(n8123), .ZN(n8000)
         );
  AOI211_X1 U9585 ( .C1(n9269), .C2(n8002), .A(n8001), .B(n8000), .ZN(n8003)
         );
  OAI211_X1 U9586 ( .C1(n9965), .C2(n9903), .A(n8004), .B(n8003), .ZN(P1_U3231) );
  INV_X1 U9587 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8010) );
  AOI22_X1 U9588 ( .A1(n8005), .A2(n9813), .B1(n9956), .B2(n8115), .ZN(n8006)
         );
  OAI211_X1 U9589 ( .C1(n8008), .C2(n9804), .A(n8007), .B(n8006), .ZN(n8011)
         );
  NAND2_X1 U9590 ( .A1(n8011), .A2(n9860), .ZN(n8009) );
  OAI21_X1 U9591 ( .B1(n9860), .B2(n8010), .A(n8009), .ZN(P1_U3486) );
  NAND2_X1 U9592 ( .A1(n8011), .A2(n9988), .ZN(n8012) );
  OAI21_X1 U9593 ( .B1(n9988), .B2(n6956), .A(n8012), .ZN(P1_U3533) );
  XOR2_X1 U9594 ( .A(n8014), .B(n8013), .Z(n8164) );
  INV_X1 U9595 ( .A(n8164), .ZN(n8024) );
  INV_X1 U9596 ( .A(n8014), .ZN(n8015) );
  XNOR2_X1 U9597 ( .A(n8016), .B(n8015), .ZN(n8017) );
  NAND2_X1 U9598 ( .A1(n8017), .A2(n9724), .ZN(n8019) );
  AOI22_X1 U9599 ( .A1(n9728), .A2(n9726), .B1(n9295), .B2(n9727), .ZN(n8018)
         );
  NAND2_X1 U9600 ( .A1(n8019), .A2(n8018), .ZN(n8162) );
  AOI211_X1 U9601 ( .C1(n8212), .C2(n4589), .A(n9969), .B(n8155), .ZN(n8163)
         );
  NAND2_X1 U9602 ( .A1(n8163), .A2(n9950), .ZN(n8021) );
  AOI22_X1 U9603 ( .A1(n9612), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9237), .B2(
        n9942), .ZN(n8020) );
  OAI211_X1 U9604 ( .C1(n9240), .C2(n9945), .A(n8021), .B(n8020), .ZN(n8022)
         );
  AOI21_X1 U9605 ( .B1(n9714), .B2(n8162), .A(n8022), .ZN(n8023) );
  OAI21_X1 U9606 ( .B1(n8024), .B2(n9741), .A(n8023), .ZN(P1_U3280) );
  INV_X1 U9607 ( .A(n8025), .ZN(n8049) );
  OAI222_X1 U9608 ( .A1(n9117), .A2(n8049), .B1(P2_U3151), .B2(n6749), .C1(
        n8026), .C2(n9105), .ZN(P2_U3271) );
  INV_X1 U9609 ( .A(n8029), .ZN(n8027) );
  XNOR2_X1 U9610 ( .A(n8028), .B(n8027), .ZN(n10068) );
  XNOR2_X1 U9611 ( .A(n8030), .B(n8029), .ZN(n8032) );
  OAI22_X1 U9612 ( .A1(n8133), .A2(n8930), .B1(n8191), .B2(n8928), .ZN(n8031)
         );
  AOI21_X1 U9613 ( .B1(n8032), .B2(n8914), .A(n8031), .ZN(n8033) );
  OAI21_X1 U9614 ( .B1(n10068), .B2(n8927), .A(n8033), .ZN(n10069) );
  NAND2_X1 U9615 ( .A1(n10069), .A2(n8942), .ZN(n8036) );
  OAI22_X1 U9616 ( .A1(n8942), .A2(n6421), .B1(n8187), .B2(n8899), .ZN(n8034)
         );
  AOI21_X1 U9617 ( .B1(n8890), .B2(n10071), .A(n8034), .ZN(n8035) );
  OAI211_X1 U9618 ( .C1(n10068), .C2(n8327), .A(n8036), .B(n8035), .ZN(
        P2_U3223) );
  NAND2_X1 U9619 ( .A1(n8037), .A2(n8199), .ZN(n8038) );
  NAND3_X1 U9620 ( .A1(n8039), .A2(n8914), .A3(n8038), .ZN(n8041) );
  AOI22_X1 U9621 ( .A1(n8557), .A2(n8911), .B1(n8909), .B2(n8912), .ZN(n8040)
         );
  NAND2_X1 U9622 ( .A1(n8041), .A2(n8040), .ZN(n10075) );
  INV_X1 U9623 ( .A(n10075), .ZN(n8048) );
  OAI21_X1 U9624 ( .B1(n8043), .B2(n8199), .A(n8042), .ZN(n10077) );
  INV_X1 U9625 ( .A(n8923), .ZN(n8822) );
  INV_X1 U9626 ( .A(n8208), .ZN(n10074) );
  INV_X1 U9627 ( .A(n8044), .ZN(n8203) );
  AOI22_X1 U9628 ( .A1(n8920), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8937), .B2(
        n8203), .ZN(n8045) );
  OAI21_X1 U9629 ( .B1(n10074), .B2(n8820), .A(n8045), .ZN(n8046) );
  AOI21_X1 U9630 ( .B1(n10077), .B2(n8822), .A(n8046), .ZN(n8047) );
  OAI21_X1 U9631 ( .B1(n8048), .B2(n8920), .A(n8047), .ZN(P2_U3222) );
  OAI222_X1 U9632 ( .A1(n8050), .A2(P1_U3086), .B1(n9884), .B2(n8049), .C1(
        n10495), .C2(n9882), .ZN(P1_U3331) );
  NOR2_X1 U9633 ( .A1(n8097), .A2(n8052), .ZN(n8053) );
  INV_X1 U9634 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8054) );
  MUX2_X1 U9635 ( .A(n8054), .B(P2_REG2_REG_12__SCAN_IN), .S(n8080), .Z(n8055)
         );
  INV_X1 U9636 ( .A(n8055), .ZN(n8056) );
  AOI21_X1 U9637 ( .B1(n4582), .B2(n8056), .A(n8569), .ZN(n8083) );
  MUX2_X1 U9638 ( .A(n8058), .B(n8057), .S(n8699), .Z(n8061) );
  AND2_X1 U9639 ( .A1(n8061), .A2(n8097), .ZN(n8065) );
  INV_X1 U9640 ( .A(n8061), .ZN(n8063) );
  AND2_X1 U9641 ( .A1(n8063), .A2(n8062), .ZN(n8064) );
  OR2_X1 U9642 ( .A1(n8065), .A2(n8064), .ZN(n8088) );
  MUX2_X1 U9643 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8699), .Z(n8066) );
  AND2_X1 U9644 ( .A1(n8066), .A2(n8570), .ZN(n8577) );
  INV_X1 U9645 ( .A(n8577), .ZN(n8069) );
  MUX2_X1 U9646 ( .A(n8054), .B(n8067), .S(n8699), .Z(n8068) );
  NAND2_X1 U9647 ( .A1(n8068), .A2(n8080), .ZN(n8578) );
  NAND2_X1 U9648 ( .A1(n8069), .A2(n8578), .ZN(n8070) );
  XNOR2_X1 U9649 ( .A(n8579), .B(n8070), .ZN(n8078) );
  NOR2_X1 U9650 ( .A1(n8097), .A2(n8073), .ZN(n8074) );
  AOI22_X1 U9651 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8080), .B1(n8570), .B2(
        n8067), .ZN(n8075) );
  AOI21_X1 U9652 ( .B1(n4585), .B2(n8075), .A(n8567), .ZN(n8076) );
  NOR2_X1 U9653 ( .A1(n8076), .A2(n10022), .ZN(n8077) );
  AOI21_X1 U9654 ( .B1(n8078), .B2(n10020), .A(n8077), .ZN(n8082) );
  INV_X1 U9655 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10345) );
  NOR2_X1 U9656 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10345), .ZN(n8441) );
  INV_X1 U9657 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10134) );
  NOR2_X1 U9658 ( .A1(n10011), .A2(n10134), .ZN(n8079) );
  AOI211_X1 U9659 ( .C1(n10014), .C2(n8080), .A(n8441), .B(n8079), .ZN(n8081)
         );
  OAI211_X1 U9660 ( .C1(n8083), .C2(n10026), .A(n8082), .B(n8081), .ZN(
        P2_U3194) );
  AOI21_X1 U9661 ( .B1(n8057), .B2(n8085), .A(n8084), .ZN(n8099) );
  AOI21_X1 U9662 ( .B1(n8088), .B2(n8087), .A(n8086), .ZN(n8091) );
  INV_X1 U9663 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10130) );
  OR2_X1 U9664 ( .A1(n10011), .A2(n10130), .ZN(n8090) );
  INV_X1 U9665 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10523) );
  NOR2_X1 U9666 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10523), .ZN(n8202) );
  INV_X1 U9667 ( .A(n8202), .ZN(n8089) );
  OAI211_X1 U9668 ( .C1(n8091), .C2(n8707), .A(n8090), .B(n8089), .ZN(n8096)
         );
  AOI21_X1 U9669 ( .B1(n8058), .B2(n8093), .A(n8092), .ZN(n8094) );
  NOR2_X1 U9670 ( .A1(n8094), .A2(n10026), .ZN(n8095) );
  AOI211_X1 U9671 ( .C1(n10014), .C2(n8097), .A(n8096), .B(n8095), .ZN(n8098)
         );
  OAI21_X1 U9672 ( .B1(n8099), .B2(n10022), .A(n8098), .ZN(P2_U3193) );
  AOI22_X1 U9673 ( .A1(n8109), .A2(n8233), .B1(n9148), .B2(n9297), .ZN(n8105)
         );
  XOR2_X1 U9674 ( .A(n8277), .B(n8105), .Z(n8106) );
  NOR2_X1 U9675 ( .A1(n8110), .A2(n8108), .ZN(n9897) );
  AOI22_X1 U9676 ( .A1(n8109), .A2(n8306), .B1(n9149), .B2(n9297), .ZN(n9898)
         );
  NAND2_X1 U9677 ( .A1(n8115), .A2(n8233), .ZN(n8112) );
  NAND2_X1 U9678 ( .A1(n9296), .A2(n8306), .ZN(n8111) );
  NAND2_X1 U9679 ( .A1(n8112), .A2(n8111), .ZN(n8113) );
  XNOR2_X1 U9680 ( .A(n8113), .B(n9152), .ZN(n8116) );
  AND2_X1 U9681 ( .A1(n9296), .A2(n9149), .ZN(n8114) );
  AOI21_X1 U9682 ( .B1(n8115), .B2(n9148), .A(n8114), .ZN(n8117) );
  NAND2_X1 U9683 ( .A1(n8116), .A2(n8117), .ZN(n8216) );
  INV_X1 U9684 ( .A(n8116), .ZN(n8119) );
  INV_X1 U9685 ( .A(n8117), .ZN(n8118) );
  NAND2_X1 U9686 ( .A1(n8119), .A2(n8118), .ZN(n8120) );
  NAND2_X1 U9687 ( .A1(n8216), .A2(n8120), .ZN(n8121) );
  OAI21_X1 U9688 ( .B1(n4581), .B2(n8122), .A(n9906), .ZN(n8127) );
  AND2_X1 U9689 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9393) );
  OAI22_X1 U9690 ( .A1(n8123), .A2(n9279), .B1(n9890), .B2(n6023), .ZN(n8124)
         );
  AOI211_X1 U9691 ( .C1(n8125), .C2(n9269), .A(n9393), .B(n8124), .ZN(n8126)
         );
  OAI211_X1 U9692 ( .C1(n4715), .C2(n9903), .A(n8127), .B(n8126), .ZN(P1_U3236) );
  AOI21_X1 U9693 ( .B1(n8548), .B2(n8559), .A(n8128), .ZN(n8132) );
  INV_X1 U9694 ( .A(n8129), .ZN(n8130) );
  NAND2_X1 U9695 ( .A1(n8533), .A2(n8130), .ZN(n8131) );
  OAI211_X1 U9696 ( .C1(n8196), .C2(n8544), .A(n8132), .B(n8131), .ZN(n8144)
         );
  XNOR2_X1 U9697 ( .A(n10067), .B(n8198), .ZN(n8179) );
  XNOR2_X1 U9698 ( .A(n8179), .B(n8133), .ZN(n8142) );
  INV_X1 U9699 ( .A(n8134), .ZN(n8136) );
  NAND2_X1 U9700 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  INV_X1 U9701 ( .A(n8182), .ZN(n8140) );
  AOI211_X1 U9702 ( .C1(n8142), .C2(n8141), .A(n8538), .B(n8140), .ZN(n8143)
         );
  AOI211_X1 U9703 ( .C1(n10067), .C2(n8534), .A(n8144), .B(n8143), .ZN(n8145)
         );
  INV_X1 U9704 ( .A(n8145), .ZN(P2_U3171) );
  XNOR2_X1 U9705 ( .A(n8146), .B(n4874), .ZN(n9980) );
  INV_X1 U9706 ( .A(n9980), .ZN(n8161) );
  NAND2_X1 U9707 ( .A1(n8148), .A2(n8147), .ZN(n8149) );
  NAND2_X1 U9708 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  NAND2_X1 U9709 ( .A1(n8151), .A2(n9724), .ZN(n8153) );
  AOI22_X1 U9710 ( .A1(n9727), .A2(n9294), .B1(n9701), .B2(n9728), .ZN(n8152)
         );
  NAND2_X1 U9711 ( .A1(n8153), .A2(n8152), .ZN(n9978) );
  INV_X1 U9712 ( .A(n8154), .ZN(n9733) );
  OAI211_X1 U9713 ( .C1(n9976), .C2(n8155), .A(n9733), .B(n9813), .ZN(n9975)
         );
  INV_X1 U9714 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8156) );
  OAI22_X1 U9715 ( .A1(n9714), .A2(n8156), .B1(n9131), .B2(n9711), .ZN(n8157)
         );
  AOI21_X1 U9716 ( .B1(n9134), .B2(n9642), .A(n8157), .ZN(n8158) );
  OAI21_X1 U9717 ( .B1(n9975), .B2(n9646), .A(n8158), .ZN(n8159) );
  AOI21_X1 U9718 ( .B1(n9978), .B2(n9714), .A(n8159), .ZN(n8160) );
  OAI21_X1 U9719 ( .B1(n8161), .B2(n9741), .A(n8160), .ZN(P1_U3279) );
  AOI211_X1 U9720 ( .C1(n8164), .C2(n9979), .A(n8163), .B(n8162), .ZN(n8167)
         );
  MUX2_X1 U9721 ( .A(n8165), .B(n8167), .S(n9988), .Z(n8166) );
  OAI21_X1 U9722 ( .B1(n9240), .B2(n9823), .A(n8166), .ZN(P1_U3535) );
  INV_X1 U9723 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8168) );
  MUX2_X1 U9724 ( .A(n8168), .B(n8167), .S(n9860), .Z(n8169) );
  OAI21_X1 U9725 ( .B1(n9240), .B2(n9864), .A(n8169), .ZN(P1_U3492) );
  OAI21_X1 U9726 ( .B1(n8172), .B2(n8171), .A(n8170), .ZN(n10081) );
  INV_X1 U9727 ( .A(n8914), .ZN(n8932) );
  XNOR2_X1 U9728 ( .A(n8173), .B(n8174), .ZN(n8175) );
  OAI222_X1 U9729 ( .A1(n8928), .A2(n8439), .B1(n8930), .B2(n8191), .C1(n8932), 
        .C2(n8175), .ZN(n10082) );
  NAND2_X1 U9730 ( .A1(n10082), .A2(n8942), .ZN(n8178) );
  OAI22_X1 U9731 ( .A1(n8942), .A2(n8054), .B1(n8443), .B2(n8899), .ZN(n8176)
         );
  AOI21_X1 U9732 ( .B1(n10084), .B2(n8890), .A(n8176), .ZN(n8177) );
  OAI211_X1 U9733 ( .C1(n8923), .C2(n10081), .A(n8178), .B(n8177), .ZN(
        P2_U3221) );
  INV_X1 U9734 ( .A(n8179), .ZN(n8180) );
  NAND2_X1 U9735 ( .A1(n8180), .A2(n8558), .ZN(n8181) );
  XNOR2_X1 U9736 ( .A(n10071), .B(n8198), .ZN(n8183) );
  OAI21_X1 U9737 ( .B1(n8184), .B2(n8183), .A(n8200), .ZN(n8185) );
  NAND2_X1 U9738 ( .A1(n8185), .A2(n8515), .ZN(n8194) );
  AOI21_X1 U9739 ( .B1(n8548), .B2(n8558), .A(n8186), .ZN(n8190) );
  INV_X1 U9740 ( .A(n8187), .ZN(n8188) );
  NAND2_X1 U9741 ( .A1(n8533), .A2(n8188), .ZN(n8189) );
  OAI211_X1 U9742 ( .C1(n8191), .C2(n8544), .A(n8190), .B(n8189), .ZN(n8192)
         );
  AOI21_X1 U9743 ( .B1(n10071), .B2(n8534), .A(n8192), .ZN(n8193) );
  NAND2_X1 U9744 ( .A1(n8194), .A2(n8193), .ZN(P2_U3157) );
  INV_X1 U9745 ( .A(n8195), .ZN(n8197) );
  NAND2_X1 U9746 ( .A1(n8197), .A2(n8196), .ZN(n8201) );
  XNOR2_X1 U9747 ( .A(n8199), .B(n8198), .ZN(n8347) );
  NAND2_X1 U9748 ( .A1(n8350), .A2(n8515), .ZN(n8211) );
  AOI21_X1 U9749 ( .B1(n8200), .B2(n8201), .A(n8347), .ZN(n8210) );
  AOI21_X1 U9750 ( .B1(n8548), .B2(n8557), .A(n8202), .ZN(n8205) );
  NAND2_X1 U9751 ( .A1(n8533), .A2(n8203), .ZN(n8204) );
  OAI211_X1 U9752 ( .C1(n8206), .C2(n8544), .A(n8205), .B(n8204), .ZN(n8207)
         );
  AOI21_X1 U9753 ( .B1(n8208), .B2(n8534), .A(n8207), .ZN(n8209) );
  OAI21_X1 U9754 ( .B1(n8211), .B2(n8210), .A(n8209), .ZN(P2_U3176) );
  OAI22_X1 U9755 ( .A1(n9240), .A2(n8284), .B1(n9179), .B2(n8310), .ZN(n8229)
         );
  NAND2_X1 U9756 ( .A1(n8212), .A2(n8233), .ZN(n8214) );
  NAND2_X1 U9757 ( .A1(n9294), .A2(n8306), .ZN(n8213) );
  NAND2_X1 U9758 ( .A1(n8214), .A2(n8213), .ZN(n8215) );
  XNOR2_X1 U9759 ( .A(n8215), .B(n8277), .ZN(n8228) );
  INV_X1 U9760 ( .A(n8216), .ZN(n9175) );
  NAND2_X1 U9761 ( .A1(n8221), .A2(n8233), .ZN(n8218) );
  NAND2_X1 U9762 ( .A1(n9295), .A2(n8306), .ZN(n8217) );
  NAND2_X1 U9763 ( .A1(n8218), .A2(n8217), .ZN(n8219) );
  XNOR2_X1 U9764 ( .A(n8219), .B(n9152), .ZN(n8222) );
  AND2_X1 U9765 ( .A1(n9295), .A2(n9149), .ZN(n8220) );
  AOI21_X1 U9766 ( .B1(n8221), .B2(n8306), .A(n8220), .ZN(n8223) );
  NAND2_X1 U9767 ( .A1(n8222), .A2(n8223), .ZN(n8227) );
  INV_X1 U9768 ( .A(n8222), .ZN(n8225) );
  INV_X1 U9769 ( .A(n8223), .ZN(n8224) );
  NAND2_X1 U9770 ( .A1(n8225), .A2(n8224), .ZN(n8226) );
  AND2_X1 U9771 ( .A1(n8227), .A2(n8226), .ZN(n9174) );
  XOR2_X1 U9772 ( .A(n8229), .B(n8228), .Z(n9234) );
  AOI22_X1 U9773 ( .A1(n9134), .A2(n8233), .B1(n9148), .B2(n9726), .ZN(n8230)
         );
  XNOR2_X1 U9774 ( .A(n8230), .B(n8277), .ZN(n8232) );
  OAI22_X1 U9775 ( .A1(n9976), .A2(n8284), .B1(n9280), .B2(n8310), .ZN(n9129)
         );
  NAND2_X1 U9776 ( .A1(n9734), .A2(n8233), .ZN(n8235) );
  NAND2_X1 U9777 ( .A1(n9701), .A2(n8306), .ZN(n8234) );
  NAND2_X1 U9778 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  XNOR2_X1 U9779 ( .A(n8236), .B(n9152), .ZN(n8237) );
  OAI22_X1 U9780 ( .A1(n9865), .A2(n8284), .B1(n9199), .B2(n8310), .ZN(n9275)
         );
  NAND3_X1 U9781 ( .A1(n8238), .A2(n8237), .A3(n9127), .ZN(n9272) );
  OAI21_X1 U9782 ( .B1(n9273), .B2(n9275), .A(n9272), .ZN(n9197) );
  NAND2_X1 U9783 ( .A1(n9812), .A2(n8233), .ZN(n8240) );
  NAND2_X1 U9784 ( .A1(n4793), .A2(n8306), .ZN(n8239) );
  NAND2_X1 U9785 ( .A1(n8240), .A2(n8239), .ZN(n8241) );
  XNOR2_X1 U9786 ( .A(n8241), .B(n9152), .ZN(n8244) );
  NOR2_X1 U9787 ( .A1(n9278), .A2(n8310), .ZN(n8242) );
  AOI21_X1 U9788 ( .B1(n9812), .B2(n9148), .A(n8242), .ZN(n8243) );
  OR2_X1 U9789 ( .A1(n8244), .A2(n8243), .ZN(n9195) );
  NAND2_X1 U9790 ( .A1(n9197), .A2(n9195), .ZN(n8245) );
  NAND2_X1 U9791 ( .A1(n8244), .A2(n8243), .ZN(n9194) );
  NAND2_X1 U9792 ( .A1(n8245), .A2(n9194), .ZN(n9204) );
  OAI22_X1 U9793 ( .A1(n9858), .A2(n8293), .B1(n9256), .B2(n8284), .ZN(n8246)
         );
  XNOR2_X1 U9794 ( .A(n8246), .B(n8277), .ZN(n8249) );
  OR2_X1 U9795 ( .A1(n9858), .A2(n8284), .ZN(n8248) );
  NAND2_X1 U9796 ( .A1(n9702), .A2(n9149), .ZN(n8247) );
  NAND2_X1 U9797 ( .A1(n8248), .A2(n8247), .ZN(n8250) );
  NAND2_X1 U9798 ( .A1(n8249), .A2(n8250), .ZN(n9205) );
  INV_X1 U9799 ( .A(n8249), .ZN(n8252) );
  INV_X1 U9800 ( .A(n8250), .ZN(n8251) );
  NAND2_X1 U9801 ( .A1(n8252), .A2(n8251), .ZN(n9206) );
  AOI22_X1 U9802 ( .A1(n4719), .A2(n8233), .B1(n9148), .B2(n9293), .ZN(n8253)
         );
  XNOR2_X1 U9803 ( .A(n8253), .B(n8277), .ZN(n8255) );
  AOI22_X1 U9804 ( .A1(n4719), .A2(n8306), .B1(n9149), .B2(n9293), .ZN(n9253)
         );
  OAI22_X1 U9805 ( .A1(n9652), .A2(n8293), .B1(n9292), .B2(n8284), .ZN(n8257)
         );
  XNOR2_X1 U9806 ( .A(n8257), .B(n8277), .ZN(n8259) );
  OAI22_X1 U9807 ( .A1(n9652), .A2(n8284), .B1(n9292), .B2(n8310), .ZN(n8258)
         );
  XNOR2_X1 U9808 ( .A(n8259), .B(n8258), .ZN(n9143) );
  NAND2_X1 U9809 ( .A1(n8259), .A2(n8258), .ZN(n8260) );
  NAND2_X1 U9810 ( .A1(n9643), .A2(n8233), .ZN(n8262) );
  NAND2_X1 U9811 ( .A1(n9291), .A2(n8306), .ZN(n8261) );
  NAND2_X1 U9812 ( .A1(n8262), .A2(n8261), .ZN(n8263) );
  XNOR2_X1 U9813 ( .A(n8263), .B(n9152), .ZN(n8265) );
  AND2_X1 U9814 ( .A1(n9291), .A2(n9149), .ZN(n8264) );
  AOI21_X1 U9815 ( .B1(n9643), .B2(n8306), .A(n8264), .ZN(n8266) );
  NAND2_X1 U9816 ( .A1(n8265), .A2(n8266), .ZN(n9223) );
  INV_X1 U9817 ( .A(n8265), .ZN(n8268) );
  INV_X1 U9818 ( .A(n8266), .ZN(n8267) );
  NAND2_X1 U9819 ( .A1(n8268), .A2(n8267), .ZN(n9224) );
  NAND2_X1 U9820 ( .A1(n8269), .A2(n9224), .ZN(n9164) );
  INV_X1 U9821 ( .A(n9164), .ZN(n8275) );
  OAI22_X1 U9822 ( .A1(n9848), .A2(n8293), .B1(n9246), .B2(n8284), .ZN(n8270)
         );
  XNOR2_X1 U9823 ( .A(n8270), .B(n8277), .ZN(n9165) );
  OR2_X1 U9824 ( .A1(n9848), .A2(n8284), .ZN(n8272) );
  NAND2_X1 U9825 ( .A1(n9610), .A2(n9149), .ZN(n8271) );
  NAND2_X1 U9826 ( .A1(n8272), .A2(n8271), .ZN(n9166) );
  NAND2_X1 U9827 ( .A1(n9165), .A2(n9166), .ZN(n8273) );
  AOI22_X1 U9828 ( .A1(n9782), .A2(n8233), .B1(n9148), .B2(n9290), .ZN(n8276)
         );
  XOR2_X1 U9829 ( .A(n8277), .B(n8276), .Z(n9241) );
  OAI22_X1 U9830 ( .A1(n9605), .A2(n8284), .B1(n9584), .B2(n8310), .ZN(n9242)
         );
  OAI22_X1 U9831 ( .A1(n9843), .A2(n8293), .B1(n9569), .B2(n8284), .ZN(n8278)
         );
  XNOR2_X1 U9832 ( .A(n8278), .B(n9152), .ZN(n8282) );
  OR2_X1 U9833 ( .A1(n9843), .A2(n8284), .ZN(n8280) );
  NAND2_X1 U9834 ( .A1(n9609), .A2(n9149), .ZN(n8279) );
  NAND2_X1 U9835 ( .A1(n8282), .A2(n8281), .ZN(n9215) );
  OAI21_X1 U9836 ( .B1(n8282), .B2(n8281), .A(n9215), .ZN(n9137) );
  OAI22_X1 U9837 ( .A1(n9576), .A2(n8293), .B1(n9585), .B2(n8284), .ZN(n8283)
         );
  XNOR2_X1 U9838 ( .A(n8283), .B(n9152), .ZN(n8287) );
  OR2_X1 U9839 ( .A1(n9576), .A2(n8284), .ZN(n8286) );
  NAND2_X1 U9840 ( .A1(n9289), .A2(n9149), .ZN(n8285) );
  NAND2_X1 U9841 ( .A1(n8287), .A2(n8288), .ZN(n8292) );
  INV_X1 U9842 ( .A(n8287), .ZN(n8290) );
  INV_X1 U9843 ( .A(n8288), .ZN(n8289) );
  NAND2_X1 U9844 ( .A1(n8290), .A2(n8289), .ZN(n8291) );
  OAI22_X1 U9845 ( .A1(n9838), .A2(n8284), .B1(n9570), .B2(n8310), .ZN(n8299)
         );
  OAI22_X1 U9846 ( .A1(n9838), .A2(n8293), .B1(n9570), .B2(n8284), .ZN(n8294)
         );
  XNOR2_X1 U9847 ( .A(n8294), .B(n8277), .ZN(n8300) );
  XOR2_X1 U9848 ( .A(n8299), .B(n8300), .Z(n9188) );
  NAND2_X1 U9849 ( .A1(n9187), .A2(n9188), .ZN(n9186) );
  NAND2_X1 U9850 ( .A1(n9763), .A2(n8233), .ZN(n8296) );
  NAND2_X1 U9851 ( .A1(n9288), .A2(n8306), .ZN(n8295) );
  NAND2_X1 U9852 ( .A1(n8296), .A2(n8295), .ZN(n8297) );
  XNOR2_X1 U9853 ( .A(n8297), .B(n9152), .ZN(n8302) );
  AND2_X1 U9854 ( .A1(n9288), .A2(n9149), .ZN(n8298) );
  AOI21_X1 U9855 ( .B1(n9763), .B2(n9148), .A(n8298), .ZN(n8303) );
  XNOR2_X1 U9856 ( .A(n8302), .B(n8303), .ZN(n9261) );
  NOR2_X1 U9857 ( .A1(n8300), .A2(n8299), .ZN(n9262) );
  NOR2_X1 U9858 ( .A1(n9261), .A2(n9262), .ZN(n8301) );
  INV_X1 U9859 ( .A(n8302), .ZN(n8305) );
  INV_X1 U9860 ( .A(n8303), .ZN(n8304) );
  NAND2_X1 U9861 ( .A1(n9529), .A2(n8233), .ZN(n8308) );
  INV_X1 U9862 ( .A(n9537), .ZN(n9498) );
  NAND2_X1 U9863 ( .A1(n9498), .A2(n8306), .ZN(n8307) );
  NAND2_X1 U9864 ( .A1(n8308), .A2(n8307), .ZN(n8309) );
  XNOR2_X1 U9865 ( .A(n8309), .B(n9152), .ZN(n8313) );
  INV_X1 U9866 ( .A(n8313), .ZN(n8315) );
  NOR2_X1 U9867 ( .A1(n9537), .A2(n8310), .ZN(n8311) );
  AOI21_X1 U9868 ( .B1(n9529), .B2(n9148), .A(n8311), .ZN(n8312) );
  INV_X1 U9869 ( .A(n8312), .ZN(n8314) );
  AOI21_X1 U9870 ( .B1(n8315), .B2(n8314), .A(n9161), .ZN(n8316) );
  INV_X1 U9871 ( .A(n8316), .ZN(n8317) );
  NOR2_X1 U9872 ( .A1(n8317), .A2(n4530), .ZN(n8318) );
  NOR2_X1 U9873 ( .A1(n9923), .A2(n9518), .ZN(n8320) );
  OAI22_X1 U9874 ( .A1(n9524), .A2(n9279), .B1(n9890), .B2(n9525), .ZN(n8319)
         );
  AOI211_X1 U9875 ( .C1(P1_REG3_REG_27__SCAN_IN), .C2(P1_U3086), .A(n8320), 
        .B(n8319), .ZN(n8321) );
  AND2_X1 U9876 ( .A1(n8323), .A2(n8937), .ZN(n8714) );
  NOR2_X1 U9877 ( .A1(n8324), .A2(n8820), .ZN(n8325) );
  AOI211_X1 U9878 ( .C1(n8920), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8714), .B(
        n8325), .ZN(n8326) );
  OAI222_X1 U9879 ( .A1(n9117), .A2(n9876), .B1(n8330), .B2(P2_U3151), .C1(
        n8329), .C2(n9122), .ZN(P2_U3266) );
  OAI21_X1 U9880 ( .B1(n8332), .B2(n4597), .A(n8331), .ZN(n8333) );
  NAND2_X1 U9881 ( .A1(n8333), .A2(n9906), .ZN(n8337) );
  AOI22_X1 U9882 ( .A1(n8335), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n9900), .B2(
        n8334), .ZN(n8336) );
  OAI211_X1 U9883 ( .C1(n8338), .C2(n9903), .A(n8337), .B(n8336), .ZN(P1_U3237) );
  AOI22_X1 U9884 ( .A1(n8340), .A2(n8515), .B1(n8339), .B2(n8534), .ZN(n8343)
         );
  NAND2_X1 U9885 ( .A1(n8341), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8342) );
  OAI211_X1 U9886 ( .C1(n6678), .C2(n8544), .A(n8343), .B(n8342), .ZN(P2_U3172) );
  INV_X1 U9887 ( .A(n8344), .ZN(n9875) );
  OAI222_X1 U9888 ( .A1(n9105), .A2(n8346), .B1(n9117), .B2(n9875), .C1(
        P2_U3151), .C2(n8345), .ZN(P2_U3265) );
  INV_X1 U9889 ( .A(n8347), .ZN(n8348) );
  NAND2_X1 U9890 ( .A1(n8348), .A2(n8556), .ZN(n8349) );
  XNOR2_X1 U9891 ( .A(n10084), .B(n8421), .ZN(n8351) );
  XNOR2_X1 U9892 ( .A(n8351), .B(n8912), .ZN(n8437) );
  INV_X1 U9893 ( .A(n8351), .ZN(n8352) );
  NAND2_X1 U9894 ( .A1(n8352), .A2(n8912), .ZN(n8353) );
  NAND2_X1 U9895 ( .A1(n8354), .A2(n8353), .ZN(n8494) );
  XNOR2_X1 U9896 ( .A(n9097), .B(n8421), .ZN(n8355) );
  NAND2_X1 U9897 ( .A1(n8355), .A2(n8439), .ZN(n8492) );
  NAND2_X1 U9898 ( .A1(n8494), .A2(n8492), .ZN(n8357) );
  INV_X1 U9899 ( .A(n8355), .ZN(n8356) );
  NAND2_X1 U9900 ( .A1(n8356), .A2(n8896), .ZN(n8493) );
  XNOR2_X1 U9901 ( .A(n9090), .B(n8421), .ZN(n8358) );
  XNOR2_X1 U9902 ( .A(n8358), .B(n8496), .ZN(n8398) );
  NAND2_X1 U9903 ( .A1(n8358), .A2(n8496), .ZN(n8359) );
  XNOR2_X1 U9904 ( .A(n9084), .B(n8421), .ZN(n8362) );
  XNOR2_X1 U9905 ( .A(n8362), .B(n8399), .ZN(n8539) );
  INV_X1 U9906 ( .A(n8539), .ZN(n8360) );
  NAND2_X1 U9907 ( .A1(n8361), .A2(n8360), .ZN(n8541) );
  INV_X1 U9908 ( .A(n8362), .ZN(n8363) );
  NAND2_X1 U9909 ( .A1(n8363), .A2(n8897), .ZN(n8364) );
  NAND2_X1 U9910 ( .A1(n8541), .A2(n8364), .ZN(n8456) );
  XNOR2_X1 U9911 ( .A(n8461), .B(n8421), .ZN(n8365) );
  XNOR2_X1 U9912 ( .A(n8365), .B(n8543), .ZN(n8455) );
  NAND2_X1 U9913 ( .A1(n8365), .A2(n8885), .ZN(n8366) );
  XNOR2_X1 U9914 ( .A(n9072), .B(n8421), .ZN(n8368) );
  XNOR2_X1 U9915 ( .A(n8368), .B(n8855), .ZN(n8464) );
  NAND2_X1 U9916 ( .A1(n8368), .A2(n8855), .ZN(n8510) );
  NAND2_X1 U9917 ( .A1(n8462), .A2(n8510), .ZN(n8369) );
  XNOR2_X1 U9918 ( .A(n8988), .B(n8421), .ZN(n8370) );
  XNOR2_X1 U9919 ( .A(n8370), .B(n8864), .ZN(n8511) );
  NAND2_X1 U9920 ( .A1(n8370), .A2(n8466), .ZN(n8371) );
  XNOR2_X1 U9921 ( .A(n9062), .B(n7199), .ZN(n8372) );
  XNOR2_X1 U9922 ( .A(n8372), .B(n8854), .ZN(n8411) );
  INV_X1 U9923 ( .A(n8372), .ZN(n8373) );
  NAND2_X1 U9924 ( .A1(n8373), .A2(n8854), .ZN(n8374) );
  XNOR2_X1 U9925 ( .A(n9056), .B(n8421), .ZN(n8375) );
  XNOR2_X1 U9926 ( .A(n8375), .B(n8841), .ZN(n8486) );
  NAND2_X1 U9927 ( .A1(n8485), .A2(n8486), .ZN(n8377) );
  NAND2_X1 U9928 ( .A1(n8375), .A2(n8808), .ZN(n8376) );
  NAND2_X1 U9929 ( .A1(n8377), .A2(n8376), .ZN(n8429) );
  XNOR2_X1 U9930 ( .A(n8817), .B(n8421), .ZN(n8378) );
  XNOR2_X1 U9931 ( .A(n8378), .B(n8831), .ZN(n8430) );
  NAND2_X1 U9932 ( .A1(n8429), .A2(n8430), .ZN(n8380) );
  NAND2_X1 U9933 ( .A1(n8378), .A2(n8798), .ZN(n8379) );
  NAND2_X1 U9934 ( .A1(n8380), .A2(n8379), .ZN(n8502) );
  XNOR2_X1 U9935 ( .A(n8507), .B(n8421), .ZN(n8381) );
  XNOR2_X1 U9936 ( .A(n8381), .B(n8788), .ZN(n8503) );
  AND2_X1 U9937 ( .A1(n8381), .A2(n8809), .ZN(n8382) );
  XNOR2_X1 U9938 ( .A(n9035), .B(n8421), .ZN(n8476) );
  XNOR2_X1 U9939 ( .A(n9041), .B(n7199), .ZN(n8472) );
  INV_X1 U9940 ( .A(n8472), .ZN(n8383) );
  OAI22_X1 U9941 ( .A1(n8476), .A2(n8475), .B1(n8799), .B2(n8383), .ZN(n8387)
         );
  OAI21_X1 U9942 ( .B1(n8472), .B2(n8776), .A(n8789), .ZN(n8385) );
  NOR2_X1 U9943 ( .A1(n8789), .A2(n8776), .ZN(n8384) );
  AOI22_X1 U9944 ( .A1(n8385), .A2(n8476), .B1(n8384), .B2(n8383), .ZN(n8386)
         );
  XNOR2_X1 U9945 ( .A(n9029), .B(n8421), .ZN(n8388) );
  XNOR2_X1 U9946 ( .A(n8388), .B(n8777), .ZN(n8448) );
  XNOR2_X1 U9947 ( .A(n9023), .B(n8421), .ZN(n8390) );
  NOR2_X1 U9948 ( .A1(n8390), .A2(n8389), .ZN(n8525) );
  NAND2_X1 U9949 ( .A1(n8390), .A2(n8389), .ZN(n8523) );
  XNOR2_X1 U9950 ( .A(n8743), .B(n8421), .ZN(n8418) );
  XNOR2_X1 U9951 ( .A(n8418), .B(n8530), .ZN(n8419) );
  XNOR2_X1 U9952 ( .A(n8420), .B(n8419), .ZN(n8396) );
  AOI22_X1 U9953 ( .A1(n8760), .A2(n8548), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8392) );
  NAND2_X1 U9954 ( .A1(n8739), .A2(n8533), .ZN(n8391) );
  OAI211_X1 U9955 ( .C1(n8393), .C2(n8544), .A(n8392), .B(n8391), .ZN(n8394)
         );
  AOI21_X1 U9956 ( .B1(n8743), .B2(n8534), .A(n8394), .ZN(n8395) );
  OAI21_X1 U9957 ( .B1(n8396), .B2(n8538), .A(n8395), .ZN(P2_U3154) );
  XOR2_X1 U9958 ( .A(n8398), .B(n8397), .Z(n8404) );
  NAND2_X1 U9959 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8597) );
  OAI21_X1 U9960 ( .B1(n8544), .B2(n8399), .A(n8597), .ZN(n8400) );
  AOI21_X1 U9961 ( .B1(n8548), .B2(n8896), .A(n8400), .ZN(n8401) );
  OAI21_X1 U9962 ( .B1(n8900), .B2(n8545), .A(n8401), .ZN(n8402) );
  AOI21_X1 U9963 ( .B1(n9090), .B2(n8534), .A(n8402), .ZN(n8403) );
  OAI21_X1 U9964 ( .B1(n8404), .B2(n8538), .A(n8403), .ZN(P2_U3155) );
  XNOR2_X1 U9965 ( .A(n8473), .B(n8472), .ZN(n8474) );
  XNOR2_X1 U9966 ( .A(n8474), .B(n8799), .ZN(n8409) );
  AOI22_X1 U9967 ( .A1(n8548), .A2(n8788), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8406) );
  NAND2_X1 U9968 ( .A1(n8533), .A2(n8792), .ZN(n8405) );
  OAI211_X1 U9969 ( .C1(n8475), .C2(n8544), .A(n8406), .B(n8405), .ZN(n8407)
         );
  AOI21_X1 U9970 ( .B1(n9041), .B2(n8534), .A(n8407), .ZN(n8408) );
  OAI21_X1 U9971 ( .B1(n8409), .B2(n8538), .A(n8408), .ZN(P2_U3156) );
  XOR2_X1 U9972 ( .A(n8411), .B(n8410), .Z(n8417) );
  INV_X1 U9973 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8412) );
  OAI22_X1 U9974 ( .A1(n8544), .A2(n8808), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8412), .ZN(n8413) );
  AOI21_X1 U9975 ( .B1(n8548), .B2(n8864), .A(n8413), .ZN(n8414) );
  OAI21_X1 U9976 ( .B1(n8844), .B2(n8545), .A(n8414), .ZN(n8415) );
  AOI21_X1 U9977 ( .B1(n9062), .B2(n8534), .A(n8415), .ZN(n8416) );
  OAI21_X1 U9978 ( .B1(n8417), .B2(n8538), .A(n8416), .ZN(P2_U3159) );
  XNOR2_X1 U9979 ( .A(n8718), .B(n8421), .ZN(n8422) );
  XNOR2_X1 U9980 ( .A(n8423), .B(n8422), .ZN(n8428) );
  AOI22_X1 U9981 ( .A1(n8750), .A2(n8548), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8425) );
  NAND2_X1 U9982 ( .A1(n8728), .A2(n8533), .ZN(n8424) );
  OAI211_X1 U9983 ( .C1(n8555), .C2(n8544), .A(n8425), .B(n8424), .ZN(n8426)
         );
  AOI21_X1 U9984 ( .B1(n9016), .B2(n8534), .A(n8426), .ZN(n8427) );
  OAI21_X1 U9985 ( .B1(n8428), .B2(n8538), .A(n8427), .ZN(P2_U3160) );
  XOR2_X1 U9986 ( .A(n8430), .B(n8429), .Z(n8436) );
  OAI22_X1 U9987 ( .A1(n8544), .A2(n8809), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8431), .ZN(n8433) );
  INV_X1 U9988 ( .A(n8548), .ZN(n8528) );
  NOR2_X1 U9989 ( .A1(n8528), .A2(n8808), .ZN(n8432) );
  AOI211_X1 U9990 ( .C1(n8818), .C2(n8533), .A(n8433), .B(n8432), .ZN(n8435)
         );
  NAND2_X1 U9991 ( .A1(n8817), .A2(n8534), .ZN(n8434) );
  OAI211_X1 U9992 ( .C1(n8436), .C2(n8538), .A(n8435), .B(n8434), .ZN(P2_U3163) );
  XNOR2_X1 U9993 ( .A(n8438), .B(n8437), .ZN(n8446) );
  NOR2_X1 U9994 ( .A1(n8544), .A2(n8439), .ZN(n8440) );
  AOI211_X1 U9995 ( .C1(n8548), .C2(n8556), .A(n8441), .B(n8440), .ZN(n8442)
         );
  OAI21_X1 U9996 ( .B1(n8443), .B2(n8545), .A(n8442), .ZN(n8444) );
  AOI21_X1 U9997 ( .B1(n10084), .B2(n8534), .A(n8444), .ZN(n8445) );
  OAI21_X1 U9998 ( .B1(n8446), .B2(n8538), .A(n8445), .ZN(P2_U3164) );
  XOR2_X1 U9999 ( .A(n8448), .B(n8447), .Z(n8453) );
  INV_X1 U10000 ( .A(n8544), .ZN(n8479) );
  AOI22_X1 U10001 ( .A1(n8760), .A2(n8479), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8450) );
  NAND2_X1 U10002 ( .A1(n8533), .A2(n8762), .ZN(n8449) );
  OAI211_X1 U10003 ( .C1(n8475), .C2(n8528), .A(n8450), .B(n8449), .ZN(n8451)
         );
  AOI21_X1 U10004 ( .B1(n9029), .B2(n8534), .A(n8451), .ZN(n8452) );
  OAI21_X1 U10005 ( .B1(n8453), .B2(n8538), .A(n8452), .ZN(P2_U3165) );
  OAI211_X1 U10006 ( .C1(n8456), .C2(n8455), .A(n8454), .B(n8515), .ZN(n8460)
         );
  NAND2_X1 U10007 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8639) );
  OAI21_X1 U10008 ( .B1(n8544), .B2(n8855), .A(n8639), .ZN(n8458) );
  NOR2_X1 U10009 ( .A1(n8545), .A2(n8877), .ZN(n8457) );
  AOI211_X1 U10010 ( .C1(n8548), .C2(n8897), .A(n8458), .B(n8457), .ZN(n8459)
         );
  OAI211_X1 U10011 ( .C1(n8461), .C2(n8551), .A(n8460), .B(n8459), .ZN(
        P2_U3166) );
  INV_X1 U10012 ( .A(n8462), .ZN(n8513) );
  AOI21_X1 U10013 ( .B1(n8464), .B2(n8463), .A(n8513), .ZN(n8471) );
  OAI22_X1 U10014 ( .A1(n8544), .A2(n8466), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8465), .ZN(n8467) );
  AOI21_X1 U10015 ( .B1(n8548), .B2(n8885), .A(n8467), .ZN(n8468) );
  OAI21_X1 U10016 ( .B1(n8867), .B2(n8545), .A(n8468), .ZN(n8469) );
  AOI21_X1 U10017 ( .B1(n9072), .B2(n8534), .A(n8469), .ZN(n8470) );
  OAI21_X1 U10018 ( .B1(n8471), .B2(n8538), .A(n8470), .ZN(P2_U3168) );
  OAI22_X1 U10019 ( .A1(n8474), .A2(n8776), .B1(n8473), .B2(n8472), .ZN(n8478)
         );
  XNOR2_X1 U10020 ( .A(n8476), .B(n8475), .ZN(n8477) );
  XNOR2_X1 U10021 ( .A(n8478), .B(n8477), .ZN(n8484) );
  AOI22_X1 U10022 ( .A1(n8777), .A2(n8479), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8481) );
  NAND2_X1 U10023 ( .A1(n8533), .A2(n8779), .ZN(n8480) );
  OAI211_X1 U10024 ( .C1(n8799), .C2(n8528), .A(n8481), .B(n8480), .ZN(n8482)
         );
  AOI21_X1 U10025 ( .B1(n9035), .B2(n8534), .A(n8482), .ZN(n8483) );
  OAI21_X1 U10026 ( .B1(n8484), .B2(n8538), .A(n8483), .ZN(P2_U3169) );
  XOR2_X1 U10027 ( .A(n8486), .B(n8485), .Z(n8491) );
  OAI22_X1 U10028 ( .A1(n8544), .A2(n8798), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10380), .ZN(n8488) );
  NOR2_X1 U10029 ( .A1(n8528), .A2(n8854), .ZN(n8487) );
  AOI211_X1 U10030 ( .C1(n8834), .C2(n8533), .A(n8488), .B(n8487), .ZN(n8490)
         );
  NAND2_X1 U10031 ( .A1(n9056), .A2(n8534), .ZN(n8489) );
  OAI211_X1 U10032 ( .C1(n8491), .C2(n8538), .A(n8490), .B(n8489), .ZN(
        P2_U3173) );
  NAND2_X1 U10033 ( .A1(n8493), .A2(n8492), .ZN(n8495) );
  XOR2_X1 U10034 ( .A(n8495), .B(n8494), .Z(n8501) );
  OR2_X1 U10035 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10480), .ZN(n8573) );
  OAI21_X1 U10036 ( .B1(n8544), .B2(n8496), .A(n8573), .ZN(n8497) );
  AOI21_X1 U10037 ( .B1(n8548), .B2(n8912), .A(n8497), .ZN(n8498) );
  OAI21_X1 U10038 ( .B1(n8918), .B2(n8545), .A(n8498), .ZN(n8499) );
  AOI21_X1 U10039 ( .B1(n9097), .B2(n8534), .A(n8499), .ZN(n8500) );
  OAI21_X1 U10040 ( .B1(n8501), .B2(n8538), .A(n8500), .ZN(P2_U3174) );
  XOR2_X1 U10041 ( .A(n8503), .B(n8502), .Z(n8509) );
  AOI22_X1 U10042 ( .A1(n8548), .A2(n8831), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8505) );
  NAND2_X1 U10043 ( .A1(n8533), .A2(n8802), .ZN(n8504) );
  OAI211_X1 U10044 ( .C1(n8799), .C2(n8544), .A(n8505), .B(n8504), .ZN(n8506)
         );
  AOI21_X1 U10045 ( .B1(n8507), .B2(n8534), .A(n8506), .ZN(n8508) );
  OAI21_X1 U10046 ( .B1(n8509), .B2(n8538), .A(n8508), .ZN(P2_U3175) );
  INV_X1 U10047 ( .A(n8510), .ZN(n8512) );
  NOR3_X1 U10048 ( .A1(n8513), .A2(n8512), .A3(n8511), .ZN(n8517) );
  INV_X1 U10049 ( .A(n8514), .ZN(n8516) );
  OAI21_X1 U10050 ( .B1(n8517), .B2(n8516), .A(n8515), .ZN(n8521) );
  NAND2_X1 U10051 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8682) );
  OAI21_X1 U10052 ( .B1(n8544), .B2(n8854), .A(n8682), .ZN(n8519) );
  NOR2_X1 U10053 ( .A1(n8545), .A2(n8856), .ZN(n8518) );
  AOI211_X1 U10054 ( .C1(n8548), .C2(n8874), .A(n8519), .B(n8518), .ZN(n8520)
         );
  OAI211_X1 U10055 ( .C1(n8522), .C2(n8551), .A(n8521), .B(n8520), .ZN(
        P2_U3178) );
  INV_X1 U10056 ( .A(n8523), .ZN(n8524) );
  NOR2_X1 U10057 ( .A1(n8525), .A2(n8524), .ZN(n8526) );
  XNOR2_X1 U10058 ( .A(n8527), .B(n8526), .ZN(n8537) );
  INV_X1 U10059 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10274) );
  OAI22_X1 U10060 ( .A1(n8529), .A2(n8528), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10274), .ZN(n8532) );
  NOR2_X1 U10061 ( .A1(n8530), .A2(n8544), .ZN(n8531) );
  AOI211_X1 U10062 ( .C1(n8753), .C2(n8533), .A(n8532), .B(n8531), .ZN(n8536)
         );
  NAND2_X1 U10063 ( .A1(n9023), .A2(n8534), .ZN(n8535) );
  OAI211_X1 U10064 ( .C1(n8537), .C2(n8538), .A(n8536), .B(n8535), .ZN(
        P2_U3180) );
  INV_X1 U10065 ( .A(n9084), .ZN(n8552) );
  AOI21_X1 U10066 ( .B1(n8540), .B2(n8539), .A(n8538), .ZN(n8542) );
  NAND2_X1 U10067 ( .A1(n8542), .A2(n8541), .ZN(n8550) );
  NAND2_X1 U10068 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8617) );
  OAI21_X1 U10069 ( .B1(n8544), .B2(n8543), .A(n8617), .ZN(n8547) );
  NOR2_X1 U10070 ( .A1(n8545), .A2(n8888), .ZN(n8546) );
  AOI211_X1 U10071 ( .C1(n8548), .C2(n8910), .A(n8547), .B(n8546), .ZN(n8549)
         );
  OAI211_X1 U10072 ( .C1(n8552), .C2(n8551), .A(n8550), .B(n8549), .ZN(
        P2_U3181) );
  INV_X1 U10073 ( .A(n8553), .ZN(n8713) );
  MUX2_X1 U10074 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8713), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10075 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8554), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10076 ( .A(n8555), .ZN(n8722) );
  MUX2_X1 U10077 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8722), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10078 ( .A(n8736), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8680), .Z(
        P2_U3519) );
  MUX2_X1 U10079 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8750), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10080 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8760), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10081 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8777), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10082 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8789), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10083 ( .A(n8776), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8680), .Z(
        P2_U3514) );
  MUX2_X1 U10084 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8788), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10085 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8831), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10086 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8841), .S(P2_U3893), .Z(
        P2_U3511) );
  INV_X1 U10087 ( .A(n8854), .ZN(n8830) );
  MUX2_X1 U10088 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8830), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10089 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8864), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8874), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10091 ( .A(n8885), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8680), .Z(
        P2_U3507) );
  MUX2_X1 U10092 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8897), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10093 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8910), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10094 ( .A(n8896), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8680), .Z(
        P2_U3504) );
  MUX2_X1 U10095 ( .A(n8912), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8680), .Z(
        P2_U3503) );
  MUX2_X1 U10096 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8556), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10097 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8557), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10098 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8558), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10099 ( .A(n8559), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8680), .Z(
        P2_U3499) );
  MUX2_X1 U10100 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8560), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10101 ( .A(n8561), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8680), .Z(
        P2_U3497) );
  MUX2_X1 U10102 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8562), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10103 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n6526), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10104 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8563), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10105 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8564), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10106 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8565), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10107 ( .A(n8566), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8680), .Z(
        P2_U3491) );
  AOI21_X1 U10108 ( .B1(n9003), .B2(n8568), .A(n8600), .ZN(n8585) );
  AOI21_X1 U10109 ( .B1(n8572), .B2(n8571), .A(n8587), .ZN(n8574) );
  OAI21_X1 U10110 ( .B1(n10026), .B2(n8574), .A(n8573), .ZN(n8576) );
  INV_X1 U10111 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10138) );
  NOR2_X1 U10112 ( .A1(n10011), .A2(n10138), .ZN(n8575) );
  AOI211_X1 U10113 ( .C1(n10014), .C2(n8599), .A(n8576), .B(n8575), .ZN(n8584)
         );
  AOI21_X1 U10114 ( .B1(n8579), .B2(n8578), .A(n8577), .ZN(n8581) );
  MUX2_X1 U10115 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8699), .Z(n8590) );
  XNOR2_X1 U10116 ( .A(n8590), .B(n8599), .ZN(n8580) );
  NAND2_X1 U10117 ( .A1(n8581), .A2(n8580), .ZN(n8592) );
  OAI21_X1 U10118 ( .B1(n8581), .B2(n8580), .A(n8592), .ZN(n8582) );
  NAND2_X1 U10119 ( .A1(n8582), .A2(n10020), .ZN(n8583) );
  OAI211_X1 U10120 ( .C1(n8585), .C2(n10022), .A(n8584), .B(n8583), .ZN(
        P2_U3195) );
  NOR2_X1 U10121 ( .A1(n8599), .A2(n8586), .ZN(n8588) );
  AOI22_X1 U10122 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8602), .B1(n8619), .B2(
        n6273), .ZN(n8589) );
  AOI21_X1 U10123 ( .B1(n4583), .B2(n8589), .A(n8610), .ZN(n8609) );
  MUX2_X1 U10124 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8699), .Z(n8612) );
  XNOR2_X1 U10125 ( .A(n8612), .B(n8602), .ZN(n8595) );
  INV_X1 U10126 ( .A(n8590), .ZN(n8591) );
  NAND2_X1 U10127 ( .A1(n8599), .A2(n8591), .ZN(n8593) );
  NAND2_X1 U10128 ( .A1(n8593), .A2(n8592), .ZN(n8594) );
  NAND2_X1 U10129 ( .A1(n8595), .A2(n8594), .ZN(n8613) );
  OAI21_X1 U10130 ( .B1(n8595), .B2(n8594), .A(n8613), .ZN(n8607) );
  NAND2_X1 U10131 ( .A1(n10018), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8596) );
  OAI211_X1 U10132 ( .C1(n8679), .C2(n8619), .A(n8597), .B(n8596), .ZN(n8606)
         );
  NOR2_X1 U10133 ( .A1(n8599), .A2(n8598), .ZN(n8601) );
  AOI22_X1 U10134 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8602), .B1(n8619), .B2(
        n9000), .ZN(n8603) );
  AOI21_X1 U10135 ( .B1(n4588), .B2(n8603), .A(n8620), .ZN(n8604) );
  NOR2_X1 U10136 ( .A1(n8604), .A2(n10022), .ZN(n8605) );
  AOI211_X1 U10137 ( .C1(n10020), .C2(n8607), .A(n8606), .B(n8605), .ZN(n8608)
         );
  OAI21_X1 U10138 ( .B1(n8609), .B2(n10026), .A(n8608), .ZN(P2_U3196) );
  AOI21_X1 U10139 ( .B1(n8611), .B2(n8887), .A(n8629), .ZN(n8627) );
  MUX2_X1 U10140 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8699), .Z(n8634) );
  XNOR2_X1 U10141 ( .A(n8634), .B(n8641), .ZN(n8616) );
  OR2_X1 U10142 ( .A1(n8612), .A2(n8619), .ZN(n8614) );
  NAND2_X1 U10143 ( .A1(n8614), .A2(n8613), .ZN(n8615) );
  NAND2_X1 U10144 ( .A1(n8616), .A2(n8615), .ZN(n8635) );
  OAI21_X1 U10145 ( .B1(n8616), .B2(n8615), .A(n8635), .ZN(n8625) );
  INV_X1 U10146 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U10147 ( .A1(n10014), .A2(n8641), .ZN(n8618) );
  OAI211_X1 U10148 ( .C1(n10144), .C2(n10011), .A(n8618), .B(n8617), .ZN(n8624) );
  XOR2_X1 U10149 ( .A(n4525), .B(n8633), .Z(n8621) );
  NOR2_X1 U10150 ( .A1(n8997), .A2(n8621), .ZN(n8642) );
  AOI21_X1 U10151 ( .B1(n8997), .B2(n8621), .A(n8642), .ZN(n8622) );
  NOR2_X1 U10152 ( .A1(n8622), .A2(n10022), .ZN(n8623) );
  AOI211_X1 U10153 ( .C1(n10020), .C2(n8625), .A(n8624), .B(n8623), .ZN(n8626)
         );
  OAI21_X1 U10154 ( .B1(n8627), .B2(n10026), .A(n8626), .ZN(P2_U3197) );
  NOR2_X1 U10155 ( .A1(n8641), .A2(n8628), .ZN(n8630) );
  NAND2_X1 U10156 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8658), .ZN(n8631) );
  OAI21_X1 U10157 ( .B1(n8658), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8631), .ZN(
        n8632) );
  AOI21_X1 U10158 ( .B1(n4552), .B2(n8632), .A(n8657), .ZN(n8652) );
  MUX2_X1 U10159 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8699), .Z(n8656) );
  XNOR2_X1 U10160 ( .A(n8656), .B(n8644), .ZN(n8638) );
  OR2_X1 U10161 ( .A1(n8634), .A2(n8633), .ZN(n8636) );
  NAND2_X1 U10162 ( .A1(n8636), .A2(n8635), .ZN(n8637) );
  NAND2_X1 U10163 ( .A1(n8638), .A2(n8637), .ZN(n8655) );
  OAI21_X1 U10164 ( .B1(n8638), .B2(n8637), .A(n8655), .ZN(n8650) );
  INV_X1 U10165 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10148) );
  NAND2_X1 U10166 ( .A1(n10014), .A2(n8644), .ZN(n8640) );
  OAI211_X1 U10167 ( .C1(n10148), .C2(n10011), .A(n8640), .B(n8639), .ZN(n8649) );
  NOR2_X1 U10168 ( .A1(n8641), .A2(n4525), .ZN(n8643) );
  NOR2_X1 U10169 ( .A1(n8643), .A2(n8642), .ZN(n8646) );
  AOI22_X1 U10170 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8644), .B1(n8658), .B2(
        n8994), .ZN(n8645) );
  NOR2_X1 U10171 ( .A1(n8646), .A2(n8645), .ZN(n8653) );
  AOI21_X1 U10172 ( .B1(n8646), .B2(n8645), .A(n8653), .ZN(n8647) );
  NOR2_X1 U10173 ( .A1(n8647), .A2(n10022), .ZN(n8648) );
  AOI211_X1 U10174 ( .C1(n10020), .C2(n8650), .A(n8649), .B(n8648), .ZN(n8651)
         );
  OAI21_X1 U10175 ( .B1(n8652), .B2(n10026), .A(n8651), .ZN(P2_U3198) );
  AOI21_X1 U10176 ( .B1(n8991), .B2(n8654), .A(n8686), .ZN(n8666) );
  MUX2_X1 U10177 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8699), .Z(n8672) );
  XNOR2_X1 U10178 ( .A(n8672), .B(n8685), .ZN(n8675) );
  XNOR2_X1 U10179 ( .A(n8675), .B(n8674), .ZN(n8665) );
  NOR2_X1 U10180 ( .A1(n8866), .A2(n8659), .ZN(n8668) );
  INV_X2 U10181 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  OAI21_X1 U10182 ( .B1(n8666), .B2(n10022), .A(n4573), .ZN(P2_U3199) );
  NOR2_X1 U10183 ( .A1(n8685), .A2(n8667), .ZN(n8669) );
  NOR2_X1 U10184 ( .A1(n8669), .A2(n8668), .ZN(n8671) );
  NAND2_X1 U10185 ( .A1(n8687), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8691) );
  OAI21_X1 U10186 ( .B1(n8687), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8691), .ZN(
        n8670) );
  NOR2_X1 U10187 ( .A1(n8671), .A2(n8670), .ZN(n8693) );
  AOI21_X1 U10188 ( .B1(n8671), .B2(n8670), .A(n8693), .ZN(n8690) );
  INV_X1 U10189 ( .A(n8672), .ZN(n8673) );
  MUX2_X1 U10190 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8699), .Z(n8676) );
  INV_X1 U10191 ( .A(n8698), .ZN(n8678) );
  NAND2_X1 U10192 ( .A1(n8677), .A2(n8676), .ZN(n8696) );
  NAND2_X1 U10193 ( .A1(n8678), .A2(n8696), .ZN(n8681) );
  OAI21_X1 U10194 ( .B1(n8681), .B2(n8680), .A(n8679), .ZN(n8689) );
  INV_X1 U10195 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U10196 ( .A1(n8687), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8695) );
  OAI21_X1 U10197 ( .B1(n8687), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8695), .ZN(
        n8688) );
  INV_X1 U10198 ( .A(n8691), .ZN(n8692) );
  NOR2_X1 U10199 ( .A1(n8693), .A2(n8692), .ZN(n8694) );
  MUX2_X1 U10200 ( .A(n8843), .B(P2_REG2_REG_19__SCAN_IN), .S(n8705), .Z(n8700) );
  XNOR2_X1 U10201 ( .A(n8694), .B(n8700), .ZN(n8711) );
  OAI21_X1 U10202 ( .B1(n8698), .B2(n8697), .A(n8696), .ZN(n8702) );
  MUX2_X1 U10203 ( .A(n8700), .B(n4593), .S(n8699), .Z(n8701) );
  XNOR2_X1 U10204 ( .A(n8702), .B(n8701), .ZN(n8708) );
  NAND2_X1 U10205 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8703) );
  OAI21_X1 U10206 ( .B1(n10011), .B2(n10551), .A(n8703), .ZN(n8704) );
  AOI21_X1 U10207 ( .B1(n8705), .B2(n10014), .A(n8704), .ZN(n8706) );
  OAI21_X1 U10208 ( .B1(n8708), .B2(n8707), .A(n8706), .ZN(n8709) );
  OAI21_X1 U10209 ( .B1(n8711), .B2(n10026), .A(n8710), .ZN(P2_U3201) );
  INV_X1 U10210 ( .A(n9008), .ZN(n8946) );
  NAND2_X1 U10211 ( .A1(n8713), .A2(n8712), .ZN(n8944) );
  INV_X1 U10212 ( .A(n8944), .ZN(n9009) );
  AOI21_X1 U10213 ( .B1(n9009), .B2(n8942), .A(n8714), .ZN(n8717) );
  NAND2_X1 U10214 ( .A1(n8920), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8715) );
  OAI211_X1 U10215 ( .C1(n8946), .C2(n8820), .A(n8717), .B(n8715), .ZN(
        P2_U3202) );
  NAND2_X1 U10216 ( .A1(n8920), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8716) );
  OAI211_X1 U10217 ( .C1(n8949), .C2(n8820), .A(n8717), .B(n8716), .ZN(
        P2_U3203) );
  XNOR2_X1 U10218 ( .A(n8719), .B(n8718), .ZN(n9019) );
  INV_X1 U10219 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8727) );
  XNOR2_X1 U10220 ( .A(n8721), .B(n8720), .ZN(n8726) );
  NAND2_X1 U10221 ( .A1(n8722), .A2(n8909), .ZN(n8724) );
  NAND2_X1 U10222 ( .A1(n8750), .A2(n8911), .ZN(n8723) );
  MUX2_X1 U10223 ( .A(n8727), .B(n9014), .S(n8942), .Z(n8730) );
  AOI22_X1 U10224 ( .A1(n9016), .A2(n8890), .B1(n8937), .B2(n8728), .ZN(n8729)
         );
  OAI211_X1 U10225 ( .C1(n9019), .C2(n8923), .A(n8730), .B(n8729), .ZN(
        P2_U3205) );
  XNOR2_X1 U10226 ( .A(n8732), .B(n8731), .ZN(n8956) );
  XNOR2_X1 U10227 ( .A(n8733), .B(n8734), .ZN(n8735) );
  NAND2_X1 U10228 ( .A1(n8735), .A2(n8914), .ZN(n8738) );
  AOI22_X1 U10229 ( .A1(n8736), .A2(n8909), .B1(n8911), .B2(n8760), .ZN(n8737)
         );
  NAND2_X1 U10230 ( .A1(n8738), .A2(n8737), .ZN(n8958) );
  NAND2_X1 U10231 ( .A1(n8958), .A2(n8942), .ZN(n8745) );
  INV_X1 U10232 ( .A(n8739), .ZN(n8741) );
  INV_X1 U10233 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8740) );
  OAI22_X1 U10234 ( .A1(n8741), .A2(n8899), .B1(n8942), .B2(n8740), .ZN(n8742)
         );
  AOI21_X1 U10235 ( .B1(n8743), .B2(n8890), .A(n8742), .ZN(n8744) );
  OAI211_X1 U10236 ( .C1(n8956), .C2(n8923), .A(n8745), .B(n8744), .ZN(
        P2_U3206) );
  XNOR2_X1 U10237 ( .A(n8746), .B(n8749), .ZN(n9026) );
  INV_X1 U10238 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U10239 ( .A1(n8759), .A2(n8758), .ZN(n8748) );
  AOI222_X1 U10240 ( .A1(n8914), .A2(n8751), .B1(n8777), .B2(n8911), .C1(n8750), .C2(n8909), .ZN(n9021) );
  MUX2_X1 U10241 ( .A(n8752), .B(n9021), .S(n8942), .Z(n8755) );
  AOI22_X1 U10242 ( .A1(n9023), .A2(n8890), .B1(n8937), .B2(n8753), .ZN(n8754)
         );
  OAI211_X1 U10243 ( .C1(n9026), .C2(n8923), .A(n8755), .B(n8754), .ZN(
        P2_U3207) );
  XNOR2_X1 U10244 ( .A(n8759), .B(n8758), .ZN(n8761) );
  AOI222_X1 U10245 ( .A1(n8914), .A2(n8761), .B1(n8789), .B2(n8911), .C1(n8760), .C2(n8909), .ZN(n9027) );
  INV_X1 U10246 ( .A(n9027), .ZN(n8766) );
  INV_X1 U10247 ( .A(n9029), .ZN(n8764) );
  INV_X1 U10248 ( .A(n8762), .ZN(n8763) );
  OAI22_X1 U10249 ( .A1(n8764), .A2(n8915), .B1(n8763), .B2(n8899), .ZN(n8765)
         );
  OAI21_X1 U10250 ( .B1(n8766), .B2(n8765), .A(n8942), .ZN(n8768) );
  NAND2_X1 U10251 ( .A1(n8920), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8767) );
  OAI211_X1 U10252 ( .C1(n9032), .C2(n8923), .A(n8768), .B(n8767), .ZN(
        P2_U3208) );
  OR2_X1 U10253 ( .A1(n8769), .A2(n8770), .ZN(n8772) );
  NAND2_X1 U10254 ( .A1(n8772), .A2(n8771), .ZN(n8773) );
  XNOR2_X1 U10255 ( .A(n8774), .B(n8775), .ZN(n8778) );
  AOI222_X1 U10256 ( .A1(n8914), .A2(n8778), .B1(n8777), .B2(n8909), .C1(n8776), .C2(n8911), .ZN(n9033) );
  INV_X1 U10257 ( .A(n9033), .ZN(n8783) );
  INV_X1 U10258 ( .A(n9035), .ZN(n8781) );
  INV_X1 U10259 ( .A(n8779), .ZN(n8780) );
  OAI22_X1 U10260 ( .A1(n8781), .A2(n8915), .B1(n8780), .B2(n8899), .ZN(n8782)
         );
  OAI21_X1 U10261 ( .B1(n8783), .B2(n8782), .A(n8942), .ZN(n8785) );
  NAND2_X1 U10262 ( .A1(n8920), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8784) );
  OAI211_X1 U10263 ( .C1(n9038), .C2(n8923), .A(n8785), .B(n8784), .ZN(
        P2_U3209) );
  XOR2_X1 U10264 ( .A(n8769), .B(n8786), .Z(n9044) );
  INV_X1 U10265 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8791) );
  XNOR2_X1 U10266 ( .A(n8787), .B(n8786), .ZN(n8790) );
  AOI222_X1 U10267 ( .A1(n8914), .A2(n8790), .B1(n8789), .B2(n8909), .C1(n8788), .C2(n8911), .ZN(n9039) );
  MUX2_X1 U10268 ( .A(n8791), .B(n9039), .S(n8942), .Z(n8794) );
  AOI22_X1 U10269 ( .A1(n9041), .A2(n8890), .B1(n8937), .B2(n8792), .ZN(n8793)
         );
  OAI211_X1 U10270 ( .C1(n9044), .C2(n8923), .A(n8794), .B(n8793), .ZN(
        P2_U3210) );
  XNOR2_X1 U10271 ( .A(n8796), .B(n8795), .ZN(n8797) );
  OAI222_X1 U10272 ( .A1(n8928), .A2(n8799), .B1(n8930), .B2(n8798), .C1(n8932), .C2(n8797), .ZN(n8971) );
  INV_X1 U10273 ( .A(n8971), .ZN(n8806) );
  XNOR2_X1 U10274 ( .A(n8800), .B(n8801), .ZN(n8972) );
  AOI22_X1 U10275 ( .A1(n8920), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8937), .B2(
        n8802), .ZN(n8803) );
  OAI21_X1 U10276 ( .B1(n9048), .B2(n8820), .A(n8803), .ZN(n8804) );
  AOI21_X1 U10277 ( .B1(n8972), .B2(n8822), .A(n8804), .ZN(n8805) );
  OAI21_X1 U10278 ( .B1(n8806), .B2(n8920), .A(n8805), .ZN(P2_U3211) );
  XNOR2_X1 U10279 ( .A(n8807), .B(n8814), .ZN(n8811) );
  OAI22_X1 U10280 ( .A1(n8809), .A2(n8928), .B1(n8808), .B2(n8930), .ZN(n8810)
         );
  AOI21_X1 U10281 ( .B1(n8811), .B2(n8914), .A(n8810), .ZN(n8976) );
  NAND2_X1 U10282 ( .A1(n8812), .A2(n8813), .ZN(n8816) );
  INV_X1 U10283 ( .A(n8814), .ZN(n8815) );
  XNOR2_X1 U10284 ( .A(n8816), .B(n8815), .ZN(n8975) );
  INV_X1 U10285 ( .A(n8817), .ZN(n9053) );
  AOI22_X1 U10286 ( .A1(n8920), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8937), .B2(
        n8818), .ZN(n8819) );
  OAI21_X1 U10287 ( .B1(n9053), .B2(n8820), .A(n8819), .ZN(n8821) );
  AOI21_X1 U10288 ( .B1(n8975), .B2(n8822), .A(n8821), .ZN(n8823) );
  OAI21_X1 U10289 ( .B1(n8976), .B2(n8920), .A(n8823), .ZN(P2_U3212) );
  XNOR2_X1 U10290 ( .A(n8824), .B(n8826), .ZN(n9059) );
  INV_X1 U10291 ( .A(n8825), .ZN(n8829) );
  INV_X1 U10292 ( .A(n8826), .ZN(n8828) );
  OAI21_X1 U10293 ( .B1(n8829), .B2(n8828), .A(n8827), .ZN(n8832) );
  AOI222_X1 U10294 ( .A1(n8914), .A2(n8832), .B1(n8831), .B2(n8909), .C1(n8830), .C2(n8911), .ZN(n9054) );
  MUX2_X1 U10295 ( .A(n8833), .B(n9054), .S(n8942), .Z(n8836) );
  AOI22_X1 U10296 ( .A1(n9056), .A2(n8890), .B1(n8937), .B2(n8834), .ZN(n8835)
         );
  OAI211_X1 U10297 ( .C1(n9059), .C2(n8923), .A(n8836), .B(n8835), .ZN(
        P2_U3213) );
  OAI21_X1 U10298 ( .B1(n8838), .B2(n8839), .A(n8837), .ZN(n9065) );
  XOR2_X1 U10299 ( .A(n8840), .B(n8839), .Z(n8842) );
  AOI222_X1 U10300 ( .A1(n8914), .A2(n8842), .B1(n8841), .B2(n8909), .C1(n8864), .C2(n8911), .ZN(n9060) );
  MUX2_X1 U10301 ( .A(n8843), .B(n9060), .S(n8942), .Z(n8847) );
  INV_X1 U10302 ( .A(n8844), .ZN(n8845) );
  AOI22_X1 U10303 ( .A1(n9062), .A2(n8890), .B1(n8937), .B2(n8845), .ZN(n8846)
         );
  OAI211_X1 U10304 ( .C1(n8923), .C2(n9065), .A(n8847), .B(n8846), .ZN(
        P2_U3214) );
  OAI21_X1 U10305 ( .B1(n8850), .B2(n8849), .A(n8848), .ZN(n9069) );
  XNOR2_X1 U10306 ( .A(n8851), .B(n8852), .ZN(n8853) );
  OAI222_X1 U10307 ( .A1(n8930), .A2(n8855), .B1(n8928), .B2(n8854), .C1(n8853), .C2(n8932), .ZN(n8987) );
  NAND2_X1 U10308 ( .A1(n8987), .A2(n8942), .ZN(n8860) );
  INV_X1 U10309 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8857) );
  OAI22_X1 U10310 ( .A1(n8942), .A2(n8857), .B1(n8856), .B2(n8899), .ZN(n8858)
         );
  AOI21_X1 U10311 ( .B1(n8988), .B2(n8890), .A(n8858), .ZN(n8859) );
  OAI211_X1 U10312 ( .C1(n9069), .C2(n8923), .A(n8860), .B(n8859), .ZN(
        P2_U3215) );
  XNOR2_X1 U10313 ( .A(n8861), .B(n8863), .ZN(n9075) );
  XOR2_X1 U10314 ( .A(n8862), .B(n8863), .Z(n8865) );
  AOI222_X1 U10315 ( .A1(n8914), .A2(n8865), .B1(n8885), .B2(n8911), .C1(n8864), .C2(n8909), .ZN(n9070) );
  MUX2_X1 U10316 ( .A(n8866), .B(n9070), .S(n8942), .Z(n8870) );
  INV_X1 U10317 ( .A(n8867), .ZN(n8868) );
  AOI22_X1 U10318 ( .A1(n9072), .A2(n8890), .B1(n8937), .B2(n8868), .ZN(n8869)
         );
  OAI211_X1 U10319 ( .C1(n9075), .C2(n8923), .A(n8870), .B(n8869), .ZN(
        P2_U3216) );
  XOR2_X1 U10320 ( .A(n8873), .B(n8871), .Z(n9081) );
  XOR2_X1 U10321 ( .A(n8872), .B(n8873), .Z(n8875) );
  AOI222_X1 U10322 ( .A1(n8914), .A2(n8875), .B1(n8897), .B2(n8911), .C1(n8874), .C2(n8909), .ZN(n9076) );
  MUX2_X1 U10323 ( .A(n8876), .B(n9076), .S(n8942), .Z(n8880) );
  INV_X1 U10324 ( .A(n8877), .ZN(n8878) );
  AOI22_X1 U10325 ( .A1(n9078), .A2(n8890), .B1(n8937), .B2(n8878), .ZN(n8879)
         );
  OAI211_X1 U10326 ( .C1(n9081), .C2(n8923), .A(n8880), .B(n8879), .ZN(
        P2_U3217) );
  XNOR2_X1 U10327 ( .A(n8882), .B(n8881), .ZN(n9087) );
  XNOR2_X1 U10328 ( .A(n8884), .B(n8883), .ZN(n8886) );
  AOI222_X1 U10329 ( .A1(n8914), .A2(n8886), .B1(n8885), .B2(n8909), .C1(n8910), .C2(n8911), .ZN(n9082) );
  MUX2_X1 U10330 ( .A(n8887), .B(n9082), .S(n8942), .Z(n8892) );
  INV_X1 U10331 ( .A(n8888), .ZN(n8889) );
  AOI22_X1 U10332 ( .A1(n9084), .A2(n8890), .B1(n8937), .B2(n8889), .ZN(n8891)
         );
  OAI211_X1 U10333 ( .C1(n9087), .C2(n8923), .A(n8892), .B(n8891), .ZN(
        P2_U3218) );
  XOR2_X1 U10334 ( .A(n8893), .B(n8895), .Z(n9093) );
  XOR2_X1 U10335 ( .A(n8894), .B(n8895), .Z(n8898) );
  AOI222_X1 U10336 ( .A1(n8914), .A2(n8898), .B1(n8897), .B2(n8909), .C1(n8896), .C2(n8911), .ZN(n9088) );
  INV_X1 U10337 ( .A(n9088), .ZN(n8903) );
  INV_X1 U10338 ( .A(n9090), .ZN(n8901) );
  OAI22_X1 U10339 ( .A1(n8901), .A2(n8915), .B1(n8900), .B2(n8899), .ZN(n8902)
         );
  OAI21_X1 U10340 ( .B1(n8903), .B2(n8902), .A(n8942), .ZN(n8905) );
  NAND2_X1 U10341 ( .A1(n8920), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8904) );
  OAI211_X1 U10342 ( .C1(n9093), .C2(n8923), .A(n8905), .B(n8904), .ZN(
        P2_U3219) );
  XNOR2_X1 U10343 ( .A(n8906), .B(n8908), .ZN(n9101) );
  XNOR2_X1 U10344 ( .A(n8907), .B(n8908), .ZN(n8913) );
  AOI222_X1 U10345 ( .A1(n8914), .A2(n8913), .B1(n8912), .B2(n8911), .C1(n8910), .C2(n8909), .ZN(n9094) );
  OAI21_X1 U10346 ( .B1(n8916), .B2(n8915), .A(n9094), .ZN(n8917) );
  NAND2_X1 U10347 ( .A1(n8917), .A2(n8942), .ZN(n8922) );
  INV_X1 U10348 ( .A(n8918), .ZN(n8919) );
  AOI22_X1 U10349 ( .A1(n8920), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8937), .B2(
        n8919), .ZN(n8921) );
  OAI211_X1 U10350 ( .C1(n9101), .C2(n8923), .A(n8922), .B(n8921), .ZN(
        P2_U3220) );
  NAND2_X1 U10351 ( .A1(n8925), .A2(n8924), .ZN(n8926) );
  NAND2_X1 U10352 ( .A1(n8926), .A2(n7440), .ZN(n10034) );
  INV_X1 U10353 ( .A(n10034), .ZN(n8941) );
  INV_X1 U10354 ( .A(n8927), .ZN(n8936) );
  OAI22_X1 U10355 ( .A1(n6678), .A2(n8930), .B1(n8929), .B2(n8928), .ZN(n8935)
         );
  XNOR2_X1 U10356 ( .A(n8931), .B(n6465), .ZN(n8933) );
  NOR2_X1 U10357 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  AOI211_X1 U10358 ( .C1(n8936), .C2(n10034), .A(n8935), .B(n8934), .ZN(n10036) );
  AOI22_X1 U10359 ( .A1(n10032), .A2(n8938), .B1(n8937), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8939) );
  OAI211_X1 U10360 ( .C1(n8941), .C2(n8940), .A(n10036), .B(n8939), .ZN(n8943)
         );
  MUX2_X1 U10361 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8943), .S(n8942), .Z(
        P2_U3231) );
  NOR2_X1 U10362 ( .A1(n8944), .A2(n10097), .ZN(n8947) );
  AOI21_X1 U10363 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10097), .A(n8947), .ZN(
        n8945) );
  OAI21_X1 U10364 ( .B1(n8946), .B2(n8980), .A(n8945), .ZN(P2_U3490) );
  AOI21_X1 U10365 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10097), .A(n8947), .ZN(
        n8948) );
  OAI21_X1 U10366 ( .B1(n8949), .B2(n8980), .A(n8948), .ZN(P2_U3489) );
  INV_X1 U10367 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U10368 ( .A1(n10097), .A2(n8950), .ZN(n8951) );
  NAND2_X1 U10369 ( .A1(n9016), .A2(n9004), .ZN(n8953) );
  OAI211_X1 U10370 ( .C1(n9019), .C2(n9007), .A(n8954), .B(n8953), .ZN(
        P2_U3487) );
  OAI22_X1 U10371 ( .A1(n8956), .A2(n10080), .B1(n8955), .B2(n10073), .ZN(
        n8957) );
  MUX2_X1 U10372 ( .A(n9020), .B(P2_REG1_REG_27__SCAN_IN), .S(n10097), .Z(
        P2_U3486) );
  INV_X1 U10373 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8959) );
  MUX2_X1 U10374 ( .A(n8959), .B(n9021), .S(n10099), .Z(n8961) );
  NAND2_X1 U10375 ( .A1(n9023), .A2(n9004), .ZN(n8960) );
  OAI211_X1 U10376 ( .C1(n9026), .C2(n9007), .A(n8961), .B(n8960), .ZN(
        P2_U3485) );
  INV_X1 U10377 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8962) );
  MUX2_X1 U10378 ( .A(n8962), .B(n9027), .S(n10099), .Z(n8964) );
  NAND2_X1 U10379 ( .A1(n9029), .A2(n9004), .ZN(n8963) );
  OAI211_X1 U10380 ( .C1(n9032), .C2(n9007), .A(n8964), .B(n8963), .ZN(
        P2_U3484) );
  INV_X1 U10381 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8965) );
  MUX2_X1 U10382 ( .A(n8965), .B(n9033), .S(n10099), .Z(n8967) );
  NAND2_X1 U10383 ( .A1(n9035), .A2(n9004), .ZN(n8966) );
  OAI211_X1 U10384 ( .C1(n9007), .C2(n9038), .A(n8967), .B(n8966), .ZN(
        P2_U3483) );
  INV_X1 U10385 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8968) );
  MUX2_X1 U10386 ( .A(n8968), .B(n9039), .S(n10099), .Z(n8970) );
  NAND2_X1 U10387 ( .A1(n9041), .A2(n9004), .ZN(n8969) );
  OAI211_X1 U10388 ( .C1(n9044), .C2(n9007), .A(n8970), .B(n8969), .ZN(
        P2_U3482) );
  INV_X1 U10389 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8973) );
  AOI21_X1 U10390 ( .B1(n10078), .B2(n8972), .A(n8971), .ZN(n9045) );
  MUX2_X1 U10391 ( .A(n8973), .B(n9045), .S(n10099), .Z(n8974) );
  OAI21_X1 U10392 ( .B1(n9048), .B2(n8980), .A(n8974), .ZN(P2_U3481) );
  INV_X1 U10393 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U10394 ( .A1(n8975), .A2(n10078), .ZN(n8977) );
  AND2_X1 U10395 ( .A1(n8977), .A2(n8976), .ZN(n9049) );
  MUX2_X1 U10396 ( .A(n8978), .B(n9049), .S(n10099), .Z(n8979) );
  OAI21_X1 U10397 ( .B1(n9053), .B2(n8980), .A(n8979), .ZN(P2_U3480) );
  MUX2_X1 U10398 ( .A(n8981), .B(n9054), .S(n10099), .Z(n8983) );
  NAND2_X1 U10399 ( .A1(n9056), .A2(n9004), .ZN(n8982) );
  OAI211_X1 U10400 ( .C1(n9059), .C2(n9007), .A(n8983), .B(n8982), .ZN(
        P2_U3479) );
  MUX2_X1 U10401 ( .A(n8984), .B(n9060), .S(n10099), .Z(n8986) );
  NAND2_X1 U10402 ( .A1(n9062), .A2(n9004), .ZN(n8985) );
  OAI211_X1 U10403 ( .C1(n9065), .C2(n9007), .A(n8986), .B(n8985), .ZN(
        P2_U3478) );
  AOI21_X1 U10404 ( .B1(n10085), .B2(n8988), .A(n8987), .ZN(n9066) );
  MUX2_X1 U10405 ( .A(n8989), .B(n9066), .S(n10099), .Z(n8990) );
  OAI21_X1 U10406 ( .B1(n9007), .B2(n9069), .A(n8990), .ZN(P2_U3477) );
  MUX2_X1 U10407 ( .A(n8991), .B(n9070), .S(n10099), .Z(n8993) );
  NAND2_X1 U10408 ( .A1(n9072), .A2(n9004), .ZN(n8992) );
  OAI211_X1 U10409 ( .C1(n9007), .C2(n9075), .A(n8993), .B(n8992), .ZN(
        P2_U3476) );
  MUX2_X1 U10410 ( .A(n8994), .B(n9076), .S(n10099), .Z(n8996) );
  NAND2_X1 U10411 ( .A1(n9078), .A2(n9004), .ZN(n8995) );
  OAI211_X1 U10412 ( .C1(n9081), .C2(n9007), .A(n8996), .B(n8995), .ZN(
        P2_U3475) );
  MUX2_X1 U10413 ( .A(n8997), .B(n9082), .S(n10099), .Z(n8999) );
  NAND2_X1 U10414 ( .A1(n9084), .A2(n9004), .ZN(n8998) );
  OAI211_X1 U10415 ( .C1(n9007), .C2(n9087), .A(n8999), .B(n8998), .ZN(
        P2_U3474) );
  MUX2_X1 U10416 ( .A(n9000), .B(n9088), .S(n10099), .Z(n9002) );
  NAND2_X1 U10417 ( .A1(n9090), .A2(n9004), .ZN(n9001) );
  OAI211_X1 U10418 ( .C1(n9007), .C2(n9093), .A(n9002), .B(n9001), .ZN(
        P2_U3473) );
  MUX2_X1 U10419 ( .A(n9003), .B(n9094), .S(n10099), .Z(n9006) );
  NAND2_X1 U10420 ( .A1(n9097), .A2(n9004), .ZN(n9005) );
  OAI211_X1 U10421 ( .C1(n9007), .C2(n9101), .A(n9006), .B(n9005), .ZN(
        P2_U3472) );
  NAND2_X1 U10422 ( .A1(n9008), .A2(n9096), .ZN(n9010) );
  NAND2_X1 U10423 ( .A1(n9009), .A2(n10086), .ZN(n9012) );
  OAI211_X1 U10424 ( .C1(n6103), .C2(n10086), .A(n9010), .B(n9012), .ZN(
        P2_U3458) );
  NAND2_X1 U10425 ( .A1(n9011), .A2(n9096), .ZN(n9013) );
  OAI211_X1 U10426 ( .C1(n6109), .C2(n10086), .A(n9013), .B(n9012), .ZN(
        P2_U3457) );
  MUX2_X1 U10427 ( .A(n9015), .B(n9014), .S(n10086), .Z(n9018) );
  NAND2_X1 U10428 ( .A1(n9016), .A2(n9096), .ZN(n9017) );
  OAI211_X1 U10429 ( .C1(n9019), .C2(n9100), .A(n9018), .B(n9017), .ZN(
        P2_U3455) );
  MUX2_X1 U10430 ( .A(n9020), .B(P2_REG0_REG_27__SCAN_IN), .S(n10087), .Z(
        P2_U3454) );
  MUX2_X1 U10431 ( .A(n9022), .B(n9021), .S(n10086), .Z(n9025) );
  NAND2_X1 U10432 ( .A1(n9023), .A2(n9096), .ZN(n9024) );
  OAI211_X1 U10433 ( .C1(n9026), .C2(n9100), .A(n9025), .B(n9024), .ZN(
        P2_U3453) );
  MUX2_X1 U10434 ( .A(n9028), .B(n9027), .S(n10086), .Z(n9031) );
  NAND2_X1 U10435 ( .A1(n9029), .A2(n9096), .ZN(n9030) );
  OAI211_X1 U10436 ( .C1(n9032), .C2(n9100), .A(n9031), .B(n9030), .ZN(
        P2_U3452) );
  MUX2_X1 U10437 ( .A(n9034), .B(n9033), .S(n10086), .Z(n9037) );
  NAND2_X1 U10438 ( .A1(n9035), .A2(n9096), .ZN(n9036) );
  OAI211_X1 U10439 ( .C1(n9038), .C2(n9100), .A(n9037), .B(n9036), .ZN(
        P2_U3451) );
  INV_X1 U10440 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9040) );
  MUX2_X1 U10441 ( .A(n9040), .B(n9039), .S(n10086), .Z(n9043) );
  NAND2_X1 U10442 ( .A1(n9041), .A2(n9096), .ZN(n9042) );
  OAI211_X1 U10443 ( .C1(n9044), .C2(n9100), .A(n9043), .B(n9042), .ZN(
        P2_U3450) );
  INV_X1 U10444 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9046) );
  MUX2_X1 U10445 ( .A(n9046), .B(n9045), .S(n10086), .Z(n9047) );
  OAI21_X1 U10446 ( .B1(n9048), .B2(n9052), .A(n9047), .ZN(P2_U3449) );
  INV_X1 U10447 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9050) );
  MUX2_X1 U10448 ( .A(n9050), .B(n9049), .S(n10086), .Z(n9051) );
  OAI21_X1 U10449 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(P2_U3448) );
  MUX2_X1 U10450 ( .A(n9055), .B(n9054), .S(n10086), .Z(n9058) );
  NAND2_X1 U10451 ( .A1(n9056), .A2(n9096), .ZN(n9057) );
  OAI211_X1 U10452 ( .C1(n9059), .C2(n9100), .A(n9058), .B(n9057), .ZN(
        P2_U3447) );
  INV_X1 U10453 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9061) );
  MUX2_X1 U10454 ( .A(n9061), .B(n9060), .S(n10086), .Z(n9064) );
  NAND2_X1 U10455 ( .A1(n9062), .A2(n9096), .ZN(n9063) );
  OAI211_X1 U10456 ( .C1(n9065), .C2(n9100), .A(n9064), .B(n9063), .ZN(
        P2_U3446) );
  MUX2_X1 U10457 ( .A(n9067), .B(n9066), .S(n10086), .Z(n9068) );
  OAI21_X1 U10458 ( .B1(n9069), .B2(n9100), .A(n9068), .ZN(P2_U3444) );
  INV_X1 U10459 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9071) );
  MUX2_X1 U10460 ( .A(n9071), .B(n9070), .S(n10086), .Z(n9074) );
  NAND2_X1 U10461 ( .A1(n9072), .A2(n9096), .ZN(n9073) );
  OAI211_X1 U10462 ( .C1(n9075), .C2(n9100), .A(n9074), .B(n9073), .ZN(
        P2_U3441) );
  INV_X1 U10463 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9077) );
  MUX2_X1 U10464 ( .A(n9077), .B(n9076), .S(n10086), .Z(n9080) );
  NAND2_X1 U10465 ( .A1(n9078), .A2(n9096), .ZN(n9079) );
  OAI211_X1 U10466 ( .C1(n9081), .C2(n9100), .A(n9080), .B(n9079), .ZN(
        P2_U3438) );
  INV_X1 U10467 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9083) );
  MUX2_X1 U10468 ( .A(n9083), .B(n9082), .S(n10086), .Z(n9086) );
  NAND2_X1 U10469 ( .A1(n9084), .A2(n9096), .ZN(n9085) );
  OAI211_X1 U10470 ( .C1(n9087), .C2(n9100), .A(n9086), .B(n9085), .ZN(
        P2_U3435) );
  INV_X1 U10471 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9089) );
  MUX2_X1 U10472 ( .A(n9089), .B(n9088), .S(n10086), .Z(n9092) );
  NAND2_X1 U10473 ( .A1(n9090), .A2(n9096), .ZN(n9091) );
  OAI211_X1 U10474 ( .C1(n9093), .C2(n9100), .A(n9092), .B(n9091), .ZN(
        P2_U3432) );
  INV_X1 U10475 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9095) );
  MUX2_X1 U10476 ( .A(n9095), .B(n9094), .S(n10086), .Z(n9099) );
  NAND2_X1 U10477 ( .A1(n9097), .A2(n9096), .ZN(n9098) );
  OAI211_X1 U10478 ( .C1(n9101), .C2(n9100), .A(n9099), .B(n9098), .ZN(
        P2_U3429) );
  MUX2_X1 U10479 ( .A(n9103), .B(P2_D_REG_1__SCAN_IN), .S(n9102), .Z(P2_U3377)
         );
  NAND3_X1 U10480 ( .A1(n6094), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9107) );
  OAI22_X1 U10481 ( .A1(n9104), .A2(n9107), .B1(n9106), .B2(n9105), .ZN(n9108)
         );
  AOI21_X1 U10482 ( .B1(n6066), .B2(n9109), .A(n9108), .ZN(n9110) );
  INV_X1 U10483 ( .A(n9110), .ZN(P2_U3264) );
  INV_X1 U10484 ( .A(n6132), .ZN(n9878) );
  AOI21_X1 U10485 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9115), .A(n9111), .ZN(
        n9112) );
  OAI21_X1 U10486 ( .B1(n9878), .B2(n9117), .A(n9112), .ZN(P2_U3267) );
  INV_X1 U10487 ( .A(n9113), .ZN(n9879) );
  AOI21_X1 U10488 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n9115), .A(n9114), .ZN(
        n9116) );
  OAI21_X1 U10489 ( .B1(n9879), .B2(n9117), .A(n9116), .ZN(P2_U3268) );
  INV_X1 U10490 ( .A(n9118), .ZN(n9880) );
  OAI222_X1 U10491 ( .A1(n9117), .A2(n9880), .B1(P2_U3151), .B2(n9120), .C1(
        n9119), .C2(n9122), .ZN(P2_U3269) );
  INV_X1 U10492 ( .A(n9121), .ZN(n9883) );
  OAI222_X1 U10493 ( .A1(n9117), .A2(n9883), .B1(P2_U3151), .B2(n5078), .C1(
        n9123), .C2(n9122), .ZN(P2_U3270) );
  INV_X1 U10494 ( .A(n9124), .ZN(n9125) );
  MUX2_X1 U10495 ( .A(n9125), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10496 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  XOR2_X1 U10497 ( .A(n9129), .B(n9128), .Z(n9136) );
  OAI22_X1 U10498 ( .A1(n9923), .A2(n9131), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9130), .ZN(n9133) );
  OAI22_X1 U10499 ( .A1(n9179), .A2(n9279), .B1(n9890), .B2(n9199), .ZN(n9132)
         );
  AOI211_X1 U10500 ( .C1(n9134), .C2(n9920), .A(n9133), .B(n9132), .ZN(n9135)
         );
  OAI21_X1 U10501 ( .B1(n9136), .B2(n9916), .A(n9135), .ZN(P1_U3215) );
  AOI21_X1 U10502 ( .B1(n9137), .B2(n4549), .A(n4520), .ZN(n9142) );
  OAI22_X1 U10503 ( .A1(n9923), .A2(n9591), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9138), .ZN(n9140) );
  OAI22_X1 U10504 ( .A1(n9585), .A2(n9890), .B1(n9584), .B2(n9279), .ZN(n9139)
         );
  AOI211_X1 U10505 ( .C1(n9590), .C2(n9920), .A(n9140), .B(n9139), .ZN(n9141)
         );
  OAI21_X1 U10506 ( .B1(n9142), .B2(n9916), .A(n9141), .ZN(P1_U3216) );
  NAND2_X1 U10507 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9470) );
  OAI21_X1 U10508 ( .B1(n9923), .B2(n9653), .A(n9470), .ZN(n9145) );
  OAI22_X1 U10509 ( .A1(n9661), .A2(n9279), .B1(n9890), .B2(n9663), .ZN(n9144)
         );
  AOI211_X1 U10510 ( .C1(n9798), .C2(n9920), .A(n9145), .B(n9144), .ZN(n9146)
         );
  OAI21_X1 U10511 ( .B1(n9147), .B2(n9916), .A(n9146), .ZN(P1_U3219) );
  NAND2_X1 U10512 ( .A1(n9752), .A2(n9148), .ZN(n9151) );
  NAND2_X1 U10513 ( .A1(n9287), .A2(n9149), .ZN(n9150) );
  NAND2_X1 U10514 ( .A1(n9151), .A2(n9150), .ZN(n9153) );
  XNOR2_X1 U10515 ( .A(n9153), .B(n9152), .ZN(n9156) );
  NAND2_X1 U10516 ( .A1(n9752), .A2(n8233), .ZN(n9154) );
  OAI21_X1 U10517 ( .B1(n9525), .B2(n8284), .A(n9154), .ZN(n9155) );
  XNOR2_X1 U10518 ( .A(n9156), .B(n9155), .ZN(n9162) );
  OAI22_X1 U10519 ( .A1(n9923), .A2(n9510), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9157), .ZN(n9160) );
  OAI22_X1 U10520 ( .A1(n9537), .A2(n9279), .B1(n9890), .B2(n9158), .ZN(n9159)
         );
  AOI211_X1 U10521 ( .C1(n9752), .C2(n9920), .A(n9160), .B(n9159), .ZN(n9163)
         );
  XOR2_X1 U10522 ( .A(n9166), .B(n9165), .Z(n9167) );
  XNOR2_X1 U10523 ( .A(n9164), .B(n9167), .ZN(n9172) );
  NOR2_X1 U10524 ( .A1(n9923), .A2(n9627), .ZN(n9170) );
  AOI22_X1 U10525 ( .A1(n9290), .A2(n9728), .B1(n9727), .B2(n9291), .ZN(n9623)
         );
  OAI22_X1 U10526 ( .A1(n9623), .A2(n9911), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9168), .ZN(n9169) );
  AOI211_X1 U10527 ( .C1(n9626), .C2(n9920), .A(n9170), .B(n9169), .ZN(n9171)
         );
  OAI21_X1 U10528 ( .B1(n9172), .B2(n9916), .A(n9171), .ZN(P1_U3223) );
  INV_X1 U10529 ( .A(n9173), .ZN(n9177) );
  NOR3_X1 U10530 ( .A1(n4581), .A2(n9175), .A3(n9174), .ZN(n9176) );
  OAI21_X1 U10531 ( .B1(n9177), .B2(n9176), .A(n9906), .ZN(n9185) );
  INV_X1 U10532 ( .A(n9178), .ZN(n9183) );
  OAI22_X1 U10533 ( .A1(n9180), .A2(n9279), .B1(n9890), .B2(n9179), .ZN(n9181)
         );
  AOI211_X1 U10534 ( .C1(n9269), .C2(n9183), .A(n9182), .B(n9181), .ZN(n9184)
         );
  OAI211_X1 U10535 ( .C1(n6024), .C2(n9903), .A(n9185), .B(n9184), .ZN(
        P1_U3224) );
  OAI21_X1 U10536 ( .B1(n9188), .B2(n9187), .A(n9186), .ZN(n9192) );
  OAI22_X1 U10537 ( .A1(n9585), .A2(n9662), .B1(n9524), .B2(n9664), .ZN(n9552)
         );
  AOI22_X1 U10538 ( .A1(n9552), .A2(n9900), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9190) );
  NAND2_X1 U10539 ( .A1(n9558), .A2(n9269), .ZN(n9189) );
  OAI211_X1 U10540 ( .C1(n9838), .C2(n9903), .A(n9190), .B(n9189), .ZN(n9191)
         );
  AOI21_X1 U10541 ( .B1(n9192), .B2(n9906), .A(n9191), .ZN(n9193) );
  INV_X1 U10542 ( .A(n9193), .ZN(P1_U3225) );
  NAND2_X1 U10543 ( .A1(n9195), .A2(n9194), .ZN(n9196) );
  XNOR2_X1 U10544 ( .A(n9197), .B(n9196), .ZN(n9203) );
  INV_X1 U10545 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9198) );
  OAI22_X1 U10546 ( .A1(n9923), .A2(n9712), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9198), .ZN(n9201) );
  OAI22_X1 U10547 ( .A1(n9199), .A2(n9279), .B1(n9890), .B2(n9256), .ZN(n9200)
         );
  AOI211_X1 U10548 ( .C1(n9812), .C2(n9920), .A(n9201), .B(n9200), .ZN(n9202)
         );
  OAI21_X1 U10549 ( .B1(n9203), .B2(n9916), .A(n9202), .ZN(P1_U3226) );
  NAND2_X1 U10550 ( .A1(n9206), .A2(n9205), .ZN(n9207) );
  XNOR2_X1 U10551 ( .A(n9204), .B(n9207), .ZN(n9214) );
  NOR2_X1 U10552 ( .A1(n9923), .A2(n9691), .ZN(n9212) );
  NAND2_X1 U10553 ( .A1(n4793), .A2(n9727), .ZN(n9209) );
  NAND2_X1 U10554 ( .A1(n9293), .A2(n9728), .ZN(n9208) );
  AND2_X1 U10555 ( .A1(n9209), .A2(n9208), .ZN(n9686) );
  OAI21_X1 U10556 ( .B1(n9686), .B2(n9911), .A(n9210), .ZN(n9211) );
  AOI211_X1 U10557 ( .C1(n9690), .C2(n9920), .A(n9212), .B(n9211), .ZN(n9213)
         );
  OAI21_X1 U10558 ( .B1(n9214), .B2(n9916), .A(n9213), .ZN(P1_U3228) );
  OAI21_X1 U10559 ( .B1(n9217), .B2(n4558), .A(n9906), .ZN(n9222) );
  NOR2_X1 U10560 ( .A1(n9218), .A2(n9923), .ZN(n9220) );
  OAI22_X1 U10561 ( .A1(n9570), .A2(n9890), .B1(n9569), .B2(n9279), .ZN(n9219)
         );
  AOI211_X1 U10562 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n9220), 
        .B(n9219), .ZN(n9221) );
  OAI211_X1 U10563 ( .C1(n9576), .C2(n9903), .A(n9222), .B(n9221), .ZN(
        P1_U3229) );
  NAND2_X1 U10564 ( .A1(n9224), .A2(n9223), .ZN(n9226) );
  XOR2_X1 U10565 ( .A(n9226), .B(n9225), .Z(n9231) );
  INV_X1 U10566 ( .A(n9641), .ZN(n9228) );
  OAI22_X1 U10567 ( .A1(n9246), .A2(n9664), .B1(n9292), .B2(n9662), .ZN(n9638)
         );
  AOI22_X1 U10568 ( .A1(n9638), .A2(n9900), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9227) );
  OAI21_X1 U10569 ( .B1(n9228), .B2(n9923), .A(n9227), .ZN(n9229) );
  AOI21_X1 U10570 ( .B1(n9643), .B2(n9920), .A(n9229), .ZN(n9230) );
  OAI21_X1 U10571 ( .B1(n9231), .B2(n9916), .A(n9230), .ZN(P1_U3233) );
  OAI21_X1 U10572 ( .B1(n9234), .B2(n9233), .A(n9232), .ZN(n9235) );
  NAND2_X1 U10573 ( .A1(n9235), .A2(n9906), .ZN(n9239) );
  AND2_X1 U10574 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9406) );
  OAI22_X1 U10575 ( .A1(n9280), .A2(n9890), .B1(n9279), .B2(n6023), .ZN(n9236)
         );
  AOI211_X1 U10576 ( .C1(n9237), .C2(n9269), .A(n9406), .B(n9236), .ZN(n9238)
         );
  OAI211_X1 U10577 ( .C1(n9240), .C2(n9903), .A(n9239), .B(n9238), .ZN(
        P1_U3234) );
  XOR2_X1 U10578 ( .A(n9242), .B(n9241), .Z(n9243) );
  XNOR2_X1 U10579 ( .A(n9244), .B(n9243), .ZN(n9250) );
  OAI22_X1 U10580 ( .A1(n9923), .A2(n9602), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9245), .ZN(n9248) );
  OAI22_X1 U10581 ( .A1(n9569), .A2(n9890), .B1(n9246), .B2(n9279), .ZN(n9247)
         );
  AOI211_X1 U10582 ( .C1(n9782), .C2(n9920), .A(n9248), .B(n9247), .ZN(n9249)
         );
  OAI21_X1 U10583 ( .B1(n9250), .B2(n9916), .A(n9249), .ZN(P1_U3235) );
  NAND2_X1 U10584 ( .A1(n9252), .A2(n9251), .ZN(n9254) );
  XNOR2_X1 U10585 ( .A(n9254), .B(n9253), .ZN(n9260) );
  OAI22_X1 U10586 ( .A1(n9923), .A2(n9671), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9255), .ZN(n9258) );
  OAI22_X1 U10587 ( .A1(n9256), .A2(n9279), .B1(n9890), .B2(n9292), .ZN(n9257)
         );
  AOI211_X1 U10588 ( .C1(n4719), .C2(n9920), .A(n9258), .B(n9257), .ZN(n9259)
         );
  OAI21_X1 U10589 ( .B1(n9260), .B2(n9916), .A(n9259), .ZN(P1_U3238) );
  INV_X1 U10590 ( .A(n9186), .ZN(n9263) );
  OAI21_X1 U10591 ( .B1(n9263), .B2(n9262), .A(n9261), .ZN(n9265) );
  NAND3_X1 U10592 ( .A1(n9265), .A2(n9906), .A3(n9264), .ZN(n9271) );
  NOR2_X1 U10593 ( .A1(n9266), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9268) );
  OAI22_X1 U10594 ( .A1(n9570), .A2(n9279), .B1(n9537), .B2(n9890), .ZN(n9267)
         );
  AOI211_X1 U10595 ( .C1(n9269), .C2(n9541), .A(n9268), .B(n9267), .ZN(n9270)
         );
  OAI211_X1 U10596 ( .C1(n9544), .C2(n9903), .A(n9271), .B(n9270), .ZN(
        P1_U3240) );
  INV_X1 U10597 ( .A(n9272), .ZN(n9274) );
  NOR2_X1 U10598 ( .A1(n9274), .A2(n9273), .ZN(n9276) );
  XNOR2_X1 U10599 ( .A(n9276), .B(n9275), .ZN(n9284) );
  OAI22_X1 U10600 ( .A1(n9923), .A2(n9735), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9277), .ZN(n9282) );
  OAI22_X1 U10601 ( .A1(n9280), .A2(n9279), .B1(n9890), .B2(n9278), .ZN(n9281)
         );
  AOI211_X1 U10602 ( .C1(n9734), .C2(n9920), .A(n9282), .B(n9281), .ZN(n9283)
         );
  OAI21_X1 U10603 ( .B1(n9284), .B2(n9916), .A(n9283), .ZN(P1_U3241) );
  MUX2_X1 U10604 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9285), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10605 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9286), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10606 ( .A(n9499), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9306), .Z(
        P1_U3583) );
  MUX2_X1 U10607 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9287), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10608 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9498), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10609 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9288), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10610 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9289), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10611 ( .A(n9609), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9306), .Z(
        P1_U3577) );
  MUX2_X1 U10612 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9290), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10613 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9610), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10614 ( .A(n9291), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9306), .Z(
        P1_U3574) );
  INV_X1 U10615 ( .A(n9292), .ZN(n9677) );
  MUX2_X1 U10616 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9677), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10617 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9293), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10618 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9702), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10619 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n4793), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10620 ( .A(n9701), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9306), .Z(
        P1_U3569) );
  MUX2_X1 U10621 ( .A(n9726), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9306), .Z(
        P1_U3568) );
  MUX2_X1 U10622 ( .A(n9294), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9306), .Z(
        P1_U3567) );
  MUX2_X1 U10623 ( .A(n9295), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9306), .Z(
        P1_U3566) );
  MUX2_X1 U10624 ( .A(n9296), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9306), .Z(
        P1_U3565) );
  MUX2_X1 U10625 ( .A(n9297), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9306), .Z(
        P1_U3564) );
  MUX2_X1 U10626 ( .A(n9298), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9306), .Z(
        P1_U3563) );
  MUX2_X1 U10627 ( .A(n9299), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9306), .Z(
        P1_U3562) );
  MUX2_X1 U10628 ( .A(n9300), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9306), .Z(
        P1_U3561) );
  MUX2_X1 U10629 ( .A(n9301), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9306), .Z(
        P1_U3560) );
  MUX2_X1 U10630 ( .A(n9302), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9306), .Z(
        P1_U3559) );
  MUX2_X1 U10631 ( .A(n9303), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9306), .Z(
        P1_U3558) );
  MUX2_X1 U10632 ( .A(n9304), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9306), .Z(
        P1_U3557) );
  MUX2_X1 U10633 ( .A(n9305), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9306), .Z(
        P1_U3556) );
  MUX2_X1 U10634 ( .A(n4512), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9306), .Z(
        P1_U3555) );
  MUX2_X1 U10635 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n7038), .S(P1_U3973), .Z(
        P1_U3554) );
  INV_X1 U10636 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10101) );
  INV_X1 U10637 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9307) );
  OAI22_X1 U10638 ( .A1(n9472), .A2(n10101), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9307), .ZN(n9308) );
  AOI21_X1 U10639 ( .B1(n9309), .B2(n9373), .A(n9308), .ZN(n9318) );
  OAI211_X1 U10640 ( .C1(n9312), .C2(n9311), .A(n9439), .B(n9310), .ZN(n9317)
         );
  OAI211_X1 U10641 ( .C1(n9315), .C2(n9314), .A(n9445), .B(n9313), .ZN(n9316)
         );
  NAND3_X1 U10642 ( .A1(n9318), .A2(n9317), .A3(n9316), .ZN(P1_U3244) );
  OAI211_X1 U10643 ( .C1(n9321), .C2(n9320), .A(n9445), .B(n9319), .ZN(n9333)
         );
  MUX2_X1 U10644 ( .A(n6891), .B(P1_REG1_REG_3__SCAN_IN), .S(n9327), .Z(n9323)
         );
  NAND3_X1 U10645 ( .A1(n9324), .A2(n9323), .A3(n9322), .ZN(n9325) );
  NAND3_X1 U10646 ( .A1(n9439), .A2(n9326), .A3(n9325), .ZN(n9332) );
  NAND2_X1 U10647 ( .A1(n9373), .A2(n9327), .ZN(n9331) );
  NOR2_X1 U10648 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9328), .ZN(n9329) );
  AOI21_X1 U10649 ( .B1(n9933), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9329), .ZN(
        n9330) );
  NAND4_X1 U10650 ( .A1(n9333), .A2(n9332), .A3(n9331), .A4(n9330), .ZN(
        P1_U3246) );
  INV_X1 U10651 ( .A(n9334), .ZN(n9337) );
  NOR2_X1 U10652 ( .A1(n9459), .A2(n9335), .ZN(n9336) );
  AOI211_X1 U10653 ( .C1(n9933), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9337), .B(
        n9336), .ZN(n9347) );
  OAI211_X1 U10654 ( .C1(n9340), .C2(n9339), .A(n9445), .B(n9338), .ZN(n9346)
         );
  NAND3_X1 U10655 ( .A1(n9343), .A2(n9342), .A3(n9341), .ZN(n9344) );
  NAND3_X1 U10656 ( .A1(n9439), .A2(n9356), .A3(n9344), .ZN(n9345) );
  NAND3_X1 U10657 ( .A1(n9347), .A2(n9346), .A3(n9345), .ZN(P1_U3248) );
  NOR2_X1 U10658 ( .A1(n9459), .A2(n9348), .ZN(n9349) );
  AOI211_X1 U10659 ( .C1(n9933), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9350), .B(
        n9349), .ZN(n9361) );
  OAI211_X1 U10660 ( .C1(n9353), .C2(n9352), .A(n9445), .B(n9351), .ZN(n9360)
         );
  INV_X1 U10661 ( .A(n9370), .ZN(n9358) );
  NAND3_X1 U10662 ( .A1(n9356), .A2(n9355), .A3(n9354), .ZN(n9357) );
  NAND3_X1 U10663 ( .A1(n9439), .A2(n9358), .A3(n9357), .ZN(n9359) );
  NAND3_X1 U10664 ( .A1(n9361), .A2(n9360), .A3(n9359), .ZN(P1_U3249) );
  OAI211_X1 U10665 ( .C1(n9364), .C2(n9363), .A(n9445), .B(n9362), .ZN(n9377)
         );
  MUX2_X1 U10666 ( .A(n6899), .B(P1_REG1_REG_7__SCAN_IN), .S(n9372), .Z(n9367)
         );
  INV_X1 U10667 ( .A(n9365), .ZN(n9366) );
  NAND2_X1 U10668 ( .A1(n9367), .A2(n9366), .ZN(n9369) );
  OAI211_X1 U10669 ( .C1(n9370), .C2(n9369), .A(n9439), .B(n9368), .ZN(n9376)
         );
  AOI21_X1 U10670 ( .B1(n9933), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9371), .ZN(
        n9375) );
  NAND2_X1 U10671 ( .A1(n9373), .A2(n9372), .ZN(n9374) );
  NAND4_X1 U10672 ( .A1(n9377), .A2(n9376), .A3(n9375), .A4(n9374), .ZN(
        P1_U3250) );
  NOR2_X1 U10673 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9378), .ZN(n9899) );
  NOR2_X1 U10674 ( .A1(n9459), .A2(n9379), .ZN(n9380) );
  AOI211_X1 U10675 ( .C1(n9933), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n9899), .B(
        n9380), .ZN(n9390) );
  AOI211_X1 U10676 ( .C1(n9383), .C2(n9382), .A(n9381), .B(n9465), .ZN(n9384)
         );
  INV_X1 U10677 ( .A(n9384), .ZN(n9389) );
  OAI211_X1 U10678 ( .C1(n9387), .C2(n9386), .A(n9439), .B(n9385), .ZN(n9388)
         );
  NAND3_X1 U10679 ( .A1(n9390), .A2(n9389), .A3(n9388), .ZN(P1_U3253) );
  NOR2_X1 U10680 ( .A1(n9459), .A2(n9391), .ZN(n9392) );
  AOI211_X1 U10681 ( .C1(n9933), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9393), .B(
        n9392), .ZN(n9403) );
  OAI211_X1 U10682 ( .C1(n9396), .C2(n9395), .A(n9439), .B(n9394), .ZN(n9402)
         );
  AOI211_X1 U10683 ( .C1(n9399), .C2(n9398), .A(n9397), .B(n9465), .ZN(n9400)
         );
  INV_X1 U10684 ( .A(n9400), .ZN(n9401) );
  NAND3_X1 U10685 ( .A1(n9403), .A2(n9402), .A3(n9401), .ZN(P1_U3254) );
  NOR2_X1 U10686 ( .A1(n9459), .A2(n9404), .ZN(n9405) );
  AOI211_X1 U10687 ( .C1(n9933), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n9406), .B(
        n9405), .ZN(n9416) );
  OAI211_X1 U10688 ( .C1(n9409), .C2(n9408), .A(n9439), .B(n9407), .ZN(n9415)
         );
  AOI211_X1 U10689 ( .C1(n9412), .C2(n9411), .A(n9410), .B(n9465), .ZN(n9413)
         );
  INV_X1 U10690 ( .A(n9413), .ZN(n9414) );
  NAND3_X1 U10691 ( .A1(n9416), .A2(n9415), .A3(n9414), .ZN(P1_U3256) );
  AND2_X1 U10692 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9419) );
  NOR2_X1 U10693 ( .A1(n9459), .A2(n9417), .ZN(n9418) );
  AOI211_X1 U10694 ( .C1(n9933), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9419), .B(
        n9418), .ZN(n9429) );
  OAI211_X1 U10695 ( .C1(n9422), .C2(n9421), .A(n9439), .B(n9420), .ZN(n9428)
         );
  AOI211_X1 U10696 ( .C1(n9425), .C2(n9424), .A(n9423), .B(n9465), .ZN(n9426)
         );
  INV_X1 U10697 ( .A(n9426), .ZN(n9427) );
  NAND3_X1 U10698 ( .A1(n9429), .A2(n9428), .A3(n9427), .ZN(P1_U3257) );
  AND2_X1 U10699 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9432) );
  NOR2_X1 U10700 ( .A1(n9459), .A2(n9430), .ZN(n9431) );
  AOI211_X1 U10701 ( .C1(n9933), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9432), .B(
        n9431), .ZN(n9450) );
  OR2_X1 U10702 ( .A1(n9433), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U10703 ( .A1(n9435), .A2(n9434), .ZN(n9437) );
  XNOR2_X1 U10704 ( .A(n9454), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U10705 ( .A1(n9437), .A2(n9436), .ZN(n9438) );
  NAND3_X1 U10706 ( .A1(n9439), .A2(n9456), .A3(n9438), .ZN(n9449) );
  INV_X1 U10707 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9442) );
  OR2_X1 U10708 ( .A1(n9454), .A2(n9442), .ZN(n9444) );
  NAND2_X1 U10709 ( .A1(n9454), .A2(n9442), .ZN(n9443) );
  NAND2_X1 U10710 ( .A1(n9444), .A2(n9443), .ZN(n9446) );
  NAND2_X1 U10711 ( .A1(n9447), .A2(n9446), .ZN(n9452) );
  OAI211_X1 U10712 ( .C1(n9447), .C2(n9446), .A(n9445), .B(n9452), .ZN(n9448)
         );
  NAND3_X1 U10713 ( .A1(n9450), .A2(n9449), .A3(n9448), .ZN(P1_U3261) );
  NAND2_X1 U10714 ( .A1(n9454), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U10715 ( .A1(n9452), .A2(n9451), .ZN(n9453) );
  XNOR2_X1 U10716 ( .A(n9453), .B(n9654), .ZN(n9461) );
  NAND2_X1 U10717 ( .A1(n9454), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U10718 ( .A1(n9456), .A2(n9455), .ZN(n9458) );
  XNOR2_X1 U10719 ( .A(n9458), .B(n9457), .ZN(n9462) );
  OR2_X1 U10720 ( .A1(n9464), .A2(n9462), .ZN(n9460) );
  OAI211_X1 U10721 ( .C1(n9465), .C2(n9461), .A(n9460), .B(n9459), .ZN(n9468)
         );
  INV_X1 U10722 ( .A(n9461), .ZN(n9466) );
  INV_X1 U10723 ( .A(n9462), .ZN(n9463) );
  OAI22_X1 U10724 ( .A1(n9466), .A2(n9465), .B1(n9464), .B2(n9463), .ZN(n9467)
         );
  MUX2_X1 U10725 ( .A(n9468), .B(n9467), .S(n7033), .Z(n9469) );
  INV_X1 U10726 ( .A(n9469), .ZN(n9471) );
  OAI211_X1 U10727 ( .C1(n9473), .C2(n9472), .A(n9471), .B(n9470), .ZN(
        P1_U3262) );
  NOR2_X1 U10728 ( .A1(n9612), .A2(n9746), .ZN(n9479) );
  NOR2_X1 U10729 ( .A1(n9745), .A2(n9945), .ZN(n9474) );
  AOI211_X1 U10730 ( .C1(n9612), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9479), .B(
        n9474), .ZN(n9475) );
  OAI21_X1 U10731 ( .B1(n9476), .B2(n9646), .A(n9475), .ZN(P1_U3263) );
  OAI211_X1 U10732 ( .C1(n9828), .C2(n9478), .A(n9813), .B(n9477), .ZN(n9747)
         );
  NAND2_X1 U10733 ( .A1(n9612), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9481) );
  INV_X1 U10734 ( .A(n9479), .ZN(n9480) );
  OAI211_X1 U10735 ( .C1(n9828), .C2(n9945), .A(n9481), .B(n9480), .ZN(n9482)
         );
  INV_X1 U10736 ( .A(n9482), .ZN(n9483) );
  OAI21_X1 U10737 ( .B1(n9747), .B2(n9646), .A(n9483), .ZN(P1_U3264) );
  INV_X1 U10738 ( .A(n9484), .ZN(n9495) );
  INV_X1 U10739 ( .A(n9485), .ZN(n9486) );
  AOI22_X1 U10740 ( .A1(n9612), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9486), .B2(
        n9942), .ZN(n9489) );
  NAND2_X1 U10741 ( .A1(n9487), .A2(n9642), .ZN(n9488) );
  OAI211_X1 U10742 ( .C1(n9491), .C2(n9490), .A(n9489), .B(n9488), .ZN(n9492)
         );
  AOI21_X1 U10743 ( .B1(n9493), .B2(n9714), .A(n9492), .ZN(n9494) );
  OAI21_X1 U10744 ( .B1(n9495), .B2(n9741), .A(n9494), .ZN(P1_U3356) );
  NAND2_X1 U10745 ( .A1(n9499), .A2(n9728), .ZN(n9500) );
  NAND2_X1 U10746 ( .A1(n9504), .A2(n9503), .ZN(n9506) );
  NAND2_X1 U10747 ( .A1(n9506), .A2(n9505), .ZN(n9507) );
  NAND2_X1 U10748 ( .A1(n9750), .A2(n9707), .ZN(n9515) );
  AOI211_X1 U10749 ( .C1(n9752), .C2(n9516), .A(n9969), .B(n9509), .ZN(n9751)
         );
  NOR2_X1 U10750 ( .A1(n4707), .A2(n9945), .ZN(n9513) );
  OAI22_X1 U10751 ( .A1(n9714), .A2(n9511), .B1(n9510), .B2(n9711), .ZN(n9512)
         );
  AOI211_X1 U10752 ( .C1(n9751), .C2(n9950), .A(n9513), .B(n9512), .ZN(n9514)
         );
  OAI211_X1 U10753 ( .C1(n9612), .C2(n9754), .A(n9515), .B(n9514), .ZN(
        P1_U3265) );
  AOI21_X1 U10754 ( .B1(n9529), .B2(n9538), .A(n9969), .ZN(n9517) );
  NOR2_X1 U10755 ( .A1(n9711), .A2(n9518), .ZN(n9526) );
  INV_X1 U10756 ( .A(n9519), .ZN(n9522) );
  NOR3_X1 U10757 ( .A1(n4541), .A2(n9520), .A3(n9527), .ZN(n9521) );
  OAI222_X1 U10758 ( .A1(n9664), .A2(n9525), .B1(n9662), .B2(n9524), .C1(n9659), .C2(n9523), .ZN(n9756) );
  AOI211_X1 U10759 ( .C1(n9757), .C2(n7033), .A(n9526), .B(n9756), .ZN(n9532)
         );
  XNOR2_X1 U10760 ( .A(n9528), .B(n9527), .ZN(n9758) );
  NAND2_X1 U10761 ( .A1(n9758), .A2(n9707), .ZN(n9531) );
  AOI22_X1 U10762 ( .A1(n9529), .A2(n9642), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9612), .ZN(n9530) );
  OAI211_X1 U10763 ( .C1(n9612), .C2(n9532), .A(n9531), .B(n9530), .ZN(
        P1_U3266) );
  XOR2_X1 U10764 ( .A(n9534), .B(n9533), .Z(n9765) );
  AOI21_X1 U10765 ( .B1(n9535), .B2(n9534), .A(n4541), .ZN(n9536) );
  OAI222_X1 U10766 ( .A1(n9664), .A2(n9537), .B1(n9662), .B2(n9570), .C1(n9659), .C2(n9536), .ZN(n9761) );
  INV_X1 U10767 ( .A(n9555), .ZN(n9540) );
  INV_X1 U10768 ( .A(n9538), .ZN(n9539) );
  AOI211_X1 U10769 ( .C1(n9763), .C2(n9540), .A(n9969), .B(n9539), .ZN(n9762)
         );
  NAND2_X1 U10770 ( .A1(n9762), .A2(n9950), .ZN(n9543) );
  AOI22_X1 U10771 ( .A1(n9612), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9541), .B2(
        n9942), .ZN(n9542) );
  OAI211_X1 U10772 ( .C1(n9544), .C2(n9945), .A(n9543), .B(n9542), .ZN(n9545)
         );
  AOI21_X1 U10773 ( .B1(n9761), .B2(n9714), .A(n9545), .ZN(n9546) );
  OAI21_X1 U10774 ( .B1(n9765), .B2(n9741), .A(n9546), .ZN(P1_U3267) );
  XOR2_X1 U10775 ( .A(n9547), .B(n9548), .Z(n9768) );
  INV_X1 U10776 ( .A(n9768), .ZN(n9563) );
  INV_X1 U10777 ( .A(n9548), .ZN(n9549) );
  XNOR2_X1 U10778 ( .A(n9550), .B(n9549), .ZN(n9551) );
  NAND2_X1 U10779 ( .A1(n9551), .A2(n9724), .ZN(n9554) );
  INV_X1 U10780 ( .A(n9552), .ZN(n9553) );
  NAND2_X1 U10781 ( .A1(n9554), .A2(n9553), .ZN(n9766) );
  INV_X1 U10782 ( .A(n9571), .ZN(n9556) );
  AOI211_X1 U10783 ( .C1(n9557), .C2(n9556), .A(n9969), .B(n9555), .ZN(n9767)
         );
  NAND2_X1 U10784 ( .A1(n9767), .A2(n9950), .ZN(n9560) );
  AOI22_X1 U10785 ( .A1(n9558), .A2(n9942), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9612), .ZN(n9559) );
  OAI211_X1 U10786 ( .C1(n9838), .C2(n9945), .A(n9560), .B(n9559), .ZN(n9561)
         );
  AOI21_X1 U10787 ( .B1(n9714), .B2(n9766), .A(n9561), .ZN(n9562) );
  OAI21_X1 U10788 ( .B1(n9563), .B2(n9741), .A(n9562), .ZN(P1_U3268) );
  XNOR2_X1 U10789 ( .A(n9564), .B(n9566), .ZN(n9775) );
  NAND2_X1 U10790 ( .A1(n9580), .A2(n9565), .ZN(n9567) );
  XNOR2_X1 U10791 ( .A(n9567), .B(n9566), .ZN(n9568) );
  OAI222_X1 U10792 ( .A1(n9664), .A2(n9570), .B1(n9662), .B2(n9569), .C1(n9568), .C2(n9659), .ZN(n9771) );
  INV_X1 U10793 ( .A(n9589), .ZN(n9572) );
  AOI211_X1 U10794 ( .C1(n9773), .C2(n9572), .A(n9969), .B(n9571), .ZN(n9772)
         );
  NAND2_X1 U10795 ( .A1(n9772), .A2(n9950), .ZN(n9575) );
  AOI22_X1 U10796 ( .A1(n9573), .A2(n9942), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9612), .ZN(n9574) );
  OAI211_X1 U10797 ( .C1(n9576), .C2(n9945), .A(n9575), .B(n9574), .ZN(n9577)
         );
  AOI21_X1 U10798 ( .B1(n9771), .B2(n9714), .A(n9577), .ZN(n9578) );
  OAI21_X1 U10799 ( .B1(n9775), .B2(n9741), .A(n9578), .ZN(P1_U3269) );
  XNOR2_X1 U10800 ( .A(n9579), .B(n9582), .ZN(n9778) );
  INV_X1 U10801 ( .A(n9778), .ZN(n9597) );
  OAI21_X1 U10802 ( .B1(n9582), .B2(n9581), .A(n9580), .ZN(n9583) );
  NAND2_X1 U10803 ( .A1(n9583), .A2(n9724), .ZN(n9588) );
  OAI22_X1 U10804 ( .A1(n9585), .A2(n9664), .B1(n9584), .B2(n9662), .ZN(n9586)
         );
  INV_X1 U10805 ( .A(n9586), .ZN(n9587) );
  NAND2_X1 U10806 ( .A1(n9588), .A2(n9587), .ZN(n9776) );
  AOI211_X1 U10807 ( .C1(n9590), .C2(n9600), .A(n9969), .B(n9589), .ZN(n9777)
         );
  NAND2_X1 U10808 ( .A1(n9777), .A2(n9950), .ZN(n9594) );
  INV_X1 U10809 ( .A(n9591), .ZN(n9592) );
  AOI22_X1 U10810 ( .A1(n9592), .A2(n9942), .B1(n9612), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9593) );
  OAI211_X1 U10811 ( .C1(n9843), .C2(n9945), .A(n9594), .B(n9593), .ZN(n9595)
         );
  AOI21_X1 U10812 ( .B1(n9714), .B2(n9776), .A(n9595), .ZN(n9596) );
  OAI21_X1 U10813 ( .B1(n9597), .B2(n9741), .A(n9596), .ZN(P1_U3270) );
  XNOR2_X1 U10814 ( .A(n9598), .B(n9607), .ZN(n9785) );
  INV_X1 U10815 ( .A(n9600), .ZN(n9601) );
  AOI211_X1 U10816 ( .C1(n9782), .C2(n9625), .A(n9969), .B(n9601), .ZN(n9781)
         );
  INV_X1 U10817 ( .A(n9602), .ZN(n9603) );
  AOI22_X1 U10818 ( .A1(n9612), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9603), .B2(
        n9942), .ZN(n9604) );
  OAI21_X1 U10819 ( .B1(n9605), .B2(n9945), .A(n9604), .ZN(n9614) );
  OAI21_X1 U10820 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(n9611) );
  AOI222_X1 U10821 ( .A1(n9724), .A2(n9611), .B1(n9610), .B2(n9727), .C1(n9609), .C2(n9728), .ZN(n9784) );
  NOR2_X1 U10822 ( .A1(n9784), .A2(n9612), .ZN(n9613) );
  AOI211_X1 U10823 ( .C1(n9781), .C2(n9950), .A(n9614), .B(n9613), .ZN(n9615)
         );
  OAI21_X1 U10824 ( .B1(n9785), .B2(n9741), .A(n9615), .ZN(P1_U3271) );
  XOR2_X1 U10825 ( .A(n9622), .B(n9616), .Z(n9788) );
  INV_X1 U10826 ( .A(n9788), .ZN(n9633) );
  NAND2_X1 U10827 ( .A1(n9618), .A2(n9617), .ZN(n9621) );
  INV_X1 U10828 ( .A(n9619), .ZN(n9620) );
  AOI21_X1 U10829 ( .B1(n9622), .B2(n9621), .A(n9620), .ZN(n9624) );
  OAI21_X1 U10830 ( .B1(n9624), .B2(n9659), .A(n9623), .ZN(n9786) );
  AOI211_X1 U10831 ( .C1(n9626), .C2(n9640), .A(n9969), .B(n9599), .ZN(n9787)
         );
  NAND2_X1 U10832 ( .A1(n9787), .A2(n9950), .ZN(n9630) );
  INV_X1 U10833 ( .A(n9627), .ZN(n9628) );
  AOI22_X1 U10834 ( .A1(n9612), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9628), .B2(
        n9942), .ZN(n9629) );
  OAI211_X1 U10835 ( .C1(n9848), .C2(n9945), .A(n9630), .B(n9629), .ZN(n9631)
         );
  AOI21_X1 U10836 ( .B1(n9786), .B2(n9714), .A(n9631), .ZN(n9632) );
  OAI21_X1 U10837 ( .B1(n9633), .B2(n9741), .A(n9632), .ZN(P1_U3272) );
  XNOR2_X1 U10838 ( .A(n9634), .B(n9635), .ZN(n9793) );
  XNOR2_X1 U10839 ( .A(n9637), .B(n9636), .ZN(n9639) );
  AOI21_X1 U10840 ( .B1(n9639), .B2(n9724), .A(n9638), .ZN(n9792) );
  INV_X1 U10841 ( .A(n9792), .ZN(n9648) );
  OAI211_X1 U10842 ( .C1(n9852), .C2(n9651), .A(n9813), .B(n9640), .ZN(n9791)
         );
  AOI22_X1 U10843 ( .A1(n9612), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9641), .B2(
        n9942), .ZN(n9645) );
  NAND2_X1 U10844 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  OAI211_X1 U10845 ( .C1(n9791), .C2(n9646), .A(n9645), .B(n9644), .ZN(n9647)
         );
  AOI21_X1 U10846 ( .B1(n9648), .B2(n9714), .A(n9647), .ZN(n9649) );
  OAI21_X1 U10847 ( .B1(n9793), .B2(n9741), .A(n9649), .ZN(P1_U3273) );
  XOR2_X1 U10848 ( .A(n9650), .B(n9657), .Z(n9800) );
  AOI211_X1 U10849 ( .C1(n9798), .C2(n9669), .A(n9969), .B(n9651), .ZN(n9797)
         );
  NOR2_X1 U10850 ( .A1(n9652), .A2(n9945), .ZN(n9656) );
  OAI22_X1 U10851 ( .A1(n9714), .A2(n9654), .B1(n9653), .B2(n9711), .ZN(n9655)
         );
  AOI211_X1 U10852 ( .C1(n9797), .C2(n9950), .A(n9656), .B(n9655), .ZN(n9666)
         );
  XNOR2_X1 U10853 ( .A(n9658), .B(n9657), .ZN(n9660) );
  OAI222_X1 U10854 ( .A1(n9664), .A2(n9663), .B1(n9662), .B2(n9661), .C1(n9660), .C2(n9659), .ZN(n9796) );
  NAND2_X1 U10855 ( .A1(n9796), .A2(n9714), .ZN(n9665) );
  OAI211_X1 U10856 ( .C1(n9800), .C2(n9741), .A(n9666), .B(n9665), .ZN(
        P1_U3274) );
  INV_X1 U10857 ( .A(n9667), .ZN(n9668) );
  XNOR2_X1 U10858 ( .A(n9668), .B(n9676), .ZN(n9805) );
  INV_X1 U10859 ( .A(n9669), .ZN(n9670) );
  AOI211_X1 U10860 ( .C1(n4719), .C2(n4720), .A(n9969), .B(n9670), .ZN(n9801)
         );
  INV_X1 U10861 ( .A(n9671), .ZN(n9672) );
  AOI22_X1 U10862 ( .A1(n9612), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9672), .B2(
        n9942), .ZN(n9673) );
  OAI21_X1 U10863 ( .B1(n9674), .B2(n9945), .A(n9673), .ZN(n9680) );
  OAI21_X1 U10864 ( .B1(n9676), .B2(n4572), .A(n9675), .ZN(n9678) );
  AOI222_X1 U10865 ( .A1(n9724), .A2(n9678), .B1(n9677), .B2(n9728), .C1(n9702), .C2(n9727), .ZN(n9803) );
  NOR2_X1 U10866 ( .A1(n9803), .A2(n9612), .ZN(n9679) );
  AOI211_X1 U10867 ( .C1(n9801), .C2(n9950), .A(n9680), .B(n9679), .ZN(n9681)
         );
  OAI21_X1 U10868 ( .B1(n9805), .B2(n9741), .A(n9681), .ZN(P1_U3275) );
  NAND2_X1 U10869 ( .A1(n9683), .A2(n9682), .ZN(n9684) );
  NAND3_X1 U10870 ( .A1(n9685), .A2(n9724), .A3(n9684), .ZN(n9687) );
  NAND2_X1 U10871 ( .A1(n9687), .A2(n9686), .ZN(n9806) );
  INV_X1 U10872 ( .A(n9806), .ZN(n9697) );
  XNOR2_X1 U10873 ( .A(n9688), .B(n5566), .ZN(n9808) );
  NAND2_X1 U10874 ( .A1(n9808), .A2(n9707), .ZN(n9696) );
  AOI211_X1 U10875 ( .C1(n9690), .C2(n9708), .A(n9969), .B(n9689), .ZN(n9807)
         );
  NOR2_X1 U10876 ( .A1(n9858), .A2(n9945), .ZN(n9694) );
  OAI22_X1 U10877 ( .A1(n9714), .A2(n9692), .B1(n9691), .B2(n9711), .ZN(n9693)
         );
  AOI211_X1 U10878 ( .C1(n9807), .C2(n9950), .A(n9694), .B(n9693), .ZN(n9695)
         );
  OAI211_X1 U10879 ( .C1(n9612), .C2(n9697), .A(n9696), .B(n9695), .ZN(
        P1_U3276) );
  OAI21_X1 U10880 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9703) );
  AOI222_X1 U10881 ( .A1(n9724), .A2(n9703), .B1(n9702), .B2(n9728), .C1(n9701), .C2(n9727), .ZN(n9816) );
  OR2_X1 U10882 ( .A1(n9705), .A2(n9704), .ZN(n9811) );
  NAND3_X1 U10883 ( .A1(n9811), .A2(n9706), .A3(n9707), .ZN(n9719) );
  INV_X1 U10884 ( .A(n9708), .ZN(n9709) );
  AOI21_X1 U10885 ( .B1(n9812), .B2(n9731), .A(n9709), .ZN(n9814) );
  NOR2_X1 U10886 ( .A1(n9710), .A2(n9945), .ZN(n9716) );
  OAI22_X1 U10887 ( .A1(n9714), .A2(n9713), .B1(n9712), .B2(n9711), .ZN(n9715)
         );
  AOI211_X1 U10888 ( .C1(n9814), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9718)
         );
  OAI211_X1 U10889 ( .C1(n9612), .C2(n9816), .A(n9719), .B(n9718), .ZN(
        P1_U3277) );
  XNOR2_X1 U10890 ( .A(n9720), .B(n9723), .ZN(n9820) );
  INV_X1 U10891 ( .A(n9820), .ZN(n9742) );
  OAI21_X1 U10892 ( .B1(n9723), .B2(n9722), .A(n9721), .ZN(n9725) );
  NAND2_X1 U10893 ( .A1(n9725), .A2(n9724), .ZN(n9730) );
  AOI22_X1 U10894 ( .A1(n4793), .A2(n9728), .B1(n9727), .B2(n9726), .ZN(n9729)
         );
  NAND2_X1 U10895 ( .A1(n9730), .A2(n9729), .ZN(n9818) );
  INV_X1 U10896 ( .A(n9731), .ZN(n9732) );
  AOI211_X1 U10897 ( .C1(n9734), .C2(n9733), .A(n9969), .B(n9732), .ZN(n9819)
         );
  NAND2_X1 U10898 ( .A1(n9819), .A2(n9950), .ZN(n9738) );
  INV_X1 U10899 ( .A(n9735), .ZN(n9736) );
  AOI22_X1 U10900 ( .A1(n9612), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9736), .B2(
        n9942), .ZN(n9737) );
  OAI211_X1 U10901 ( .C1(n9865), .C2(n9945), .A(n9738), .B(n9737), .ZN(n9739)
         );
  AOI21_X1 U10902 ( .B1(n9714), .B2(n9818), .A(n9739), .ZN(n9740) );
  OAI21_X1 U10903 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(P1_U3278) );
  INV_X1 U10904 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9744) );
  AND2_X1 U10905 ( .A1(n9747), .A2(n9746), .ZN(n9826) );
  INV_X1 U10906 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9748) );
  MUX2_X1 U10907 ( .A(n9826), .B(n9748), .S(n9985), .Z(n9749) );
  OAI21_X1 U10908 ( .B1(n9828), .B2(n9823), .A(n9749), .ZN(P1_U3552) );
  NAND2_X1 U10909 ( .A1(n9750), .A2(n9979), .ZN(n9755) );
  AOI21_X1 U10910 ( .B1(n9956), .B2(n9752), .A(n9751), .ZN(n9753) );
  NAND3_X1 U10911 ( .A1(n9755), .A2(n9754), .A3(n9753), .ZN(n9829) );
  MUX2_X1 U10912 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9829), .S(n9988), .Z(
        P1_U3550) );
  AOI211_X1 U10913 ( .C1(n9758), .C2(n9979), .A(n9757), .B(n9756), .ZN(n9830)
         );
  MUX2_X1 U10914 ( .A(n9759), .B(n9830), .S(n9988), .Z(n9760) );
  OAI21_X1 U10915 ( .B1(n9833), .B2(n9823), .A(n9760), .ZN(P1_U3549) );
  AOI211_X1 U10916 ( .C1(n9956), .C2(n9763), .A(n9762), .B(n9761), .ZN(n9764)
         );
  OAI21_X1 U10917 ( .B1(n9765), .B2(n9804), .A(n9764), .ZN(n9834) );
  MUX2_X1 U10918 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9834), .S(n9988), .Z(
        P1_U3548) );
  INV_X1 U10919 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9769) );
  AOI211_X1 U10920 ( .C1(n9768), .C2(n9979), .A(n9767), .B(n9766), .ZN(n9835)
         );
  MUX2_X1 U10921 ( .A(n9769), .B(n9835), .S(n9988), .Z(n9770) );
  OAI21_X1 U10922 ( .B1(n9838), .B2(n9823), .A(n9770), .ZN(P1_U3547) );
  AOI211_X1 U10923 ( .C1(n9956), .C2(n9773), .A(n9772), .B(n9771), .ZN(n9774)
         );
  OAI21_X1 U10924 ( .B1(n9775), .B2(n9804), .A(n9774), .ZN(n9839) );
  MUX2_X1 U10925 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9839), .S(n9988), .Z(
        P1_U3546) );
  INV_X1 U10926 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9779) );
  AOI211_X1 U10927 ( .C1(n9778), .C2(n9979), .A(n9777), .B(n9776), .ZN(n9840)
         );
  MUX2_X1 U10928 ( .A(n9779), .B(n9840), .S(n9988), .Z(n9780) );
  OAI21_X1 U10929 ( .B1(n9843), .B2(n9823), .A(n9780), .ZN(P1_U3545) );
  AOI21_X1 U10930 ( .B1(n9956), .B2(n9782), .A(n9781), .ZN(n9783) );
  OAI211_X1 U10931 ( .C1(n9785), .C2(n9804), .A(n9784), .B(n9783), .ZN(n9844)
         );
  MUX2_X1 U10932 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9844), .S(n9988), .Z(
        P1_U3544) );
  INV_X1 U10933 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9789) );
  AOI211_X1 U10934 ( .C1(n9788), .C2(n9979), .A(n9787), .B(n9786), .ZN(n9845)
         );
  MUX2_X1 U10935 ( .A(n9789), .B(n9845), .S(n9988), .Z(n9790) );
  OAI21_X1 U10936 ( .B1(n9848), .B2(n9823), .A(n9790), .ZN(P1_U3543) );
  OAI211_X1 U10937 ( .C1(n9793), .C2(n9804), .A(n9792), .B(n9791), .ZN(n9849)
         );
  MUX2_X1 U10938 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9849), .S(n9988), .Z(n9794) );
  INV_X1 U10939 ( .A(n9794), .ZN(n9795) );
  OAI21_X1 U10940 ( .B1(n9852), .B2(n9823), .A(n9795), .ZN(P1_U3542) );
  AOI211_X1 U10941 ( .C1(n9956), .C2(n9798), .A(n9797), .B(n9796), .ZN(n9799)
         );
  OAI21_X1 U10942 ( .B1(n9800), .B2(n9804), .A(n9799), .ZN(n9853) );
  MUX2_X1 U10943 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9853), .S(n9988), .Z(
        P1_U3541) );
  AOI21_X1 U10944 ( .B1(n9956), .B2(n4719), .A(n9801), .ZN(n9802) );
  OAI211_X1 U10945 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9854)
         );
  MUX2_X1 U10946 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9854), .S(n9988), .Z(
        P1_U3540) );
  AOI211_X1 U10947 ( .C1(n9808), .C2(n9979), .A(n9807), .B(n9806), .ZN(n9855)
         );
  MUX2_X1 U10948 ( .A(n9809), .B(n9855), .S(n9988), .Z(n9810) );
  OAI21_X1 U10949 ( .B1(n9858), .B2(n9823), .A(n9810), .ZN(P1_U3539) );
  NAND3_X1 U10950 ( .A1(n9811), .A2(n9706), .A3(n9979), .ZN(n9817) );
  AOI22_X1 U10951 ( .A1(n9814), .A2(n9813), .B1(n9956), .B2(n9812), .ZN(n9815)
         );
  NAND3_X1 U10952 ( .A1(n9817), .A2(n9816), .A3(n9815), .ZN(n9859) );
  MUX2_X1 U10953 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9859), .S(n9988), .Z(
        P1_U3538) );
  INV_X1 U10954 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9821) );
  AOI211_X1 U10955 ( .C1(n9820), .C2(n9979), .A(n9819), .B(n9818), .ZN(n9861)
         );
  MUX2_X1 U10956 ( .A(n9821), .B(n9861), .S(n9988), .Z(n9822) );
  OAI21_X1 U10957 ( .B1(n9865), .B2(n9823), .A(n9822), .ZN(P1_U3537) );
  MUX2_X1 U10958 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9824), .S(n9988), .Z(
        P1_U3522) );
  MUX2_X1 U10959 ( .A(n9826), .B(n9825), .S(n6057), .Z(n9827) );
  OAI21_X1 U10960 ( .B1(n9828), .B2(n9864), .A(n9827), .ZN(P1_U3520) );
  MUX2_X1 U10961 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9829), .S(n9860), .Z(
        P1_U3518) );
  MUX2_X1 U10962 ( .A(n9831), .B(n9830), .S(n9860), .Z(n9832) );
  OAI21_X1 U10963 ( .B1(n9833), .B2(n9864), .A(n9832), .ZN(P1_U3517) );
  MUX2_X1 U10964 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9834), .S(n9860), .Z(
        P1_U3516) );
  MUX2_X1 U10965 ( .A(n9836), .B(n9835), .S(n9860), .Z(n9837) );
  OAI21_X1 U10966 ( .B1(n9838), .B2(n9864), .A(n9837), .ZN(P1_U3515) );
  MUX2_X1 U10967 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9839), .S(n9860), .Z(
        P1_U3514) );
  INV_X1 U10968 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9841) );
  MUX2_X1 U10969 ( .A(n9841), .B(n9840), .S(n9860), .Z(n9842) );
  OAI21_X1 U10970 ( .B1(n9843), .B2(n9864), .A(n9842), .ZN(P1_U3513) );
  MUX2_X1 U10971 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9844), .S(n9860), .Z(
        P1_U3512) );
  INV_X1 U10972 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9846) );
  MUX2_X1 U10973 ( .A(n9846), .B(n9845), .S(n9860), .Z(n9847) );
  OAI21_X1 U10974 ( .B1(n9848), .B2(n9864), .A(n9847), .ZN(P1_U3511) );
  MUX2_X1 U10975 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9849), .S(n9860), .Z(n9850) );
  INV_X1 U10976 ( .A(n9850), .ZN(n9851) );
  OAI21_X1 U10977 ( .B1(n9852), .B2(n9864), .A(n9851), .ZN(P1_U3510) );
  MUX2_X1 U10978 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9853), .S(n9860), .Z(
        P1_U3509) );
  MUX2_X1 U10979 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9854), .S(n9860), .Z(
        P1_U3507) );
  INV_X1 U10980 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9856) );
  MUX2_X1 U10981 ( .A(n9856), .B(n9855), .S(n9860), .Z(n9857) );
  OAI21_X1 U10982 ( .B1(n9858), .B2(n9864), .A(n9857), .ZN(P1_U3504) );
  MUX2_X1 U10983 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9859), .S(n9860), .Z(
        P1_U3501) );
  INV_X1 U10984 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9862) );
  MUX2_X1 U10985 ( .A(n9862), .B(n9861), .S(n9860), .Z(n9863) );
  OAI21_X1 U10986 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(P1_U3498) );
  MUX2_X1 U10987 ( .A(P1_D_REG_0__SCAN_IN), .B(n9867), .S(n9866), .Z(P1_U3439)
         );
  INV_X1 U10988 ( .A(n6066), .ZN(n9873) );
  INV_X1 U10989 ( .A(n9868), .ZN(n9869) );
  NOR4_X1 U10990 ( .A1(n9869), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n4641), .ZN(n9870) );
  AOI21_X1 U10991 ( .B1(n9871), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9870), .ZN(
        n9872) );
  OAI21_X1 U10992 ( .B1(n9873), .B2(n9884), .A(n9872), .ZN(P1_U3324) );
  OAI222_X1 U10993 ( .A1(n9874), .A2(P1_U3086), .B1(n9884), .B2(n9875), .C1(
        n10522), .C2(n9882), .ZN(P1_U3325) );
  OAI222_X1 U10994 ( .A1(P1_U3086), .A2(n9877), .B1(n9884), .B2(n9876), .C1(
        n10247), .C2(n9882), .ZN(P1_U3326) );
  OAI222_X1 U10995 ( .A1(P1_U3086), .A2(n5966), .B1(n9884), .B2(n9878), .C1(
        n10244), .C2(n9882), .ZN(P1_U3327) );
  OAI222_X1 U10996 ( .A1(P1_U3086), .A2(n9927), .B1(n9884), .B2(n9879), .C1(
        n10265), .C2(n9882), .ZN(P1_U3328) );
  OAI222_X1 U10997 ( .A1(n9881), .A2(P1_U3086), .B1(n9884), .B2(n9880), .C1(
        n10246), .C2(n9882), .ZN(P1_U3329) );
  OAI222_X1 U10998 ( .A1(n9885), .A2(P1_U3086), .B1(n9884), .B2(n9883), .C1(
        n10221), .C2(n9882), .ZN(P1_U3330) );
  MUX2_X1 U10999 ( .A(n9886), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11000 ( .A(n9887), .ZN(n9892) );
  OAI22_X1 U11001 ( .A1(n9890), .A2(n9889), .B1(n9903), .B2(n9888), .ZN(n9891)
         );
  AOI21_X1 U11002 ( .B1(n9892), .B2(n9906), .A(n9891), .ZN(n9893) );
  OAI21_X1 U11003 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(P1_U3232) );
  OAI21_X1 U11004 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(n9907) );
  AOI21_X1 U11005 ( .B1(n9901), .B2(n9900), .A(n9899), .ZN(n9902) );
  OAI21_X1 U11006 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(n9905) );
  AOI21_X1 U11007 ( .B1(n9907), .B2(n9906), .A(n9905), .ZN(n9908) );
  OAI21_X1 U11008 ( .B1(n9909), .B2(n9923), .A(n9908), .ZN(P1_U3217) );
  XNOR2_X1 U11009 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11010 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11011 ( .B1(n9912), .B2(n9911), .A(n9910), .ZN(n9919) );
  AOI21_X1 U11012 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9917) );
  NOR2_X1 U11013 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  AOI211_X1 U11014 ( .C1(n9921), .C2(n9920), .A(n9919), .B(n9918), .ZN(n9922)
         );
  OAI21_X1 U11015 ( .B1(n9924), .B2(n9923), .A(n9922), .ZN(P1_U3221) );
  INV_X1 U11016 ( .A(n9925), .ZN(n9932) );
  NAND2_X1 U11017 ( .A1(n9927), .A2(n9926), .ZN(n9930) );
  NAND2_X1 U11018 ( .A1(n9928), .A2(n9930), .ZN(n9929) );
  MUX2_X1 U11019 ( .A(n9930), .B(n9929), .S(P1_IR_REG_0__SCAN_IN), .Z(n9931)
         );
  NAND2_X1 U11020 ( .A1(n9932), .A2(n9931), .ZN(n9935) );
  AOI22_X1 U11021 ( .A1(n9933), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9934) );
  OAI21_X1 U11022 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(P1_U3243) );
  INV_X1 U11023 ( .A(n9937), .ZN(n9938) );
  AOI21_X1 U11024 ( .B1(n9940), .B2(n9939), .A(n9938), .ZN(n9953) );
  INV_X1 U11025 ( .A(n9941), .ZN(n9951) );
  AOI22_X1 U11026 ( .A1(n9612), .A2(P1_REG2_REG_1__SCAN_IN), .B1(n9942), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n9943) );
  OAI21_X1 U11027 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(n9949) );
  NOR3_X1 U11028 ( .A1(n9947), .A2(n9612), .A3(n9946), .ZN(n9948) );
  AOI211_X1 U11029 ( .C1(n9951), .C2(n9950), .A(n9949), .B(n9948), .ZN(n9952)
         );
  OAI21_X1 U11030 ( .B1(n9612), .B2(n9953), .A(n9952), .ZN(P1_U3292) );
  AND2_X1 U11031 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9954), .ZN(P1_U3294) );
  AND2_X1 U11032 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9954), .ZN(P1_U3295) );
  AND2_X1 U11033 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9954), .ZN(P1_U3296) );
  AND2_X1 U11034 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9954), .ZN(P1_U3297) );
  AND2_X1 U11035 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9954), .ZN(P1_U3298) );
  AND2_X1 U11036 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9954), .ZN(P1_U3299) );
  AND2_X1 U11037 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9954), .ZN(P1_U3300) );
  AND2_X1 U11038 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9954), .ZN(P1_U3301) );
  AND2_X1 U11039 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9954), .ZN(P1_U3302) );
  AND2_X1 U11040 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9954), .ZN(P1_U3303) );
  AND2_X1 U11041 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9954), .ZN(P1_U3304) );
  AND2_X1 U11042 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9954), .ZN(P1_U3305) );
  AND2_X1 U11043 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9954), .ZN(P1_U3306) );
  AND2_X1 U11044 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9954), .ZN(P1_U3307) );
  AND2_X1 U11045 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9954), .ZN(P1_U3308) );
  AND2_X1 U11046 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9954), .ZN(P1_U3309) );
  AND2_X1 U11047 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9954), .ZN(P1_U3310) );
  AND2_X1 U11048 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9954), .ZN(P1_U3311) );
  AND2_X1 U11049 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9954), .ZN(P1_U3312) );
  AND2_X1 U11050 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9954), .ZN(P1_U3313) );
  AND2_X1 U11051 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9954), .ZN(P1_U3314) );
  AND2_X1 U11052 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9954), .ZN(P1_U3315) );
  AND2_X1 U11053 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9954), .ZN(P1_U3316) );
  AND2_X1 U11054 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9954), .ZN(P1_U3317) );
  AND2_X1 U11055 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9954), .ZN(P1_U3318) );
  AND2_X1 U11056 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9954), .ZN(P1_U3319) );
  NOR2_X1 U11057 ( .A1(n9955), .A2(n10498), .ZN(P1_U3320) );
  NOR2_X1 U11058 ( .A1(n9955), .A2(n10211), .ZN(P1_U3321) );
  NOR2_X1 U11059 ( .A1(n9955), .A2(n10368), .ZN(P1_U3322) );
  NOR2_X1 U11060 ( .A1(n9955), .A2(n10524), .ZN(P1_U3323) );
  OAI22_X1 U11061 ( .A1(n9958), .A2(n9969), .B1(n9957), .B2(n6011), .ZN(n9960)
         );
  AOI211_X1 U11062 ( .C1(n9979), .C2(n9961), .A(n9960), .B(n9959), .ZN(n9982)
         );
  INV_X1 U11063 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U11064 ( .A1(n9860), .A2(n9982), .B1(n9962), .B2(n6057), .ZN(
        P1_U3465) );
  OAI211_X1 U11065 ( .C1(n9965), .C2(n6011), .A(n9964), .B(n9963), .ZN(n9966)
         );
  AOI21_X1 U11066 ( .B1(n9979), .B2(n9967), .A(n9966), .ZN(n9983) );
  INV_X1 U11067 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9968) );
  AOI22_X1 U11068 ( .A1(n9860), .A2(n9983), .B1(n9968), .B2(n6057), .ZN(
        P1_U3480) );
  OAI22_X1 U11069 ( .A1(n9970), .A2(n9969), .B1(n6024), .B2(n6011), .ZN(n9971)
         );
  AOI211_X1 U11070 ( .C1(n9973), .C2(n9979), .A(n9972), .B(n9971), .ZN(n9984)
         );
  INV_X1 U11071 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11072 ( .A1(n9860), .A2(n9984), .B1(n9974), .B2(n6057), .ZN(
        P1_U3489) );
  OAI21_X1 U11073 ( .B1(n9976), .B2(n6011), .A(n9975), .ZN(n9977) );
  AOI211_X1 U11074 ( .C1(n9980), .C2(n9979), .A(n9978), .B(n9977), .ZN(n9987)
         );
  INV_X1 U11075 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U11076 ( .A1(n9860), .A2(n9987), .B1(n9981), .B2(n6057), .ZN(
        P1_U3495) );
  AOI22_X1 U11077 ( .A1(n9988), .A2(n9982), .B1(n6894), .B2(n9985), .ZN(
        P1_U3526) );
  AOI22_X1 U11078 ( .A1(n9988), .A2(n9983), .B1(n6904), .B2(n9985), .ZN(
        P1_U3531) );
  AOI22_X1 U11079 ( .A1(n9988), .A2(n9984), .B1(n6954), .B2(n9985), .ZN(
        P1_U3534) );
  AOI22_X1 U11080 ( .A1(n9988), .A2(n9987), .B1(n9986), .B2(n9985), .ZN(
        P1_U3536) );
  INV_X1 U11081 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10102) );
  OAI21_X1 U11082 ( .B1(n9990), .B2(n9989), .A(n10020), .ZN(n10003) );
  NAND2_X1 U11083 ( .A1(n9991), .A2(n6799), .ZN(n9992) );
  NAND2_X1 U11084 ( .A1(n9993), .A2(n9992), .ZN(n9996) );
  NOR2_X1 U11085 ( .A1(n9994), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9995) );
  AOI21_X1 U11086 ( .B1(n9997), .B2(n9996), .A(n9995), .ZN(n10001) );
  INV_X1 U11087 ( .A(n9998), .ZN(n9999) );
  NAND2_X1 U11088 ( .A1(n10014), .A2(n9999), .ZN(n10000) );
  OAI211_X1 U11089 ( .C1(n10003), .C2(n10002), .A(n10001), .B(n10000), .ZN(
        n10004) );
  INV_X1 U11090 ( .A(n10004), .ZN(n10010) );
  INV_X1 U11091 ( .A(n10005), .ZN(n10006) );
  AOI21_X1 U11092 ( .B1(n7305), .B2(n10007), .A(n10006), .ZN(n10008) );
  OR2_X1 U11093 ( .A1(n10026), .A2(n10008), .ZN(n10009) );
  OAI211_X1 U11094 ( .C1(n10102), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        P2_U3183) );
  AOI21_X1 U11095 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(n10031) );
  OAI21_X1 U11096 ( .B1(n10017), .B2(n10016), .A(n10015), .ZN(n10019) );
  AOI22_X1 U11097 ( .A1(n10020), .A2(n10019), .B1(n10018), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n10030) );
  AOI21_X1 U11098 ( .B1(n10021), .B2(n6360), .A(n4594), .ZN(n10023) );
  OR2_X1 U11099 ( .A1(n10023), .A2(n10022), .ZN(n10029) );
  AOI21_X1 U11100 ( .B1(n10025), .B2(n7796), .A(n10024), .ZN(n10027) );
  OR2_X1 U11101 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  NAND4_X1 U11102 ( .A1(n10031), .A2(n10030), .A3(n10029), .A4(n10028), .ZN(
        P2_U3189) );
  AOI22_X1 U11103 ( .A1(n10034), .A2(n10033), .B1(n10085), .B2(n10032), .ZN(
        n10035) );
  AND2_X1 U11104 ( .A1(n10036), .A2(n10035), .ZN(n10088) );
  AOI22_X1 U11105 ( .A1(n10087), .A2(n6303), .B1(n10088), .B2(n10086), .ZN(
        P2_U3396) );
  INV_X1 U11106 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10042) );
  INV_X1 U11107 ( .A(n10037), .ZN(n10041) );
  OAI22_X1 U11108 ( .A1(n10039), .A2(n10080), .B1(n10038), .B2(n10073), .ZN(
        n10040) );
  NOR2_X1 U11109 ( .A1(n10041), .A2(n10040), .ZN(n10089) );
  AOI22_X1 U11110 ( .A1(n10087), .A2(n10042), .B1(n10089), .B2(n10086), .ZN(
        P2_U3399) );
  INV_X1 U11111 ( .A(n10043), .ZN(n10047) );
  OAI22_X1 U11112 ( .A1(n10045), .A2(n10080), .B1(n10044), .B2(n10073), .ZN(
        n10046) );
  NOR2_X1 U11113 ( .A1(n10047), .A2(n10046), .ZN(n10090) );
  AOI22_X1 U11114 ( .A1(n10087), .A2(n6325), .B1(n10090), .B2(n10086), .ZN(
        P2_U3402) );
  INV_X1 U11115 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10052) );
  OAI22_X1 U11116 ( .A1(n10049), .A2(n6746), .B1(n10048), .B2(n10073), .ZN(
        n10050) );
  NOR2_X1 U11117 ( .A1(n10051), .A2(n10050), .ZN(n10091) );
  AOI22_X1 U11118 ( .A1(n10087), .A2(n10052), .B1(n10091), .B2(n10086), .ZN(
        P2_U3405) );
  INV_X1 U11119 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10057) );
  OAI22_X1 U11120 ( .A1(n10054), .A2(n6746), .B1(n10053), .B2(n10073), .ZN(
        n10055) );
  NOR2_X1 U11121 ( .A1(n10056), .A2(n10055), .ZN(n10092) );
  AOI22_X1 U11122 ( .A1(n10087), .A2(n10057), .B1(n10092), .B2(n10086), .ZN(
        P2_U3411) );
  INV_X1 U11123 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10063) );
  INV_X1 U11124 ( .A(n10058), .ZN(n10062) );
  OAI22_X1 U11125 ( .A1(n10060), .A2(n10080), .B1(n10059), .B2(n10073), .ZN(
        n10061) );
  NOR2_X1 U11126 ( .A1(n10062), .A2(n10061), .ZN(n10093) );
  AOI22_X1 U11127 ( .A1(n10087), .A2(n10063), .B1(n10093), .B2(n10086), .ZN(
        P2_U3414) );
  NOR2_X1 U11128 ( .A1(n10064), .A2(n6746), .ZN(n10066) );
  AOI211_X1 U11129 ( .C1(n10085), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        n10094) );
  AOI22_X1 U11130 ( .A1(n10087), .A2(n6410), .B1(n10094), .B2(n10086), .ZN(
        P2_U3417) );
  INV_X1 U11131 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10072) );
  NOR2_X1 U11132 ( .A1(n10068), .A2(n6746), .ZN(n10070) );
  AOI211_X1 U11133 ( .C1(n10085), .C2(n10071), .A(n10070), .B(n10069), .ZN(
        n10095) );
  AOI22_X1 U11134 ( .A1(n10087), .A2(n10072), .B1(n10095), .B2(n10086), .ZN(
        P2_U3420) );
  INV_X1 U11135 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10079) );
  NOR2_X1 U11136 ( .A1(n10074), .A2(n10073), .ZN(n10076) );
  AOI211_X1 U11137 ( .C1(n10078), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        n10096) );
  AOI22_X1 U11138 ( .A1(n10087), .A2(n10079), .B1(n10096), .B2(n10086), .ZN(
        P2_U3423) );
  NOR2_X1 U11139 ( .A1(n10081), .A2(n10080), .ZN(n10083) );
  AOI211_X1 U11140 ( .C1(n10085), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10098) );
  AOI22_X1 U11141 ( .A1(n10087), .A2(n6439), .B1(n10098), .B2(n10086), .ZN(
        P2_U3426) );
  AOI22_X1 U11142 ( .A1(n10099), .A2(n10088), .B1(n6301), .B2(n10097), .ZN(
        P2_U3461) );
  AOI22_X1 U11143 ( .A1(n10099), .A2(n10089), .B1(n6798), .B2(n10097), .ZN(
        P2_U3462) );
  AOI22_X1 U11144 ( .A1(n10099), .A2(n10090), .B1(n6326), .B2(n10097), .ZN(
        P2_U3463) );
  AOI22_X1 U11145 ( .A1(n10099), .A2(n10091), .B1(n6280), .B2(n10097), .ZN(
        P2_U3464) );
  AOI22_X1 U11146 ( .A1(n10099), .A2(n10092), .B1(n6360), .B2(n10097), .ZN(
        P2_U3466) );
  AOI22_X1 U11147 ( .A1(n10099), .A2(n10093), .B1(n6348), .B2(n10097), .ZN(
        P2_U3467) );
  AOI22_X1 U11148 ( .A1(n10099), .A2(n10094), .B1(n6407), .B2(n10097), .ZN(
        P2_U3468) );
  AOI22_X1 U11149 ( .A1(n10099), .A2(n10095), .B1(n6420), .B2(n10097), .ZN(
        P2_U3469) );
  AOI22_X1 U11150 ( .A1(n10099), .A2(n10096), .B1(n8057), .B2(n10097), .ZN(
        P2_U3470) );
  AOI22_X1 U11151 ( .A1(n10099), .A2(n10098), .B1(n8067), .B2(n10097), .ZN(
        P2_U3471) );
  NAND2_X1 U11152 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10100) );
  NOR2_X1 U11153 ( .A1(n10101), .A2(n10100), .ZN(n10104) );
  AOI21_X1 U11154 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10106) );
  NOR2_X1 U11155 ( .A1(n10104), .A2(n10106), .ZN(n10103) );
  XNOR2_X1 U11156 ( .A(n10103), .B(n10102), .ZN(ADD_1068_U5) );
  XOR2_X1 U11157 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11158 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10153) );
  NOR2_X1 U11159 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10151) );
  NOR2_X1 U11160 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10147) );
  NOR2_X1 U11161 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10143) );
  NOR2_X1 U11162 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10141) );
  NOR2_X1 U11163 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10137) );
  NOR2_X1 U11164 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10133) );
  NOR2_X1 U11165 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10129) );
  NOR2_X1 U11166 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10125) );
  NOR2_X1 U11167 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10121) );
  NOR2_X1 U11168 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10118) );
  NOR2_X1 U11169 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10116) );
  NOR2_X1 U11170 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10114) );
  NOR2_X1 U11171 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10112) );
  NAND2_X1 U11172 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10110) );
  XOR2_X1 U11173 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10569) );
  NAND2_X1 U11174 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10108) );
  NOR2_X1 U11175 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10104), .ZN(n10105) );
  NOR2_X1 U11176 ( .A1(n10106), .A2(n10105), .ZN(n10559) );
  XOR2_X1 U11177 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10558) );
  NAND2_X1 U11178 ( .A1(n10559), .A2(n10558), .ZN(n10107) );
  NAND2_X1 U11179 ( .A1(n10108), .A2(n10107), .ZN(n10568) );
  NAND2_X1 U11180 ( .A1(n10569), .A2(n10568), .ZN(n10109) );
  NAND2_X1 U11181 ( .A1(n10110), .A2(n10109), .ZN(n10571) );
  XNOR2_X1 U11182 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10570) );
  NOR2_X1 U11183 ( .A1(n10571), .A2(n10570), .ZN(n10111) );
  NOR2_X1 U11184 ( .A1(n10112), .A2(n10111), .ZN(n10561) );
  XNOR2_X1 U11185 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10560) );
  NOR2_X1 U11186 ( .A1(n10561), .A2(n10560), .ZN(n10113) );
  NOR2_X1 U11187 ( .A1(n10114), .A2(n10113), .ZN(n10567) );
  XNOR2_X1 U11188 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10566) );
  NOR2_X1 U11189 ( .A1(n10567), .A2(n10566), .ZN(n10115) );
  NOR2_X1 U11190 ( .A1(n10116), .A2(n10115), .ZN(n10563) );
  XNOR2_X1 U11191 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10562) );
  NOR2_X1 U11192 ( .A1(n10563), .A2(n10562), .ZN(n10117) );
  NOR2_X1 U11193 ( .A1(n10118), .A2(n10117), .ZN(n10565) );
  INV_X1 U11194 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10119) );
  AOI22_X1 U11195 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n6934), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10119), .ZN(n10564) );
  NOR2_X1 U11196 ( .A1(n10565), .A2(n10564), .ZN(n10120) );
  NOR2_X1 U11197 ( .A1(n10121), .A2(n10120), .ZN(n10557) );
  INV_X1 U11198 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10123) );
  AOI22_X1 U11199 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10123), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10122), .ZN(n10556) );
  NOR2_X1 U11200 ( .A1(n10557), .A2(n10556), .ZN(n10124) );
  NOR2_X1 U11201 ( .A1(n10125), .A2(n10124), .ZN(n10171) );
  INV_X1 U11202 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U11203 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10127), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10126), .ZN(n10170) );
  NOR2_X1 U11204 ( .A1(n10171), .A2(n10170), .ZN(n10128) );
  NOR2_X1 U11205 ( .A1(n10129), .A2(n10128), .ZN(n10169) );
  INV_X1 U11206 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U11207 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10131), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10130), .ZN(n10168) );
  NOR2_X1 U11208 ( .A1(n10169), .A2(n10168), .ZN(n10132) );
  NOR2_X1 U11209 ( .A1(n10133), .A2(n10132), .ZN(n10167) );
  INV_X1 U11210 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U11211 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10135), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10134), .ZN(n10166) );
  NOR2_X1 U11212 ( .A1(n10167), .A2(n10166), .ZN(n10136) );
  NOR2_X1 U11213 ( .A1(n10137), .A2(n10136), .ZN(n10165) );
  INV_X1 U11214 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10139) );
  AOI22_X1 U11215 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10139), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10138), .ZN(n10164) );
  NOR2_X1 U11216 ( .A1(n10165), .A2(n10164), .ZN(n10140) );
  NOR2_X1 U11217 ( .A1(n10141), .A2(n10140), .ZN(n10163) );
  XNOR2_X1 U11218 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10162) );
  NOR2_X1 U11219 ( .A1(n10163), .A2(n10162), .ZN(n10142) );
  NOR2_X1 U11220 ( .A1(n10143), .A2(n10142), .ZN(n10161) );
  INV_X1 U11221 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U11222 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n10145), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10144), .ZN(n10160) );
  NOR2_X1 U11223 ( .A1(n10161), .A2(n10160), .ZN(n10146) );
  NOR2_X1 U11224 ( .A1(n10147), .A2(n10146), .ZN(n10159) );
  INV_X1 U11225 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U11226 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n10149), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n10148), .ZN(n10158) );
  NOR2_X1 U11227 ( .A1(n10159), .A2(n10158), .ZN(n10150) );
  NOR2_X1 U11228 ( .A1(n10151), .A2(n10150), .ZN(n10157) );
  XNOR2_X1 U11229 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10156) );
  NOR2_X1 U11230 ( .A1(n10157), .A2(n10156), .ZN(n10152) );
  NOR2_X1 U11231 ( .A1(n10153), .A2(n10152), .ZN(n10154) );
  NOR2_X1 U11232 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10154), .ZN(n10174) );
  AND2_X1 U11233 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10154), .ZN(n10172) );
  NOR2_X1 U11234 ( .A1(n10174), .A2(n10172), .ZN(n10155) );
  XOR2_X1 U11235 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10155), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11236 ( .A(n10157), .B(n10156), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11237 ( .A(n10159), .B(n10158), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11238 ( .A(n10161), .B(n10160), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11239 ( .A(n10163), .B(n10162), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11240 ( .A(n10165), .B(n10164), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11241 ( .A(n10167), .B(n10166), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11242 ( .A(n10169), .B(n10168), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11243 ( .A(n10171), .B(n10170), .ZN(ADD_1068_U63) );
  NOR2_X1 U11244 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10172), .ZN(n10173) );
  NOR2_X1 U11245 ( .A1(n10174), .A2(n10173), .ZN(n10555) );
  OAI22_X1 U11246 ( .A1(SI_18_), .A2(keyinput_g14), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n10175) );
  AOI221_X1 U11247 ( .B1(SI_18_), .B2(keyinput_g14), .C1(keyinput_g17), .C2(
        SI_15_), .A(n10175), .ZN(n10182) );
  OAI22_X1 U11248 ( .A1(SI_6_), .A2(keyinput_g26), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_g66), .ZN(n10176) );
  AOI221_X1 U11249 ( .B1(SI_6_), .B2(keyinput_g26), .C1(keyinput_g66), .C2(
        P2_DATAO_REG_30__SCAN_IN), .A(n10176), .ZN(n10181) );
  OAI22_X1 U11250 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput_g85), .B1(
        keyinput_g114), .B2(P1_IR_REG_24__SCAN_IN), .ZN(n10177) );
  AOI221_X1 U11251 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput_g114), .A(n10177), .ZN(n10180) );
  OAI22_X1 U11252 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        keyinput_g52), .B2(P2_REG3_REG_4__SCAN_IN), .ZN(n10178) );
  AOI221_X1 U11253 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_g52), .A(n10178), .ZN(n10179) );
  NAND4_X1 U11254 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10316) );
  OAI22_X1 U11255 ( .A1(SI_25_), .A2(keyinput_g7), .B1(keyinput_g105), .B2(
        P1_IR_REG_15__SCAN_IN), .ZN(n10183) );
  AOI221_X1 U11256 ( .B1(SI_25_), .B2(keyinput_g7), .C1(P1_IR_REG_15__SCAN_IN), 
        .C2(keyinput_g105), .A(n10183), .ZN(n10209) );
  INV_X1 U11257 ( .A(SI_16_), .ZN(n10189) );
  OAI22_X1 U11258 ( .A1(SI_2_), .A2(keyinput_g30), .B1(P1_IR_REG_9__SCAN_IN), 
        .B2(keyinput_g99), .ZN(n10184) );
  AOI221_X1 U11259 ( .B1(SI_2_), .B2(keyinput_g30), .C1(keyinput_g99), .C2(
        P1_IR_REG_9__SCAN_IN), .A(n10184), .ZN(n10187) );
  OAI22_X1 U11260 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_g82), .B1(
        keyinput_g107), .B2(P1_IR_REG_17__SCAN_IN), .ZN(n10185) );
  AOI221_X1 U11261 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_g107), .A(n10185), .ZN(n10186) );
  OAI211_X1 U11262 ( .C1(n10189), .C2(keyinput_g16), .A(n10187), .B(n10186), 
        .ZN(n10188) );
  AOI21_X1 U11263 ( .B1(n10189), .B2(keyinput_g16), .A(n10188), .ZN(n10208) );
  AOI22_X1 U11264 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_g90), .B1(SI_11_), 
        .B2(keyinput_g21), .ZN(n10190) );
  OAI221_X1 U11265 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_g90), .C1(SI_11_), 
        .C2(keyinput_g21), .A(n10190), .ZN(n10197) );
  AOI22_X1 U11266 ( .A1(SI_29_), .A2(keyinput_g3), .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n10191) );
  OAI221_X1 U11267 ( .B1(SI_29_), .B2(keyinput_g3), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n10191), .ZN(n10196)
         );
  AOI22_X1 U11268 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .ZN(n10192) );
  OAI221_X1 U11269 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_g51), .A(n10192), .ZN(n10195)
         );
  AOI22_X1 U11270 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_g112), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n10193) );
  OAI221_X1 U11271 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_g112), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n10193), .ZN(n10194)
         );
  NOR4_X1 U11272 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10207) );
  AOI22_X1 U11273 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(keyinput_g35), .ZN(n10198) );
  OAI221_X1 U11274 ( .B1(SI_4_), .B2(keyinput_g28), .C1(P2_REG3_REG_7__SCAN_IN), .C2(keyinput_g35), .A(n10198), .ZN(n10205) );
  AOI22_X1 U11275 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_g106), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .ZN(n10199) );
  OAI221_X1 U11276 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_g106), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_g76), .A(n10199), .ZN(n10204)
         );
  AOI22_X1 U11277 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n10200) );
  OAI221_X1 U11278 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n10200), .ZN(n10203) );
  AOI22_X1 U11279 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_g110), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .ZN(n10201) );
  OAI221_X1 U11280 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_g110), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_g75), .A(n10201), .ZN(n10202)
         );
  NOR4_X1 U11281 ( .A1(n10205), .A2(n10204), .A3(n10203), .A4(n10202), .ZN(
        n10206) );
  NAND4_X1 U11282 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10315) );
  AOI22_X1 U11283 ( .A1(n5410), .A2(keyinput_g98), .B1(keyinput_g126), .B2(
        n10211), .ZN(n10210) );
  OAI221_X1 U11284 ( .B1(n5410), .B2(keyinput_g98), .C1(n10211), .C2(
        keyinput_g126), .A(n10210), .ZN(n10219) );
  AOI22_X1 U11285 ( .A1(P2_U3151), .A2(keyinput_g34), .B1(keyinput_g81), .B2(
        n10403), .ZN(n10212) );
  OAI221_X1 U11286 ( .B1(P2_U3151), .B2(keyinput_g34), .C1(n10403), .C2(
        keyinput_g81), .A(n10212), .ZN(n10218) );
  INV_X1 U11287 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10364) );
  XOR2_X1 U11288 ( .A(n10364), .B(keyinput_g38), .Z(n10216) );
  XNOR2_X1 U11289 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_g72), .ZN(n10215) );
  XNOR2_X1 U11290 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g91), .ZN(n10214) );
  XNOR2_X1 U11291 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_g115), .ZN(n10213)
         );
  NAND4_X1 U11292 ( .A1(n10216), .A2(n10215), .A3(n10214), .A4(n10213), .ZN(
        n10217) );
  NOR3_X1 U11293 ( .A1(n10219), .A2(n10218), .A3(n10217), .ZN(n10258) );
  AOI22_X1 U11294 ( .A1(n10221), .A2(keyinput_g71), .B1(keyinput_g122), .B2(
        n10387), .ZN(n10220) );
  OAI221_X1 U11295 ( .B1(n10221), .B2(keyinput_g71), .C1(n10387), .C2(
        keyinput_g122), .A(n10220), .ZN(n10225) );
  XNOR2_X1 U11296 ( .A(n10368), .B(keyinput_g125), .ZN(n10224) );
  XNOR2_X1 U11297 ( .A(n10222), .B(keyinput_g31), .ZN(n10223) );
  OR3_X1 U11298 ( .A1(n10225), .A2(n10224), .A3(n10223), .ZN(n10233) );
  AOI22_X1 U11299 ( .A1(n10227), .A2(keyinput_g9), .B1(n6087), .B2(
        keyinput_g49), .ZN(n10226) );
  OAI221_X1 U11300 ( .B1(n10227), .B2(keyinput_g9), .C1(n6087), .C2(
        keyinput_g49), .A(n10226), .ZN(n10232) );
  INV_X1 U11301 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10230) );
  AOI22_X1 U11302 ( .A1(n10230), .A2(keyinput_g37), .B1(keyinput_g15), .B2(
        n10229), .ZN(n10228) );
  OAI221_X1 U11303 ( .B1(n10230), .B2(keyinput_g37), .C1(n10229), .C2(
        keyinput_g15), .A(n10228), .ZN(n10231) );
  NOR3_X1 U11304 ( .A1(n10233), .A2(n10232), .A3(n10231), .ZN(n10257) );
  AOI22_X1 U11305 ( .A1(n10512), .A2(keyinput_g123), .B1(n8412), .B2(
        keyinput_g41), .ZN(n10234) );
  OAI221_X1 U11306 ( .B1(n10512), .B2(keyinput_g123), .C1(n8412), .C2(
        keyinput_g41), .A(n10234), .ZN(n10242) );
  INV_X1 U11307 ( .A(SI_30_), .ZN(n10370) );
  AOI22_X1 U11308 ( .A1(n10370), .A2(keyinput_g2), .B1(n10481), .B2(
        keyinput_g19), .ZN(n10235) );
  OAI221_X1 U11309 ( .B1(n10370), .B2(keyinput_g2), .C1(n10481), .C2(
        keyinput_g19), .A(n10235), .ZN(n10241) );
  XNOR2_X1 U11310 ( .A(SI_3_), .B(keyinput_g29), .ZN(n10239) );
  XNOR2_X1 U11311 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_g80), .ZN(n10238) );
  XNOR2_X1 U11312 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g92), .ZN(n10237) );
  XNOR2_X1 U11313 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_g55), .ZN(n10236)
         );
  NAND4_X1 U11314 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10240) );
  NOR3_X1 U11315 ( .A1(n10242), .A2(n10241), .A3(n10240), .ZN(n10256) );
  AOI22_X1 U11316 ( .A1(n10494), .A2(keyinput_g39), .B1(keyinput_g68), .B2(
        n10244), .ZN(n10243) );
  OAI221_X1 U11317 ( .B1(n10494), .B2(keyinput_g39), .C1(n10244), .C2(
        keyinput_g68), .A(n10243), .ZN(n10254) );
  AOI22_X1 U11318 ( .A1(n10247), .A2(keyinput_g67), .B1(keyinput_g70), .B2(
        n10246), .ZN(n10245) );
  OAI221_X1 U11319 ( .B1(n10247), .B2(keyinput_g67), .C1(n10246), .C2(
        keyinput_g70), .A(n10245), .ZN(n10253) );
  XOR2_X1 U11320 ( .A(n5172), .B(keyinput_g116), .Z(n10251) );
  XOR2_X1 U11321 ( .A(n6091), .B(keyinput_g42), .Z(n10250) );
  XNOR2_X1 U11322 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g101), .ZN(n10249)
         );
  XNOR2_X1 U11323 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g97), .ZN(n10248) );
  NAND4_X1 U11324 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10252) );
  NOR3_X1 U11325 ( .A1(n10254), .A2(n10253), .A3(n10252), .ZN(n10255) );
  NAND4_X1 U11326 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10314) );
  INV_X1 U11327 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U11328 ( .A1(n10260), .A2(keyinput_g36), .B1(keyinput_g4), .B2(
        n10520), .ZN(n10259) );
  OAI221_X1 U11329 ( .B1(n10260), .B2(keyinput_g36), .C1(n10520), .C2(
        keyinput_g4), .A(n10259), .ZN(n10263) );
  INV_X1 U11330 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10261) );
  XNOR2_X1 U11331 ( .A(n10261), .B(keyinput_g0), .ZN(n10262) );
  NOR2_X1 U11332 ( .A1(n10263), .A2(n10262), .ZN(n10272) );
  AOI22_X1 U11333 ( .A1(n10483), .A2(keyinput_g27), .B1(n10265), .B2(
        keyinput_g69), .ZN(n10264) );
  OAI221_X1 U11334 ( .B1(n10483), .B2(keyinput_g27), .C1(n10265), .C2(
        keyinput_g69), .A(n10264), .ZN(n10266) );
  INV_X1 U11335 ( .A(n10266), .ZN(n10271) );
  AOI22_X1 U11336 ( .A1(n6302), .A2(keyinput_g59), .B1(n10404), .B2(
        keyinput_g6), .ZN(n10267) );
  OAI221_X1 U11337 ( .B1(n6302), .B2(keyinput_g59), .C1(n10404), .C2(
        keyinput_g6), .A(n10267), .ZN(n10268) );
  INV_X1 U11338 ( .A(n10268), .ZN(n10270) );
  XNOR2_X1 U11339 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_g117), .ZN(n10269)
         );
  AND4_X1 U11340 ( .A1(n10272), .A2(n10271), .A3(n10270), .A4(n10269), .ZN(
        n10312) );
  AOI22_X1 U11341 ( .A1(n10498), .A2(keyinput_g127), .B1(n10274), .B2(
        keyinput_g62), .ZN(n10273) );
  OAI221_X1 U11342 ( .B1(n10498), .B2(keyinput_g127), .C1(n10274), .C2(
        keyinput_g62), .A(n10273), .ZN(n10286) );
  INV_X1 U11343 ( .A(SI_12_), .ZN(n10276) );
  AOI22_X1 U11344 ( .A1(n6088), .A2(keyinput_g43), .B1(keyinput_g20), .B2(
        n10276), .ZN(n10275) );
  OAI221_X1 U11345 ( .B1(n6088), .B2(keyinput_g43), .C1(n10276), .C2(
        keyinput_g20), .A(n10275), .ZN(n10285) );
  INV_X1 U11346 ( .A(SI_14_), .ZN(n10279) );
  AOI22_X1 U11347 ( .A1(n10279), .A2(keyinput_g18), .B1(n10278), .B2(
        keyinput_g74), .ZN(n10277) );
  OAI221_X1 U11348 ( .B1(n10279), .B2(keyinput_g18), .C1(n10278), .C2(
        keyinput_g74), .A(n10277), .ZN(n10284) );
  INV_X1 U11349 ( .A(SI_0_), .ZN(n10280) );
  XOR2_X1 U11350 ( .A(n10280), .B(keyinput_g32), .Z(n10282) );
  XNOR2_X1 U11351 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g102), .ZN(n10281)
         );
  NAND2_X1 U11352 ( .A1(n10282), .A2(n10281), .ZN(n10283) );
  NOR4_X1 U11353 ( .A1(n10286), .A2(n10285), .A3(n10284), .A4(n10283), .ZN(
        n10311) );
  INV_X1 U11354 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U11355 ( .A1(n5582), .A2(keyinput_g108), .B1(n10288), .B2(
        keyinput_g60), .ZN(n10287) );
  OAI221_X1 U11356 ( .B1(n5582), .B2(keyinput_g108), .C1(n10288), .C2(
        keyinput_g60), .A(n10287), .ZN(n10298) );
  AOI22_X1 U11357 ( .A1(n5175), .A2(keyinput_g118), .B1(n10290), .B2(
        keyinput_g23), .ZN(n10289) );
  OAI221_X1 U11358 ( .B1(n5175), .B2(keyinput_g118), .C1(n10290), .C2(
        keyinput_g23), .A(n10289), .ZN(n10297) );
  INV_X1 U11359 ( .A(SI_10_), .ZN(n10292) );
  AOI22_X1 U11360 ( .A1(n10394), .A2(keyinput_g53), .B1(keyinput_g22), .B2(
        n10292), .ZN(n10291) );
  OAI221_X1 U11361 ( .B1(n10394), .B2(keyinput_g53), .C1(n10292), .C2(
        keyinput_g22), .A(n10291), .ZN(n10296) );
  XNOR2_X1 U11362 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g121), .ZN(n10294)
         );
  XNOR2_X1 U11363 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_g64), .ZN(n10293) );
  NAND2_X1 U11364 ( .A1(n10294), .A2(n10293), .ZN(n10295) );
  NOR4_X1 U11365 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10310) );
  AOI22_X1 U11366 ( .A1(n10508), .A2(keyinput_g77), .B1(n10300), .B2(
        keyinput_g73), .ZN(n10299) );
  OAI221_X1 U11367 ( .B1(n10508), .B2(keyinput_g77), .C1(n10300), .C2(
        keyinput_g73), .A(n10299), .ZN(n10308) );
  INV_X1 U11368 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U11369 ( .A1(n10379), .A2(keyinput_g5), .B1(n10497), .B2(
        keyinput_g63), .ZN(n10301) );
  OAI221_X1 U11370 ( .B1(n10379), .B2(keyinput_g5), .C1(n10497), .C2(
        keyinput_g63), .A(n10301), .ZN(n10307) );
  XOR2_X1 U11371 ( .A(n5584), .B(keyinput_g109), .Z(n10305) );
  XNOR2_X1 U11372 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g96), .ZN(n10304) );
  XNOR2_X1 U11373 ( .A(SI_22_), .B(keyinput_g10), .ZN(n10303) );
  XNOR2_X1 U11374 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_g103), .ZN(n10302)
         );
  NAND4_X1 U11375 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10306) );
  NOR3_X1 U11376 ( .A1(n10308), .A2(n10307), .A3(n10306), .ZN(n10309) );
  NAND4_X1 U11377 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n10309), .ZN(
        n10313) );
  NOR4_X1 U11378 ( .A1(n10316), .A2(n10315), .A3(n10314), .A4(n10313), .ZN(
        n10550) );
  OAI22_X1 U11379 ( .A1(SI_20_), .A2(keyinput_g12), .B1(keyinput_g78), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n10317) );
  AOI221_X1 U11380 ( .B1(SI_20_), .B2(keyinput_g12), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput_g78), .A(n10317), .ZN(n10324)
         );
  OAI22_X1 U11381 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_g94), .B1(
        keyinput_g1), .B2(SI_31_), .ZN(n10318) );
  AOI221_X1 U11382 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_g94), .C1(SI_31_), 
        .C2(keyinput_g1), .A(n10318), .ZN(n10323) );
  OAI22_X1 U11383 ( .A1(SI_24_), .A2(keyinput_g8), .B1(keyinput_g100), .B2(
        P1_IR_REG_10__SCAN_IN), .ZN(n10319) );
  AOI221_X1 U11384 ( .B1(SI_24_), .B2(keyinput_g8), .C1(P1_IR_REG_10__SCAN_IN), 
        .C2(keyinput_g100), .A(n10319), .ZN(n10322) );
  OAI22_X1 U11385 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        keyinput_g120), .B2(P1_IR_REG_30__SCAN_IN), .ZN(n10320) );
  AOI221_X1 U11386 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P1_IR_REG_30__SCAN_IN), .C2(keyinput_g120), .A(n10320), .ZN(n10321) );
  NAND4_X1 U11387 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10353) );
  OAI22_X1 U11388 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_g48), .B1(
        keyinput_g95), .B2(P1_IR_REG_5__SCAN_IN), .ZN(n10325) );
  AOI221_X1 U11389 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_g95), .A(n10325), .ZN(n10332) );
  OAI22_X1 U11390 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(SI_21_), .B2(keyinput_g11), .ZN(n10326) );
  AOI221_X1 U11391 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        keyinput_g11), .C2(SI_21_), .A(n10326), .ZN(n10331) );
  OAI22_X1 U11392 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_g58), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .ZN(n10327) );
  AOI221_X1 U11393 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .C1(
        keyinput_g65), .C2(P2_DATAO_REG_31__SCAN_IN), .A(n10327), .ZN(n10330)
         );
  OAI22_X1 U11394 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(keyinput_g83), .B1(
        keyinput_g24), .B2(SI_8_), .ZN(n10328) );
  AOI221_X1 U11395 ( .B1(P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_g83), .C1(
        SI_8_), .C2(keyinput_g24), .A(n10328), .ZN(n10329) );
  NAND4_X1 U11396 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10352) );
  OAI22_X1 U11397 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        keyinput_g44), .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n10333) );
  AOI221_X1 U11398 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_g44), .A(n10333), .ZN(n10340) );
  OAI22_X1 U11399 ( .A1(SI_19_), .A2(keyinput_g13), .B1(keyinput_g88), .B2(
        P2_DATAO_REG_8__SCAN_IN), .ZN(n10334) );
  AOI221_X1 U11400 ( .B1(SI_19_), .B2(keyinput_g13), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_g88), .A(n10334), .ZN(n10339)
         );
  OAI22_X1 U11401 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_g89), .B1(
        keyinput_g104), .B2(P1_IR_REG_14__SCAN_IN), .ZN(n10335) );
  AOI221_X1 U11402 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_g89), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_g104), .A(n10335), .ZN(n10338) );
  OAI22_X1 U11403 ( .A1(SI_7_), .A2(keyinput_g25), .B1(keyinput_g119), .B2(
        P1_IR_REG_29__SCAN_IN), .ZN(n10336) );
  AOI221_X1 U11404 ( .B1(SI_7_), .B2(keyinput_g25), .C1(P1_IR_REG_29__SCAN_IN), 
        .C2(keyinput_g119), .A(n10336), .ZN(n10337) );
  NAND4_X1 U11405 ( .A1(n10340), .A2(n10339), .A3(n10338), .A4(n10337), .ZN(
        n10351) );
  OAI22_X1 U11406 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_g47), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .ZN(n10341) );
  AOI221_X1 U11407 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .C1(
        keyinput_g84), .C2(P2_DATAO_REG_12__SCAN_IN), .A(n10341), .ZN(n10349)
         );
  OAI22_X1 U11408 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_g111), .B1(
        keyinput_g93), .B2(P1_IR_REG_3__SCAN_IN), .ZN(n10342) );
  AOI221_X1 U11409 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_g111), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput_g93), .A(n10342), .ZN(n10348) );
  OAI22_X1 U11410 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_g113), .B1(
        P1_D_REG_2__SCAN_IN), .B2(keyinput_g124), .ZN(n10343) );
  AOI221_X1 U11411 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_g113), .C1(
        keyinput_g124), .C2(P1_D_REG_2__SCAN_IN), .A(n10343), .ZN(n10347) );
  OAI22_X1 U11412 ( .A1(n10345), .A2(keyinput_g46), .B1(keyinput_g79), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n10344) );
  AOI221_X1 U11413 ( .B1(n10345), .B2(keyinput_g46), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_g79), .A(n10344), .ZN(n10346)
         );
  NAND4_X1 U11414 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n10350) );
  NOR4_X1 U11415 ( .A1(n10353), .A2(n10352), .A3(n10351), .A4(n10350), .ZN(
        n10549) );
  AOI22_X1 U11416 ( .A1(n8412), .A2(keyinput_f41), .B1(keyinput_f33), .B2(
        n5037), .ZN(n10354) );
  OAI221_X1 U11417 ( .B1(n8412), .B2(keyinput_f41), .C1(n5037), .C2(
        keyinput_f33), .A(n10354), .ZN(n10362) );
  XOR2_X1 U11418 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_f100), .Z(n10361) );
  XNOR2_X1 U11419 ( .A(keyinput_f50), .B(n8465), .ZN(n10360) );
  XNOR2_X1 U11420 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_f93), .ZN(n10358) );
  XNOR2_X1 U11421 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_f74), .ZN(n10357) );
  XNOR2_X1 U11422 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_f34), .ZN(n10356) );
  XNOR2_X1 U11423 ( .A(SI_1_), .B(keyinput_f31), .ZN(n10355) );
  NAND4_X1 U11424 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10359) );
  NOR4_X1 U11425 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n10543) );
  AOI22_X1 U11426 ( .A1(n10365), .A2(keyinput_f7), .B1(n10364), .B2(
        keyinput_f38), .ZN(n10363) );
  OAI221_X1 U11427 ( .B1(n10365), .B2(keyinput_f7), .C1(n10364), .C2(
        keyinput_f38), .A(n10363), .ZN(n10377) );
  AOI22_X1 U11428 ( .A1(n10368), .A2(keyinput_f125), .B1(n10367), .B2(
        keyinput_f85), .ZN(n10366) );
  OAI221_X1 U11429 ( .B1(n10368), .B2(keyinput_f125), .C1(n10367), .C2(
        keyinput_f85), .A(n10366), .ZN(n10376) );
  AOI22_X1 U11430 ( .A1(n10371), .A2(keyinput_f78), .B1(keyinput_f2), .B2(
        n10370), .ZN(n10369) );
  OAI221_X1 U11431 ( .B1(n10371), .B2(keyinput_f78), .C1(n10370), .C2(
        keyinput_f2), .A(n10369), .ZN(n10375) );
  XNOR2_X1 U11432 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_f75), .ZN(n10373) );
  XNOR2_X1 U11433 ( .A(SI_4_), .B(keyinput_f28), .ZN(n10372) );
  NAND2_X1 U11434 ( .A1(n10373), .A2(n10372), .ZN(n10374) );
  NOR4_X1 U11435 ( .A1(n10377), .A2(n10376), .A3(n10375), .A4(n10374), .ZN(
        n10542) );
  OAI22_X1 U11436 ( .A1(n10380), .A2(keyinput_f55), .B1(n10379), .B2(
        keyinput_f5), .ZN(n10378) );
  AOI221_X1 U11437 ( .B1(n10380), .B2(keyinput_f55), .C1(keyinput_f5), .C2(
        n10379), .A(n10378), .ZN(n10392) );
  OAI22_X1 U11438 ( .A1(n10382), .A2(keyinput_f89), .B1(n5582), .B2(
        keyinput_f108), .ZN(n10381) );
  AOI221_X1 U11439 ( .B1(n10382), .B2(keyinput_f89), .C1(keyinput_f108), .C2(
        n5582), .A(n10381), .ZN(n10391) );
  OAI22_X1 U11440 ( .A1(n10385), .A2(keyinput_f83), .B1(n10384), .B2(
        keyinput_f54), .ZN(n10383) );
  AOI221_X1 U11441 ( .B1(n10385), .B2(keyinput_f83), .C1(keyinput_f54), .C2(
        n10384), .A(n10383), .ZN(n10390) );
  OAI22_X1 U11442 ( .A1(n10388), .A2(keyinput_f8), .B1(n10387), .B2(
        keyinput_f122), .ZN(n10386) );
  AOI221_X1 U11443 ( .B1(n10388), .B2(keyinput_f8), .C1(keyinput_f122), .C2(
        n10387), .A(n10386), .ZN(n10389) );
  NAND4_X1 U11444 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10408) );
  AOI22_X1 U11445 ( .A1(n10394), .A2(keyinput_f53), .B1(keyinput_f43), .B2(
        n6088), .ZN(n10393) );
  OAI221_X1 U11446 ( .B1(n10394), .B2(keyinput_f53), .C1(n6088), .C2(
        keyinput_f43), .A(n10393), .ZN(n10398) );
  XOR2_X1 U11447 ( .A(keyinput_f0), .B(P2_WR_REG_SCAN_IN), .Z(n10397) );
  XNOR2_X1 U11448 ( .A(n10395), .B(keyinput_f30), .ZN(n10396) );
  OR3_X1 U11449 ( .A1(n10398), .A2(n10397), .A3(n10396), .ZN(n10407) );
  AOI22_X1 U11450 ( .A1(n10401), .A2(keyinput_f80), .B1(n10400), .B2(
        keyinput_f35), .ZN(n10399) );
  OAI221_X1 U11451 ( .B1(n10401), .B2(keyinput_f80), .C1(n10400), .C2(
        keyinput_f35), .A(n10399), .ZN(n10406) );
  AOI22_X1 U11452 ( .A1(n10404), .A2(keyinput_f6), .B1(keyinput_f81), .B2(
        n10403), .ZN(n10402) );
  OAI221_X1 U11453 ( .B1(n10404), .B2(keyinput_f6), .C1(n10403), .C2(
        keyinput_f81), .A(n10402), .ZN(n10405) );
  NOR4_X1 U11454 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10541) );
  OAI22_X1 U11455 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput_f64), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_f95), .ZN(n10409) );
  AOI221_X1 U11456 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput_f64), .C1(
        keyinput_f95), .C2(P1_IR_REG_5__SCAN_IN), .A(n10409), .ZN(n10416) );
  OAI22_X1 U11457 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_f71), .ZN(n10410) );
  AOI221_X1 U11458 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        keyinput_f71), .C2(P2_DATAO_REG_25__SCAN_IN), .A(n10410), .ZN(n10415)
         );
  OAI22_X1 U11459 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        keyinput_f113), .B2(P1_IR_REG_23__SCAN_IN), .ZN(n10411) );
  AOI221_X1 U11460 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_f113), .A(n10411), .ZN(n10414) );
  OAI22_X1 U11461 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_f111), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(keyinput_f120), .ZN(n10412) );
  AOI221_X1 U11462 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_f111), .C1(
        keyinput_f120), .C2(P1_IR_REG_30__SCAN_IN), .A(n10412), .ZN(n10413) );
  NAND4_X1 U11463 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10539) );
  AOI22_X1 U11464 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f91), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .ZN(n10417) );
  OAI221_X1 U11465 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f91), .C1(
        P2_DATAO_REG_20__SCAN_IN), .C2(keyinput_f76), .A(n10417), .ZN(n10424)
         );
  AOI22_X1 U11466 ( .A1(SI_7_), .A2(keyinput_f25), .B1(SI_21_), .B2(
        keyinput_f11), .ZN(n10418) );
  OAI221_X1 U11467 ( .B1(SI_7_), .B2(keyinput_f25), .C1(SI_21_), .C2(
        keyinput_f11), .A(n10418), .ZN(n10423) );
  AOI22_X1 U11468 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_f102), .B1(SI_20_), .B2(keyinput_f12), .ZN(n10419) );
  OAI221_X1 U11469 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_f102), .C1(
        SI_20_), .C2(keyinput_f12), .A(n10419), .ZN(n10422) );
  AOI22_X1 U11470 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .ZN(n10420) );
  OAI221_X1 U11471 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput_f86), .A(n10420), .ZN(n10421)
         );
  NOR4_X1 U11472 ( .A1(n10424), .A2(n10423), .A3(n10422), .A4(n10421), .ZN(
        n10442) );
  AOI22_X1 U11473 ( .A1(SI_10_), .A2(keyinput_f22), .B1(SI_17_), .B2(
        keyinput_f15), .ZN(n10425) );
  OAI221_X1 U11474 ( .B1(SI_10_), .B2(keyinput_f22), .C1(SI_17_), .C2(
        keyinput_f15), .A(n10425), .ZN(n10432) );
  AOI22_X1 U11475 ( .A1(SI_19_), .A2(keyinput_f13), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n10426) );
  OAI221_X1 U11476 ( .B1(SI_19_), .B2(keyinput_f13), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n10426), .ZN(n10431)
         );
  AOI22_X1 U11477 ( .A1(SI_16_), .A2(keyinput_f16), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n10427) );
  OAI221_X1 U11478 ( .B1(SI_16_), .B2(keyinput_f16), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n10427), .ZN(n10430)
         );
  AOI22_X1 U11479 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_f88), .B1(SI_8_), .B2(keyinput_f24), .ZN(n10428) );
  OAI221_X1 U11480 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .C1(
        SI_8_), .C2(keyinput_f24), .A(n10428), .ZN(n10429) );
  NOR4_X1 U11481 ( .A1(n10432), .A2(n10431), .A3(n10430), .A4(n10429), .ZN(
        n10441) );
  OAI22_X1 U11482 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        keyinput_f57), .B2(P2_REG3_REG_22__SCAN_IN), .ZN(n10433) );
  AOI221_X1 U11483 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n10433), .ZN(n10439)
         );
  OAI22_X1 U11484 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_f82), .B1(
        keyinput_f1), .B2(SI_31_), .ZN(n10434) );
  AOI221_X1 U11485 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .C1(
        SI_31_), .C2(keyinput_f1), .A(n10434), .ZN(n10438) );
  OAI22_X1 U11486 ( .A1(SI_15_), .A2(keyinput_f17), .B1(P1_D_REG_4__SCAN_IN), 
        .B2(keyinput_f126), .ZN(n10435) );
  AOI221_X1 U11487 ( .B1(SI_15_), .B2(keyinput_f17), .C1(keyinput_f126), .C2(
        P1_D_REG_4__SCAN_IN), .A(n10435), .ZN(n10437) );
  XNOR2_X1 U11488 ( .A(SI_3_), .B(keyinput_f29), .ZN(n10436) );
  AND4_X1 U11489 ( .A1(n10439), .A2(n10438), .A3(n10437), .A4(n10436), .ZN(
        n10440) );
  NAND3_X1 U11490 ( .A1(n10442), .A2(n10441), .A3(n10440), .ZN(n10538) );
  AOI22_X1 U11491 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_f116), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_f97), .ZN(n10443) );
  OAI221_X1 U11492 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_f116), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput_f97), .A(n10443), .ZN(n10450) );
  AOI22_X1 U11493 ( .A1(SI_9_), .A2(keyinput_f23), .B1(SI_12_), .B2(
        keyinput_f20), .ZN(n10444) );
  OAI221_X1 U11494 ( .B1(SI_9_), .B2(keyinput_f23), .C1(SI_12_), .C2(
        keyinput_f20), .A(n10444), .ZN(n10449) );
  AOI22_X1 U11495 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_f109), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .ZN(n10445) );
  OAI221_X1 U11496 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_f109), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n10445), .ZN(n10448) );
  AOI22_X1 U11497 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_f94), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n10446) );
  OAI221_X1 U11498 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_f94), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n10446), .ZN(n10447)
         );
  NOR4_X1 U11499 ( .A1(n10450), .A2(n10449), .A3(n10448), .A4(n10447), .ZN(
        n10478) );
  AOI22_X1 U11500 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_f99), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .ZN(n10451) );
  OAI221_X1 U11501 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_f99), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_f69), .A(n10451), .ZN(n10458)
         );
  AOI22_X1 U11502 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_f117), .B1(SI_14_), .B2(keyinput_f18), .ZN(n10452) );
  OAI221_X1 U11503 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_f117), .C1(
        SI_14_), .C2(keyinput_f18), .A(n10452), .ZN(n10457) );
  AOI22_X1 U11504 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f118), .B1(SI_11_), .B2(keyinput_f21), .ZN(n10453) );
  OAI221_X1 U11505 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f118), .C1(
        SI_11_), .C2(keyinput_f21), .A(n10453), .ZN(n10456) );
  AOI22_X1 U11506 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_f98), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .ZN(n10454) );
  OAI221_X1 U11507 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput_f98), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput_f67), .A(n10454), .ZN(n10455)
         );
  NOR4_X1 U11508 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10477) );
  AOI22_X1 U11509 ( .A1(SI_18_), .A2(keyinput_f14), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .ZN(n10459) );
  OAI221_X1 U11510 ( .B1(SI_18_), .B2(keyinput_f14), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n10459), .ZN(n10466)
         );
  AOI22_X1 U11511 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_f68), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n10460) );
  OAI221_X1 U11512 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_f68), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n10460), .ZN(n10465)
         );
  AOI22_X1 U11513 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_f114), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_f106), .ZN(n10461) );
  OAI221_X1 U11514 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_f114), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_f106), .A(n10461), .ZN(n10464) );
  AOI22_X1 U11515 ( .A1(SI_0_), .A2(keyinput_f32), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .ZN(n10462) );
  OAI221_X1 U11516 ( .B1(SI_0_), .B2(keyinput_f32), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_f70), .A(n10462), .ZN(n10463)
         );
  NOR4_X1 U11517 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10476) );
  AOI22_X1 U11518 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_f79), .B1(
        P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .ZN(n10467) );
  OAI221_X1 U11519 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_f79), .C1(
        P2_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n10467), .ZN(n10474) );
  AOI22_X1 U11520 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput_f96), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n10468) );
  OAI221_X1 U11521 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput_f96), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n10468), .ZN(n10473)
         );
  AOI22_X1 U11522 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_f87), .B1(
        SI_23_), .B2(keyinput_f9), .ZN(n10469) );
  OAI221_X1 U11523 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .C1(
        SI_23_), .C2(keyinput_f9), .A(n10469), .ZN(n10472) );
  AOI22_X1 U11524 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f103), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_f107), .ZN(n10470) );
  OAI221_X1 U11525 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f103), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_f107), .A(n10470), .ZN(n10471) );
  NOR4_X1 U11526 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10475) );
  NAND4_X1 U11527 ( .A1(n10478), .A2(n10477), .A3(n10476), .A4(n10475), .ZN(
        n10537) );
  AOI22_X1 U11528 ( .A1(n10481), .A2(keyinput_f19), .B1(n10480), .B2(
        keyinput_f56), .ZN(n10479) );
  OAI221_X1 U11529 ( .B1(n10481), .B2(keyinput_f19), .C1(n10480), .C2(
        keyinput_f56), .A(n10479), .ZN(n10492) );
  AOI22_X1 U11530 ( .A1(n10484), .A2(keyinput_f10), .B1(keyinput_f27), .B2(
        n10483), .ZN(n10482) );
  OAI221_X1 U11531 ( .B1(n10484), .B2(keyinput_f10), .C1(n10483), .C2(
        keyinput_f27), .A(n10482), .ZN(n10491) );
  AOI22_X1 U11532 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_f73), .B1(
        n10486), .B2(keyinput_f52), .ZN(n10485) );
  OAI221_X1 U11533 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .C1(
        n10486), .C2(keyinput_f52), .A(n10485), .ZN(n10490) );
  XNOR2_X1 U11534 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_f101), .ZN(n10488)
         );
  XNOR2_X1 U11535 ( .A(SI_6_), .B(keyinput_f26), .ZN(n10487) );
  NAND2_X1 U11536 ( .A1(n10488), .A2(n10487), .ZN(n10489) );
  NOR4_X1 U11537 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10535) );
  AOI22_X1 U11538 ( .A1(n10495), .A2(keyinput_f72), .B1(n10494), .B2(
        keyinput_f39), .ZN(n10493) );
  OAI221_X1 U11539 ( .B1(n10495), .B2(keyinput_f72), .C1(n10494), .C2(
        keyinput_f39), .A(n10493), .ZN(n10505) );
  AOI22_X1 U11540 ( .A1(n10498), .A2(keyinput_f127), .B1(n10497), .B2(
        keyinput_f63), .ZN(n10496) );
  OAI221_X1 U11541 ( .B1(n10498), .B2(keyinput_f127), .C1(n10497), .C2(
        keyinput_f63), .A(n10496), .ZN(n10504) );
  XNOR2_X1 U11542 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_f90), .ZN(n10502) );
  XNOR2_X1 U11543 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f110), .ZN(n10501)
         );
  XNOR2_X1 U11544 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_f119), .ZN(n10500)
         );
  XNOR2_X1 U11545 ( .A(keyinput_f59), .B(P2_REG3_REG_2__SCAN_IN), .ZN(n10499)
         );
  NAND4_X1 U11546 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10503) );
  NOR3_X1 U11547 ( .A1(n10505), .A2(n10504), .A3(n10503), .ZN(n10534) );
  INV_X1 U11548 ( .A(SI_29_), .ZN(n10507) );
  AOI22_X1 U11549 ( .A1(n10508), .A2(keyinput_f77), .B1(n10507), .B2(
        keyinput_f3), .ZN(n10506) );
  OAI221_X1 U11550 ( .B1(n10508), .B2(keyinput_f77), .C1(n10507), .C2(
        keyinput_f3), .A(n10506), .ZN(n10518) );
  AOI22_X1 U11551 ( .A1(n5169), .A2(keyinput_f104), .B1(keyinput_f105), .B2(
        n4919), .ZN(n10509) );
  OAI221_X1 U11552 ( .B1(n5169), .B2(keyinput_f104), .C1(n4919), .C2(
        keyinput_f105), .A(n10509), .ZN(n10517) );
  AOI22_X1 U11553 ( .A1(n5949), .A2(keyinput_f112), .B1(n10511), .B2(
        keyinput_f84), .ZN(n10510) );
  OAI221_X1 U11554 ( .B1(n5949), .B2(keyinput_f112), .C1(n10511), .C2(
        keyinput_f84), .A(n10510), .ZN(n10516) );
  XOR2_X1 U11555 ( .A(n10512), .B(keyinput_f123), .Z(n10514) );
  XNOR2_X1 U11556 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f121), .ZN(n10513)
         );
  NAND2_X1 U11557 ( .A1(n10514), .A2(n10513), .ZN(n10515) );
  NOR4_X1 U11558 ( .A1(n10518), .A2(n10517), .A3(n10516), .A4(n10515), .ZN(
        n10533) );
  AOI22_X1 U11559 ( .A1(n10520), .A2(keyinput_f4), .B1(keyinput_f44), .B2(
        n9994), .ZN(n10519) );
  OAI221_X1 U11560 ( .B1(n10520), .B2(keyinput_f4), .C1(n9994), .C2(
        keyinput_f44), .A(n10519), .ZN(n10531) );
  AOI22_X1 U11561 ( .A1(n10523), .A2(keyinput_f58), .B1(keyinput_f66), .B2(
        n10522), .ZN(n10521) );
  OAI221_X1 U11562 ( .B1(n10523), .B2(keyinput_f58), .C1(n10522), .C2(
        keyinput_f66), .A(n10521), .ZN(n10530) );
  XNOR2_X1 U11563 ( .A(n10524), .B(keyinput_f124), .ZN(n10529) );
  XNOR2_X1 U11564 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_f115), .ZN(n10527)
         );
  XNOR2_X1 U11565 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_f51), .ZN(n10526)
         );
  XNOR2_X1 U11566 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_f92), .ZN(n10525) );
  NAND3_X1 U11567 ( .A1(n10527), .A2(n10526), .A3(n10525), .ZN(n10528) );
  NOR4_X1 U11568 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10532) );
  NAND4_X1 U11569 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10536) );
  NOR4_X1 U11570 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10540) );
  NAND4_X1 U11571 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10545) );
  AOI21_X1 U11572 ( .B1(keyinput_f45), .B2(n10545), .A(keyinput_g45), .ZN(
        n10547) );
  INV_X1 U11573 ( .A(keyinput_f45), .ZN(n10544) );
  AOI21_X1 U11574 ( .B1(n10545), .B2(n10544), .A(n8431), .ZN(n10546) );
  AOI22_X1 U11575 ( .A1(n8431), .A2(n10547), .B1(keyinput_g45), .B2(n10546), 
        .ZN(n10548) );
  AOI21_X1 U11576 ( .B1(n10550), .B2(n10549), .A(n10548), .ZN(n10553) );
  XNOR2_X1 U11577 ( .A(n10551), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n10552) );
  XNOR2_X1 U11578 ( .A(n10553), .B(n10552), .ZN(n10554) );
  XNOR2_X1 U11579 ( .A(n10555), .B(n10554), .ZN(ADD_1068_U4) );
  XNOR2_X1 U11580 ( .A(n10557), .B(n10556), .ZN(ADD_1068_U47) );
  XOR2_X1 U11581 ( .A(n10559), .B(n10558), .Z(ADD_1068_U54) );
  XNOR2_X1 U11582 ( .A(n10561), .B(n10560), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11583 ( .A(n10563), .B(n10562), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11584 ( .A(n10565), .B(n10564), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11585 ( .A(n10567), .B(n10566), .ZN(ADD_1068_U50) );
  XOR2_X1 U11586 ( .A(n10569), .B(n10568), .Z(ADD_1068_U53) );
  XNOR2_X1 U11587 ( .A(n10571), .B(n10570), .ZN(ADD_1068_U52) );
  INV_X2 U5062 ( .A(n8277), .ZN(n9152) );
  NAND2_X1 U5144 ( .A1(n8565), .A2(n6679), .ZN(n6502) );
endmodule

