

module b21_C_SARLock_k_64_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10043;

  NOR2_X1 U4769 ( .A1(n8144), .A2(n8145), .ZN(n8143) );
  INV_X2 U4770 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X2 U4771 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  CLKBUF_X2 U4772 ( .A(n5763), .Z(n8041) );
  INV_X1 U4773 ( .A(n8009), .ZN(n7989) );
  CLKBUF_X1 U4774 ( .A(n6512), .Z(n4264) );
  NAND2_X2 U4775 ( .A1(n9810), .A2(n8236), .ZN(n5763) );
  CLKBUF_X2 U4776 ( .A(n5686), .Z(n8732) );
  AND4_X1 U4778 ( .A1(n5579), .A2(n6003), .A3(n5128), .A4(n4825), .ZN(n4306)
         );
  INV_X1 U4780 ( .A(n8043), .ZN(n7439) );
  NAND2_X1 U4781 ( .A1(n7581), .A2(n7583), .ZN(n7715) );
  INV_X1 U4782 ( .A(n5691), .ZN(n4275) );
  AND2_X1 U4784 ( .A1(n4433), .A2(n4429), .ZN(n4430) );
  OR3_X2 U4785 ( .A1(n9125), .A2(n9238), .A3(n4482), .ZN(n4300) );
  AND2_X1 U4786 ( .A1(n9047), .A2(n8871), .ZN(n9022) );
  INV_X1 U4787 ( .A(n9584), .ZN(n9655) );
  NAND2_X1 U4788 ( .A1(n4304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5013) );
  AND4_X1 U4789 ( .A1(n5476), .A2(n5475), .A3(n5474), .A4(n5473), .ZN(n6023)
         );
  NOR2_X2 U4790 ( .A1(n9235), .A2(n4300), .ZN(n9056) );
  NAND4_X1 U4791 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n8158)
         );
  INV_X1 U4792 ( .A(n5118), .ZN(n7747) );
  INV_X1 U4793 ( .A(n8932), .ZN(n6395) );
  NAND2_X2 U4794 ( .A1(n5127), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U4795 ( .A1(n5742), .A2(n6106), .ZN(n4263) );
  OR2_X2 U4796 ( .A1(n5593), .A2(n9774), .ZN(n7580) );
  NAND4_X2 U4797 ( .A1(n5114), .A2(n5113), .A3(n5112), .A4(n5111), .ZN(n5593)
         );
  OAI22_X2 U4798 ( .A1(n9004), .A2(n9003), .B1(n9002), .B2(n9001), .ZN(n9212)
         );
  AOI21_X2 U4799 ( .B1(n4569), .B2(n4571), .A(n4568), .ZN(n9004) );
  AOI21_X2 U4800 ( .B1(n6974), .B2(n6973), .A(n6972), .ZN(n7127) );
  NAND2_X2 U4801 ( .A1(n4733), .A2(n4731), .ZN(n6974) );
  INV_X1 U4802 ( .A(n5609), .ZN(n7458) );
  OAI211_X1 U4803 ( .C1(n5364), .C2(n6044), .A(n6043), .B(n6042), .ZN(n6512)
         );
  OR2_X2 U4804 ( .A1(n8418), .A2(n6109), .ZN(n7581) );
  XNOR2_X2 U4805 ( .A(n5013), .B(n5012), .ZN(n7756) );
  CLKBUF_X1 U4806 ( .A(n9107), .Z(n4273) );
  NAND2_X1 U4807 ( .A1(n8639), .A2(n8642), .ZN(n7820) );
  NAND2_X1 U4808 ( .A1(n9275), .A2(n4341), .ZN(n9152) );
  NAND2_X1 U4809 ( .A1(n7512), .A2(n7511), .ZN(n8435) );
  OAI21_X1 U4810 ( .B1(n7127), .B2(n7126), .A(n7125), .ZN(n4419) );
  NOR2_X1 U4811 ( .A1(n4266), .A2(n4774), .ZN(n4773) );
  INV_X1 U4812 ( .A(n6233), .ZN(n4266) );
  OR2_X1 U4813 ( .A1(n7246), .A2(n8603), .ZN(n7278) );
  NAND2_X2 U4814 ( .A1(n7567), .A2(n7589), .ZN(n6140) );
  INV_X1 U4815 ( .A(n9609), .ZN(n8952) );
  INV_X2 U4816 ( .A(n7900), .ZN(n6561) );
  INV_X4 U4817 ( .A(n6180), .ZN(n4265) );
  NAND2_X1 U4818 ( .A1(n7757), .A2(n8253), .ZN(n5740) );
  AND3_X1 U4819 ( .A1(n5135), .A2(n6395), .A3(n4450), .ZN(n5676) );
  INV_X1 U4820 ( .A(n6022), .ZN(n6028) );
  INV_X2 U4821 ( .A(n7697), .ZN(n7710) );
  XNOR2_X1 U4822 ( .A(n5097), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8253) );
  BUF_X2 U4823 ( .A(n5775), .Z(n7518) );
  AND2_X1 U4824 ( .A1(n5029), .A2(n5030), .ZN(n5038) );
  OAI21_X1 U4825 ( .B1(n4923), .B2(n4596), .A(n4931), .ZN(n4595) );
  CLKBUF_X2 U4826 ( .A(n4834), .Z(n5340) );
  NAND2_X1 U4827 ( .A1(n4748), .A2(n4747), .ZN(n8653) );
  NOR2_X1 U4828 ( .A1(n4432), .A2(n4430), .ZN(n8610) );
  AND2_X1 U4829 ( .A1(n4422), .A2(n7939), .ZN(n4421) );
  OR2_X1 U4830 ( .A1(n8445), .A2(n4385), .ZN(n8523) );
  NOR2_X1 U4831 ( .A1(n9080), .A2(n9022), .ZN(n9023) );
  OR2_X1 U4832 ( .A1(n8063), .A2(n7416), .ZN(n7422) );
  NAND2_X1 U4833 ( .A1(n8130), .A2(n7393), .ZN(n7417) );
  AOI211_X1 U4834 ( .C1(n9632), .C2(n9373), .A(n9372), .B(n9371), .ZN(n9416)
         );
  OAI21_X1 U4835 ( .B1(n7337), .B2(n4674), .A(n4672), .ZN(n7390) );
  NAND2_X1 U4836 ( .A1(n4556), .A2(n4311), .ZN(n9275) );
  INV_X1 U4837 ( .A(n9022), .ZN(n9082) );
  NAND2_X1 U4838 ( .A1(n9238), .A2(n8941), .ZN(n9024) );
  NAND2_X1 U4839 ( .A1(n7138), .A2(n7137), .ZN(n7163) );
  NAND2_X1 U4840 ( .A1(n7982), .A2(n7981), .ZN(n9245) );
  AND2_X1 U4841 ( .A1(n7161), .A2(n7160), .ZN(n7162) );
  XNOR2_X1 U4842 ( .A(n7510), .B(n7509), .ZN(n9324) );
  NAND2_X1 U4843 ( .A1(n7131), .A2(n7132), .ZN(n7161) );
  OAI21_X1 U4844 ( .B1(n7182), .B2(n4373), .A(n4371), .ZN(n8372) );
  NOR2_X1 U4845 ( .A1(n6822), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U4846 ( .A1(n6532), .A2(n6531), .ZN(n6657) );
  AOI21_X1 U4847 ( .B1(n6689), .B2(n6690), .A(n4314), .ZN(n4734) );
  AND2_X1 U4848 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  AND2_X1 U4849 ( .A1(n8701), .A2(n8675), .ZN(n8903) );
  NOR2_X1 U4850 ( .A1(n6196), .A2(n4741), .ZN(n4740) );
  INV_X2 U4851 ( .A(n9825), .ZN(n4267) );
  INV_X2 U4852 ( .A(n9833), .ZN(n4268) );
  NAND2_X1 U4853 ( .A1(n6366), .A2(n6365), .ZN(n6562) );
  AND2_X1 U4854 ( .A1(n8809), .A2(n8754), .ZN(n8904) );
  OAI21_X1 U4855 ( .B1(n5631), .B2(n5630), .A(n5629), .ZN(n5845) );
  NAND2_X1 U4856 ( .A1(n6371), .A2(n6370), .ZN(n6595) );
  INV_X2 U4857 ( .A(n9697), .ZN(n4269) );
  AND3_X1 U4858 ( .A1(n5928), .A2(n5927), .A3(n5926), .ZN(n9790) );
  INV_X1 U4859 ( .A(n7974), .ZN(n8012) );
  INV_X2 U4860 ( .A(n5663), .ZN(n8009) );
  INV_X1 U4861 ( .A(n6415), .ZN(n8951) );
  OR2_X1 U4862 ( .A1(n6931), .A2(n6930), .ZN(n7100) );
  AND3_X1 U4863 ( .A1(n5774), .A2(n5773), .A3(n5772), .ZN(n6118) );
  NAND2_X1 U4864 ( .A1(n5465), .A2(n5464), .ZN(n6083) );
  AND4_X1 U4865 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n9609)
         );
  AND4_X1 U4866 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n6415)
         );
  AND4_X1 U4867 ( .A1(n6052), .A2(n6051), .A3(n6050), .A4(n6049), .ZN(n9593)
         );
  NAND2_X1 U4868 ( .A1(n4592), .A2(n4590), .ZN(n4950) );
  AND2_X1 U4869 ( .A1(n5463), .A2(n5984), .ZN(n5465) );
  INV_X1 U4870 ( .A(n6031), .ZN(n9641) );
  NAND2_X1 U4871 ( .A1(n5614), .A2(n5613), .ZN(n8159) );
  INV_X1 U4872 ( .A(n5469), .ZN(n8682) );
  CLKBUF_X1 U4873 ( .A(n5356), .Z(n8931) );
  INV_X2 U4874 ( .A(n5691), .ZN(n7826) );
  NAND2_X1 U4875 ( .A1(n4924), .A2(n4593), .ZN(n4592) );
  INV_X1 U4876 ( .A(n5741), .ZN(n5617) );
  AND4_X1 U4877 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(n6663)
         );
  NAND2_X1 U4878 ( .A1(n4377), .A2(n4912), .ZN(n4924) );
  NAND4_X1 U4879 ( .A1(n5599), .A2(n5598), .A3(n5597), .A4(n5596), .ZN(n8418)
         );
  AND3_X2 U4880 ( .A1(n5461), .A2(n5460), .A3(n5459), .ZN(n5469) );
  INV_X1 U4881 ( .A(n5472), .ZN(n5691) );
  AND2_X1 U4882 ( .A1(n5135), .A2(n5134), .ZN(n5356) );
  AND3_X2 U4883 ( .A1(n5592), .A2(n5591), .A3(n5590), .ZN(n9774) );
  AND3_X1 U4884 ( .A1(n5605), .A2(n5604), .A3(n5603), .ZN(n6109) );
  OR2_X1 U4885 ( .A1(n5685), .A2(n5671), .ZN(n5674) );
  NAND2_X1 U4886 ( .A1(n4652), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U4887 ( .A1(n4902), .A2(n4901), .ZN(n4909) );
  INV_X1 U4888 ( .A(n5970), .ZN(n5108) );
  INV_X2 U4889 ( .A(n7445), .ZN(n7320) );
  AOI21_X1 U4890 ( .B1(n4959), .B2(n4636), .A(n4634), .ZN(n4633) );
  OAI21_X1 U4891 ( .B1(n4595), .B2(n4927), .A(n4325), .ZN(n4591) );
  NAND2_X1 U4892 ( .A1(n4854), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5016) );
  AND2_X2 U4893 ( .A1(n5101), .A2(n8057), .ZN(n5595) );
  INV_X1 U4894 ( .A(n8058), .ZN(n5032) );
  INV_X1 U4895 ( .A(n4927), .ZN(n4596) );
  NAND2_X1 U4896 ( .A1(n5092), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6008) );
  NOR2_X1 U4897 ( .A1(n5092), .A2(n4852), .ZN(n5017) );
  XNOR2_X1 U4898 ( .A(n5031), .B(n4487), .ZN(n8058) );
  MUX2_X1 U4899 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5026), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5029) );
  NAND2_X1 U4900 ( .A1(n4911), .A2(SI_3_), .ZN(n4912) );
  XNOR2_X1 U4901 ( .A(n5368), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9588) );
  XNOR2_X1 U4902 ( .A(n4987), .B(n9995), .ZN(n8057) );
  NAND2_X1 U4903 ( .A1(n5030), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5031) );
  OR2_X1 U4904 ( .A1(n8537), .A2(n4853), .ZN(n4985) );
  XNOR2_X1 U4905 ( .A(n4933), .B(SI_5_), .ZN(n4930) );
  INV_X2 U4906 ( .A(n9323), .ZN(n8059) );
  NAND2_X1 U4907 ( .A1(n5587), .A2(P1_U3084), .ZN(n9328) );
  AND3_X1 U4908 ( .A1(n4870), .A2(n4869), .A3(n4334), .ZN(n5009) );
  INV_X2 U4909 ( .A(n6728), .ZN(n4270) );
  NOR2_X1 U4910 ( .A1(n4920), .A2(n4847), .ZN(n4870) );
  NAND2_X1 U4911 ( .A1(n4875), .A2(n4805), .ZN(n4804) );
  AND2_X1 U4912 ( .A1(n4884), .A2(n4818), .ZN(n4913) );
  INV_X1 U4913 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5128) );
  NOR2_X1 U4914 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4818) );
  OR2_X1 U4915 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4272) );
  INV_X1 U4916 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U4917 ( .A1(n4486), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4271) );
  INV_X1 U4918 ( .A(n7094), .ZN(n4274) );
  NOR2_X1 U4919 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4884) );
  AOI21_X1 U4920 ( .B1(n6942), .B2(n6941), .A(n6940), .ZN(n7091) );
  NAND2_X1 U4921 ( .A1(n9131), .A2(n9130), .ZN(n9258) );
  AOI22_X1 U4922 ( .A1(n9136), .A2(n9013), .B1(n9012), .B2(n9149), .ZN(n9131)
         );
  NAND2_X1 U4923 ( .A1(n6090), .A2(n6089), .ZN(n9580) );
  NAND2_X2 U4924 ( .A1(n5356), .A2(n6395), .ZN(n5359) );
  NOR2_X2 U4925 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4890) );
  NAND2_X1 U4926 ( .A1(n6083), .A2(n6082), .ZN(n6427) );
  AOI22_X2 U4927 ( .A1(n9212), .A2(n9211), .B1(n9205), .B2(n9292), .ZN(n9194)
         );
  OR2_X1 U4928 ( .A1(n5685), .A2(n6034), .ZN(n6037) );
  INV_X4 U4929 ( .A(n5587), .ZN(n4276) );
  NAND4_X2 U4930 ( .A1(n5398), .A2(n5397), .A3(n5396), .A4(n5395), .ZN(n5462)
         );
  OAI21_X1 U4931 ( .B1(n6427), .B2(n8897), .A(n6084), .ZN(n9599) );
  NAND2_X2 U4932 ( .A1(n6614), .A2(n8824), .ZN(n6877) );
  INV_X1 U4933 ( .A(n7445), .ZN(n4277) );
  AND2_X1 U4934 ( .A1(n5101), .A2(n8057), .ZN(n4278) );
  AND2_X1 U4935 ( .A1(n5101), .A2(n8057), .ZN(n4279) );
  NOR2_X1 U4936 ( .A1(n6433), .A2(n6022), .ZN(n9601) );
  AND2_X1 U4937 ( .A1(n5032), .A2(n5038), .ZN(n4280) );
  AND2_X1 U4938 ( .A1(n5032), .A2(n5038), .ZN(n4281) );
  AND2_X1 U4939 ( .A1(n5032), .A2(n5038), .ZN(n5712) );
  XNOR2_X2 U4940 ( .A(n4985), .B(n4984), .ZN(n4988) );
  AOI21_X1 U4941 ( .B1(n5355), .B2(n5128), .A(n4915), .ZN(n5133) );
  NAND2_X1 U4942 ( .A1(n4619), .A2(n4618), .ZN(n7515) );
  AOI21_X1 U4943 ( .B1(n4621), .B2(n4623), .A(n4354), .ZN(n4618) );
  OAI21_X1 U4944 ( .B1(n7058), .B2(n7057), .A(n7056), .ZN(n7117) );
  NAND2_X1 U4945 ( .A1(n4597), .A2(n4598), .ZN(n5631) );
  INV_X1 U4946 ( .A(n4599), .ZN(n4598) );
  OAI21_X1 U4947 ( .B1(n4602), .B2(n4600), .A(n5572), .ZN(n4599) );
  NOR3_X1 U4948 ( .A1(n8233), .A2(n8435), .A3(n4547), .ZN(n8184) );
  NAND2_X1 U4949 ( .A1(n7787), .A2(n7507), .ZN(n4547) );
  NAND2_X1 U4950 ( .A1(n4767), .A2(n4766), .ZN(n8206) );
  AOI21_X1 U4951 ( .B1(n4768), .B2(n4730), .A(n8214), .ZN(n4766) );
  INV_X1 U4952 ( .A(n8732), .ZN(n7823) );
  INV_X1 U4953 ( .A(n5364), .ZN(n7822) );
  OR2_X1 U4954 ( .A1(n7376), .A2(n4418), .ZN(n4674) );
  OR2_X1 U4955 ( .A1(n8124), .A2(n4676), .ZN(n4418) );
  INV_X1 U4956 ( .A(n7347), .ZN(n4676) );
  INV_X1 U4957 ( .A(n7605), .ZN(n4700) );
  AND2_X1 U4958 ( .A1(n4633), .A2(n4414), .ZN(n4411) );
  NAND2_X1 U4959 ( .A1(n4948), .A2(n4952), .ZN(n4414) );
  NOR2_X1 U4960 ( .A1(n4995), .A2(n4637), .ZN(n4636) );
  INV_X1 U4961 ( .A(n4963), .ZN(n4637) );
  NAND2_X1 U4962 ( .A1(n4966), .A2(n4965), .ZN(n4994) );
  NAND2_X1 U4963 ( .A1(n7544), .A2(n7543), .ZN(n7709) );
  INV_X1 U4964 ( .A(n8427), .ZN(n7544) );
  INV_X1 U4965 ( .A(n7782), .ZN(n7788) );
  NOR2_X1 U4966 ( .A1(n8451), .A2(n8119), .ZN(n8227) );
  INV_X1 U4967 ( .A(n7617), .ZN(n4360) );
  OR2_X1 U4968 ( .A1(n9800), .A2(n6239), .ZN(n7597) );
  OR2_X1 U4969 ( .A1(n8158), .A2(n6118), .ZN(n7567) );
  NAND2_X1 U4970 ( .A1(n7568), .A2(n7588), .ZN(n7719) );
  OR2_X1 U4971 ( .A1(n5661), .A2(n8009), .ZN(n5668) );
  AND2_X1 U4972 ( .A1(n5652), .A2(n5134), .ZN(n4450) );
  AND2_X1 U4973 ( .A1(n4454), .A2(n4453), .ZN(n8972) );
  NAND2_X1 U4974 ( .A1(n9506), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4453) );
  OR2_X1 U4975 ( .A1(n9245), .A2(n9075), .ZN(n9047) );
  NOR2_X1 U4976 ( .A1(n9046), .A2(n4538), .ZN(n4537) );
  NAND2_X1 U4977 ( .A1(n9253), .A2(n9017), .ZN(n8889) );
  NAND2_X1 U4978 ( .A1(n9191), .A2(n9009), .ZN(n4561) );
  NAND2_X1 U4979 ( .A1(n4489), .A2(n4307), .ZN(n6926) );
  NAND2_X1 U4980 ( .A1(n4490), .A2(n8819), .ZN(n4488) );
  AND2_X1 U4981 ( .A1(n8841), .A2(n8840), .ZN(n7263) );
  NAND2_X1 U4982 ( .A1(n4835), .A2(n4825), .ZN(n4447) );
  NAND2_X1 U4983 ( .A1(n4405), .A2(n4404), .ZN(n5161) );
  AOI21_X1 U4984 ( .B1(n4286), .B2(n4410), .A(n4323), .ZN(n4404) );
  NAND2_X1 U4985 ( .A1(n4413), .A2(n4952), .ZN(n4961) );
  NOR2_X1 U4986 ( .A1(n4668), .A2(n7310), .ZN(n4667) );
  INV_X1 U4987 ( .A(n4670), .ZN(n4668) );
  AND4_X1 U4988 ( .A1(n6500), .A2(n6499), .A3(n6498), .A4(n6497), .ZN(n6844)
         );
  AND2_X1 U4989 ( .A1(n7698), .A2(n7699), .ZN(n7782) );
  OR2_X1 U4990 ( .A1(n8451), .A2(n8269), .ZN(n7775) );
  NAND2_X1 U4991 ( .A1(n8266), .A2(n4726), .ZN(n4723) );
  NOR2_X1 U4992 ( .A1(n4728), .A2(n4727), .ZN(n4726) );
  INV_X1 U4993 ( .A(n8246), .ZN(n4727) );
  OR2_X1 U4994 ( .A1(n4728), .A2(n7737), .ZN(n4725) );
  OR2_X1 U4995 ( .A1(n8454), .A2(n7414), .ZN(n7774) );
  NAND2_X1 U4996 ( .A1(n8268), .A2(n8267), .ZN(n8266) );
  AOI21_X1 U4997 ( .B1(n4365), .B2(n4308), .A(n4364), .ZN(n8304) );
  INV_X1 U4998 ( .A(n4366), .ZN(n4364) );
  INV_X1 U4999 ( .A(n8357), .ZN(n4365) );
  NAND2_X1 U5000 ( .A1(n8357), .A2(n4702), .ZN(n8333) );
  NAND2_X1 U5001 ( .A1(n4780), .A2(n4312), .ZN(n7008) );
  INV_X1 U5002 ( .A(n7540), .ZN(n7339) );
  INV_X1 U5003 ( .A(n5602), .ZN(n7338) );
  NAND2_X1 U5004 ( .A1(n6657), .A2(n4309), .ZN(n6541) );
  INV_X1 U5005 ( .A(n6222), .ZN(n4774) );
  OR2_X1 U5006 ( .A1(n9716), .A2(n9800), .ZN(n6222) );
  NAND2_X1 U5007 ( .A1(n5854), .A2(n5853), .ZN(n7568) );
  NAND2_X1 U5008 ( .A1(n7976), .A2(n7978), .ZN(n7979) );
  INV_X1 U5009 ( .A(n7977), .ZN(n7978) );
  INV_X1 U5010 ( .A(n7979), .ZN(n4746) );
  NAND2_X1 U5011 ( .A1(n5458), .A2(n5587), .ZN(n5686) );
  AND2_X1 U5012 ( .A1(n9235), .A2(n9074), .ZN(n8878) );
  OR2_X1 U5013 ( .A1(n5557), .A2(n5556), .ZN(n4393) );
  OR2_X1 U5014 ( .A1(n9238), .A2(n9084), .ZN(n9048) );
  NAND2_X1 U5015 ( .A1(n9238), .A2(n9084), .ZN(n9050) );
  NAND2_X1 U5016 ( .A1(n9391), .A2(n7129), .ZN(n7092) );
  NOR2_X1 U5017 ( .A1(n9391), .A2(n7129), .ZN(n7093) );
  INV_X1 U5018 ( .A(n9591), .ZN(n9612) );
  AND2_X1 U5019 ( .A1(n6880), .A2(n6879), .ZN(n9396) );
  XNOR2_X1 U5020 ( .A(n7515), .B(n7514), .ZN(n8664) );
  NAND2_X1 U5021 ( .A1(n7152), .A2(n7151), .ZN(n7494) );
  XNOR2_X1 U5022 ( .A(n7494), .B(n7493), .ZN(n7980) );
  XNOR2_X1 U5023 ( .A(n7117), .B(n7116), .ZN(n7940) );
  NAND2_X1 U5024 ( .A1(n9324), .A2(n5954), .ZN(n7512) );
  INV_X1 U5025 ( .A(n4930), .ZN(n4931) );
  INV_X1 U5026 ( .A(n5844), .ZN(n4585) );
  INV_X1 U5027 ( .A(n4603), .ZN(n4602) );
  AOI21_X1 U5028 ( .B1(n5160), .B2(n5159), .A(n4608), .ZN(n4607) );
  INV_X1 U5029 ( .A(n4814), .ZN(n4608) );
  AOI21_X1 U5030 ( .B1(n4675), .B2(n4673), .A(n4320), .ZN(n4672) );
  INV_X1 U5031 ( .A(n4303), .ZN(n4673) );
  AOI21_X1 U5032 ( .B1(n8190), .B2(n4710), .A(n4708), .ZN(n4707) );
  INV_X1 U5033 ( .A(n7699), .ZN(n4708) );
  OR2_X1 U5034 ( .A1(n8435), .A2(n7779), .ZN(n7695) );
  INV_X1 U5035 ( .A(n4800), .ZN(n4796) );
  NOR2_X1 U5036 ( .A1(n8303), .A2(n4801), .ZN(n4800) );
  INV_X1 U5037 ( .A(n7772), .ZN(n4801) );
  OR2_X1 U5038 ( .A1(n8466), .A2(n8283), .ZN(n7668) );
  AND2_X1 U5039 ( .A1(n4552), .A2(n4553), .ZN(n4551) );
  NOR2_X1 U5040 ( .A1(n8471), .A2(n8477), .ZN(n4553) );
  INV_X1 U5041 ( .A(n4338), .ZN(n4791) );
  AND2_X1 U5042 ( .A1(n4298), .A2(n4793), .ZN(n4790) );
  NOR2_X1 U5043 ( .A1(n8335), .A2(n7645), .ZN(n4702) );
  INV_X1 U5044 ( .A(n7639), .ZN(n4375) );
  INV_X1 U5045 ( .A(n4302), .ZN(n4372) );
  NAND2_X1 U5046 ( .A1(n7175), .A2(n4802), .ZN(n7765) );
  AND2_X1 U5047 ( .A1(n7733), .A2(n7174), .ZN(n4802) );
  NOR2_X1 U5048 ( .A1(n8508), .A2(n8503), .ZN(n4546) );
  OR2_X1 U5049 ( .A1(n8508), .A2(n7077), .ZN(n7629) );
  NOR2_X1 U5050 ( .A1(n6959), .A2(n8513), .ZN(n7014) );
  OAI21_X1 U5051 ( .B1(n7724), .B2(n4700), .A(n7559), .ZN(n4698) );
  INV_X1 U5052 ( .A(n7603), .ZN(n4381) );
  INV_X1 U5053 ( .A(n7591), .ZN(n6144) );
  NOR2_X1 U5054 ( .A1(n8451), .A2(n8260), .ZN(n8251) );
  NAND2_X1 U5055 ( .A1(n8410), .A2(n7580), .ZN(n8413) );
  AND2_X1 U5056 ( .A1(n5123), .A2(n4848), .ZN(n5335) );
  INV_X1 U5057 ( .A(n8560), .ZN(n4435) );
  AOI21_X1 U5058 ( .B1(n4441), .B2(n4444), .A(n4440), .ZN(n4439) );
  INV_X1 U5059 ( .A(n8585), .ZN(n4440) );
  XNOR2_X1 U5060 ( .A(n4448), .B(n8009), .ZN(n5682) );
  INV_X1 U5061 ( .A(n4449), .ZN(n4448) );
  OAI22_X1 U5062 ( .A1(n6180), .A2(n6023), .B1(n6028), .B2(n7900), .ZN(n4449)
         );
  NAND2_X1 U5063 ( .A1(n8599), .A2(n7807), .ZN(n7816) );
  NOR2_X1 U5064 ( .A1(n9514), .A2(n8974), .ZN(n8975) );
  NOR2_X1 U5065 ( .A1(n9235), .A2(n9074), .ZN(n8879) );
  NAND2_X1 U5066 ( .A1(n9091), .A2(n4483), .ZN(n4482) );
  INV_X1 U5067 ( .A(n4484), .ZN(n4483) );
  AND2_X1 U5068 ( .A1(n9098), .A2(n9114), .ZN(n9046) );
  OR2_X1 U5069 ( .A1(n9248), .A2(n9114), .ZN(n9020) );
  OR2_X1 U5070 ( .A1(n9270), .A2(n9141), .ZN(n9037) );
  NOR2_X1 U5071 ( .A1(n9292), .A2(n9299), .ZN(n4480) );
  INV_X1 U5072 ( .A(n8798), .ZN(n4490) );
  NOR2_X1 U5073 ( .A1(n6824), .A2(n4474), .ZN(n4472) );
  OAI21_X1 U5074 ( .B1(n6601), .B2(n4566), .A(n8823), .ZN(n4565) );
  OR2_X1 U5075 ( .A1(n6876), .A2(n6982), .ZN(n8798) );
  OR2_X1 U5076 ( .A1(n6702), .A2(n6595), .ZN(n4474) );
  INV_X1 U5077 ( .A(n7262), .ZN(n4572) );
  NAND2_X1 U5078 ( .A1(n7260), .A2(n7259), .ZN(n4573) );
  OAI211_X1 U5079 ( .C1(n5364), .C2(n9330), .A(n5689), .B(n5688), .ZN(n6031)
         );
  OR2_X1 U5080 ( .A1(n8732), .A2(n5687), .ZN(n5688) );
  INV_X1 U5081 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4836) );
  OAI21_X1 U5082 ( .B1(n7515), .B2(n7500), .A(n7499), .ZN(n7535) );
  XNOR2_X1 U5083 ( .A(n5141), .B(P1_IR_REG_28__SCAN_IN), .ZN(n5144) );
  OAI21_X1 U5084 ( .B1(n7117), .B2(n7116), .A(n7115), .ZN(n7150) );
  INV_X1 U5085 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4581) );
  NAND2_X1 U5086 ( .A1(n4611), .A2(n4609), .ZN(n7058) );
  AOI21_X1 U5087 ( .B1(n4613), .B2(n4615), .A(n4610), .ZN(n4609) );
  INV_X1 U5088 ( .A(n6924), .ZN(n4610) );
  OAI21_X1 U5089 ( .B1(n6354), .B2(n6353), .A(n6352), .ZN(n6456) );
  OAI21_X1 U5090 ( .B1(n5845), .B2(n4586), .A(n4584), .ZN(n6125) );
  INV_X1 U5091 ( .A(n4587), .ZN(n4586) );
  AOI21_X1 U5092 ( .B1(n4587), .B2(n4585), .A(n4345), .ZN(n4584) );
  NOR2_X1 U5093 ( .A1(n6001), .A2(n4588), .ZN(n4587) );
  AOI21_X1 U5094 ( .B1(n4607), .B2(n4605), .A(n4604), .ZN(n4603) );
  INV_X1 U5095 ( .A(n5339), .ZN(n4604) );
  INV_X1 U5096 ( .A(n5159), .ZN(n4605) );
  INV_X1 U5097 ( .A(n4607), .ZN(n4606) );
  AOI21_X1 U5098 ( .B1(n4815), .B2(n4409), .A(n4408), .ZN(n4407) );
  INV_X1 U5099 ( .A(n5044), .ZN(n4409) );
  INV_X1 U5100 ( .A(n5059), .ZN(n4408) );
  INV_X1 U5101 ( .A(n4815), .ZN(n4410) );
  AOI21_X1 U5102 ( .B1(n4633), .B2(n4635), .A(n4632), .ZN(n4631) );
  INV_X1 U5103 ( .A(n4813), .ZN(n4632) );
  NAND2_X1 U5104 ( .A1(n4994), .A2(n4968), .ZN(n4995) );
  NAND2_X1 U5105 ( .A1(n5362), .A2(n4880), .ZN(n4882) );
  NOR2_X1 U5106 ( .A1(n4647), .A2(n4643), .ZN(n4642) );
  INV_X1 U5107 ( .A(n9726), .ZN(n4643) );
  INV_X1 U5108 ( .A(n5934), .ZN(n4647) );
  INV_X1 U5109 ( .A(n5952), .ZN(n4645) );
  INV_X1 U5110 ( .A(n8040), .ZN(n4691) );
  NAND2_X1 U5111 ( .A1(n5959), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6340) );
  OR2_X1 U5112 ( .A1(n7318), .A2(n7317), .ZN(n7352) );
  NOR2_X1 U5113 ( .A1(n9700), .A2(n4662), .ZN(n4661) );
  INV_X1 U5114 ( .A(n6473), .ZN(n4662) );
  AND2_X1 U5115 ( .A1(n5755), .A2(n5756), .ZN(n5832) );
  NOR2_X1 U5116 ( .A1(n7310), .A2(n7211), .ZN(n4666) );
  AOI21_X1 U5117 ( .B1(n7211), .B2(n7205), .A(n4288), .ZN(n4670) );
  AOI21_X1 U5118 ( .B1(n4682), .B2(n4680), .A(n4679), .ZN(n4678) );
  INV_X1 U5119 ( .A(n4682), .ZN(n4681) );
  INV_X1 U5120 ( .A(n7204), .ZN(n4679) );
  INV_X1 U5121 ( .A(n9343), .ZN(n8185) );
  NAND2_X1 U5122 ( .A1(n7507), .A2(n8200), .ZN(n7508) );
  AND2_X1 U5123 ( .A1(n4725), .A2(n7682), .ZN(n4724) );
  AND2_X1 U5124 ( .A1(n4769), .A2(n7776), .ZN(n4768) );
  NAND2_X1 U5125 ( .A1(n8240), .A2(n7506), .ZN(n7776) );
  NAND2_X1 U5126 ( .A1(n8230), .A2(n4770), .ZN(n4769) );
  INV_X1 U5127 ( .A(n7775), .ZN(n4770) );
  OR2_X1 U5128 ( .A1(n8454), .A2(n8284), .ZN(n8246) );
  INV_X1 U5129 ( .A(n4713), .ZN(n8268) );
  AOI21_X1 U5130 ( .B1(n4717), .B2(n4715), .A(n7674), .ZN(n4714) );
  INV_X1 U5131 ( .A(n4717), .ZN(n4716) );
  AND2_X1 U5132 ( .A1(n8246), .A2(n7676), .ZN(n8267) );
  OR2_X1 U5133 ( .A1(n8289), .A2(n8454), .ZN(n8260) );
  AND2_X1 U5134 ( .A1(n8279), .A2(n4283), .ZN(n4798) );
  NAND2_X1 U5135 ( .A1(n7773), .A2(n4800), .ZN(n4799) );
  NAND2_X1 U5136 ( .A1(n8304), .A2(n8303), .ZN(n8302) );
  OR2_X1 U5137 ( .A1(n8477), .A2(n8085), .ZN(n7656) );
  NAND2_X1 U5138 ( .A1(n8370), .A2(n7504), .ZN(n8357) );
  NAND2_X1 U5139 ( .A1(n8372), .A2(n8371), .ZN(n8370) );
  NOR2_X1 U5140 ( .A1(n8394), .A2(n8487), .ZN(n8365) );
  NAND2_X1 U5141 ( .A1(n7014), .A2(n4542), .ZN(n8394) );
  AND2_X1 U5142 ( .A1(n4544), .A2(n4543), .ZN(n4542) );
  INV_X1 U5143 ( .A(n8493), .ZN(n4543) );
  NAND2_X1 U5144 ( .A1(n6954), .A2(n4359), .ZN(n4357) );
  AOI21_X1 U5145 ( .B1(n4359), .B2(n4363), .A(n7623), .ZN(n4358) );
  AND4_X1 U5146 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n7046)
         );
  NAND2_X1 U5147 ( .A1(n4362), .A2(n4301), .ZN(n4361) );
  AND2_X1 U5148 ( .A1(n7617), .A2(n4301), .ZN(n7729) );
  NAND2_X1 U5149 ( .A1(n4776), .A2(n6229), .ZN(n4775) );
  AOI21_X1 U5150 ( .B1(n6140), .B2(n4778), .A(n4316), .ZN(n4777) );
  INV_X1 U5151 ( .A(n6140), .ZN(n4779) );
  INV_X1 U5152 ( .A(n5882), .ZN(n4376) );
  NAND2_X1 U5153 ( .A1(n8403), .A2(n5594), .ZN(n4764) );
  OR2_X1 U5154 ( .A1(n5593), .A2(n8405), .ZN(n5594) );
  OR2_X1 U5155 ( .A1(n6099), .A2(n9763), .ZN(n6149) );
  AND2_X1 U5156 ( .A1(n5617), .A2(n7755), .ZN(n9809) );
  INV_X1 U5157 ( .A(n4804), .ZN(n4803) );
  INV_X1 U5158 ( .A(n4654), .ZN(n4653) );
  OAI21_X1 U5159 ( .B1(n5093), .B2(n4853), .A(n5094), .ZN(n4654) );
  AND2_X1 U5160 ( .A1(n4849), .A2(n4848), .ZN(n4649) );
  INV_X1 U5161 ( .A(n4740), .ZN(n4739) );
  NOR2_X1 U5162 ( .A1(n4746), .A2(n4744), .ZN(n4743) );
  OR2_X1 U5163 ( .A1(n8549), .A2(n8016), .ZN(n7992) );
  NAND2_X1 U5164 ( .A1(n6059), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6070) );
  INV_X1 U5165 ( .A(n6061), .ZN(n6059) );
  NAND2_X1 U5166 ( .A1(n7098), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7246) );
  INV_X1 U5167 ( .A(n4425), .ZN(n4428) );
  NAND2_X1 U5168 ( .A1(n7827), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n7848) );
  INV_X1 U5169 ( .A(n7829), .ZN(n7827) );
  INV_X1 U5170 ( .A(n7891), .ZN(n7889) );
  AND2_X1 U5171 ( .A1(n7899), .A2(n7898), .ZN(n7903) );
  INV_X1 U5172 ( .A(n5668), .ZN(n4753) );
  AND2_X1 U5173 ( .A1(n8654), .A2(n4346), .ZN(n4747) );
  NAND2_X1 U5174 ( .A1(n7943), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U5175 ( .A1(n5447), .A2(n5184), .ZN(n5448) );
  AND2_X1 U5176 ( .A1(n4393), .A2(n4392), .ZN(n5447) );
  NAND2_X1 U5177 ( .A1(n5885), .A2(n5183), .ZN(n4392) );
  NOR2_X1 U5178 ( .A1(n5283), .A2(n5284), .ZN(n5547) );
  INV_X1 U5179 ( .A(n5297), .ZN(n4461) );
  NOR2_X1 U5180 ( .A1(n5547), .A2(n5546), .ZN(n5545) );
  OR2_X1 U5181 ( .A1(n9483), .A2(n9482), .ZN(n9480) );
  OR2_X1 U5182 ( .A1(n9488), .A2(n4457), .ZN(n4456) );
  NOR2_X1 U5183 ( .A1(n4459), .A2(n4458), .ZN(n4457) );
  INV_X1 U5184 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n4458) );
  NAND2_X1 U5185 ( .A1(n4456), .A2(n4455), .ZN(n4454) );
  INV_X1 U5186 ( .A(n9502), .ZN(n4455) );
  OR2_X1 U5187 ( .A1(n9521), .A2(n9522), .ZN(n4397) );
  XNOR2_X1 U5188 ( .A(n8975), .B(n4470), .ZN(n9528) );
  OR2_X1 U5189 ( .A1(n9528), .A2(n9529), .ZN(n4469) );
  NAND2_X1 U5190 ( .A1(n4397), .A2(n4396), .ZN(n4395) );
  NAND2_X1 U5191 ( .A1(n8973), .A2(n9394), .ZN(n4396) );
  XNOR2_X1 U5192 ( .A(n4465), .B(n7833), .ZN(n8985) );
  NOR2_X1 U5193 ( .A1(n9565), .A2(n4466), .ZN(n4465) );
  AND2_X1 U5194 ( .A1(n9571), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4466) );
  XNOR2_X1 U5195 ( .A(n4389), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U5196 ( .A1(n4391), .A2(n4390), .ZN(n4389) );
  NAND2_X1 U5197 ( .A1(n8966), .A2(n8967), .ZN(n4390) );
  NAND2_X1 U5198 ( .A1(n4525), .A2(n4528), .ZN(n9073) );
  AOI21_X1 U5199 ( .B1(n4533), .B2(n4530), .A(n4529), .ZN(n4528) );
  INV_X1 U5200 ( .A(n9047), .ZN(n4529) );
  NAND2_X1 U5201 ( .A1(n9048), .A2(n9050), .ZN(n9072) );
  OAI21_X1 U5202 ( .B1(n9046), .B2(n4536), .A(n9045), .ZN(n4535) );
  NAND2_X1 U5203 ( .A1(n9044), .A2(n9043), .ZN(n4536) );
  NAND2_X1 U5204 ( .A1(n9112), .A2(n4537), .ZN(n4534) );
  AOI21_X1 U5205 ( .B1(n4577), .B2(n9113), .A(n4575), .ZN(n4574) );
  INV_X1 U5206 ( .A(n9021), .ZN(n4575) );
  INV_X1 U5207 ( .A(n8889), .ZN(n9044) );
  OR2_X1 U5208 ( .A1(n9267), .A2(n9012), .ZN(n9119) );
  AND2_X1 U5209 ( .A1(n9270), .A2(n9167), .ZN(n9010) );
  NAND2_X1 U5210 ( .A1(n4561), .A2(n4559), .ZN(n4558) );
  INV_X1 U5211 ( .A(n9007), .ZN(n4559) );
  NAND2_X1 U5212 ( .A1(n4326), .A2(n4561), .ZN(n4557) );
  AND2_X1 U5213 ( .A1(n9284), .A2(n9204), .ZN(n9008) );
  NAND2_X1 U5214 ( .A1(n8892), .A2(n9035), .ZN(n9169) );
  AND2_X1 U5215 ( .A1(n7876), .A2(n7875), .ZN(n9184) );
  INV_X1 U5216 ( .A(n9031), .ZN(n4501) );
  AOI21_X1 U5217 ( .B1(n9203), .B2(n4504), .A(n4503), .ZN(n4502) );
  INV_X1 U5218 ( .A(n9030), .ZN(n4504) );
  NAND2_X1 U5219 ( .A1(n4506), .A2(n4505), .ZN(n9221) );
  AOI21_X1 U5220 ( .B1(n4507), .B2(n4513), .A(n7272), .ZN(n4506) );
  NOR2_X1 U5221 ( .A1(n7273), .A2(n9299), .ZN(n9213) );
  AOI21_X1 U5222 ( .B1(n4514), .B2(n4512), .A(n4319), .ZN(n4511) );
  INV_X1 U5223 ( .A(n8805), .ZN(n4512) );
  AND2_X1 U5224 ( .A1(n6984), .A2(n8945), .ZN(n6940) );
  NAND2_X1 U5225 ( .A1(n6617), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6628) );
  INV_X1 U5226 ( .A(n6618), .ZN(n6617) );
  AND2_X1 U5227 ( .A1(n8815), .A2(n8820), .ZN(n8896) );
  AND2_X1 U5228 ( .A1(n4524), .A2(n8701), .ZN(n4522) );
  AND4_X1 U5229 ( .A1(n6385), .A2(n6384), .A3(n6383), .A4(n6382), .ZN(n6678)
         );
  INV_X1 U5230 ( .A(n6399), .ZN(n4517) );
  NAND2_X1 U5231 ( .A1(n4495), .A2(n8692), .ZN(n6514) );
  INV_X1 U5232 ( .A(n9589), .ZN(n4495) );
  OR2_X1 U5233 ( .A1(n4494), .A2(n6039), .ZN(n4493) );
  OR2_X1 U5234 ( .A1(n6040), .A2(n5685), .ZN(n6043) );
  AND2_X1 U5235 ( .A1(n5479), .A2(n5478), .ZN(n9591) );
  AND2_X1 U5236 ( .A1(n8923), .A2(n5145), .ZN(n9357) );
  NAND2_X1 U5237 ( .A1(n7825), .A2(n7824), .ZN(n9288) );
  AND2_X1 U5238 ( .A1(n4819), .A2(n4928), .ZN(n4763) );
  XNOR2_X1 U5239 ( .A(n7535), .B(n7534), .ZN(n7533) );
  XNOR2_X1 U5240 ( .A(n5142), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5146) );
  XNOR2_X1 U5241 ( .A(n5131), .B(n5130), .ZN(n5386) );
  NAND2_X1 U5242 ( .A1(n5134), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5131) );
  NAND2_X1 U5243 ( .A1(n6716), .A2(n6715), .ZN(n7330) );
  XNOR2_X1 U5244 ( .A(n6710), .B(n6711), .ZN(n7864) );
  INV_X1 U5245 ( .A(n4447), .ZN(n4445) );
  NAND2_X1 U5246 ( .A1(n4589), .A2(n5846), .ZN(n6002) );
  NAND2_X1 U5247 ( .A1(n5845), .A2(n5844), .ZN(n4589) );
  OAI21_X1 U5248 ( .B1(n5161), .B2(n5160), .A(n5159), .ZN(n5338) );
  NAND2_X1 U5249 ( .A1(n4272), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4886) );
  INV_X1 U5250 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U5251 ( .A1(n4886), .A2(n4885), .ZN(n4905) );
  NAND2_X1 U5252 ( .A1(n5956), .A2(n5955), .ZN(n9800) );
  AND2_X1 U5253 ( .A1(n4694), .A2(n4693), .ZN(n4692) );
  NAND2_X1 U5254 ( .A1(n8145), .A2(n7451), .ZN(n4693) );
  INV_X1 U5255 ( .A(n7465), .ZN(n4694) );
  NAND2_X1 U5256 ( .A1(n7980), .A2(n5954), .ZN(n7455) );
  NAND2_X1 U5257 ( .A1(n7341), .A2(n7340), .ZN(n8483) );
  NAND2_X1 U5258 ( .A1(n6736), .A2(n6735), .ZN(n6950) );
  AND4_X1 U5259 ( .A1(n7029), .A2(n7028), .A3(n7027), .A4(n7026), .ZN(n8106)
         );
  NAND2_X1 U5260 ( .A1(n6324), .A2(n6323), .ZN(n9808) );
  NAND2_X1 U5261 ( .A1(n8144), .A2(n8145), .ZN(n4417) );
  AND2_X1 U5262 ( .A1(n5822), .A2(n5799), .ZN(n8147) );
  NOR2_X1 U5263 ( .A1(n5612), .A2(n4809), .ZN(n5613) );
  NAND2_X1 U5264 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  NAND2_X1 U5265 ( .A1(n7542), .A2(n7541), .ZN(n8427) );
  AOI21_X1 U5266 ( .B1(n8664), .B2(n5954), .A(n7516), .ZN(n7787) );
  AND2_X1 U5267 ( .A1(n7794), .A2(n7793), .ZN(n8432) );
  NAND2_X1 U5268 ( .A1(n7780), .A2(n7779), .ZN(n7781) );
  NAND2_X1 U5269 ( .A1(n8224), .A2(n8230), .ZN(n8223) );
  NAND2_X1 U5270 ( .A1(n8244), .A2(n7775), .ZN(n8224) );
  NAND2_X1 U5271 ( .A1(n4387), .A2(n8231), .ZN(n8445) );
  OR2_X1 U5272 ( .A1(n8232), .A2(n8326), .ZN(n4387) );
  NAND2_X1 U5273 ( .A1(n4723), .A2(n4725), .ZN(n8228) );
  NAND2_X1 U5274 ( .A1(n4780), .A2(n4783), .ZN(n6952) );
  CLKBUF_X1 U5275 ( .A(n6958), .Z(n8422) );
  NAND2_X1 U5276 ( .A1(n9324), .A2(n6363), .ZN(n7994) );
  NAND2_X1 U5277 ( .A1(n7940), .A2(n6363), .ZN(n7942) );
  NAND2_X1 U5278 ( .A1(n7243), .A2(n7242), .ZN(n7302) );
  AND4_X1 U5279 ( .A1(n6075), .A2(n6074), .A3(n6073), .A4(n6072), .ZN(n6588)
         );
  INV_X1 U5280 ( .A(n9157), .ZN(n9270) );
  AOI21_X1 U5281 ( .B1(n8929), .B2(n9128), .A(n6395), .ZN(n4628) );
  NAND2_X1 U5282 ( .A1(n8930), .A2(n8931), .ZN(n4629) );
  NAND2_X1 U5283 ( .A1(n8928), .A2(n9588), .ZN(n4627) );
  AOI21_X1 U5284 ( .B1(n8933), .B2(n6395), .A(n8938), .ZN(n4625) );
  INV_X1 U5285 ( .A(n9593), .ZN(n8950) );
  XNOR2_X1 U5286 ( .A(n4395), .B(n9532), .ZN(n9533) );
  OAI22_X1 U5287 ( .A1(n8985), .A2(n9564), .B1(n8984), .B2(n9576), .ZN(n4464)
         );
  INV_X1 U5288 ( .A(n8983), .ZN(n8984) );
  OAI21_X1 U5289 ( .B1(n9579), .B2(n4722), .A(n8987), .ZN(n4401) );
  AOI21_X1 U5290 ( .B1(n8743), .B2(n6363), .A(n8742), .ZN(n8993) );
  NOR2_X1 U5291 ( .A1(n8082), .A2(n7369), .ZN(n7376) );
  INV_X1 U5292 ( .A(n4674), .ZN(n4675) );
  INV_X1 U5293 ( .A(n4622), .ZN(n4621) );
  OAI21_X1 U5294 ( .B1(n7493), .B2(n4623), .A(n7509), .ZN(n4622) );
  INV_X1 U5295 ( .A(n7495), .ZN(n4623) );
  INV_X1 U5296 ( .A(n4614), .ZN(n4613) );
  OAI21_X1 U5297 ( .B1(n4616), .B2(n4615), .A(n6922), .ZN(n4614) );
  INV_X1 U5298 ( .A(n6721), .ZN(n4615) );
  INV_X1 U5299 ( .A(n5846), .ZN(n4588) );
  NAND2_X1 U5300 ( .A1(n4606), .A2(n5569), .ZN(n4600) );
  NOR2_X1 U5301 ( .A1(n4602), .A2(n5573), .ZN(n4601) );
  INV_X1 U5302 ( .A(n4591), .ZN(n4590) );
  INV_X1 U5303 ( .A(n4595), .ZN(n4593) );
  NAND2_X1 U5304 ( .A1(n4878), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4721) );
  INV_X1 U5305 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4878) );
  NOR2_X1 U5306 ( .A1(n7042), .A2(n4687), .ZN(n4686) );
  INV_X1 U5307 ( .A(n6831), .ZN(n4687) );
  INV_X1 U5308 ( .A(n8073), .ZN(n4677) );
  INV_X1 U5309 ( .A(n4686), .ZN(n4680) );
  INV_X1 U5310 ( .A(n4707), .ZN(n4705) );
  NOR2_X1 U5311 ( .A1(n7543), .A2(n7747), .ZN(n4712) );
  INV_X1 U5312 ( .A(n7695), .ZN(n4711) );
  NAND2_X1 U5313 ( .A1(n4730), .A2(n4729), .ZN(n4728) );
  INV_X1 U5314 ( .A(n8227), .ZN(n4729) );
  NAND2_X1 U5315 ( .A1(n8240), .A2(n8216), .ZN(n7681) );
  NOR2_X1 U5316 ( .A1(n8279), .A2(n4718), .ZN(n4717) );
  INV_X1 U5317 ( .A(n7668), .ZN(n4718) );
  AOI21_X1 U5318 ( .B1(n4370), .B2(n4368), .A(n4367), .ZN(n4366) );
  INV_X1 U5319 ( .A(n7665), .ZN(n4367) );
  NOR2_X1 U5320 ( .A1(n4702), .A2(n4369), .ZN(n4368) );
  INV_X1 U5321 ( .A(n7656), .ZN(n4369) );
  INV_X1 U5322 ( .A(n8318), .ZN(n4370) );
  NOR2_X1 U5323 ( .A1(n7763), .A2(n4545), .ZN(n4544) );
  INV_X1 U5324 ( .A(n4546), .ZN(n4545) );
  INV_X1 U5325 ( .A(n7625), .ZN(n7021) );
  OR2_X1 U5326 ( .A1(n6495), .A2(n6494), .ZN(n6745) );
  AND2_X1 U5327 ( .A1(n6244), .A2(n4539), .ZN(n6737) );
  AND2_X1 U5328 ( .A1(n9821), .A2(n4299), .ZN(n4539) );
  NOR2_X1 U5329 ( .A1(n6529), .A2(n9808), .ZN(n4541) );
  NAND2_X1 U5330 ( .A1(n4382), .A2(n4266), .ZN(n6523) );
  INV_X1 U5331 ( .A(n6232), .ZN(n4382) );
  AND2_X1 U5332 ( .A1(n5912), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5935) );
  INV_X1 U5333 ( .A(n5855), .ZN(n4778) );
  NOR2_X1 U5334 ( .A1(n6443), .A2(n5853), .ZN(n5860) );
  NAND2_X1 U5335 ( .A1(n8413), .A2(n8404), .ZN(n8403) );
  INV_X1 U5336 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4875) );
  INV_X1 U5337 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4805) );
  NOR2_X1 U5338 ( .A1(n4531), .A2(n4527), .ZN(n4526) );
  INV_X1 U5339 ( .A(n4533), .ZN(n4531) );
  INV_X1 U5340 ( .A(n4537), .ZN(n4530) );
  NOR2_X1 U5341 ( .A1(n4578), .A2(n9019), .ZN(n4577) );
  INV_X1 U5342 ( .A(n9020), .ZN(n4578) );
  NAND2_X1 U5343 ( .A1(n9098), .A2(n4485), .ZN(n4484) );
  OR2_X1 U5344 ( .A1(n9261), .A2(n9140), .ZN(n8890) );
  NAND2_X1 U5345 ( .A1(n4480), .A2(n9200), .ZN(n4479) );
  AND2_X1 U5346 ( .A1(n4511), .A2(n4508), .ZN(n4507) );
  NAND2_X1 U5347 ( .A1(n6360), .A2(n6359), .ZN(n4562) );
  INV_X1 U5348 ( .A(n8809), .ZN(n4494) );
  NAND2_X1 U5349 ( .A1(n6045), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6061) );
  AND2_X1 U5350 ( .A1(n6395), .A2(n9128), .ZN(n5466) );
  NAND2_X1 U5351 ( .A1(n8793), .A2(n8675), .ZN(n4518) );
  INV_X1 U5352 ( .A(n4520), .ZN(n4519) );
  OAI21_X1 U5353 ( .B1(n4522), .B2(n4521), .A(n8815), .ZN(n4520) );
  NAND2_X1 U5354 ( .A1(n8886), .A2(n9588), .ZN(n8877) );
  INV_X1 U5355 ( .A(n5133), .ZN(n5132) );
  NAND2_X1 U5356 ( .A1(n6128), .A2(n6127), .ZN(n6354) );
  NAND2_X1 U5357 ( .A1(n6125), .A2(n6124), .ZN(n6128) );
  AND2_X1 U5358 ( .A1(n5846), .A2(n5637), .ZN(n5844) );
  NAND2_X1 U5359 ( .A1(n5000), .A2(n4999), .ZN(n5044) );
  INV_X1 U5360 ( .A(n4994), .ZN(n4634) );
  INV_X1 U5361 ( .A(n4636), .ZN(n4635) );
  NOR2_X1 U5362 ( .A1(n7045), .A2(n4683), .ZN(n4682) );
  INV_X1 U5363 ( .A(n4685), .ZN(n4683) );
  NAND2_X1 U5364 ( .A1(n7040), .A2(n7041), .ZN(n4685) );
  NAND2_X1 U5365 ( .A1(n6832), .A2(n4686), .ZN(n4684) );
  INV_X1 U5366 ( .A(n4659), .ZN(n4658) );
  OAI21_X1 U5367 ( .B1(n4660), .B2(n4661), .A(n6792), .ZN(n4659) );
  NAND2_X1 U5368 ( .A1(n4658), .A2(n4660), .ZN(n4656) );
  OR2_X1 U5369 ( .A1(n7407), .A2(n8065), .ZN(n7409) );
  OR2_X1 U5370 ( .A1(n7359), .A2(n9905), .ZN(n7382) );
  INV_X1 U5371 ( .A(n7187), .ZN(n7186) );
  NOR2_X1 U5372 ( .A1(n7713), .A2(n7712), .ZN(n7745) );
  AND2_X1 U5373 ( .A1(n7711), .A2(n7710), .ZN(n7712) );
  INV_X1 U5374 ( .A(n4703), .ZN(n7531) );
  OAI21_X1 U5375 ( .B1(n8198), .B2(n4706), .A(n4704), .ZN(n4703) );
  NAND2_X1 U5376 ( .A1(n7706), .A2(n4710), .ZN(n4706) );
  AOI21_X1 U5377 ( .B1(n4705), .B2(n7706), .A(n4712), .ZN(n4704) );
  AND4_X1 U5378 ( .A1(n6843), .A2(n6842), .A3(n6841), .A4(n6840), .ZN(n7077)
         );
  NAND2_X1 U5379 ( .A1(n5775), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U5380 ( .A1(n8196), .A2(n7695), .ZN(n7789) );
  NOR3_X1 U5381 ( .A1(n8233), .A2(n8435), .A3(n8440), .ZN(n8193) );
  AOI21_X1 U5382 ( .B1(n8266), .B2(n8246), .A(n8247), .ZN(n8226) );
  OAI21_X1 U5383 ( .B1(n7773), .B2(n4797), .A(n4795), .ZN(n8259) );
  INV_X1 U5384 ( .A(n4798), .ZN(n4797) );
  AOI21_X1 U5385 ( .B1(n4798), .B2(n4796), .A(n4317), .ZN(n4795) );
  NOR2_X1 U5386 ( .A1(n8293), .A2(n4550), .ZN(n4549) );
  INV_X1 U5387 ( .A(n4551), .ZN(n4550) );
  AND2_X1 U5388 ( .A1(n8302), .A2(n4717), .ZN(n8282) );
  NAND2_X1 U5389 ( .A1(n8349), .A2(n4553), .ZN(n8313) );
  NAND2_X1 U5390 ( .A1(n4347), .A2(n4298), .ZN(n4789) );
  NAND2_X1 U5391 ( .A1(n8349), .A2(n8344), .ZN(n8338) );
  AND2_X1 U5392 ( .A1(n8353), .A2(n8365), .ZN(n8349) );
  INV_X1 U5393 ( .A(n4374), .ZN(n4373) );
  AOI21_X1 U5394 ( .B1(n4372), .B2(n4374), .A(n7641), .ZN(n4371) );
  NOR2_X1 U5395 ( .A1(n7766), .A2(n4375), .ZN(n4374) );
  NAND2_X1 U5396 ( .A1(n7014), .A2(n4544), .ZN(n8393) );
  OR2_X1 U5397 ( .A1(n7079), .A2(n7078), .ZN(n7187) );
  NAND2_X1 U5398 ( .A1(n7182), .A2(n7553), .ZN(n7184) );
  NAND2_X1 U5399 ( .A1(n7175), .A2(n7174), .ZN(n7179) );
  AND2_X1 U5400 ( .A1(n7553), .A2(n7552), .ZN(n7632) );
  INV_X1 U5401 ( .A(n7632), .ZN(n7732) );
  NAND2_X1 U5402 ( .A1(n7014), .A2(n7013), .ZN(n7072) );
  INV_X1 U5403 ( .A(n4784), .ZN(n4783) );
  OAI22_X1 U5404 ( .A1(n7729), .A2(n4785), .B1(n8152), .B2(n6950), .ZN(n4784)
         );
  NAND2_X1 U5405 ( .A1(n4786), .A2(n6732), .ZN(n4785) );
  INV_X1 U5406 ( .A(n7727), .ZN(n4786) );
  NAND2_X1 U5407 ( .A1(n4781), .A2(n4310), .ZN(n4780) );
  INV_X1 U5408 ( .A(n7729), .ZN(n4787) );
  NAND2_X1 U5409 ( .A1(n6233), .A2(n4380), .ZN(n4378) );
  NAND2_X1 U5410 ( .A1(n6660), .A2(n7605), .ZN(n6537) );
  AND4_X1 U5411 ( .A1(n6491), .A2(n6490), .A3(n6489), .A4(n6488), .ZN(n9702)
         );
  OAI21_X1 U5412 ( .B1(n4776), .B2(n4772), .A(n4771), .ZN(n6659) );
  AOI21_X1 U5413 ( .B1(n4773), .B2(n7722), .A(n4287), .ZN(n4771) );
  INV_X1 U5414 ( .A(n4773), .ZN(n4772) );
  NAND2_X1 U5415 ( .A1(n6244), .A2(n4541), .ZN(n6667) );
  AND2_X1 U5416 ( .A1(n7560), .A2(n7605), .ZN(n7724) );
  NAND2_X1 U5417 ( .A1(n6523), .A2(n7603), .ZN(n6661) );
  NAND2_X1 U5418 ( .A1(n6661), .A2(n7724), .ZN(n6660) );
  AND4_X1 U5419 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(n9713)
         );
  NAND2_X1 U5420 ( .A1(n6244), .A2(n9719), .ZN(n6669) );
  NAND2_X1 U5421 ( .A1(n4355), .A2(n9790), .ZN(n6215) );
  NOR2_X1 U5422 ( .A1(n6215), .A2(n9793), .ZN(n6162) );
  NAND2_X1 U5423 ( .A1(n4695), .A2(n7569), .ZN(n6145) );
  NOR2_X1 U5424 ( .A1(n6144), .A2(n4697), .ZN(n4696) );
  INV_X1 U5425 ( .A(n7589), .ZN(n4697) );
  AND4_X1 U5426 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(n6239)
         );
  NAND2_X1 U5427 ( .A1(n7569), .A2(n7591), .ZN(n7718) );
  NAND2_X1 U5428 ( .A1(n4764), .A2(n7715), .ZN(n5852) );
  AND2_X1 U5429 ( .A1(n7572), .A2(n8410), .ZN(n5607) );
  NAND2_X1 U5430 ( .A1(n5607), .A2(n5608), .ZN(n5857) );
  AND3_X1 U5431 ( .A1(n5762), .A2(n5761), .A3(n5760), .ZN(n9780) );
  OR2_X1 U5432 ( .A1(n5602), .A2(n5589), .ZN(n5590) );
  INV_X1 U5433 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5010) );
  INV_X1 U5434 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4648) );
  AND2_X1 U5435 ( .A1(n4842), .A2(n4903), .ZN(n4765) );
  OR2_X1 U5436 ( .A1(n6380), .A2(n6693), .ZN(n6608) );
  INV_X1 U5437 ( .A(n5682), .ZN(n5679) );
  AND2_X1 U5438 ( .A1(n7840), .A2(n7841), .ZN(n8569) );
  AND2_X1 U5439 ( .A1(n4442), .A2(n7863), .ZN(n4441) );
  NAND2_X1 U5440 ( .A1(n8619), .A2(n4443), .ZN(n4442) );
  INV_X1 U5441 ( .A(n8619), .ZN(n4444) );
  OR2_X1 U5442 ( .A1(n7928), .A2(n7927), .ZN(n7944) );
  INV_X1 U5443 ( .A(n8611), .ZN(n4431) );
  NAND2_X1 U5444 ( .A1(n4420), .A2(n4436), .ZN(n4425) );
  INV_X1 U5445 ( .A(n8631), .ZN(n4420) );
  NAND2_X1 U5446 ( .A1(n4427), .A2(n4297), .ZN(n4426) );
  NOR2_X1 U5447 ( .A1(n8602), .A2(n4755), .ZN(n4754) );
  INV_X1 U5448 ( .A(n4757), .ZN(n4755) );
  NAND2_X1 U5449 ( .A1(n7799), .A2(n7798), .ZN(n4757) );
  NAND2_X1 U5450 ( .A1(n7800), .A2(n4758), .ZN(n4756) );
  OR2_X1 U5451 ( .A1(n7799), .A2(n7798), .ZN(n4758) );
  INV_X1 U5452 ( .A(n6070), .ZN(n6069) );
  OR2_X1 U5453 ( .A1(n7848), .A2(n8621), .ZN(n7869) );
  NAND2_X1 U5454 ( .A1(n6557), .A2(n6689), .ZN(n4733) );
  NAND2_X1 U5455 ( .A1(n7277), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U5456 ( .A1(n7816), .A2(n7817), .ZN(n8639) );
  INV_X1 U5457 ( .A(n6176), .ZN(n4741) );
  INV_X1 U5458 ( .A(n6885), .ZN(n6884) );
  OR2_X1 U5459 ( .A1(n9229), .A2(n8991), .ZN(n8924) );
  INV_X1 U5460 ( .A(n7983), .ZN(n8024) );
  NOR2_X1 U5461 ( .A1(n9439), .A2(n4398), .ZN(n9438) );
  NAND2_X1 U5462 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n4398) );
  NAND2_X1 U5463 ( .A1(n5448), .A2(n5185), .ZN(n5189) );
  NAND2_X1 U5464 ( .A1(n4460), .A2(n4318), .ZN(n9449) );
  NOR2_X1 U5465 ( .A1(n9476), .A2(n9475), .ZN(n9474) );
  NOR2_X1 U5466 ( .A1(n9474), .A2(n4452), .ZN(n5304) );
  AND2_X1 U5467 ( .A1(n9479), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U5468 ( .A1(n5304), .A2(n5303), .ZN(n8969) );
  NAND2_X1 U5469 ( .A1(n8969), .A2(n4451), .ZN(n9490) );
  OR2_X1 U5470 ( .A1(n8970), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4451) );
  XNOR2_X1 U5471 ( .A(n8972), .B(n8973), .ZN(n9516) );
  AND2_X1 U5472 ( .A1(n4469), .A2(n4468), .ZN(n9540) );
  NAND2_X1 U5473 ( .A1(n8976), .A2(n9532), .ZN(n4468) );
  OR2_X1 U5474 ( .A1(n9573), .A2(n9574), .ZN(n4391) );
  NOR2_X1 U5475 ( .A1(n8879), .A2(n8878), .ZN(n9025) );
  NOR2_X1 U5476 ( .A1(n9125), .A2(n4484), .ZN(n9094) );
  NOR2_X1 U5477 ( .A1(n9018), .A2(n9253), .ZN(n9019) );
  NOR2_X1 U5478 ( .A1(n9125), .A2(n9253), .ZN(n9108) );
  NAND2_X1 U5479 ( .A1(n9261), .A2(n9015), .ZN(n9016) );
  AND2_X1 U5480 ( .A1(n9043), .A2(n8889), .ZN(n9113) );
  NOR2_X1 U5481 ( .A1(n4273), .A2(n9113), .ZN(n9106) );
  NAND2_X1 U5482 ( .A1(n8890), .A2(n9042), .ZN(n9130) );
  OR2_X1 U5483 ( .A1(n9137), .A2(n9138), .ZN(n9120) );
  AND2_X1 U5484 ( .A1(n7897), .A2(n7896), .ZN(n9141) );
  AOI21_X1 U5485 ( .B1(n4284), .B2(n4499), .A(n4498), .ZN(n4497) );
  INV_X1 U5486 ( .A(n9203), .ZN(n4499) );
  NOR2_X1 U5487 ( .A1(n7273), .A2(n4478), .ZN(n9214) );
  INV_X1 U5488 ( .A(n4480), .ZN(n4478) );
  INV_X1 U5489 ( .A(n4570), .ZN(n4568) );
  AOI21_X1 U5490 ( .B1(n4571), .B2(n7258), .A(n4291), .ZN(n4570) );
  OAI21_X1 U5491 ( .B1(n6881), .B2(n4490), .A(n8819), .ZN(n6882) );
  NAND2_X1 U5492 ( .A1(n6606), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6618) );
  INV_X1 U5493 ( .A(n6608), .ZN(n6606) );
  NAND2_X1 U5494 ( .A1(n4473), .A2(n4472), .ZN(n9352) );
  NAND2_X1 U5495 ( .A1(n4473), .A2(n4289), .ZN(n6895) );
  INV_X1 U5496 ( .A(n4565), .ZN(n4564) );
  NOR2_X1 U5497 ( .A1(n6406), .A2(n4474), .ZN(n9350) );
  CLKBUF_X1 U5498 ( .A(n6650), .Z(n6651) );
  NOR2_X1 U5499 ( .A1(n6406), .A2(n6595), .ZN(n6646) );
  NOR2_X1 U5500 ( .A1(n4447), .A2(n4322), .ZN(n4446) );
  AND4_X1 U5501 ( .A1(n5695), .A2(n5694), .A3(n5693), .A4(n5692), .ZN(n6414)
         );
  NAND2_X1 U5502 ( .A1(n8734), .A2(n8733), .ZN(n9373) );
  NAND2_X1 U5503 ( .A1(n8666), .A2(n8665), .ZN(n9235) );
  NAND2_X1 U5504 ( .A1(n7962), .A2(n7961), .ZN(n9248) );
  NAND2_X1 U5505 ( .A1(n7959), .A2(n6363), .ZN(n7962) );
  NAND2_X1 U5506 ( .A1(n7847), .A2(n7846), .ZN(n9284) );
  NAND2_X1 U5507 ( .A1(n4573), .A2(n7262), .ZN(n7264) );
  AND3_X1 U5508 ( .A1(n6058), .A2(n6057), .A3(n6056), .ZN(n9668) );
  NAND2_X1 U5509 ( .A1(n9615), .A2(n9638), .ZN(n9684) );
  INV_X1 U5510 ( .A(n9632), .ZN(n9678) );
  AND2_X1 U5511 ( .A1(n5536), .A2(n5981), .ZN(n9632) );
  NOR2_X1 U5512 ( .A1(n4812), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4762) );
  INV_X1 U5513 ( .A(SI_30_), .ZN(n4583) );
  CLKBUF_X1 U5514 ( .A(n5144), .Z(n5145) );
  XNOR2_X1 U5515 ( .A(n7150), .B(n7149), .ZN(n7959) );
  NOR2_X1 U5516 ( .A1(n4580), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4579) );
  NOR2_X1 U5517 ( .A1(n7329), .A2(n4617), .ZN(n4616) );
  INV_X1 U5518 ( .A(n6715), .ZN(n4617) );
  OAI21_X1 U5519 ( .B1(n5161), .B2(n4606), .A(n4603), .ZN(n5574) );
  NAND2_X1 U5520 ( .A1(n4406), .A2(n4407), .ZN(n5070) );
  OR2_X1 U5521 ( .A1(n5045), .A2(n4410), .ZN(n4406) );
  NAND2_X1 U5522 ( .A1(n4638), .A2(n4963), .ZN(n4996) );
  NAND2_X1 U5523 ( .A1(n4961), .A2(n4960), .ZN(n4638) );
  XNOR2_X1 U5524 ( .A(n4961), .B(n4959), .ZN(n6053) );
  NAND2_X1 U5525 ( .A1(n4594), .A2(n4927), .ZN(n4932) );
  INV_X1 U5526 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4928) );
  AND2_X1 U5527 ( .A1(n4913), .A2(n4819), .ZN(n4917) );
  NAND2_X1 U5528 ( .A1(n4888), .A2(n4887), .ZN(n4388) );
  XNOR2_X1 U5529 ( .A(n4899), .B(SI_2_), .ZN(n4897) );
  AOI21_X1 U5530 ( .B1(n5934), .B2(n4646), .A(n4645), .ZN(n4644) );
  INV_X1 U5531 ( .A(n5932), .ZN(n4646) );
  NAND2_X1 U5532 ( .A1(n8144), .A2(n7451), .ZN(n4689) );
  XNOR2_X1 U5533 ( .A(n7417), .B(n4816), .ZN(n8063) );
  NOR2_X1 U5534 ( .A1(n4691), .A2(n7452), .ZN(n4690) );
  NAND2_X1 U5535 ( .A1(n4305), .A2(n5749), .ZN(n5820) );
  NAND2_X1 U5536 ( .A1(n4403), .A2(n7358), .ZN(n8471) );
  AND4_X1 U5537 ( .A1(n7192), .A2(n7191), .A3(n7190), .A4(n7189), .ZN(n8105)
         );
  NAND2_X1 U5538 ( .A1(n7207), .A2(n7206), .ZN(n4669) );
  OAI21_X1 U5539 ( .B1(n7207), .B2(n4671), .A(n4670), .ZN(n7311) );
  NAND2_X1 U5540 ( .A1(n7217), .A2(n7216), .ZN(n8493) );
  NAND2_X1 U5541 ( .A1(n7399), .A2(n7398), .ZN(n8454) );
  INV_X1 U5542 ( .A(n5110), .ZN(n5109) );
  NAND2_X1 U5543 ( .A1(n6832), .A2(n6831), .ZN(n7043) );
  NAND2_X1 U5544 ( .A1(n6835), .A2(n6834), .ZN(n8513) );
  AOI21_X1 U5545 ( .B1(n6474), .B2(n4661), .A(n4660), .ZN(n4657) );
  AOI21_X1 U5546 ( .B1(n4666), .B2(n4670), .A(n4665), .ZN(n4664) );
  NOR2_X1 U5547 ( .A1(n7309), .A2(n7308), .ZN(n4665) );
  NAND2_X1 U5548 ( .A1(n7314), .A2(n7313), .ZN(n8487) );
  NAND2_X1 U5549 ( .A1(n9724), .A2(n5932), .ZN(n5933) );
  NAND2_X1 U5550 ( .A1(n5933), .A2(n5934), .ZN(n5953) );
  NAND2_X1 U5551 ( .A1(n7069), .A2(n7068), .ZN(n8503) );
  NAND2_X1 U5552 ( .A1(n5775), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U5553 ( .A1(n5609), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U5554 ( .A1(n5775), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5112) );
  AND2_X1 U5555 ( .A1(n7502), .A2(n7501), .ZN(n9343) );
  AND2_X1 U5556 ( .A1(n8202), .A2(n8201), .ZN(n8438) );
  AND2_X1 U5557 ( .A1(n8219), .A2(n8218), .ZN(n8443) );
  AND2_X1 U5558 ( .A1(n4724), .A2(n4723), .ZN(n8215) );
  OAI21_X1 U5559 ( .B1(n8244), .B2(n4730), .A(n4768), .ZN(n8208) );
  NAND2_X1 U5560 ( .A1(n7425), .A2(n7424), .ZN(n8451) );
  NAND2_X1 U5561 ( .A1(n7940), .A2(n5954), .ZN(n7425) );
  AND2_X1 U5562 ( .A1(n8271), .A2(n8270), .ZN(n8457) );
  NAND2_X1 U5563 ( .A1(n4799), .A2(n4798), .ZN(n8278) );
  NAND2_X1 U5564 ( .A1(n4799), .A2(n4283), .ZN(n8276) );
  AND2_X1 U5565 ( .A1(n8308), .A2(n8307), .ZN(n8469) );
  NAND2_X1 U5566 ( .A1(n8333), .A2(n7656), .ZN(n8317) );
  NAND2_X1 U5567 ( .A1(n8357), .A2(n7654), .ZN(n8327) );
  NAND2_X1 U5568 ( .A1(n8385), .A2(n4793), .ZN(n4792) );
  NAND2_X1 U5569 ( .A1(n7503), .A2(n7639), .ZN(n8380) );
  NAND2_X1 U5570 ( .A1(n4357), .A2(n4358), .ZN(n7020) );
  NAND2_X1 U5571 ( .A1(n4361), .A2(n7617), .ZN(n7019) );
  NAND2_X1 U5572 ( .A1(n4782), .A2(n6732), .ZN(n6951) );
  NAND2_X1 U5573 ( .A1(n6730), .A2(n7727), .ZN(n4782) );
  NAND2_X1 U5574 ( .A1(n6657), .A2(n6533), .ZN(n6539) );
  NAND2_X1 U5575 ( .A1(n4775), .A2(n4773), .ZN(n6530) );
  NAND2_X1 U5576 ( .A1(n4775), .A2(n6222), .ZN(n6227) );
  OR2_X1 U5577 ( .A1(n9763), .A2(n6100), .ZN(n8389) );
  NAND2_X1 U5578 ( .A1(n5856), .A2(n6140), .ZN(n6136) );
  NAND2_X1 U5579 ( .A1(n6440), .A2(n5855), .ZN(n5856) );
  NAND2_X1 U5580 ( .A1(n4376), .A2(n5954), .ZN(n5774) );
  INV_X1 U5581 ( .A(n9780), .ZN(n5853) );
  OR2_X1 U5582 ( .A1(n5585), .A2(n6098), .ZN(n9833) );
  OAI21_X1 U5583 ( .B1(n8448), .B2(n9804), .A(n4315), .ZN(n4385) );
  AND2_X1 U5584 ( .A1(n8447), .A2(n9809), .ZN(n4386) );
  NAND2_X1 U5585 ( .A1(n4651), .A2(n4650), .ZN(n5096) );
  AOI21_X1 U5586 ( .B1(n4653), .B2(n4853), .A(n4853), .ZN(n4650) );
  NAND2_X1 U5587 ( .A1(n8653), .A2(n7979), .ZN(n8551) );
  AND4_X1 U5588 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n7144)
         );
  OR2_X1 U5589 ( .A1(n4437), .A2(n4436), .ZN(n8558) );
  NOR2_X1 U5590 ( .A1(n8629), .A2(n8631), .ZN(n4437) );
  NAND2_X1 U5591 ( .A1(n7909), .A2(n7908), .ZN(n9267) );
  OAI21_X1 U5592 ( .B1(n6557), .B2(n6690), .A(n6689), .ZN(n6819) );
  NAND2_X1 U5593 ( .A1(n4742), .A2(n4313), .ZN(n8037) );
  OR2_X1 U5594 ( .A1(n4747), .A2(n4746), .ZN(n4745) );
  AND2_X1 U5595 ( .A1(n7484), .A2(n5669), .ZN(n8577) );
  OAI21_X1 U5596 ( .B1(n8571), .B2(n4444), .A(n4441), .ZN(n8584) );
  NAND2_X1 U5597 ( .A1(n7867), .A2(n7866), .ZN(n9277) );
  NAND2_X1 U5598 ( .A1(n7291), .A2(n7290), .ZN(n7800) );
  NAND2_X1 U5599 ( .A1(n4756), .A2(n4757), .ZN(n8601) );
  NAND2_X1 U5600 ( .A1(n7271), .A2(n7270), .ZN(n9299) );
  NAND2_X1 U5601 ( .A1(n8618), .A2(n8619), .ZN(n8617) );
  NAND2_X1 U5602 ( .A1(n8571), .A2(n8567), .ZN(n8618) );
  AND4_X1 U5603 ( .A1(n6623), .A2(n6622), .A3(n6621), .A4(n6620), .ZN(n6982)
         );
  INV_X1 U5604 ( .A(n9396), .ZN(n6984) );
  NAND2_X1 U5605 ( .A1(n4733), .A2(n4734), .ZN(n6821) );
  INV_X1 U5606 ( .A(n8657), .ZN(n8644) );
  AND2_X1 U5607 ( .A1(n7997), .A2(n7964), .ZN(n9096) );
  NAND2_X1 U5608 ( .A1(n7983), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U5609 ( .A1(n5472), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4760) );
  INV_X1 U5610 ( .A(n4393), .ZN(n5555) );
  NAND2_X1 U5611 ( .A1(n4462), .A2(n5297), .ZN(n5542) );
  NAND2_X1 U5612 ( .A1(n5296), .A2(n5295), .ZN(n4462) );
  NOR2_X1 U5613 ( .A1(n5545), .A2(n5285), .ZN(n9458) );
  NAND2_X1 U5614 ( .A1(n9458), .A2(n9457), .ZN(n9456) );
  AND2_X1 U5615 ( .A1(n9480), .A2(n5290), .ZN(n5292) );
  INV_X1 U5616 ( .A(n4456), .ZN(n9503) );
  INV_X1 U5617 ( .A(n4454), .ZN(n9501) );
  INV_X1 U5618 ( .A(n4397), .ZN(n9520) );
  INV_X1 U5619 ( .A(n4469), .ZN(n9527) );
  AOI21_X1 U5620 ( .B1(n9533), .B2(P1_REG1_REG_15__SCAN_IN), .A(n4394), .ZN(
        n8962) );
  NOR2_X1 U5621 ( .A1(n4395), .A2(n4470), .ZN(n4394) );
  INV_X1 U5622 ( .A(n4391), .ZN(n9572) );
  INV_X1 U5623 ( .A(n9373), .ZN(n8996) );
  AND2_X1 U5624 ( .A1(n4300), .A2(n9067), .ZN(n9239) );
  AOI21_X1 U5625 ( .B1(n9077), .B2(n9612), .A(n9076), .ZN(n9241) );
  INV_X1 U5626 ( .A(n9245), .ZN(n9091) );
  INV_X1 U5627 ( .A(n4535), .ZN(n4532) );
  OAI21_X1 U5628 ( .B1(n9112), .B2(n9044), .A(n9043), .ZN(n9099) );
  INV_X1 U5629 ( .A(n9248), .ZN(n9098) );
  INV_X1 U5630 ( .A(n9267), .ZN(n9149) );
  AND2_X1 U5631 ( .A1(n7888), .A2(n7887), .ZN(n9157) );
  NAND2_X1 U5632 ( .A1(n4557), .A2(n4558), .ZN(n4555) );
  NAND2_X1 U5633 ( .A1(n4554), .A2(n4557), .ZN(n9170) );
  OR2_X1 U5634 ( .A1(n9194), .A2(n4558), .ZN(n4554) );
  NAND2_X1 U5635 ( .A1(n4500), .A2(n4502), .ZN(n9181) );
  NAND2_X1 U5636 ( .A1(n4501), .A2(n9203), .ZN(n4500) );
  NAND2_X1 U5637 ( .A1(n4560), .A2(n9006), .ZN(n9180) );
  OR2_X1 U5638 ( .A1(n9194), .A2(n9007), .ZN(n4560) );
  NAND2_X1 U5639 ( .A1(n9202), .A2(n9203), .ZN(n9201) );
  NAND2_X1 U5640 ( .A1(n9031), .A2(n9030), .ZN(n9202) );
  NAND2_X1 U5641 ( .A1(n4510), .A2(n4514), .ZN(n4509) );
  NAND2_X1 U5642 ( .A1(n6652), .A2(n6602), .ZN(n9349) );
  NAND2_X1 U5643 ( .A1(n4523), .A2(n4522), .ZN(n6643) );
  NAND2_X1 U5644 ( .A1(n4523), .A2(n8701), .ZN(n6625) );
  NAND2_X1 U5645 ( .A1(n6514), .A2(n8697), .ZN(n6067) );
  INV_X1 U5646 ( .A(n9619), .ZN(n9132) );
  OR2_X1 U5647 ( .A1(n5625), .A2(n5977), .ZN(n9697) );
  OAI21_X1 U5648 ( .B1(n7533), .B2(n4583), .A(n7536), .ZN(n4582) );
  NAND2_X1 U5649 ( .A1(n4620), .A2(n7495), .ZN(n7510) );
  XNOR2_X1 U5650 ( .A(n6923), .B(n6922), .ZN(n7906) );
  NAND2_X1 U5651 ( .A1(n4612), .A2(n6721), .ZN(n6923) );
  NAND2_X1 U5652 ( .A1(n6716), .A2(n4616), .ZN(n4612) );
  CLKBUF_X1 U5653 ( .A(n5386), .Z(n8886) );
  NAND2_X1 U5654 ( .A1(n5340), .A2(n4835), .ZN(n5638) );
  NOR2_X1 U5655 ( .A1(n5076), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5167) );
  XNOR2_X1 U5656 ( .A(n4924), .B(n4923), .ZN(n5882) );
  INV_X1 U5657 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10001) );
  INV_X1 U5658 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5687) );
  XNOR2_X1 U5659 ( .A(n4471), .B(n4906), .ZN(n9330) );
  NAND2_X1 U5660 ( .A1(n4905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4471) );
  INV_X1 U5661 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5672) );
  OAI21_X1 U5662 ( .B1(n4886), .B2(n4885), .A(n4905), .ZN(n5675) );
  XNOR2_X1 U5663 ( .A(n4399), .B(n4907), .ZN(n9430) );
  NAND2_X1 U5664 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4399) );
  OAI21_X1 U5665 ( .B1(n8143), .B2(n4416), .A(n4415), .ZN(P2_U3242) );
  AOI21_X1 U5666 ( .B1(n8447), .B2(n8147), .A(n8146), .ZN(n4415) );
  NAND2_X1 U5667 ( .A1(n4417), .A2(n9733), .ZN(n4416) );
  AOI211_X1 U5668 ( .C1(n8431), .C2(n8409), .A(n7796), .B(n7795), .ZN(n7797)
         );
  NAND2_X1 U5669 ( .A1(n4384), .A2(n4383), .ZN(P2_U3514) );
  NAND2_X1 U5670 ( .A1(n9825), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n4383) );
  NAND2_X1 U5671 ( .A1(n8523), .A2(n4267), .ZN(n4384) );
  NAND2_X1 U5672 ( .A1(n4624), .A2(n8937), .ZN(P1_U3240) );
  NAND2_X1 U5673 ( .A1(n4626), .A2(n4625), .ZN(n4624) );
  INV_X1 U5674 ( .A(n4401), .ZN(n4400) );
  NAND2_X1 U5675 ( .A1(n4464), .A2(n9128), .ZN(n4402) );
  NAND2_X1 U5676 ( .A1(n8986), .A2(n9588), .ZN(n4467) );
  AND4_X1 U5677 ( .A1(n4822), .A2(n4821), .A3(n4938), .A4(n4820), .ZN(n4282)
         );
  INV_X2 U5678 ( .A(n5907), .ZN(n5954) );
  OR2_X1 U5679 ( .A1(n8466), .A2(n8319), .ZN(n4283) );
  AND2_X1 U5680 ( .A1(n4502), .A2(n8893), .ZN(n4284) );
  AND4_X2 U5681 ( .A1(n4306), .A2(n4828), .A3(n4827), .A4(n4826), .ZN(n4285)
         );
  AND2_X1 U5682 ( .A1(n4407), .A2(n5067), .ZN(n4286) );
  NAND2_X1 U5683 ( .A1(n6616), .A2(n6615), .ZN(n6876) );
  INV_X1 U5684 ( .A(n6876), .ZN(n4475) );
  NAND2_X1 U5685 ( .A1(n7681), .A2(n7682), .ZN(n8230) );
  INV_X1 U5686 ( .A(n8230), .ZN(n4730) );
  AND2_X1 U5687 ( .A1(n6529), .A2(n8155), .ZN(n4287) );
  AND2_X1 U5688 ( .A1(n7668), .A2(n7667), .ZN(n8303) );
  INV_X1 U5689 ( .A(n8303), .ZN(n4715) );
  AND2_X1 U5690 ( .A1(n7214), .A2(n7213), .ZN(n4288) );
  AND2_X1 U5691 ( .A1(n4475), .A2(n4472), .ZN(n4289) );
  AND2_X1 U5692 ( .A1(n6367), .A2(n6362), .ZN(n4290) );
  INV_X1 U5693 ( .A(n4301), .ZN(n4363) );
  AND2_X1 U5694 ( .A1(n7302), .A2(n8942), .ZN(n4291) );
  NOR2_X1 U5695 ( .A1(n5543), .A2(n4461), .ZN(n4292) );
  AND3_X1 U5696 ( .A1(n4823), .A2(n4336), .A3(n4282), .ZN(n4293) );
  AND2_X1 U5697 ( .A1(n4649), .A2(n4648), .ZN(n4294) );
  AND2_X1 U5698 ( .A1(n4656), .A2(n6797), .ZN(n4295) );
  NAND2_X1 U5699 ( .A1(n6157), .A2(n9793), .ZN(n4296) );
  OR2_X1 U5700 ( .A1(n7923), .A2(n4435), .ZN(n4297) );
  NAND2_X1 U5701 ( .A1(n4517), .A2(n8675), .ZN(n4523) );
  AND2_X1 U5702 ( .A1(n8837), .A2(n4515), .ZN(n4514) );
  AND2_X1 U5703 ( .A1(n8006), .A2(n8005), .ZN(n9084) );
  AND4_X1 U5704 ( .A1(n6890), .A2(n6889), .A3(n6888), .A4(n6887), .ZN(n7129)
         );
  OR2_X1 U5705 ( .A1(n8483), .A2(n8374), .ZN(n4298) );
  NAND2_X1 U5706 ( .A1(n4684), .A2(n4685), .ZN(n7044) );
  NAND2_X1 U5707 ( .A1(n7337), .A2(n7336), .ZN(n8070) );
  AND2_X1 U5708 ( .A1(n4541), .A2(n4540), .ZN(n4299) );
  OR3_X1 U5709 ( .A1(n5792), .A2(n5791), .A3(n9809), .ZN(n8128) );
  INV_X1 U5710 ( .A(n5359), .ZN(n5357) );
  NAND2_X1 U5711 ( .A1(n6950), .A2(n6844), .ZN(n4301) );
  NAND2_X1 U5712 ( .A1(n4765), .A2(n4890), .ZN(n4920) );
  NAND2_X1 U5713 ( .A1(n4890), .A2(n4842), .ZN(n4895) );
  AND2_X1 U5714 ( .A1(n7183), .A2(n7553), .ZN(n4302) );
  AND2_X1 U5715 ( .A1(n4677), .A2(n7336), .ZN(n4303) );
  NAND2_X1 U5716 ( .A1(n7597), .A2(n7598), .ZN(n6229) );
  NOR2_X1 U5717 ( .A1(n7018), .A2(n4360), .ZN(n4359) );
  INV_X1 U5718 ( .A(n4823), .ZN(n4937) );
  XNOR2_X1 U5719 ( .A(n8451), .B(n8119), .ZN(n8247) );
  XNOR2_X1 U5720 ( .A(n5016), .B(n5015), .ZN(n5119) );
  NAND2_X1 U5721 ( .A1(n4534), .A2(n4532), .ZN(n9081) );
  OR2_X1 U5722 ( .A1(n4872), .A2(n4804), .ZN(n4304) );
  NAND2_X1 U5723 ( .A1(n9261), .A2(n9140), .ZN(n9042) );
  INV_X1 U5724 ( .A(n9042), .ZN(n4527) );
  INV_X1 U5725 ( .A(n9028), .ZN(n4508) );
  OR2_X1 U5726 ( .A1(n5744), .A2(n5743), .ZN(n4305) );
  NAND2_X1 U5727 ( .A1(n7580), .A2(n8411), .ZN(n7572) );
  NAND2_X1 U5728 ( .A1(n7820), .A2(n8640), .ZN(n8568) );
  NAND2_X2 U5729 ( .A1(n5359), .A2(n5652), .ZN(n7900) );
  NOR2_X1 U5730 ( .A1(n7263), .A2(n4572), .ZN(n4571) );
  AND2_X1 U5731 ( .A1(n8626), .A2(n8630), .ZN(n8629) );
  NAND2_X1 U5732 ( .A1(n7810), .A2(n7809), .ZN(n9292) );
  AND2_X1 U5733 ( .A1(n8909), .A2(n4488), .ZN(n4307) );
  INV_X1 U5734 ( .A(n7018), .ZN(n7730) );
  NAND2_X1 U5735 ( .A1(n6605), .A2(n6604), .ZN(n6824) );
  AND2_X1 U5736 ( .A1(n4370), .A2(n7656), .ZN(n4308) );
  AND2_X1 U5737 ( .A1(n7726), .A2(n6533), .ZN(n4309) );
  NAND2_X1 U5738 ( .A1(n7350), .A2(n7349), .ZN(n8477) );
  INV_X1 U5739 ( .A(n4710), .ZN(n4709) );
  NOR2_X1 U5740 ( .A1(n7693), .A2(n4711), .ZN(n4710) );
  AND2_X1 U5741 ( .A1(n4787), .A2(n6732), .ZN(n4310) );
  INV_X1 U5742 ( .A(n6229), .ZN(n7722) );
  INV_X1 U5743 ( .A(n8293), .ZN(n8460) );
  NAND2_X1 U5744 ( .A1(n7396), .A2(n7395), .ZN(n8293) );
  XNOR2_X1 U5745 ( .A(n5068), .B(SI_11_), .ZN(n5067) );
  INV_X1 U5746 ( .A(n7211), .ZN(n4671) );
  INV_X1 U5747 ( .A(n4481), .ZN(n9086) );
  NOR2_X1 U5748 ( .A1(n9125), .A2(n4482), .ZN(n4481) );
  INV_X1 U5749 ( .A(n5298), .ZN(n4463) );
  INV_X1 U5750 ( .A(n4514), .ZN(n4513) );
  INV_X1 U5751 ( .A(n9383), .ZN(n7261) );
  AND2_X1 U5752 ( .A1(n7097), .A2(n7096), .ZN(n9383) );
  AND2_X1 U5753 ( .A1(n4555), .A2(n9169), .ZN(n4311) );
  XNOR2_X1 U5754 ( .A(n8440), .B(n8200), .ZN(n8214) );
  XNOR2_X1 U5755 ( .A(n4962), .B(SI_7_), .ZN(n4959) );
  AND2_X1 U5756 ( .A1(n4783), .A2(n7018), .ZN(n4312) );
  AND2_X1 U5757 ( .A1(n4745), .A2(n7992), .ZN(n4313) );
  AND2_X1 U5758 ( .A1(n6818), .A2(n6817), .ZN(n4314) );
  NOR2_X1 U5759 ( .A1(n8446), .A2(n4386), .ZN(n4315) );
  NOR2_X1 U5760 ( .A1(n8158), .A2(n6135), .ZN(n4316) );
  NOR2_X1 U5761 ( .A1(n8460), .A2(n8134), .ZN(n4317) );
  INV_X1 U5762 ( .A(n4548), .ZN(n8210) );
  NOR2_X1 U5763 ( .A1(n8233), .A2(n8440), .ZN(n4548) );
  OR2_X1 U5764 ( .A1(n4292), .A2(n5298), .ZN(n4318) );
  AND2_X1 U5765 ( .A1(n8835), .A2(n8840), .ZN(n4319) );
  NOR2_X1 U5766 ( .A1(n7376), .A2(n7375), .ZN(n4320) );
  NAND2_X1 U5767 ( .A1(n4834), .A2(n4285), .ZN(n4321) );
  AND2_X1 U5768 ( .A1(n7695), .A2(n7694), .ZN(n8197) );
  OR2_X1 U5769 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4322) );
  AND2_X1 U5770 ( .A1(n5069), .A2(SI_11_), .ZN(n4323) );
  AND2_X1 U5771 ( .A1(n4689), .A2(n4692), .ZN(n4324) );
  NAND2_X1 U5772 ( .A1(n4933), .A2(SI_5_), .ZN(n4325) );
  INV_X1 U5773 ( .A(n4948), .ZN(n4949) );
  XNOR2_X1 U5774 ( .A(n4951), .B(SI_6_), .ZN(n4948) );
  INV_X1 U5775 ( .A(n8793), .ZN(n4521) );
  OR2_X1 U5776 ( .A1(n9008), .A2(n9005), .ZN(n4326) );
  AND2_X1 U5777 ( .A1(n4285), .A2(n4762), .ZN(n4327) );
  NOR2_X1 U5778 ( .A1(n9106), .A2(n9019), .ZN(n4328) );
  OR2_X1 U5779 ( .A1(n8503), .A2(n8106), .ZN(n7553) );
  OR2_X1 U5780 ( .A1(n8493), .A2(n8105), .ZN(n7637) );
  AND3_X1 U5781 ( .A1(n4296), .A2(n7598), .A3(n7597), .ZN(n4329) );
  AND2_X1 U5782 ( .A1(n4358), .A2(n7021), .ZN(n4330) );
  INV_X1 U5783 ( .A(n8814), .ZN(n4524) );
  NAND2_X1 U5784 ( .A1(n7773), .A2(n7772), .ZN(n8298) );
  NOR2_X1 U5785 ( .A1(n8143), .A2(n7452), .ZN(n4331) );
  NAND2_X1 U5786 ( .A1(n4824), .A2(n4581), .ZN(n4580) );
  INV_X1 U5787 ( .A(n4580), .ZN(n4516) );
  AND2_X1 U5788 ( .A1(n5295), .A2(n4463), .ZN(n4332) );
  NOR2_X1 U5789 ( .A1(n4700), .A2(n4381), .ZN(n4380) );
  INV_X1 U5790 ( .A(n6602), .ZN(n4566) );
  NAND2_X1 U5791 ( .A1(n8447), .A2(n7506), .ZN(n7682) );
  AND2_X1 U5792 ( .A1(n8900), .A2(n4491), .ZN(n4333) );
  AND2_X1 U5793 ( .A1(n4803), .A2(n5012), .ZN(n4334) );
  AND2_X1 U5794 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n4335) );
  AND2_X1 U5795 ( .A1(n4516), .A2(n5027), .ZN(n4336) );
  INV_X1 U5796 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U5797 ( .A1(n4988), .A2(n8057), .ZN(n7445) );
  XNOR2_X1 U5798 ( .A(n4582), .B(n7539), .ZN(n8743) );
  AND2_X1 U5799 ( .A1(n4573), .A2(n4571), .ZN(n4337) );
  NAND2_X1 U5800 ( .A1(n8071), .A2(n7347), .ZN(n8079) );
  NAND2_X1 U5801 ( .A1(n6556), .A2(n6555), .ZN(n6557) );
  NAND2_X1 U5802 ( .A1(n7942), .A2(n7941), .ZN(n9253) );
  INV_X1 U5803 ( .A(n9253), .ZN(n4485) );
  OR2_X1 U5804 ( .A1(n8369), .A2(n8074), .ZN(n4338) );
  AND2_X1 U5805 ( .A1(n7951), .A2(n7950), .ZN(n9017) );
  INV_X1 U5806 ( .A(n9391), .ZN(n7106) );
  AND2_X1 U5807 ( .A1(n6928), .A2(n6927), .ZN(n9391) );
  AND2_X1 U5808 ( .A1(n8349), .A2(n4551), .ZN(n4339) );
  NAND2_X1 U5809 ( .A1(n4509), .A2(n4511), .ZN(n9029) );
  NAND2_X1 U5810 ( .A1(n4792), .A2(n4338), .ZN(n8348) );
  INV_X1 U5811 ( .A(n9032), .ZN(n4503) );
  NAND2_X1 U5812 ( .A1(n4567), .A2(n6601), .ZN(n6652) );
  NAND2_X1 U5813 ( .A1(n4756), .A2(n4754), .ZN(n8599) );
  OR2_X1 U5814 ( .A1(n9253), .A2(n9017), .ZN(n9043) );
  INV_X1 U5815 ( .A(n9043), .ZN(n4538) );
  NAND2_X1 U5816 ( .A1(n5340), .A2(n4445), .ZN(n4340) );
  INV_X1 U5817 ( .A(n9033), .ZN(n4498) );
  NAND2_X1 U5818 ( .A1(n7455), .A2(n7454), .ZN(n8440) );
  INV_X1 U5819 ( .A(n8440), .ZN(n7507) );
  NAND2_X1 U5820 ( .A1(n7012), .A2(n7011), .ZN(n8508) );
  NAND2_X1 U5821 ( .A1(n4823), .A2(n4282), .ZN(n5076) );
  NAND2_X1 U5822 ( .A1(n7182), .A2(n4302), .ZN(n7503) );
  NOR3_X1 U5823 ( .A1(n7273), .A2(n9284), .A3(n4479), .ZN(n4476) );
  NAND2_X1 U5824 ( .A1(n5123), .A2(n4649), .ZN(n5641) );
  XNOR2_X1 U5825 ( .A(n7679), .B(n8043), .ZN(n8091) );
  NOR2_X1 U5826 ( .A1(n7257), .A2(n9383), .ZN(n7258) );
  NAND2_X1 U5827 ( .A1(n7178), .A2(n7177), .ZN(n7763) );
  OR2_X1 U5828 ( .A1(n9176), .A2(n9184), .ZN(n4341) );
  AND2_X1 U5829 ( .A1(n4684), .A2(n4682), .ZN(n4342) );
  INV_X1 U5830 ( .A(n4477), .ZN(n9195) );
  NOR2_X1 U5831 ( .A1(n7273), .A2(n4479), .ZN(n4477) );
  INV_X1 U5832 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U5833 ( .A1(n7337), .A2(n4303), .ZN(n8071) );
  NAND2_X1 U5834 ( .A1(n7656), .A2(n7655), .ZN(n8335) );
  INV_X1 U5835 ( .A(n7923), .ZN(n4436) );
  AND2_X1 U5836 ( .A1(n8483), .A2(n8374), .ZN(n4343) );
  AND2_X1 U5837 ( .A1(n4669), .A2(n7211), .ZN(n4344) );
  AND2_X1 U5838 ( .A1(n6000), .A2(SI_17_), .ZN(n4345) );
  NAND2_X1 U5839 ( .A1(n7958), .A2(n7957), .ZN(n4346) );
  NAND2_X1 U5840 ( .A1(n7994), .A2(n7993), .ZN(n9238) );
  INV_X1 U5841 ( .A(n9261), .ZN(n9014) );
  NAND2_X1 U5842 ( .A1(n7926), .A2(n7925), .ZN(n9261) );
  INV_X1 U5843 ( .A(n8240), .ZN(n8447) );
  AND2_X1 U5844 ( .A1(n7438), .A2(n7437), .ZN(n8240) );
  OR2_X1 U5845 ( .A1(n4343), .A2(n4791), .ZN(n4347) );
  NAND2_X1 U5846 ( .A1(n6484), .A2(n6483), .ZN(n6731) );
  OR2_X1 U5847 ( .A1(n4692), .A2(n4691), .ZN(n4348) );
  NOR2_X1 U5848 ( .A1(n5982), .A2(n6395), .ZN(n4349) );
  INV_X1 U5849 ( .A(n9493), .ZN(n4459) );
  OR2_X1 U5850 ( .A1(n5585), .A2(n5584), .ZN(n9825) );
  NAND2_X1 U5851 ( .A1(n6145), .A2(n7721), .ZN(n6230) );
  AND2_X1 U5852 ( .A1(n6177), .A2(n6176), .ZN(n4350) );
  NAND2_X1 U5853 ( .A1(n7379), .A2(n7378), .ZN(n8466) );
  INV_X1 U5854 ( .A(n8466), .ZN(n4552) );
  INV_X1 U5855 ( .A(n8567), .ZN(n4443) );
  AND2_X1 U5856 ( .A1(n7014), .A2(n4546), .ZN(n4351) );
  OAI21_X1 U5857 ( .B1(n6399), .B2(n4518), .A(n4519), .ZN(n9354) );
  NAND2_X1 U5858 ( .A1(n6143), .A2(n7589), .ZN(n6211) );
  NAND2_X1 U5859 ( .A1(n4641), .A2(n4644), .ZN(n6309) );
  INV_X1 U5860 ( .A(n4657), .ZN(n6793) );
  NAND2_X1 U5861 ( .A1(n9725), .A2(n9726), .ZN(n9724) );
  NAND2_X1 U5862 ( .A1(n4562), .A2(n6362), .ZN(n6397) );
  OR2_X1 U5863 ( .A1(n4872), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4352) );
  OR2_X1 U5864 ( .A1(n6404), .A2(n6562), .ZN(n6406) );
  INV_X1 U5865 ( .A(n6406), .ZN(n4473) );
  AND2_X1 U5866 ( .A1(n6244), .A2(n4299), .ZN(n4353) );
  AND2_X1 U5867 ( .A1(n7497), .A2(n7496), .ZN(n4354) );
  INV_X1 U5868 ( .A(n9532), .ZN(n4470) );
  XNOR2_X1 U5869 ( .A(n5011), .B(n5010), .ZN(n5115) );
  NAND2_X1 U5870 ( .A1(n6477), .A2(n6476), .ZN(n6911) );
  INV_X1 U5871 ( .A(n6911), .ZN(n4540) );
  AND2_X1 U5872 ( .A1(n5860), .A2(n6118), .ZN(n4355) );
  OAI21_X1 U5873 ( .B1(n6440), .B2(n4779), .A(n4777), .ZN(n6210) );
  OR2_X1 U5874 ( .A1(n5372), .A2(n5659), .ZN(n5666) );
  AND2_X1 U5875 ( .A1(n4462), .A2(n4292), .ZN(n4356) );
  XNOR2_X1 U5876 ( .A(n5355), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8932) );
  INV_X1 U5877 ( .A(n8253), .ZN(n8236) );
  INV_X1 U5878 ( .A(n9588), .ZN(n9128) );
  XNOR2_X1 U5879 ( .A(n5096), .B(n5095), .ZN(n6358) );
  INV_X1 U5880 ( .A(n5038), .ZN(n9319) );
  NOR2_X1 U5881 ( .A1(n4986), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8537) );
  INV_X1 U5882 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4722) );
  OR2_X1 U5883 ( .A1(n6581), .A2(n6580), .ZN(n6685) );
  NAND3_X2 U5884 ( .A1(n7820), .A2(n7839), .A3(n8640), .ZN(n8571) );
  INV_X1 U5885 ( .A(n4734), .ZN(n4732) );
  NOR2_X2 U5886 ( .A1(n6279), .A2(n6194), .ZN(n6195) );
  OAI21_X1 U5887 ( .B1(n4961), .B2(n4635), .A(n4633), .ZN(n5043) );
  NAND2_X1 U5888 ( .A1(n4909), .A2(n4908), .ZN(n4377) );
  NAND2_X1 U5889 ( .A1(n4926), .A2(SI_4_), .ZN(n4927) );
  NAND2_X1 U5890 ( .A1(n4950), .A2(n4949), .ZN(n4413) );
  INV_X1 U5891 ( .A(n8903), .ZN(n6367) );
  NAND2_X1 U5892 ( .A1(n4576), .A2(n4574), .ZN(n9080) );
  OAI22_X1 U5893 ( .A1(n6877), .A2(n8908), .B1(n6982), .B2(n4475), .ZN(n6942)
         );
  OAI21_X4 U5894 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n4722), .ZN(n4720) );
  NAND2_X1 U5895 ( .A1(n4357), .A2(n4330), .ZN(n7075) );
  INV_X1 U5896 ( .A(n6954), .ZN(n4362) );
  NAND2_X1 U5897 ( .A1(n6232), .A2(n4380), .ZN(n4379) );
  NAND3_X1 U5898 ( .A1(n4379), .A2(n4699), .A3(n4378), .ZN(n4701) );
  NAND2_X1 U5899 ( .A1(n4388), .A2(n4883), .ZN(n4898) );
  MUX2_X1 U5900 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5587), .Z(n4887) );
  MUX2_X1 U5901 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n5487), .S(n9430), .Z(n9439)
         );
  NAND3_X1 U5902 ( .A1(n4402), .A2(n4467), .A3(n4400), .ZN(P1_U3260) );
  NAND2_X1 U5903 ( .A1(n7864), .A2(n5954), .ZN(n4403) );
  NAND2_X1 U5904 ( .A1(n6458), .A2(n6457), .ZN(n6710) );
  NAND2_X1 U5905 ( .A1(n5045), .A2(n4286), .ZN(n4405) );
  NAND2_X1 U5906 ( .A1(n5045), .A2(n5044), .ZN(n5058) );
  NAND3_X1 U5907 ( .A1(n4592), .A2(n4952), .A3(n4590), .ZN(n4412) );
  NAND2_X1 U5908 ( .A1(n4412), .A2(n4411), .ZN(n4630) );
  NAND2_X2 U5909 ( .A1(n4721), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4719) );
  NAND2_X4 U5910 ( .A1(n4719), .A2(n4720), .ZN(n5587) );
  NAND2_X1 U5911 ( .A1(n5587), .A2(n4335), .ZN(n4880) );
  AND3_X2 U5912 ( .A1(n4823), .A2(n4516), .A3(n4282), .ZN(n4834) );
  AND2_X2 U5913 ( .A1(n4913), .A2(n4763), .ZN(n4823) );
  NAND2_X1 U5914 ( .A1(n7128), .A2(n4419), .ZN(n7131) );
  NAND2_X2 U5915 ( .A1(n4423), .A2(n4421), .ZN(n8591) );
  NAND3_X1 U5916 ( .A1(n4433), .A2(n4431), .A3(n4434), .ZN(n4422) );
  NAND3_X1 U5917 ( .A1(n4426), .A2(n4424), .A3(n4431), .ZN(n4423) );
  NAND2_X1 U5918 ( .A1(n4425), .A2(n4297), .ZN(n4424) );
  INV_X1 U5919 ( .A(n4434), .ZN(n4427) );
  NAND2_X1 U5920 ( .A1(n8559), .A2(n4297), .ZN(n4432) );
  NAND2_X1 U5921 ( .A1(n4428), .A2(n4434), .ZN(n8559) );
  INV_X2 U5922 ( .A(n8629), .ZN(n4434) );
  CLKBUF_X1 U5923 ( .A(n4434), .Z(n4429) );
  NOR2_X2 U5924 ( .A1(n8631), .A2(n4435), .ZN(n4433) );
  NAND2_X1 U5925 ( .A1(n8571), .A2(n4441), .ZN(n4438) );
  NAND2_X1 U5926 ( .A1(n4438), .A2(n4439), .ZN(n7885) );
  NAND2_X1 U5927 ( .A1(n5340), .A2(n4446), .ZN(n5367) );
  INV_X1 U5928 ( .A(n5367), .ZN(n4837) );
  NAND2_X1 U5929 ( .A1(n5296), .A2(n4332), .ZN(n4460) );
  INV_X1 U5930 ( .A(n4476), .ZN(n9186) );
  NAND2_X1 U5931 ( .A1(n4486), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5139) );
  NAND4_X1 U5932 ( .A1(n4285), .A2(n4823), .A3(n4579), .A4(n4282), .ZN(n4486)
         );
  AND2_X4 U5933 ( .A1(n5038), .A2(n8058), .ZN(n7983) );
  INV_X1 U5934 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4487) );
  NAND2_X1 U5935 ( .A1(n6881), .A2(n8819), .ZN(n4489) );
  INV_X1 U5936 ( .A(n5464), .ZN(n6025) );
  OAI21_X1 U5937 ( .B1(n5464), .B2(n5465), .A(n6083), .ZN(n5997) );
  XNOR2_X1 U5938 ( .A(n6024), .B(n5464), .ZN(n5480) );
  NOR2_X1 U5939 ( .A1(n8901), .A2(n5464), .ZN(n4491) );
  OR2_X1 U5940 ( .A1(n8697), .A2(n4494), .ZN(n4492) );
  OAI211_X1 U5941 ( .C1(n9589), .C2(n4493), .A(n8902), .B(n4492), .ZN(n6386)
         );
  NAND2_X1 U5942 ( .A1(n9031), .A2(n4284), .ZN(n4496) );
  NAND2_X1 U5943 ( .A1(n4496), .A2(n4497), .ZN(n9166) );
  NAND2_X1 U5944 ( .A1(n7107), .A2(n4507), .ZN(n4505) );
  INV_X1 U5945 ( .A(n7107), .ZN(n4510) );
  OAI21_X1 U5946 ( .B1(n7107), .B2(n8912), .A(n8805), .ZN(n7285) );
  NAND2_X1 U5947 ( .A1(n8912), .A2(n8805), .ZN(n4515) );
  AND2_X1 U5948 ( .A1(n4327), .A2(n4834), .ZN(n5028) );
  NAND2_X1 U5949 ( .A1(n4327), .A2(n4293), .ZN(n5030) );
  NAND2_X1 U5950 ( .A1(n9121), .A2(n9042), .ZN(n9112) );
  NAND2_X1 U5951 ( .A1(n9121), .A2(n4526), .ZN(n4525) );
  NOR2_X2 U5952 ( .A1(n9082), .A2(n4535), .ZN(n4533) );
  AOI21_X1 U5953 ( .B1(n7784), .B2(n8430), .A(n8184), .ZN(n8431) );
  NAND2_X1 U5954 ( .A1(n8349), .A2(n4549), .ZN(n8289) );
  NAND2_X1 U5955 ( .A1(n9194), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U5956 ( .A1(n4562), .A2(n4290), .ZN(n6396) );
  INV_X1 U5957 ( .A(n6651), .ZN(n4567) );
  NAND2_X1 U5958 ( .A1(n4563), .A2(n4564), .ZN(n6614) );
  NAND2_X1 U5959 ( .A1(n6650), .A2(n6602), .ZN(n4563) );
  INV_X1 U5960 ( .A(n7260), .ZN(n4569) );
  NAND2_X1 U5961 ( .A1(n9107), .A2(n4577), .ZN(n4576) );
  NAND2_X1 U5962 ( .A1(n4924), .A2(n4923), .ZN(n4594) );
  NAND2_X1 U5963 ( .A1(n5161), .A2(n4601), .ZN(n4597) );
  NAND2_X1 U5964 ( .A1(n6716), .A2(n4613), .ZN(n4611) );
  NAND2_X1 U5965 ( .A1(n7494), .A2(n4621), .ZN(n4619) );
  NAND2_X1 U5966 ( .A1(n7494), .A2(n7493), .ZN(n4620) );
  NAND3_X1 U5967 ( .A1(n4629), .A2(n4628), .A3(n4627), .ZN(n4626) );
  NAND2_X1 U5968 ( .A1(n4630), .A2(n4631), .ZN(n5045) );
  OAI211_X1 U5969 ( .C1(n4720), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n4639), .B(
        n4640), .ZN(n4899) );
  NAND3_X1 U5970 ( .A1(n4720), .A2(n4719), .A3(n5672), .ZN(n4639) );
  NAND3_X1 U5971 ( .A1(n4721), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(n5600), .ZN(
        n4640) );
  NAND3_X1 U5972 ( .A1(n4305), .A2(n5749), .A3(n5748), .ZN(n5817) );
  NAND2_X1 U5973 ( .A1(n5743), .A2(n5744), .ZN(n5749) );
  NAND2_X1 U5974 ( .A1(n9725), .A2(n4642), .ZN(n4641) );
  NAND2_X1 U5975 ( .A1(n5123), .A2(n4294), .ZN(n5643) );
  NAND2_X1 U5976 ( .A1(n6008), .A2(n4653), .ZN(n4651) );
  NAND2_X1 U5977 ( .A1(n6008), .A2(n5093), .ZN(n4652) );
  NAND2_X1 U5978 ( .A1(n6474), .A2(n4658), .ZN(n4655) );
  NAND2_X1 U5979 ( .A1(n4655), .A2(n4295), .ZN(n6798) );
  NAND2_X1 U5980 ( .A1(n6474), .A2(n6473), .ZN(n9699) );
  NOR2_X1 U5981 ( .A1(n6481), .A2(n6480), .ZN(n4660) );
  NAND2_X1 U5982 ( .A1(n4663), .A2(n4664), .ZN(n7332) );
  NAND2_X1 U5983 ( .A1(n7207), .A2(n4667), .ZN(n4663) );
  OAI21_X1 U5984 ( .B1(n6832), .B2(n4681), .A(n4678), .ZN(n7228) );
  NAND2_X1 U5985 ( .A1(n8144), .A2(n4690), .ZN(n4688) );
  NAND2_X1 U5986 ( .A1(n4688), .A2(n4348), .ZN(n8046) );
  NAND2_X1 U5987 ( .A1(n6230), .A2(n4329), .ZN(n6231) );
  NAND2_X1 U5988 ( .A1(n6143), .A2(n4696), .ZN(n4695) );
  INV_X1 U5989 ( .A(n4698), .ZN(n4699) );
  NAND2_X1 U5990 ( .A1(n4701), .A2(n7561), .ZN(n6742) );
  OAI21_X1 U5991 ( .B1(n8198), .B2(n4709), .A(n4707), .ZN(n7530) );
  NAND2_X1 U5992 ( .A1(n8198), .A2(n8197), .ZN(n8196) );
  OAI21_X1 U5993 ( .B1(n8304), .B2(n4716), .A(n4714), .ZN(n4713) );
  NAND2_X1 U5994 ( .A1(n8302), .A2(n7668), .ZN(n8280) );
  NAND3_X1 U5995 ( .A1(n4720), .A2(n4719), .A3(n4879), .ZN(n5362) );
  NAND3_X1 U5996 ( .A1(n4724), .A2(n8214), .A3(n4723), .ZN(n8213) );
  NAND2_X1 U5997 ( .A1(n5892), .A2(n5893), .ZN(n6177) );
  NAND2_X1 U5998 ( .A1(n4736), .A2(n4735), .ZN(n6198) );
  NAND3_X1 U5999 ( .A1(n5892), .A2(n5893), .A3(n6195), .ZN(n4735) );
  AOI21_X1 U6000 ( .B1(n6195), .B2(n4739), .A(n4738), .ZN(n4736) );
  NAND2_X1 U6001 ( .A1(n4737), .A2(n6195), .ZN(n6281) );
  NAND2_X1 U6002 ( .A1(n6177), .A2(n4740), .ZN(n4737) );
  INV_X1 U6003 ( .A(n6197), .ZN(n4738) );
  NAND2_X1 U6004 ( .A1(n8591), .A2(n8592), .ZN(n4748) );
  NAND2_X1 U6005 ( .A1(n8591), .A2(n4743), .ZN(n4742) );
  INV_X1 U6006 ( .A(n8592), .ZN(n4744) );
  AND2_X1 U6007 ( .A1(n4748), .A2(n4346), .ZN(n8655) );
  NAND2_X1 U6008 ( .A1(n4749), .A2(n5665), .ZN(n7484) );
  NAND2_X1 U6009 ( .A1(n5668), .A2(n5666), .ZN(n4749) );
  NAND4_X1 U6010 ( .A1(n5669), .A2(n4752), .A3(n4750), .A4(n8578), .ZN(n7487)
         );
  NAND2_X1 U6011 ( .A1(n4751), .A2(n5665), .ZN(n4750) );
  INV_X1 U6012 ( .A(n5666), .ZN(n4751) );
  NAND2_X1 U6013 ( .A1(n4753), .A2(n5665), .ZN(n4752) );
  AND2_X1 U6014 ( .A1(n5040), .A2(n4759), .ZN(n4761) );
  NAND3_X1 U6015 ( .A1(n9319), .A2(n8058), .A3(P1_REG0_REG_0__SCAN_IN), .ZN(
        n4759) );
  NAND3_X1 U6016 ( .A1(n4761), .A2(n5039), .A3(n4760), .ZN(n5463) );
  AND2_X2 U6017 ( .A1(n9319), .A2(n5032), .ZN(n5472) );
  AND2_X2 U6018 ( .A1(n9319), .A2(n8058), .ZN(n5471) );
  OAI21_X1 U6019 ( .B1(n7715), .B2(n4764), .A(n5852), .ZN(n5606) );
  NAND2_X1 U6020 ( .A1(n8244), .A2(n4768), .ZN(n4767) );
  INV_X1 U6021 ( .A(n6223), .ZN(n4776) );
  NAND2_X1 U6022 ( .A1(n6210), .A2(n7718), .ZN(n6138) );
  NAND2_X1 U6023 ( .A1(n8157), .A2(n9790), .ZN(n7591) );
  INV_X1 U6024 ( .A(n6730), .ZN(n4781) );
  NAND2_X1 U6025 ( .A1(n8385), .A2(n4790), .ZN(n4788) );
  NAND2_X1 U6026 ( .A1(n4788), .A2(n4789), .ZN(n8336) );
  NAND2_X1 U6027 ( .A1(n8385), .A2(n7768), .ZN(n8364) );
  NOR2_X1 U6028 ( .A1(n7769), .A2(n4794), .ZN(n4793) );
  INV_X1 U6029 ( .A(n7768), .ZN(n4794) );
  NAND2_X2 U6030 ( .A1(n7070), .A2(n7732), .ZN(n7175) );
  NAND2_X1 U6031 ( .A1(n4870), .A2(n4869), .ZN(n4872) );
  XNOR2_X1 U6032 ( .A(n7533), .B(SI_30_), .ZN(n8730) );
  OR2_X1 U6033 ( .A1(n5009), .A2(n4853), .ZN(n5011) );
  NAND2_X1 U6034 ( .A1(n5458), .A2(n7537), .ZN(n5685) );
  NAND2_X1 U6035 ( .A1(n7790), .A2(n8384), .ZN(n7794) );
  INV_X1 U6036 ( .A(n6023), .ZN(n6029) );
  CLKBUF_X1 U6037 ( .A(n5146), .Z(n8055) );
  NAND2_X1 U6038 ( .A1(n4851), .A2(n4850), .ZN(n5092) );
  OR2_X1 U6039 ( .A1(n9166), .A2(n9169), .ZN(n9036) );
  NAND2_X1 U6040 ( .A1(n5745), .A2(n5763), .ZN(n5747) );
  NAND2_X1 U6041 ( .A1(n10043), .A2(n8091), .ZN(n7434) );
  NAND2_X1 U6042 ( .A1(n7747), .A2(n5119), .ZN(n5741) );
  NAND2_X1 U6043 ( .A1(n7166), .A2(n7165), .ZN(n7291) );
  NAND2_X1 U6044 ( .A1(n7163), .A2(n7162), .ZN(n7166) );
  NAND2_X1 U6045 ( .A1(n6541), .A2(n6534), .ZN(n6730) );
  NAND2_X1 U6046 ( .A1(n4837), .A2(n4836), .ZN(n5127) );
  OR2_X1 U6047 ( .A1(n7540), .A2(n5586), .ZN(n5592) );
  NAND2_X1 U6048 ( .A1(n5852), .A2(n5851), .ZN(n6441) );
  NAND2_X1 U6049 ( .A1(n5763), .A2(n5593), .ZN(n5743) );
  NAND2_X2 U6050 ( .A1(n5602), .A2(n7537), .ZN(n7540) );
  INV_X1 U6051 ( .A(n7715), .ZN(n5608) );
  AND2_X2 U6052 ( .A1(n5101), .A2(n5100), .ZN(n5775) );
  INV_X1 U6053 ( .A(n4988), .ZN(n5101) );
  OR2_X1 U6054 ( .A1(n5028), .A2(n4915), .ZN(n5026) );
  NAND2_X1 U6055 ( .A1(n6685), .A2(n6684), .ZN(n4806) );
  AND2_X1 U6056 ( .A1(n5767), .A2(n5766), .ZN(n4807) );
  AND4_X1 U6057 ( .A1(n6936), .A2(n6935), .A3(n6934), .A4(n6933), .ZN(n7257)
         );
  AND2_X1 U6058 ( .A1(n9091), .A2(n9075), .ZN(n4808) );
  AND2_X1 U6059 ( .A1(n7320), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4809) );
  INV_X1 U6060 ( .A(n5471), .ZN(n5690) );
  NAND2_X1 U6061 ( .A1(n5386), .A2(n5466), .ZN(n4810) );
  NAND2_X1 U6062 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n4811) );
  NAND2_X1 U6063 ( .A1(n5025), .A2(n5024), .ZN(n4812) );
  AND2_X1 U6064 ( .A1(n5044), .A2(n5002), .ZN(n4813) );
  AND2_X1 U6065 ( .A1(n5339), .A2(n5166), .ZN(n4814) );
  AND2_X1 U6066 ( .A1(n5059), .A2(n5050), .ZN(n4815) );
  INV_X1 U6067 ( .A(n8650), .ZN(n8652) );
  AND2_X1 U6068 ( .A1(n7478), .A2(n7477), .ZN(n7779) );
  INV_X1 U6069 ( .A(n8200), .ZN(n7777) );
  XOR2_X1 U6070 ( .A(n8293), .B(n8043), .Z(n4816) );
  INV_X1 U6071 ( .A(n8896), .ZN(n6601) );
  AND2_X1 U6072 ( .A1(n7406), .A2(n7405), .ZN(n8284) );
  AND2_X1 U6073 ( .A1(n8433), .A2(n8432), .ZN(n4817) );
  INV_X1 U6074 ( .A(n8435), .ZN(n7780) );
  INV_X1 U6075 ( .A(n8508), .ZN(n7013) );
  OAI21_X1 U6076 ( .B1(n8259), .B2(n8267), .A(n7774), .ZN(n8243) );
  XNOR2_X1 U6078 ( .A(n8454), .B(n7439), .ZN(n8116) );
  NAND2_X1 U6079 ( .A1(n8336), .A2(n8335), .ZN(n8337) );
  INV_X1 U6080 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4820) );
  INV_X1 U6081 ( .A(n7546), .ZN(n7543) );
  INV_X1 U6082 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4819) );
  INV_X1 U6083 ( .A(n6335), .ZN(n6332) );
  AND2_X1 U6084 ( .A1(n7415), .A2(n8115), .ZN(n7419) );
  AND2_X1 U6085 ( .A1(n5512), .A2(n5511), .ZN(n5722) );
  AND2_X1 U6086 ( .A1(n8181), .A2(n8148), .ZN(n7792) );
  INV_X1 U6087 ( .A(n7733), .ZN(n7183) );
  INV_X1 U6088 ( .A(n7719), .ZN(n7576) );
  INV_X1 U6089 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U6090 ( .A1(n7974), .A2(n5463), .ZN(n5371) );
  NAND2_X1 U6091 ( .A1(n4806), .A2(n6681), .ZN(n6688) );
  INV_X1 U6092 ( .A(n7278), .ZN(n7277) );
  INV_X1 U6093 ( .A(n7944), .ZN(n7943) );
  INV_X1 U6094 ( .A(n7912), .ZN(n7910) );
  OR2_X1 U6095 ( .A1(n7869), .A2(n7868), .ZN(n7891) );
  NAND2_X1 U6096 ( .A1(n8684), .A2(n6030), .ZN(n9606) );
  INV_X1 U6097 ( .A(n4959), .ZN(n4960) );
  OR2_X1 U6098 ( .A1(n6745), .A2(n6744), .ZN(n6838) );
  INV_X1 U6099 ( .A(n8041), .ZN(n6325) );
  INV_X1 U6100 ( .A(n8451), .ZN(n7679) );
  OR2_X1 U6101 ( .A1(n6098), .A2(n5790), .ZN(n5793) );
  OR2_X1 U6102 ( .A1(n7441), .A2(n7440), .ZN(n7470) );
  AOI21_X1 U6103 ( .B1(n8217), .B2(n8419), .A(n7792), .ZN(n7793) );
  OR2_X1 U6104 ( .A1(n7426), .A2(n8095), .ZN(n7441) );
  INV_X1 U6105 ( .A(n7724), .ZN(n6531) );
  OR2_X1 U6106 ( .A1(n6628), .A2(n6627), .ZN(n6885) );
  INV_X1 U6107 ( .A(n7100), .ZN(n7098) );
  NAND2_X1 U6108 ( .A1(n7889), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7912) );
  INV_X1 U6109 ( .A(n7816), .ZN(n7819) );
  NAND2_X1 U6110 ( .A1(n7910), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7928) );
  AOI21_X1 U6111 ( .B1(n9073), .B2(n9050), .A(n9049), .ZN(n9052) );
  NOR2_X1 U6112 ( .A1(n9200), .A2(n9185), .ZN(n9005) );
  AND2_X1 U6113 ( .A1(n8798), .A2(n8819), .ZN(n8908) );
  NAND2_X1 U6114 ( .A1(n6456), .A2(n6455), .ZN(n6458) );
  NAND2_X1 U6115 ( .A1(n5048), .A2(n5047), .ZN(n5059) );
  NAND2_X1 U6116 ( .A1(n5830), .A2(n5832), .ZN(n5831) );
  AND3_X1 U6117 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U6118 ( .A1(n7186), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7318) );
  INV_X1 U6119 ( .A(n8214), .ZN(n8207) );
  INV_X1 U6120 ( .A(n8279), .ZN(n8275) );
  INV_X1 U6121 ( .A(n7726), .ZN(n6538) );
  INV_X1 U6122 ( .A(n7766), .ZN(n8388) );
  NAND2_X1 U6123 ( .A1(n7980), .A2(n6363), .ZN(n7982) );
  NAND2_X1 U6124 ( .A1(n6884), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U6125 ( .A1(n6069), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6373) );
  OR2_X1 U6126 ( .A1(n7938), .A2(n7937), .ZN(n7939) );
  OR2_X1 U6127 ( .A1(n6373), .A2(n6372), .ZN(n6380) );
  INV_X1 U6128 ( .A(n5386), .ZN(n5393) );
  OR2_X1 U6129 ( .A1(n9109), .A2(n8020), .ZN(n7951) );
  INV_X1 U6130 ( .A(n9005), .ZN(n9006) );
  AND2_X1 U6131 ( .A1(n8804), .A2(n8828), .ZN(n8909) );
  OR2_X1 U6132 ( .A1(n8877), .A2(n8932), .ZN(n9638) );
  AND2_X1 U6133 ( .A1(n4942), .A2(n4941), .ZN(n9624) );
  NAND2_X1 U6134 ( .A1(n4900), .A2(SI_2_), .ZN(n4901) );
  OR3_X1 U6135 ( .A1(n6925), .A2(n7063), .A3(n7122), .ZN(n5796) );
  AND2_X1 U6136 ( .A1(n5935), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U6138 ( .A1(n8041), .A2(n7549), .ZN(n7753) );
  AND2_X1 U6139 ( .A1(n7432), .A2(n7431), .ZN(n8119) );
  AND4_X1 U6140 ( .A1(n6347), .A2(n6346), .A3(n6345), .A4(n6344), .ZN(n6662)
         );
  AND2_X1 U6141 ( .A1(n5244), .A2(n5615), .ZN(n9749) );
  NOR2_X1 U6142 ( .A1(n8432), .A2(n8402), .ZN(n7795) );
  AND2_X1 U6143 ( .A1(n7646), .A2(n7652), .ZN(n8371) );
  OR2_X1 U6144 ( .A1(n9766), .A2(n5099), .ZN(n6098) );
  AND2_X1 U6145 ( .A1(n8376), .A2(n8375), .ZN(n8490) );
  AND2_X1 U6146 ( .A1(n5081), .A2(n5080), .ZN(n9762) );
  AND2_X1 U6147 ( .A1(n8027), .A2(n8026), .ZN(n9074) );
  AND4_X1 U6148 ( .A1(n7105), .A2(n7104), .A3(n7103), .A4(n7102), .ZN(n7294)
         );
  NOR2_X1 U6149 ( .A1(n5292), .A2(n5291), .ZN(n8956) );
  INV_X1 U6150 ( .A(n8993), .ZN(n9229) );
  AND2_X1 U6151 ( .A1(n8894), .A2(n9032), .ZN(n9203) );
  INV_X1 U6152 ( .A(n9608), .ZN(n9359) );
  OR2_X1 U6153 ( .A1(n9638), .A2(n5391), .ZN(n9618) );
  NOR2_X1 U6154 ( .A1(n9370), .A2(n9680), .ZN(n9371) );
  OR2_X1 U6155 ( .A1(n5486), .A2(n5979), .ZN(n5625) );
  INV_X1 U6156 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4938) );
  XNOR2_X1 U6157 ( .A(n4910), .B(SI_3_), .ZN(n4908) );
  INV_X1 U6158 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6784) );
  OR2_X1 U6159 ( .A1(n8142), .A2(n8330), .ZN(n9714) );
  INV_X1 U6160 ( .A(n9717), .ZN(n8135) );
  AND2_X1 U6161 ( .A1(n7196), .A2(n7195), .ZN(n8502) );
  INV_X1 U6162 ( .A(n9764), .ZN(n9767) );
  INV_X1 U6163 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5758) );
  INV_X1 U6164 ( .A(n9288), .ZN(n9200) );
  INV_X1 U6165 ( .A(n8648), .ZN(n8663) );
  NAND2_X1 U6166 ( .A1(n7970), .A2(n7969), .ZN(n9114) );
  INV_X1 U6167 ( .A(n9454), .ZN(n9564) );
  OAI21_X1 U6168 ( .B1(n9066), .B2(n9072), .A(n9065), .ZN(n9242) );
  NAND2_X1 U6169 ( .A1(n6079), .A2(n9618), .ZN(n9617) );
  OR2_X1 U6170 ( .A1(n5625), .A2(n9628), .ZN(n9686) );
  INV_X1 U6171 ( .A(n9626), .ZN(n9627) );
  AND3_X1 U6172 ( .A1(n5651), .A2(n5652), .A3(P1_STATE_REG_SCAN_IN), .ZN(n9630) );
  NOR2_X1 U6173 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4822) );
  NOR2_X1 U6174 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4821) );
  INV_X1 U6175 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4824) );
  INV_X1 U6176 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5579) );
  INV_X1 U6177 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6003) );
  INV_X1 U6178 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4825) );
  NOR2_X1 U6179 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4828) );
  NOR2_X1 U6180 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4827) );
  NOR2_X1 U6181 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4826) );
  INV_X1 U6182 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4830) );
  INV_X1 U6183 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U6184 ( .A1(n5139), .A2(n5022), .ZN(n4833) );
  NAND2_X1 U6185 ( .A1(n4833), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4829) );
  INV_X1 U6186 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5023) );
  XNOR2_X1 U6187 ( .A(n4829), .B(n5023), .ZN(n7124) );
  NAND2_X1 U6188 ( .A1(n4321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4831) );
  XNOR2_X1 U6189 ( .A(n4831), .B(n4830), .ZN(n6988) );
  OR2_X1 U6190 ( .A1(n5139), .A2(n5022), .ZN(n4832) );
  NAND2_X1 U6191 ( .A1(n4833), .A2(n4832), .ZN(n7064) );
  OR3_X2 U6192 ( .A1(n7124), .A2(n6988), .A3(n7064), .ZN(n5652) );
  INV_X1 U6193 ( .A(n5652), .ZN(n4841) );
  NOR2_X1 U6194 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4835) );
  INV_X1 U6195 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5129) );
  INV_X1 U6196 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5130) );
  NAND3_X1 U6197 ( .A1(n5129), .A2(n5128), .A3(n5130), .ZN(n4838) );
  OAI21_X1 U6198 ( .B1(n5127), .B2(n4838), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4840) );
  INV_X1 U6199 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4839) );
  XNOR2_X1 U6200 ( .A(n4840), .B(n4839), .ZN(n5651) );
  NAND2_X1 U6201 ( .A1(n4841), .A2(n5651), .ZN(n5423) );
  OR2_X2 U6202 ( .A1(n5423), .A2(P1_U3084), .ZN(n8954) );
  INV_X1 U6203 ( .A(n8954), .ZN(P1_U4006) );
  NOR2_X1 U6204 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4846) );
  NOR2_X1 U6205 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4845) );
  NOR2_X1 U6206 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4844) );
  NOR2_X1 U6207 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4843) );
  NAND4_X1 U6208 ( .A1(n4846), .A2(n4845), .A3(n4844), .A4(n4843), .ZN(n4847)
         );
  BUF_X1 U6209 ( .A(n4870), .Z(n5123) );
  INV_X1 U6210 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4848) );
  INV_X1 U6211 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5413) );
  INV_X1 U6212 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4864) );
  AND3_X1 U6213 ( .A1(n5416), .A2(n5413), .A3(n4864), .ZN(n4849) );
  INV_X1 U6214 ( .A(n5643), .ZN(n4851) );
  INV_X1 U6215 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4850) );
  INV_X1 U6216 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5093) );
  INV_X1 U6217 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5094) );
  INV_X1 U6218 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5095) );
  NAND3_X1 U6219 ( .A1(n5093), .A2(n5094), .A3(n5095), .ZN(n4852) );
  INV_X1 U6220 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U6221 ( .A1(n5017), .A2(n4865), .ZN(n4854) );
  INV_X1 U6222 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4853) );
  INV_X1 U6223 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U6224 ( .A1(n5016), .A2(n5015), .ZN(n4855) );
  NAND2_X1 U6225 ( .A1(n4855), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4877) );
  INV_X1 U6226 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4856) );
  NAND2_X1 U6227 ( .A1(n4877), .A2(n4856), .ZN(n4857) );
  NAND2_X1 U6228 ( .A1(n4857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4859) );
  INV_X1 U6229 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4858) );
  XNOR2_X1 U6230 ( .A(n4859), .B(n4858), .ZN(n6925) );
  NOR2_X1 U6231 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4863) );
  NOR2_X1 U6232 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4862) );
  NOR2_X1 U6233 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4861) );
  NOR2_X1 U6234 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n4860) );
  NAND4_X1 U6235 ( .A1(n4863), .A2(n4862), .A3(n4861), .A4(n4860), .ZN(n4868)
         );
  NOR2_X1 U6236 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4866) );
  NAND4_X1 U6237 ( .A1(n4866), .A2(n4865), .A3(n4864), .A4(n5416), .ZN(n4867)
         );
  NOR2_X1 U6238 ( .A1(n4868), .A2(n4867), .ZN(n4869) );
  NAND2_X1 U6239 ( .A1(n4872), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4871) );
  MUX2_X1 U6240 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4871), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n4873) );
  NAND2_X1 U6241 ( .A1(n4873), .A2(n4352), .ZN(n7063) );
  NAND2_X1 U6242 ( .A1(n4352), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4874) );
  MUX2_X1 U6243 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4874), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n4876) );
  NAND2_X1 U6244 ( .A1(n4876), .A2(n4304), .ZN(n7122) );
  INV_X1 U6245 ( .A(n5796), .ZN(n5199) );
  XNOR2_X1 U6246 ( .A(n4877), .B(P2_IR_REG_23__SCAN_IN), .ZN(n5794) );
  NOR2_X1 U6247 ( .A1(n5794), .A2(P2_U3152), .ZN(n9769) );
  AND2_X1 U6248 ( .A1(n5199), .A2(n9769), .ZN(P2_U3966) );
  NOR2_X1 U6249 ( .A1(n5587), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9323) );
  AND2_X1 U6250 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4879) );
  INV_X1 U6251 ( .A(SI_1_), .ZN(n4881) );
  XNOR2_X1 U6252 ( .A(n4882), .B(n4881), .ZN(n4888) );
  NAND2_X1 U6253 ( .A1(n4882), .A2(SI_1_), .ZN(n4883) );
  XNOR2_X1 U6254 ( .A(n4898), .B(n4897), .ZN(n5671) );
  OAI222_X1 U6255 ( .A1(n9328), .A2(n5672), .B1(n8059), .B2(n5671), .C1(
        P1_U3084), .C2(n5675), .ZN(P1_U3351) );
  NOR2_X1 U6256 ( .A1(n5587), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8540) );
  INV_X1 U6257 ( .A(n8540), .ZN(n8545) );
  INV_X1 U6258 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5586) );
  AND2_X1 U6259 ( .A1(n5587), .A2(P2_U3152), .ZN(n6728) );
  XNOR2_X1 U6260 ( .A(n4888), .B(n4887), .ZN(n5588) );
  NAND2_X1 U6261 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4889) );
  MUX2_X1 U6262 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4889), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n4892) );
  INV_X1 U6263 ( .A(n4890), .ZN(n4891) );
  NAND2_X1 U6264 ( .A1(n4892), .A2(n4891), .ZN(n5589) );
  OAI222_X1 U6265 ( .A1(n8545), .A2(n5586), .B1(n4270), .B2(n5588), .C1(
        P2_U3152), .C2(n5589), .ZN(P2_U3357) );
  NOR2_X1 U6266 ( .A1(n4890), .A2(n4853), .ZN(n4893) );
  MUX2_X1 U6267 ( .A(n4853), .B(n4893), .S(P2_IR_REG_2__SCAN_IN), .Z(n4894) );
  INV_X1 U6268 ( .A(n4894), .ZN(n4896) );
  NAND2_X1 U6269 ( .A1(n4896), .A2(n4895), .ZN(n5601) );
  OAI222_X1 U6270 ( .A1(n8545), .A2(n5600), .B1(n4270), .B2(n5671), .C1(
        P2_U3152), .C2(n5601), .ZN(P2_U3356) );
  NAND2_X1 U6271 ( .A1(n4898), .A2(n4897), .ZN(n4902) );
  INV_X1 U6272 ( .A(n4899), .ZN(n4900) );
  MUX2_X1 U6273 ( .A(n5758), .B(n5687), .S(n4276), .Z(n4910) );
  XNOR2_X1 U6274 ( .A(n4909), .B(n4908), .ZN(n5757) );
  NAND2_X1 U6275 ( .A1(n4895), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4904) );
  INV_X1 U6276 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4903) );
  XNOR2_X1 U6277 ( .A(n4904), .B(n4903), .ZN(n5759) );
  OAI222_X1 U6278 ( .A1(n8545), .A2(n5758), .B1(n4270), .B2(n5757), .C1(
        P2_U3152), .C2(n5759), .ZN(P2_U3355) );
  INV_X1 U6279 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4906) );
  OAI222_X1 U6280 ( .A1(n9328), .A2(n5687), .B1(n8059), .B2(n5757), .C1(
        P1_U3084), .C2(n9330), .ZN(P1_U3350) );
  INV_X1 U6281 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5457) );
  INV_X1 U6282 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4907) );
  OAI222_X1 U6283 ( .A1(n9328), .A2(n5457), .B1(n8059), .B2(n5588), .C1(
        P1_U3084), .C2(n9430), .ZN(P1_U3352) );
  INV_X1 U6284 ( .A(n4910), .ZN(n4911) );
  INV_X1 U6285 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5770) );
  INV_X4 U6286 ( .A(n5587), .ZN(n7537) );
  MUX2_X1 U6287 ( .A(n5770), .B(n10001), .S(n7537), .Z(n4925) );
  XNOR2_X2 U6288 ( .A(n4925), .B(SI_4_), .ZN(n4923) );
  INV_X1 U6289 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4915) );
  NOR2_X1 U6290 ( .A1(n4913), .A2(n4915), .ZN(n4914) );
  MUX2_X1 U6291 ( .A(n4915), .B(n4914), .S(P1_IR_REG_4__SCAN_IN), .Z(n4916) );
  INV_X1 U6292 ( .A(n4916), .ZN(n4919) );
  INV_X1 U6293 ( .A(n4917), .ZN(n4918) );
  NAND2_X1 U6294 ( .A1(n4919), .A2(n4918), .ZN(n5885) );
  OAI222_X1 U6295 ( .A1(n9328), .A2(n10001), .B1(n8059), .B2(n5882), .C1(
        P1_U3084), .C2(n5885), .ZN(P1_U3349) );
  NAND2_X1 U6296 ( .A1(n4920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4922) );
  INV_X1 U6297 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4921) );
  XNOR2_X1 U6298 ( .A(n4922), .B(n4921), .ZN(n5771) );
  OAI222_X1 U6299 ( .A1(n8545), .A2(n5770), .B1(n4270), .B2(n5882), .C1(
        P2_U3152), .C2(n5771), .ZN(P2_U3354) );
  INV_X1 U6300 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6035) );
  INV_X1 U6301 ( .A(n4925), .ZN(n4926) );
  MUX2_X1 U6302 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4276), .Z(n4933) );
  XNOR2_X1 U6303 ( .A(n4932), .B(n4930), .ZN(n5923) );
  INV_X1 U6304 ( .A(n5923), .ZN(n6034) );
  OR2_X1 U6305 ( .A1(n4917), .A2(n4915), .ZN(n4929) );
  XNOR2_X1 U6306 ( .A(n4929), .B(n4928), .ZN(n6038) );
  OAI222_X1 U6307 ( .A1(n9328), .A2(n6035), .B1(n8059), .B2(n6034), .C1(
        P1_U3084), .C2(n6038), .ZN(P1_U3348) );
  INV_X1 U6308 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5925) );
  NOR2_X1 U6309 ( .A1(n4920), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n4973) );
  OR2_X1 U6310 ( .A1(n4973), .A2(n4853), .ZN(n4934) );
  XNOR2_X1 U6311 ( .A(n4934), .B(P2_IR_REG_5__SCAN_IN), .ZN(n5529) );
  INV_X1 U6312 ( .A(n5529), .ZN(n5924) );
  OAI222_X1 U6313 ( .A1(n8545), .A2(n5925), .B1(n4270), .B2(n6034), .C1(
        P2_U3152), .C2(n5924), .ZN(P2_U3353) );
  MUX2_X1 U6314 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4276), .Z(n4951) );
  XNOR2_X1 U6315 ( .A(n4950), .B(n4948), .ZN(n5908) );
  INV_X1 U6316 ( .A(n5908), .ZN(n6040) );
  INV_X1 U6317 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U6318 ( .A1(n4934), .A2(n4971), .ZN(n4935) );
  NAND2_X1 U6319 ( .A1(n4935), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4953) );
  XNOR2_X1 U6320 ( .A(n4953), .B(P2_IR_REG_6__SCAN_IN), .ZN(n5909) );
  AOI22_X1 U6321 ( .A1(n5909), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8540), .ZN(n4936) );
  OAI21_X1 U6322 ( .B1(n6040), .B2(n4270), .A(n4936), .ZN(P2_U3352) );
  INV_X1 U6323 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U6324 ( .A1(n4937), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4939) );
  XNOR2_X1 U6325 ( .A(n4939), .B(n4938), .ZN(n6044) );
  OAI222_X1 U6326 ( .A1(n9328), .A2(n6041), .B1(n8059), .B2(n6040), .C1(
        P1_U3084), .C2(n6044), .ZN(P1_U3347) );
  INV_X1 U6327 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U6328 ( .A1(n7064), .A2(P1_B_REG_SCAN_IN), .ZN(n4940) );
  MUX2_X1 U6329 ( .A(P1_B_REG_SCAN_IN), .B(n4940), .S(n6988), .Z(n4942) );
  INV_X1 U6330 ( .A(n7124), .ZN(n4941) );
  NAND2_X1 U6331 ( .A1(n9624), .A2(n4947), .ZN(n4944) );
  NAND2_X1 U6332 ( .A1(n7124), .A2(n7064), .ZN(n4943) );
  NAND2_X1 U6333 ( .A1(n4944), .A2(n4943), .ZN(n5485) );
  INV_X1 U6334 ( .A(n5485), .ZN(n4945) );
  NAND2_X1 U6335 ( .A1(n4945), .A2(n9630), .ZN(n4946) );
  OAI21_X1 U6336 ( .B1(n9630), .B2(n4947), .A(n4946), .ZN(P1_U3441) );
  NAND2_X1 U6337 ( .A1(n4951), .A2(SI_6_), .ZN(n4952) );
  MUX2_X1 U6338 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4276), .Z(n4962) );
  INV_X1 U6339 ( .A(n6053), .ZN(n4958) );
  INV_X1 U6340 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6341 ( .A1(n4953), .A2(n4970), .ZN(n4954) );
  NAND2_X1 U6342 ( .A1(n4954), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4955) );
  XNOR2_X1 U6343 ( .A(n4955), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9756) );
  AOI22_X1 U6344 ( .A1(n9756), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n8540), .ZN(n4956) );
  OAI21_X1 U6345 ( .B1(n4958), .B2(n4270), .A(n4956), .ZN(P2_U3351) );
  INV_X1 U6346 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6055) );
  OR2_X1 U6347 ( .A1(n4937), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6348 ( .A1(n4976), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4957) );
  XNOR2_X1 U6349 ( .A(n4957), .B(P1_IR_REG_7__SCAN_IN), .ZN(n5544) );
  INV_X1 U6350 ( .A(n5544), .ZN(n6054) );
  OAI222_X1 U6351 ( .A1(n9328), .A2(n6055), .B1(n8059), .B2(n4958), .C1(
        P1_U3084), .C2(n6054), .ZN(P1_U3346) );
  NAND2_X1 U6352 ( .A1(n4962), .A2(SI_7_), .ZN(n4963) );
  INV_X1 U6353 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n4964) );
  INV_X1 U6354 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n4983) );
  MUX2_X1 U6355 ( .A(n4964), .B(n4983), .S(n4276), .Z(n4966) );
  INV_X1 U6356 ( .A(SI_8_), .ZN(n4965) );
  INV_X1 U6357 ( .A(n4966), .ZN(n4967) );
  NAND2_X1 U6358 ( .A1(n4967), .A2(SI_8_), .ZN(n4968) );
  XNOR2_X1 U6359 ( .A(n4996), .B(n4995), .ZN(n6364) );
  INV_X1 U6360 ( .A(n6364), .ZN(n4982) );
  INV_X1 U6361 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4969) );
  AND3_X1 U6362 ( .A1(n4971), .A2(n4970), .A3(n4969), .ZN(n4972) );
  NAND2_X1 U6363 ( .A1(n4973), .A2(n4972), .ZN(n5003) );
  NAND2_X1 U6364 ( .A1(n5003), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4974) );
  XNOR2_X1 U6365 ( .A(n4974), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6224) );
  AOI22_X1 U6366 ( .A1(n6224), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n8540), .ZN(n4975) );
  OAI21_X1 U6367 ( .B1(n4982), .B2(n4270), .A(n4975), .ZN(P2_U3350) );
  NOR2_X1 U6368 ( .A1(n4976), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n4979) );
  NOR2_X1 U6369 ( .A1(n4979), .A2(n4915), .ZN(n4977) );
  MUX2_X1 U6370 ( .A(n4915), .B(n4977), .S(P1_IR_REG_8__SCAN_IN), .Z(n4981) );
  INV_X1 U6371 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U6372 ( .A1(n4979), .A2(n4978), .ZN(n5051) );
  INV_X1 U6373 ( .A(n5051), .ZN(n4980) );
  OR2_X1 U6374 ( .A1(n4981), .A2(n4980), .ZN(n9451) );
  OAI222_X1 U6375 ( .A1(n9328), .A2(n4983), .B1(n8059), .B2(n4982), .C1(
        P1_U3084), .C2(n9451), .ZN(P1_U3345) );
  INV_X1 U6376 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6377 ( .A1(n5009), .A2(n5010), .ZN(n4986) );
  INV_X1 U6378 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6379 ( .A1(n4986), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4987) );
  INV_X1 U6380 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9995) );
  INV_X1 U6381 ( .A(n8057), .ZN(n5100) );
  AND2_X4 U6382 ( .A1(n4988), .A2(n5100), .ZN(n5609) );
  NAND2_X1 U6383 ( .A1(n5609), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U6384 ( .A1(n5595), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U6385 ( .A1(n7525), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n4989) );
  AND3_X1 U6386 ( .A1(n4991), .A2(n4990), .A3(n4989), .ZN(n7546) );
  NAND2_X1 U6387 ( .A1(P2_U3966), .A2(n7543), .ZN(n4992) );
  OAI21_X1 U6388 ( .B1(P2_U3966), .B2(n4993), .A(n4992), .ZN(P2_U3583) );
  INV_X1 U6389 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n4998) );
  INV_X1 U6390 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4997) );
  MUX2_X1 U6391 ( .A(n4998), .B(n4997), .S(n4276), .Z(n5000) );
  INV_X1 U6392 ( .A(SI_9_), .ZN(n4999) );
  INV_X1 U6393 ( .A(n5000), .ZN(n5001) );
  NAND2_X1 U6394 ( .A1(n5001), .A2(SI_9_), .ZN(n5002) );
  XNOR2_X1 U6395 ( .A(n5043), .B(n4813), .ZN(n6369) );
  INV_X1 U6396 ( .A(n6369), .ZN(n5008) );
  OR2_X1 U6397 ( .A1(n5003), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6398 ( .A1(n5054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5004) );
  XNOR2_X1 U6399 ( .A(n5004), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6322) );
  AOI22_X1 U6400 ( .A1(n6322), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n8540), .ZN(n5005) );
  OAI21_X1 U6401 ( .B1(n5008), .B2(n4270), .A(n5005), .ZN(P2_U3349) );
  NAND2_X1 U6402 ( .A1(n5051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5006) );
  XNOR2_X1 U6403 ( .A(n5006), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9467) );
  INV_X1 U6404 ( .A(n9328), .ZN(n5848) );
  AOI22_X1 U6405 ( .A1(n9467), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n5848), .ZN(n5007) );
  OAI21_X1 U6406 ( .B1(n5008), .B2(n8059), .A(n5007), .ZN(P1_U3344) );
  NAND2_X1 U6407 ( .A1(n5796), .A2(n9769), .ZN(n9763) );
  NAND2_X1 U6408 ( .A1(n5794), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7760) );
  NAND2_X1 U6409 ( .A1(n9763), .A2(n7760), .ZN(n5014) );
  INV_X1 U6410 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5012) );
  NAND2_X2 U6411 ( .A1(n5115), .A2(n7756), .ZN(n5602) );
  NAND2_X1 U6412 ( .A1(n5014), .A2(n7338), .ZN(n5021) );
  INV_X1 U6413 ( .A(n5119), .ZN(n7757) );
  OR2_X1 U6414 ( .A1(n5017), .A2(n4853), .ZN(n5018) );
  XNOR2_X1 U6415 ( .A(n5018), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5118) );
  AND2_X1 U6416 ( .A1(n7757), .A2(n5118), .ZN(n5791) );
  INV_X1 U6417 ( .A(n5791), .ZN(n5019) );
  OR2_X1 U6418 ( .A1(n9763), .A2(n5019), .ZN(n5020) );
  NAND2_X1 U6419 ( .A1(n5021), .A2(n5020), .ZN(n9747) );
  NOR2_X1 U6420 ( .A1(P2_U3966), .A2(n9747), .ZN(P2_U3151) );
  INV_X1 U6421 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6422 ( .A1(n5023), .A2(n5022), .ZN(n5137) );
  INV_X1 U6423 ( .A(n5137), .ZN(n5025) );
  NOR2_X1 U6424 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5024) );
  INV_X1 U6425 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6426 ( .A1(n7983), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U6427 ( .A1(n4275), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5034) );
  INV_X2 U6428 ( .A(n5690), .ZN(n8735) );
  NAND2_X1 U6429 ( .A1(n8735), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5033) );
  NAND3_X1 U6430 ( .A1(n5035), .A2(n5034), .A3(n5033), .ZN(n8771) );
  NAND2_X1 U6431 ( .A1(P1_U4006), .A2(n8771), .ZN(n5036) );
  OAI21_X1 U6432 ( .B1(P1_U4006), .B2(n5037), .A(n5036), .ZN(P1_U3586) );
  INV_X1 U6433 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6434 ( .A1(n4281), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U6435 ( .A1(n7983), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5039) );
  NAND2_X1 U6436 ( .A1(P1_U4006), .A2(n5463), .ZN(n5041) );
  OAI21_X1 U6437 ( .B1(P1_U4006), .B2(n5042), .A(n5041), .ZN(P1_U3555) );
  INV_X1 U6438 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5056) );
  INV_X1 U6439 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5046) );
  MUX2_X1 U6440 ( .A(n5056), .B(n5046), .S(n4276), .Z(n5048) );
  INV_X1 U6441 ( .A(SI_10_), .ZN(n5047) );
  INV_X1 U6442 ( .A(n5048), .ZN(n5049) );
  NAND2_X1 U6443 ( .A1(n5049), .A2(SI_10_), .ZN(n5050) );
  XNOR2_X1 U6444 ( .A(n5058), .B(n4815), .ZN(n6598) );
  INV_X1 U6445 ( .A(n6598), .ZN(n5057) );
  OR2_X1 U6446 ( .A1(n5051), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6447 ( .A1(n5060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5052) );
  XNOR2_X1 U6448 ( .A(n5052), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9479) );
  AOI22_X1 U6449 ( .A1(n9479), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n5848), .ZN(n5053) );
  OAI21_X1 U6450 ( .B1(n5057), .B2(n8059), .A(n5053), .ZN(P1_U3343) );
  OR2_X1 U6451 ( .A1(n5054), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U6452 ( .A1(n5063), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5055) );
  XNOR2_X1 U6453 ( .A(n5055), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6475) );
  INV_X1 U6454 ( .A(n6475), .ZN(n5334) );
  OAI222_X1 U6455 ( .A1(P2_U3152), .A2(n5334), .B1(n4270), .B2(n5057), .C1(
        n5056), .C2(n8545), .ZN(P2_U3348) );
  INV_X1 U6456 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5066) );
  INV_X1 U6457 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5062) );
  MUX2_X1 U6458 ( .A(n5066), .B(n5062), .S(n7537), .Z(n5068) );
  XNOR2_X1 U6459 ( .A(n5070), .B(n5067), .ZN(n6603) );
  INV_X1 U6460 ( .A(n6603), .ZN(n5065) );
  OAI21_X1 U6461 ( .B1(n5060), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5061) );
  XNOR2_X1 U6462 ( .A(n5061), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8970) );
  INV_X1 U6463 ( .A(n8970), .ZN(n8957) );
  OAI222_X1 U6464 ( .A1(n8059), .A2(n5065), .B1(n8957), .B2(P1_U3084), .C1(
        n5062), .C2(n9328), .ZN(P1_U3342) );
  OAI21_X1 U6465 ( .B1(n5063), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5064) );
  XNOR2_X1 U6466 ( .A(n5064), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6482) );
  INV_X1 U6467 ( .A(n6482), .ZN(n5508) );
  OAI222_X1 U6468 ( .A1(n8545), .A2(n5066), .B1(n4270), .B2(n5065), .C1(n5508), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U6469 ( .A(n5068), .ZN(n5069) );
  INV_X1 U6470 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5126) );
  INV_X1 U6471 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5071) );
  MUX2_X1 U6472 ( .A(n5126), .B(n5071), .S(n4276), .Z(n5073) );
  INV_X1 U6473 ( .A(SI_12_), .ZN(n5072) );
  NAND2_X1 U6474 ( .A1(n5073), .A2(n5072), .ZN(n5159) );
  INV_X1 U6475 ( .A(n5073), .ZN(n5074) );
  NAND2_X1 U6476 ( .A1(n5074), .A2(SI_12_), .ZN(n5075) );
  NAND2_X1 U6477 ( .A1(n5159), .A2(n5075), .ZN(n5160) );
  XNOR2_X1 U6478 ( .A(n5161), .B(n5160), .ZN(n6733) );
  INV_X1 U6479 ( .A(n6733), .ZN(n5125) );
  NAND2_X1 U6480 ( .A1(n5076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5077) );
  XNOR2_X1 U6481 ( .A(n5077), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9493) );
  AOI22_X1 U6482 ( .A1(n9493), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n5848), .ZN(n5078) );
  OAI21_X1 U6483 ( .B1(n5125), .B2(n8059), .A(n5078), .ZN(P1_U3341) );
  INV_X1 U6484 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9768) );
  INV_X1 U6485 ( .A(n7122), .ZN(n5081) );
  XNOR2_X1 U6486 ( .A(n6925), .B(P2_B_REG_SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6487 ( .A1(n7063), .A2(n5079), .ZN(n5080) );
  AND2_X1 U6488 ( .A1(n7063), .A2(n7122), .ZN(n9770) );
  AOI21_X1 U6489 ( .B1(n9768), .B2(n9762), .A(n9770), .ZN(n5788) );
  NOR4_X1 U6490 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5090) );
  INV_X1 U6491 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9963) );
  INV_X1 U6492 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10003) );
  INV_X1 U6493 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9996) );
  INV_X1 U6494 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9983) );
  NAND4_X1 U6495 ( .A1(n9963), .A2(n10003), .A3(n9996), .A4(n9983), .ZN(n5087)
         );
  NOR4_X1 U6496 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5085) );
  NOR4_X1 U6497 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5084) );
  NOR4_X1 U6498 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5083) );
  NOR4_X1 U6499 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5082) );
  NAND4_X1 U6500 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), .ZN(n5086)
         );
  NOR4_X1 U6501 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5087), .A4(n5086), .ZN(n5089) );
  NOR4_X1 U6502 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5088) );
  NAND3_X1 U6503 ( .A1(n5090), .A2(n5089), .A3(n5088), .ZN(n5091) );
  NAND2_X1 U6504 ( .A1(n5091), .A2(n9762), .ZN(n5789) );
  INV_X1 U6505 ( .A(n9763), .ZN(n5821) );
  NAND2_X1 U6506 ( .A1(n6358), .A2(n8236), .ZN(n7755) );
  NAND2_X1 U6507 ( .A1(n5791), .A2(n7755), .ZN(n6096) );
  NAND3_X1 U6508 ( .A1(n6358), .A2(n8253), .A3(n5119), .ZN(n9814) );
  OR2_X1 U6509 ( .A1(n9814), .A2(n5118), .ZN(n6100) );
  NAND4_X1 U6510 ( .A1(n5789), .A2(n5821), .A3(n6096), .A4(n6100), .ZN(n5098)
         );
  OR2_X1 U6511 ( .A1(n5788), .A2(n5098), .ZN(n5585) );
  AND2_X1 U6512 ( .A1(n6925), .A2(n7122), .ZN(n9766) );
  INV_X1 U6513 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9765) );
  AND2_X1 U6514 ( .A1(n9762), .A2(n9765), .ZN(n5099) );
  NAND2_X1 U6515 ( .A1(n4279), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5102) );
  AND2_X1 U6516 ( .A1(n5103), .A2(n5102), .ZN(n5106) );
  NAND2_X1 U6517 ( .A1(n5609), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6518 ( .A1(n7320), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5104) );
  NAND3_X1 U6519 ( .A1(n5106), .A2(n5105), .A3(n5104), .ZN(n5110) );
  INV_X1 U6520 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U6521 ( .A1(n5587), .A2(SI_0_), .ZN(n5107) );
  XNOR2_X1 U6522 ( .A(n5107), .B(n5042), .ZN(n8546) );
  MUX2_X1 U6523 ( .A(n9745), .B(n8546), .S(n5602), .Z(n5970) );
  NAND2_X1 U6524 ( .A1(n5109), .A2(n5108), .ZN(n8411) );
  NAND2_X1 U6525 ( .A1(n5110), .A2(n5970), .ZN(n7716) );
  NAND2_X1 U6526 ( .A1(n8411), .A2(n7716), .ZN(n6269) );
  INV_X1 U6527 ( .A(n6358), .ZN(n7744) );
  NAND2_X1 U6528 ( .A1(n7744), .A2(n5118), .ZN(n7549) );
  NAND2_X1 U6529 ( .A1(n7549), .A2(n5740), .ZN(n8414) );
  NAND2_X1 U6530 ( .A1(n5609), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U6531 ( .A1(n4278), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6532 ( .A1(n4277), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5111) );
  INV_X1 U6533 ( .A(n5115), .ZN(n5615) );
  NAND2_X1 U6534 ( .A1(n5791), .A2(n5115), .ZN(n8330) );
  INV_X1 U6535 ( .A(n8330), .ZN(n8417) );
  AND2_X1 U6536 ( .A1(n5593), .A2(n8417), .ZN(n5116) );
  AOI21_X1 U6537 ( .B1(n6269), .B2(n8414), .A(n5116), .ZN(n6270) );
  NAND2_X1 U6538 ( .A1(n6358), .A2(n5118), .ZN(n6106) );
  XNOR2_X1 U6539 ( .A(n6106), .B(n7757), .ZN(n5117) );
  NAND2_X1 U6540 ( .A1(n5117), .A2(n8236), .ZN(n7181) );
  AND2_X1 U6541 ( .A1(n7181), .A2(n9814), .ZN(n9804) );
  INV_X1 U6542 ( .A(n9804), .ZN(n9823) );
  NAND2_X1 U6543 ( .A1(n9823), .A2(n6269), .ZN(n5121) );
  NAND2_X1 U6544 ( .A1(n5108), .A2(n5617), .ZN(n5120) );
  AND3_X1 U6545 ( .A1(n6270), .A2(n5121), .A3(n5120), .ZN(n9772) );
  NAND2_X1 U6546 ( .A1(n9833), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5122) );
  OAI21_X1 U6547 ( .B1(n9833), .B2(n9772), .A(n5122), .ZN(P2_U3520) );
  OR2_X1 U6548 ( .A1(n5123), .A2(n4853), .ZN(n5124) );
  XNOR2_X1 U6549 ( .A(n5124), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6734) );
  INV_X1 U6550 ( .A(n6734), .ZN(n5723) );
  OAI222_X1 U6551 ( .A1(n8545), .A2(n5126), .B1(n4270), .B2(n5125), .C1(
        P2_U3152), .C2(n5723), .ZN(P2_U3346) );
  NAND2_X1 U6552 ( .A1(n5132), .A2(n5129), .ZN(n5134) );
  NAND2_X1 U6553 ( .A1(n5133), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5135) );
  NAND2_X1 U6554 ( .A1(n5393), .A2(n8931), .ZN(n5477) );
  INV_X1 U6555 ( .A(n5651), .ZN(n6726) );
  OR2_X1 U6556 ( .A1(n5477), .A2(n6726), .ZN(n5136) );
  NAND2_X1 U6557 ( .A1(n5136), .A2(n5423), .ZN(n5192) );
  NAND2_X1 U6558 ( .A1(n5137), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6559 ( .A1(n4271), .A2(n5138), .ZN(n5142) );
  INV_X1 U6560 ( .A(n5142), .ZN(n5140) );
  NAND2_X1 U6561 ( .A1(n5140), .A2(n4811), .ZN(n5141) );
  NAND2_X2 U6562 ( .A1(n5144), .A2(n5146), .ZN(n5458) );
  OR2_X1 U6563 ( .A1(n5192), .A2(n7822), .ZN(n5154) );
  NAND2_X1 U6564 ( .A1(n5154), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U6565 ( .A(P1_U3083), .ZN(n5143) );
  NAND2_X1 U6566 ( .A1(n5143), .A2(n5423), .ZN(n9579) );
  INV_X1 U6567 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n5158) );
  OR2_X1 U6568 ( .A1(n5145), .A2(P1_U3084), .ZN(n9325) );
  OR2_X1 U6569 ( .A1(n5192), .A2(n9325), .ZN(n5170) );
  INV_X1 U6570 ( .A(n5170), .ZN(n5147) );
  NAND2_X1 U6571 ( .A1(n5147), .A2(n8055), .ZN(n9576) );
  INV_X1 U6572 ( .A(n9576), .ZN(n9557) );
  INV_X1 U6573 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9441) );
  NAND3_X1 U6574 ( .A1(n9557), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9441), .ZN(
        n5157) );
  NAND2_X1 U6575 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n5171) );
  INV_X1 U6576 ( .A(n5171), .ZN(n5148) );
  NOR2_X1 U6577 ( .A1(n8055), .A2(n5148), .ZN(n5149) );
  NOR2_X1 U6578 ( .A1(n5149), .A2(n5145), .ZN(n5421) );
  OAI21_X1 U6579 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9441), .A(n5421), .ZN(n5151) );
  NOR2_X1 U6580 ( .A1(n8055), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5150) );
  OAI22_X1 U6581 ( .A1(n9325), .A2(n5150), .B1(P1_U3084), .B2(n9440), .ZN(
        n5424) );
  NAND2_X1 U6582 ( .A1(n5151), .A2(n5424), .ZN(n5153) );
  INV_X1 U6583 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5152) );
  OAI22_X1 U6584 ( .A1(n5154), .A2(n5153), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5152), .ZN(n5155) );
  INV_X1 U6585 ( .A(n5155), .ZN(n5156) );
  OAI211_X1 U6586 ( .C1(n9579), .C2(n5158), .A(n5157), .B(n5156), .ZN(P1_U3241) );
  INV_X1 U6587 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5337) );
  INV_X1 U6588 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5162) );
  MUX2_X1 U6589 ( .A(n5337), .B(n5162), .S(n7537), .Z(n5164) );
  INV_X1 U6590 ( .A(SI_13_), .ZN(n5163) );
  NAND2_X1 U6591 ( .A1(n5164), .A2(n5163), .ZN(n5339) );
  INV_X1 U6592 ( .A(n5164), .ZN(n5165) );
  NAND2_X1 U6593 ( .A1(n5165), .A2(SI_13_), .ZN(n5166) );
  XNOR2_X1 U6594 ( .A(n5338), .B(n4814), .ZN(n6878) );
  INV_X1 U6595 ( .A(n6878), .ZN(n5336) );
  OR2_X1 U6596 ( .A1(n5167), .A2(n4915), .ZN(n5168) );
  XNOR2_X1 U6597 ( .A(n5168), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9506) );
  AOI22_X1 U6598 ( .A1(n9506), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n5848), .ZN(n5169) );
  OAI21_X1 U6599 ( .B1(n5336), .B2(n8059), .A(n5169), .ZN(P1_U3340) );
  INV_X1 U6600 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n5198) );
  NOR2_X1 U6601 ( .A1(n5170), .A2(n8055), .ZN(n9454) );
  INV_X1 U6602 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U6603 ( .A1(n5885), .A2(n6420), .ZN(n5175) );
  INV_X1 U6604 ( .A(n5175), .ZN(n5176) );
  INV_X1 U6605 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5174) );
  INV_X1 U6606 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5433) );
  INV_X1 U6607 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5990) );
  MUX2_X1 U6608 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n5990), .S(n9430), .Z(n9434)
         );
  NOR2_X1 U6609 ( .A1(n9434), .A2(n5171), .ZN(n9433) );
  NOR2_X1 U6610 ( .A1(n9430), .A2(n5990), .ZN(n5434) );
  MUX2_X1 U6611 ( .A(n5433), .B(P1_REG2_REG_2__SCAN_IN), .S(n5675), .Z(n5172)
         );
  OAI21_X1 U6612 ( .B1(n9433), .B2(n5434), .A(n5172), .ZN(n5437) );
  OAI21_X1 U6613 ( .B1(n5433), .B2(n5675), .A(n5437), .ZN(n9338) );
  MUX2_X1 U6614 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n5174), .S(n9330), .Z(n5173)
         );
  INV_X1 U6615 ( .A(n5173), .ZN(n9337) );
  NAND2_X1 U6616 ( .A1(n9338), .A2(n9337), .ZN(n9336) );
  OAI21_X1 U6617 ( .B1(n9330), .B2(n5174), .A(n9336), .ZN(n5561) );
  OAI21_X1 U6618 ( .B1(n5885), .B2(n6420), .A(n5175), .ZN(n5560) );
  NOR2_X1 U6619 ( .A1(n5561), .A2(n5560), .ZN(n5559) );
  NOR2_X1 U6620 ( .A1(n5176), .A2(n5559), .ZN(n5446) );
  INV_X1 U6621 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9597) );
  NAND2_X1 U6622 ( .A1(n6038), .A2(n9597), .ZN(n5177) );
  OAI21_X1 U6623 ( .B1(n6038), .B2(n9597), .A(n5177), .ZN(n5445) );
  NOR2_X1 U6624 ( .A1(n5446), .A2(n5445), .ZN(n5444) );
  INV_X1 U6625 ( .A(n5177), .ZN(n5178) );
  NOR2_X1 U6626 ( .A1(n5444), .A2(n5178), .ZN(n5296) );
  INV_X1 U6627 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5179) );
  MUX2_X1 U6628 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n5179), .S(n6044), .Z(n5294)
         );
  XNOR2_X1 U6629 ( .A(n5296), .B(n5294), .ZN(n5196) );
  INV_X1 U6630 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5180) );
  MUX2_X1 U6631 ( .A(n5180), .B(P1_REG1_REG_5__SCAN_IN), .S(n6038), .Z(n5184)
         );
  INV_X1 U6632 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5183) );
  MUX2_X1 U6633 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n5183), .S(n5885), .Z(n5556)
         );
  INV_X1 U6634 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5182) );
  INV_X1 U6635 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9688) );
  INV_X1 U6636 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5487) );
  NOR2_X1 U6637 ( .A1(n9430), .A2(n5487), .ZN(n5427) );
  MUX2_X1 U6638 ( .A(n9688), .B(P1_REG1_REG_2__SCAN_IN), .S(n5675), .Z(n5181)
         );
  OAI21_X1 U6639 ( .B1(n9438), .B2(n5427), .A(n5181), .ZN(n5430) );
  OAI21_X1 U6640 ( .B1(n9688), .B2(n5675), .A(n5430), .ZN(n9335) );
  MUX2_X1 U6641 ( .A(n5182), .B(P1_REG1_REG_3__SCAN_IN), .S(n9330), .Z(n9334)
         );
  NAND2_X1 U6642 ( .A1(n9335), .A2(n9334), .ZN(n9333) );
  OAI21_X1 U6643 ( .B1(n9330), .B2(n5182), .A(n9333), .ZN(n5557) );
  INV_X1 U6644 ( .A(n6038), .ZN(n5453) );
  NAND2_X1 U6645 ( .A1(n5453), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5185) );
  INV_X1 U6646 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5186) );
  AND2_X1 U6647 ( .A1(n6044), .A2(n5186), .ZN(n5284) );
  NOR2_X1 U6648 ( .A1(n6044), .A2(n5186), .ZN(n5187) );
  OR2_X1 U6649 ( .A1(n5284), .A2(n5187), .ZN(n5188) );
  NOR2_X1 U6650 ( .A1(n5189), .A2(n5188), .ZN(n5283) );
  AOI21_X1 U6651 ( .B1(n5189), .B2(n5188), .A(n5283), .ZN(n5194) );
  NOR2_X1 U6652 ( .A1(n8055), .A2(P1_U3084), .ZN(n5190) );
  NAND2_X1 U6653 ( .A1(n5190), .A2(n5145), .ZN(n5191) );
  OR2_X1 U6654 ( .A1(n5192), .A2(n5191), .ZN(n9452) );
  INV_X1 U6655 ( .A(n9452), .ZN(n9570) );
  INV_X1 U6656 ( .A(n6044), .ZN(n5293) );
  INV_X1 U6657 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6046) );
  NOR2_X1 U6658 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6046), .ZN(n6283) );
  AOI21_X1 U6659 ( .B1(n9570), .B2(n5293), .A(n6283), .ZN(n5193) );
  OAI21_X1 U6660 ( .B1(n9576), .B2(n5194), .A(n5193), .ZN(n5195) );
  AOI21_X1 U6661 ( .B1(n9454), .B2(n5196), .A(n5195), .ZN(n5197) );
  OAI21_X1 U6662 ( .B1(n9579), .B2(n5198), .A(n5197), .ZN(P1_U3247) );
  INV_X2 U6663 ( .A(P2_U3966), .ZN(n8160) );
  NAND2_X1 U6664 ( .A1(n5199), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5200) );
  OAI211_X1 U6665 ( .C1(n9763), .C2(n5791), .A(n7760), .B(n5200), .ZN(n5201)
         );
  NAND2_X1 U6666 ( .A1(n5201), .A2(n5602), .ZN(n5220) );
  NAND2_X1 U6667 ( .A1(n8160), .A2(n5220), .ZN(n5243) );
  AND2_X1 U6668 ( .A1(n5243), .A2(n5115), .ZN(n9757) );
  INV_X1 U6669 ( .A(n9747), .ZN(n6298) );
  INV_X1 U6670 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6671 ( .A1(n6224), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5218) );
  INV_X1 U6672 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5202) );
  MUX2_X1 U6673 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n5202), .S(n6224), .Z(n5250)
         );
  NAND2_X1 U6674 ( .A1(n9756), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5217) );
  INV_X1 U6675 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5203) );
  MUX2_X1 U6676 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n5203), .S(n9756), .Z(n9754)
         );
  NAND2_X1 U6677 ( .A1(n5909), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5216) );
  INV_X1 U6678 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5204) );
  MUX2_X1 U6679 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n5204), .S(n5909), .Z(n5261)
         );
  NAND2_X1 U6680 ( .A1(n5529), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5215) );
  INV_X1 U6681 ( .A(n5771), .ZN(n5213) );
  INV_X1 U6682 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5205) );
  MUX2_X1 U6683 ( .A(n5205), .B(P2_REG1_REG_1__SCAN_IN), .S(n5589), .Z(n5310)
         );
  AND2_X1 U6684 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n5206) );
  NAND2_X1 U6685 ( .A1(n5310), .A2(n5206), .ZN(n5345) );
  INV_X1 U6686 ( .A(n5589), .ZN(n5316) );
  NAND2_X1 U6687 ( .A1(n5316), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6688 ( .A1(n5345), .A2(n5344), .ZN(n5209) );
  INV_X1 U6689 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5207) );
  MUX2_X1 U6690 ( .A(n5207), .B(P2_REG1_REG_2__SCAN_IN), .S(n5601), .Z(n5208)
         );
  AND2_X1 U6691 ( .A1(n5209), .A2(n5208), .ZN(n5497) );
  NOR2_X1 U6692 ( .A1(n5601), .A2(n5207), .ZN(n5492) );
  INV_X1 U6693 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5210) );
  MUX2_X1 U6694 ( .A(n5210), .B(P2_REG1_REG_3__SCAN_IN), .S(n5759), .Z(n5211)
         );
  OAI21_X1 U6695 ( .B1(n5497), .B2(n5492), .A(n5211), .ZN(n5495) );
  INV_X1 U6696 ( .A(n5759), .ZN(n5212) );
  NAND2_X1 U6697 ( .A1(n5212), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5272) );
  INV_X1 U6698 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5867) );
  MUX2_X1 U6699 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5867), .S(n5771), .Z(n5271)
         );
  AOI21_X1 U6700 ( .B1(n5495), .B2(n5272), .A(n5271), .ZN(n5274) );
  AOI21_X1 U6701 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n5213), .A(n5274), .ZN(
        n5519) );
  INV_X1 U6702 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9828) );
  MUX2_X1 U6703 ( .A(n9828), .B(P2_REG1_REG_5__SCAN_IN), .S(n5529), .Z(n5214)
         );
  OR2_X1 U6704 ( .A1(n5519), .A2(n5214), .ZN(n5522) );
  NAND2_X1 U6705 ( .A1(n5215), .A2(n5522), .ZN(n5262) );
  NAND2_X1 U6706 ( .A1(n5261), .A2(n5262), .ZN(n5260) );
  NAND2_X1 U6707 ( .A1(n5216), .A2(n5260), .ZN(n9755) );
  NAND2_X1 U6708 ( .A1(n9754), .A2(n9755), .ZN(n9752) );
  NAND2_X1 U6709 ( .A1(n5217), .A2(n9752), .ZN(n5251) );
  NAND2_X1 U6710 ( .A1(n5250), .A2(n5251), .ZN(n5249) );
  NAND2_X1 U6711 ( .A1(n5218), .A2(n5249), .ZN(n5223) );
  INV_X1 U6712 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5219) );
  MUX2_X1 U6713 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n5219), .S(n6322), .Z(n5222)
         );
  INV_X1 U6714 ( .A(n5220), .ZN(n5221) );
  AND2_X1 U6715 ( .A1(n5221), .A2(n7756), .ZN(n9753) );
  NAND2_X1 U6716 ( .A1(n5222), .A2(n5223), .ZN(n5321) );
  OAI211_X1 U6717 ( .C1(n5223), .C2(n5222), .A(n9753), .B(n5321), .ZN(n5224)
         );
  NAND2_X1 U6718 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6337) );
  OAI211_X1 U6719 ( .C1(n6298), .C2(n5225), .A(n5224), .B(n6337), .ZN(n5226)
         );
  AOI21_X1 U6720 ( .B1(n6322), .B2(n9757), .A(n5226), .ZN(n5248) );
  NAND2_X1 U6721 ( .A1(n6224), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5240) );
  INV_X1 U6722 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5227) );
  MUX2_X1 U6723 ( .A(n5227), .B(P2_REG2_REG_8__SCAN_IN), .S(n6224), .Z(n5228)
         );
  INV_X1 U6724 ( .A(n5228), .ZN(n5256) );
  NAND2_X1 U6725 ( .A1(n9756), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5239) );
  INV_X1 U6726 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5229) );
  MUX2_X1 U6727 ( .A(n5229), .B(P2_REG2_REG_7__SCAN_IN), .S(n9756), .Z(n5230)
         );
  INV_X1 U6728 ( .A(n5230), .ZN(n9750) );
  NAND2_X1 U6729 ( .A1(n5909), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5238) );
  INV_X1 U6730 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5231) );
  MUX2_X1 U6731 ( .A(n5231), .B(P2_REG2_REG_6__SCAN_IN), .S(n5909), .Z(n5232)
         );
  INV_X1 U6732 ( .A(n5232), .ZN(n5267) );
  NAND2_X1 U6733 ( .A1(n5529), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5237) );
  INV_X1 U6734 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5234) );
  XNOR2_X1 U6735 ( .A(n5601), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n5343) );
  XNOR2_X1 U6736 ( .A(n5589), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n5313) );
  AND2_X1 U6737 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n5312) );
  NAND2_X1 U6738 ( .A1(n5313), .A2(n5312), .ZN(n5311) );
  NAND2_X1 U6739 ( .A1(n5316), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6740 ( .A1(n5311), .A2(n5233), .ZN(n5342) );
  INV_X1 U6741 ( .A(n5601), .ZN(n5352) );
  AOI22_X1 U6742 ( .A1(n5343), .A2(n5342), .B1(n5352), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n5491) );
  INV_X1 U6743 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6442) );
  MUX2_X1 U6744 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6442), .S(n5759), .Z(n5490)
         );
  NOR2_X1 U6745 ( .A1(n5491), .A2(n5490), .ZN(n5489) );
  NOR2_X1 U6746 ( .A1(n5759), .A2(n6442), .ZN(n5278) );
  MUX2_X1 U6747 ( .A(n5234), .B(P2_REG2_REG_4__SCAN_IN), .S(n5771), .Z(n5277)
         );
  OAI21_X1 U6748 ( .B1(n5489), .B2(n5278), .A(n5277), .ZN(n5280) );
  OAI21_X1 U6749 ( .B1(n5234), .B2(n5771), .A(n5280), .ZN(n5531) );
  INV_X1 U6750 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5235) );
  MUX2_X1 U6751 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n5235), .S(n5529), .Z(n5236)
         );
  NAND2_X1 U6752 ( .A1(n5531), .A2(n5236), .ZN(n5530) );
  NAND2_X1 U6753 ( .A1(n5237), .A2(n5530), .ZN(n5268) );
  NAND2_X1 U6754 ( .A1(n5267), .A2(n5268), .ZN(n5266) );
  NAND2_X1 U6755 ( .A1(n5238), .A2(n5266), .ZN(n9751) );
  NAND2_X1 U6756 ( .A1(n9750), .A2(n9751), .ZN(n9748) );
  NAND2_X1 U6757 ( .A1(n5239), .A2(n9748), .ZN(n5257) );
  NAND2_X1 U6758 ( .A1(n5256), .A2(n5257), .ZN(n5255) );
  NAND2_X1 U6759 ( .A1(n5240), .A2(n5255), .ZN(n5246) );
  INV_X1 U6760 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5241) );
  MUX2_X1 U6761 ( .A(n5241), .B(P2_REG2_REG_9__SCAN_IN), .S(n6322), .Z(n5242)
         );
  INV_X1 U6762 ( .A(n5242), .ZN(n5245) );
  INV_X1 U6763 ( .A(n7756), .ZN(n7791) );
  NAND2_X1 U6764 ( .A1(n5243), .A2(n7791), .ZN(n8171) );
  INV_X1 U6765 ( .A(n8171), .ZN(n5244) );
  NAND2_X1 U6766 ( .A1(n5245), .A2(n5246), .ZN(n5327) );
  OAI211_X1 U6767 ( .C1(n5246), .C2(n5245), .A(n9749), .B(n5327), .ZN(n5247)
         );
  NAND2_X1 U6768 ( .A1(n5248), .A2(n5247), .ZN(P2_U3254) );
  INV_X1 U6769 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n5253) );
  OAI211_X1 U6770 ( .C1(n5251), .C2(n5250), .A(n9753), .B(n5249), .ZN(n5252)
         );
  NAND2_X1 U6771 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n9712) );
  OAI211_X1 U6772 ( .C1(n6298), .C2(n5253), .A(n5252), .B(n9712), .ZN(n5254)
         );
  AOI21_X1 U6773 ( .B1(n6224), .B2(n9757), .A(n5254), .ZN(n5259) );
  OAI211_X1 U6774 ( .C1(n5257), .C2(n5256), .A(n9749), .B(n5255), .ZN(n5258)
         );
  NAND2_X1 U6775 ( .A1(n5259), .A2(n5258), .ZN(P2_U3253) );
  INV_X1 U6776 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n5264) );
  OAI211_X1 U6777 ( .C1(n5262), .C2(n5261), .A(n9753), .B(n5260), .ZN(n5263)
         );
  NAND2_X1 U6778 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n5944) );
  OAI211_X1 U6779 ( .C1(n6298), .C2(n5264), .A(n5263), .B(n5944), .ZN(n5265)
         );
  AOI21_X1 U6780 ( .B1(n5909), .B2(n9757), .A(n5265), .ZN(n5270) );
  OAI211_X1 U6781 ( .C1(n5268), .C2(n5267), .A(n9749), .B(n5266), .ZN(n5269)
         );
  NAND2_X1 U6782 ( .A1(n5270), .A2(n5269), .ZN(P2_U3251) );
  INV_X1 U6783 ( .A(n9757), .ZN(n9739) );
  NAND2_X1 U6784 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n5801) );
  INV_X1 U6785 ( .A(n5801), .ZN(n5276) );
  INV_X1 U6786 ( .A(n9753), .ZN(n9740) );
  AND3_X1 U6787 ( .A1(n5495), .A2(n5272), .A3(n5271), .ZN(n5273) );
  NOR3_X1 U6788 ( .A1(n9740), .A2(n5274), .A3(n5273), .ZN(n5275) );
  AOI211_X1 U6789 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9747), .A(n5276), .B(
        n5275), .ZN(n5282) );
  OR3_X1 U6790 ( .A1(n5489), .A2(n5278), .A3(n5277), .ZN(n5279) );
  NAND3_X1 U6791 ( .A1(n9749), .A2(n5280), .A3(n5279), .ZN(n5281) );
  OAI211_X1 U6792 ( .C1(n9739), .C2(n5771), .A(n5282), .B(n5281), .ZN(P2_U3249) );
  NOR2_X1 U6793 ( .A1(n9467), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5288) );
  INV_X1 U6794 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5286) );
  NOR2_X1 U6795 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n5544), .ZN(n5285) );
  INV_X1 U6796 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9694) );
  AOI22_X1 U6797 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6054), .B1(n5544), .B2(
        n9694), .ZN(n5546) );
  MUX2_X1 U6798 ( .A(n5286), .B(P1_REG1_REG_8__SCAN_IN), .S(n9451), .Z(n9457)
         );
  OAI21_X1 U6799 ( .B1(n9451), .B2(n5286), .A(n9456), .ZN(n9470) );
  INV_X1 U6800 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5287) );
  MUX2_X1 U6801 ( .A(n5287), .B(P1_REG1_REG_9__SCAN_IN), .S(n9467), .Z(n9469)
         );
  NOR2_X1 U6802 ( .A1(n9470), .A2(n9469), .ZN(n9468) );
  NOR2_X1 U6803 ( .A1(n5288), .A2(n9468), .ZN(n9483) );
  INV_X1 U6804 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5289) );
  MUX2_X1 U6805 ( .A(n5289), .B(P1_REG1_REG_10__SCAN_IN), .S(n9479), .Z(n9482)
         );
  OR2_X1 U6806 ( .A1(n9479), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5290) );
  INV_X1 U6807 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9414) );
  AOI22_X1 U6808 ( .A1(n8970), .A2(n9414), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n8957), .ZN(n5291) );
  AOI21_X1 U6809 ( .B1(n5292), .B2(n5291), .A(n8956), .ZN(n5309) );
  NOR2_X1 U6810 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n5544), .ZN(n5298) );
  INV_X1 U6811 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6078) );
  AOI22_X1 U6812 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6054), .B1(n5544), .B2(
        n6078), .ZN(n5543) );
  NAND2_X1 U6813 ( .A1(n5293), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5297) );
  INV_X1 U6814 ( .A(n5294), .ZN(n5295) );
  AND2_X1 U6815 ( .A1(n9449), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5299) );
  INV_X1 U6816 ( .A(n9451), .ZN(n9447) );
  OAI22_X1 U6817 ( .A1(n5299), .A2(n9447), .B1(n9449), .B2(
        P1_REG2_REG_8__SCAN_IN), .ZN(n9464) );
  OR2_X1 U6818 ( .A1(n9467), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6819 ( .A1(n9467), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6820 ( .A1(n5301), .A2(n5300), .ZN(n9463) );
  NOR2_X1 U6821 ( .A1(n9464), .A2(n9463), .ZN(n9462) );
  AOI21_X1 U6822 ( .B1(n9467), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9462), .ZN(
        n9476) );
  XNOR2_X1 U6823 ( .A(n9479), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9475) );
  NOR2_X1 U6824 ( .A1(n8970), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5302) );
  AOI21_X1 U6825 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n8970), .A(n5302), .ZN(
        n5303) );
  OAI21_X1 U6826 ( .B1(n5304), .B2(n5303), .A(n8969), .ZN(n5305) );
  NAND2_X1 U6827 ( .A1(n5305), .A2(n9454), .ZN(n5308) );
  INV_X1 U6828 ( .A(n9579), .ZN(n9432) );
  AND2_X1 U6829 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6823) );
  NOR2_X1 U6830 ( .A1(n9452), .A2(n8957), .ZN(n5306) );
  AOI211_X1 U6831 ( .C1(n9432), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n6823), .B(
        n5306), .ZN(n5307) );
  OAI211_X1 U6832 ( .C1(n5309), .C2(n9576), .A(n5308), .B(n5307), .ZN(P1_U3252) );
  AND2_X1 U6833 ( .A1(n9753), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9738) );
  AOI22_X1 U6834 ( .A1(n9738), .A2(P2_IR_REG_0__SCAN_IN), .B1(n9753), .B2(
        n5310), .ZN(n5320) );
  INV_X1 U6835 ( .A(n5345), .ZN(n5319) );
  OAI211_X1 U6836 ( .C1(n5313), .C2(n5312), .A(n9749), .B(n5311), .ZN(n5318)
         );
  INV_X1 U6837 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n5314) );
  INV_X1 U6838 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5823) );
  OAI22_X1 U6839 ( .A1(n6298), .A2(n5314), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5823), .ZN(n5315) );
  AOI21_X1 U6840 ( .B1(n9757), .B2(n5316), .A(n5315), .ZN(n5317) );
  OAI211_X1 U6841 ( .C1(n5320), .C2(n5319), .A(n5318), .B(n5317), .ZN(P2_U3246) );
  NAND2_X1 U6842 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n9701) );
  INV_X1 U6843 ( .A(n9701), .ZN(n5326) );
  INV_X1 U6844 ( .A(n5321), .ZN(n5322) );
  AOI21_X1 U6845 ( .B1(n6322), .B2(P2_REG1_REG_9__SCAN_IN), .A(n5322), .ZN(
        n5324) );
  INV_X1 U6846 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6921) );
  MUX2_X1 U6847 ( .A(n6921), .B(P2_REG1_REG_10__SCAN_IN), .S(n6475), .Z(n5323)
         );
  NOR2_X1 U6848 ( .A1(n5323), .A2(n5324), .ZN(n5406) );
  AOI211_X1 U6849 ( .C1(n5324), .C2(n5323), .A(n5406), .B(n9740), .ZN(n5325)
         );
  AOI211_X1 U6850 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9747), .A(n5326), .B(
        n5325), .ZN(n5333) );
  NAND2_X1 U6851 ( .A1(n6322), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6852 ( .A1(n5328), .A2(n5327), .ZN(n5331) );
  INV_X1 U6853 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5329) );
  MUX2_X1 U6854 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n5329), .S(n6475), .Z(n5330)
         );
  NAND2_X1 U6855 ( .A1(n6475), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5402) );
  OAI211_X1 U6856 ( .C1(n6475), .C2(P2_REG2_REG_10__SCAN_IN), .A(n5331), .B(
        n5402), .ZN(n5401) );
  OAI211_X1 U6857 ( .C1(n5331), .C2(n5330), .A(n9749), .B(n5401), .ZN(n5332)
         );
  OAI211_X1 U6858 ( .C1(n9739), .C2(n5334), .A(n5333), .B(n5332), .ZN(P2_U3255) );
  OR2_X1 U6859 ( .A1(n5335), .A2(n4853), .ZN(n5414) );
  XNOR2_X1 U6860 ( .A(n5414), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6833) );
  INV_X1 U6861 ( .A(n6833), .ZN(n5880) );
  OAI222_X1 U6862 ( .A1(n8545), .A2(n5337), .B1(n4270), .B2(n5336), .C1(n5880), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U6863 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5420) );
  INV_X1 U6864 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5341) );
  MUX2_X1 U6865 ( .A(n5420), .B(n5341), .S(n4276), .Z(n5570) );
  XNOR2_X1 U6866 ( .A(n5570), .B(SI_14_), .ZN(n5569) );
  XNOR2_X1 U6867 ( .A(n5574), .B(n5569), .ZN(n7009) );
  INV_X1 U6868 ( .A(n7009), .ZN(n5419) );
  OR2_X1 U6869 ( .A1(n5340), .A2(n4915), .ZN(n5580) );
  XNOR2_X1 U6870 ( .A(n5580), .B(n5579), .ZN(n8973) );
  OAI222_X1 U6871 ( .A1(n8059), .A2(n5419), .B1(n8973), .B2(P1_U3084), .C1(
        n5341), .C2(n9328), .ZN(P1_U3339) );
  INV_X1 U6872 ( .A(n9749), .ZN(n6466) );
  XNOR2_X1 U6873 ( .A(n5343), .B(n5342), .ZN(n5354) );
  INV_X1 U6874 ( .A(n5497), .ZN(n5348) );
  MUX2_X1 U6875 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5207), .S(n5601), .Z(n5346)
         );
  NAND3_X1 U6876 ( .A1(n5346), .A2(n5345), .A3(n5344), .ZN(n5347) );
  NAND3_X1 U6877 ( .A1(n9753), .A2(n5348), .A3(n5347), .ZN(n5350) );
  AOI22_X1 U6878 ( .A1(n9747), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n5349) );
  NAND2_X1 U6879 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  AOI21_X1 U6880 ( .B1(n5352), .B2(n9757), .A(n5351), .ZN(n5353) );
  OAI21_X1 U6881 ( .B1(n6466), .B2(n5354), .A(n5353), .ZN(P2_U3247) );
  NOR2_X1 U6882 ( .A1(n5652), .A2(n9441), .ZN(n5358) );
  AOI21_X1 U6883 ( .B1(n5676), .B2(n5463), .A(n5358), .ZN(n5366) );
  INV_X1 U6884 ( .A(SI_0_), .ZN(n5361) );
  INV_X1 U6885 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5360) );
  OAI21_X1 U6886 ( .B1(n5587), .B2(n5361), .A(n5360), .ZN(n5363) );
  AND2_X1 U6887 ( .A1(n5363), .A2(n5362), .ZN(n9329) );
  BUF_X1 U6888 ( .A(n5458), .Z(n5364) );
  MUX2_X1 U6889 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9329), .S(n5364), .Z(n5984) );
  NAND2_X1 U6890 ( .A1(n6561), .A2(n5984), .ZN(n5365) );
  AND2_X1 U6891 ( .A1(n5366), .A2(n5365), .ZN(n5659) );
  NAND2_X1 U6892 ( .A1(n5367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5368) );
  AND2_X4 U6893 ( .A1(n4810), .A2(n6561), .ZN(n7974) );
  NOR2_X1 U6894 ( .A1(n5652), .A2(n9440), .ZN(n5369) );
  AOI21_X1 U6895 ( .B1(n5676), .B2(n5984), .A(n5369), .ZN(n5370) );
  NAND2_X1 U6896 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  AOI21_X1 U6897 ( .B1(n5659), .B2(n5372), .A(n4751), .ZN(n5422) );
  NOR4_X1 U6898 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5376) );
  NOR4_X1 U6899 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5375) );
  NOR4_X1 U6900 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5374) );
  NOR4_X1 U6901 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5373) );
  NAND4_X1 U6902 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), .ZN(n5382)
         );
  NOR2_X1 U6903 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .ZN(
        n5380) );
  NOR4_X1 U6904 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5379) );
  NOR4_X1 U6905 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5378) );
  NOR4_X1 U6906 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5377) );
  NAND4_X1 U6907 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), .ZN(n5381)
         );
  OAI21_X1 U6908 ( .B1(n5382), .B2(n5381), .A(n9624), .ZN(n5484) );
  INV_X1 U6909 ( .A(n5484), .ZN(n5383) );
  OR2_X1 U6910 ( .A1(n5383), .A2(n5485), .ZN(n5976) );
  INV_X1 U6911 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U6912 ( .A1(n9624), .A2(n9631), .ZN(n5385) );
  NAND2_X1 U6913 ( .A1(n7124), .A2(n6988), .ZN(n5384) );
  NAND2_X1 U6914 ( .A1(n5385), .A2(n5384), .ZN(n5977) );
  NOR2_X1 U6915 ( .A1(n5976), .A2(n5977), .ZN(n5389) );
  AND2_X1 U6916 ( .A1(n5389), .A2(n9630), .ZN(n5394) );
  INV_X1 U6917 ( .A(n8931), .ZN(n6522) );
  NAND2_X1 U6918 ( .A1(n8886), .A2(n6522), .ZN(n5982) );
  INV_X1 U6919 ( .A(n5982), .ZN(n5536) );
  INV_X1 U6920 ( .A(n5466), .ZN(n5981) );
  INV_X1 U6921 ( .A(n5477), .ZN(n8923) );
  NOR2_X1 U6922 ( .A1(n9632), .A2(n8923), .ZN(n5387) );
  NAND2_X1 U6923 ( .A1(n5394), .A2(n5387), .ZN(n8650) );
  INV_X1 U6924 ( .A(n5389), .ZN(n5388) );
  NAND3_X1 U6925 ( .A1(n4349), .A2(n5388), .A3(n9630), .ZN(n5657) );
  OR2_X1 U6926 ( .A1(n5389), .A2(n9632), .ZN(n5654) );
  OR2_X1 U6927 ( .A1(n5477), .A2(n5466), .ZN(n5653) );
  NAND2_X1 U6928 ( .A1(n5653), .A2(n9630), .ZN(n5979) );
  INV_X1 U6929 ( .A(n5979), .ZN(n5390) );
  NAND3_X1 U6930 ( .A1(n5657), .A2(n5654), .A3(n5390), .ZN(n8580) );
  NAND2_X1 U6931 ( .A1(n5394), .A2(n4349), .ZN(n5392) );
  NAND2_X1 U6932 ( .A1(n6522), .A2(n9630), .ZN(n5391) );
  NAND2_X1 U6933 ( .A1(n5392), .A2(n9618), .ZN(n8648) );
  INV_X1 U6934 ( .A(n5984), .ZN(n5540) );
  NAND2_X1 U6935 ( .A1(n5393), .A2(n9128), .ZN(n5660) );
  OR2_X1 U6936 ( .A1(n5359), .A2(n5660), .ZN(n5989) );
  INV_X1 U6937 ( .A(n5989), .ZN(n8935) );
  NAND2_X1 U6938 ( .A1(n5394), .A2(n8935), .ZN(n5718) );
  INV_X1 U6939 ( .A(n5145), .ZN(n8934) );
  OR2_X1 U6940 ( .A1(n5718), .A2(n8934), .ZN(n8657) );
  NAND2_X1 U6941 ( .A1(n4280), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6942 ( .A1(n5471), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6943 ( .A1(n5472), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5395) );
  INV_X1 U6944 ( .A(n5462), .ZN(n8681) );
  OAI22_X1 U6945 ( .A1(n8663), .A2(n5540), .B1(n8657), .B2(n8681), .ZN(n5399)
         );
  AOI21_X1 U6946 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n8580), .A(n5399), .ZN(
        n5400) );
  OAI21_X1 U6947 ( .B1(n5422), .B2(n8650), .A(n5400), .ZN(P1_U3230) );
  NAND2_X1 U6948 ( .A1(n5402), .A2(n5401), .ZN(n5405) );
  INV_X1 U6949 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5403) );
  AOI22_X1 U6950 ( .A1(n6482), .A2(n5403), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n5508), .ZN(n5404) );
  NOR2_X1 U6951 ( .A1(n5405), .A2(n5404), .ZN(n5502) );
  AOI21_X1 U6952 ( .B1(n5405), .B2(n5404), .A(n5502), .ZN(n5412) );
  AOI21_X1 U6953 ( .B1(n6475), .B2(P2_REG1_REG_10__SCAN_IN), .A(n5406), .ZN(
        n5506) );
  INV_X1 U6954 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9952) );
  MUX2_X1 U6955 ( .A(n9952), .B(P2_REG1_REG_11__SCAN_IN), .S(n6482), .Z(n5505)
         );
  XNOR2_X1 U6956 ( .A(n5506), .B(n5505), .ZN(n5409) );
  INV_X1 U6957 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6493) );
  NOR2_X1 U6958 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6493), .ZN(n5407) );
  AOI21_X1 U6959 ( .B1(n9747), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n5407), .ZN(
        n5408) );
  OAI21_X1 U6960 ( .B1(n9740), .B2(n5409), .A(n5408), .ZN(n5410) );
  AOI21_X1 U6961 ( .B1(n6482), .B2(n9757), .A(n5410), .ZN(n5411) );
  OAI21_X1 U6962 ( .B1(n5412), .B2(n6466), .A(n5411), .ZN(P2_U3256) );
  NAND2_X1 U6963 ( .A1(n5414), .A2(n5413), .ZN(n5415) );
  NAND2_X1 U6964 ( .A1(n5415), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5417) );
  OR2_X1 U6965 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  NAND2_X1 U6966 ( .A1(n5417), .A2(n5416), .ZN(n5647) );
  AND2_X1 U6967 ( .A1(n5418), .A2(n5647), .ZN(n7010) );
  INV_X1 U6968 ( .A(n7010), .ZN(n6013) );
  OAI222_X1 U6969 ( .A1(n8545), .A2(n5420), .B1(n4270), .B2(n5419), .C1(n6013), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U6970 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n5443) );
  INV_X1 U6971 ( .A(n8055), .ZN(n8989) );
  OAI21_X1 U6972 ( .B1(n5422), .B2(n8989), .A(n5421), .ZN(n5426) );
  INV_X1 U6973 ( .A(n5423), .ZN(n5425) );
  NAND3_X1 U6974 ( .A1(n5426), .A2(n5425), .A3(n5424), .ZN(n5567) );
  MUX2_X1 U6975 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9688), .S(n5675), .Z(n5429)
         );
  INV_X1 U6976 ( .A(n5427), .ZN(n5428) );
  NAND2_X1 U6977 ( .A1(n5429), .A2(n5428), .ZN(n5431) );
  OAI211_X1 U6978 ( .C1(n9438), .C2(n5431), .A(n9557), .B(n5430), .ZN(n5441)
         );
  INV_X1 U6979 ( .A(n5675), .ZN(n5432) );
  AOI22_X1 U6980 ( .A1(n9570), .A2(n5432), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n5440) );
  MUX2_X1 U6981 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n5433), .S(n5675), .Z(n5436)
         );
  INV_X1 U6982 ( .A(n5434), .ZN(n5435) );
  NAND2_X1 U6983 ( .A1(n5436), .A2(n5435), .ZN(n5438) );
  OAI211_X1 U6984 ( .C1(n9433), .C2(n5438), .A(n9454), .B(n5437), .ZN(n5439)
         );
  AND3_X1 U6985 ( .A1(n5441), .A2(n5440), .A3(n5439), .ZN(n5442) );
  OAI211_X1 U6986 ( .C1(n9579), .C2(n5443), .A(n5567), .B(n5442), .ZN(P1_U3243) );
  AOI21_X1 U6987 ( .B1(n5446), .B2(n5445), .A(n5444), .ZN(n5456) );
  AND2_X1 U6988 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6257) );
  INV_X1 U6989 ( .A(n5447), .ZN(n5451) );
  MUX2_X1 U6990 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5180), .S(n6038), .Z(n5450)
         );
  INV_X1 U6991 ( .A(n5448), .ZN(n5449) );
  AOI211_X1 U6992 ( .C1(n5451), .C2(n5450), .A(n5449), .B(n9576), .ZN(n5452)
         );
  AOI211_X1 U6993 ( .C1(n9570), .C2(n5453), .A(n6257), .B(n5452), .ZN(n5455)
         );
  NAND2_X1 U6994 ( .A1(n9432), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n5454) );
  OAI211_X1 U6995 ( .C1(n5456), .C2(n9564), .A(n5455), .B(n5454), .ZN(P1_U3246) );
  OR2_X1 U6996 ( .A1(n5685), .A2(n5588), .ZN(n5461) );
  OR2_X1 U6997 ( .A1(n5686), .A2(n5457), .ZN(n5460) );
  OR2_X1 U6998 ( .A1(n5458), .A2(n9430), .ZN(n5459) );
  XNOR2_X2 U6999 ( .A(n5462), .B(n5469), .ZN(n5464) );
  INV_X1 U7000 ( .A(n5997), .ZN(n5483) );
  OR2_X1 U7001 ( .A1(n5660), .A2(n5357), .ZN(n5468) );
  NAND3_X1 U7002 ( .A1(n8886), .A2(n8931), .A3(n5466), .ZN(n5467) );
  AND2_X1 U7003 ( .A1(n5468), .A2(n5467), .ZN(n9615) );
  NAND2_X1 U7004 ( .A1(n8682), .A2(n5984), .ZN(n5991) );
  OR2_X1 U7005 ( .A1(n5982), .A2(n8932), .ZN(n9680) );
  INV_X1 U7006 ( .A(n9680), .ZN(n9633) );
  OR2_X1 U7007 ( .A1(n8682), .A2(n5984), .ZN(n6433) );
  NAND3_X1 U7008 ( .A1(n5991), .A2(n9633), .A3(n6433), .ZN(n5470) );
  OAI21_X1 U7009 ( .B1(n9678), .B2(n5469), .A(n5470), .ZN(n5482) );
  INV_X1 U7010 ( .A(n9357), .ZN(n9610) );
  NAND2_X1 U7011 ( .A1(n7983), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U7012 ( .A1(n4281), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U7013 ( .A1(n5471), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U7014 ( .A1(n5472), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5473) );
  OR2_X1 U7015 ( .A1(n5477), .A2(n5145), .ZN(n9608) );
  INV_X1 U7016 ( .A(n5463), .ZN(n5481) );
  NOR2_X1 U7017 ( .A1(n5463), .A2(n5540), .ZN(n6024) );
  NAND2_X1 U7018 ( .A1(n5393), .A2(n9588), .ZN(n5479) );
  OR2_X1 U7019 ( .A1(n6522), .A2(n6395), .ZN(n5478) );
  OAI222_X1 U7020 ( .A1(n9610), .A2(n6023), .B1(n9608), .B2(n5481), .C1(n5480), 
        .C2(n9591), .ZN(n5994) );
  AOI211_X1 U7021 ( .C1(n5483), .C2(n9684), .A(n5482), .B(n5994), .ZN(n10015)
         );
  OAI211_X1 U7022 ( .C1(n9638), .C2(n8931), .A(n5485), .B(n5484), .ZN(n5486)
         );
  NAND2_X1 U7023 ( .A1(n9697), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5488) );
  OAI21_X1 U7024 ( .B1(n10015), .B2(n9697), .A(n5488), .ZN(P1_U3524) );
  AOI211_X1 U7025 ( .C1(n5491), .C2(n5490), .A(n5489), .B(n6466), .ZN(n5501)
         );
  AOI22_X1 U7026 ( .A1(n9747), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n5499) );
  INV_X1 U7027 ( .A(n5492), .ZN(n5494) );
  MUX2_X1 U7028 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n5210), .S(n5759), .Z(n5493)
         );
  NAND2_X1 U7029 ( .A1(n5494), .A2(n5493), .ZN(n5496) );
  OAI211_X1 U7030 ( .C1(n5497), .C2(n5496), .A(n9753), .B(n5495), .ZN(n5498)
         );
  OAI211_X1 U7031 ( .C1(n9739), .C2(n5759), .A(n5499), .B(n5498), .ZN(n5500)
         );
  OR2_X1 U7032 ( .A1(n5501), .A2(n5500), .ZN(P2_U3248) );
  NOR2_X1 U7033 ( .A1(n6482), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5503) );
  NOR2_X1 U7034 ( .A1(n5503), .A2(n5502), .ZN(n5730) );
  INV_X1 U7035 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5728) );
  XNOR2_X1 U7036 ( .A(n6734), .B(n5728), .ZN(n5504) );
  XNOR2_X1 U7037 ( .A(n5730), .B(n5504), .ZN(n5518) );
  INV_X1 U7038 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n5515) );
  INV_X1 U7039 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6910) );
  MUX2_X1 U7040 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6910), .S(n6734), .Z(n5512)
         );
  OR2_X1 U7041 ( .A1(n5506), .A2(n5505), .ZN(n5507) );
  OAI21_X1 U7042 ( .B1(n9952), .B2(n5508), .A(n5507), .ZN(n5509) );
  INV_X1 U7043 ( .A(n5509), .ZN(n5511) );
  INV_X1 U7044 ( .A(n5722), .ZN(n5510) );
  OAI21_X1 U7045 ( .B1(n5512), .B2(n5511), .A(n5510), .ZN(n5513) );
  NAND2_X1 U7046 ( .A1(n9753), .A2(n5513), .ZN(n5514) );
  NAND2_X1 U7047 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6805) );
  OAI211_X1 U7048 ( .C1(n6298), .C2(n5515), .A(n5514), .B(n6805), .ZN(n5516)
         );
  AOI21_X1 U7049 ( .B1(n6734), .B2(n9757), .A(n5516), .ZN(n5517) );
  OAI21_X1 U7050 ( .B1(n5518), .B2(n6466), .A(n5517), .ZN(P2_U3257) );
  NOR3_X1 U7051 ( .A1(n6466), .A2(P2_REG2_REG_5__SCAN_IN), .A3(n5531), .ZN(
        n5521) );
  INV_X1 U7052 ( .A(n5519), .ZN(n5523) );
  NOR3_X1 U7053 ( .A1(n9740), .A2(P2_REG1_REG_5__SCAN_IN), .A3(n5523), .ZN(
        n5520) );
  NOR3_X1 U7054 ( .A1(n5521), .A2(n9757), .A3(n5520), .ZN(n5535) );
  INV_X1 U7055 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n5527) );
  NOR2_X1 U7056 ( .A1(n5529), .A2(n9828), .ZN(n5524) );
  OAI211_X1 U7057 ( .C1(n5524), .C2(n5523), .A(n9753), .B(n5522), .ZN(n5526)
         );
  AND2_X1 U7058 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9727) );
  INV_X1 U7059 ( .A(n9727), .ZN(n5525) );
  OAI211_X1 U7060 ( .C1(n6298), .C2(n5527), .A(n5526), .B(n5525), .ZN(n5528)
         );
  INV_X1 U7061 ( .A(n5528), .ZN(n5534) );
  NOR2_X1 U7062 ( .A1(n5529), .A2(n5235), .ZN(n5532) );
  OAI211_X1 U7063 ( .C1(n5532), .C2(n5531), .A(n9749), .B(n5530), .ZN(n5533)
         );
  OAI211_X1 U7064 ( .C1(n5535), .C2(n5924), .A(n5534), .B(n5533), .ZN(P2_U3250) );
  AND2_X1 U7065 ( .A1(n5540), .A2(n5463), .ZN(n8679) );
  NOR2_X1 U7066 ( .A1(n8679), .A2(n6024), .ZN(n8899) );
  OR3_X1 U7067 ( .A1(n8899), .A2(n8935), .A3(n5536), .ZN(n5538) );
  NAND2_X1 U7068 ( .A1(n9357), .A2(n5462), .ZN(n5537) );
  NAND2_X1 U7069 ( .A1(n5538), .A2(n5537), .ZN(n5986) );
  INV_X1 U7070 ( .A(n5986), .ZN(n5539) );
  OAI21_X1 U7071 ( .B1(n5540), .B2(n5982), .A(n5539), .ZN(n5626) );
  NAND2_X1 U7072 ( .A1(n5626), .A2(n4269), .ZN(n5541) );
  OAI21_X1 U7073 ( .B1(n4269), .B2(n9441), .A(n5541), .ZN(P1_U3523) );
  INV_X1 U7074 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n5554) );
  AOI21_X1 U7075 ( .B1(n5543), .B2(n5542), .A(n4356), .ZN(n5551) );
  AND2_X1 U7076 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6200) );
  AOI21_X1 U7077 ( .B1(n9570), .B2(n5544), .A(n6200), .ZN(n5550) );
  AOI21_X1 U7078 ( .B1(n5547), .B2(n5546), .A(n5545), .ZN(n5548) );
  OR2_X1 U7079 ( .A1(n9576), .A2(n5548), .ZN(n5549) );
  OAI211_X1 U7080 ( .C1(n9564), .C2(n5551), .A(n5550), .B(n5549), .ZN(n5552)
         );
  INV_X1 U7081 ( .A(n5552), .ZN(n5553) );
  OAI21_X1 U7082 ( .B1(n5554), .B2(n9579), .A(n5553), .ZN(P1_U3248) );
  AOI21_X1 U7083 ( .B1(n5557), .B2(n5556), .A(n5555), .ZN(n5558) );
  NOR2_X1 U7084 ( .A1(n9576), .A2(n5558), .ZN(n5566) );
  AOI21_X1 U7085 ( .B1(n5561), .B2(n5560), .A(n5559), .ZN(n5564) );
  NAND2_X1 U7086 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n5902) );
  INV_X1 U7087 ( .A(n5885), .ZN(n5562) );
  NAND2_X1 U7088 ( .A1(n9570), .A2(n5562), .ZN(n5563) );
  OAI211_X1 U7089 ( .C1(n9564), .C2(n5564), .A(n5902), .B(n5563), .ZN(n5565)
         );
  AOI211_X1 U7090 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9432), .A(n5566), .B(
        n5565), .ZN(n5568) );
  NAND2_X1 U7091 ( .A1(n5568), .A2(n5567), .ZN(P1_U3245) );
  INV_X1 U7092 ( .A(n5569), .ZN(n5573) );
  INV_X1 U7093 ( .A(n5570), .ZN(n5571) );
  NAND2_X1 U7094 ( .A1(n5571), .A2(SI_14_), .ZN(n5572) );
  INV_X1 U7095 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5650) );
  INV_X1 U7096 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5575) );
  MUX2_X1 U7097 ( .A(n5650), .B(n5575), .S(n7537), .Z(n5576) );
  INV_X1 U7098 ( .A(SI_15_), .ZN(n9923) );
  NAND2_X1 U7099 ( .A1(n5576), .A2(n9923), .ZN(n5629) );
  INV_X1 U7100 ( .A(n5576), .ZN(n5577) );
  NAND2_X1 U7101 ( .A1(n5577), .A2(SI_15_), .ZN(n5578) );
  NAND2_X1 U7102 ( .A1(n5629), .A2(n5578), .ZN(n5630) );
  XNOR2_X1 U7103 ( .A(n5631), .B(n5630), .ZN(n7095) );
  INV_X1 U7104 ( .A(n7095), .ZN(n5649) );
  NAND2_X1 U7105 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  NAND2_X1 U7106 ( .A1(n5581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5582) );
  XNOR2_X1 U7107 ( .A(n5582), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9532) );
  AOI22_X1 U7108 ( .A1(n9532), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n5848), .ZN(n5583) );
  OAI21_X1 U7109 ( .B1(n5649), .B2(n8059), .A(n5583), .ZN(P1_U3338) );
  INV_X1 U7110 ( .A(n6098), .ZN(n5584) );
  INV_X1 U7111 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7112 ( .A1(n5602), .A2(n5587), .ZN(n5907) );
  OR2_X1 U7113 ( .A1(n5907), .A2(n5588), .ZN(n5591) );
  NAND2_X1 U7114 ( .A1(n5593), .A2(n9774), .ZN(n8410) );
  NAND2_X1 U7115 ( .A1(n5110), .A2(n5108), .ZN(n8404) );
  INV_X1 U7116 ( .A(n9774), .ZN(n8405) );
  NAND2_X1 U7117 ( .A1(n5595), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7118 ( .A1(n7320), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5596) );
  OR2_X1 U7119 ( .A1(n5907), .A2(n5671), .ZN(n5605) );
  OR2_X1 U7120 ( .A1(n7540), .A2(n5600), .ZN(n5604) );
  OR2_X1 U7121 ( .A1(n5602), .A2(n5601), .ZN(n5603) );
  NAND2_X1 U7122 ( .A1(n8418), .A2(n6109), .ZN(n7583) );
  INV_X1 U7123 ( .A(n5606), .ZN(n6110) );
  INV_X1 U7124 ( .A(n8414), .ZN(n8326) );
  INV_X1 U7125 ( .A(n8326), .ZN(n8384) );
  OAI21_X1 U7126 ( .B1(n5608), .B2(n5607), .A(n5857), .ZN(n5616) );
  NAND2_X1 U7127 ( .A1(n5595), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7128 ( .A1(n5609), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5611) );
  INV_X1 U7129 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7130 ( .A1(n5775), .A2(n5839), .ZN(n5610) );
  NAND2_X1 U7131 ( .A1(n5791), .A2(n5615), .ZN(n8328) );
  INV_X1 U7132 ( .A(n8328), .ZN(n8419) );
  AOI222_X1 U7133 ( .A1(n8384), .A2(n5616), .B1(n8159), .B2(n8417), .C1(n5593), 
        .C2(n8419), .ZN(n6105) );
  INV_X1 U7134 ( .A(n6109), .ZN(n5850) );
  NAND2_X1 U7135 ( .A1(n9774), .A2(n5970), .ZN(n5618) );
  OR2_X1 U7136 ( .A1(n5618), .A2(n5850), .ZN(n6443) );
  AND2_X4 U7137 ( .A1(n5617), .A2(n6358), .ZN(n9810) );
  NAND2_X1 U7138 ( .A1(n5618), .A2(n5850), .ZN(n5619) );
  AND3_X1 U7139 ( .A1(n6443), .A2(n9810), .A3(n5619), .ZN(n6102) );
  AOI21_X1 U7140 ( .B1(n9809), .B2(n5850), .A(n6102), .ZN(n5620) );
  OAI211_X1 U7141 ( .C1(n9804), .C2(n6110), .A(n6105), .B(n5620), .ZN(n5623)
         );
  NAND2_X1 U7142 ( .A1(n4267), .A2(n5623), .ZN(n5621) );
  OAI21_X1 U7143 ( .B1(n4267), .B2(n5622), .A(n5621), .ZN(P2_U3457) );
  NAND2_X1 U7144 ( .A1(n4268), .A2(n5623), .ZN(n5624) );
  OAI21_X1 U7145 ( .B1(n4268), .B2(n5207), .A(n5624), .ZN(P2_U3522) );
  INV_X1 U7146 ( .A(n5977), .ZN(n9628) );
  INV_X2 U7147 ( .A(n9686), .ZN(n10017) );
  INV_X1 U7148 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7149 ( .A1(n5626), .A2(n10017), .ZN(n5627) );
  OAI21_X1 U7150 ( .B1(n10017), .B2(n5628), .A(n5627), .ZN(P1_U3454) );
  INV_X1 U7151 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5633) );
  INV_X1 U7152 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5632) );
  MUX2_X1 U7153 ( .A(n5633), .B(n5632), .S(n4276), .Z(n5635) );
  INV_X1 U7154 ( .A(SI_16_), .ZN(n5634) );
  NAND2_X1 U7155 ( .A1(n5635), .A2(n5634), .ZN(n5846) );
  INV_X1 U7156 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U7157 ( .A1(n5636), .A2(SI_16_), .ZN(n5637) );
  XNOR2_X1 U7158 ( .A(n5845), .B(n5844), .ZN(n7241) );
  INV_X1 U7159 ( .A(n7241), .ZN(n5646) );
  NAND2_X1 U7160 ( .A1(n5638), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5639) );
  XNOR2_X1 U7161 ( .A(n5639), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9543) );
  AOI22_X1 U7162 ( .A1(n9543), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n5848), .ZN(n5640) );
  OAI21_X1 U7163 ( .B1(n5646), .B2(n8059), .A(n5640), .ZN(P1_U3337) );
  NAND2_X1 U7164 ( .A1(n5641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5642) );
  MUX2_X1 U7165 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5642), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5644) );
  AND2_X1 U7166 ( .A1(n5644), .A2(n5643), .ZN(n7176) );
  AOI22_X1 U7167 ( .A1(n7176), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8540), .ZN(n5645) );
  OAI21_X1 U7168 ( .B1(n5646), .B2(n4270), .A(n5645), .ZN(P2_U3342) );
  NAND2_X1 U7169 ( .A1(n5647), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5648) );
  XNOR2_X1 U7170 ( .A(n5648), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7067) );
  INV_X1 U7171 ( .A(n7067), .ZN(n6300) );
  OAI222_X1 U7172 ( .A1(n8545), .A2(n5650), .B1(n4270), .B2(n5649), .C1(
        P2_U3152), .C2(n6300), .ZN(P2_U3343) );
  AND3_X1 U7173 ( .A1(n5653), .A2(n5652), .A3(n5651), .ZN(n5655) );
  NAND2_X1 U7174 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  NAND2_X1 U7175 ( .A1(n5656), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7176 ( .A1(n5658), .A2(n5657), .ZN(n8660) );
  INV_X1 U7177 ( .A(n8660), .ZN(n8646) );
  INV_X1 U7178 ( .A(n5659), .ZN(n5661) );
  NAND2_X1 U7179 ( .A1(n5660), .A2(n5359), .ZN(n5663) );
  NAND2_X1 U7180 ( .A1(n5676), .A2(n5462), .ZN(n5662) );
  OAI21_X1 U7181 ( .B1(n5469), .B2(n7900), .A(n5662), .ZN(n5664) );
  XNOR2_X1 U7182 ( .A(n5664), .B(n5663), .ZN(n5667) );
  INV_X1 U7183 ( .A(n5667), .ZN(n5665) );
  NAND3_X1 U7184 ( .A1(n5668), .A2(n5667), .A3(n5666), .ZN(n5669) );
  INV_X2 U7185 ( .A(n5676), .ZN(n6180) );
  NOR2_X1 U7186 ( .A1(n5469), .A2(n6180), .ZN(n5670) );
  AOI21_X1 U7187 ( .B1(n7974), .B2(n5462), .A(n5670), .ZN(n8578) );
  NAND2_X1 U7188 ( .A1(n7487), .A2(n7484), .ZN(n5684) );
  OR2_X1 U7189 ( .A1(n5686), .A2(n5672), .ZN(n5673) );
  OAI211_X2 U7190 ( .C1(n5364), .C2(n5675), .A(n5674), .B(n5673), .ZN(n6022)
         );
  NAND2_X1 U7191 ( .A1(n7974), .A2(n6029), .ZN(n5678) );
  NAND2_X1 U7192 ( .A1(n4265), .A2(n6022), .ZN(n5677) );
  AND2_X1 U7193 ( .A1(n5678), .A2(n5677), .ZN(n5680) );
  NAND2_X1 U7194 ( .A1(n5679), .A2(n5680), .ZN(n5706) );
  INV_X1 U7195 ( .A(n5680), .ZN(n5681) );
  NAND2_X1 U7196 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  AND2_X1 U7197 ( .A1(n5706), .A2(n5683), .ZN(n7485) );
  NAND2_X1 U7198 ( .A1(n5684), .A2(n7485), .ZN(n5707) );
  INV_X1 U7199 ( .A(n5707), .ZN(n7488) );
  INV_X1 U7200 ( .A(n5706), .ZN(n5705) );
  OR2_X1 U7201 ( .A1(n5685), .A2(n5757), .ZN(n5689) );
  INV_X1 U7202 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5713) );
  NAND2_X1 U7203 ( .A1(n4281), .A2(n5713), .ZN(n5695) );
  NAND2_X1 U7204 ( .A1(n7983), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7205 ( .A1(n5471), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U7206 ( .A1(n4275), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5692) );
  OR2_X1 U7207 ( .A1(n6414), .A2(n6180), .ZN(n5696) );
  OAI21_X1 U7208 ( .B1(n9641), .B2(n7900), .A(n5696), .ZN(n5697) );
  XNOR2_X1 U7209 ( .A(n5697), .B(n8009), .ZN(n5700) );
  INV_X1 U7210 ( .A(n6414), .ZN(n8953) );
  NAND2_X1 U7211 ( .A1(n7974), .A2(n8953), .ZN(n5699) );
  NAND2_X1 U7212 ( .A1(n4265), .A2(n6031), .ZN(n5698) );
  AND2_X1 U7213 ( .A1(n5699), .A2(n5698), .ZN(n5701) );
  NAND2_X1 U7214 ( .A1(n5700), .A2(n5701), .ZN(n5890) );
  INV_X1 U7215 ( .A(n5700), .ZN(n5703) );
  INV_X1 U7216 ( .A(n5701), .ZN(n5702) );
  NAND2_X1 U7217 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  AND2_X1 U7218 ( .A1(n5890), .A2(n5704), .ZN(n5708) );
  NOR3_X1 U7219 ( .A1(n7488), .A2(n5705), .A3(n5708), .ZN(n5711) );
  NAND2_X1 U7220 ( .A1(n5707), .A2(n5706), .ZN(n5709) );
  NAND2_X1 U7221 ( .A1(n5709), .A2(n5708), .ZN(n5891) );
  INV_X1 U7222 ( .A(n5891), .ZN(n5710) );
  OAI21_X1 U7223 ( .B1(n5711), .B2(n5710), .A(n8652), .ZN(n5721) );
  NAND2_X1 U7224 ( .A1(n7983), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5717) );
  XNOR2_X1 U7225 ( .A(n5713), .B(P1_REG3_REG_4__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7226 ( .A1(n4281), .A2(n5881), .ZN(n5716) );
  NAND2_X1 U7227 ( .A1(n7826), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7228 ( .A1(n5471), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5714) );
  AND2_X1 U7229 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9332) );
  OR2_X1 U7230 ( .A1(n5718), .A2(n5145), .ZN(n8656) );
  OAI22_X1 U7231 ( .A1(n8663), .A2(n9641), .B1(n8656), .B2(n6023), .ZN(n5719)
         );
  AOI211_X1 U7232 ( .C1(n8644), .C2(n8952), .A(n9332), .B(n5719), .ZN(n5720)
         );
  OAI211_X1 U7233 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8646), .A(n5721), .B(
        n5720), .ZN(P1_U3216) );
  INV_X1 U7234 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5724) );
  AOI21_X1 U7235 ( .B1(n6910), .B2(n5723), .A(n5722), .ZN(n5874) );
  AOI22_X1 U7236 ( .A1(n6833), .A2(n5724), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n5880), .ZN(n5873) );
  NOR2_X1 U7237 ( .A1(n5874), .A2(n5873), .ZN(n5872) );
  AOI21_X1 U7238 ( .B1(n5880), .B2(n5724), .A(n5872), .ZN(n5726) );
  INV_X1 U7239 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6012) );
  AOI22_X1 U7240 ( .A1(n7010), .A2(n6012), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n6013), .ZN(n5725) );
  NOR2_X1 U7241 ( .A1(n5726), .A2(n5725), .ZN(n6011) );
  AOI21_X1 U7242 ( .B1(n5726), .B2(n5725), .A(n6011), .ZN(n5739) );
  INV_X1 U7243 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5727) );
  AOI22_X1 U7244 ( .A1(n7010), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n5727), .B2(
        n6013), .ZN(n5734) );
  INV_X1 U7245 ( .A(n5730), .ZN(n5729) );
  NOR2_X1 U7246 ( .A1(n5729), .A2(n5728), .ZN(n5731) );
  OAI22_X1 U7247 ( .A1(n5731), .A2(n6734), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n5730), .ZN(n5870) );
  NOR2_X1 U7248 ( .A1(n6833), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5732) );
  AOI21_X1 U7249 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n6833), .A(n5732), .ZN(
        n5869) );
  NAND2_X1 U7250 ( .A1(n5870), .A2(n5869), .ZN(n5868) );
  OAI21_X1 U7251 ( .B1(n6833), .B2(P2_REG2_REG_13__SCAN_IN), .A(n5868), .ZN(
        n5733) );
  NAND2_X1 U7252 ( .A1(n5734), .A2(n5733), .ZN(n6015) );
  OAI21_X1 U7253 ( .B1(n5734), .B2(n5733), .A(n6015), .ZN(n5737) );
  AND2_X1 U7254 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7048) );
  AOI21_X1 U7255 ( .B1(n9747), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7048), .ZN(
        n5735) );
  OAI21_X1 U7256 ( .B1(n9739), .B2(n6013), .A(n5735), .ZN(n5736) );
  AOI21_X1 U7257 ( .B1(n5737), .B2(n9749), .A(n5736), .ZN(n5738) );
  OAI21_X1 U7258 ( .B1(n5739), .B2(n9740), .A(n5738), .ZN(P2_U3259) );
  NAND3_X1 U7259 ( .A1(n5741), .A2(n7747), .A3(n5740), .ZN(n5742) );
  NAND2_X1 U7260 ( .A1(n5742), .A2(n6106), .ZN(n5750) );
  XNOR2_X1 U7261 ( .A(n5750), .B(n9774), .ZN(n5744) );
  INV_X1 U7262 ( .A(n8404), .ZN(n5745) );
  OR2_X1 U7263 ( .A1(n4263), .A2(n5108), .ZN(n5746) );
  NAND2_X1 U7264 ( .A1(n5747), .A2(n5746), .ZN(n5819) );
  INV_X1 U7265 ( .A(n5819), .ZN(n5748) );
  NAND2_X1 U7266 ( .A1(n5817), .A2(n5749), .ZN(n5830) );
  XNOR2_X1 U7267 ( .A(n4263), .B(n6109), .ZN(n5754) );
  INV_X1 U7268 ( .A(n5754), .ZN(n5752) );
  NAND2_X1 U7269 ( .A1(n5763), .A2(n8418), .ZN(n5753) );
  INV_X1 U7270 ( .A(n5753), .ZN(n5751) );
  NAND2_X1 U7271 ( .A1(n5752), .A2(n5751), .ZN(n5755) );
  NAND2_X1 U7272 ( .A1(n5754), .A2(n5753), .ZN(n5756) );
  NAND2_X1 U7273 ( .A1(n5831), .A2(n5756), .ZN(n5837) );
  INV_X1 U7274 ( .A(n5837), .ZN(n5769) );
  OR2_X1 U7275 ( .A1(n5907), .A2(n5757), .ZN(n5762) );
  OR2_X1 U7276 ( .A1(n7540), .A2(n5758), .ZN(n5761) );
  OR2_X1 U7277 ( .A1(n5602), .A2(n5759), .ZN(n5760) );
  XNOR2_X1 U7278 ( .A(n4263), .B(n9780), .ZN(n5764) );
  NAND2_X1 U7279 ( .A1(n8041), .A2(n8159), .ZN(n5765) );
  XNOR2_X1 U7280 ( .A(n5764), .B(n5765), .ZN(n5836) );
  INV_X1 U7281 ( .A(n5836), .ZN(n5768) );
  INV_X1 U7282 ( .A(n5764), .ZN(n5767) );
  INV_X1 U7283 ( .A(n5765), .ZN(n5766) );
  AOI21_X1 U7284 ( .B1(n5769), .B2(n5768), .A(n4807), .ZN(n5787) );
  OR2_X1 U7285 ( .A1(n7540), .A2(n5770), .ZN(n5773) );
  OR2_X1 U7286 ( .A1(n5602), .A2(n5771), .ZN(n5772) );
  XNOR2_X1 U7287 ( .A(n8043), .B(n6118), .ZN(n5781) );
  NAND2_X1 U7288 ( .A1(n7320), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7289 ( .A1(n5595), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5779) );
  XNOR2_X1 U7290 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6113) );
  INV_X1 U7291 ( .A(n6113), .ZN(n5776) );
  NAND2_X1 U7292 ( .A1(n7518), .A2(n5776), .ZN(n5778) );
  OR2_X1 U7293 ( .A1(n7458), .A2(n5867), .ZN(n5777) );
  NAND2_X1 U7294 ( .A1(n8041), .A2(n8158), .ZN(n5782) );
  NAND2_X1 U7295 ( .A1(n5781), .A2(n5782), .ZN(n5921) );
  INV_X1 U7296 ( .A(n5781), .ZN(n5784) );
  INV_X1 U7297 ( .A(n5782), .ZN(n5783) );
  NAND2_X1 U7298 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  AND2_X1 U7299 ( .A1(n5921), .A2(n5785), .ZN(n5786) );
  NAND2_X1 U7300 ( .A1(n5787), .A2(n5786), .ZN(n5922) );
  OAI21_X1 U7301 ( .B1(n5787), .B2(n5786), .A(n5922), .ZN(n5815) );
  AND2_X1 U7302 ( .A1(n5789), .A2(n5788), .ZN(n6097) );
  INV_X1 U7303 ( .A(n6097), .ZN(n5790) );
  NOR2_X1 U7304 ( .A1(n5793), .A2(n9763), .ZN(n5803) );
  INV_X1 U7305 ( .A(n5803), .ZN(n5792) );
  INV_X1 U7306 ( .A(n8128), .ZN(n9733) );
  NAND2_X1 U7307 ( .A1(n5793), .A2(n6100), .ZN(n5822) );
  INV_X1 U7308 ( .A(n5794), .ZN(n5795) );
  AND3_X1 U7309 ( .A1(n5796), .A2(n5795), .A3(n6096), .ZN(n5797) );
  NAND2_X1 U7310 ( .A1(n5822), .A2(n5797), .ZN(n5798) );
  NAND2_X1 U7311 ( .A1(n5798), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9737) );
  INV_X1 U7312 ( .A(n9809), .ZN(n9820) );
  NOR2_X1 U7313 ( .A1(n9763), .A2(n9820), .ZN(n5799) );
  INV_X1 U7314 ( .A(n6118), .ZN(n6135) );
  NAND2_X1 U7315 ( .A1(n8147), .A2(n6135), .ZN(n5800) );
  OAI211_X1 U7316 ( .C1(n9737), .C2(n6113), .A(n5801), .B(n5800), .ZN(n5814)
         );
  INV_X1 U7317 ( .A(n7755), .ZN(n5802) );
  NAND2_X1 U7318 ( .A1(n5803), .A2(n5802), .ZN(n8142) );
  NOR2_X1 U7319 ( .A1(n8142), .A2(n8328), .ZN(n9717) );
  INV_X1 U7320 ( .A(n8159), .ZN(n5854) );
  NAND2_X1 U7321 ( .A1(n5609), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7322 ( .A1(n7320), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5811) );
  INV_X1 U7323 ( .A(n5912), .ZN(n5807) );
  INV_X1 U7324 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7325 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5804) );
  NAND2_X1 U7326 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  NAND2_X1 U7327 ( .A1(n5807), .A2(n5806), .ZN(n9736) );
  INV_X1 U7328 ( .A(n9736), .ZN(n5808) );
  NAND2_X1 U7329 ( .A1(n7518), .A2(n5808), .ZN(n5810) );
  NAND2_X1 U7330 ( .A1(n5595), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5809) );
  NAND4_X1 U7331 ( .A1(n5812), .A2(n5811), .A3(n5810), .A4(n5809), .ZN(n8157)
         );
  INV_X1 U7332 ( .A(n8157), .ZN(n5941) );
  OAI22_X1 U7333 ( .A1(n8135), .A2(n5854), .B1(n5941), .B2(n9714), .ZN(n5813)
         );
  AOI211_X1 U7334 ( .C1(n5815), .C2(n9733), .A(n5814), .B(n5813), .ZN(n5816)
         );
  INV_X1 U7335 ( .A(n5816), .ZN(P2_U3232) );
  INV_X1 U7336 ( .A(n5817), .ZN(n5818) );
  AOI21_X1 U7337 ( .B1(n5820), .B2(n5819), .A(n5818), .ZN(n5827) );
  INV_X1 U7338 ( .A(n9714), .ZN(n5840) );
  INV_X1 U7339 ( .A(n8147), .ZN(n9731) );
  AND3_X1 U7340 ( .A1(n5822), .A2(n5821), .A3(n6096), .ZN(n5969) );
  OAI22_X1 U7341 ( .A1(n9731), .A2(n9774), .B1(n5969), .B2(n5823), .ZN(n5824)
         );
  AOI21_X1 U7342 ( .B1(n5840), .B2(n8418), .A(n5824), .ZN(n5826) );
  NAND2_X1 U7343 ( .A1(n9717), .A2(n5110), .ZN(n5825) );
  OAI211_X1 U7344 ( .C1(n5827), .C2(n8128), .A(n5826), .B(n5825), .ZN(P2_U3224) );
  INV_X1 U7345 ( .A(n5593), .ZN(n5975) );
  INV_X1 U7346 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5828) );
  OAI22_X1 U7347 ( .A1(n9731), .A2(n6109), .B1(n5969), .B2(n5828), .ZN(n5829)
         );
  AOI21_X1 U7348 ( .B1(n5840), .B2(n8159), .A(n5829), .ZN(n5835) );
  OAI21_X1 U7349 ( .B1(n5832), .B2(n5830), .A(n5831), .ZN(n5833) );
  NAND2_X1 U7350 ( .A1(n5833), .A2(n9733), .ZN(n5834) );
  OAI211_X1 U7351 ( .C1(n5975), .C2(n8135), .A(n5835), .B(n5834), .ZN(P2_U3239) );
  XNOR2_X1 U7352 ( .A(n5837), .B(n5836), .ZN(n5843) );
  INV_X1 U7353 ( .A(n9737), .ZN(n8140) );
  OAI22_X1 U7354 ( .A1(n9731), .A2(n9780), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5839), .ZN(n5838) );
  AOI21_X1 U7355 ( .B1(n8140), .B2(n5839), .A(n5838), .ZN(n5842) );
  AOI22_X1 U7356 ( .A1(n9717), .A2(n8418), .B1(n5840), .B2(n8158), .ZN(n5841)
         );
  OAI211_X1 U7357 ( .C1(n5843), .C2(n8128), .A(n5842), .B(n5841), .ZN(P2_U3220) );
  INV_X1 U7358 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5951) );
  INV_X1 U7359 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5847) );
  MUX2_X1 U7360 ( .A(n5951), .B(n5847), .S(n4276), .Z(n5999) );
  XNOR2_X1 U7361 ( .A(n5999), .B(SI_17_), .ZN(n5998) );
  XNOR2_X1 U7362 ( .A(n6002), .B(n5998), .ZN(n7269) );
  INV_X1 U7363 ( .A(n7269), .ZN(n5950) );
  NAND2_X1 U7364 ( .A1(n4340), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6004) );
  XNOR2_X1 U7365 ( .A(n6004), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9555) );
  AOI22_X1 U7366 ( .A1(n9555), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n5848), .ZN(n5849) );
  OAI21_X1 U7367 ( .B1(n5950), .B2(n8059), .A(n5849), .ZN(P1_U3336) );
  INV_X1 U7368 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5864) );
  OR2_X1 U7369 ( .A1(n8418), .A2(n5850), .ZN(n5851) );
  NAND2_X1 U7370 ( .A1(n8159), .A2(n9780), .ZN(n7588) );
  NAND2_X1 U7371 ( .A1(n6441), .A2(n7719), .ZN(n6440) );
  OR2_X1 U7372 ( .A1(n8159), .A2(n5853), .ZN(n5855) );
  NAND2_X1 U7373 ( .A1(n8158), .A2(n6118), .ZN(n7589) );
  OAI21_X1 U7374 ( .B1(n5856), .B2(n6140), .A(n6136), .ZN(n6120) );
  INV_X1 U7375 ( .A(n6120), .ZN(n5862) );
  NAND2_X1 U7376 ( .A1(n5857), .A2(n7581), .ZN(n6448) );
  NAND2_X1 U7377 ( .A1(n6448), .A2(n7576), .ZN(n6142) );
  NAND2_X1 U7378 ( .A1(n6142), .A2(n7568), .ZN(n5858) );
  XOR2_X1 U7379 ( .A(n6140), .B(n5858), .Z(n5859) );
  AOI222_X1 U7380 ( .A1(n8384), .A2(n5859), .B1(n8157), .B2(n8417), .C1(n8159), 
        .C2(n8419), .ZN(n6122) );
  INV_X1 U7381 ( .A(n5860), .ZN(n6444) );
  INV_X1 U7382 ( .A(n9810), .ZN(n9781) );
  AOI211_X1 U7383 ( .C1(n6135), .C2(n6444), .A(n9781), .B(n4355), .ZN(n6116)
         );
  AOI21_X1 U7384 ( .B1(n9809), .B2(n6135), .A(n6116), .ZN(n5861) );
  OAI211_X1 U7385 ( .C1(n9804), .C2(n5862), .A(n6122), .B(n5861), .ZN(n5865)
         );
  NAND2_X1 U7386 ( .A1(n5865), .A2(n4267), .ZN(n5863) );
  OAI21_X1 U7387 ( .B1(n4267), .B2(n5864), .A(n5863), .ZN(P2_U3463) );
  NAND2_X1 U7388 ( .A1(n5865), .A2(n4268), .ZN(n5866) );
  OAI21_X1 U7389 ( .B1(n4268), .B2(n5867), .A(n5866), .ZN(P2_U3524) );
  OAI21_X1 U7390 ( .B1(n5870), .B2(n5869), .A(n5868), .ZN(n5871) );
  NAND2_X1 U7391 ( .A1(n5871), .A2(n9749), .ZN(n5879) );
  NAND2_X1 U7392 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6847) );
  INV_X1 U7393 ( .A(n6847), .ZN(n5877) );
  AOI21_X1 U7394 ( .B1(n5874), .B2(n5873), .A(n5872), .ZN(n5875) );
  NOR2_X1 U7395 ( .A1(n9740), .A2(n5875), .ZN(n5876) );
  AOI211_X1 U7396 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n9747), .A(n5877), .B(
        n5876), .ZN(n5878) );
  OAI211_X1 U7397 ( .C1(n9739), .C2(n5880), .A(n5879), .B(n5878), .ZN(P2_U3258) );
  INV_X1 U7398 ( .A(n5881), .ZN(n6419) );
  OR2_X1 U7399 ( .A1(n5685), .A2(n5882), .ZN(n5884) );
  OR2_X1 U7400 ( .A1(n8732), .A2(n10001), .ZN(n5883) );
  OAI211_X1 U7401 ( .C1(n5364), .C2(n5885), .A(n5884), .B(n5883), .ZN(n6424)
         );
  INV_X1 U7402 ( .A(n6424), .ZN(n9648) );
  OR2_X1 U7403 ( .A1(n9609), .A2(n6180), .ZN(n5886) );
  OAI21_X1 U7404 ( .B1(n9648), .B2(n7900), .A(n5886), .ZN(n5887) );
  XNOR2_X1 U7405 ( .A(n5887), .B(n8009), .ZN(n6174) );
  NAND2_X1 U7406 ( .A1(n7974), .A2(n8952), .ZN(n5889) );
  NAND2_X1 U7407 ( .A1(n4265), .A2(n6424), .ZN(n5888) );
  NAND2_X1 U7408 ( .A1(n5889), .A2(n5888), .ZN(n6173) );
  XNOR2_X1 U7409 ( .A(n6174), .B(n6173), .ZN(n5893) );
  NAND2_X1 U7410 ( .A1(n5891), .A2(n5890), .ZN(n5892) );
  OAI21_X1 U7411 ( .B1(n5893), .B2(n5892), .A(n6177), .ZN(n5894) );
  NAND2_X1 U7412 ( .A1(n5894), .A2(n8652), .ZN(n5906) );
  NAND2_X1 U7413 ( .A1(n7983), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5901) );
  NAND3_X1 U7414 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6047) );
  INV_X1 U7415 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7416 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5895) );
  NAND2_X1 U7417 ( .A1(n5896), .A2(n5895), .ZN(n5897) );
  AND2_X1 U7418 ( .A1(n6047), .A2(n5897), .ZN(n9585) );
  NAND2_X1 U7419 ( .A1(n4280), .A2(n9585), .ZN(n5900) );
  NAND2_X1 U7420 ( .A1(n7826), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7421 ( .A1(n5471), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5898) );
  INV_X1 U7422 ( .A(n5902), .ZN(n5904) );
  OAI22_X1 U7423 ( .A1(n8663), .A2(n9648), .B1(n8656), .B2(n6414), .ZN(n5903)
         );
  AOI211_X1 U7424 ( .C1(n8644), .C2(n8951), .A(n5904), .B(n5903), .ZN(n5905)
         );
  OAI211_X1 U7425 ( .C1(n8646), .C2(n6419), .A(n5906), .B(n5905), .ZN(P1_U3228) );
  NAND2_X1 U7426 ( .A1(n5908), .A2(n5954), .ZN(n5911) );
  AOI22_X1 U7427 ( .A1(n7339), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7338), .B2(
        n5909), .ZN(n5910) );
  NAND2_X1 U7428 ( .A1(n5911), .A2(n5910), .ZN(n9793) );
  XNOR2_X1 U7429 ( .A(n8043), .B(n9793), .ZN(n5919) );
  NAND2_X1 U7430 ( .A1(n5609), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7431 ( .A1(n7320), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5916) );
  NOR2_X1 U7432 ( .A1(n5912), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5913) );
  NOR2_X1 U7433 ( .A1(n5935), .A2(n5913), .ZN(n5942) );
  NAND2_X1 U7434 ( .A1(n7518), .A2(n5942), .ZN(n5915) );
  NAND2_X1 U7435 ( .A1(n5595), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5914) );
  NAND4_X1 U7436 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n8156)
         );
  AND2_X1 U7437 ( .A1(n8041), .A2(n8156), .ZN(n5918) );
  OR2_X1 U7438 ( .A1(n5919), .A2(n5918), .ZN(n5952) );
  NAND2_X1 U7439 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  AND2_X1 U7440 ( .A1(n5952), .A2(n5920), .ZN(n5934) );
  NAND2_X1 U7441 ( .A1(n5922), .A2(n5921), .ZN(n9725) );
  NAND2_X1 U7442 ( .A1(n5923), .A2(n5954), .ZN(n5928) );
  OR2_X1 U7443 ( .A1(n5602), .A2(n5924), .ZN(n5927) );
  OR2_X1 U7444 ( .A1(n7540), .A2(n5925), .ZN(n5926) );
  XNOR2_X1 U7445 ( .A(n8043), .B(n9790), .ZN(n5930) );
  NAND2_X1 U7446 ( .A1(n8041), .A2(n8157), .ZN(n5929) );
  NAND2_X1 U7447 ( .A1(n5930), .A2(n5929), .ZN(n5932) );
  OR2_X1 U7448 ( .A1(n5930), .A2(n5929), .ZN(n5931) );
  AND2_X1 U7449 ( .A1(n5932), .A2(n5931), .ZN(n9726) );
  OAI21_X1 U7450 ( .B1(n5934), .B2(n5933), .A(n5953), .ZN(n5947) );
  NAND2_X1 U7451 ( .A1(n7320), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7452 ( .A1(n5595), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5939) );
  NOR2_X1 U7453 ( .A1(n5935), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5936) );
  NOR2_X1 U7454 ( .A1(n5959), .A2(n5936), .ZN(n5957) );
  NAND2_X1 U7455 ( .A1(n7518), .A2(n5957), .ZN(n5938) );
  NAND2_X1 U7456 ( .A1(n5609), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5937) );
  OAI22_X1 U7457 ( .A1(n8135), .A2(n5941), .B1(n6239), .B2(n9714), .ZN(n5946)
         );
  INV_X1 U7458 ( .A(n5942), .ZN(n6150) );
  NAND2_X1 U7459 ( .A1(n8147), .A2(n9793), .ZN(n5943) );
  OAI211_X1 U7460 ( .C1(n9737), .C2(n6150), .A(n5944), .B(n5943), .ZN(n5945)
         );
  AOI211_X1 U7461 ( .C1(n5947), .C2(n9733), .A(n5946), .B(n5945), .ZN(n5948)
         );
  INV_X1 U7462 ( .A(n5948), .ZN(P2_U3241) );
  NAND2_X1 U7463 ( .A1(n5643), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U7464 ( .A(n5949), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7215) );
  INV_X1 U7465 ( .A(n7215), .ZN(n6999) );
  OAI222_X1 U7466 ( .A1(n8545), .A2(n5951), .B1(n4270), .B2(n5950), .C1(n6999), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U7467 ( .A1(n6053), .A2(n5954), .ZN(n5956) );
  AOI22_X1 U7468 ( .A1(n7339), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7338), .B2(
        n9756), .ZN(n5955) );
  XNOR2_X1 U7469 ( .A(n9800), .B(n8043), .ZN(n6314) );
  NOR2_X1 U7470 ( .A1(n6325), .A2(n6239), .ZN(n6313) );
  XNOR2_X1 U7471 ( .A(n6314), .B(n6313), .ZN(n6310) );
  XNOR2_X1 U7472 ( .A(n6309), .B(n6310), .ZN(n5968) );
  INV_X1 U7473 ( .A(n5957), .ZN(n6164) );
  INV_X1 U7474 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5958) );
  OAI22_X1 U7475 ( .A1(n9737), .A2(n6164), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5958), .ZN(n5966) );
  INV_X1 U7476 ( .A(n8156), .ZN(n6157) );
  NAND2_X1 U7477 ( .A1(n7320), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7478 ( .A1(n5595), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5963) );
  OAI21_X1 U7479 ( .B1(n5959), .B2(P2_REG3_REG_8__SCAN_IN), .A(n6340), .ZN(
        n9723) );
  INV_X1 U7480 ( .A(n9723), .ZN(n5960) );
  NAND2_X1 U7481 ( .A1(n7518), .A2(n5960), .ZN(n5962) );
  NAND2_X1 U7482 ( .A1(n5609), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5961) );
  OAI22_X1 U7483 ( .A1(n8135), .A2(n6157), .B1(n6663), .B2(n9714), .ZN(n5965)
         );
  AOI211_X1 U7484 ( .C1(n8147), .C2(n9800), .A(n5966), .B(n5965), .ZN(n5967)
         );
  OAI21_X1 U7485 ( .B1(n5968), .B2(n8128), .A(n5967), .ZN(P2_U3215) );
  INV_X1 U7486 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6271) );
  NOR2_X1 U7487 ( .A1(n5969), .A2(n6271), .ZN(n5973) );
  MUX2_X1 U7488 ( .A(n5970), .B(n7716), .S(n8041), .Z(n5971) );
  AOI21_X1 U7489 ( .B1(n8411), .B2(n5971), .A(n8128), .ZN(n5972) );
  AOI211_X1 U7490 ( .C1(n8147), .C2(n5108), .A(n5973), .B(n5972), .ZN(n5974)
         );
  OAI21_X1 U7491 ( .B1(n5975), .B2(n9714), .A(n5974), .ZN(P2_U3234) );
  INV_X1 U7492 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9435) );
  INV_X1 U7493 ( .A(n5976), .ZN(n5978) );
  NAND2_X1 U7494 ( .A1(n5978), .A2(n5977), .ZN(n5980) );
  OR2_X1 U7495 ( .A1(n5980), .A2(n5979), .ZN(n6079) );
  NAND2_X1 U7496 ( .A1(n9617), .A2(n4349), .ZN(n9619) );
  NOR2_X1 U7497 ( .A1(n5982), .A2(n5981), .ZN(n5983) );
  AND2_X1 U7498 ( .A1(n9617), .A2(n5983), .ZN(n9603) );
  OAI21_X1 U7499 ( .B1(n9132), .B2(n9603), .A(n5984), .ZN(n5988) );
  NOR2_X1 U7500 ( .A1(n9618), .A2(n5152), .ZN(n5985) );
  OAI21_X1 U7501 ( .B1(n5986), .B2(n5985), .A(n9617), .ZN(n5987) );
  OAI211_X1 U7502 ( .C1(n9435), .C2(n9617), .A(n5988), .B(n5987), .ZN(P1_U3291) );
  AND2_X1 U7503 ( .A1(n7989), .A2(n5989), .ZN(n9595) );
  NAND2_X1 U7504 ( .A1(n9617), .A2(n9595), .ZN(n9228) );
  INV_X1 U7505 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9429) );
  OAI22_X1 U7506 ( .A1(n9617), .A2(n5990), .B1(n9429), .B2(n9618), .ZN(n5993)
         );
  AND3_X1 U7507 ( .A1(n9603), .A2(n6433), .A3(n5991), .ZN(n5992) );
  AOI211_X1 U7508 ( .C1(n9132), .C2(n8682), .A(n5993), .B(n5992), .ZN(n5996)
         );
  NAND2_X1 U7509 ( .A1(n5994), .A2(n9617), .ZN(n5995) );
  OAI211_X1 U7510 ( .C1(n9228), .C2(n5997), .A(n5996), .B(n5995), .ZN(P1_U3290) );
  INV_X1 U7511 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6007) );
  INV_X1 U7512 ( .A(n5998), .ZN(n6001) );
  INV_X1 U7513 ( .A(n5999), .ZN(n6000) );
  MUX2_X1 U7514 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4276), .Z(n6126) );
  XNOR2_X1 U7515 ( .A(n6126), .B(SI_18_), .ZN(n6123) );
  XNOR2_X1 U7516 ( .A(n6125), .B(n6123), .ZN(n7808) );
  INV_X1 U7517 ( .A(n7808), .ZN(n6009) );
  NAND2_X1 U7518 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  NAND2_X1 U7519 ( .A1(n6005), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6006) );
  XNOR2_X1 U7520 ( .A(n6006), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9571) );
  INV_X1 U7521 ( .A(n9571), .ZN(n8966) );
  OAI222_X1 U7522 ( .A1(n9328), .A2(n6007), .B1(n8059), .B2(n6009), .C1(
        P1_U3084), .C2(n8966), .ZN(P1_U3335) );
  INV_X1 U7523 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7524 ( .A(n6008), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7312) );
  INV_X1 U7525 ( .A(n7312), .ZN(n8161) );
  OAI222_X1 U7526 ( .A1(n8545), .A2(n6010), .B1(n4270), .B2(n6009), .C1(
        P2_U3152), .C2(n8161), .ZN(P2_U3340) );
  AOI21_X1 U7527 ( .B1(n6013), .B2(n6012), .A(n6011), .ZN(n6290) );
  XNOR2_X1 U7528 ( .A(n6290), .B(n6300), .ZN(n6014) );
  NAND2_X1 U7529 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n6014), .ZN(n6291) );
  OAI211_X1 U7530 ( .C1(n6014), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9753), .B(
        n6291), .ZN(n6021) );
  OAI21_X1 U7531 ( .B1(n7010), .B2(P2_REG2_REG_14__SCAN_IN), .A(n6015), .ZN(
        n6299) );
  XNOR2_X1 U7532 ( .A(n6299), .B(n7067), .ZN(n6016) );
  INV_X1 U7533 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U7534 ( .A1(n6016), .A2(n9964), .ZN(n6301) );
  OAI21_X1 U7535 ( .B1(n6016), .B2(n9964), .A(n6301), .ZN(n6019) );
  AND2_X1 U7536 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7235) );
  AOI21_X1 U7537 ( .B1(n9747), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7235), .ZN(
        n6017) );
  OAI21_X1 U7538 ( .B1(n9739), .B2(n6300), .A(n6017), .ZN(n6018) );
  AOI21_X1 U7539 ( .B1(n6019), .B2(n9749), .A(n6018), .ZN(n6020) );
  NAND2_X1 U7540 ( .A1(n6021), .A2(n6020), .ZN(P2_U3260) );
  NAND2_X1 U7541 ( .A1(n6023), .A2(n6022), .ZN(n8684) );
  NAND2_X1 U7542 ( .A1(n6025), .A2(n6024), .ZN(n6027) );
  NAND2_X1 U7543 ( .A1(n8681), .A2(n8682), .ZN(n6026) );
  NAND2_X1 U7544 ( .A1(n6027), .A2(n6026), .ZN(n6428) );
  NAND2_X1 U7545 ( .A1(n6029), .A2(n6028), .ZN(n8688) );
  AND2_X2 U7546 ( .A1(n8688), .A2(n8684), .ZN(n8897) );
  NAND2_X1 U7547 ( .A1(n6428), .A2(n8897), .ZN(n6030) );
  NAND2_X1 U7548 ( .A1(n9641), .A2(n8953), .ZN(n8690) );
  NAND2_X1 U7549 ( .A1(n6414), .A2(n6031), .ZN(n8686) );
  NAND2_X1 U7550 ( .A1(n8690), .A2(n8686), .ZN(n6085) );
  INV_X1 U7551 ( .A(n6085), .ZN(n9607) );
  NAND2_X1 U7552 ( .A1(n9606), .A2(n9607), .ZN(n9605) );
  NAND2_X1 U7553 ( .A1(n9605), .A2(n8686), .ZN(n6413) );
  NAND2_X1 U7554 ( .A1(n9609), .A2(n6424), .ZN(n8693) );
  NAND2_X1 U7555 ( .A1(n9648), .A2(n8952), .ZN(n8691) );
  NAND2_X1 U7556 ( .A1(n8693), .A2(n8691), .ZN(n6088) );
  INV_X1 U7557 ( .A(n6088), .ZN(n8898) );
  NAND2_X1 U7558 ( .A1(n6413), .A2(n8898), .ZN(n6033) );
  NAND2_X1 U7559 ( .A1(n8686), .A2(n8693), .ZN(n6032) );
  NAND2_X1 U7560 ( .A1(n6032), .A2(n8691), .ZN(n8750) );
  NAND2_X1 U7561 ( .A1(n6033), .A2(n8750), .ZN(n9589) );
  OR2_X1 U7562 ( .A1(n8732), .A2(n6035), .ZN(n6036) );
  OAI211_X2 U7563 ( .C1(n5364), .C2(n6038), .A(n6037), .B(n6036), .ZN(n9584)
         );
  NAND2_X1 U7564 ( .A1(n6415), .A2(n9584), .ZN(n8692) );
  INV_X1 U7565 ( .A(n8692), .ZN(n6039) );
  OR2_X1 U7566 ( .A1(n8732), .A2(n6041), .ZN(n6042) );
  INV_X1 U7567 ( .A(n6512), .ZN(n9660) );
  NAND2_X1 U7568 ( .A1(n7983), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6052) );
  INV_X1 U7569 ( .A(n6047), .ZN(n6045) );
  NAND2_X1 U7570 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  AND2_X1 U7571 ( .A1(n6061), .A2(n6048), .ZN(n6511) );
  NAND2_X1 U7572 ( .A1(n5712), .A2(n6511), .ZN(n6051) );
  NAND2_X1 U7573 ( .A1(n7826), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7574 ( .A1(n8735), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7575 ( .A1(n9660), .A2(n8950), .ZN(n8754) );
  NAND2_X1 U7576 ( .A1(n9655), .A2(n8951), .ZN(n8752) );
  AND2_X1 U7577 ( .A1(n8754), .A2(n8752), .ZN(n8697) );
  NAND2_X1 U7578 ( .A1(n9593), .A2(n4264), .ZN(n8809) );
  INV_X2 U7579 ( .A(n5685), .ZN(n6363) );
  NAND2_X1 U7580 ( .A1(n6053), .A2(n6363), .ZN(n6058) );
  OR2_X1 U7581 ( .A1(n5364), .A2(n6054), .ZN(n6057) );
  OR2_X1 U7582 ( .A1(n8732), .A2(n6055), .ZN(n6056) );
  NAND2_X1 U7583 ( .A1(n7983), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6066) );
  INV_X1 U7584 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7585 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  AND2_X1 U7586 ( .A1(n6070), .A2(n6062), .ZN(n6202) );
  NAND2_X1 U7587 ( .A1(n5712), .A2(n6202), .ZN(n6065) );
  NAND2_X1 U7588 ( .A1(n7826), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7589 ( .A1(n8735), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6063) );
  NAND4_X1 U7590 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n8949)
         );
  NAND2_X1 U7591 ( .A1(n9668), .A2(n8949), .ZN(n8811) );
  INV_X1 U7592 ( .A(n8949), .ZN(n6361) );
  INV_X1 U7593 ( .A(n9668), .ZN(n6201) );
  NAND2_X1 U7594 ( .A1(n6361), .A2(n6201), .ZN(n8808) );
  NAND2_X1 U7595 ( .A1(n8811), .A2(n8808), .ZN(n6359) );
  INV_X1 U7596 ( .A(n6359), .ZN(n8902) );
  NAND3_X1 U7597 ( .A1(n6067), .A2(n8809), .A3(n6359), .ZN(n6068) );
  NAND2_X1 U7598 ( .A1(n6386), .A2(n6068), .ZN(n6076) );
  NAND2_X1 U7599 ( .A1(n7983), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6075) );
  INV_X1 U7600 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U7601 ( .A1(n6070), .A2(n6571), .ZN(n6071) );
  AND2_X1 U7602 ( .A1(n6373), .A2(n6071), .ZN(n6574) );
  NAND2_X1 U7603 ( .A1(n5712), .A2(n6574), .ZN(n6074) );
  NAND2_X1 U7604 ( .A1(n8735), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7605 ( .A1(n7826), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6072) );
  INV_X1 U7606 ( .A(n6588), .ZN(n8948) );
  AOI222_X1 U7607 ( .A1(n9612), .A2(n6076), .B1(n8948), .B2(n9357), .C1(n8950), 
        .C2(n9359), .ZN(n9667) );
  INV_X2 U7608 ( .A(n9617), .ZN(n9598) );
  INV_X1 U7609 ( .A(n6202), .ZN(n6077) );
  OAI22_X1 U7610 ( .A1(n9617), .A2(n6078), .B1(n6077), .B2(n9618), .ZN(n6081)
         );
  NAND2_X1 U7611 ( .A1(n9601), .A2(n9641), .ZN(n9600) );
  OR2_X2 U7612 ( .A1(n9600), .A2(n6424), .ZN(n9581) );
  OR2_X2 U7613 ( .A1(n9581), .A2(n9584), .ZN(n9582) );
  NOR2_X2 U7614 ( .A1(n9582), .A2(n4264), .ZN(n6508) );
  NAND2_X1 U7615 ( .A1(n6508), .A2(n9668), .ZN(n6404) );
  OAI211_X1 U7616 ( .C1(n6508), .C2(n9668), .A(n6404), .B(n9633), .ZN(n9666)
         );
  NOR2_X1 U7617 ( .A1(n6079), .A2(n9588), .ZN(n9209) );
  INV_X1 U7618 ( .A(n9209), .ZN(n6899) );
  NOR2_X1 U7619 ( .A1(n9666), .A2(n6899), .ZN(n6080) );
  AOI211_X1 U7620 ( .C1(n9132), .C2(n6201), .A(n6081), .B(n6080), .ZN(n6095)
         );
  NAND2_X1 U7621 ( .A1(n5462), .A2(n8682), .ZN(n6082) );
  NAND2_X1 U7622 ( .A1(n6023), .A2(n6028), .ZN(n6084) );
  NAND2_X1 U7623 ( .A1(n9599), .A2(n6085), .ZN(n6087) );
  NAND2_X1 U7624 ( .A1(n6414), .A2(n9641), .ZN(n6086) );
  NAND2_X1 U7625 ( .A1(n6087), .A2(n6086), .ZN(n6412) );
  NAND2_X1 U7626 ( .A1(n6412), .A2(n6088), .ZN(n6090) );
  NAND2_X1 U7627 ( .A1(n9609), .A2(n9648), .ZN(n6089) );
  AND2_X1 U7628 ( .A1(n8692), .A2(n8752), .ZN(n8900) );
  OAI22_X1 U7629 ( .A1(n9580), .A2(n8900), .B1(n6415), .B2(n9655), .ZN(n6506)
         );
  INV_X1 U7630 ( .A(n6506), .ZN(n6092) );
  INV_X1 U7631 ( .A(n8904), .ZN(n6091) );
  NAND2_X1 U7632 ( .A1(n6092), .A2(n6091), .ZN(n6505) );
  NAND2_X1 U7633 ( .A1(n9593), .A2(n9660), .ZN(n6093) );
  NAND2_X1 U7634 ( .A1(n6505), .A2(n6093), .ZN(n6360) );
  XNOR2_X1 U7635 ( .A(n6360), .B(n6359), .ZN(n9670) );
  INV_X1 U7636 ( .A(n9228), .ZN(n9171) );
  NAND2_X1 U7637 ( .A1(n9670), .A2(n9171), .ZN(n6094) );
  OAI211_X1 U7638 ( .C1(n9667), .C2(n9598), .A(n6095), .B(n6094), .ZN(P1_U3284) );
  NAND3_X1 U7639 ( .A1(n6098), .A2(n6097), .A3(n6096), .ZN(n6099) );
  NAND2_X1 U7640 ( .A1(n6149), .A2(n8389), .ZN(n6958) );
  INV_X2 U7641 ( .A(n6958), .ZN(n8402) );
  INV_X1 U7642 ( .A(n6149), .ZN(n6101) );
  NAND2_X1 U7643 ( .A1(n6101), .A2(n8236), .ZN(n6526) );
  INV_X1 U7644 ( .A(n6526), .ZN(n6115) );
  INV_X1 U7645 ( .A(n8389), .ZN(n8408) );
  AOI22_X1 U7646 ( .A1(n6115), .A2(n6102), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8408), .ZN(n6104) );
  NAND2_X1 U7647 ( .A1(n8402), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6103) );
  OAI211_X1 U7648 ( .C1(n6105), .C2(n8402), .A(n6104), .B(n6103), .ZN(n6112)
         );
  INV_X1 U7649 ( .A(n7181), .ZN(n6107) );
  NOR2_X1 U7650 ( .A1(n6106), .A2(n8236), .ZN(n6261) );
  OAI21_X2 U7651 ( .B1(n6107), .B2(n6261), .A(n8422), .ZN(n8399) );
  AND2_X1 U7652 ( .A1(n5617), .A2(n7744), .ZN(n6108) );
  NAND2_X1 U7653 ( .A1(n8422), .A2(n6108), .ZN(n8368) );
  OAI22_X1 U7654 ( .A1(n6110), .A2(n8399), .B1(n6109), .B2(n8368), .ZN(n6111)
         );
  OR2_X1 U7655 ( .A1(n6112), .A2(n6111), .ZN(P2_U3294) );
  INV_X1 U7656 ( .A(n8399), .ZN(n8407) );
  OAI22_X1 U7657 ( .A1(n5234), .A2(n8422), .B1(n6113), .B2(n8389), .ZN(n6114)
         );
  AOI21_X1 U7658 ( .B1(n6116), .B2(n6115), .A(n6114), .ZN(n6117) );
  OAI21_X1 U7659 ( .B1(n6118), .B2(n8368), .A(n6117), .ZN(n6119) );
  AOI21_X1 U7660 ( .B1(n8407), .B2(n6120), .A(n6119), .ZN(n6121) );
  OAI21_X1 U7661 ( .B1(n6122), .B2(n8402), .A(n6121), .ZN(P2_U3292) );
  INV_X1 U7662 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6132) );
  INV_X1 U7663 ( .A(n6123), .ZN(n6124) );
  NAND2_X1 U7664 ( .A1(n6126), .A2(SI_18_), .ZN(n6127) );
  INV_X1 U7665 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6134) );
  MUX2_X1 U7666 ( .A(n6132), .B(n6134), .S(n7537), .Z(n6129) );
  INV_X1 U7667 ( .A(SI_19_), .ZN(n9937) );
  NAND2_X1 U7668 ( .A1(n6129), .A2(n9937), .ZN(n6352) );
  INV_X1 U7669 ( .A(n6129), .ZN(n6130) );
  NAND2_X1 U7670 ( .A1(n6130), .A2(SI_19_), .ZN(n6131) );
  NAND2_X1 U7671 ( .A1(n6352), .A2(n6131), .ZN(n6353) );
  XNOR2_X1 U7672 ( .A(n6354), .B(n6353), .ZN(n7821) );
  INV_X1 U7673 ( .A(n7821), .ZN(n6133) );
  OAI222_X1 U7674 ( .A1(n8545), .A2(n6132), .B1(n4270), .B2(n6133), .C1(
        P2_U3152), .C2(n8236), .ZN(P2_U3339) );
  OAI222_X1 U7675 ( .A1(n9328), .A2(n6134), .B1(n8059), .B2(n6133), .C1(n9128), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OR2_X1 U7676 ( .A1(n8157), .A2(n9790), .ZN(n7569) );
  INV_X1 U7677 ( .A(n9790), .ZN(n6218) );
  OR2_X1 U7678 ( .A1(n8157), .A2(n6218), .ZN(n6137) );
  NAND2_X1 U7679 ( .A1(n6138), .A2(n6137), .ZN(n6156) );
  XNOR2_X1 U7680 ( .A(n8156), .B(n9793), .ZN(n7721) );
  XNOR2_X1 U7681 ( .A(n6156), .B(n7721), .ZN(n9797) );
  INV_X1 U7682 ( .A(n7568), .ZN(n6139) );
  NOR2_X1 U7683 ( .A1(n6140), .A2(n6139), .ZN(n6141) );
  NAND2_X1 U7684 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  OAI21_X1 U7685 ( .B1(n7721), .B2(n6145), .A(n6230), .ZN(n6148) );
  NAND2_X1 U7686 ( .A1(n8157), .A2(n8419), .ZN(n6146) );
  OAI21_X1 U7687 ( .B1(n6239), .B2(n8330), .A(n6146), .ZN(n6147) );
  AOI21_X1 U7688 ( .B1(n6148), .B2(n8414), .A(n6147), .ZN(n9796) );
  MUX2_X1 U7689 ( .A(n5231), .B(n9796), .S(n8422), .Z(n6153) );
  AOI21_X1 U7690 ( .B1(n9793), .B2(n6215), .A(n6162), .ZN(n9794) );
  NOR2_X2 U7691 ( .A1(n6149), .A2(n8041), .ZN(n8409) );
  INV_X1 U7692 ( .A(n9793), .ZN(n7584) );
  OAI22_X1 U7693 ( .A1(n8368), .A2(n7584), .B1(n8389), .B2(n6150), .ZN(n6151)
         );
  AOI21_X1 U7694 ( .B1(n9794), .B2(n8409), .A(n6151), .ZN(n6152) );
  OAI211_X1 U7695 ( .C1(n8399), .C2(n9797), .A(n6153), .B(n6152), .ZN(P2_U3290) );
  NOR2_X1 U7696 ( .A1(n8156), .A2(n9793), .ZN(n6155) );
  NAND2_X1 U7697 ( .A1(n8156), .A2(n9793), .ZN(n6154) );
  OAI21_X1 U7698 ( .B1(n6156), .B2(n6155), .A(n6154), .ZN(n6223) );
  NAND2_X1 U7699 ( .A1(n9800), .A2(n6239), .ZN(n7598) );
  XNOR2_X1 U7700 ( .A(n6223), .B(n6229), .ZN(n9805) );
  NAND2_X1 U7701 ( .A1(n6230), .A2(n4296), .ZN(n6158) );
  XNOR2_X1 U7702 ( .A(n6158), .B(n7722), .ZN(n6161) );
  NAND2_X1 U7703 ( .A1(n8156), .A2(n8419), .ZN(n6159) );
  OAI21_X1 U7704 ( .B1(n6663), .B2(n8330), .A(n6159), .ZN(n6160) );
  AOI21_X1 U7705 ( .B1(n6161), .B2(n8414), .A(n6160), .ZN(n9803) );
  MUX2_X1 U7706 ( .A(n5229), .B(n9803), .S(n8422), .Z(n6168) );
  INV_X1 U7707 ( .A(n6162), .ZN(n6163) );
  INV_X1 U7708 ( .A(n9800), .ZN(n6165) );
  AND2_X1 U7709 ( .A1(n6162), .A2(n6165), .ZN(n6244) );
  AOI21_X1 U7710 ( .B1(n9800), .B2(n6163), .A(n6244), .ZN(n9801) );
  OAI22_X1 U7711 ( .A1(n8368), .A2(n6165), .B1(n8389), .B2(n6164), .ZN(n6166)
         );
  AOI21_X1 U7712 ( .B1(n9801), .B2(n8409), .A(n6166), .ZN(n6167) );
  OAI211_X1 U7713 ( .C1(n8399), .C2(n9805), .A(n6168), .B(n6167), .ZN(P2_U3289) );
  NAND2_X1 U7714 ( .A1(n4265), .A2(n8949), .ZN(n6169) );
  OAI21_X1 U7715 ( .B1(n9668), .B2(n7900), .A(n6169), .ZN(n6170) );
  XNOR2_X1 U7716 ( .A(n6170), .B(n8009), .ZN(n6554) );
  NAND2_X1 U7717 ( .A1(n7974), .A2(n8949), .ZN(n6172) );
  OR2_X1 U7718 ( .A1(n9668), .A2(n6180), .ZN(n6171) );
  NAND2_X1 U7719 ( .A1(n6172), .A2(n6171), .ZN(n6552) );
  XNOR2_X1 U7720 ( .A(n6554), .B(n6552), .ZN(n6199) );
  INV_X1 U7721 ( .A(n6173), .ZN(n6175) );
  NAND2_X1 U7722 ( .A1(n6175), .A2(n6174), .ZN(n6176) );
  OR2_X1 U7723 ( .A1(n6415), .A2(n6180), .ZN(n6178) );
  OAI21_X1 U7724 ( .B1(n9655), .B2(n7900), .A(n6178), .ZN(n6179) );
  XNOR2_X1 U7725 ( .A(n6179), .B(n8009), .ZN(n6192) );
  NAND2_X1 U7726 ( .A1(n7974), .A2(n8951), .ZN(n6182) );
  NAND2_X1 U7727 ( .A1(n4265), .A2(n9584), .ZN(n6181) );
  AND2_X1 U7728 ( .A1(n6182), .A2(n6181), .ZN(n6254) );
  AND2_X1 U7729 ( .A1(n6192), .A2(n6254), .ZN(n6196) );
  OR2_X1 U7730 ( .A1(n9593), .A2(n6180), .ZN(n6183) );
  OAI21_X1 U7731 ( .B1(n9660), .B2(n7900), .A(n6183), .ZN(n6184) );
  XNOR2_X1 U7732 ( .A(n6184), .B(n8009), .ZN(n6187) );
  NAND2_X1 U7733 ( .A1(n7974), .A2(n8950), .ZN(n6186) );
  NAND2_X1 U7734 ( .A1(n4265), .A2(n4264), .ZN(n6185) );
  AND2_X1 U7735 ( .A1(n6186), .A2(n6185), .ZN(n6188) );
  NAND2_X1 U7736 ( .A1(n6187), .A2(n6188), .ZN(n6197) );
  INV_X1 U7737 ( .A(n6187), .ZN(n6190) );
  INV_X1 U7738 ( .A(n6188), .ZN(n6189) );
  NAND2_X1 U7739 ( .A1(n6190), .A2(n6189), .ZN(n6191) );
  NAND2_X1 U7740 ( .A1(n6197), .A2(n6191), .ZN(n6279) );
  INV_X1 U7741 ( .A(n6192), .ZN(n6252) );
  INV_X1 U7742 ( .A(n6254), .ZN(n6193) );
  AND2_X1 U7743 ( .A1(n6252), .A2(n6193), .ZN(n6194) );
  NAND2_X1 U7744 ( .A1(n6198), .A2(n6199), .ZN(n6556) );
  OAI21_X1 U7745 ( .B1(n6199), .B2(n6198), .A(n6556), .ZN(n6208) );
  INV_X1 U7746 ( .A(n8656), .ZN(n8633) );
  AOI21_X1 U7747 ( .B1(n8633), .B2(n8950), .A(n6200), .ZN(n6206) );
  NAND2_X1 U7748 ( .A1(n8648), .A2(n6201), .ZN(n6205) );
  NAND2_X1 U7749 ( .A1(n8660), .A2(n6202), .ZN(n6204) );
  NAND2_X1 U7750 ( .A1(n8644), .A2(n8948), .ZN(n6203) );
  NAND4_X1 U7751 ( .A1(n6206), .A2(n6205), .A3(n6204), .A4(n6203), .ZN(n6207)
         );
  AOI21_X1 U7752 ( .B1(n6208), .B2(n8652), .A(n6207), .ZN(n6209) );
  INV_X1 U7753 ( .A(n6209), .ZN(P1_U3211) );
  XNOR2_X1 U7754 ( .A(n6210), .B(n7718), .ZN(n9792) );
  INV_X1 U7755 ( .A(n9792), .ZN(n6221) );
  XNOR2_X1 U7756 ( .A(n6211), .B(n7718), .ZN(n6214) );
  NAND2_X1 U7757 ( .A1(n8158), .A2(n8419), .ZN(n6213) );
  NAND2_X1 U7758 ( .A1(n8156), .A2(n8417), .ZN(n6212) );
  NAND2_X1 U7759 ( .A1(n6213), .A2(n6212), .ZN(n9728) );
  AOI21_X1 U7760 ( .B1(n6214), .B2(n8414), .A(n9728), .ZN(n9789) );
  INV_X1 U7761 ( .A(n9789), .ZN(n6217) );
  OAI211_X1 U7762 ( .C1(n4355), .C2(n9790), .A(n9810), .B(n6215), .ZN(n9788)
         );
  OAI22_X1 U7763 ( .A1(n9788), .A2(n8253), .B1(n8389), .B2(n9736), .ZN(n6216)
         );
  OAI21_X1 U7764 ( .B1(n6217), .B2(n6216), .A(n8422), .ZN(n6220) );
  INV_X1 U7765 ( .A(n8368), .ZN(n8406) );
  AOI22_X1 U7766 ( .A1(n8406), .A2(n6218), .B1(n8402), .B2(
        P2_REG2_REG_5__SCAN_IN), .ZN(n6219) );
  OAI211_X1 U7767 ( .C1(n6221), .C2(n8399), .A(n6220), .B(n6219), .ZN(P2_U3291) );
  INV_X1 U7768 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6249) );
  INV_X1 U7769 ( .A(n6239), .ZN(n9716) );
  NAND2_X1 U7770 ( .A1(n6364), .A2(n5954), .ZN(n6226) );
  AOI22_X1 U7771 ( .A1(n7339), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7338), .B2(
        n6224), .ZN(n6225) );
  NAND2_X1 U7772 ( .A1(n6226), .A2(n6225), .ZN(n6529) );
  OR2_X1 U7773 ( .A1(n6529), .A2(n6663), .ZN(n7602) );
  NAND2_X1 U7774 ( .A1(n6529), .A2(n6663), .ZN(n7603) );
  NAND2_X1 U7775 ( .A1(n7602), .A2(n7603), .ZN(n6233) );
  NAND2_X1 U7776 ( .A1(n6227), .A2(n4266), .ZN(n6228) );
  NAND2_X1 U7777 ( .A1(n6530), .A2(n6228), .ZN(n6268) );
  OR2_X1 U7778 ( .A1(n6268), .A2(n7181), .ZN(n6243) );
  NAND2_X1 U7779 ( .A1(n6231), .A2(n7597), .ZN(n6232) );
  NAND2_X1 U7780 ( .A1(n6232), .A2(n6233), .ZN(n6234) );
  NAND2_X1 U7781 ( .A1(n6523), .A2(n6234), .ZN(n6241) );
  NAND2_X1 U7782 ( .A1(n5609), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7783 ( .A1(n7320), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6237) );
  XNOR2_X1 U7784 ( .A(n6340), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7785 ( .A1(n7518), .A2(n6336), .ZN(n6236) );
  NAND2_X1 U7786 ( .A1(n5595), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6235) );
  OAI22_X1 U7787 ( .A1(n6239), .A2(n8328), .B1(n9713), .B2(n8330), .ZN(n6240)
         );
  AOI21_X1 U7788 ( .B1(n6241), .B2(n8414), .A(n6240), .ZN(n6242) );
  NAND2_X1 U7789 ( .A1(n6243), .A2(n6242), .ZN(n6262) );
  INV_X1 U7790 ( .A(n6262), .ZN(n6247) );
  INV_X1 U7791 ( .A(n6529), .ZN(n9719) );
  OR2_X1 U7792 ( .A1(n6244), .A2(n9719), .ZN(n6245) );
  AND2_X1 U7793 ( .A1(n6669), .A2(n6245), .ZN(n6265) );
  AOI22_X1 U7794 ( .A1(n6265), .A2(n9810), .B1(n9809), .B2(n6529), .ZN(n6246)
         );
  OAI211_X1 U7795 ( .C1(n9814), .C2(n6268), .A(n6247), .B(n6246), .ZN(n6250)
         );
  NAND2_X1 U7796 ( .A1(n6250), .A2(n4267), .ZN(n6248) );
  OAI21_X1 U7797 ( .B1(n4267), .B2(n6249), .A(n6248), .ZN(P2_U3475) );
  NAND2_X1 U7798 ( .A1(n6250), .A2(n4268), .ZN(n6251) );
  OAI21_X1 U7799 ( .B1(n4268), .B2(n5202), .A(n6251), .ZN(P2_U3528) );
  INV_X1 U7800 ( .A(n9585), .ZN(n6260) );
  NOR2_X1 U7801 ( .A1(n4350), .A2(n6252), .ZN(n6277) );
  AOI21_X1 U7802 ( .B1(n4350), .B2(n6252), .A(n6277), .ZN(n6253) );
  NAND2_X1 U7803 ( .A1(n6253), .A2(n6254), .ZN(n6280) );
  OAI21_X1 U7804 ( .B1(n6254), .B2(n6253), .A(n6280), .ZN(n6255) );
  NAND2_X1 U7805 ( .A1(n6255), .A2(n8652), .ZN(n6259) );
  OAI22_X1 U7806 ( .A1(n8663), .A2(n9655), .B1(n8657), .B2(n9593), .ZN(n6256)
         );
  AOI211_X1 U7807 ( .C1(n8633), .C2(n8952), .A(n6257), .B(n6256), .ZN(n6258)
         );
  OAI211_X1 U7808 ( .C1(n8646), .C2(n6260), .A(n6259), .B(n6258), .ZN(P1_U3225) );
  AND2_X1 U7809 ( .A1(n8422), .A2(n6261), .ZN(n7202) );
  INV_X1 U7810 ( .A(n7202), .ZN(n6968) );
  MUX2_X1 U7811 ( .A(n6262), .B(P2_REG2_REG_8__SCAN_IN), .S(n8402), .Z(n6263)
         );
  INV_X1 U7812 ( .A(n6263), .ZN(n6267) );
  OAI22_X1 U7813 ( .A1(n8368), .A2(n9719), .B1(n8389), .B2(n9723), .ZN(n6264)
         );
  AOI21_X1 U7814 ( .B1(n6265), .B2(n8409), .A(n6264), .ZN(n6266) );
  OAI211_X1 U7815 ( .C1(n6268), .C2(n6968), .A(n6267), .B(n6266), .ZN(P2_U3288) );
  INV_X1 U7816 ( .A(n6269), .ZN(n6276) );
  OAI21_X1 U7817 ( .B1(n6271), .B2(n8389), .A(n6270), .ZN(n6273) );
  INV_X1 U7818 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9742) );
  NOR2_X1 U7819 ( .A1(n8422), .A2(n9742), .ZN(n6272) );
  AOI21_X1 U7820 ( .B1(n8422), .B2(n6273), .A(n6272), .ZN(n6275) );
  OAI21_X1 U7821 ( .B1(n8406), .B2(n8409), .A(n5108), .ZN(n6274) );
  OAI211_X1 U7822 ( .C1(n6276), .C2(n8399), .A(n6275), .B(n6274), .ZN(P2_U3296) );
  INV_X1 U7823 ( .A(n6277), .ZN(n6278) );
  NAND3_X1 U7824 ( .A1(n6280), .A2(n6279), .A3(n6278), .ZN(n6282) );
  AOI21_X1 U7825 ( .B1(n6282), .B2(n6281), .A(n8650), .ZN(n6289) );
  AOI21_X1 U7826 ( .B1(n8633), .B2(n8951), .A(n6283), .ZN(n6287) );
  NAND2_X1 U7827 ( .A1(n8660), .A2(n6511), .ZN(n6286) );
  NAND2_X1 U7828 ( .A1(n8648), .A2(n4264), .ZN(n6285) );
  NAND2_X1 U7829 ( .A1(n8644), .A2(n8949), .ZN(n6284) );
  NAND4_X1 U7830 ( .A1(n6287), .A2(n6286), .A3(n6285), .A4(n6284), .ZN(n6288)
         );
  OR2_X1 U7831 ( .A1(n6289), .A2(n6288), .ZN(P1_U3237) );
  NAND2_X1 U7832 ( .A1(n7067), .A2(n6290), .ZN(n6292) );
  NAND2_X1 U7833 ( .A1(n6292), .A2(n6291), .ZN(n6295) );
  OR2_X1 U7834 ( .A1(n7176), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U7835 ( .A1(n7176), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7836 ( .A1(n6459), .A2(n6293), .ZN(n6294) );
  NOR2_X1 U7837 ( .A1(n6295), .A2(n6294), .ZN(n6461) );
  AOI21_X1 U7838 ( .B1(n6295), .B2(n6294), .A(n6461), .ZN(n6308) );
  INV_X1 U7839 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6297) );
  INV_X1 U7840 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7078) );
  NOR2_X1 U7841 ( .A1(n7078), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8108) );
  INV_X1 U7842 ( .A(n8108), .ZN(n6296) );
  OAI21_X1 U7843 ( .B1(n6298), .B2(n6297), .A(n6296), .ZN(n6306) );
  NAND2_X1 U7844 ( .A1(n6300), .A2(n6299), .ZN(n6302) );
  NAND2_X1 U7845 ( .A1(n6302), .A2(n6301), .ZN(n6304) );
  XNOR2_X1 U7846 ( .A(n7176), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n6303) );
  NOR2_X1 U7847 ( .A1(n6304), .A2(n6303), .ZN(n6464) );
  AOI211_X1 U7848 ( .C1(n6304), .C2(n6303), .A(n6466), .B(n6464), .ZN(n6305)
         );
  AOI211_X1 U7849 ( .C1(n9757), .C2(n7176), .A(n6306), .B(n6305), .ZN(n6307)
         );
  OAI21_X1 U7850 ( .B1(n6308), .B2(n9740), .A(n6307), .ZN(P2_U3261) );
  INV_X1 U7851 ( .A(n6309), .ZN(n6312) );
  INV_X1 U7852 ( .A(n6310), .ZN(n6311) );
  NAND2_X1 U7853 ( .A1(n6312), .A2(n6311), .ZN(n6316) );
  NAND2_X1 U7854 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  NAND2_X1 U7855 ( .A1(n6316), .A2(n6315), .ZN(n9710) );
  XNOR2_X1 U7856 ( .A(n6529), .B(n7439), .ZN(n6317) );
  NOR2_X1 U7857 ( .A1(n6325), .A2(n6663), .ZN(n6318) );
  XNOR2_X1 U7858 ( .A(n6317), .B(n6318), .ZN(n9711) );
  NAND2_X1 U7859 ( .A1(n9710), .A2(n9711), .ZN(n6321) );
  INV_X1 U7860 ( .A(n6317), .ZN(n6319) );
  NAND2_X1 U7861 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  NAND2_X1 U7862 ( .A1(n6321), .A2(n6320), .ZN(n6331) );
  NAND2_X1 U7863 ( .A1(n6369), .A2(n5954), .ZN(n6324) );
  AOI22_X1 U7864 ( .A1(n7339), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7338), .B2(
        n6322), .ZN(n6323) );
  XNOR2_X1 U7865 ( .A(n9808), .B(n7439), .ZN(n6326) );
  OR2_X1 U7866 ( .A1(n6325), .A2(n9713), .ZN(n6327) );
  NAND2_X1 U7867 ( .A1(n6326), .A2(n6327), .ZN(n6473) );
  INV_X1 U7868 ( .A(n6326), .ZN(n6329) );
  INV_X1 U7869 ( .A(n6327), .ZN(n6328) );
  NAND2_X1 U7870 ( .A1(n6329), .A2(n6328), .ZN(n6330) );
  NAND2_X1 U7871 ( .A1(n6473), .A2(n6330), .ZN(n6335) );
  INV_X1 U7872 ( .A(n6331), .ZN(n6333) );
  NAND2_X1 U7873 ( .A1(n6333), .A2(n6332), .ZN(n6474) );
  INV_X1 U7874 ( .A(n6474), .ZN(n6334) );
  AOI21_X1 U7875 ( .B1(n6331), .B2(n6335), .A(n6334), .ZN(n6351) );
  INV_X1 U7876 ( .A(n6336), .ZN(n6670) );
  OAI21_X1 U7877 ( .B1(n9737), .B2(n6670), .A(n6337), .ZN(n6349) );
  NAND2_X1 U7878 ( .A1(n7320), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U7879 ( .A1(n5609), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6346) );
  INV_X1 U7880 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6339) );
  INV_X1 U7881 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U7882 ( .B1(n6340), .B2(n6339), .A(n6338), .ZN(n6343) );
  INV_X1 U7883 ( .A(n6340), .ZN(n6342) );
  AND2_X1 U7884 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n6341) );
  NAND2_X1 U7885 ( .A1(n6342), .A2(n6341), .ZN(n6486) );
  NAND2_X1 U7886 ( .A1(n6343), .A2(n6486), .ZN(n9709) );
  INV_X1 U7887 ( .A(n9709), .ZN(n6546) );
  NAND2_X1 U7888 ( .A1(n7518), .A2(n6546), .ZN(n6345) );
  NAND2_X1 U7889 ( .A1(n5595), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6344) );
  OAI22_X1 U7890 ( .A1(n8135), .A2(n6663), .B1(n6662), .B2(n9714), .ZN(n6348)
         );
  AOI211_X1 U7891 ( .C1(n8147), .C2(n9808), .A(n6349), .B(n6348), .ZN(n6350)
         );
  OAI21_X1 U7892 ( .B1(n6351), .B2(n8128), .A(n6350), .ZN(P2_U3233) );
  INV_X1 U7893 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7348) );
  INV_X1 U7894 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7845) );
  MUX2_X1 U7895 ( .A(n7348), .B(n7845), .S(n7537), .Z(n6355) );
  INV_X1 U7896 ( .A(SI_20_), .ZN(n9941) );
  NAND2_X1 U7897 ( .A1(n6355), .A2(n9941), .ZN(n6457) );
  INV_X1 U7898 ( .A(n6355), .ZN(n6356) );
  NAND2_X1 U7899 ( .A1(n6356), .A2(SI_20_), .ZN(n6357) );
  AND2_X1 U7900 ( .A1(n6457), .A2(n6357), .ZN(n6455) );
  XNOR2_X1 U7901 ( .A(n6456), .B(n6455), .ZN(n7844) );
  INV_X1 U7902 ( .A(n7844), .ZN(n6394) );
  OAI222_X1 U7903 ( .A1(n8545), .A2(n7348), .B1(n4270), .B2(n6394), .C1(n6358), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NAND2_X1 U7904 ( .A1(n9668), .A2(n6361), .ZN(n6362) );
  NAND2_X1 U7905 ( .A1(n6364), .A2(n6363), .ZN(n6366) );
  AOI22_X1 U7906 ( .A1(n7823), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7822), .B2(
        n9447), .ZN(n6365) );
  OR2_X1 U7907 ( .A1(n6562), .A2(n6588), .ZN(n8701) );
  NAND2_X1 U7908 ( .A1(n6562), .A2(n6588), .ZN(n8675) );
  NAND2_X1 U7909 ( .A1(n6562), .A2(n8948), .ZN(n6368) );
  NAND2_X1 U7910 ( .A1(n6396), .A2(n6368), .ZN(n6594) );
  NAND2_X1 U7911 ( .A1(n6369), .A2(n6363), .ZN(n6371) );
  AOI22_X1 U7912 ( .A1(n7823), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7822), .B2(
        n9467), .ZN(n6370) );
  INV_X1 U7913 ( .A(n6595), .ZN(n9679) );
  NAND2_X1 U7914 ( .A1(n7983), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6378) );
  INV_X1 U7915 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U7916 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  AND2_X1 U7917 ( .A1(n6380), .A2(n6374), .ZN(n6590) );
  NAND2_X1 U7918 ( .A1(n5712), .A2(n6590), .ZN(n6377) );
  NAND2_X1 U7919 ( .A1(n7826), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U7920 ( .A1(n8735), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6375) );
  NAND4_X1 U7921 ( .A1(n6378), .A2(n6377), .A3(n6376), .A4(n6375), .ZN(n8947)
         );
  AND2_X1 U7922 ( .A1(n9679), .A2(n8947), .ZN(n8814) );
  INV_X1 U7923 ( .A(n8947), .ZN(n6695) );
  NAND2_X1 U7924 ( .A1(n6595), .A2(n6695), .ZN(n6642) );
  INV_X1 U7925 ( .A(n6642), .ZN(n8817) );
  OR2_X1 U7926 ( .A1(n8814), .A2(n8817), .ZN(n8905) );
  INV_X1 U7927 ( .A(n8905), .ZN(n6379) );
  XNOR2_X1 U7928 ( .A(n6594), .B(n6379), .ZN(n9685) );
  INV_X1 U7929 ( .A(n9685), .ZN(n6393) );
  INV_X1 U7930 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U7931 ( .A1(n6380), .A2(n6693), .ZN(n6381) );
  AND2_X1 U7932 ( .A1(n6608), .A2(n6381), .ZN(n6697) );
  NAND2_X1 U7933 ( .A1(n5712), .A2(n6697), .ZN(n6385) );
  NAND2_X1 U7934 ( .A1(n7983), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U7935 ( .A1(n8735), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U7936 ( .A1(n7826), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U7937 ( .A1(n6386), .A2(n8808), .ZN(n6399) );
  INV_X1 U7938 ( .A(n8675), .ZN(n8816) );
  XOR2_X1 U7939 ( .A(n6625), .B(n8905), .Z(n6387) );
  OAI222_X1 U7940 ( .A1(n9610), .A2(n6678), .B1(n9608), .B2(n6588), .C1(n9591), 
        .C2(n6387), .ZN(n9682) );
  INV_X1 U7941 ( .A(n6646), .ZN(n6388) );
  OAI21_X1 U7942 ( .B1(n9679), .B2(n4473), .A(n6388), .ZN(n9681) );
  INV_X1 U7943 ( .A(n9603), .ZN(n9000) );
  INV_X1 U7944 ( .A(n9618), .ZN(n9586) );
  AOI22_X1 U7945 ( .A1(n9598), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6590), .B2(
        n9586), .ZN(n6390) );
  NAND2_X1 U7946 ( .A1(n9132), .A2(n6595), .ZN(n6389) );
  OAI211_X1 U7947 ( .C1(n9681), .C2(n9000), .A(n6390), .B(n6389), .ZN(n6391)
         );
  AOI21_X1 U7948 ( .B1(n9682), .B2(n9617), .A(n6391), .ZN(n6392) );
  OAI21_X1 U7949 ( .B1(n9228), .B2(n6393), .A(n6392), .ZN(P1_U3282) );
  OAI222_X1 U7950 ( .A1(n9328), .A2(n7845), .B1(P1_U3084), .B2(n6395), .C1(
        n8059), .C2(n6394), .ZN(P1_U3333) );
  NAND2_X1 U7951 ( .A1(n6397), .A2(n8903), .ZN(n6398) );
  NAND2_X1 U7952 ( .A1(n6396), .A2(n6398), .ZN(n6403) );
  AOI22_X1 U7953 ( .A1(n9359), .A2(n8949), .B1(n9357), .B2(n8947), .ZN(n6402)
         );
  XNOR2_X1 U7954 ( .A(n6399), .B(n8903), .ZN(n6400) );
  NAND2_X1 U7955 ( .A1(n6400), .A2(n9612), .ZN(n6401) );
  OAI211_X1 U7956 ( .C1(n6403), .C2(n9615), .A(n6402), .B(n6401), .ZN(n9674)
         );
  INV_X1 U7957 ( .A(n9674), .ZN(n6411) );
  INV_X1 U7958 ( .A(n6403), .ZN(n9676) );
  NOR3_X1 U7959 ( .A1(n9598), .A2(n5359), .A3(n9128), .ZN(n9604) );
  NAND2_X1 U7960 ( .A1(n6404), .A2(n6562), .ZN(n6405) );
  NAND2_X1 U7961 ( .A1(n6406), .A2(n6405), .ZN(n9673) );
  AOI22_X1 U7962 ( .A1(n9598), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6574), .B2(
        n9586), .ZN(n6408) );
  NAND2_X1 U7963 ( .A1(n9132), .A2(n6562), .ZN(n6407) );
  OAI211_X1 U7964 ( .C1(n9673), .C2(n9000), .A(n6408), .B(n6407), .ZN(n6409)
         );
  AOI21_X1 U7965 ( .B1(n9676), .B2(n9604), .A(n6409), .ZN(n6410) );
  OAI21_X1 U7966 ( .B1(n6411), .B2(n9598), .A(n6410), .ZN(P1_U3283) );
  XNOR2_X1 U7967 ( .A(n6412), .B(n8898), .ZN(n9647) );
  INV_X1 U7968 ( .A(n9604), .ZN(n6439) );
  XNOR2_X1 U7969 ( .A(n6413), .B(n8898), .ZN(n6417) );
  OAI22_X1 U7970 ( .A1(n9610), .A2(n6415), .B1(n6414), .B2(n9608), .ZN(n6416)
         );
  AOI21_X1 U7971 ( .B1(n6417), .B2(n9612), .A(n6416), .ZN(n6418) );
  OAI21_X1 U7972 ( .B1(n9647), .B2(n9615), .A(n6418), .ZN(n9650) );
  NAND2_X1 U7973 ( .A1(n9650), .A2(n9617), .ZN(n6426) );
  OAI22_X1 U7974 ( .A1(n9617), .A2(n6420), .B1(n6419), .B2(n9618), .ZN(n6423)
         );
  INV_X1 U7975 ( .A(n9600), .ZN(n6421) );
  OAI21_X1 U7976 ( .B1(n6421), .B2(n9648), .A(n9581), .ZN(n9649) );
  NOR2_X1 U7977 ( .A1(n9649), .A2(n9000), .ZN(n6422) );
  AOI211_X1 U7978 ( .C1(n9132), .C2(n6424), .A(n6423), .B(n6422), .ZN(n6425)
         );
  OAI211_X1 U7979 ( .C1(n9647), .C2(n6439), .A(n6426), .B(n6425), .ZN(P1_U3287) );
  XNOR2_X1 U7980 ( .A(n6427), .B(n8897), .ZN(n6432) );
  INV_X1 U7981 ( .A(n6432), .ZN(n9637) );
  INV_X1 U7982 ( .A(n9615), .ZN(n9363) );
  INV_X1 U7983 ( .A(n6428), .ZN(n8685) );
  XNOR2_X1 U7984 ( .A(n8685), .B(n8897), .ZN(n6430) );
  AOI22_X1 U7985 ( .A1(n9359), .A2(n5462), .B1(n9357), .B2(n8953), .ZN(n6429)
         );
  OAI21_X1 U7986 ( .B1(n6430), .B2(n9591), .A(n6429), .ZN(n6431) );
  AOI21_X1 U7987 ( .B1(n6432), .B2(n9363), .A(n6431), .ZN(n9636) );
  MUX2_X1 U7988 ( .A(n5433), .B(n9636), .S(n9617), .Z(n6438) );
  AND2_X1 U7989 ( .A1(n6433), .A2(n6022), .ZN(n6434) );
  NOR2_X1 U7990 ( .A1(n9601), .A2(n6434), .ZN(n9634) );
  INV_X1 U7991 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6435) );
  OAI22_X1 U7992 ( .A1(n9619), .A2(n6028), .B1(n6435), .B2(n9618), .ZN(n6436)
         );
  AOI21_X1 U7993 ( .B1(n9603), .B2(n9634), .A(n6436), .ZN(n6437) );
  OAI211_X1 U7994 ( .C1(n9637), .C2(n6439), .A(n6438), .B(n6437), .ZN(P1_U3289) );
  OAI21_X1 U7995 ( .B1(n6441), .B2(n7719), .A(n6440), .ZN(n9785) );
  INV_X1 U7996 ( .A(n9785), .ZN(n6454) );
  OAI22_X1 U7997 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n8389), .B1(n8422), .B2(
        n6442), .ZN(n6447) );
  INV_X1 U7998 ( .A(n8409), .ZN(n8295) );
  INV_X1 U7999 ( .A(n6443), .ZN(n6445) );
  OAI21_X1 U8000 ( .B1(n9780), .B2(n6445), .A(n6444), .ZN(n9782) );
  NOR2_X1 U8001 ( .A1(n8295), .A2(n9782), .ZN(n6446) );
  AOI211_X1 U8002 ( .C1(n8406), .C2(n5853), .A(n6447), .B(n6446), .ZN(n6453)
         );
  AOI22_X1 U8003 ( .A1(n8419), .A2(n8418), .B1(n8158), .B2(n8417), .ZN(n6451)
         );
  OAI21_X1 U8004 ( .B1(n7576), .B2(n6448), .A(n6142), .ZN(n6449) );
  NAND2_X1 U8005 ( .A1(n6449), .A2(n8414), .ZN(n6450) );
  OAI211_X1 U8006 ( .C1(n6454), .C2(n7181), .A(n6451), .B(n6450), .ZN(n9783)
         );
  NAND2_X1 U8007 ( .A1(n9783), .A2(n8422), .ZN(n6452) );
  OAI211_X1 U8008 ( .C1(n6454), .C2(n6968), .A(n6453), .B(n6452), .ZN(P2_U3293) );
  INV_X1 U8009 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7357) );
  INV_X1 U8010 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7865) );
  MUX2_X1 U8011 ( .A(n7357), .B(n7865), .S(n7537), .Z(n6713) );
  XNOR2_X1 U8012 ( .A(n6713), .B(SI_21_), .ZN(n6711) );
  INV_X1 U8013 ( .A(n7864), .ZN(n6521) );
  OAI222_X1 U8014 ( .A1(n8545), .A2(n7357), .B1(n4270), .B2(n6521), .C1(n7747), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U8015 ( .A(n6459), .ZN(n6460) );
  NOR2_X1 U8016 ( .A1(n6461), .A2(n6460), .ZN(n6997) );
  XNOR2_X1 U8017 ( .A(n7215), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n6995) );
  XNOR2_X1 U8018 ( .A(n6997), .B(n6995), .ZN(n6471) );
  INV_X1 U8019 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7218) );
  NOR2_X1 U8020 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7218), .ZN(n6462) );
  AOI21_X1 U8021 ( .B1(n9747), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n6462), .ZN(
        n6463) );
  OAI21_X1 U8022 ( .B1(n9739), .B2(n6999), .A(n6463), .ZN(n6470) );
  AOI21_X1 U8023 ( .B1(n7176), .B2(P2_REG2_REG_16__SCAN_IN), .A(n6464), .ZN(
        n6468) );
  NAND2_X1 U8024 ( .A1(n7215), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6465) );
  OAI21_X1 U8025 ( .B1(n7215), .B2(P2_REG2_REG_17__SCAN_IN), .A(n6465), .ZN(
        n6467) );
  NOR2_X1 U8026 ( .A1(n6468), .A2(n6467), .ZN(n6989) );
  AOI211_X1 U8027 ( .C1(n6468), .C2(n6467), .A(n6466), .B(n6989), .ZN(n6469)
         );
  AOI211_X1 U8028 ( .C1(n6471), .C2(n9753), .A(n6470), .B(n6469), .ZN(n6472)
         );
  INV_X1 U8029 ( .A(n6472), .ZN(P2_U3262) );
  NAND2_X1 U8030 ( .A1(n6598), .A2(n5954), .ZN(n6477) );
  AOI22_X1 U8031 ( .A1(n7339), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7338), .B2(
        n6475), .ZN(n6476) );
  XNOR2_X1 U8032 ( .A(n6911), .B(n8043), .ZN(n6478) );
  NOR2_X1 U8033 ( .A1(n6325), .A2(n6662), .ZN(n6479) );
  XNOR2_X1 U8034 ( .A(n6478), .B(n6479), .ZN(n9700) );
  INV_X1 U8035 ( .A(n6478), .ZN(n6481) );
  INV_X1 U8036 ( .A(n6479), .ZN(n6480) );
  NAND2_X1 U8037 ( .A1(n6603), .A2(n5954), .ZN(n6484) );
  AOI22_X1 U8038 ( .A1(n7339), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7338), .B2(
        n6482), .ZN(n6483) );
  XNOR2_X1 U8039 ( .A(n6731), .B(n7439), .ZN(n6794) );
  NAND2_X1 U8040 ( .A1(n7320), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U8041 ( .A1(n5595), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6490) );
  INV_X1 U8042 ( .A(n6486), .ZN(n6485) );
  NAND2_X1 U8043 ( .A1(n6485), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U8044 ( .A1(n6486), .A2(n6493), .ZN(n6487) );
  AND2_X1 U8045 ( .A1(n6495), .A2(n6487), .ZN(n6492) );
  NAND2_X1 U8046 ( .A1(n7518), .A2(n6492), .ZN(n6489) );
  NAND2_X1 U8047 ( .A1(n5609), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6488) );
  NOR2_X1 U8048 ( .A1(n6325), .A2(n9702), .ZN(n6795) );
  XNOR2_X1 U8049 ( .A(n6794), .B(n6795), .ZN(n6792) );
  XNOR2_X1 U8050 ( .A(n6793), .B(n6792), .ZN(n6504) );
  INV_X1 U8051 ( .A(n6492), .ZN(n6525) );
  OAI22_X1 U8052 ( .A1(n9737), .A2(n6525), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6493), .ZN(n6502) );
  NAND2_X1 U8053 ( .A1(n7320), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U8054 ( .A1(n5609), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6499) );
  INV_X1 U8055 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6494) );
  NAND2_X1 U8056 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  AND2_X1 U8057 ( .A1(n6745), .A2(n6496), .ZN(n6803) );
  NAND2_X1 U8058 ( .A1(n7518), .A2(n6803), .ZN(n6498) );
  NAND2_X1 U8059 ( .A1(n5595), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6497) );
  OAI22_X1 U8060 ( .A1(n8135), .A2(n6662), .B1(n6844), .B2(n9714), .ZN(n6501)
         );
  AOI211_X1 U8061 ( .C1(n8147), .C2(n6731), .A(n6502), .B(n6501), .ZN(n6503)
         );
  OAI21_X1 U8062 ( .B1(n6504), .B2(n8128), .A(n6503), .ZN(P2_U3238) );
  NAND2_X1 U8063 ( .A1(n6506), .A2(n8904), .ZN(n6507) );
  NAND2_X1 U8064 ( .A1(n6505), .A2(n6507), .ZN(n9664) );
  INV_X1 U8065 ( .A(n6508), .ZN(n6510) );
  NAND2_X1 U8066 ( .A1(n9582), .A2(n4264), .ZN(n6509) );
  NAND2_X1 U8067 ( .A1(n6510), .A2(n6509), .ZN(n9661) );
  AOI22_X1 U8068 ( .A1(n9132), .A2(n4264), .B1(n6511), .B2(n9586), .ZN(n6513)
         );
  OAI21_X1 U8069 ( .B1(n9661), .B2(n9000), .A(n6513), .ZN(n6519) );
  NAND2_X1 U8070 ( .A1(n6514), .A2(n8752), .ZN(n8788) );
  XNOR2_X1 U8071 ( .A(n8788), .B(n8904), .ZN(n6517) );
  NAND2_X1 U8072 ( .A1(n9664), .A2(n9363), .ZN(n6516) );
  AOI22_X1 U8073 ( .A1(n9359), .A2(n8951), .B1(n9357), .B2(n8949), .ZN(n6515)
         );
  OAI211_X1 U8074 ( .C1(n9591), .C2(n6517), .A(n6516), .B(n6515), .ZN(n9662)
         );
  MUX2_X1 U8075 ( .A(n9662), .B(P1_REG2_REG_6__SCAN_IN), .S(n9598), .Z(n6518)
         );
  AOI211_X1 U8076 ( .C1(n9604), .C2(n9664), .A(n6519), .B(n6518), .ZN(n6520)
         );
  INV_X1 U8077 ( .A(n6520), .ZN(P1_U3285) );
  OAI222_X1 U8078 ( .A1(n9328), .A2(n7865), .B1(P1_U3084), .B2(n6522), .C1(
        n8059), .C2(n6521), .ZN(P1_U3332) );
  OR2_X1 U8079 ( .A1(n9808), .A2(n9713), .ZN(n7560) );
  NAND2_X1 U8080 ( .A1(n9808), .A2(n9713), .ZN(n7605) );
  OR2_X1 U8081 ( .A1(n6911), .A2(n6662), .ZN(n7559) );
  NAND2_X1 U8082 ( .A1(n6911), .A2(n6662), .ZN(n7561) );
  OR2_X1 U8083 ( .A1(n6731), .A2(n9702), .ZN(n7610) );
  NAND2_X1 U8084 ( .A1(n6731), .A2(n9702), .ZN(n7609) );
  NAND2_X1 U8085 ( .A1(n7610), .A2(n7609), .ZN(n7727) );
  XOR2_X1 U8086 ( .A(n6742), .B(n7727), .Z(n6524) );
  INV_X1 U8087 ( .A(n6844), .ZN(n8152) );
  INV_X1 U8088 ( .A(n6662), .ZN(n8154) );
  AOI222_X1 U8089 ( .A1(n8384), .A2(n6524), .B1(n8152), .B2(n8417), .C1(n8154), 
        .C2(n8419), .ZN(n9819) );
  OAI22_X1 U8090 ( .A1(n8422), .A2(n5403), .B1(n6525), .B2(n8389), .ZN(n6528)
         );
  INV_X1 U8091 ( .A(n6731), .ZN(n9821) );
  INV_X1 U8092 ( .A(n6737), .ZN(n6739) );
  OAI211_X1 U8093 ( .C1(n9821), .C2(n4353), .A(n6739), .B(n9810), .ZN(n9818)
         );
  NOR2_X1 U8094 ( .A1(n9818), .A2(n6526), .ZN(n6527) );
  AOI211_X1 U8095 ( .C1(n8406), .C2(n6731), .A(n6528), .B(n6527), .ZN(n6536)
         );
  INV_X1 U8096 ( .A(n6663), .ZN(n8155) );
  INV_X1 U8097 ( .A(n6659), .ZN(n6532) );
  INV_X1 U8098 ( .A(n9713), .ZN(n9704) );
  OR2_X1 U8099 ( .A1(n9808), .A2(n9704), .ZN(n6533) );
  NAND2_X1 U8100 ( .A1(n7559), .A2(n7561), .ZN(n7726) );
  NAND2_X1 U8101 ( .A1(n6911), .A2(n8154), .ZN(n6534) );
  XOR2_X1 U8102 ( .A(n6730), .B(n7727), .Z(n9824) );
  NAND2_X1 U8103 ( .A1(n9824), .A2(n8407), .ZN(n6535) );
  OAI211_X1 U8104 ( .C1(n9819), .C2(n8402), .A(n6536), .B(n6535), .ZN(P2_U3285) );
  XNOR2_X1 U8105 ( .A(n6537), .B(n6538), .ZN(n6544) );
  OAI22_X1 U8106 ( .A1(n9713), .A2(n8328), .B1(n9702), .B2(n8330), .ZN(n6543)
         );
  NAND2_X1 U8107 ( .A1(n6539), .A2(n6538), .ZN(n6540) );
  NAND2_X1 U8108 ( .A1(n6541), .A2(n6540), .ZN(n6916) );
  NOR2_X1 U8109 ( .A1(n6916), .A2(n7181), .ZN(n6542) );
  AOI211_X1 U8110 ( .C1(n6544), .C2(n8414), .A(n6543), .B(n6542), .ZN(n6915)
         );
  INV_X1 U8111 ( .A(n6916), .ZN(n6550) );
  AND2_X1 U8112 ( .A1(n6667), .A2(n6911), .ZN(n6545) );
  OR2_X1 U8113 ( .A1(n6545), .A2(n4353), .ZN(n6912) );
  AOI22_X1 U8114 ( .A1(n8402), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n6546), .B2(
        n8408), .ZN(n6548) );
  NAND2_X1 U8115 ( .A1(n8406), .A2(n6911), .ZN(n6547) );
  OAI211_X1 U8116 ( .C1(n6912), .C2(n8295), .A(n6548), .B(n6547), .ZN(n6549)
         );
  AOI21_X1 U8117 ( .B1(n6550), .B2(n7202), .A(n6549), .ZN(n6551) );
  OAI21_X1 U8118 ( .B1(n6915), .B2(n8402), .A(n6551), .ZN(P2_U3286) );
  INV_X1 U8119 ( .A(n6562), .ZN(n9672) );
  INV_X1 U8120 ( .A(n6552), .ZN(n6553) );
  NAND2_X1 U8121 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  INV_X1 U8122 ( .A(n6557), .ZN(n6560) );
  NAND2_X1 U8123 ( .A1(n7974), .A2(n8948), .ZN(n6559) );
  NAND2_X1 U8124 ( .A1(n6562), .A2(n4265), .ZN(n6558) );
  NAND2_X1 U8125 ( .A1(n6559), .A2(n6558), .ZN(n6682) );
  NOR2_X1 U8126 ( .A1(n6560), .A2(n6682), .ZN(n6568) );
  NAND2_X1 U8127 ( .A1(n6562), .A2(n7995), .ZN(n6564) );
  OR2_X1 U8128 ( .A1(n6588), .A2(n6180), .ZN(n6563) );
  NAND2_X1 U8129 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  XNOR2_X1 U8130 ( .A(n6565), .B(n7989), .ZN(n6683) );
  INV_X1 U8131 ( .A(n6683), .ZN(n6567) );
  NOR2_X1 U8132 ( .A1(n6568), .A2(n6567), .ZN(n6584) );
  INV_X1 U8133 ( .A(n6584), .ZN(n6570) );
  INV_X1 U8134 ( .A(n6682), .ZN(n6566) );
  NOR2_X1 U8135 ( .A1(n6557), .A2(n6566), .ZN(n6583) );
  OAI21_X1 U8136 ( .B1(n6568), .B2(n6583), .A(n6567), .ZN(n6569) );
  OAI211_X1 U8137 ( .C1(n6570), .C2(n6583), .A(n8652), .B(n6569), .ZN(n6576)
         );
  NAND2_X1 U8138 ( .A1(n8633), .A2(n8949), .ZN(n6572) );
  OR2_X1 U8139 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6571), .ZN(n9450) );
  OAI211_X1 U8140 ( .C1(n6695), .C2(n8657), .A(n6572), .B(n9450), .ZN(n6573)
         );
  AOI21_X1 U8141 ( .B1(n6574), .B2(n8660), .A(n6573), .ZN(n6575) );
  OAI211_X1 U8142 ( .C1(n9672), .C2(n8663), .A(n6576), .B(n6575), .ZN(P1_U3219) );
  NAND2_X1 U8143 ( .A1(n6595), .A2(n7995), .ZN(n6578) );
  NAND2_X1 U8144 ( .A1(n4265), .A2(n8947), .ZN(n6577) );
  NAND2_X1 U8145 ( .A1(n6578), .A2(n6577), .ZN(n6579) );
  XNOR2_X1 U8146 ( .A(n6579), .B(n8009), .ZN(n6581) );
  AOI22_X1 U8147 ( .A1(n6595), .A2(n4265), .B1(n7974), .B2(n8947), .ZN(n6580)
         );
  NAND2_X1 U8148 ( .A1(n6581), .A2(n6580), .ZN(n6681) );
  NAND2_X1 U8149 ( .A1(n6681), .A2(n6685), .ZN(n6582) );
  NOR3_X1 U8150 ( .A1(n6584), .A2(n6583), .A3(n6582), .ZN(n6680) );
  OAI21_X1 U8151 ( .B1(n6584), .B2(n6583), .A(n6582), .ZN(n6585) );
  INV_X1 U8152 ( .A(n6585), .ZN(n6586) );
  OAI21_X1 U8153 ( .B1(n6680), .B2(n6586), .A(n8652), .ZN(n6592) );
  INV_X1 U8154 ( .A(n6678), .ZN(n9358) );
  AND2_X1 U8155 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9466) );
  AOI21_X1 U8156 ( .B1(n8644), .B2(n9358), .A(n9466), .ZN(n6587) );
  OAI21_X1 U8157 ( .B1(n6588), .B2(n8656), .A(n6587), .ZN(n6589) );
  AOI21_X1 U8158 ( .B1(n6590), .B2(n8660), .A(n6589), .ZN(n6591) );
  OAI211_X1 U8159 ( .C1(n9679), .C2(n8663), .A(n6592), .B(n6591), .ZN(P1_U3229) );
  OR2_X1 U8160 ( .A1(n6595), .A2(n8947), .ZN(n6593) );
  NAND2_X1 U8161 ( .A1(n6594), .A2(n6593), .ZN(n6597) );
  NAND2_X1 U8162 ( .A1(n6595), .A2(n8947), .ZN(n6596) );
  NAND2_X1 U8163 ( .A1(n6597), .A2(n6596), .ZN(n6650) );
  NAND2_X1 U8164 ( .A1(n6598), .A2(n6363), .ZN(n6600) );
  AOI22_X1 U8165 ( .A1(n7823), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7822), .B2(
        n9479), .ZN(n6599) );
  NAND2_X1 U8166 ( .A1(n6600), .A2(n6599), .ZN(n6702) );
  OR2_X1 U8167 ( .A1(n6702), .A2(n6678), .ZN(n8815) );
  NAND2_X1 U8168 ( .A1(n6702), .A2(n6678), .ZN(n8820) );
  OR2_X1 U8169 ( .A1(n6702), .A2(n9358), .ZN(n6602) );
  NAND2_X1 U8170 ( .A1(n6603), .A2(n6363), .ZN(n6605) );
  AOI22_X1 U8171 ( .A1(n7823), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7822), .B2(
        n8970), .ZN(n6604) );
  NAND2_X1 U8172 ( .A1(n7983), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6613) );
  INV_X1 U8173 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U8174 ( .A1(n6608), .A2(n6607), .ZN(n6609) );
  AND2_X1 U8175 ( .A1(n6618), .A2(n6609), .ZN(n9364) );
  NAND2_X1 U8176 ( .A1(n5712), .A2(n9364), .ZN(n6612) );
  NAND2_X1 U8177 ( .A1(n7826), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U8178 ( .A1(n8735), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6610) );
  NAND4_X1 U8179 ( .A1(n6613), .A2(n6612), .A3(n6611), .A4(n6610), .ZN(n8946)
         );
  NAND2_X1 U8180 ( .A1(n6824), .A2(n8946), .ZN(n8823) );
  OR2_X1 U8181 ( .A1(n6824), .A2(n8946), .ZN(n8824) );
  NAND2_X1 U8182 ( .A1(n6733), .A2(n6363), .ZN(n6616) );
  AOI22_X1 U8183 ( .A1(n7823), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7822), .B2(
        n9493), .ZN(n6615) );
  NAND2_X1 U8184 ( .A1(n7826), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6623) );
  NAND2_X1 U8185 ( .A1(n7983), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6622) );
  INV_X1 U8186 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U8187 ( .A1(n6618), .A2(n6868), .ZN(n6619) );
  AND2_X1 U8188 ( .A1(n6628), .A2(n6619), .ZN(n6867) );
  NAND2_X1 U8189 ( .A1(n5712), .A2(n6867), .ZN(n6621) );
  NAND2_X1 U8190 ( .A1(n8735), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U8191 ( .A1(n6876), .A2(n6982), .ZN(n8819) );
  INV_X1 U8192 ( .A(n8908), .ZN(n6624) );
  XNOR2_X1 U8193 ( .A(n6877), .B(n6624), .ZN(n9404) );
  AND2_X1 U8194 ( .A1(n8820), .A2(n6642), .ZN(n8793) );
  INV_X1 U8195 ( .A(n8946), .ZN(n6814) );
  NAND2_X1 U8196 ( .A1(n6824), .A2(n6814), .ZN(n8671) );
  NAND2_X1 U8197 ( .A1(n9354), .A2(n8671), .ZN(n6626) );
  OR2_X1 U8198 ( .A1(n6824), .A2(n6814), .ZN(n8703) );
  NAND2_X1 U8199 ( .A1(n6626), .A2(n8703), .ZN(n6881) );
  XNOR2_X1 U8200 ( .A(n6881), .B(n8908), .ZN(n6635) );
  NAND2_X1 U8201 ( .A1(n7826), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U8202 ( .A1(n7983), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6632) );
  INV_X1 U8203 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U8204 ( .A1(n6628), .A2(n6627), .ZN(n6629) );
  AND2_X1 U8205 ( .A1(n6885), .A2(n6629), .ZN(n6979) );
  NAND2_X1 U8206 ( .A1(n5712), .A2(n6979), .ZN(n6631) );
  NAND2_X1 U8207 ( .A1(n8735), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6630) );
  INV_X1 U8208 ( .A(n7144), .ZN(n8945) );
  AOI22_X1 U8209 ( .A1(n9359), .A2(n8946), .B1(n9357), .B2(n8945), .ZN(n6634)
         );
  OAI21_X1 U8210 ( .B1(n6635), .B2(n9591), .A(n6634), .ZN(n6636) );
  AOI21_X1 U8211 ( .B1(n9404), .B2(n9363), .A(n6636), .ZN(n9406) );
  INV_X1 U8212 ( .A(n6702), .ZN(n6700) );
  INV_X1 U8213 ( .A(n6824), .ZN(n9408) );
  AOI21_X1 U8214 ( .B1(n9352), .B2(n6876), .A(n9680), .ZN(n6637) );
  NAND2_X1 U8215 ( .A1(n6637), .A2(n6895), .ZN(n9402) );
  AOI22_X1 U8216 ( .A1(n9598), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n6867), .B2(
        n9586), .ZN(n6639) );
  NAND2_X1 U8217 ( .A1(n6876), .A2(n9132), .ZN(n6638) );
  OAI211_X1 U8218 ( .C1(n9402), .C2(n6899), .A(n6639), .B(n6638), .ZN(n6640)
         );
  AOI21_X1 U8219 ( .B1(n9404), .B2(n9604), .A(n6640), .ZN(n6641) );
  OAI21_X1 U8220 ( .B1(n9406), .B2(n9598), .A(n6641), .ZN(P1_U3279) );
  NAND2_X1 U8221 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  XNOR2_X1 U8222 ( .A(n6644), .B(n8896), .ZN(n6645) );
  AOI222_X1 U8223 ( .A1(n9612), .A2(n6645), .B1(n8947), .B2(n9359), .C1(n8946), 
        .C2(n9357), .ZN(n6704) );
  OAI21_X1 U8224 ( .B1(n6646), .B2(n6700), .A(n9633), .ZN(n6647) );
  NOR2_X1 U8225 ( .A1(n6647), .A2(n9350), .ZN(n6701) );
  NAND2_X1 U8226 ( .A1(n9598), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U8227 ( .A1(n9586), .A2(n6697), .ZN(n6648) );
  OAI211_X1 U8228 ( .C1(n6700), .C2(n9619), .A(n6649), .B(n6648), .ZN(n6655)
         );
  INV_X1 U8229 ( .A(n6652), .ZN(n6653) );
  AOI21_X1 U8230 ( .B1(n8896), .B2(n6651), .A(n6653), .ZN(n6705) );
  NOR2_X1 U8231 ( .A1(n6705), .A2(n9228), .ZN(n6654) );
  AOI211_X1 U8232 ( .C1(n6701), .C2(n9209), .A(n6655), .B(n6654), .ZN(n6656)
         );
  OAI21_X1 U8233 ( .B1(n9598), .B2(n6704), .A(n6656), .ZN(P1_U3281) );
  INV_X1 U8234 ( .A(n6657), .ZN(n6658) );
  AOI21_X1 U8235 ( .B1(n7724), .B2(n6659), .A(n6658), .ZN(n9815) );
  OAI21_X1 U8236 ( .B1(n7724), .B2(n6661), .A(n6660), .ZN(n6666) );
  OAI22_X1 U8237 ( .A1(n6663), .A2(n8328), .B1(n6662), .B2(n8330), .ZN(n6665)
         );
  NOR2_X1 U8238 ( .A1(n9815), .A2(n7181), .ZN(n6664) );
  AOI211_X1 U8239 ( .C1(n8384), .C2(n6666), .A(n6665), .B(n6664), .ZN(n9813)
         );
  MUX2_X1 U8240 ( .A(n5241), .B(n9813), .S(n8422), .Z(n6674) );
  INV_X1 U8241 ( .A(n6667), .ZN(n6668) );
  AOI21_X1 U8242 ( .B1(n9808), .B2(n6669), .A(n6668), .ZN(n9811) );
  INV_X1 U8243 ( .A(n9808), .ZN(n6671) );
  OAI22_X1 U8244 ( .A1(n8368), .A2(n6671), .B1(n8389), .B2(n6670), .ZN(n6672)
         );
  AOI21_X1 U8245 ( .B1(n9811), .B2(n8409), .A(n6672), .ZN(n6673) );
  OAI211_X1 U8246 ( .C1(n9815), .C2(n6968), .A(n6674), .B(n6673), .ZN(P2_U3287) );
  NAND2_X1 U8247 ( .A1(n6702), .A2(n7995), .ZN(n6676) );
  OR2_X1 U8248 ( .A1(n6678), .A2(n6180), .ZN(n6675) );
  NAND2_X1 U8249 ( .A1(n6676), .A2(n6675), .ZN(n6677) );
  XNOR2_X1 U8250 ( .A(n6677), .B(n7989), .ZN(n6816) );
  NOR2_X1 U8251 ( .A1(n8012), .A2(n6678), .ZN(n6679) );
  AOI21_X1 U8252 ( .B1(n6702), .B2(n4265), .A(n6679), .ZN(n6817) );
  XNOR2_X1 U8253 ( .A(n6816), .B(n6817), .ZN(n6687) );
  INV_X1 U8254 ( .A(n6681), .ZN(n6686) );
  NOR3_X1 U8255 ( .A1(n6680), .A2(n6687), .A3(n6686), .ZN(n6692) );
  OAI21_X1 U8256 ( .B1(n6683), .B2(n6682), .A(n6681), .ZN(n6690) );
  NAND2_X1 U8257 ( .A1(n6683), .A2(n6682), .ZN(n6684) );
  INV_X1 U8258 ( .A(n6819), .ZN(n6691) );
  OAI21_X1 U8259 ( .B1(n6692), .B2(n6691), .A(n8652), .ZN(n6699) );
  NOR2_X1 U8260 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6693), .ZN(n9478) );
  AOI21_X1 U8261 ( .B1(n8644), .B2(n8946), .A(n9478), .ZN(n6694) );
  OAI21_X1 U8262 ( .B1(n6695), .B2(n8656), .A(n6694), .ZN(n6696) );
  AOI21_X1 U8263 ( .B1(n6697), .B2(n8660), .A(n6696), .ZN(n6698) );
  OAI211_X1 U8264 ( .C1(n6700), .C2(n8663), .A(n6699), .B(n6698), .ZN(P1_U3215) );
  INV_X1 U8265 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6707) );
  INV_X1 U8266 ( .A(n9684), .ZN(n9375) );
  AOI21_X1 U8267 ( .B1(n9632), .B2(n6702), .A(n6701), .ZN(n6703) );
  OAI211_X1 U8268 ( .C1(n6705), .C2(n9375), .A(n6704), .B(n6703), .ZN(n6708)
         );
  NAND2_X1 U8269 ( .A1(n6708), .A2(n10017), .ZN(n6706) );
  OAI21_X1 U8270 ( .B1(n10017), .B2(n6707), .A(n6706), .ZN(P1_U3484) );
  NAND2_X1 U8271 ( .A1(n6708), .A2(n4269), .ZN(n6709) );
  OAI21_X1 U8272 ( .B1(n4269), .B2(n5289), .A(n6709), .ZN(P1_U3533) );
  INV_X1 U8273 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7907) );
  INV_X1 U8274 ( .A(n6710), .ZN(n6712) );
  NAND2_X1 U8275 ( .A1(n6712), .A2(n6711), .ZN(n6716) );
  INV_X1 U8276 ( .A(n6713), .ZN(n6714) );
  NAND2_X1 U8277 ( .A1(n6714), .A2(SI_21_), .ZN(n6715) );
  INV_X1 U8278 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7377) );
  INV_X1 U8279 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8039) );
  MUX2_X1 U8280 ( .A(n7377), .B(n8039), .S(n4276), .Z(n6718) );
  INV_X1 U8281 ( .A(SI_22_), .ZN(n6717) );
  NAND2_X1 U8282 ( .A1(n6718), .A2(n6717), .ZN(n6721) );
  INV_X1 U8283 ( .A(n6718), .ZN(n6719) );
  NAND2_X1 U8284 ( .A1(n6719), .A2(SI_22_), .ZN(n6720) );
  NAND2_X1 U8285 ( .A1(n6721), .A2(n6720), .ZN(n7329) );
  INV_X1 U8286 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7394) );
  MUX2_X1 U8287 ( .A(n7394), .B(n7907), .S(n7537), .Z(n6723) );
  INV_X1 U8288 ( .A(SI_23_), .ZN(n6722) );
  NAND2_X1 U8289 ( .A1(n6723), .A2(n6722), .ZN(n6924) );
  INV_X1 U8290 ( .A(n6723), .ZN(n6724) );
  NAND2_X1 U8291 ( .A1(n6724), .A2(SI_23_), .ZN(n6725) );
  AND2_X1 U8292 ( .A1(n6924), .A2(n6725), .ZN(n6922) );
  NAND2_X1 U8293 ( .A1(n7906), .A2(n9323), .ZN(n6727) );
  NAND2_X1 U8294 ( .A1(n6726), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8938) );
  OAI211_X1 U8295 ( .C1(n7907), .C2(n9328), .A(n6727), .B(n8938), .ZN(P1_U3330) );
  NAND2_X1 U8296 ( .A1(n7906), .A2(n6728), .ZN(n6729) );
  OAI211_X1 U8297 ( .C1(n7394), .C2(n8545), .A(n6729), .B(n7760), .ZN(P2_U3335) );
  INV_X1 U8298 ( .A(n9702), .ZN(n8153) );
  NAND2_X1 U8299 ( .A1(n6731), .A2(n8153), .ZN(n6732) );
  NAND2_X1 U8300 ( .A1(n6733), .A2(n5954), .ZN(n6736) );
  AOI22_X1 U8301 ( .A1(n7339), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7338), .B2(
        n6734), .ZN(n6735) );
  OR2_X1 U8302 ( .A1(n6950), .A2(n6844), .ZN(n7617) );
  XOR2_X1 U8303 ( .A(n6951), .B(n7729), .Z(n6905) );
  INV_X1 U8304 ( .A(n6950), .ZN(n6741) );
  NAND2_X1 U8305 ( .A1(n6737), .A2(n6741), .ZN(n6959) );
  INV_X1 U8306 ( .A(n6959), .ZN(n6738) );
  AOI21_X1 U8307 ( .B1(n6950), .B2(n6739), .A(n6738), .ZN(n6902) );
  AOI22_X1 U8308 ( .A1(n8402), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n6803), .B2(
        n8408), .ZN(n6740) );
  OAI21_X1 U8309 ( .B1(n6741), .B2(n8368), .A(n6740), .ZN(n6755) );
  NAND2_X1 U8310 ( .A1(n6742), .A2(n7610), .ZN(n6743) );
  NAND2_X1 U8311 ( .A1(n6743), .A2(n7609), .ZN(n6954) );
  XNOR2_X1 U8312 ( .A(n6954), .B(n7729), .ZN(n6753) );
  NAND2_X1 U8313 ( .A1(n5609), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6750) );
  NAND2_X1 U8314 ( .A1(n7320), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6749) );
  INV_X1 U8315 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U8316 ( .A1(n6745), .A2(n6744), .ZN(n6746) );
  AND2_X1 U8317 ( .A1(n6838), .A2(n6746), .ZN(n6961) );
  NAND2_X1 U8318 ( .A1(n7518), .A2(n6961), .ZN(n6748) );
  NAND2_X1 U8319 ( .A1(n5595), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6747) );
  OR2_X1 U8320 ( .A1(n7046), .A2(n8330), .ZN(n6752) );
  OR2_X1 U8321 ( .A1(n9702), .A2(n8328), .ZN(n6751) );
  NAND2_X1 U8322 ( .A1(n6752), .A2(n6751), .ZN(n6804) );
  AOI21_X1 U8323 ( .B1(n6753), .B2(n8384), .A(n6804), .ZN(n6904) );
  NOR2_X1 U8324 ( .A1(n6904), .A2(n8402), .ZN(n6754) );
  AOI211_X1 U8325 ( .C1(n6902), .C2(n8409), .A(n6755), .B(n6754), .ZN(n6756)
         );
  OAI21_X1 U8326 ( .B1(n8399), .B2(n6905), .A(n6756), .ZN(P2_U3284) );
  INV_X1 U8327 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10026) );
  NOR2_X1 U8328 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6757) );
  AOI21_X1 U8329 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6757), .ZN(n9841) );
  NOR2_X1 U8330 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6758) );
  AOI21_X1 U8331 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6758), .ZN(n9844) );
  NOR2_X1 U8332 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6759) );
  AOI21_X1 U8333 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6759), .ZN(n9847) );
  NOR2_X1 U8334 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6760) );
  AOI21_X1 U8335 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6760), .ZN(n9850) );
  NOR2_X1 U8336 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6761) );
  AOI21_X1 U8337 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6761), .ZN(n9853) );
  NOR2_X1 U8338 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6767) );
  XNOR2_X1 U8339 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10039) );
  NAND2_X1 U8340 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6765) );
  XOR2_X1 U8341 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10037) );
  NAND2_X1 U8342 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n6763) );
  XOR2_X1 U8343 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10035) );
  AOI21_X1 U8344 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9835) );
  NAND3_X1 U8345 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9837) );
  OAI21_X1 U8346 ( .B1(n9835), .B2(n5314), .A(n9837), .ZN(n10034) );
  NAND2_X1 U8347 ( .A1(n10035), .A2(n10034), .ZN(n6762) );
  NAND2_X1 U8348 ( .A1(n6763), .A2(n6762), .ZN(n10036) );
  NAND2_X1 U8349 ( .A1(n10037), .A2(n10036), .ZN(n6764) );
  NAND2_X1 U8350 ( .A1(n6765), .A2(n6764), .ZN(n10038) );
  NOR2_X1 U8351 ( .A1(n10039), .A2(n10038), .ZN(n6766) );
  NOR2_X1 U8352 ( .A1(n6767), .A2(n6766), .ZN(n6768) );
  NOR2_X1 U8353 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6768), .ZN(n10022) );
  AND2_X1 U8354 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6768), .ZN(n10021) );
  NOR2_X1 U8355 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10021), .ZN(n6769) );
  NOR2_X1 U8356 ( .A1(n10022), .A2(n6769), .ZN(n6770) );
  NAND2_X1 U8357 ( .A1(n6770), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6772) );
  XOR2_X1 U8358 ( .A(n6770), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10020) );
  NAND2_X1 U8359 ( .A1(n10020), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U8360 ( .A1(n6772), .A2(n6771), .ZN(n6773) );
  NAND2_X1 U8361 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n6773), .ZN(n6775) );
  XOR2_X1 U8362 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n6773), .Z(n10033) );
  NAND2_X1 U8363 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10033), .ZN(n6774) );
  NAND2_X1 U8364 ( .A1(n6775), .A2(n6774), .ZN(n6776) );
  AND2_X1 U8365 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n6776), .ZN(n6777) );
  XNOR2_X1 U8366 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n6776), .ZN(n10032) );
  NOR2_X1 U8367 ( .A1(n5253), .A2(n10032), .ZN(n10031) );
  NOR2_X1 U8368 ( .A1(n6777), .A2(n10031), .ZN(n6778) );
  NOR2_X1 U8369 ( .A1(n6778), .A2(n5225), .ZN(n6779) );
  INV_X1 U8370 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10030) );
  XNOR2_X1 U8371 ( .A(n5225), .B(n6778), .ZN(n10029) );
  NOR2_X1 U8372 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  NOR2_X1 U8373 ( .A1(n6779), .A2(n10028), .ZN(n9862) );
  NAND2_X1 U8374 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n6780) );
  OAI21_X1 U8375 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n6780), .ZN(n9861) );
  NOR2_X1 U8376 ( .A1(n9862), .A2(n9861), .ZN(n9860) );
  AOI21_X1 U8377 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9860), .ZN(n9859) );
  NAND2_X1 U8378 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n6781) );
  OAI21_X1 U8379 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6781), .ZN(n9858) );
  NOR2_X1 U8380 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  AOI21_X1 U8381 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9857), .ZN(n9856) );
  NOR2_X1 U8382 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6782) );
  AOI21_X1 U8383 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6782), .ZN(n9855) );
  NAND2_X1 U8384 ( .A1(n9856), .A2(n9855), .ZN(n9854) );
  OAI21_X1 U8385 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9854), .ZN(n9852) );
  NAND2_X1 U8386 ( .A1(n9853), .A2(n9852), .ZN(n9851) );
  OAI21_X1 U8387 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9851), .ZN(n9849) );
  NAND2_X1 U8388 ( .A1(n9850), .A2(n9849), .ZN(n9848) );
  OAI21_X1 U8389 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9848), .ZN(n9846) );
  NAND2_X1 U8390 ( .A1(n9847), .A2(n9846), .ZN(n9845) );
  OAI21_X1 U8391 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9845), .ZN(n9843) );
  NAND2_X1 U8392 ( .A1(n9844), .A2(n9843), .ZN(n9842) );
  OAI21_X1 U8393 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9842), .ZN(n9840) );
  NAND2_X1 U8394 ( .A1(n9841), .A2(n9840), .ZN(n9839) );
  OAI21_X1 U8395 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9839), .ZN(n10025) );
  NOR2_X1 U8396 ( .A1(n10026), .A2(n10025), .ZN(n6783) );
  NAND2_X1 U8397 ( .A1(n10026), .A2(n10025), .ZN(n10024) );
  OAI21_X1 U8398 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n6783), .A(n10024), .ZN(
        n6786) );
  XNOR2_X1 U8399 ( .A(n6784), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n6785) );
  XNOR2_X1 U8400 ( .A(n6786), .B(n6785), .ZN(ADD_1071_U4) );
  XNOR2_X1 U8401 ( .A(n6950), .B(n7439), .ZN(n6787) );
  OR2_X1 U8402 ( .A1(n6325), .A2(n6844), .ZN(n6788) );
  NAND2_X1 U8403 ( .A1(n6787), .A2(n6788), .ZN(n6831) );
  INV_X1 U8404 ( .A(n6787), .ZN(n6790) );
  INV_X1 U8405 ( .A(n6788), .ZN(n6789) );
  NAND2_X1 U8406 ( .A1(n6790), .A2(n6789), .ZN(n6791) );
  NAND2_X1 U8407 ( .A1(n6831), .A2(n6791), .ZN(n6802) );
  INV_X1 U8408 ( .A(n6794), .ZN(n6796) );
  NAND2_X1 U8409 ( .A1(n6796), .A2(n6795), .ZN(n6797) );
  INV_X1 U8410 ( .A(n6798), .ZN(n6800) );
  INV_X1 U8411 ( .A(n6802), .ZN(n6799) );
  NAND2_X1 U8412 ( .A1(n6800), .A2(n6799), .ZN(n6832) );
  INV_X1 U8413 ( .A(n6832), .ZN(n6801) );
  AOI21_X1 U8414 ( .B1(n6802), .B2(n6798), .A(n6801), .ZN(n6810) );
  INV_X1 U8415 ( .A(n6803), .ZN(n6807) );
  INV_X1 U8416 ( .A(n8142), .ZN(n9729) );
  NAND2_X1 U8417 ( .A1(n9729), .A2(n6804), .ZN(n6806) );
  OAI211_X1 U8418 ( .C1(n9737), .C2(n6807), .A(n6806), .B(n6805), .ZN(n6808)
         );
  AOI21_X1 U8419 ( .B1(n6950), .B2(n8147), .A(n6808), .ZN(n6809) );
  OAI21_X1 U8420 ( .B1(n6810), .B2(n8128), .A(n6809), .ZN(P2_U3226) );
  NAND2_X1 U8421 ( .A1(n6824), .A2(n7995), .ZN(n6812) );
  NAND2_X1 U8422 ( .A1(n4265), .A2(n8946), .ZN(n6811) );
  NAND2_X1 U8423 ( .A1(n6812), .A2(n6811), .ZN(n6813) );
  XNOR2_X1 U8424 ( .A(n6813), .B(n8009), .ZN(n6861) );
  NOR2_X1 U8425 ( .A1(n8012), .A2(n6814), .ZN(n6815) );
  AOI21_X1 U8426 ( .B1(n6824), .B2(n4265), .A(n6815), .ZN(n6862) );
  XNOR2_X1 U8427 ( .A(n6861), .B(n6862), .ZN(n6822) );
  INV_X1 U8428 ( .A(n6816), .ZN(n6818) );
  INV_X1 U8429 ( .A(n6974), .ZN(n6820) );
  AOI211_X1 U8430 ( .C1(n6822), .C2(n6821), .A(n8650), .B(n6820), .ZN(n6830)
         );
  AOI21_X1 U8431 ( .B1(n8633), .B2(n9358), .A(n6823), .ZN(n6828) );
  NAND2_X1 U8432 ( .A1(n6824), .A2(n8648), .ZN(n6827) );
  NAND2_X1 U8433 ( .A1(n8660), .A2(n9364), .ZN(n6826) );
  INV_X1 U8434 ( .A(n6982), .ZN(n9356) );
  NAND2_X1 U8435 ( .A1(n8644), .A2(n9356), .ZN(n6825) );
  NAND4_X1 U8436 ( .A1(n6828), .A2(n6827), .A3(n6826), .A4(n6825), .ZN(n6829)
         );
  OR2_X1 U8437 ( .A1(n6830), .A2(n6829), .ZN(P1_U3234) );
  NAND2_X1 U8438 ( .A1(n6878), .A2(n5954), .ZN(n6835) );
  AOI22_X1 U8439 ( .A1(n7339), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7338), .B2(
        n6833), .ZN(n6834) );
  XNOR2_X1 U8440 ( .A(n8513), .B(n8043), .ZN(n7040) );
  NOR2_X1 U8441 ( .A1(n6325), .A2(n7046), .ZN(n7041) );
  XNOR2_X1 U8442 ( .A(n7040), .B(n7041), .ZN(n7042) );
  XNOR2_X1 U8443 ( .A(n7043), .B(n7042), .ZN(n6852) );
  INV_X1 U8444 ( .A(n6961), .ZN(n6849) );
  NAND2_X1 U8445 ( .A1(n7320), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U8446 ( .A1(n5595), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6842) );
  INV_X1 U8447 ( .A(n6838), .ZN(n6836) );
  NAND2_X1 U8448 ( .A1(n6836), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7024) );
  INV_X1 U8449 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U8450 ( .A1(n6838), .A2(n6837), .ZN(n6839) );
  AND2_X1 U8451 ( .A1(n7024), .A2(n6839), .ZN(n7049) );
  NAND2_X1 U8452 ( .A1(n7518), .A2(n7049), .ZN(n6841) );
  NAND2_X1 U8453 ( .A1(n5609), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6840) );
  OR2_X1 U8454 ( .A1(n7077), .A2(n8330), .ZN(n6846) );
  OR2_X1 U8455 ( .A1(n6844), .A2(n8328), .ZN(n6845) );
  NAND2_X1 U8456 ( .A1(n6846), .A2(n6845), .ZN(n6955) );
  NAND2_X1 U8457 ( .A1(n9729), .A2(n6955), .ZN(n6848) );
  OAI211_X1 U8458 ( .C1(n9737), .C2(n6849), .A(n6848), .B(n6847), .ZN(n6850)
         );
  AOI21_X1 U8459 ( .B1(n8513), .B2(n8147), .A(n6850), .ZN(n6851) );
  OAI21_X1 U8460 ( .B1(n6852), .B2(n8128), .A(n6851), .ZN(P2_U3236) );
  NAND2_X1 U8461 ( .A1(n6876), .A2(n7995), .ZN(n6854) );
  OR2_X1 U8462 ( .A1(n6982), .A2(n6180), .ZN(n6853) );
  NAND2_X1 U8463 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  XNOR2_X1 U8464 ( .A(n6855), .B(n8009), .ZN(n6860) );
  INV_X1 U8465 ( .A(n6860), .ZN(n6858) );
  NOR2_X1 U8466 ( .A1(n8012), .A2(n6982), .ZN(n6856) );
  AOI21_X1 U8467 ( .B1(n6876), .B2(n4265), .A(n6856), .ZN(n6859) );
  INV_X1 U8468 ( .A(n6859), .ZN(n6857) );
  NAND2_X1 U8469 ( .A1(n6858), .A2(n6857), .ZN(n6969) );
  NAND2_X1 U8470 ( .A1(n6860), .A2(n6859), .ZN(n6971) );
  NAND2_X1 U8471 ( .A1(n6969), .A2(n6971), .ZN(n6866) );
  INV_X1 U8472 ( .A(n6861), .ZN(n6864) );
  INV_X1 U8473 ( .A(n6862), .ZN(n6863) );
  NAND2_X1 U8474 ( .A1(n6864), .A2(n6863), .ZN(n6970) );
  NAND2_X1 U8475 ( .A1(n6974), .A2(n6970), .ZN(n6865) );
  XOR2_X1 U8476 ( .A(n6866), .B(n6865), .Z(n6875) );
  NAND2_X1 U8477 ( .A1(n8633), .A2(n8946), .ZN(n6872) );
  NAND2_X1 U8478 ( .A1(n8644), .A2(n8945), .ZN(n6871) );
  NAND2_X1 U8479 ( .A1(n8660), .A2(n6867), .ZN(n6870) );
  NOR2_X1 U8480 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6868), .ZN(n9492) );
  INV_X1 U8481 ( .A(n9492), .ZN(n6869) );
  NAND4_X1 U8482 ( .A1(n6872), .A2(n6871), .A3(n6870), .A4(n6869), .ZN(n6873)
         );
  AOI21_X1 U8483 ( .B1(n6876), .B2(n8648), .A(n6873), .ZN(n6874) );
  OAI21_X1 U8484 ( .B1(n6875), .B2(n8650), .A(n6874), .ZN(P1_U3222) );
  NAND2_X1 U8485 ( .A1(n6878), .A2(n6363), .ZN(n6880) );
  AOI22_X1 U8486 ( .A1(n7823), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7822), .B2(
        n9506), .ZN(n6879) );
  OR2_X1 U8487 ( .A1(n6984), .A2(n7144), .ZN(n8804) );
  NAND2_X1 U8488 ( .A1(n6984), .A2(n7144), .ZN(n8828) );
  XNOR2_X1 U8489 ( .A(n6942), .B(n8909), .ZN(n9398) );
  OAI21_X1 U8490 ( .B1(n8909), .B2(n6882), .A(n6926), .ZN(n6883) );
  NAND2_X1 U8491 ( .A1(n6883), .A2(n9612), .ZN(n6892) );
  NAND2_X1 U8492 ( .A1(n7826), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U8493 ( .A1(n7983), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6889) );
  INV_X1 U8494 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7142) );
  NAND2_X1 U8495 ( .A1(n6885), .A2(n7142), .ZN(n6886) );
  AND2_X1 U8496 ( .A1(n6931), .A2(n6886), .ZN(n7146) );
  NAND2_X1 U8497 ( .A1(n5712), .A2(n7146), .ZN(n6888) );
  NAND2_X1 U8498 ( .A1(n8735), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6887) );
  INV_X1 U8499 ( .A(n7129), .ZN(n8944) );
  AOI22_X1 U8500 ( .A1(n9359), .A2(n9356), .B1(n9357), .B2(n8944), .ZN(n6891)
         );
  NAND2_X1 U8501 ( .A1(n6892), .A2(n6891), .ZN(n6893) );
  AOI21_X1 U8502 ( .B1(n9398), .B2(n9363), .A(n6893), .ZN(n9400) );
  NAND2_X1 U8503 ( .A1(n6895), .A2(n6984), .ZN(n6894) );
  NAND2_X1 U8504 ( .A1(n6894), .A2(n9633), .ZN(n6896) );
  NOR2_X2 U8505 ( .A1(n6895), .A2(n6984), .ZN(n6944) );
  OR2_X1 U8506 ( .A1(n6896), .A2(n6944), .ZN(n9395) );
  AOI22_X1 U8507 ( .A1(n9598), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n6979), .B2(
        n9586), .ZN(n6898) );
  NAND2_X1 U8508 ( .A1(n6984), .A2(n9132), .ZN(n6897) );
  OAI211_X1 U8509 ( .C1(n9395), .C2(n6899), .A(n6898), .B(n6897), .ZN(n6900)
         );
  AOI21_X1 U8510 ( .B1(n9398), .B2(n9604), .A(n6900), .ZN(n6901) );
  OAI21_X1 U8511 ( .B1(n9400), .B2(n9598), .A(n6901), .ZN(P1_U3278) );
  INV_X1 U8512 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6907) );
  AOI22_X1 U8513 ( .A1(n6902), .A2(n9810), .B1(n9809), .B2(n6950), .ZN(n6903)
         );
  OAI211_X1 U8514 ( .C1(n6905), .C2(n9804), .A(n6904), .B(n6903), .ZN(n6908)
         );
  NAND2_X1 U8515 ( .A1(n6908), .A2(n4267), .ZN(n6906) );
  OAI21_X1 U8516 ( .B1(n4267), .B2(n6907), .A(n6906), .ZN(P2_U3487) );
  NAND2_X1 U8517 ( .A1(n6908), .A2(n4268), .ZN(n6909) );
  OAI21_X1 U8518 ( .B1(n4268), .B2(n6910), .A(n6909), .ZN(P2_U3532) );
  INV_X1 U8519 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6918) );
  OAI22_X1 U8520 ( .A1(n6912), .A2(n9781), .B1(n4540), .B2(n9820), .ZN(n6913)
         );
  INV_X1 U8521 ( .A(n6913), .ZN(n6914) );
  OAI211_X1 U8522 ( .C1(n9814), .C2(n6916), .A(n6915), .B(n6914), .ZN(n6919)
         );
  NAND2_X1 U8523 ( .A1(n6919), .A2(n4267), .ZN(n6917) );
  OAI21_X1 U8524 ( .B1(n4267), .B2(n6918), .A(n6917), .ZN(P2_U3481) );
  NAND2_X1 U8525 ( .A1(n6919), .A2(n4268), .ZN(n6920) );
  OAI21_X1 U8526 ( .B1(n4268), .B2(n6921), .A(n6920), .ZN(P2_U3530) );
  INV_X1 U8527 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7397) );
  INV_X1 U8528 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9920) );
  MUX2_X1 U8529 ( .A(n7397), .B(n9920), .S(n7537), .Z(n7054) );
  XNOR2_X1 U8530 ( .A(n7054), .B(SI_24_), .ZN(n7053) );
  XNOR2_X1 U8531 ( .A(n7058), .B(n7053), .ZN(n7924) );
  INV_X1 U8532 ( .A(n7924), .ZN(n6987) );
  OAI222_X1 U8533 ( .A1(P2_U3152), .A2(n6925), .B1(n4270), .B2(n6987), .C1(
        n7397), .C2(n8545), .ZN(P2_U3334) );
  NAND2_X1 U8534 ( .A1(n6926), .A2(n8828), .ZN(n7107) );
  NAND2_X1 U8535 ( .A1(n7009), .A2(n6363), .ZN(n6928) );
  INV_X1 U8536 ( .A(n8973), .ZN(n9519) );
  AOI22_X1 U8537 ( .A1(n7823), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7822), .B2(
        n9519), .ZN(n6927) );
  XNOR2_X1 U8538 ( .A(n7106), .B(n7129), .ZN(n8912) );
  INV_X1 U8539 ( .A(n8912), .ZN(n6929) );
  XNOR2_X1 U8540 ( .A(n7107), .B(n6929), .ZN(n6939) );
  NAND2_X1 U8541 ( .A1(n7983), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6936) );
  NAND2_X1 U8542 ( .A1(n8735), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6935) );
  INV_X1 U8543 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U8544 ( .A1(n6931), .A2(n6930), .ZN(n6932) );
  AND2_X1 U8545 ( .A1(n7100), .A2(n6932), .ZN(n7170) );
  NAND2_X1 U8546 ( .A1(n5712), .A2(n7170), .ZN(n6934) );
  NAND2_X1 U8547 ( .A1(n7826), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6933) );
  INV_X1 U8548 ( .A(n7257), .ZN(n8943) );
  NAND2_X1 U8549 ( .A1(n9357), .A2(n8943), .ZN(n6937) );
  OAI21_X1 U8550 ( .B1(n7144), .B2(n9608), .A(n6937), .ZN(n6938) );
  AOI21_X1 U8551 ( .B1(n6939), .B2(n9612), .A(n6938), .ZN(n9390) );
  NAND2_X1 U8552 ( .A1(n9396), .A2(n7144), .ZN(n6941) );
  XNOR2_X1 U8553 ( .A(n4274), .B(n8912), .ZN(n9393) );
  NAND2_X1 U8554 ( .A1(n9393), .A2(n9171), .ZN(n6949) );
  AND2_X2 U8555 ( .A1(n6944), .A2(n9391), .ZN(n7109) );
  INV_X1 U8556 ( .A(n7109), .ZN(n6943) );
  OAI211_X1 U8557 ( .C1(n9391), .C2(n6944), .A(n6943), .B(n9633), .ZN(n9389)
         );
  INV_X1 U8558 ( .A(n9389), .ZN(n6947) );
  AOI22_X1 U8559 ( .A1(n9598), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7146), .B2(
        n9586), .ZN(n6945) );
  OAI21_X1 U8560 ( .B1(n9391), .B2(n9619), .A(n6945), .ZN(n6946) );
  AOI21_X1 U8561 ( .B1(n6947), .B2(n9209), .A(n6946), .ZN(n6948) );
  OAI211_X1 U8562 ( .C1(n9598), .C2(n9390), .A(n6949), .B(n6948), .ZN(P1_U3277) );
  OR2_X1 U8563 ( .A1(n8513), .A2(n7046), .ZN(n7621) );
  NAND2_X1 U8564 ( .A1(n8513), .A2(n7046), .ZN(n7620) );
  NAND2_X1 U8565 ( .A1(n7621), .A2(n7620), .ZN(n7018) );
  NAND2_X1 U8566 ( .A1(n6952), .A2(n7730), .ZN(n6953) );
  NAND2_X1 U8567 ( .A1(n7008), .A2(n6953), .ZN(n8516) );
  XNOR2_X1 U8568 ( .A(n7019), .B(n7018), .ZN(n6956) );
  AOI21_X1 U8569 ( .B1(n6956), .B2(n8414), .A(n6955), .ZN(n6957) );
  OAI21_X1 U8570 ( .B1(n8516), .B2(n7181), .A(n6957), .ZN(n8518) );
  NAND2_X1 U8571 ( .A1(n8518), .A2(n6958), .ZN(n6967) );
  INV_X1 U8572 ( .A(n7014), .ZN(n7016) );
  NAND2_X1 U8573 ( .A1(n6959), .A2(n8513), .ZN(n6960) );
  AND2_X1 U8574 ( .A1(n7016), .A2(n6960), .ZN(n8514) );
  INV_X1 U8575 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U8576 ( .A1(n8513), .A2(n8406), .ZN(n6963) );
  NAND2_X1 U8577 ( .A1(n8408), .A2(n6961), .ZN(n6962) );
  OAI211_X1 U8578 ( .C1(n8422), .C2(n6964), .A(n6963), .B(n6962), .ZN(n6965)
         );
  AOI21_X1 U8579 ( .B1(n8514), .B2(n8409), .A(n6965), .ZN(n6966) );
  OAI211_X1 U8580 ( .C1(n8516), .C2(n6968), .A(n6967), .B(n6966), .ZN(P2_U3283) );
  AND2_X1 U8581 ( .A1(n6970), .A2(n6969), .ZN(n6973) );
  INV_X1 U8582 ( .A(n6971), .ZN(n6972) );
  OR2_X1 U8583 ( .A1(n9396), .A2(n6180), .ZN(n6976) );
  NAND2_X1 U8584 ( .A1(n7974), .A2(n8945), .ZN(n6975) );
  NAND2_X1 U8585 ( .A1(n6976), .A2(n6975), .ZN(n7125) );
  OAI22_X1 U8586 ( .A1(n9396), .A2(n7900), .B1(n7144), .B2(n6180), .ZN(n6977)
         );
  XNOR2_X1 U8587 ( .A(n6977), .B(n7989), .ZN(n7126) );
  XOR2_X1 U8588 ( .A(n7125), .B(n7126), .Z(n6978) );
  XNOR2_X1 U8589 ( .A(n7127), .B(n6978), .ZN(n6986) );
  AND2_X1 U8590 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9505) );
  AOI21_X1 U8591 ( .B1(n8644), .B2(n8944), .A(n9505), .ZN(n6981) );
  NAND2_X1 U8592 ( .A1(n8660), .A2(n6979), .ZN(n6980) );
  OAI211_X1 U8593 ( .C1(n6982), .C2(n8656), .A(n6981), .B(n6980), .ZN(n6983)
         );
  AOI21_X1 U8594 ( .B1(n6984), .B2(n8648), .A(n6983), .ZN(n6985) );
  OAI21_X1 U8595 ( .B1(n6986), .B2(n8650), .A(n6985), .ZN(P1_U3232) );
  OAI222_X1 U8596 ( .A1(n9328), .A2(n9920), .B1(P1_U3084), .B2(n6988), .C1(
        n8059), .C2(n6987), .ZN(P1_U3329) );
  AOI21_X1 U8597 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n7215), .A(n6989), .ZN(
        n8162) );
  XNOR2_X1 U8598 ( .A(n8162), .B(n7312), .ZN(n6991) );
  INV_X1 U8599 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U8600 ( .A1(n6991), .A2(n6990), .ZN(n8164) );
  OAI21_X1 U8601 ( .B1(n6991), .B2(n6990), .A(n8164), .ZN(n6992) );
  NAND2_X1 U8602 ( .A1(n6992), .A2(n9749), .ZN(n7006) );
  AND2_X1 U8603 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7325) );
  INV_X1 U8604 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6993) );
  NAND2_X1 U8605 ( .A1(n8161), .A2(n6993), .ZN(n8166) );
  NAND2_X1 U8606 ( .A1(n7312), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6994) );
  NAND2_X1 U8607 ( .A1(n8166), .A2(n6994), .ZN(n7002) );
  INV_X1 U8608 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7000) );
  INV_X1 U8609 ( .A(n6995), .ZN(n6996) );
  NAND2_X1 U8610 ( .A1(n6997), .A2(n6996), .ZN(n6998) );
  OAI21_X1 U8611 ( .B1(n7000), .B2(n6999), .A(n6998), .ZN(n7001) );
  OR2_X1 U8612 ( .A1(n7002), .A2(n7001), .ZN(n8167) );
  NAND2_X1 U8613 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  AOI21_X1 U8614 ( .B1(n8167), .B2(n7003), .A(n9740), .ZN(n7004) );
  AOI211_X1 U8615 ( .C1(n9747), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n7325), .B(
        n7004), .ZN(n7005) );
  OAI211_X1 U8616 ( .C1(n9739), .C2(n8161), .A(n7006), .B(n7005), .ZN(P2_U3263) );
  INV_X1 U8617 ( .A(n7046), .ZN(n8151) );
  NAND2_X1 U8618 ( .A1(n8513), .A2(n8151), .ZN(n7007) );
  NAND2_X1 U8619 ( .A1(n7008), .A2(n7007), .ZN(n7066) );
  NAND2_X1 U8620 ( .A1(n7009), .A2(n5954), .ZN(n7012) );
  AOI22_X1 U8621 ( .A1(n7339), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7338), .B2(
        n7010), .ZN(n7011) );
  NAND2_X1 U8622 ( .A1(n8508), .A2(n7077), .ZN(n7628) );
  NAND2_X1 U8623 ( .A1(n7629), .A2(n7628), .ZN(n7625) );
  XNOR2_X1 U8624 ( .A(n7066), .B(n7625), .ZN(n8512) );
  INV_X1 U8625 ( .A(n7072), .ZN(n7015) );
  AOI21_X1 U8626 ( .B1(n8508), .B2(n7016), .A(n7015), .ZN(n8509) );
  AOI22_X1 U8627 ( .A1(n8402), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7049), .B2(
        n8408), .ZN(n7017) );
  OAI21_X1 U8628 ( .B1(n7013), .B2(n8368), .A(n7017), .ZN(n7033) );
  AOI21_X1 U8629 ( .B1(n7020), .B2(n7625), .A(n8326), .ZN(n7031) );
  NAND2_X1 U8630 ( .A1(n5609), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7029) );
  NAND2_X1 U8631 ( .A1(n7320), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7028) );
  INV_X1 U8632 ( .A(n7024), .ZN(n7022) );
  NAND2_X1 U8633 ( .A1(n7022), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7079) );
  INV_X1 U8634 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7023) );
  NAND2_X1 U8635 ( .A1(n7024), .A2(n7023), .ZN(n7025) );
  AND2_X1 U8636 ( .A1(n7079), .A2(n7025), .ZN(n7236) );
  NAND2_X1 U8637 ( .A1(n7518), .A2(n7236), .ZN(n7027) );
  NAND2_X1 U8638 ( .A1(n5595), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7026) );
  OAI22_X1 U8639 ( .A1(n7046), .A2(n8328), .B1(n8106), .B2(n8330), .ZN(n7030)
         );
  AOI21_X1 U8640 ( .B1(n7031), .B2(n7075), .A(n7030), .ZN(n8511) );
  NOR2_X1 U8641 ( .A1(n8511), .A2(n8402), .ZN(n7032) );
  AOI211_X1 U8642 ( .C1(n8509), .C2(n8409), .A(n7033), .B(n7032), .ZN(n7034)
         );
  OAI21_X1 U8643 ( .B1(n8399), .B2(n8512), .A(n7034), .ZN(P2_U3282) );
  XNOR2_X1 U8644 ( .A(n8508), .B(n7439), .ZN(n7035) );
  OR2_X1 U8645 ( .A1(n6325), .A2(n7077), .ZN(n7036) );
  NAND2_X1 U8646 ( .A1(n7035), .A2(n7036), .ZN(n7204) );
  INV_X1 U8647 ( .A(n7035), .ZN(n7038) );
  INV_X1 U8648 ( .A(n7036), .ZN(n7037) );
  NAND2_X1 U8649 ( .A1(n7038), .A2(n7037), .ZN(n7039) );
  NAND2_X1 U8650 ( .A1(n7204), .A2(n7039), .ZN(n7045) );
  AOI21_X1 U8651 ( .B1(n7045), .B2(n7044), .A(n4342), .ZN(n7052) );
  OAI22_X1 U8652 ( .A1(n8135), .A2(n7046), .B1(n8106), .B2(n9714), .ZN(n7047)
         );
  AOI211_X1 U8653 ( .C1(n8140), .C2(n7049), .A(n7048), .B(n7047), .ZN(n7051)
         );
  NAND2_X1 U8654 ( .A1(n8508), .A2(n8147), .ZN(n7050) );
  OAI211_X1 U8655 ( .C1(n7052), .C2(n8128), .A(n7051), .B(n7050), .ZN(P2_U3217) );
  INV_X1 U8656 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7423) );
  INV_X1 U8657 ( .A(n7053), .ZN(n7057) );
  INV_X1 U8658 ( .A(n7054), .ZN(n7055) );
  NAND2_X1 U8659 ( .A1(n7055), .A2(SI_24_), .ZN(n7056) );
  INV_X1 U8660 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9970) );
  MUX2_X1 U8661 ( .A(n7423), .B(n9970), .S(n7537), .Z(n7060) );
  INV_X1 U8662 ( .A(SI_25_), .ZN(n7059) );
  NAND2_X1 U8663 ( .A1(n7060), .A2(n7059), .ZN(n7115) );
  INV_X1 U8664 ( .A(n7060), .ZN(n7061) );
  NAND2_X1 U8665 ( .A1(n7061), .A2(SI_25_), .ZN(n7062) );
  NAND2_X1 U8666 ( .A1(n7115), .A2(n7062), .ZN(n7116) );
  INV_X1 U8667 ( .A(n7940), .ZN(n7065) );
  OAI222_X1 U8668 ( .A1(n8545), .A2(n7423), .B1(n4270), .B2(n7065), .C1(
        P2_U3152), .C2(n7063), .ZN(P2_U3333) );
  OAI222_X1 U8669 ( .A1(n9328), .A2(n9970), .B1(n8059), .B2(n7065), .C1(n7064), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U8670 ( .A(n7077), .ZN(n8150) );
  OAI22_X2 U8671 ( .A1(n7066), .A2(n7021), .B1(n8508), .B2(n8150), .ZN(n7070)
         );
  NAND2_X1 U8672 ( .A1(n7095), .A2(n5954), .ZN(n7069) );
  AOI22_X1 U8673 ( .A1(n7339), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7338), .B2(
        n7067), .ZN(n7068) );
  NAND2_X1 U8674 ( .A1(n8503), .A2(n8106), .ZN(n7552) );
  OAI21_X1 U8675 ( .B1(n7070), .B2(n7732), .A(n7175), .ZN(n7071) );
  INV_X1 U8676 ( .A(n7071), .ZN(n8507) );
  AOI21_X1 U8677 ( .B1(n8503), .B2(n7072), .A(n4351), .ZN(n8504) );
  INV_X1 U8678 ( .A(n8503), .ZN(n7074) );
  AOI22_X1 U8679 ( .A1(n8402), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7236), .B2(
        n8408), .ZN(n7073) );
  OAI21_X1 U8680 ( .B1(n7074), .B2(n8368), .A(n7073), .ZN(n7089) );
  NAND2_X1 U8681 ( .A1(n7075), .A2(n7629), .ZN(n7076) );
  NAND2_X1 U8682 ( .A1(n7076), .A2(n7632), .ZN(n7182) );
  OAI211_X1 U8683 ( .C1(n7076), .C2(n7632), .A(n7182), .B(n8384), .ZN(n7087)
         );
  OR2_X1 U8684 ( .A1(n7077), .A2(n8328), .ZN(n7086) );
  NAND2_X1 U8685 ( .A1(n7525), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7084) );
  NAND2_X1 U8686 ( .A1(n5609), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U8687 ( .A1(n7079), .A2(n7078), .ZN(n7080) );
  AND2_X1 U8688 ( .A1(n7187), .A2(n7080), .ZN(n8109) );
  NAND2_X1 U8689 ( .A1(n7518), .A2(n8109), .ZN(n7082) );
  NAND2_X1 U8690 ( .A1(n5595), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7081) );
  AND4_X1 U8691 ( .A1(n7084), .A2(n7083), .A3(n7082), .A4(n7081), .ZN(n7762)
         );
  OR2_X1 U8692 ( .A1(n7762), .A2(n8330), .ZN(n7085) );
  AND2_X1 U8693 ( .A1(n7086), .A2(n7085), .ZN(n7233) );
  AND2_X1 U8694 ( .A1(n7087), .A2(n7233), .ZN(n8506) );
  NOR2_X1 U8695 ( .A1(n8506), .A2(n8402), .ZN(n7088) );
  AOI211_X1 U8696 ( .C1(n8504), .C2(n8409), .A(n7089), .B(n7088), .ZN(n7090)
         );
  OAI21_X1 U8697 ( .B1(n8507), .B2(n8399), .A(n7090), .ZN(P2_U3281) );
  INV_X1 U8698 ( .A(n7091), .ZN(n7094) );
  OAI21_X2 U8699 ( .B1(n7094), .B2(n7093), .A(n7092), .ZN(n7260) );
  NAND2_X1 U8700 ( .A1(n7095), .A2(n6363), .ZN(n7097) );
  AOI22_X1 U8701 ( .A1(n7823), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7822), .B2(
        n9532), .ZN(n7096) );
  OR2_X1 U8702 ( .A1(n7261), .A2(n7257), .ZN(n7286) );
  NAND2_X1 U8703 ( .A1(n7261), .A2(n7257), .ZN(n8709) );
  NAND2_X1 U8704 ( .A1(n7286), .A2(n8709), .ZN(n8830) );
  XNOR2_X1 U8705 ( .A(n7260), .B(n8830), .ZN(n9387) );
  INV_X1 U8706 ( .A(n9387), .ZN(n7114) );
  NAND2_X1 U8707 ( .A1(n7983), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7105) );
  INV_X1 U8708 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7099) );
  NAND2_X1 U8709 ( .A1(n7100), .A2(n7099), .ZN(n7101) );
  AND2_X1 U8710 ( .A1(n7246), .A2(n7101), .ZN(n7301) );
  NAND2_X1 U8711 ( .A1(n5712), .A2(n7301), .ZN(n7104) );
  NAND2_X1 U8712 ( .A1(n8735), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7103) );
  NAND2_X1 U8713 ( .A1(n7826), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7102) );
  OR2_X1 U8714 ( .A1(n7106), .A2(n7129), .ZN(n8805) );
  INV_X1 U8715 ( .A(n8830), .ZN(n8910) );
  XNOR2_X1 U8716 ( .A(n7285), .B(n8910), .ZN(n7108) );
  OAI222_X1 U8717 ( .A1(n9610), .A2(n7294), .B1(n9608), .B2(n7129), .C1(n9591), 
        .C2(n7108), .ZN(n9385) );
  NAND2_X1 U8718 ( .A1(n7109), .A2(n9383), .ZN(n7255) );
  OAI21_X1 U8719 ( .B1(n7109), .B2(n9383), .A(n7255), .ZN(n9384) );
  AOI22_X1 U8720 ( .A1(n9598), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7170), .B2(
        n9586), .ZN(n7111) );
  NAND2_X1 U8721 ( .A1(n7261), .A2(n9132), .ZN(n7110) );
  OAI211_X1 U8722 ( .C1(n9384), .C2(n9000), .A(n7111), .B(n7110), .ZN(n7112)
         );
  AOI21_X1 U8723 ( .B1(n9385), .B2(n9617), .A(n7112), .ZN(n7113) );
  OAI21_X1 U8724 ( .B1(n7114), .B2(n9228), .A(n7113), .ZN(P1_U3276) );
  INV_X1 U8725 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7436) );
  INV_X1 U8726 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7960) );
  MUX2_X1 U8727 ( .A(n7436), .B(n7960), .S(n4276), .Z(n7119) );
  INV_X1 U8728 ( .A(SI_26_), .ZN(n7118) );
  NAND2_X1 U8729 ( .A1(n7119), .A2(n7118), .ZN(n7151) );
  INV_X1 U8730 ( .A(n7119), .ZN(n7120) );
  NAND2_X1 U8731 ( .A1(n7120), .A2(SI_26_), .ZN(n7121) );
  AND2_X1 U8732 ( .A1(n7151), .A2(n7121), .ZN(n7149) );
  INV_X1 U8733 ( .A(n7959), .ZN(n7123) );
  OAI222_X1 U8734 ( .A1(P2_U3152), .A2(n7122), .B1(n4270), .B2(n7123), .C1(
        n7436), .C2(n8545), .ZN(P2_U3332) );
  OAI222_X1 U8735 ( .A1(n9328), .A2(n7960), .B1(P1_U3084), .B2(n7124), .C1(
        n8059), .C2(n7123), .ZN(P1_U3327) );
  NAND2_X1 U8736 ( .A1(n7127), .A2(n7126), .ZN(n7128) );
  OAI22_X1 U8737 ( .A1(n9391), .A2(n7900), .B1(n7129), .B2(n6180), .ZN(n7130)
         );
  XNOR2_X1 U8738 ( .A(n7130), .B(n7989), .ZN(n7132) );
  INV_X1 U8739 ( .A(n7161), .ZN(n7141) );
  INV_X1 U8740 ( .A(n7131), .ZN(n7134) );
  INV_X1 U8741 ( .A(n7132), .ZN(n7133) );
  NAND2_X1 U8742 ( .A1(n7134), .A2(n7133), .ZN(n7138) );
  OR2_X1 U8743 ( .A1(n9391), .A2(n6180), .ZN(n7136) );
  NAND2_X1 U8744 ( .A1(n7974), .A2(n8944), .ZN(n7135) );
  NAND2_X1 U8745 ( .A1(n7136), .A2(n7135), .ZN(n7137) );
  AOI21_X1 U8746 ( .B1(n7138), .B2(n7161), .A(n7137), .ZN(n7139) );
  NOR2_X1 U8747 ( .A1(n7139), .A2(n8650), .ZN(n7140) );
  OAI21_X1 U8748 ( .B1(n7141), .B2(n7163), .A(n7140), .ZN(n7148) );
  NOR2_X1 U8749 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7142), .ZN(n9518) );
  AOI21_X1 U8750 ( .B1(n8644), .B2(n8943), .A(n9518), .ZN(n7143) );
  OAI21_X1 U8751 ( .B1(n7144), .B2(n8656), .A(n7143), .ZN(n7145) );
  AOI21_X1 U8752 ( .B1(n7146), .B2(n8660), .A(n7145), .ZN(n7147) );
  OAI211_X1 U8753 ( .C1(n9391), .C2(n8663), .A(n7148), .B(n7147), .ZN(P1_U3213) );
  INV_X1 U8754 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7453) );
  NAND2_X1 U8755 ( .A1(n7150), .A2(n7149), .ZN(n7152) );
  INV_X1 U8756 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8056) );
  MUX2_X1 U8757 ( .A(n7453), .B(n8056), .S(n7537), .Z(n7154) );
  INV_X1 U8758 ( .A(SI_27_), .ZN(n7153) );
  NAND2_X1 U8759 ( .A1(n7154), .A2(n7153), .ZN(n7495) );
  INV_X1 U8760 ( .A(n7154), .ZN(n7155) );
  NAND2_X1 U8761 ( .A1(n7155), .A2(SI_27_), .ZN(n7156) );
  AND2_X1 U8762 ( .A1(n7495), .A2(n7156), .ZN(n7493) );
  INV_X1 U8763 ( .A(n7980), .ZN(n8054) );
  OAI222_X1 U8764 ( .A1(n8545), .A2(n7453), .B1(n4270), .B2(n8054), .C1(n7756), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  NAND2_X1 U8765 ( .A1(n7163), .A2(n7161), .ZN(n7159) );
  OAI22_X1 U8766 ( .A1(n9383), .A2(n7900), .B1(n7257), .B2(n6180), .ZN(n7157)
         );
  XNOR2_X1 U8767 ( .A(n7157), .B(n8009), .ZN(n7160) );
  INV_X1 U8768 ( .A(n7160), .ZN(n7158) );
  NAND2_X1 U8769 ( .A1(n7159), .A2(n7158), .ZN(n7290) );
  INV_X1 U8770 ( .A(n7290), .ZN(n7164) );
  OAI22_X1 U8771 ( .A1(n9383), .A2(n6180), .B1(n7257), .B2(n8012), .ZN(n7165)
         );
  OAI21_X1 U8772 ( .B1(n7164), .B2(n7291), .A(n8652), .ZN(n7173) );
  AOI21_X1 U8773 ( .B1(n7290), .B2(n7166), .A(n7165), .ZN(n7172) );
  NAND2_X1 U8774 ( .A1(n8633), .A2(n8944), .ZN(n7167) );
  NAND2_X1 U8775 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9526) );
  OAI211_X1 U8776 ( .C1(n7294), .C2(n8657), .A(n7167), .B(n9526), .ZN(n7169)
         );
  NOR2_X1 U8777 ( .A1(n9383), .A2(n8663), .ZN(n7168) );
  AOI211_X1 U8778 ( .C1(n7170), .C2(n8660), .A(n7169), .B(n7168), .ZN(n7171)
         );
  OAI21_X1 U8779 ( .B1(n7173), .B2(n7172), .A(n7171), .ZN(P1_U3239) );
  INV_X1 U8780 ( .A(n8106), .ZN(n8149) );
  OR2_X1 U8781 ( .A1(n8503), .A2(n8149), .ZN(n7174) );
  NAND2_X1 U8782 ( .A1(n7241), .A2(n5954), .ZN(n7178) );
  AOI22_X1 U8783 ( .A1(n7339), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7338), .B2(
        n7176), .ZN(n7177) );
  OR2_X1 U8784 ( .A1(n7763), .A2(n7762), .ZN(n7633) );
  NAND2_X1 U8785 ( .A1(n7763), .A2(n7762), .ZN(n7639) );
  NAND2_X1 U8786 ( .A1(n7633), .A2(n7639), .ZN(n7733) );
  NAND2_X1 U8787 ( .A1(n7179), .A2(n7183), .ZN(n7180) );
  NAND2_X1 U8788 ( .A1(n7765), .A2(n7180), .ZN(n7197) );
  OR2_X1 U8789 ( .A1(n7197), .A2(n7181), .ZN(n7196) );
  NAND2_X1 U8790 ( .A1(n7184), .A2(n7733), .ZN(n7185) );
  NAND2_X1 U8791 ( .A1(n7503), .A2(n7185), .ZN(n7194) );
  NAND2_X1 U8792 ( .A1(n7187), .A2(n7218), .ZN(n7188) );
  NAND2_X1 U8793 ( .A1(n7318), .A2(n7188), .ZN(n8390) );
  INV_X1 U8794 ( .A(n7518), .ZN(n7472) );
  OR2_X1 U8795 ( .A1(n8390), .A2(n7472), .ZN(n7192) );
  NAND2_X1 U8796 ( .A1(n7320), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U8797 ( .A1(n5609), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7190) );
  NAND2_X1 U8798 ( .A1(n5595), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7189) );
  OAI22_X1 U8799 ( .A1(n8105), .A2(n8330), .B1(n8106), .B2(n8328), .ZN(n7193)
         );
  AOI21_X1 U8800 ( .B1(n7194), .B2(n8384), .A(n7193), .ZN(n7195) );
  INV_X1 U8801 ( .A(n7197), .ZN(n8500) );
  INV_X1 U8802 ( .A(n7763), .ZN(n8497) );
  OR2_X1 U8803 ( .A1(n4351), .A2(n8497), .ZN(n7198) );
  NAND2_X1 U8804 ( .A1(n8393), .A2(n7198), .ZN(n8498) );
  AOI22_X1 U8805 ( .A1(n8402), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8109), .B2(
        n8408), .ZN(n7200) );
  NAND2_X1 U8806 ( .A1(n7763), .A2(n8406), .ZN(n7199) );
  OAI211_X1 U8807 ( .C1(n8498), .C2(n8295), .A(n7200), .B(n7199), .ZN(n7201)
         );
  AOI21_X1 U8808 ( .B1(n8500), .B2(n7202), .A(n7201), .ZN(n7203) );
  OAI21_X1 U8809 ( .B1(n8502), .B2(n8402), .A(n7203), .ZN(P2_U3280) );
  INV_X1 U8810 ( .A(n7228), .ZN(n7207) );
  XNOR2_X1 U8811 ( .A(n8503), .B(n7439), .ZN(n7229) );
  OR2_X1 U8812 ( .A1(n6325), .A2(n8106), .ZN(n7208) );
  AND2_X1 U8813 ( .A1(n7229), .A2(n7208), .ZN(n7205) );
  INV_X1 U8814 ( .A(n7205), .ZN(n7206) );
  XNOR2_X1 U8815 ( .A(n7763), .B(n7439), .ZN(n7214) );
  NOR2_X1 U8816 ( .A1(n6325), .A2(n7762), .ZN(n7212) );
  XNOR2_X1 U8817 ( .A(n7214), .B(n7212), .ZN(n8101) );
  INV_X1 U8818 ( .A(n7229), .ZN(n7209) );
  INV_X1 U8819 ( .A(n7208), .ZN(n7232) );
  NAND2_X1 U8820 ( .A1(n7209), .A2(n7232), .ZN(n7210) );
  AND2_X1 U8821 ( .A1(n8101), .A2(n7210), .ZN(n7211) );
  INV_X1 U8822 ( .A(n7212), .ZN(n7213) );
  NAND2_X1 U8823 ( .A1(n7269), .A2(n5954), .ZN(n7217) );
  AOI22_X1 U8824 ( .A1(n7339), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7338), .B2(
        n7215), .ZN(n7216) );
  XNOR2_X1 U8825 ( .A(n8493), .B(n8043), .ZN(n7306) );
  NOR2_X1 U8826 ( .A1(n6325), .A2(n8105), .ZN(n7307) );
  XNOR2_X1 U8827 ( .A(n7306), .B(n7307), .ZN(n7310) );
  XNOR2_X1 U8828 ( .A(n7311), .B(n7310), .ZN(n7227) );
  OAI22_X1 U8829 ( .A1(n9737), .A2(n8390), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7218), .ZN(n7225) );
  INV_X1 U8830 ( .A(n5595), .ZN(n7529) );
  NAND2_X1 U8831 ( .A1(n5609), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7220) );
  NAND2_X1 U8832 ( .A1(n7320), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7219) );
  OAI211_X1 U8833 ( .C1(n6990), .C2(n7529), .A(n7220), .B(n7219), .ZN(n7221)
         );
  INV_X1 U8834 ( .A(n7221), .ZN(n7223) );
  XNOR2_X1 U8835 ( .A(n7318), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U8836 ( .A1(n8366), .A2(n7518), .ZN(n7222) );
  AND2_X1 U8837 ( .A1(n7223), .A2(n7222), .ZN(n8074) );
  OAI22_X1 U8838 ( .A1(n8135), .A2(n7762), .B1(n8074), .B2(n9714), .ZN(n7224)
         );
  AOI211_X1 U8839 ( .C1(n8493), .C2(n8147), .A(n7225), .B(n7224), .ZN(n7226)
         );
  OAI21_X1 U8840 ( .B1(n7227), .B2(n8128), .A(n7226), .ZN(P2_U3230) );
  NAND2_X1 U8841 ( .A1(n7228), .A2(n7229), .ZN(n8100) );
  OR2_X1 U8842 ( .A1(n7228), .A2(n7229), .ZN(n7230) );
  NAND2_X1 U8843 ( .A1(n8100), .A2(n7230), .ZN(n7231) );
  NOR2_X1 U8844 ( .A1(n7231), .A2(n7232), .ZN(n8103) );
  AOI21_X1 U8845 ( .B1(n7232), .B2(n7231), .A(n8103), .ZN(n7239) );
  NOR2_X1 U8846 ( .A1(n8142), .A2(n7233), .ZN(n7234) );
  AOI211_X1 U8847 ( .C1(n8140), .C2(n7236), .A(n7235), .B(n7234), .ZN(n7238)
         );
  NAND2_X1 U8848 ( .A1(n8503), .A2(n8147), .ZN(n7237) );
  OAI211_X1 U8849 ( .C1(n7239), .C2(n8128), .A(n7238), .B(n7237), .ZN(P2_U3243) );
  NAND2_X1 U8850 ( .A1(n7285), .A2(n8709), .ZN(n7240) );
  NAND2_X1 U8851 ( .A1(n7240), .A2(n7286), .ZN(n7244) );
  NAND2_X1 U8852 ( .A1(n7241), .A2(n6363), .ZN(n7243) );
  AOI22_X1 U8853 ( .A1(n7823), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7822), .B2(
        n9543), .ZN(n7242) );
  OR2_X1 U8854 ( .A1(n7302), .A2(n7294), .ZN(n8841) );
  NAND2_X1 U8855 ( .A1(n7302), .A2(n7294), .ZN(n8840) );
  INV_X1 U8856 ( .A(n7263), .ZN(n8913) );
  XNOR2_X1 U8857 ( .A(n7244), .B(n8913), .ZN(n7245) );
  NAND2_X1 U8858 ( .A1(n7245), .A2(n9612), .ZN(n7253) );
  NAND2_X1 U8859 ( .A1(n7983), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7251) );
  INV_X1 U8860 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U8861 ( .A1(n7246), .A2(n8603), .ZN(n7247) );
  AND2_X1 U8862 ( .A1(n7278), .A2(n7247), .ZN(n8604) );
  NAND2_X1 U8863 ( .A1(n5712), .A2(n8604), .ZN(n7250) );
  NAND2_X1 U8864 ( .A1(n7826), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7249) );
  NAND2_X1 U8865 ( .A1(n8735), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7248) );
  NAND4_X1 U8866 ( .A1(n7251), .A2(n7250), .A3(n7249), .A4(n7248), .ZN(n9223)
         );
  AOI22_X1 U8867 ( .A1(n9359), .A2(n8943), .B1(n9357), .B2(n9223), .ZN(n7252)
         );
  NAND2_X1 U8868 ( .A1(n7253), .A2(n7252), .ZN(n9378) );
  INV_X1 U8869 ( .A(n9378), .ZN(n7268) );
  OR2_X2 U8870 ( .A1(n7255), .A2(n7302), .ZN(n7273) );
  INV_X1 U8871 ( .A(n7273), .ZN(n7254) );
  AOI211_X1 U8872 ( .C1(n7302), .C2(n7255), .A(n9680), .B(n7254), .ZN(n9380)
         );
  INV_X1 U8873 ( .A(n7302), .ZN(n9377) );
  AOI22_X1 U8874 ( .A1(n9598), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7301), .B2(
        n9586), .ZN(n7256) );
  OAI21_X1 U8875 ( .B1(n9377), .B2(n9619), .A(n7256), .ZN(n7266) );
  INV_X1 U8876 ( .A(n7258), .ZN(n7259) );
  NAND2_X1 U8877 ( .A1(n9383), .A2(n7257), .ZN(n7262) );
  AND2_X1 U8878 ( .A1(n7264), .A2(n7263), .ZN(n9376) );
  NOR3_X1 U8879 ( .A1(n4337), .A2(n9376), .A3(n9228), .ZN(n7265) );
  AOI211_X1 U8880 ( .C1(n9209), .C2(n9380), .A(n7266), .B(n7265), .ZN(n7267)
         );
  OAI21_X1 U8881 ( .B1(n9598), .B2(n7268), .A(n7267), .ZN(P1_U3275) );
  INV_X1 U8882 ( .A(n7294), .ZN(n8942) );
  NAND2_X1 U8883 ( .A1(n7269), .A2(n6363), .ZN(n7271) );
  AOI22_X1 U8884 ( .A1(n7823), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7822), .B2(
        n9555), .ZN(n7270) );
  INV_X1 U8885 ( .A(n9223), .ZN(n9002) );
  NOR2_X1 U8886 ( .A1(n9299), .A2(n9002), .ZN(n9028) );
  NAND2_X1 U8887 ( .A1(n9299), .A2(n9002), .ZN(n9027) );
  INV_X1 U8888 ( .A(n9027), .ZN(n7272) );
  OR2_X1 U8889 ( .A1(n9028), .A2(n7272), .ZN(n8914) );
  INV_X1 U8890 ( .A(n8914), .ZN(n8843) );
  XNOR2_X1 U8891 ( .A(n9004), .B(n8843), .ZN(n9301) );
  AOI211_X1 U8892 ( .C1(n9299), .C2(n7273), .A(n9680), .B(n9213), .ZN(n9298)
         );
  INV_X1 U8893 ( .A(n9299), .ZN(n9001) );
  NOR2_X1 U8894 ( .A1(n9001), .A2(n9619), .ZN(n7276) );
  INV_X1 U8895 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8979) );
  INV_X1 U8896 ( .A(n8604), .ZN(n7274) );
  OAI22_X1 U8897 ( .A1(n9617), .A2(n8979), .B1(n7274), .B2(n9618), .ZN(n7275)
         );
  AOI211_X1 U8898 ( .C1(n9298), .C2(n9209), .A(n7276), .B(n7275), .ZN(n7289)
         );
  INV_X1 U8899 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U8900 ( .A1(n7278), .A2(n9897), .ZN(n7279) );
  NAND2_X1 U8901 ( .A1(n7829), .A2(n7279), .ZN(n9216) );
  INV_X1 U8902 ( .A(n5712), .ZN(n8020) );
  OR2_X1 U8903 ( .A1(n9216), .A2(n8020), .ZN(n7284) );
  NAND2_X1 U8904 ( .A1(n7983), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7281) );
  NAND2_X1 U8905 ( .A1(n7826), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7280) );
  AND2_X1 U8906 ( .A1(n7281), .A2(n7280), .ZN(n7283) );
  NAND2_X1 U8907 ( .A1(n8735), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n7282) );
  AND3_X1 U8908 ( .A1(n7284), .A2(n7283), .A3(n7282), .ZN(n8718) );
  AND2_X1 U8909 ( .A1(n8840), .A2(n8709), .ZN(n8837) );
  NAND2_X1 U8910 ( .A1(n8841), .A2(n7286), .ZN(n8835) );
  XNOR2_X1 U8911 ( .A(n9029), .B(n8843), .ZN(n7287) );
  OAI222_X1 U8912 ( .A1(n9610), .A2(n8718), .B1(n9608), .B2(n7294), .C1(n9591), 
        .C2(n7287), .ZN(n9297) );
  NAND2_X1 U8913 ( .A1(n9297), .A2(n9617), .ZN(n7288) );
  OAI211_X1 U8914 ( .C1(n9301), .C2(n9228), .A(n7289), .B(n7288), .ZN(P1_U3274) );
  NAND2_X1 U8915 ( .A1(n7302), .A2(n4265), .ZN(n7293) );
  NAND2_X1 U8916 ( .A1(n7974), .A2(n8942), .ZN(n7292) );
  NAND2_X1 U8917 ( .A1(n7293), .A2(n7292), .ZN(n7798) );
  NAND2_X1 U8918 ( .A1(n7302), .A2(n7995), .ZN(n7296) );
  OR2_X1 U8919 ( .A1(n7294), .A2(n6180), .ZN(n7295) );
  NAND2_X1 U8920 ( .A1(n7296), .A2(n7295), .ZN(n7297) );
  XNOR2_X1 U8921 ( .A(n7297), .B(n7989), .ZN(n7799) );
  XOR2_X1 U8922 ( .A(n7798), .B(n7799), .Z(n7298) );
  XNOR2_X1 U8923 ( .A(n7800), .B(n7298), .ZN(n7305) );
  NAND2_X1 U8924 ( .A1(n8633), .A2(n8943), .ZN(n7299) );
  NAND2_X1 U8925 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9537) );
  OAI211_X1 U8926 ( .C1(n9002), .C2(n8657), .A(n7299), .B(n9537), .ZN(n7300)
         );
  AOI21_X1 U8927 ( .B1(n7301), .B2(n8660), .A(n7300), .ZN(n7304) );
  NAND2_X1 U8928 ( .A1(n7302), .A2(n8648), .ZN(n7303) );
  OAI211_X1 U8929 ( .C1(n7305), .C2(n8650), .A(n7304), .B(n7303), .ZN(P1_U3224) );
  INV_X1 U8930 ( .A(n7306), .ZN(n7309) );
  INV_X1 U8931 ( .A(n7307), .ZN(n7308) );
  NAND2_X1 U8932 ( .A1(n7808), .A2(n5954), .ZN(n7314) );
  AOI22_X1 U8933 ( .A1(n7339), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7338), .B2(
        n7312), .ZN(n7313) );
  XNOR2_X1 U8934 ( .A(n8487), .B(n7439), .ZN(n7333) );
  NOR2_X1 U8935 ( .A1(n8074), .A2(n6325), .ZN(n7334) );
  XNOR2_X1 U8936 ( .A(n7333), .B(n7334), .ZN(n7331) );
  XNOR2_X1 U8937 ( .A(n7332), .B(n7331), .ZN(n7328) );
  INV_X1 U8938 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7316) );
  INV_X1 U8939 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7315) );
  OAI21_X1 U8940 ( .B1(n7318), .B2(n7316), .A(n7315), .ZN(n7319) );
  NAND2_X1 U8941 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n7317) );
  AND2_X1 U8942 ( .A1(n7319), .A2(n7352), .ZN(n8351) );
  NAND2_X1 U8943 ( .A1(n8351), .A2(n7518), .ZN(n7323) );
  AOI22_X1 U8944 ( .A1(n5609), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n7525), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n7322) );
  NAND2_X1 U8945 ( .A1(n4279), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7321) );
  AND3_X1 U8946 ( .A1(n7323), .A2(n7322), .A3(n7321), .ZN(n8329) );
  OAI22_X1 U8947 ( .A1(n8135), .A2(n8105), .B1(n8329), .B2(n9714), .ZN(n7324)
         );
  AOI211_X1 U8948 ( .C1(n8140), .C2(n8366), .A(n7325), .B(n7324), .ZN(n7327)
         );
  NAND2_X1 U8949 ( .A1(n8487), .A2(n8147), .ZN(n7326) );
  OAI211_X1 U8950 ( .C1(n7328), .C2(n8128), .A(n7327), .B(n7326), .ZN(P2_U3240) );
  XNOR2_X1 U8951 ( .A(n7330), .B(n7329), .ZN(n7886) );
  INV_X1 U8952 ( .A(n7886), .ZN(n8038) );
  OAI222_X1 U8953 ( .A1(n8545), .A2(n7377), .B1(n4270), .B2(n8038), .C1(
        P2_U3152), .C2(n5119), .ZN(P2_U3336) );
  NAND2_X1 U8954 ( .A1(n7332), .A2(n7331), .ZN(n7337) );
  INV_X1 U8955 ( .A(n7333), .ZN(n7335) );
  NAND2_X1 U8956 ( .A1(n7335), .A2(n7334), .ZN(n7336) );
  NAND2_X1 U8957 ( .A1(n7821), .A2(n5954), .ZN(n7341) );
  AOI22_X1 U8958 ( .A1(n7339), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7338), .B2(
        n8253), .ZN(n7340) );
  XNOR2_X1 U8959 ( .A(n8483), .B(n7439), .ZN(n7342) );
  OR2_X1 U8960 ( .A1(n8329), .A2(n6325), .ZN(n7343) );
  NAND2_X1 U8961 ( .A1(n7342), .A2(n7343), .ZN(n7347) );
  INV_X1 U8962 ( .A(n7342), .ZN(n7345) );
  INV_X1 U8963 ( .A(n7343), .ZN(n7344) );
  NAND2_X1 U8964 ( .A1(n7345), .A2(n7344), .ZN(n7346) );
  NAND2_X1 U8965 ( .A1(n7347), .A2(n7346), .ZN(n8073) );
  NAND2_X1 U8966 ( .A1(n7844), .A2(n5954), .ZN(n7350) );
  OR2_X1 U8967 ( .A1(n7540), .A2(n7348), .ZN(n7349) );
  XNOR2_X1 U8968 ( .A(n8477), .B(n7439), .ZN(n7370) );
  INV_X1 U8969 ( .A(n7352), .ZN(n7351) );
  NAND2_X1 U8970 ( .A1(n7351), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7359) );
  INV_X1 U8971 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U8972 ( .A1(n7352), .A2(n9967), .ZN(n7353) );
  NAND2_X1 U8973 ( .A1(n7359), .A2(n7353), .ZN(n8341) );
  OR2_X1 U8974 ( .A1(n8341), .A2(n7472), .ZN(n7356) );
  AOI22_X1 U8975 ( .A1(n5609), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n7525), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U8976 ( .A1(n4279), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7354) );
  AND3_X1 U8977 ( .A1(n7356), .A2(n7355), .A3(n7354), .ZN(n8085) );
  INV_X1 U8978 ( .A(n8085), .ZN(n8359) );
  NAND2_X1 U8979 ( .A1(n8359), .A2(n8041), .ZN(n7371) );
  XNOR2_X1 U8980 ( .A(n7370), .B(n7371), .ZN(n8124) );
  OR2_X1 U8981 ( .A1(n7540), .A2(n7357), .ZN(n7358) );
  XNOR2_X1 U8982 ( .A(n8471), .B(n7439), .ZN(n7368) );
  INV_X1 U8983 ( .A(n7368), .ZN(n7366) );
  INV_X1 U8984 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U8985 ( .A1(n7359), .A2(n9905), .ZN(n7360) );
  AND2_X1 U8986 ( .A1(n7382), .A2(n7360), .ZN(n8321) );
  NAND2_X1 U8987 ( .A1(n8321), .A2(n7518), .ZN(n7365) );
  INV_X1 U8988 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U8989 ( .A1(n5609), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7362) );
  NAND2_X1 U8990 ( .A1(n7525), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7361) );
  OAI211_X1 U8991 ( .C1(n8315), .C2(n7529), .A(n7362), .B(n7361), .ZN(n7363)
         );
  INV_X1 U8992 ( .A(n7363), .ZN(n7364) );
  AND2_X1 U8993 ( .A1(n7365), .A2(n7364), .ZN(n8331) );
  NOR2_X1 U8994 ( .A1(n8331), .A2(n6325), .ZN(n7367) );
  NAND2_X1 U8995 ( .A1(n7366), .A2(n7367), .ZN(n7374) );
  INV_X1 U8996 ( .A(n7374), .ZN(n7369) );
  XNOR2_X1 U8997 ( .A(n7368), .B(n7367), .ZN(n8082) );
  INV_X1 U8998 ( .A(n7370), .ZN(n7373) );
  INV_X1 U8999 ( .A(n7371), .ZN(n7372) );
  NAND2_X1 U9000 ( .A1(n7373), .A2(n7372), .ZN(n8080) );
  AND2_X1 U9001 ( .A1(n8080), .A2(n7374), .ZN(n7375) );
  NAND2_X1 U9002 ( .A1(n7886), .A2(n5954), .ZN(n7379) );
  OR2_X1 U9003 ( .A1(n7540), .A2(n7377), .ZN(n7378) );
  XNOR2_X1 U9004 ( .A(n8466), .B(n7439), .ZN(n7391) );
  XNOR2_X1 U9005 ( .A(n7390), .B(n7391), .ZN(n8132) );
  INV_X1 U9006 ( .A(n7382), .ZN(n7380) );
  NAND2_X1 U9007 ( .A1(n7380), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n7407) );
  INV_X1 U9008 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7381) );
  NAND2_X1 U9009 ( .A1(n7382), .A2(n7381), .ZN(n7383) );
  NAND2_X1 U9010 ( .A1(n7407), .A2(n7383), .ZN(n8299) );
  OR2_X1 U9011 ( .A1(n8299), .A2(n7472), .ZN(n7389) );
  INV_X1 U9012 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U9013 ( .A1(n7525), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7385) );
  NAND2_X1 U9014 ( .A1(n5609), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7384) );
  OAI211_X1 U9015 ( .C1(n7529), .C2(n7386), .A(n7385), .B(n7384), .ZN(n7387)
         );
  INV_X1 U9016 ( .A(n7387), .ZN(n7388) );
  AND2_X1 U9017 ( .A1(n7389), .A2(n7388), .ZN(n8283) );
  INV_X1 U9018 ( .A(n8283), .ZN(n8319) );
  NAND2_X1 U9019 ( .A1(n8319), .A2(n8041), .ZN(n8131) );
  NAND2_X1 U9020 ( .A1(n8132), .A2(n8131), .ZN(n8130) );
  INV_X1 U9021 ( .A(n7390), .ZN(n7392) );
  NAND2_X1 U9022 ( .A1(n7392), .A2(n7391), .ZN(n7393) );
  NAND2_X1 U9023 ( .A1(n7906), .A2(n5954), .ZN(n7396) );
  OR2_X1 U9024 ( .A1(n7540), .A2(n7394), .ZN(n7395) );
  NAND2_X1 U9025 ( .A1(n7924), .A2(n5954), .ZN(n7399) );
  OR2_X1 U9026 ( .A1(n7540), .A2(n7397), .ZN(n7398) );
  INV_X1 U9027 ( .A(n8116), .ZN(n7415) );
  INV_X1 U9028 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8065) );
  INV_X1 U9029 ( .A(n7409), .ZN(n7400) );
  NAND2_X1 U9030 ( .A1(n7400), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7426) );
  INV_X1 U9031 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U9032 ( .A1(n7409), .A2(n9910), .ZN(n7401) );
  NAND2_X1 U9033 ( .A1(n7426), .A2(n7401), .ZN(n8262) );
  OR2_X1 U9034 ( .A1(n8262), .A2(n7472), .ZN(n7406) );
  INV_X1 U9035 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9908) );
  NAND2_X1 U9036 ( .A1(n7525), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7403) );
  NAND2_X1 U9037 ( .A1(n5595), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7402) );
  OAI211_X1 U9038 ( .C1(n7458), .C2(n9908), .A(n7403), .B(n7402), .ZN(n7404)
         );
  INV_X1 U9039 ( .A(n7404), .ZN(n7405) );
  INV_X1 U9040 ( .A(n8284), .ZN(n7414) );
  NAND2_X1 U9041 ( .A1(n7407), .A2(n8065), .ZN(n7408) );
  AND2_X1 U9042 ( .A1(n7409), .A2(n7408), .ZN(n8064) );
  INV_X1 U9043 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U9044 ( .A1(n5609), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n7411) );
  NAND2_X1 U9045 ( .A1(n7525), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7410) );
  OAI211_X1 U9046 ( .C1(n8290), .C2(n7529), .A(n7411), .B(n7410), .ZN(n7412)
         );
  AOI21_X1 U9047 ( .B1(n8064), .B2(n7518), .A(n7412), .ZN(n8134) );
  OR2_X1 U9048 ( .A1(n8134), .A2(n6325), .ZN(n8114) );
  INV_X1 U9049 ( .A(n8114), .ZN(n7413) );
  OAI21_X1 U9050 ( .B1(n7415), .B2(n7414), .A(n7413), .ZN(n7416) );
  NOR2_X1 U9051 ( .A1(n7417), .A2(n4816), .ZN(n8112) );
  NOR2_X1 U9052 ( .A1(n8284), .A2(n6325), .ZN(n8115) );
  INV_X1 U9053 ( .A(n8115), .ZN(n7418) );
  NAND2_X1 U9054 ( .A1(n8116), .A2(n7418), .ZN(n7420) );
  AOI21_X1 U9055 ( .B1(n8112), .B2(n7420), .A(n7419), .ZN(n7421) );
  OR2_X1 U9056 ( .A1(n7540), .A2(n7423), .ZN(n7424) );
  INV_X1 U9057 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U9058 ( .A1(n7426), .A2(n8095), .ZN(n7427) );
  NAND2_X1 U9059 ( .A1(n7441), .A2(n7427), .ZN(n8252) );
  OR2_X1 U9060 ( .A1(n8252), .A2(n7472), .ZN(n7432) );
  INV_X1 U9061 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U9062 ( .A1(n4279), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7429) );
  NAND2_X1 U9063 ( .A1(n7525), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7428) );
  OAI211_X1 U9064 ( .C1(n7458), .C2(n9969), .A(n7429), .B(n7428), .ZN(n7430)
         );
  INV_X1 U9065 ( .A(n7430), .ZN(n7431) );
  INV_X1 U9066 ( .A(n8119), .ZN(n8269) );
  NAND2_X1 U9067 ( .A1(n8269), .A2(n8041), .ZN(n8090) );
  OAI21_X1 U9068 ( .B1(n10043), .B2(n8091), .A(n8090), .ZN(n7435) );
  NAND2_X1 U9069 ( .A1(n7435), .A2(n7434), .ZN(n8144) );
  NAND2_X1 U9070 ( .A1(n7959), .A2(n5954), .ZN(n7438) );
  OR2_X1 U9071 ( .A1(n7540), .A2(n7436), .ZN(n7437) );
  XNOR2_X1 U9072 ( .A(n8240), .B(n7439), .ZN(n7450) );
  INV_X1 U9073 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U9074 ( .A1(n7441), .A2(n7440), .ZN(n7442) );
  AND2_X1 U9075 ( .A1(n7470), .A2(n7442), .ZN(n8237) );
  NAND2_X1 U9076 ( .A1(n8237), .A2(n7518), .ZN(n7448) );
  INV_X1 U9077 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U9078 ( .A1(n5609), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7444) );
  NAND2_X1 U9079 ( .A1(n4279), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7443) );
  OAI211_X1 U9080 ( .C1(n7445), .C2(n9984), .A(n7444), .B(n7443), .ZN(n7446)
         );
  INV_X1 U9081 ( .A(n7446), .ZN(n7447) );
  NAND2_X1 U9082 ( .A1(n7448), .A2(n7447), .ZN(n8216) );
  AND2_X1 U9083 ( .A1(n8216), .A2(n8041), .ZN(n7449) );
  NAND2_X1 U9084 ( .A1(n7450), .A2(n7449), .ZN(n7451) );
  OAI21_X1 U9085 ( .B1(n7450), .B2(n7449), .A(n7451), .ZN(n8145) );
  INV_X1 U9086 ( .A(n7451), .ZN(n7452) );
  OR2_X1 U9087 ( .A1(n7540), .A2(n7453), .ZN(n7454) );
  XNOR2_X1 U9088 ( .A(n8440), .B(n8043), .ZN(n7463) );
  XNOR2_X1 U9089 ( .A(n7470), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U9090 ( .A1(n8211), .A2(n7518), .ZN(n7461) );
  INV_X1 U9091 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U9092 ( .A1(n4279), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7457) );
  NAND2_X1 U9093 ( .A1(n7525), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7456) );
  OAI211_X1 U9094 ( .C1(n7458), .C2(n9981), .A(n7457), .B(n7456), .ZN(n7459)
         );
  INV_X1 U9095 ( .A(n7459), .ZN(n7460) );
  NAND2_X1 U9096 ( .A1(n7461), .A2(n7460), .ZN(n8200) );
  AND2_X1 U9097 ( .A1(n8200), .A2(n8041), .ZN(n7462) );
  NAND2_X1 U9098 ( .A1(n7463), .A2(n7462), .ZN(n8040) );
  OAI21_X1 U9099 ( .B1(n7463), .B2(n7462), .A(n8040), .ZN(n7465) );
  AOI21_X1 U9100 ( .B1(n4331), .B2(n7465), .A(n8128), .ZN(n7464) );
  INV_X1 U9101 ( .A(n7464), .ZN(n7483) );
  INV_X1 U9102 ( .A(n8216), .ZN(n7506) );
  INV_X1 U9103 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7469) );
  OAI22_X1 U9104 ( .A1(n7506), .A2(n8135), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7469), .ZN(n7481) );
  INV_X1 U9105 ( .A(n7470), .ZN(n7467) );
  AND2_X1 U9106 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n7466) );
  NAND2_X1 U9107 ( .A1(n7467), .A2(n7466), .ZN(n7517) );
  INV_X1 U9108 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7468) );
  OAI21_X1 U9109 ( .B1(n7470), .B2(n7469), .A(n7468), .ZN(n7471) );
  NAND2_X1 U9110 ( .A1(n7517), .A2(n7471), .ZN(n8047) );
  OR2_X1 U9111 ( .A1(n8047), .A2(n7472), .ZN(n7478) );
  INV_X1 U9112 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7475) );
  NAND2_X1 U9113 ( .A1(n5609), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U9114 ( .A1(n7525), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7473) );
  OAI211_X1 U9115 ( .C1(n7475), .C2(n7529), .A(n7474), .B(n7473), .ZN(n7476)
         );
  INV_X1 U9116 ( .A(n7476), .ZN(n7477) );
  INV_X1 U9117 ( .A(n8211), .ZN(n7479) );
  OAI22_X1 U9118 ( .A1(n7779), .A2(n9714), .B1(n7479), .B2(n9737), .ZN(n7480)
         );
  AOI211_X1 U9119 ( .C1(n8440), .C2(n8147), .A(n7481), .B(n7480), .ZN(n7482)
         );
  OAI21_X1 U9120 ( .B1(n7483), .B2(n4324), .A(n7482), .ZN(P2_U3216) );
  INV_X1 U9121 ( .A(n7484), .ZN(n7486) );
  NOR2_X1 U9122 ( .A1(n7486), .A2(n7485), .ZN(n7489) );
  AOI21_X1 U9123 ( .B1(n7489), .B2(n7487), .A(n7488), .ZN(n7492) );
  AOI22_X1 U9124 ( .A1(n8633), .A2(n5462), .B1(n8644), .B2(n8953), .ZN(n7491)
         );
  AOI22_X1 U9125 ( .A1(n8648), .A2(n6022), .B1(n8580), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7490) );
  OAI211_X1 U9126 ( .C1(n7492), .C2(n8650), .A(n7491), .B(n7490), .ZN(P1_U3235) );
  INV_X1 U9127 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8544) );
  INV_X1 U9128 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9327) );
  MUX2_X1 U9129 ( .A(n8544), .B(n9327), .S(n7537), .Z(n7497) );
  XNOR2_X1 U9130 ( .A(n7497), .B(SI_28_), .ZN(n7509) );
  INV_X1 U9131 ( .A(SI_28_), .ZN(n7496) );
  INV_X1 U9132 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9896) );
  INV_X1 U9133 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9322) );
  MUX2_X1 U9134 ( .A(n9896), .B(n9322), .S(n4276), .Z(n7513) );
  INV_X1 U9135 ( .A(n7513), .ZN(n7498) );
  NOR2_X1 U9136 ( .A1(n7498), .A2(SI_29_), .ZN(n7500) );
  NAND2_X1 U9137 ( .A1(n7498), .A2(SI_29_), .ZN(n7499) );
  MUX2_X1 U9138 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7537), .Z(n7534) );
  NAND2_X1 U9139 ( .A1(n8730), .A2(n5954), .ZN(n7502) );
  INV_X1 U9140 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8060) );
  OR2_X1 U9141 ( .A1(n7540), .A2(n8060), .ZN(n7501) );
  NAND2_X1 U9142 ( .A1(n8493), .A2(n8105), .ZN(n7638) );
  NAND2_X1 U9143 ( .A1(n7637), .A2(n7638), .ZN(n7766) );
  OR2_X1 U9144 ( .A1(n8487), .A2(n8074), .ZN(n7646) );
  NAND2_X1 U9145 ( .A1(n8487), .A2(n8074), .ZN(n7652) );
  OR2_X1 U9146 ( .A1(n8483), .A2(n8329), .ZN(n7650) );
  NAND2_X1 U9147 ( .A1(n8483), .A2(n8329), .ZN(n7654) );
  NAND2_X1 U9148 ( .A1(n7650), .A2(n7654), .ZN(n8354) );
  INV_X1 U9149 ( .A(n7646), .ZN(n8355) );
  NOR2_X1 U9150 ( .A1(n8354), .A2(n8355), .ZN(n7504) );
  NAND2_X1 U9151 ( .A1(n8477), .A2(n8085), .ZN(n7655) );
  INV_X1 U9152 ( .A(n8335), .ZN(n7505) );
  OR2_X1 U9153 ( .A1(n8471), .A2(n8331), .ZN(n7657) );
  NAND2_X1 U9154 ( .A1(n8471), .A2(n8331), .ZN(n7665) );
  NAND2_X1 U9155 ( .A1(n7657), .A2(n7665), .ZN(n8318) );
  NAND2_X1 U9156 ( .A1(n8466), .A2(n8283), .ZN(n7667) );
  XNOR2_X1 U9157 ( .A(n8293), .B(n8134), .ZN(n8279) );
  INV_X1 U9158 ( .A(n8134), .ZN(n8306) );
  NOR2_X1 U9159 ( .A1(n8460), .A2(n8306), .ZN(n7674) );
  NAND2_X1 U9160 ( .A1(n8454), .A2(n8284), .ZN(n7676) );
  NAND2_X1 U9161 ( .A1(n8213), .A2(n7508), .ZN(n8198) );
  OR2_X1 U9162 ( .A1(n7540), .A2(n8544), .ZN(n7511) );
  NAND2_X1 U9163 ( .A1(n8435), .A2(n7779), .ZN(n7694) );
  XNOR2_X1 U9164 ( .A(n7513), .B(SI_29_), .ZN(n7514) );
  NOR2_X1 U9165 ( .A1(n7540), .A2(n9896), .ZN(n7516) );
  INV_X1 U9166 ( .A(n7517), .ZN(n7785) );
  NAND2_X1 U9167 ( .A1(n7785), .A2(n7518), .ZN(n7524) );
  INV_X1 U9168 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7521) );
  NAND2_X1 U9169 ( .A1(n7525), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U9170 ( .A1(n5609), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7519) );
  OAI211_X1 U9171 ( .C1(n7521), .C2(n7529), .A(n7520), .B(n7519), .ZN(n7522)
         );
  INV_X1 U9172 ( .A(n7522), .ZN(n7523) );
  NAND2_X1 U9173 ( .A1(n7524), .A2(n7523), .ZN(n8199) );
  AND2_X1 U9174 ( .A1(n7787), .A2(n8199), .ZN(n7693) );
  INV_X1 U9175 ( .A(n7787), .ZN(n8430) );
  INV_X1 U9176 ( .A(n8199), .ZN(n8050) );
  NAND2_X1 U9177 ( .A1(n8430), .A2(n8050), .ZN(n7699) );
  INV_X1 U9178 ( .A(n7530), .ZN(n7532) );
  INV_X1 U9179 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U9180 ( .A1(n7525), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U9181 ( .A1(n5609), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7526) );
  OAI211_X1 U9182 ( .C1(n7529), .C2(n7528), .A(n7527), .B(n7526), .ZN(n8148)
         );
  NAND2_X1 U9183 ( .A1(n9343), .A2(n8148), .ZN(n7706) );
  AOI21_X1 U9184 ( .B1(n9343), .B2(n7532), .A(n7531), .ZN(n7547) );
  NAND2_X1 U9185 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  MUX2_X1 U9186 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7537), .Z(n7538) );
  XNOR2_X1 U9187 ( .A(n7538), .B(SI_31_), .ZN(n7539) );
  NAND2_X1 U9188 ( .A1(n8743), .A2(n5954), .ZN(n7542) );
  OR2_X1 U9189 ( .A1(n7540), .A2(n5037), .ZN(n7541) );
  INV_X1 U9190 ( .A(n8148), .ZN(n7545) );
  NAND2_X1 U9191 ( .A1(n8185), .A2(n7545), .ZN(n7701) );
  NAND2_X1 U9192 ( .A1(n7709), .A2(n7701), .ZN(n7550) );
  NAND2_X1 U9193 ( .A1(n8427), .A2(n7546), .ZN(n7707) );
  OAI21_X1 U9194 ( .B1(n7547), .B2(n7550), .A(n7707), .ZN(n7548) );
  XNOR2_X1 U9195 ( .A(n7548), .B(n8253), .ZN(n7754) );
  INV_X1 U9196 ( .A(n7550), .ZN(n7741) );
  AND3_X1 U9197 ( .A1(n5119), .A2(n8253), .A3(n5118), .ZN(n7697) );
  INV_X1 U9198 ( .A(n7706), .ZN(n7705) );
  OAI21_X1 U9199 ( .B1(n7697), .B2(n8246), .A(n4730), .ZN(n7688) );
  INV_X1 U9200 ( .A(n8267), .ZN(n8258) );
  NOR2_X1 U9201 ( .A1(n8293), .A2(n8134), .ZN(n7551) );
  OAI21_X1 U9202 ( .B1(n8258), .B2(n7551), .A(n7697), .ZN(n7673) );
  INV_X1 U9203 ( .A(n7552), .ZN(n7555) );
  INV_X1 U9204 ( .A(n7553), .ZN(n7554) );
  MUX2_X1 U9205 ( .A(n7555), .B(n7554), .S(n7697), .Z(n7556) );
  NOR2_X1 U9206 ( .A1(n7733), .A2(n7556), .ZN(n7636) );
  AND2_X1 U9207 ( .A1(n7559), .A2(n7560), .ZN(n7557) );
  MUX2_X1 U9208 ( .A(n7605), .B(n7557), .S(n7697), .Z(n7558) );
  NAND2_X1 U9209 ( .A1(n7558), .A2(n7561), .ZN(n7564) );
  OAI211_X1 U9210 ( .C1(n7564), .C2(n7560), .A(n7610), .B(n7559), .ZN(n7563)
         );
  NAND2_X1 U9211 ( .A1(n7609), .A2(n7561), .ZN(n7562) );
  MUX2_X1 U9212 ( .A(n7563), .B(n7562), .S(n7697), .Z(n7616) );
  INV_X1 U9213 ( .A(n7564), .ZN(n7608) );
  NAND2_X1 U9214 ( .A1(n7569), .A2(n7567), .ZN(n7566) );
  NAND2_X1 U9215 ( .A1(n7591), .A2(n7589), .ZN(n7565) );
  MUX2_X1 U9216 ( .A(n7566), .B(n7565), .S(n7710), .Z(n7593) );
  AND2_X1 U9217 ( .A1(n7568), .A2(n7567), .ZN(n7570) );
  OAI211_X1 U9218 ( .C1(n7593), .C2(n7570), .A(n7569), .B(n4296), .ZN(n7571)
         );
  NAND2_X1 U9219 ( .A1(n7571), .A2(n7710), .ZN(n7579) );
  INV_X1 U9220 ( .A(n7593), .ZN(n7577) );
  AND2_X1 U9221 ( .A1(n7716), .A2(n5118), .ZN(n7573) );
  OAI211_X1 U9222 ( .C1(n7573), .C2(n7572), .A(n7583), .B(n8410), .ZN(n7574)
         );
  NAND3_X1 U9223 ( .A1(n7574), .A2(n7581), .A3(n7710), .ZN(n7575) );
  NAND3_X1 U9224 ( .A1(n7577), .A2(n7576), .A3(n7575), .ZN(n7578) );
  NAND2_X1 U9225 ( .A1(n7579), .A2(n7578), .ZN(n7596) );
  NAND2_X1 U9226 ( .A1(n8410), .A2(n7716), .ZN(n7582) );
  NAND3_X1 U9227 ( .A1(n7582), .A2(n7581), .A3(n7580), .ZN(n7587) );
  AND2_X1 U9228 ( .A1(n7583), .A2(n7697), .ZN(n7586) );
  NAND2_X1 U9229 ( .A1(n7584), .A2(n8156), .ZN(n7590) );
  INV_X1 U9230 ( .A(n7590), .ZN(n7585) );
  AOI21_X1 U9231 ( .B1(n7587), .B2(n7586), .A(n7585), .ZN(n7595) );
  AND2_X1 U9232 ( .A1(n7589), .A2(n7588), .ZN(n7592) );
  OAI211_X1 U9233 ( .C1(n7593), .C2(n7592), .A(n7591), .B(n7590), .ZN(n7594)
         );
  AOI22_X1 U9234 ( .A1(n7596), .A2(n7595), .B1(n7697), .B2(n7594), .ZN(n7601)
         );
  OAI21_X1 U9235 ( .B1(n4296), .B2(n7710), .A(n7722), .ZN(n7600) );
  MUX2_X1 U9236 ( .A(n7598), .B(n7597), .S(n7697), .Z(n7599) );
  OAI211_X1 U9237 ( .C1(n7601), .C2(n7600), .A(n4266), .B(n7599), .ZN(n7606)
         );
  MUX2_X1 U9238 ( .A(n7603), .B(n7602), .S(n7710), .Z(n7604) );
  NAND3_X1 U9239 ( .A1(n7606), .A2(n7605), .A3(n7604), .ZN(n7607) );
  AND2_X1 U9240 ( .A1(n7608), .A2(n7607), .ZN(n7615) );
  NAND2_X1 U9241 ( .A1(n4301), .A2(n7609), .ZN(n7612) );
  NAND2_X1 U9242 ( .A1(n7617), .A2(n7610), .ZN(n7611) );
  MUX2_X1 U9243 ( .A(n7612), .B(n7611), .S(n7697), .Z(n7613) );
  INV_X1 U9244 ( .A(n7613), .ZN(n7614) );
  OAI21_X1 U9245 ( .B1(n7616), .B2(n7615), .A(n7614), .ZN(n7619) );
  MUX2_X1 U9246 ( .A(n7617), .B(n4301), .S(n7697), .Z(n7618) );
  NAND3_X1 U9247 ( .A1(n7619), .A2(n7730), .A3(n7618), .ZN(n7627) );
  INV_X1 U9248 ( .A(n7620), .ZN(n7623) );
  INV_X1 U9249 ( .A(n7621), .ZN(n7622) );
  MUX2_X1 U9250 ( .A(n7623), .B(n7622), .S(n7697), .Z(n7624) );
  NOR2_X1 U9251 ( .A1(n7625), .A2(n7624), .ZN(n7626) );
  NAND2_X1 U9252 ( .A1(n7627), .A2(n7626), .ZN(n7631) );
  MUX2_X1 U9253 ( .A(n7629), .B(n7628), .S(n7697), .Z(n7630) );
  NAND3_X1 U9254 ( .A1(n7632), .A2(n7631), .A3(n7630), .ZN(n7635) );
  INV_X1 U9255 ( .A(n7633), .ZN(n7634) );
  AOI22_X1 U9256 ( .A1(n7636), .A2(n7635), .B1(n7634), .B2(n7710), .ZN(n7644)
         );
  INV_X1 U9257 ( .A(n7637), .ZN(n7641) );
  OAI211_X1 U9258 ( .C1(n7766), .C2(n7639), .A(n7638), .B(n7652), .ZN(n7640)
         );
  MUX2_X1 U9259 ( .A(n7641), .B(n7640), .S(n7697), .Z(n7642) );
  INV_X1 U9260 ( .A(n7642), .ZN(n7643) );
  OAI21_X1 U9261 ( .B1(n7644), .B2(n7766), .A(n7643), .ZN(n7653) );
  INV_X1 U9262 ( .A(n7654), .ZN(n7645) );
  AOI21_X1 U9263 ( .B1(n7653), .B2(n7646), .A(n7645), .ZN(n7648) );
  NAND2_X1 U9264 ( .A1(n7656), .A2(n7650), .ZN(n7647) );
  OAI211_X1 U9265 ( .C1(n7648), .C2(n7647), .A(n7665), .B(n7655), .ZN(n7649)
         );
  NAND3_X1 U9266 ( .A1(n7649), .A2(n7697), .A3(n7668), .ZN(n7663) );
  INV_X1 U9267 ( .A(n7663), .ZN(n7666) );
  INV_X1 U9268 ( .A(n7657), .ZN(n7662) );
  INV_X1 U9269 ( .A(n7650), .ZN(n7651) );
  AOI211_X1 U9270 ( .C1(n7653), .C2(n7652), .A(n8355), .B(n7651), .ZN(n7659)
         );
  NAND2_X1 U9271 ( .A1(n7655), .A2(n7654), .ZN(n7658) );
  OAI211_X1 U9272 ( .C1(n7659), .C2(n7658), .A(n7657), .B(n7656), .ZN(n7660)
         );
  NAND3_X1 U9273 ( .A1(n7660), .A2(n7667), .A3(n7710), .ZN(n7661) );
  OAI21_X1 U9274 ( .B1(n7663), .B2(n7662), .A(n7661), .ZN(n7664) );
  OAI21_X1 U9275 ( .B1(n7666), .B2(n7665), .A(n7664), .ZN(n7670) );
  MUX2_X1 U9276 ( .A(n7668), .B(n7667), .S(n7697), .Z(n7669) );
  NAND3_X1 U9277 ( .A1(n7670), .A2(n8275), .A3(n7669), .ZN(n7672) );
  INV_X1 U9278 ( .A(n7676), .ZN(n7671) );
  AOI21_X1 U9279 ( .B1(n7673), .B2(n7672), .A(n7671), .ZN(n7678) );
  INV_X1 U9280 ( .A(n7674), .ZN(n7675) );
  AOI21_X1 U9281 ( .B1(n7676), .B2(n7675), .A(n7697), .ZN(n7677) );
  INV_X1 U9282 ( .A(n8247), .ZN(n7737) );
  OAI21_X1 U9283 ( .B1(n7678), .B2(n7677), .A(n7737), .ZN(n7687) );
  OAI21_X1 U9284 ( .B1(n7679), .B2(n8269), .A(n7682), .ZN(n7680) );
  NAND2_X1 U9285 ( .A1(n7680), .A2(n7681), .ZN(n7685) );
  INV_X1 U9286 ( .A(n7681), .ZN(n7683) );
  OAI21_X1 U9287 ( .B1(n7683), .B2(n8227), .A(n7682), .ZN(n7684) );
  MUX2_X1 U9288 ( .A(n7685), .B(n7684), .S(n7697), .Z(n7686) );
  OAI21_X1 U9289 ( .B1(n7688), .B2(n7687), .A(n7686), .ZN(n7692) );
  NOR2_X1 U9290 ( .A1(n7777), .A2(n7710), .ZN(n7690) );
  NOR2_X1 U9291 ( .A1(n8200), .A2(n7697), .ZN(n7689) );
  MUX2_X1 U9292 ( .A(n7690), .B(n7689), .S(n8440), .Z(n7691) );
  INV_X1 U9293 ( .A(n8197), .ZN(n8190) );
  AOI211_X1 U9294 ( .C1(n7692), .C2(n8214), .A(n7691), .B(n8190), .ZN(n7703)
         );
  INV_X1 U9295 ( .A(n7693), .ZN(n7698) );
  MUX2_X1 U9296 ( .A(n7695), .B(n7694), .S(n7697), .Z(n7696) );
  NAND2_X1 U9297 ( .A1(n7782), .A2(n7696), .ZN(n7702) );
  MUX2_X1 U9298 ( .A(n7699), .B(n7698), .S(n7697), .Z(n7700) );
  OAI211_X1 U9299 ( .C1(n7703), .C2(n7702), .A(n7701), .B(n7700), .ZN(n7704)
         );
  OAI22_X1 U9300 ( .A1(n7741), .A2(n7710), .B1(n7705), .B2(n7704), .ZN(n7708)
         );
  NAND2_X1 U9301 ( .A1(n7707), .A2(n7706), .ZN(n7714) );
  AOI22_X1 U9302 ( .A1(n7708), .A2(n7707), .B1(n7710), .B2(n7714), .ZN(n7713)
         );
  INV_X1 U9303 ( .A(n7709), .ZN(n7711) );
  INV_X1 U9304 ( .A(n7745), .ZN(n7751) );
  OAI21_X1 U9305 ( .B1(n7744), .B2(n5740), .A(n9781), .ZN(n7750) );
  INV_X1 U9306 ( .A(n7714), .ZN(n7742) );
  INV_X1 U9307 ( .A(n8354), .ZN(n7735) );
  NOR2_X1 U9308 ( .A1(n7572), .A2(n7715), .ZN(n7717) );
  NAND4_X1 U9309 ( .A1(n7717), .A2(n7744), .A3(n7716), .A4(n8410), .ZN(n7720)
         );
  NOR4_X1 U9310 ( .A1(n7720), .A2(n7719), .A3(n6140), .A4(n7718), .ZN(n7723)
         );
  NAND4_X1 U9311 ( .A1(n7723), .A2(n7722), .A3(n4266), .A4(n7721), .ZN(n7725)
         );
  NOR4_X1 U9312 ( .A1(n7727), .A2(n7726), .A3(n7725), .A4(n6531), .ZN(n7728)
         );
  NAND4_X1 U9313 ( .A1(n7021), .A2(n7730), .A3(n7729), .A4(n7728), .ZN(n7731)
         );
  NOR4_X1 U9314 ( .A1(n7766), .A2(n7733), .A3(n7732), .A4(n7731), .ZN(n7734)
         );
  NAND4_X1 U9315 ( .A1(n7505), .A2(n8371), .A3(n7735), .A4(n7734), .ZN(n7736)
         );
  NOR4_X1 U9316 ( .A1(n8258), .A2(n8318), .A3(n4715), .A4(n7736), .ZN(n7738)
         );
  NAND4_X1 U9317 ( .A1(n4730), .A2(n7738), .A3(n8275), .A4(n7737), .ZN(n7739)
         );
  NOR4_X1 U9318 ( .A1(n7788), .A2(n7739), .A3(n8190), .A4(n8207), .ZN(n7740)
         );
  NAND3_X1 U9319 ( .A1(n7742), .A2(n7741), .A3(n7740), .ZN(n7743) );
  XNOR2_X1 U9320 ( .A(n7743), .B(n8253), .ZN(n7748) );
  AOI21_X1 U9321 ( .B1(n7745), .B2(n5740), .A(n7744), .ZN(n7746) );
  AOI21_X1 U9322 ( .B1(n7748), .B2(n7747), .A(n7746), .ZN(n7749) );
  AOI21_X1 U9323 ( .B1(n7751), .B2(n7750), .A(n7749), .ZN(n7752) );
  AOI21_X1 U9324 ( .B1(n7754), .B2(n7753), .A(n7752), .ZN(n7761) );
  NOR4_X1 U9325 ( .A1(n9763), .A2(n7756), .A3(n7755), .A4(n8328), .ZN(n7759)
         );
  OAI21_X1 U9326 ( .B1(n7760), .B2(n7757), .A(P2_B_REG_SCAN_IN), .ZN(n7758) );
  OAI22_X1 U9327 ( .A1(n7761), .A2(n7760), .B1(n7759), .B2(n7758), .ZN(
        P2_U3244) );
  INV_X1 U9328 ( .A(n7762), .ZN(n8381) );
  NAND2_X1 U9329 ( .A1(n7763), .A2(n8381), .ZN(n7764) );
  NAND2_X1 U9330 ( .A1(n7765), .A2(n7764), .ZN(n8387) );
  INV_X1 U9331 ( .A(n8387), .ZN(n7767) );
  NAND2_X1 U9332 ( .A1(n7767), .A2(n7766), .ZN(n8385) );
  INV_X1 U9333 ( .A(n8105), .ZN(n8373) );
  OR2_X1 U9334 ( .A1(n8493), .A2(n8373), .ZN(n7768) );
  INV_X1 U9335 ( .A(n8074), .ZN(n8382) );
  NOR2_X1 U9336 ( .A1(n8487), .A2(n8382), .ZN(n7769) );
  INV_X1 U9337 ( .A(n8487), .ZN(n8369) );
  INV_X1 U9338 ( .A(n8329), .ZN(n8374) );
  NAND2_X1 U9339 ( .A1(n8477), .A2(n8359), .ZN(n7770) );
  NAND2_X1 U9340 ( .A1(n8337), .A2(n7770), .ZN(n8312) );
  INV_X1 U9341 ( .A(n8331), .ZN(n8305) );
  OR2_X1 U9342 ( .A1(n8471), .A2(n8305), .ZN(n7771) );
  NAND2_X1 U9343 ( .A1(n8312), .A2(n7771), .ZN(n7773) );
  NAND2_X1 U9344 ( .A1(n8471), .A2(n8305), .ZN(n7772) );
  NAND2_X1 U9345 ( .A1(n8243), .A2(n8247), .ZN(n8244) );
  NAND2_X1 U9346 ( .A1(n7507), .A2(n7777), .ZN(n7778) );
  NAND2_X1 U9347 ( .A1(n8206), .A2(n7778), .ZN(n8191) );
  NAND2_X1 U9348 ( .A1(n8191), .A2(n8190), .ZN(n8189) );
  INV_X1 U9349 ( .A(n7779), .ZN(n8217) );
  NAND2_X1 U9350 ( .A1(n8189), .A2(n7781), .ZN(n7783) );
  XNOR2_X2 U9351 ( .A(n7783), .B(n7782), .ZN(n8434) );
  INV_X1 U9352 ( .A(n8477), .ZN(n8344) );
  INV_X1 U9353 ( .A(n8483), .ZN(n8353) );
  NAND2_X1 U9354 ( .A1(n8240), .A2(n8251), .ZN(n8233) );
  INV_X1 U9355 ( .A(n8193), .ZN(n7784) );
  AOI22_X1 U9356 ( .A1(n7785), .A2(n8408), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8402), .ZN(n7786) );
  OAI21_X1 U9357 ( .B1(n7787), .B2(n8368), .A(n7786), .ZN(n7796) );
  XNOR2_X1 U9358 ( .A(n7789), .B(n7788), .ZN(n7790) );
  AOI21_X1 U9359 ( .B1(n7791), .B2(P2_B_REG_SCAN_IN), .A(n8330), .ZN(n8181) );
  OAI21_X1 U9360 ( .B1(n8434), .B2(n8399), .A(n7797), .ZN(P2_U3267) );
  NAND2_X1 U9361 ( .A1(n9299), .A2(n7995), .ZN(n7802) );
  NAND2_X1 U9362 ( .A1(n4265), .A2(n9223), .ZN(n7801) );
  NAND2_X1 U9363 ( .A1(n7802), .A2(n7801), .ZN(n7803) );
  XNOR2_X1 U9364 ( .A(n7803), .B(n8009), .ZN(n7806) );
  NOR2_X1 U9365 ( .A1(n8012), .A2(n9002), .ZN(n7804) );
  AOI21_X1 U9366 ( .B1(n9299), .B2(n4265), .A(n7804), .ZN(n7805) );
  XNOR2_X1 U9367 ( .A(n7806), .B(n7805), .ZN(n8602) );
  NAND2_X1 U9368 ( .A1(n7806), .A2(n7805), .ZN(n7807) );
  NAND2_X1 U9369 ( .A1(n7808), .A2(n6363), .ZN(n7810) );
  AOI22_X1 U9370 ( .A1(n7823), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7822), .B2(
        n9571), .ZN(n7809) );
  NAND2_X1 U9371 ( .A1(n9292), .A2(n7995), .ZN(n7812) );
  INV_X1 U9372 ( .A(n8718), .ZN(n9205) );
  NAND2_X1 U9373 ( .A1(n9205), .A2(n4265), .ZN(n7811) );
  NAND2_X1 U9374 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  XNOR2_X1 U9375 ( .A(n7813), .B(n8009), .ZN(n7817) );
  NAND2_X1 U9376 ( .A1(n9292), .A2(n4265), .ZN(n7815) );
  NAND2_X1 U9377 ( .A1(n7974), .A2(n9205), .ZN(n7814) );
  NAND2_X1 U9378 ( .A1(n7815), .A2(n7814), .ZN(n8642) );
  INV_X1 U9379 ( .A(n7817), .ZN(n7818) );
  NAND2_X1 U9381 ( .A1(n7821), .A2(n6363), .ZN(n7825) );
  AOI22_X1 U9382 ( .A1(n7823), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9588), .B2(
        n7822), .ZN(n7824) );
  NAND2_X1 U9383 ( .A1(n9288), .A2(n7995), .ZN(n7835) );
  INV_X1 U9384 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7833) );
  INV_X1 U9385 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U9386 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  NAND2_X1 U9387 ( .A1(n7848), .A2(n7830), .ZN(n9197) );
  OR2_X1 U9388 ( .A1(n9197), .A2(n8020), .ZN(n7832) );
  AOI22_X1 U9389 ( .A1(n7983), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n8735), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n7831) );
  OAI211_X1 U9390 ( .C1(n5691), .C2(n7833), .A(n7832), .B(n7831), .ZN(n9222)
         );
  NAND2_X1 U9391 ( .A1(n9222), .A2(n4265), .ZN(n7834) );
  NAND2_X1 U9392 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  XNOR2_X1 U9393 ( .A(n7836), .B(n7989), .ZN(n7840) );
  NAND2_X1 U9394 ( .A1(n9288), .A2(n4265), .ZN(n7838) );
  NAND2_X1 U9395 ( .A1(n7974), .A2(n9222), .ZN(n7837) );
  NAND2_X1 U9396 ( .A1(n7838), .A2(n7837), .ZN(n7841) );
  INV_X1 U9397 ( .A(n8569), .ZN(n7839) );
  INV_X1 U9398 ( .A(n7840), .ZN(n7843) );
  INV_X1 U9399 ( .A(n7841), .ZN(n7842) );
  NAND2_X1 U9400 ( .A1(n7843), .A2(n7842), .ZN(n8567) );
  NAND2_X1 U9401 ( .A1(n7844), .A2(n6363), .ZN(n7847) );
  OR2_X1 U9402 ( .A1(n8732), .A2(n7845), .ZN(n7846) );
  NAND2_X1 U9403 ( .A1(n9284), .A2(n7995), .ZN(n7857) );
  INV_X1 U9404 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U9405 ( .A1(n7848), .A2(n8621), .ZN(n7849) );
  NAND2_X1 U9406 ( .A1(n7869), .A2(n7849), .ZN(n9187) );
  OR2_X1 U9407 ( .A1(n9187), .A2(n8020), .ZN(n7855) );
  INV_X1 U9408 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n7852) );
  NAND2_X1 U9409 ( .A1(n7826), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7851) );
  NAND2_X1 U9410 ( .A1(n8735), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7850) );
  OAI211_X1 U9411 ( .C1(n8024), .C2(n7852), .A(n7851), .B(n7850), .ZN(n7853)
         );
  INV_X1 U9412 ( .A(n7853), .ZN(n7854) );
  NAND2_X1 U9413 ( .A1(n7855), .A2(n7854), .ZN(n9204) );
  NAND2_X1 U9414 ( .A1(n9204), .A2(n4265), .ZN(n7856) );
  NAND2_X1 U9415 ( .A1(n7857), .A2(n7856), .ZN(n7858) );
  XNOR2_X1 U9416 ( .A(n7858), .B(n7989), .ZN(n7860) );
  AND2_X1 U9417 ( .A1(n9204), .A2(n7974), .ZN(n7859) );
  AOI21_X1 U9418 ( .B1(n9284), .B2(n4265), .A(n7859), .ZN(n7861) );
  XNOR2_X1 U9419 ( .A(n7860), .B(n7861), .ZN(n8619) );
  INV_X1 U9420 ( .A(n7860), .ZN(n7862) );
  NAND2_X1 U9421 ( .A1(n7862), .A2(n7861), .ZN(n7863) );
  NAND2_X1 U9422 ( .A1(n7864), .A2(n6363), .ZN(n7867) );
  OR2_X1 U9423 ( .A1(n8732), .A2(n7865), .ZN(n7866) );
  NAND2_X1 U9424 ( .A1(n9277), .A2(n7995), .ZN(n7878) );
  INV_X1 U9425 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U9426 ( .A1(n7869), .A2(n7868), .ZN(n7870) );
  AND2_X1 U9427 ( .A1(n7891), .A2(n7870), .ZN(n9174) );
  NAND2_X1 U9428 ( .A1(n9174), .A2(n5712), .ZN(n7876) );
  INV_X1 U9429 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n7873) );
  NAND2_X1 U9430 ( .A1(n7826), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U9431 ( .A1(n8735), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n7871) );
  OAI211_X1 U9432 ( .C1(n8024), .C2(n7873), .A(n7872), .B(n7871), .ZN(n7874)
         );
  INV_X1 U9433 ( .A(n7874), .ZN(n7875) );
  INV_X1 U9434 ( .A(n9184), .ZN(n9161) );
  NAND2_X1 U9435 ( .A1(n9161), .A2(n4265), .ZN(n7877) );
  NAND2_X1 U9436 ( .A1(n7878), .A2(n7877), .ZN(n7879) );
  XNOR2_X1 U9437 ( .A(n7879), .B(n7989), .ZN(n7881) );
  NOR2_X1 U9438 ( .A1(n9184), .A2(n8012), .ZN(n7880) );
  AOI21_X1 U9439 ( .B1(n9277), .B2(n4265), .A(n7880), .ZN(n7882) );
  XNOR2_X1 U9440 ( .A(n7881), .B(n7882), .ZN(n8585) );
  INV_X1 U9441 ( .A(n7881), .ZN(n7883) );
  NAND2_X1 U9442 ( .A1(n7883), .A2(n7882), .ZN(n7884) );
  NAND2_X1 U9443 ( .A1(n7885), .A2(n7884), .ZN(n7902) );
  NAND2_X1 U9444 ( .A1(n7886), .A2(n6363), .ZN(n7888) );
  OR2_X1 U9445 ( .A1(n8732), .A2(n8039), .ZN(n7887) );
  OR2_X1 U9446 ( .A1(n9157), .A2(n6180), .ZN(n7899) );
  INV_X1 U9447 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U9448 ( .A1(n7891), .A2(n7890), .ZN(n7892) );
  NAND2_X1 U9449 ( .A1(n7912), .A2(n7892), .ZN(n9154) );
  OR2_X1 U9450 ( .A1(n9154), .A2(n8020), .ZN(n7897) );
  INV_X1 U9451 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U9452 ( .A1(n7983), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U9453 ( .A1(n4275), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n7893) );
  OAI211_X1 U9454 ( .C1(n9951), .C2(n5690), .A(n7894), .B(n7893), .ZN(n7895)
         );
  INV_X1 U9455 ( .A(n7895), .ZN(n7896) );
  INV_X1 U9456 ( .A(n9141), .ZN(n9167) );
  NAND2_X1 U9457 ( .A1(n9167), .A2(n7974), .ZN(n7898) );
  NAND2_X1 U9458 ( .A1(n7902), .A2(n7903), .ZN(n8626) );
  OAI22_X1 U9459 ( .A1(n9157), .A2(n7900), .B1(n9141), .B2(n6180), .ZN(n7901)
         );
  XNOR2_X1 U9460 ( .A(n7901), .B(n7989), .ZN(n8630) );
  INV_X1 U9461 ( .A(n7902), .ZN(n7905) );
  INV_X1 U9462 ( .A(n7903), .ZN(n7904) );
  AND2_X2 U9463 ( .A1(n7905), .A2(n7904), .ZN(n8631) );
  NAND2_X1 U9464 ( .A1(n7906), .A2(n6363), .ZN(n7909) );
  OR2_X1 U9465 ( .A1(n8732), .A2(n7907), .ZN(n7908) );
  NAND2_X1 U9466 ( .A1(n9267), .A2(n7995), .ZN(n7921) );
  INV_X1 U9467 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U9468 ( .A1(n7912), .A2(n7911), .ZN(n7913) );
  NAND2_X1 U9469 ( .A1(n7928), .A2(n7913), .ZN(n9145) );
  OR2_X1 U9470 ( .A1(n9145), .A2(n8020), .ZN(n7919) );
  INV_X1 U9471 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U9472 ( .A1(n7826), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U9473 ( .A1(n8735), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n7914) );
  OAI211_X1 U9474 ( .C1(n8024), .C2(n7916), .A(n7915), .B(n7914), .ZN(n7917)
         );
  INV_X1 U9475 ( .A(n7917), .ZN(n7918) );
  NAND2_X1 U9476 ( .A1(n7919), .A2(n7918), .ZN(n9160) );
  NAND2_X1 U9477 ( .A1(n9160), .A2(n4265), .ZN(n7920) );
  NAND2_X1 U9478 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  XNOR2_X1 U9479 ( .A(n7922), .B(n7989), .ZN(n7923) );
  AOI22_X1 U9480 ( .A1(n9267), .A2(n4265), .B1(n7974), .B2(n9160), .ZN(n8560)
         );
  NAND2_X1 U9481 ( .A1(n7924), .A2(n6363), .ZN(n7926) );
  OR2_X1 U9482 ( .A1(n8732), .A2(n9920), .ZN(n7925) );
  NAND2_X1 U9483 ( .A1(n9261), .A2(n7995), .ZN(n7935) );
  INV_X1 U9484 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n7927) );
  NAND2_X1 U9485 ( .A1(n7928), .A2(n7927), .ZN(n7929) );
  AND2_X1 U9486 ( .A1(n7944), .A2(n7929), .ZN(n9127) );
  INV_X1 U9487 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7932) );
  NAND2_X1 U9488 ( .A1(n7826), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U9489 ( .A1(n8735), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7930) );
  OAI211_X1 U9490 ( .C1(n8024), .C2(n7932), .A(n7931), .B(n7930), .ZN(n7933)
         );
  AOI21_X1 U9491 ( .B1(n9127), .B2(n5712), .A(n7933), .ZN(n9140) );
  OR2_X1 U9492 ( .A1(n9140), .A2(n6180), .ZN(n7934) );
  NAND2_X1 U9493 ( .A1(n7935), .A2(n7934), .ZN(n7936) );
  XNOR2_X1 U9494 ( .A(n7936), .B(n7989), .ZN(n7938) );
  OAI22_X1 U9495 ( .A1(n9014), .A2(n6180), .B1(n9140), .B2(n8012), .ZN(n7937)
         );
  XNOR2_X1 U9496 ( .A(n7938), .B(n7937), .ZN(n8611) );
  OR2_X1 U9497 ( .A1(n8732), .A2(n9970), .ZN(n7941) );
  INV_X1 U9498 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U9499 ( .A1(n7944), .A2(n8593), .ZN(n7945) );
  NAND2_X1 U9500 ( .A1(n7963), .A2(n7945), .ZN(n9109) );
  INV_X1 U9501 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7948) );
  NAND2_X1 U9502 ( .A1(n8735), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7947) );
  NAND2_X1 U9503 ( .A1(n4275), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n7946) );
  OAI211_X1 U9504 ( .C1(n8024), .C2(n7948), .A(n7947), .B(n7946), .ZN(n7949)
         );
  INV_X1 U9505 ( .A(n7949), .ZN(n7950) );
  OAI22_X1 U9506 ( .A1(n4485), .A2(n6180), .B1(n9017), .B2(n8012), .ZN(n7956)
         );
  NAND2_X1 U9507 ( .A1(n9253), .A2(n7995), .ZN(n7953) );
  NAND2_X1 U9508 ( .A1(n9018), .A2(n4265), .ZN(n7952) );
  NAND2_X1 U9509 ( .A1(n7953), .A2(n7952), .ZN(n7954) );
  XNOR2_X1 U9510 ( .A(n7954), .B(n7989), .ZN(n7955) );
  XOR2_X1 U9511 ( .A(n7956), .B(n7955), .Z(n8592) );
  INV_X1 U9512 ( .A(n7955), .ZN(n7958) );
  INV_X1 U9513 ( .A(n7956), .ZN(n7957) );
  OR2_X1 U9514 ( .A1(n8732), .A2(n7960), .ZN(n7961) );
  NAND2_X1 U9515 ( .A1(n9248), .A2(n7995), .ZN(n7972) );
  INV_X1 U9516 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9925) );
  OR2_X2 U9517 ( .A1(n7963), .A2(n9925), .ZN(n7997) );
  NAND2_X1 U9518 ( .A1(n7963), .A2(n9925), .ZN(n7964) );
  NAND2_X1 U9519 ( .A1(n9096), .A2(n5712), .ZN(n7970) );
  INV_X1 U9520 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U9521 ( .A1(n7826), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7966) );
  NAND2_X1 U9522 ( .A1(n8735), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7965) );
  OAI211_X1 U9523 ( .C1(n8024), .C2(n7967), .A(n7966), .B(n7965), .ZN(n7968)
         );
  INV_X1 U9524 ( .A(n7968), .ZN(n7969) );
  NAND2_X1 U9525 ( .A1(n9114), .A2(n4265), .ZN(n7971) );
  NAND2_X1 U9526 ( .A1(n7972), .A2(n7971), .ZN(n7973) );
  XNOR2_X1 U9527 ( .A(n7973), .B(n7989), .ZN(n7976) );
  AND2_X1 U9528 ( .A1(n9114), .A2(n7974), .ZN(n7975) );
  AOI21_X1 U9529 ( .B1(n9248), .B2(n4265), .A(n7975), .ZN(n7977) );
  XNOR2_X1 U9530 ( .A(n7976), .B(n7977), .ZN(n8654) );
  OR2_X1 U9531 ( .A1(n8732), .A2(n8056), .ZN(n7981) );
  NAND2_X1 U9532 ( .A1(n9245), .A2(n7995), .ZN(n7988) );
  XNOR2_X1 U9533 ( .A(n7997), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9088) );
  INV_X1 U9534 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9978) );
  NAND2_X1 U9535 ( .A1(n7983), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7985) );
  NAND2_X1 U9536 ( .A1(n7826), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7984) );
  OAI211_X1 U9537 ( .C1(n9978), .C2(n5690), .A(n7985), .B(n7984), .ZN(n7986)
         );
  AOI21_X1 U9538 ( .B1(n9088), .B2(n5712), .A(n7986), .ZN(n9075) );
  OR2_X1 U9539 ( .A1(n9075), .A2(n6180), .ZN(n7987) );
  NAND2_X1 U9540 ( .A1(n7988), .A2(n7987), .ZN(n7990) );
  XNOR2_X1 U9541 ( .A(n7990), .B(n7989), .ZN(n8549) );
  NOR2_X1 U9542 ( .A1(n9075), .A2(n8012), .ZN(n7991) );
  AOI21_X1 U9543 ( .B1(n9245), .B2(n4265), .A(n7991), .ZN(n8548) );
  INV_X1 U9544 ( .A(n8548), .ZN(n8016) );
  OR2_X1 U9545 ( .A1(n8732), .A2(n9327), .ZN(n7993) );
  NAND2_X1 U9546 ( .A1(n9238), .A2(n7995), .ZN(n8008) );
  INV_X1 U9547 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8552) );
  INV_X1 U9548 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7996) );
  OAI21_X1 U9549 ( .B1(n7997), .B2(n8552), .A(n7996), .ZN(n8000) );
  INV_X1 U9550 ( .A(n7997), .ZN(n7999) );
  AND2_X1 U9551 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n7998) );
  NAND2_X1 U9552 ( .A1(n7999), .A2(n7998), .ZN(n9057) );
  NAND2_X1 U9553 ( .A1(n8000), .A2(n9057), .ZN(n9070) );
  OR2_X1 U9554 ( .A1(n9070), .A2(n8020), .ZN(n8006) );
  INV_X1 U9555 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U9556 ( .A1(n4275), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8002) );
  NAND2_X1 U9557 ( .A1(n8735), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8001) );
  OAI211_X1 U9558 ( .C1(n8024), .C2(n8003), .A(n8002), .B(n8001), .ZN(n8004)
         );
  INV_X1 U9559 ( .A(n8004), .ZN(n8005) );
  INV_X1 U9560 ( .A(n9084), .ZN(n8941) );
  NAND2_X1 U9561 ( .A1(n8941), .A2(n4265), .ZN(n8007) );
  NAND2_X1 U9562 ( .A1(n8008), .A2(n8007), .ZN(n8010) );
  XNOR2_X1 U9563 ( .A(n8010), .B(n8009), .ZN(n8014) );
  NAND2_X1 U9564 ( .A1(n9238), .A2(n4265), .ZN(n8011) );
  OAI21_X1 U9565 ( .B1(n9084), .B2(n8012), .A(n8011), .ZN(n8013) );
  XNOR2_X1 U9566 ( .A(n8014), .B(n8013), .ZN(n8031) );
  INV_X1 U9567 ( .A(n8031), .ZN(n8015) );
  NAND2_X1 U9568 ( .A1(n8015), .A2(n8652), .ZN(n8036) );
  NAND2_X1 U9569 ( .A1(n8549), .A2(n8016), .ZN(n8030) );
  INV_X1 U9570 ( .A(n8030), .ZN(n8017) );
  NOR2_X1 U9571 ( .A1(n8017), .A2(n8650), .ZN(n8018) );
  AND2_X1 U9572 ( .A1(n8031), .A2(n8018), .ZN(n8019) );
  NAND2_X1 U9573 ( .A1(n8037), .A2(n8019), .ZN(n8035) );
  OR2_X1 U9574 ( .A1(n9057), .A2(n8020), .ZN(n8027) );
  INV_X1 U9575 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8023) );
  NAND2_X1 U9576 ( .A1(n7826), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8022) );
  NAND2_X1 U9577 ( .A1(n8735), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8021) );
  OAI211_X1 U9578 ( .C1(n8024), .C2(n8023), .A(n8022), .B(n8021), .ZN(n8025)
         );
  INV_X1 U9579 ( .A(n8025), .ZN(n8026) );
  INV_X1 U9580 ( .A(n9074), .ZN(n8940) );
  AOI22_X1 U9581 ( .A1(n8940), .A2(n8644), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8029) );
  INV_X1 U9582 ( .A(n9075), .ZN(n9101) );
  NAND2_X1 U9583 ( .A1(n9101), .A2(n8633), .ZN(n8028) );
  OAI211_X1 U9584 ( .C1(n8646), .C2(n9070), .A(n8029), .B(n8028), .ZN(n8033)
         );
  NOR3_X1 U9585 ( .A1(n8031), .A2(n8650), .A3(n8030), .ZN(n8032) );
  AOI211_X1 U9586 ( .C1(n9238), .C2(n8648), .A(n8033), .B(n8032), .ZN(n8034)
         );
  OAI211_X1 U9587 ( .C1(n8037), .C2(n8036), .A(n8035), .B(n8034), .ZN(P1_U3218) );
  OAI222_X1 U9588 ( .A1(n9328), .A2(n8039), .B1(n8059), .B2(n8038), .C1(n8886), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  NAND2_X1 U9589 ( .A1(n8217), .A2(n8041), .ZN(n8042) );
  XOR2_X1 U9590 ( .A(n8043), .B(n8042), .Z(n8044) );
  XNOR2_X1 U9591 ( .A(n8435), .B(n8044), .ZN(n8045) );
  XNOR2_X1 U9592 ( .A(n8046), .B(n8045), .ZN(n8053) );
  INV_X1 U9593 ( .A(n8047), .ZN(n8194) );
  AOI22_X1 U9594 ( .A1(n8194), .A2(n8140), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8049) );
  NAND2_X1 U9595 ( .A1(n8200), .A2(n9717), .ZN(n8048) );
  OAI211_X1 U9596 ( .C1(n8050), .C2(n9714), .A(n8049), .B(n8048), .ZN(n8051)
         );
  AOI21_X1 U9597 ( .B1(n8435), .B2(n8147), .A(n8051), .ZN(n8052) );
  OAI21_X1 U9598 ( .B1(n8053), .B2(n8128), .A(n8052), .ZN(P2_U3222) );
  OAI222_X1 U9599 ( .A1(n9328), .A2(n8056), .B1(P1_U3084), .B2(n8055), .C1(
        n8054), .C2(n8059), .ZN(P1_U3326) );
  INV_X1 U9600 ( .A(n8664), .ZN(n9320) );
  OAI222_X1 U9601 ( .A1(n8057), .A2(P2_U3152), .B1(n4270), .B2(n9320), .C1(
        n9896), .C2(n8545), .ZN(P2_U3329) );
  INV_X1 U9602 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8731) );
  INV_X1 U9603 ( .A(n8730), .ZN(n8061) );
  OAI222_X1 U9604 ( .A1(n9328), .A2(n8731), .B1(n8059), .B2(n8061), .C1(
        P1_U3084), .C2(n8058), .ZN(P1_U3323) );
  OAI222_X1 U9605 ( .A1(P2_U3152), .A2(n4988), .B1(n4270), .B2(n8061), .C1(
        n8060), .C2(n8545), .ZN(P2_U3328) );
  XNOR2_X1 U9606 ( .A(n8063), .B(n8114), .ZN(n8069) );
  INV_X1 U9607 ( .A(n8064), .ZN(n8291) );
  OAI22_X1 U9608 ( .A1(n9737), .A2(n8291), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8065), .ZN(n8067) );
  OAI22_X1 U9609 ( .A1(n8135), .A2(n8283), .B1(n8284), .B2(n9714), .ZN(n8066)
         );
  AOI211_X1 U9610 ( .C1(n8293), .C2(n8147), .A(n8067), .B(n8066), .ZN(n8068)
         );
  OAI21_X1 U9611 ( .B1(n8069), .B2(n8128), .A(n8068), .ZN(P2_U3218) );
  INV_X1 U9612 ( .A(n8071), .ZN(n8072) );
  AOI21_X1 U9613 ( .B1(n8070), .B2(n8073), .A(n8072), .ZN(n8078) );
  AND2_X1 U9614 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8177) );
  OAI22_X1 U9615 ( .A1(n8135), .A2(n8074), .B1(n8085), .B2(n9714), .ZN(n8075)
         );
  AOI211_X1 U9616 ( .C1(n8140), .C2(n8351), .A(n8177), .B(n8075), .ZN(n8077)
         );
  NAND2_X1 U9617 ( .A1(n8483), .A2(n8147), .ZN(n8076) );
  OAI211_X1 U9618 ( .C1(n8078), .C2(n8128), .A(n8077), .B(n8076), .ZN(P2_U3221) );
  OR2_X1 U9619 ( .A1(n8079), .A2(n8124), .ZN(n8081) );
  NAND2_X1 U9620 ( .A1(n8081), .A2(n8080), .ZN(n8083) );
  XNOR2_X1 U9621 ( .A(n8083), .B(n8082), .ZN(n8089) );
  INV_X1 U9622 ( .A(n8321), .ZN(n8084) );
  OAI22_X1 U9623 ( .A1(n9737), .A2(n8084), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9905), .ZN(n8087) );
  OAI22_X1 U9624 ( .A1(n8135), .A2(n8085), .B1(n8283), .B2(n9714), .ZN(n8086)
         );
  AOI211_X1 U9625 ( .C1(n8471), .C2(n8147), .A(n8087), .B(n8086), .ZN(n8088)
         );
  OAI21_X1 U9626 ( .B1(n8089), .B2(n8128), .A(n8088), .ZN(P2_U3225) );
  XNOR2_X1 U9627 ( .A(n8091), .B(n8090), .ZN(n8092) );
  XNOR2_X1 U9628 ( .A(n10043), .B(n8092), .ZN(n8099) );
  NOR2_X1 U9629 ( .A1(n8284), .A2(n8328), .ZN(n8094) );
  AOI21_X1 U9630 ( .B1(n8216), .B2(n8417), .A(n8094), .ZN(n8249) );
  NOR2_X1 U9631 ( .A1(n8249), .A2(n8142), .ZN(n8097) );
  OAI22_X1 U9632 ( .A1(n8252), .A2(n9737), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8095), .ZN(n8096) );
  AOI211_X1 U9633 ( .C1(n8451), .C2(n8147), .A(n8097), .B(n8096), .ZN(n8098)
         );
  OAI21_X1 U9634 ( .B1(n8099), .B2(n8128), .A(n8098), .ZN(P2_U3227) );
  INV_X1 U9635 ( .A(n8100), .ZN(n8102) );
  NOR3_X1 U9636 ( .A1(n8103), .A2(n8102), .A3(n8101), .ZN(n8104) );
  OAI21_X1 U9637 ( .B1(n8104), .B2(n4344), .A(n9733), .ZN(n8111) );
  OAI22_X1 U9638 ( .A1(n8135), .A2(n8106), .B1(n8105), .B2(n9714), .ZN(n8107)
         );
  AOI211_X1 U9639 ( .C1(n8140), .C2(n8109), .A(n8108), .B(n8107), .ZN(n8110)
         );
  OAI211_X1 U9640 ( .C1(n8497), .C2(n9731), .A(n8111), .B(n8110), .ZN(P2_U3228) );
  INV_X1 U9641 ( .A(n8112), .ZN(n8113) );
  OAI21_X1 U9642 ( .B1(n8063), .B2(n8114), .A(n8113), .ZN(n8118) );
  XNOR2_X1 U9643 ( .A(n8116), .B(n8115), .ZN(n8117) );
  XNOR2_X1 U9644 ( .A(n8118), .B(n8117), .ZN(n8123) );
  OAI22_X1 U9645 ( .A1(n9737), .A2(n8262), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9910), .ZN(n8121) );
  OAI22_X1 U9646 ( .A1(n8119), .A2(n9714), .B1(n8135), .B2(n8134), .ZN(n8120)
         );
  AOI211_X1 U9647 ( .C1(n8454), .C2(n8147), .A(n8121), .B(n8120), .ZN(n8122)
         );
  OAI21_X1 U9648 ( .B1(n8123), .B2(n8128), .A(n8122), .ZN(P2_U3231) );
  XNOR2_X1 U9649 ( .A(n8079), .B(n8124), .ZN(n8129) );
  OAI22_X1 U9650 ( .A1(n9737), .A2(n8341), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9967), .ZN(n8126) );
  OAI22_X1 U9651 ( .A1(n8135), .A2(n8329), .B1(n8331), .B2(n9714), .ZN(n8125)
         );
  AOI211_X1 U9652 ( .C1(n8477), .C2(n8147), .A(n8126), .B(n8125), .ZN(n8127)
         );
  OAI21_X1 U9653 ( .B1(n8129), .B2(n8128), .A(n8127), .ZN(P2_U3235) );
  OAI21_X1 U9654 ( .B1(n8132), .B2(n8131), .A(n8130), .ZN(n8133) );
  NAND2_X1 U9655 ( .A1(n8133), .A2(n9733), .ZN(n8139) );
  NOR2_X1 U9656 ( .A1(n9737), .A2(n8299), .ZN(n8137) );
  OAI22_X1 U9657 ( .A1(n8135), .A2(n8331), .B1(n8134), .B2(n9714), .ZN(n8136)
         );
  AOI211_X1 U9658 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n8137), 
        .B(n8136), .ZN(n8138) );
  OAI211_X1 U9659 ( .C1(n4552), .C2(n9731), .A(n8139), .B(n8138), .ZN(P2_U3237) );
  AOI22_X1 U9660 ( .A1(n8200), .A2(n8417), .B1(n8419), .B2(n8269), .ZN(n8231)
         );
  AOI22_X1 U9661 ( .A1(n8237), .A2(n8140), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8141) );
  OAI21_X1 U9662 ( .B1(n8231), .B2(n8142), .A(n8141), .ZN(n8146) );
  MUX2_X1 U9663 ( .A(n8148), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8160), .Z(
        P2_U3582) );
  MUX2_X1 U9664 ( .A(n8199), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8160), .Z(
        P2_U3581) );
  MUX2_X1 U9665 ( .A(n8217), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8160), .Z(
        P2_U3580) );
  MUX2_X1 U9666 ( .A(n8200), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8160), .Z(
        P2_U3579) );
  MUX2_X1 U9667 ( .A(n8216), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8160), .Z(
        P2_U3578) );
  MUX2_X1 U9668 ( .A(n8269), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8160), .Z(
        P2_U3577) );
  MUX2_X1 U9669 ( .A(n7414), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8160), .Z(
        P2_U3576) );
  MUX2_X1 U9670 ( .A(n8306), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8160), .Z(
        P2_U3575) );
  MUX2_X1 U9671 ( .A(n8319), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8160), .Z(
        P2_U3574) );
  MUX2_X1 U9672 ( .A(n8305), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8160), .Z(
        P2_U3573) );
  MUX2_X1 U9673 ( .A(n8359), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8160), .Z(
        P2_U3572) );
  MUX2_X1 U9674 ( .A(n8374), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8160), .Z(
        P2_U3571) );
  MUX2_X1 U9675 ( .A(n8382), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8160), .Z(
        P2_U3570) );
  MUX2_X1 U9676 ( .A(n8373), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8160), .Z(
        P2_U3569) );
  MUX2_X1 U9677 ( .A(n8381), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8160), .Z(
        P2_U3568) );
  MUX2_X1 U9678 ( .A(n8149), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8160), .Z(
        P2_U3567) );
  MUX2_X1 U9679 ( .A(n8150), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8160), .Z(
        P2_U3566) );
  MUX2_X1 U9680 ( .A(n8151), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8160), .Z(
        P2_U3565) );
  MUX2_X1 U9681 ( .A(n8152), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8160), .Z(
        P2_U3564) );
  MUX2_X1 U9682 ( .A(n8153), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8160), .Z(
        P2_U3563) );
  MUX2_X1 U9683 ( .A(n8154), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8160), .Z(
        P2_U3562) );
  MUX2_X1 U9684 ( .A(n9704), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8160), .Z(
        P2_U3561) );
  MUX2_X1 U9685 ( .A(n8155), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8160), .Z(
        P2_U3560) );
  MUX2_X1 U9686 ( .A(n9716), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8160), .Z(
        P2_U3559) );
  MUX2_X1 U9687 ( .A(n8156), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8160), .Z(
        P2_U3558) );
  MUX2_X1 U9688 ( .A(n8157), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8160), .Z(
        P2_U3557) );
  MUX2_X1 U9689 ( .A(n8158), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8160), .Z(
        P2_U3556) );
  MUX2_X1 U9690 ( .A(n8159), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8160), .Z(
        P2_U3555) );
  MUX2_X1 U9691 ( .A(n8418), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8160), .Z(
        P2_U3554) );
  MUX2_X1 U9692 ( .A(n5593), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8160), .Z(
        P2_U3553) );
  MUX2_X1 U9693 ( .A(n5110), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8160), .Z(
        P2_U3552) );
  NAND2_X1 U9694 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  NAND2_X1 U9695 ( .A1(n8164), .A2(n8163), .ZN(n8165) );
  XNOR2_X1 U9696 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8165), .ZN(n8172) );
  NAND2_X1 U9697 ( .A1(n8167), .A2(n8166), .ZN(n8169) );
  INV_X1 U9698 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8168) );
  XNOR2_X1 U9699 ( .A(n8169), .B(n8168), .ZN(n8174) );
  INV_X1 U9700 ( .A(n8174), .ZN(n8170) );
  AOI22_X1 U9701 ( .A1(n8172), .A2(n9749), .B1(n9753), .B2(n8170), .ZN(n8176)
         );
  NOR2_X1 U9702 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  AOI211_X1 U9703 ( .C1(n9753), .C2(n8174), .A(n9757), .B(n8173), .ZN(n8175)
         );
  MUX2_X1 U9704 ( .A(n8176), .B(n8175), .S(n8253), .Z(n8179) );
  AOI21_X1 U9705 ( .B1(n9747), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n8177), .ZN(
        n8178) );
  NAND2_X1 U9706 ( .A1(n8179), .A2(n8178), .ZN(P2_U3264) );
  NAND2_X1 U9707 ( .A1(n9343), .A2(n8184), .ZN(n8180) );
  XNOR2_X1 U9708 ( .A(n8427), .B(n8180), .ZN(n8429) );
  NAND2_X1 U9709 ( .A1(n8181), .A2(n7543), .ZN(n9342) );
  NOR2_X1 U9710 ( .A1(n8402), .A2(n9342), .ZN(n8186) );
  AOI21_X1 U9711 ( .B1(n8402), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8186), .ZN(
        n8183) );
  NAND2_X1 U9712 ( .A1(n8427), .A2(n8406), .ZN(n8182) );
  OAI211_X1 U9713 ( .C1(n8429), .C2(n8295), .A(n8183), .B(n8182), .ZN(P2_U3265) );
  XNOR2_X1 U9714 ( .A(n8185), .B(n8184), .ZN(n9345) );
  NAND2_X1 U9715 ( .A1(n9345), .A2(n8409), .ZN(n8188) );
  AOI21_X1 U9716 ( .B1(n8402), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8186), .ZN(
        n8187) );
  OAI211_X1 U9717 ( .C1(n9343), .C2(n8368), .A(n8188), .B(n8187), .ZN(P2_U3266) );
  OAI21_X1 U9718 ( .B1(n8191), .B2(n8190), .A(n8189), .ZN(n8192) );
  INV_X1 U9719 ( .A(n8192), .ZN(n8439) );
  AOI21_X1 U9720 ( .B1(n8435), .B2(n8210), .A(n8193), .ZN(n8436) );
  AOI22_X1 U9721 ( .A1(n8194), .A2(n8408), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8402), .ZN(n8195) );
  OAI21_X1 U9722 ( .B1(n7780), .B2(n8368), .A(n8195), .ZN(n8204) );
  OAI211_X1 U9723 ( .C1(n8198), .C2(n8197), .A(n8196), .B(n8414), .ZN(n8202)
         );
  AOI22_X1 U9724 ( .A1(n8200), .A2(n8419), .B1(n8199), .B2(n8417), .ZN(n8201)
         );
  NOR2_X1 U9725 ( .A1(n8438), .A2(n8402), .ZN(n8203) );
  AOI211_X1 U9726 ( .C1(n8436), .C2(n8409), .A(n8204), .B(n8203), .ZN(n8205)
         );
  OAI21_X1 U9727 ( .B1(n8439), .B2(n8399), .A(n8205), .ZN(P2_U3268) );
  OAI21_X1 U9728 ( .B1(n8208), .B2(n8207), .A(n8206), .ZN(n8209) );
  INV_X1 U9729 ( .A(n8209), .ZN(n8444) );
  AOI21_X1 U9730 ( .B1(n8440), .B2(n8233), .A(n4548), .ZN(n8441) );
  AOI22_X1 U9731 ( .A1(n8211), .A2(n8408), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8402), .ZN(n8212) );
  OAI21_X1 U9732 ( .B1(n7507), .B2(n8368), .A(n8212), .ZN(n8221) );
  OAI211_X1 U9733 ( .C1(n8215), .C2(n8214), .A(n8213), .B(n8414), .ZN(n8219)
         );
  AOI22_X1 U9734 ( .A1(n8217), .A2(n8417), .B1(n8419), .B2(n8216), .ZN(n8218)
         );
  NOR2_X1 U9735 ( .A1(n8443), .A2(n8402), .ZN(n8220) );
  AOI211_X1 U9736 ( .C1(n8441), .C2(n8409), .A(n8221), .B(n8220), .ZN(n8222)
         );
  OAI21_X1 U9737 ( .B1(n8444), .B2(n8399), .A(n8222), .ZN(P2_U3269) );
  OAI21_X1 U9738 ( .B1(n8224), .B2(n8230), .A(n8223), .ZN(n8225) );
  INV_X1 U9739 ( .A(n8225), .ZN(n8448) );
  OR2_X1 U9740 ( .A1(n8226), .A2(n8227), .ZN(n8229) );
  AOI21_X1 U9741 ( .B1(n8230), .B2(n8229), .A(n8228), .ZN(n8232) );
  INV_X1 U9742 ( .A(n8251), .ZN(n8235) );
  INV_X1 U9743 ( .A(n8233), .ZN(n8234) );
  AOI211_X1 U9744 ( .C1(n8447), .C2(n8235), .A(n9781), .B(n8234), .ZN(n8446)
         );
  AND2_X1 U9745 ( .A1(n8422), .A2(n8236), .ZN(n8396) );
  NAND2_X1 U9746 ( .A1(n8446), .A2(n8396), .ZN(n8239) );
  AOI22_X1 U9747 ( .A1(n8237), .A2(n8408), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n8402), .ZN(n8238) );
  OAI211_X1 U9748 ( .C1(n8240), .C2(n8368), .A(n8239), .B(n8238), .ZN(n8241)
         );
  AOI21_X1 U9749 ( .B1(n8445), .B2(n8422), .A(n8241), .ZN(n8242) );
  OAI21_X1 U9750 ( .B1(n8448), .B2(n8399), .A(n8242), .ZN(P2_U3270) );
  OAI21_X1 U9751 ( .B1(n8243), .B2(n8247), .A(n8244), .ZN(n8245) );
  INV_X1 U9752 ( .A(n8245), .ZN(n8453) );
  AOI22_X1 U9753 ( .A1(n8451), .A2(n8406), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8402), .ZN(n8257) );
  NAND3_X1 U9754 ( .A1(n8266), .A2(n8247), .A3(n8246), .ZN(n8248) );
  NAND2_X1 U9755 ( .A1(n8248), .A2(n8414), .ZN(n8250) );
  OAI21_X1 U9756 ( .B1(n8226), .B2(n8250), .A(n8249), .ZN(n8449) );
  AOI211_X1 U9757 ( .C1(n8451), .C2(n8260), .A(n9781), .B(n8251), .ZN(n8450)
         );
  INV_X1 U9758 ( .A(n8450), .ZN(n8254) );
  OAI22_X1 U9759 ( .A1(n8254), .A2(n8253), .B1(n8389), .B2(n8252), .ZN(n8255)
         );
  OAI21_X1 U9760 ( .B1(n8449), .B2(n8255), .A(n8422), .ZN(n8256) );
  OAI211_X1 U9761 ( .C1(n8453), .C2(n8399), .A(n8257), .B(n8256), .ZN(P2_U3271) );
  XNOR2_X1 U9762 ( .A(n8259), .B(n8258), .ZN(n8458) );
  INV_X1 U9763 ( .A(n8260), .ZN(n8261) );
  AOI21_X1 U9764 ( .B1(n8454), .B2(n8289), .A(n8261), .ZN(n8455) );
  INV_X1 U9765 ( .A(n8454), .ZN(n8265) );
  INV_X1 U9766 ( .A(n8262), .ZN(n8263) );
  AOI22_X1 U9767 ( .A1(n8263), .A2(n8408), .B1(n8402), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8264) );
  OAI21_X1 U9768 ( .B1(n8265), .B2(n8368), .A(n8264), .ZN(n8273) );
  OAI211_X1 U9769 ( .C1(n8268), .C2(n8267), .A(n8266), .B(n8414), .ZN(n8271)
         );
  AOI22_X1 U9770 ( .A1(n8269), .A2(n8417), .B1(n8419), .B2(n8306), .ZN(n8270)
         );
  NOR2_X1 U9771 ( .A1(n8457), .A2(n8402), .ZN(n8272) );
  AOI211_X1 U9772 ( .C1(n8455), .C2(n8409), .A(n8273), .B(n8272), .ZN(n8274)
         );
  OAI21_X1 U9773 ( .B1(n8399), .B2(n8458), .A(n8274), .ZN(P2_U3272) );
  NAND2_X1 U9774 ( .A1(n8276), .A2(n8275), .ZN(n8277) );
  NAND2_X1 U9775 ( .A1(n8278), .A2(n8277), .ZN(n8459) );
  AND2_X1 U9776 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  OAI21_X1 U9777 ( .B1(n8282), .B2(n8281), .A(n8414), .ZN(n8287) );
  OAI22_X1 U9778 ( .A1(n8284), .A2(n8330), .B1(n8283), .B2(n8328), .ZN(n8285)
         );
  INV_X1 U9779 ( .A(n8285), .ZN(n8286) );
  NAND2_X1 U9780 ( .A1(n8287), .A2(n8286), .ZN(n8463) );
  OR2_X1 U9781 ( .A1(n8460), .A2(n4339), .ZN(n8288) );
  NAND2_X1 U9782 ( .A1(n8289), .A2(n8288), .ZN(n8461) );
  OAI22_X1 U9783 ( .A1(n8291), .A2(n8389), .B1(n8422), .B2(n8290), .ZN(n8292)
         );
  AOI21_X1 U9784 ( .B1(n8293), .B2(n8406), .A(n8292), .ZN(n8294) );
  OAI21_X1 U9785 ( .B1(n8461), .B2(n8295), .A(n8294), .ZN(n8296) );
  AOI21_X1 U9786 ( .B1(n8463), .B2(n8422), .A(n8296), .ZN(n8297) );
  OAI21_X1 U9787 ( .B1(n8459), .B2(n8399), .A(n8297), .ZN(P2_U3273) );
  XNOR2_X1 U9788 ( .A(n8298), .B(n4715), .ZN(n8470) );
  AOI21_X1 U9789 ( .B1(n8466), .B2(n8313), .A(n4339), .ZN(n8467) );
  INV_X1 U9790 ( .A(n8299), .ZN(n8300) );
  AOI22_X1 U9791 ( .A1(n8402), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8300), .B2(
        n8408), .ZN(n8301) );
  OAI21_X1 U9792 ( .B1(n4552), .B2(n8368), .A(n8301), .ZN(n8310) );
  OAI211_X1 U9793 ( .C1(n8304), .C2(n8303), .A(n8302), .B(n8414), .ZN(n8308)
         );
  AOI22_X1 U9794 ( .A1(n8306), .A2(n8417), .B1(n8419), .B2(n8305), .ZN(n8307)
         );
  NOR2_X1 U9795 ( .A1(n8469), .A2(n8402), .ZN(n8309) );
  AOI211_X1 U9796 ( .C1(n8467), .C2(n8409), .A(n8310), .B(n8309), .ZN(n8311)
         );
  OAI21_X1 U9797 ( .B1(n8399), .B2(n8470), .A(n8311), .ZN(P2_U3274) );
  XNOR2_X1 U9798 ( .A(n8312), .B(n8318), .ZN(n8475) );
  INV_X1 U9799 ( .A(n8313), .ZN(n8314) );
  AOI21_X1 U9800 ( .B1(n8471), .B2(n8338), .A(n8314), .ZN(n8472) );
  INV_X1 U9801 ( .A(n8471), .ZN(n8316) );
  OAI22_X1 U9802 ( .A1(n8316), .A2(n8368), .B1(n8422), .B2(n8315), .ZN(n8324)
         );
  XNOR2_X1 U9803 ( .A(n8317), .B(n8318), .ZN(n8320) );
  AOI222_X1 U9804 ( .A1(n8384), .A2(n8320), .B1(n8319), .B2(n8417), .C1(n8359), 
        .C2(n8419), .ZN(n8474) );
  NAND2_X1 U9805 ( .A1(n8408), .A2(n8321), .ZN(n8322) );
  AOI21_X1 U9806 ( .B1(n8474), .B2(n8322), .A(n8402), .ZN(n8323) );
  AOI211_X1 U9807 ( .C1(n8472), .C2(n8409), .A(n8324), .B(n8323), .ZN(n8325)
         );
  OAI21_X1 U9808 ( .B1(n8399), .B2(n8475), .A(n8325), .ZN(P2_U3275) );
  AOI21_X1 U9809 ( .B1(n8327), .B2(n8335), .A(n8326), .ZN(n8334) );
  OAI22_X1 U9810 ( .A1(n8331), .A2(n8330), .B1(n8329), .B2(n8328), .ZN(n8332)
         );
  AOI21_X1 U9811 ( .B1(n8334), .B2(n8333), .A(n8332), .ZN(n8480) );
  OR2_X1 U9812 ( .A1(n8336), .A2(n8335), .ZN(n8476) );
  NAND3_X1 U9813 ( .A1(n8476), .A2(n8407), .A3(n8337), .ZN(n8347) );
  INV_X1 U9814 ( .A(n8349), .ZN(n8340) );
  INV_X1 U9815 ( .A(n8338), .ZN(n8339) );
  AOI21_X1 U9816 ( .B1(n8477), .B2(n8340), .A(n8339), .ZN(n8478) );
  INV_X1 U9817 ( .A(n8341), .ZN(n8342) );
  AOI22_X1 U9818 ( .A1(n8402), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8342), .B2(
        n8408), .ZN(n8343) );
  OAI21_X1 U9819 ( .B1(n8344), .B2(n8368), .A(n8343), .ZN(n8345) );
  AOI21_X1 U9820 ( .B1(n8478), .B2(n8409), .A(n8345), .ZN(n8346) );
  OAI211_X1 U9821 ( .C1(n8402), .C2(n8480), .A(n8347), .B(n8346), .ZN(P2_U3276) );
  XNOR2_X1 U9822 ( .A(n8348), .B(n8354), .ZN(n8486) );
  INV_X1 U9823 ( .A(n8365), .ZN(n8350) );
  AOI211_X1 U9824 ( .C1(n8483), .C2(n8350), .A(n9781), .B(n8349), .ZN(n8482)
         );
  AOI22_X1 U9825 ( .A1(n8402), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8351), .B2(
        n8408), .ZN(n8352) );
  OAI21_X1 U9826 ( .B1(n8353), .B2(n8368), .A(n8352), .ZN(n8362) );
  INV_X1 U9827 ( .A(n8370), .ZN(n8356) );
  OAI21_X1 U9828 ( .B1(n8356), .B2(n8355), .A(n8354), .ZN(n8358) );
  NAND2_X1 U9829 ( .A1(n8358), .A2(n8357), .ZN(n8360) );
  AOI222_X1 U9830 ( .A1(n8384), .A2(n8360), .B1(n8359), .B2(n8417), .C1(n8382), 
        .C2(n8419), .ZN(n8485) );
  NOR2_X1 U9831 ( .A1(n8485), .A2(n8402), .ZN(n8361) );
  AOI211_X1 U9832 ( .C1(n8482), .C2(n8396), .A(n8362), .B(n8361), .ZN(n8363)
         );
  OAI21_X1 U9833 ( .B1(n8399), .B2(n8486), .A(n8363), .ZN(P2_U3277) );
  XNOR2_X1 U9834 ( .A(n8364), .B(n8371), .ZN(n8491) );
  AOI21_X1 U9835 ( .B1(n8487), .B2(n8394), .A(n8365), .ZN(n8488) );
  AOI22_X1 U9836 ( .A1(n8402), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8366), .B2(
        n8408), .ZN(n8367) );
  OAI21_X1 U9837 ( .B1(n8369), .B2(n8368), .A(n8367), .ZN(n8378) );
  OAI211_X1 U9838 ( .C1(n8372), .C2(n8371), .A(n8370), .B(n8414), .ZN(n8376)
         );
  AOI22_X1 U9839 ( .A1(n8374), .A2(n8417), .B1(n8419), .B2(n8373), .ZN(n8375)
         );
  NOR2_X1 U9840 ( .A1(n8490), .A2(n8402), .ZN(n8377) );
  AOI211_X1 U9841 ( .C1(n8488), .C2(n8409), .A(n8378), .B(n8377), .ZN(n8379)
         );
  OAI21_X1 U9842 ( .B1(n8491), .B2(n8399), .A(n8379), .ZN(P2_U3278) );
  XNOR2_X1 U9843 ( .A(n8380), .B(n8388), .ZN(n8383) );
  AOI222_X1 U9844 ( .A1(n8384), .A2(n8383), .B1(n8382), .B2(n8417), .C1(n8381), 
        .C2(n8419), .ZN(n8495) );
  INV_X1 U9845 ( .A(n8385), .ZN(n8386) );
  AOI21_X1 U9846 ( .B1(n8388), .B2(n8387), .A(n8386), .ZN(n8496) );
  INV_X1 U9847 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8391) );
  OAI22_X1 U9848 ( .A1(n8422), .A2(n8391), .B1(n8390), .B2(n8389), .ZN(n8392)
         );
  AOI21_X1 U9849 ( .B1(n8493), .B2(n8406), .A(n8392), .ZN(n8398) );
  AOI21_X1 U9850 ( .B1(n8393), .B2(n8493), .A(n9781), .ZN(n8395) );
  AND2_X1 U9851 ( .A1(n8395), .A2(n8394), .ZN(n8492) );
  NAND2_X1 U9852 ( .A1(n8492), .A2(n8396), .ZN(n8397) );
  OAI211_X1 U9853 ( .C1(n8496), .C2(n8399), .A(n8398), .B(n8397), .ZN(n8400)
         );
  INV_X1 U9854 ( .A(n8400), .ZN(n8401) );
  OAI21_X1 U9855 ( .B1(n8402), .B2(n8495), .A(n8401), .ZN(P2_U3279) );
  OAI21_X1 U9856 ( .B1(n8413), .B2(n8404), .A(n8403), .ZN(n9778) );
  AOI22_X1 U9857 ( .A1(n8407), .A2(n9778), .B1(n8406), .B2(n8405), .ZN(n8426)
         );
  XNOR2_X1 U9858 ( .A(n5108), .B(n9774), .ZN(n9773) );
  AOI22_X1 U9859 ( .A1(n8409), .A2(n9773), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8408), .ZN(n8425) );
  NAND2_X1 U9860 ( .A1(n8402), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8424) );
  INV_X1 U9861 ( .A(n8410), .ZN(n8416) );
  INV_X1 U9862 ( .A(n8411), .ZN(n8412) );
  NAND2_X1 U9863 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  OAI211_X1 U9864 ( .C1(n7572), .C2(n8416), .A(n8415), .B(n8414), .ZN(n8421)
         );
  AOI22_X1 U9865 ( .A1(n8419), .A2(n5110), .B1(n8418), .B2(n8417), .ZN(n8420)
         );
  NAND2_X1 U9866 ( .A1(n8421), .A2(n8420), .ZN(n9776) );
  NAND2_X1 U9867 ( .A1(n8422), .A2(n9776), .ZN(n8423) );
  NAND4_X1 U9868 ( .A1(n8426), .A2(n8425), .A3(n8424), .A4(n8423), .ZN(
        P2_U3295) );
  NAND2_X1 U9869 ( .A1(n8427), .A2(n9809), .ZN(n8428) );
  OAI211_X1 U9870 ( .C1(n8429), .C2(n9781), .A(n9342), .B(n8428), .ZN(n8519)
         );
  MUX2_X1 U9871 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8519), .S(n4268), .Z(
        P2_U3551) );
  AOI22_X1 U9872 ( .A1(n8431), .A2(n9810), .B1(n9809), .B2(n8430), .ZN(n8433)
         );
  OAI21_X1 U9873 ( .B1(n8434), .B2(n9804), .A(n4817), .ZN(n8520) );
  MUX2_X1 U9874 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8520), .S(n4268), .Z(
        P2_U3549) );
  AOI22_X1 U9875 ( .A1(n8436), .A2(n9810), .B1(n9809), .B2(n8435), .ZN(n8437)
         );
  OAI211_X1 U9876 ( .C1(n8439), .C2(n9804), .A(n8438), .B(n8437), .ZN(n8521)
         );
  MUX2_X1 U9877 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8521), .S(n4268), .Z(
        P2_U3548) );
  AOI22_X1 U9878 ( .A1(n8441), .A2(n9810), .B1(n9809), .B2(n8440), .ZN(n8442)
         );
  OAI211_X1 U9879 ( .C1(n8444), .C2(n9804), .A(n8443), .B(n8442), .ZN(n8522)
         );
  MUX2_X1 U9880 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8522), .S(n4268), .Z(
        P2_U3547) );
  MUX2_X1 U9881 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8523), .S(n4268), .Z(
        P2_U3546) );
  AOI211_X1 U9882 ( .C1(n9809), .C2(n8451), .A(n8450), .B(n8449), .ZN(n8452)
         );
  OAI21_X1 U9883 ( .B1(n8453), .B2(n9804), .A(n8452), .ZN(n8524) );
  MUX2_X1 U9884 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8524), .S(n4268), .Z(
        P2_U3545) );
  AOI22_X1 U9885 ( .A1(n8455), .A2(n9810), .B1(n9809), .B2(n8454), .ZN(n8456)
         );
  OAI211_X1 U9886 ( .C1(n8458), .C2(n9804), .A(n8457), .B(n8456), .ZN(n8525)
         );
  MUX2_X1 U9887 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8525), .S(n4268), .Z(
        P2_U3544) );
  OR2_X1 U9888 ( .A1(n8459), .A2(n9804), .ZN(n8465) );
  OAI22_X1 U9889 ( .A1(n8461), .A2(n9781), .B1(n8460), .B2(n9820), .ZN(n8462)
         );
  NOR2_X1 U9890 ( .A1(n8463), .A2(n8462), .ZN(n8464) );
  NAND2_X1 U9891 ( .A1(n8465), .A2(n8464), .ZN(n8526) );
  MUX2_X1 U9892 ( .A(n8526), .B(P2_REG1_REG_23__SCAN_IN), .S(n9833), .Z(
        P2_U3543) );
  AOI22_X1 U9893 ( .A1(n8467), .A2(n9810), .B1(n9809), .B2(n8466), .ZN(n8468)
         );
  OAI211_X1 U9894 ( .C1(n8470), .C2(n9804), .A(n8469), .B(n8468), .ZN(n8527)
         );
  MUX2_X1 U9895 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8527), .S(n4268), .Z(
        P2_U3542) );
  AOI22_X1 U9896 ( .A1(n8472), .A2(n9810), .B1(n9809), .B2(n8471), .ZN(n8473)
         );
  OAI211_X1 U9897 ( .C1(n8475), .C2(n9804), .A(n8474), .B(n8473), .ZN(n8528)
         );
  MUX2_X1 U9898 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8528), .S(n4268), .Z(
        P2_U3541) );
  NAND3_X1 U9899 ( .A1(n8476), .A2(n9823), .A3(n8337), .ZN(n8481) );
  AOI22_X1 U9900 ( .A1(n8478), .A2(n9810), .B1(n9809), .B2(n8477), .ZN(n8479)
         );
  NAND3_X1 U9901 ( .A1(n8481), .A2(n8480), .A3(n8479), .ZN(n8529) );
  MUX2_X1 U9902 ( .A(n8529), .B(P2_REG1_REG_20__SCAN_IN), .S(n9833), .Z(
        P2_U3540) );
  AOI21_X1 U9903 ( .B1(n9809), .B2(n8483), .A(n8482), .ZN(n8484) );
  OAI211_X1 U9904 ( .C1(n8486), .C2(n9804), .A(n8485), .B(n8484), .ZN(n8530)
         );
  MUX2_X1 U9905 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8530), .S(n4268), .Z(
        P2_U3539) );
  AOI22_X1 U9906 ( .A1(n8488), .A2(n9810), .B1(n9809), .B2(n8487), .ZN(n8489)
         );
  OAI211_X1 U9907 ( .C1(n8491), .C2(n9804), .A(n8490), .B(n8489), .ZN(n8531)
         );
  MUX2_X1 U9908 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8531), .S(n4268), .Z(
        P2_U3538) );
  AOI21_X1 U9909 ( .B1(n9809), .B2(n8493), .A(n8492), .ZN(n8494) );
  OAI211_X1 U9910 ( .C1(n8496), .C2(n9804), .A(n8495), .B(n8494), .ZN(n8532)
         );
  MUX2_X1 U9911 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8532), .S(n4268), .Z(
        P2_U3537) );
  INV_X1 U9912 ( .A(n9814), .ZN(n9786) );
  OAI22_X1 U9913 ( .A1(n8498), .A2(n9781), .B1(n8497), .B2(n9820), .ZN(n8499)
         );
  AOI21_X1 U9914 ( .B1(n8500), .B2(n9786), .A(n8499), .ZN(n8501) );
  NAND2_X1 U9915 ( .A1(n8502), .A2(n8501), .ZN(n8533) );
  MUX2_X1 U9916 ( .A(n8533), .B(P2_REG1_REG_16__SCAN_IN), .S(n9833), .Z(
        P2_U3536) );
  AOI22_X1 U9917 ( .A1(n8504), .A2(n9810), .B1(n9809), .B2(n8503), .ZN(n8505)
         );
  OAI211_X1 U9918 ( .C1(n8507), .C2(n9804), .A(n8506), .B(n8505), .ZN(n8534)
         );
  MUX2_X1 U9919 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8534), .S(n4268), .Z(
        P2_U3535) );
  AOI22_X1 U9920 ( .A1(n8509), .A2(n9810), .B1(n9809), .B2(n8508), .ZN(n8510)
         );
  OAI211_X1 U9921 ( .C1(n8512), .C2(n9804), .A(n8511), .B(n8510), .ZN(n8535)
         );
  MUX2_X1 U9922 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8535), .S(n4268), .Z(
        P2_U3534) );
  AOI22_X1 U9923 ( .A1(n8514), .A2(n9810), .B1(n9809), .B2(n8513), .ZN(n8515)
         );
  OAI21_X1 U9924 ( .B1(n8516), .B2(n9814), .A(n8515), .ZN(n8517) );
  OR2_X1 U9925 ( .A1(n8518), .A2(n8517), .ZN(n8536) );
  MUX2_X1 U9926 ( .A(n8536), .B(P2_REG1_REG_13__SCAN_IN), .S(n9833), .Z(
        P2_U3533) );
  MUX2_X1 U9927 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8519), .S(n4267), .Z(
        P2_U3519) );
  MUX2_X1 U9928 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8520), .S(n4267), .Z(
        P2_U3517) );
  MUX2_X1 U9929 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8521), .S(n4267), .Z(
        P2_U3516) );
  MUX2_X1 U9930 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8522), .S(n4267), .Z(
        P2_U3515) );
  MUX2_X1 U9931 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8524), .S(n4267), .Z(
        P2_U3513) );
  MUX2_X1 U9932 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8525), .S(n4267), .Z(
        P2_U3512) );
  MUX2_X1 U9933 ( .A(n8526), .B(P2_REG0_REG_23__SCAN_IN), .S(n9825), .Z(
        P2_U3511) );
  MUX2_X1 U9934 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8527), .S(n4267), .Z(
        P2_U3510) );
  MUX2_X1 U9935 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8528), .S(n4267), .Z(
        P2_U3509) );
  MUX2_X1 U9936 ( .A(n8529), .B(P2_REG0_REG_20__SCAN_IN), .S(n9825), .Z(
        P2_U3508) );
  MUX2_X1 U9937 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8530), .S(n4267), .Z(
        P2_U3507) );
  MUX2_X1 U9938 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8531), .S(n4267), .Z(
        P2_U3505) );
  MUX2_X1 U9939 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8532), .S(n4267), .Z(
        P2_U3502) );
  MUX2_X1 U9940 ( .A(n8533), .B(P2_REG0_REG_16__SCAN_IN), .S(n9825), .Z(
        P2_U3499) );
  MUX2_X1 U9941 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8534), .S(n4267), .Z(
        P2_U3496) );
  MUX2_X1 U9942 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8535), .S(n4267), .Z(
        P2_U3493) );
  MUX2_X1 U9943 ( .A(n8536), .B(P2_REG0_REG_13__SCAN_IN), .S(n9825), .Z(
        P2_U3490) );
  INV_X1 U9944 ( .A(n8743), .ZN(n8542) );
  INV_X1 U9945 ( .A(n8537), .ZN(n8538) );
  NOR4_X1 U9946 ( .A1(n8538), .A2(P2_IR_REG_30__SCAN_IN), .A3(n4853), .A4(
        P2_U3152), .ZN(n8539) );
  AOI21_X1 U9947 ( .B1(n8540), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8539), .ZN(
        n8541) );
  OAI21_X1 U9948 ( .B1(n8542), .B2(n4270), .A(n8541), .ZN(P2_U3327) );
  INV_X1 U9949 ( .A(n9324), .ZN(n8543) );
  OAI222_X1 U9950 ( .A1(n8545), .A2(n8544), .B1(n4270), .B2(n8543), .C1(n5115), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  INV_X1 U9951 ( .A(n8546), .ZN(n8547) );
  MUX2_X1 U9952 ( .A(n8547), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U9953 ( .A(n8549), .B(n8548), .ZN(n8550) );
  XNOR2_X1 U9954 ( .A(n8551), .B(n8550), .ZN(n8557) );
  INV_X1 U9955 ( .A(n9114), .ZN(n9085) );
  OAI22_X1 U9956 ( .A1(n9085), .A2(n8656), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8552), .ZN(n8553) );
  AOI21_X1 U9957 ( .B1(n9088), .B2(n8660), .A(n8553), .ZN(n8554) );
  OAI21_X1 U9958 ( .B1(n9084), .B2(n8657), .A(n8554), .ZN(n8555) );
  AOI21_X1 U9959 ( .B1(n9245), .B2(n8648), .A(n8555), .ZN(n8556) );
  OAI21_X1 U9960 ( .B1(n8557), .B2(n8650), .A(n8556), .ZN(P1_U3212) );
  NAND2_X1 U9961 ( .A1(n8559), .A2(n8558), .ZN(n8561) );
  XNOR2_X1 U9962 ( .A(n8561), .B(n8560), .ZN(n8566) );
  AOI22_X1 U9963 ( .A1(n9015), .A2(n8644), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8563) );
  NAND2_X1 U9964 ( .A1(n9167), .A2(n8633), .ZN(n8562) );
  OAI211_X1 U9965 ( .C1(n8646), .C2(n9145), .A(n8563), .B(n8562), .ZN(n8564)
         );
  AOI21_X1 U9966 ( .B1(n9267), .B2(n8648), .A(n8564), .ZN(n8565) );
  OAI21_X1 U9967 ( .B1(n8566), .B2(n8650), .A(n8565), .ZN(P1_U3214) );
  OAI21_X1 U9968 ( .B1(n8569), .B2(n4443), .A(n8568), .ZN(n8570) );
  OAI21_X1 U9969 ( .B1(n8571), .B2(n4443), .A(n8570), .ZN(n8572) );
  NAND2_X1 U9970 ( .A1(n8572), .A2(n8652), .ZN(n8576) );
  INV_X1 U9971 ( .A(n9204), .ZN(n9009) );
  NAND2_X1 U9972 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8987) );
  OAI21_X1 U9973 ( .B1(n8657), .B2(n9009), .A(n8987), .ZN(n8574) );
  NOR2_X1 U9974 ( .A1(n8646), .A2(n9197), .ZN(n8573) );
  AOI211_X1 U9975 ( .C1(n8633), .C2(n9205), .A(n8574), .B(n8573), .ZN(n8575)
         );
  OAI211_X1 U9976 ( .C1(n9200), .C2(n8663), .A(n8576), .B(n8575), .ZN(P1_U3217) );
  OAI21_X1 U9977 ( .B1(n8578), .B2(n8577), .A(n7487), .ZN(n8579) );
  NAND2_X1 U9978 ( .A1(n8579), .A2(n8652), .ZN(n8583) );
  AOI22_X1 U9979 ( .A1(n8633), .A2(n5463), .B1(n8644), .B2(n6029), .ZN(n8582)
         );
  AOI22_X1 U9980 ( .A1(n8648), .A2(n8682), .B1(n8580), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n8581) );
  NAND3_X1 U9981 ( .A1(n8583), .A2(n8582), .A3(n8581), .ZN(P1_U3220) );
  XOR2_X1 U9982 ( .A(n8585), .B(n8584), .Z(n8590) );
  AOI22_X1 U9983 ( .A1(n9167), .A2(n8644), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8587) );
  NAND2_X1 U9984 ( .A1(n8660), .A2(n9174), .ZN(n8586) );
  OAI211_X1 U9985 ( .C1(n9009), .C2(n8656), .A(n8587), .B(n8586), .ZN(n8588)
         );
  AOI21_X1 U9986 ( .B1(n9277), .B2(n8648), .A(n8588), .ZN(n8589) );
  OAI21_X1 U9987 ( .B1(n8590), .B2(n8650), .A(n8589), .ZN(P1_U3221) );
  XOR2_X1 U9988 ( .A(n8592), .B(n8591), .Z(n8598) );
  OAI22_X1 U9989 ( .A1(n9140), .A2(n8656), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8593), .ZN(n8594) );
  AOI21_X1 U9990 ( .B1(n9114), .B2(n8644), .A(n8594), .ZN(n8595) );
  OAI21_X1 U9991 ( .B1(n8646), .B2(n9109), .A(n8595), .ZN(n8596) );
  AOI21_X1 U9992 ( .B1(n9253), .B2(n8648), .A(n8596), .ZN(n8597) );
  OAI21_X1 U9993 ( .B1(n8598), .B2(n8650), .A(n8597), .ZN(P1_U3223) );
  INV_X1 U9994 ( .A(n8599), .ZN(n8600) );
  AOI21_X1 U9995 ( .B1(n8602), .B2(n8601), .A(n8600), .ZN(n8609) );
  NOR2_X1 U9996 ( .A1(n8603), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9554) );
  AOI21_X1 U9997 ( .B1(n8633), .B2(n8942), .A(n9554), .ZN(n8606) );
  NAND2_X1 U9998 ( .A1(n8660), .A2(n8604), .ZN(n8605) );
  OAI211_X1 U9999 ( .C1(n8718), .C2(n8657), .A(n8606), .B(n8605), .ZN(n8607)
         );
  AOI21_X1 U10000 ( .B1(n9299), .B2(n8648), .A(n8607), .ZN(n8608) );
  OAI21_X1 U10001 ( .B1(n8609), .B2(n8650), .A(n8608), .ZN(P1_U3226) );
  XOR2_X1 U10002 ( .A(n8611), .B(n8610), .Z(n8616) );
  AOI22_X1 U10003 ( .A1(n9160), .A2(n8633), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8613) );
  NAND2_X1 U10004 ( .A1(n9127), .A2(n8660), .ZN(n8612) );
  OAI211_X1 U10005 ( .C1(n9017), .C2(n8657), .A(n8613), .B(n8612), .ZN(n8614)
         );
  AOI21_X1 U10006 ( .B1(n9261), .B2(n8648), .A(n8614), .ZN(n8615) );
  OAI21_X1 U10007 ( .B1(n8616), .B2(n8650), .A(n8615), .ZN(P1_U3227) );
  INV_X1 U10008 ( .A(n9284), .ZN(n9191) );
  OAI21_X1 U10009 ( .B1(n8619), .B2(n8618), .A(n8617), .ZN(n8620) );
  NAND2_X1 U10010 ( .A1(n8620), .A2(n8652), .ZN(n8625) );
  OAI22_X1 U10011 ( .A1(n8657), .A2(n9184), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8621), .ZN(n8623) );
  NOR2_X1 U10012 ( .A1(n8646), .A2(n9187), .ZN(n8622) );
  AOI211_X1 U10013 ( .C1(n8633), .C2(n9222), .A(n8623), .B(n8622), .ZN(n8624)
         );
  OAI211_X1 U10014 ( .C1(n9191), .C2(n8663), .A(n8625), .B(n8624), .ZN(
        P1_U3231) );
  INV_X1 U10015 ( .A(n8626), .ZN(n8628) );
  INV_X1 U10016 ( .A(n8630), .ZN(n8627) );
  OAI21_X1 U10017 ( .B1(n8631), .B2(n8628), .A(n8627), .ZN(n8632) );
  AOI22_X1 U10018 ( .A1(n8632), .A2(n4429), .B1(n8631), .B2(n8630), .ZN(n8638)
         );
  AOI22_X1 U10019 ( .A1(n9160), .A2(n8644), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8635) );
  NAND2_X1 U10020 ( .A1(n8633), .A2(n9161), .ZN(n8634) );
  OAI211_X1 U10021 ( .C1(n8646), .C2(n9154), .A(n8635), .B(n8634), .ZN(n8636)
         );
  AOI21_X1 U10022 ( .B1(n9270), .B2(n8648), .A(n8636), .ZN(n8637) );
  OAI21_X1 U10023 ( .B1(n8638), .B2(n8650), .A(n8637), .ZN(P1_U3233) );
  NAND2_X1 U10024 ( .A1(n8640), .A2(n8639), .ZN(n8641) );
  XOR2_X1 U10025 ( .A(n8642), .B(n8641), .Z(n8651) );
  NAND2_X1 U10026 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9563) );
  OAI21_X1 U10027 ( .B1(n8656), .B2(n9002), .A(n9563), .ZN(n8643) );
  AOI21_X1 U10028 ( .B1(n8644), .B2(n9222), .A(n8643), .ZN(n8645) );
  OAI21_X1 U10029 ( .B1(n8646), .B2(n9216), .A(n8645), .ZN(n8647) );
  AOI21_X1 U10030 ( .B1(n9292), .B2(n8648), .A(n8647), .ZN(n8649) );
  OAI21_X1 U10031 ( .B1(n8651), .B2(n8650), .A(n8649), .ZN(P1_U3236) );
  OAI211_X1 U10032 ( .C1(n8655), .C2(n8654), .A(n8653), .B(n8652), .ZN(n8662)
         );
  OAI22_X1 U10033 ( .A1(n9017), .A2(n8656), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9925), .ZN(n8659) );
  NOR2_X1 U10034 ( .A1(n9075), .A2(n8657), .ZN(n8658) );
  AOI211_X1 U10035 ( .C1(n9096), .C2(n8660), .A(n8659), .B(n8658), .ZN(n8661)
         );
  OAI211_X1 U10036 ( .C1(n9098), .C2(n8663), .A(n8662), .B(n8661), .ZN(
        P1_U3238) );
  NAND2_X1 U10037 ( .A1(n8664), .A2(n6363), .ZN(n8666) );
  OR2_X1 U10038 ( .A1(n8732), .A2(n9322), .ZN(n8665) );
  INV_X1 U10039 ( .A(n8879), .ZN(n8667) );
  NAND2_X1 U10040 ( .A1(n8667), .A2(n9048), .ZN(n8774) );
  INV_X1 U10041 ( .A(n8774), .ZN(n8741) );
  NAND2_X1 U10042 ( .A1(n9245), .A2(n9075), .ZN(n8871) );
  INV_X1 U10043 ( .A(n8871), .ZN(n8669) );
  NAND2_X1 U10044 ( .A1(n9248), .A2(n9085), .ZN(n9045) );
  INV_X1 U10045 ( .A(n9045), .ZN(n8668) );
  OAI21_X1 U10046 ( .B1(n8669), .B2(n8668), .A(n9047), .ZN(n8670) );
  NAND2_X1 U10047 ( .A1(n8670), .A2(n9050), .ZN(n8769) );
  INV_X1 U10048 ( .A(n8769), .ZN(n8729) );
  INV_X1 U10049 ( .A(n9160), .ZN(n9012) );
  NAND2_X1 U10050 ( .A1(n9267), .A2(n9012), .ZN(n8891) );
  AND2_X1 U10051 ( .A1(n9042), .A2(n8891), .ZN(n8749) );
  NAND2_X1 U10052 ( .A1(n9292), .A2(n8718), .ZN(n9030) );
  NAND2_X1 U10053 ( .A1(n9030), .A2(n9027), .ZN(n8785) );
  INV_X1 U10054 ( .A(n8837), .ZN(n8678) );
  OR2_X1 U10055 ( .A1(n9391), .A2(n8944), .ZN(n8827) );
  NAND2_X1 U10056 ( .A1(n8819), .A2(n8671), .ZN(n8799) );
  INV_X1 U10057 ( .A(n8815), .ZN(n8672) );
  NOR2_X1 U10058 ( .A1(n8793), .A2(n8672), .ZN(n8673) );
  NOR2_X1 U10059 ( .A1(n8799), .A2(n8673), .ZN(n8674) );
  AND2_X1 U10060 ( .A1(n8674), .A2(n8828), .ZN(n8700) );
  NAND2_X1 U10061 ( .A1(n8675), .A2(n8808), .ZN(n8790) );
  INV_X1 U10062 ( .A(n8790), .ZN(n8676) );
  NAND3_X1 U10063 ( .A1(n8827), .A2(n8700), .A3(n8676), .ZN(n8677) );
  OR3_X1 U10064 ( .A1(n8785), .A2(n8678), .A3(n8677), .ZN(n8762) );
  INV_X1 U10065 ( .A(n8762), .ZN(n8715) );
  INV_X1 U10066 ( .A(n8679), .ZN(n8680) );
  OAI211_X1 U10067 ( .C1(n8682), .C2(n8681), .A(n8931), .B(n8680), .ZN(n8683)
         );
  NAND3_X1 U10068 ( .A1(n8685), .A2(n8684), .A3(n8683), .ZN(n8689) );
  INV_X1 U10069 ( .A(n8686), .ZN(n8687) );
  AOI21_X1 U10070 ( .B1(n8689), .B2(n8688), .A(n8687), .ZN(n8696) );
  AND2_X1 U10071 ( .A1(n8691), .A2(n8690), .ZN(n8756) );
  INV_X1 U10072 ( .A(n8756), .ZN(n8695) );
  NAND2_X1 U10073 ( .A1(n8809), .A2(n8692), .ZN(n8751) );
  INV_X1 U10074 ( .A(n8751), .ZN(n8694) );
  OAI211_X1 U10075 ( .C1(n8696), .C2(n8695), .A(n8694), .B(n8693), .ZN(n8699)
         );
  INV_X1 U10076 ( .A(n8697), .ZN(n8698) );
  NAND2_X1 U10077 ( .A1(n8698), .A2(n8809), .ZN(n8755) );
  NAND3_X1 U10078 ( .A1(n8699), .A2(n8811), .A3(n8755), .ZN(n8714) );
  INV_X1 U10079 ( .A(n8840), .ZN(n8712) );
  INV_X1 U10080 ( .A(n8700), .ZN(n8707) );
  INV_X1 U10081 ( .A(n8701), .ZN(n8702) );
  NOR2_X1 U10082 ( .A1(n8814), .A2(n8702), .ZN(n8792) );
  AND2_X1 U10083 ( .A1(n8792), .A2(n8815), .ZN(n8812) );
  NAND2_X1 U10084 ( .A1(n8798), .A2(n8703), .ZN(n8704) );
  NAND2_X1 U10085 ( .A1(n8704), .A2(n8819), .ZN(n8705) );
  NAND2_X1 U10086 ( .A1(n8804), .A2(n8705), .ZN(n8797) );
  NAND2_X1 U10087 ( .A1(n8797), .A2(n8828), .ZN(n8706) );
  OAI211_X1 U10088 ( .C1(n8707), .C2(n8812), .A(n8706), .B(n8805), .ZN(n8708)
         );
  AND3_X1 U10089 ( .A1(n8709), .A2(n8708), .A3(n8827), .ZN(n8710) );
  NOR2_X1 U10090 ( .A1(n8835), .A2(n8710), .ZN(n8711) );
  OR3_X1 U10091 ( .A1(n8785), .A2(n8712), .A3(n8711), .ZN(n8760) );
  INV_X1 U10092 ( .A(n8760), .ZN(n8713) );
  AOI21_X1 U10093 ( .B1(n8715), .B2(n8714), .A(n8713), .ZN(n8725) );
  NAND2_X1 U10094 ( .A1(n9270), .A2(n9141), .ZN(n9038) );
  OR2_X1 U10095 ( .A1(n9277), .A2(n9184), .ZN(n8892) );
  AND2_X1 U10096 ( .A1(n9284), .A2(n9009), .ZN(n9034) );
  NAND2_X1 U10097 ( .A1(n8892), .A2(n9034), .ZN(n8716) );
  NAND2_X1 U10098 ( .A1(n9277), .A2(n9184), .ZN(n9035) );
  AND2_X1 U10099 ( .A1(n8716), .A2(n9035), .ZN(n8717) );
  NAND2_X1 U10100 ( .A1(n9038), .A2(n8717), .ZN(n8721) );
  INV_X1 U10101 ( .A(n9222), .ZN(n9185) );
  NAND2_X1 U10102 ( .A1(n9288), .A2(n9185), .ZN(n9032) );
  NOR2_X1 U10103 ( .A1(n8721), .A2(n4503), .ZN(n8764) );
  INV_X1 U10104 ( .A(n8764), .ZN(n8724) );
  AND2_X1 U10105 ( .A1(n9037), .A2(n8892), .ZN(n8856) );
  INV_X1 U10106 ( .A(n8856), .ZN(n8859) );
  OR2_X1 U10107 ( .A1(n9292), .A2(n8718), .ZN(n8895) );
  NAND2_X1 U10108 ( .A1(n8895), .A2(n4508), .ZN(n8786) );
  INV_X1 U10109 ( .A(n8786), .ZN(n8720) );
  AND2_X1 U10110 ( .A1(n9032), .A2(n9030), .ZN(n8848) );
  INV_X1 U10111 ( .A(n8848), .ZN(n8719) );
  OR2_X1 U10112 ( .A1(n9284), .A2(n9009), .ZN(n9033) );
  OR2_X1 U10113 ( .A1(n9288), .A2(n9185), .ZN(n8894) );
  AND2_X1 U10114 ( .A1(n9033), .A2(n8894), .ZN(n8850) );
  OAI21_X1 U10115 ( .B1(n8720), .B2(n8719), .A(n8850), .ZN(n8722) );
  NAND2_X1 U10116 ( .A1(n8721), .A2(n9037), .ZN(n8858) );
  OAI21_X1 U10117 ( .B1(n8859), .B2(n8722), .A(n8858), .ZN(n8723) );
  AND2_X1 U10118 ( .A1(n8723), .A2(n9119), .ZN(n8766) );
  OAI21_X1 U10119 ( .B1(n8725), .B2(n8724), .A(n8766), .ZN(n8726) );
  NAND2_X1 U10120 ( .A1(n9043), .A2(n8890), .ZN(n8783) );
  AOI21_X1 U10121 ( .B1(n8749), .B2(n8726), .A(n8783), .ZN(n8727) );
  INV_X1 U10122 ( .A(n9046), .ZN(n8782) );
  OAI211_X1 U10123 ( .C1(n9044), .C2(n8727), .A(n9022), .B(n8782), .ZN(n8728)
         );
  NAND2_X1 U10124 ( .A1(n8729), .A2(n8728), .ZN(n8740) );
  NAND2_X1 U10125 ( .A1(n8730), .A2(n6363), .ZN(n8734) );
  OR2_X1 U10126 ( .A1(n8732), .A2(n8731), .ZN(n8733) );
  NAND2_X1 U10127 ( .A1(n7983), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U10128 ( .A1(n4275), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8737) );
  NAND2_X1 U10129 ( .A1(n8735), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8736) );
  AND3_X1 U10130 ( .A1(n8738), .A2(n8737), .A3(n8736), .ZN(n9054) );
  NAND2_X1 U10131 ( .A1(n9373), .A2(n9054), .ZN(n8919) );
  INV_X1 U10132 ( .A(n8919), .ZN(n8739) );
  AOI211_X1 U10133 ( .C1(n8741), .C2(n8740), .A(n8878), .B(n8739), .ZN(n8745)
         );
  NOR2_X1 U10134 ( .A1(n8732), .A2(n4993), .ZN(n8742) );
  NOR2_X1 U10135 ( .A1(n8993), .A2(n8771), .ZN(n8778) );
  NOR2_X1 U10136 ( .A1(n9373), .A2(n9054), .ZN(n8747) );
  NOR2_X1 U10137 ( .A1(n8778), .A2(n8747), .ZN(n8921) );
  INV_X1 U10138 ( .A(n8921), .ZN(n8744) );
  INV_X1 U10139 ( .A(n8771), .ZN(n8991) );
  OAI21_X1 U10140 ( .B1(n8745), .B2(n8744), .A(n8924), .ZN(n8746) );
  XNOR2_X1 U10141 ( .A(n8746), .B(n9588), .ZN(n8933) );
  AOI21_X1 U10142 ( .B1(n8747), .B2(n9229), .A(n8778), .ZN(n8881) );
  INV_X1 U10143 ( .A(n8890), .ZN(n8748) );
  OAI21_X1 U10144 ( .B1(n8749), .B2(n8748), .A(n8889), .ZN(n8784) );
  INV_X1 U10145 ( .A(n8784), .ZN(n8768) );
  INV_X1 U10146 ( .A(n8750), .ZN(n8753) );
  AOI21_X1 U10147 ( .B1(n8753), .B2(n8752), .A(n8751), .ZN(n8759) );
  AND2_X1 U10148 ( .A1(n8811), .A2(n8754), .ZN(n8791) );
  INV_X1 U10149 ( .A(n8791), .ZN(n8758) );
  NAND4_X1 U10150 ( .A1(n9606), .A2(n8756), .A3(n8755), .A4(n8811), .ZN(n8757)
         );
  OAI21_X1 U10151 ( .B1(n8759), .B2(n8758), .A(n8757), .ZN(n8761) );
  OAI21_X1 U10152 ( .B1(n8762), .B2(n8761), .A(n8760), .ZN(n8763) );
  NAND2_X1 U10153 ( .A1(n8764), .A2(n8763), .ZN(n8765) );
  NAND3_X1 U10154 ( .A1(n8766), .A2(n8890), .A3(n8765), .ZN(n8767) );
  AOI211_X1 U10155 ( .C1(n8768), .C2(n8767), .A(n4538), .B(n9046), .ZN(n8770)
         );
  AOI21_X1 U10156 ( .B1(n8770), .B2(n9047), .A(n8769), .ZN(n8775) );
  INV_X1 U10157 ( .A(n9054), .ZN(n8939) );
  NAND2_X1 U10158 ( .A1(n8939), .A2(n8771), .ZN(n8772) );
  AND2_X1 U10159 ( .A1(n9373), .A2(n8772), .ZN(n8779) );
  INV_X1 U10160 ( .A(n8779), .ZN(n8880) );
  INV_X1 U10161 ( .A(n8878), .ZN(n8773) );
  OAI211_X1 U10162 ( .C1(n8775), .C2(n8774), .A(n8880), .B(n8773), .ZN(n8777)
         );
  INV_X1 U10163 ( .A(n8924), .ZN(n8776) );
  AOI21_X1 U10164 ( .B1(n8881), .B2(n8777), .A(n8776), .ZN(n8888) );
  INV_X1 U10165 ( .A(n8778), .ZN(n8780) );
  NAND2_X1 U10166 ( .A1(n8780), .A2(n8779), .ZN(n8781) );
  MUX2_X1 U10167 ( .A(n8881), .B(n8781), .S(n8877), .Z(n8885) );
  INV_X1 U10168 ( .A(n9072), .ZN(n8874) );
  MUX2_X1 U10169 ( .A(n9045), .B(n8782), .S(n8877), .Z(n8870) );
  MUX2_X1 U10170 ( .A(n8784), .B(n8783), .S(n8877), .Z(n8868) );
  INV_X1 U10171 ( .A(n8877), .ZN(n8801) );
  MUX2_X1 U10172 ( .A(n8786), .B(n8785), .S(n8801), .Z(n8787) );
  INV_X1 U10173 ( .A(n8787), .ZN(n8846) );
  XNOR2_X1 U10174 ( .A(n8788), .B(n8801), .ZN(n8789) );
  NAND2_X1 U10175 ( .A1(n8789), .A2(n8904), .ZN(n8810) );
  AOI21_X1 U10176 ( .B1(n8810), .B2(n8791), .A(n8790), .ZN(n8795) );
  INV_X1 U10177 ( .A(n8792), .ZN(n8794) );
  OAI21_X1 U10178 ( .B1(n8795), .B2(n8794), .A(n8793), .ZN(n8796) );
  NAND3_X1 U10179 ( .A1(n8796), .A2(n8815), .A3(n8798), .ZN(n8807) );
  NAND2_X1 U10180 ( .A1(n8805), .A2(n8877), .ZN(n8826) );
  OR2_X1 U10181 ( .A1(n8826), .A2(n8797), .ZN(n8803) );
  NAND2_X1 U10182 ( .A1(n8799), .A2(n8798), .ZN(n8800) );
  NAND4_X1 U10183 ( .A1(n8827), .A2(n8801), .A3(n8828), .A4(n8800), .ZN(n8802)
         );
  NAND2_X1 U10184 ( .A1(n8803), .A2(n8802), .ZN(n8831) );
  NAND2_X1 U10185 ( .A1(n8805), .A2(n8804), .ZN(n8806) );
  AOI22_X1 U10186 ( .A1(n8807), .A2(n8831), .B1(n8827), .B2(n8806), .ZN(n8834)
         );
  NAND3_X1 U10187 ( .A1(n8810), .A2(n8809), .A3(n8808), .ZN(n8813) );
  NAND3_X1 U10188 ( .A1(n8813), .A2(n8812), .A3(n8811), .ZN(n8821) );
  OAI211_X1 U10189 ( .C1(n8817), .C2(n8816), .A(n4524), .B(n8815), .ZN(n8818)
         );
  NAND4_X1 U10190 ( .A1(n8821), .A2(n8820), .A3(n8819), .A4(n8818), .ZN(n8822)
         );
  NAND2_X1 U10191 ( .A1(n8822), .A2(n8877), .ZN(n8825) );
  NAND2_X1 U10192 ( .A1(n8824), .A2(n8823), .ZN(n9355) );
  NAND2_X1 U10193 ( .A1(n8825), .A2(n9355), .ZN(n8832) );
  AOI21_X1 U10194 ( .B1(n8828), .B2(n8827), .A(n8826), .ZN(n8829) );
  AOI211_X1 U10195 ( .C1(n8832), .C2(n8831), .A(n8830), .B(n8829), .ZN(n8833)
         );
  OAI21_X1 U10196 ( .B1(n8834), .B2(n8877), .A(n8833), .ZN(n8839) );
  INV_X1 U10197 ( .A(n8835), .ZN(n8836) );
  MUX2_X1 U10198 ( .A(n8837), .B(n8836), .S(n8877), .Z(n8838) );
  NAND2_X1 U10199 ( .A1(n8839), .A2(n8838), .ZN(n8844) );
  MUX2_X1 U10200 ( .A(n8841), .B(n8840), .S(n8877), .Z(n8842) );
  NAND3_X1 U10201 ( .A1(n8844), .A2(n8843), .A3(n8842), .ZN(n8845) );
  NAND2_X1 U10202 ( .A1(n8846), .A2(n8845), .ZN(n8849) );
  NAND3_X1 U10203 ( .A1(n8849), .A2(n8895), .A3(n8894), .ZN(n8847) );
  INV_X1 U10204 ( .A(n9034), .ZN(n8893) );
  NAND3_X1 U10205 ( .A1(n8847), .A2(n9032), .A3(n8893), .ZN(n8853) );
  NAND2_X1 U10206 ( .A1(n8849), .A2(n8848), .ZN(n8851) );
  NAND2_X1 U10207 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  MUX2_X1 U10208 ( .A(n8853), .B(n8852), .S(n8877), .Z(n8860) );
  INV_X1 U10209 ( .A(n8860), .ZN(n8854) );
  OAI21_X1 U10210 ( .B1(n8854), .B2(n4498), .A(n9035), .ZN(n8857) );
  INV_X1 U10211 ( .A(n9038), .ZN(n8855) );
  AOI21_X1 U10212 ( .B1(n8857), .B2(n8856), .A(n8855), .ZN(n8862) );
  OAI211_X1 U10213 ( .C1(n8860), .C2(n8859), .A(n8858), .B(n8891), .ZN(n8861)
         );
  MUX2_X1 U10214 ( .A(n8862), .B(n8861), .S(n8877), .Z(n8865) );
  NAND2_X1 U10215 ( .A1(n8890), .A2(n9119), .ZN(n8863) );
  MUX2_X1 U10216 ( .A(n8863), .B(n4527), .S(n8877), .Z(n8864) );
  AOI21_X1 U10217 ( .B1(n8865), .B2(n9119), .A(n8864), .ZN(n8867) );
  MUX2_X1 U10218 ( .A(n9043), .B(n8889), .S(n8877), .Z(n8866) );
  NAND2_X1 U10219 ( .A1(n9248), .A2(n9114), .ZN(n9021) );
  NAND2_X1 U10220 ( .A1(n9020), .A2(n9021), .ZN(n9100) );
  OAI211_X1 U10221 ( .C1(n8868), .C2(n8867), .A(n8866), .B(n9100), .ZN(n8869)
         );
  NAND3_X1 U10222 ( .A1(n8870), .A2(n9022), .A3(n8869), .ZN(n8873) );
  MUX2_X1 U10223 ( .A(n9047), .B(n8871), .S(n8877), .Z(n8872) );
  NAND3_X1 U10224 ( .A1(n8874), .A2(n8873), .A3(n8872), .ZN(n8876) );
  MUX2_X1 U10225 ( .A(n9050), .B(n9048), .S(n8877), .Z(n8875) );
  AND3_X1 U10226 ( .A1(n9025), .A2(n8876), .A3(n8875), .ZN(n8883) );
  MUX2_X1 U10227 ( .A(n8879), .B(n8878), .S(n8877), .Z(n8882) );
  OAI211_X1 U10228 ( .C1(n8883), .C2(n8882), .A(n8881), .B(n8880), .ZN(n8884)
         );
  NAND2_X1 U10229 ( .A1(n8885), .A2(n8884), .ZN(n8927) );
  NAND3_X1 U10230 ( .A1(n8927), .A2(n8886), .A3(n8924), .ZN(n8887) );
  OAI21_X1 U10231 ( .B1(n9588), .B2(n8888), .A(n8887), .ZN(n8930) );
  INV_X1 U10232 ( .A(n9025), .ZN(n9051) );
  INV_X1 U10233 ( .A(n9130), .ZN(n9122) );
  NAND2_X1 U10234 ( .A1(n9119), .A2(n8891), .ZN(n9138) );
  NAND2_X1 U10235 ( .A1(n9037), .A2(n9038), .ZN(n9159) );
  AND2_X1 U10236 ( .A1(n8893), .A2(n9033), .ZN(n9182) );
  NAND2_X1 U10237 ( .A1(n8895), .A2(n9030), .ZN(n9211) );
  INV_X1 U10238 ( .A(n9211), .ZN(n9220) );
  INV_X1 U10239 ( .A(n9355), .ZN(n9348) );
  NAND4_X1 U10240 ( .A1(n8899), .A2(n8898), .A3(n9607), .A4(n8897), .ZN(n8901)
         );
  INV_X1 U10241 ( .A(n8900), .ZN(n9590) );
  NAND4_X1 U10242 ( .A1(n4333), .A2(n8904), .A3(n8903), .A4(n8902), .ZN(n8906)
         );
  NOR4_X1 U10243 ( .A1(n9348), .A2(n6601), .A3(n8906), .A4(n8905), .ZN(n8907)
         );
  NAND4_X1 U10244 ( .A1(n8910), .A2(n8909), .A3(n8908), .A4(n8907), .ZN(n8911)
         );
  NOR4_X1 U10245 ( .A1(n8914), .A2(n8913), .A3(n8912), .A4(n8911), .ZN(n8915)
         );
  NAND4_X1 U10246 ( .A1(n9182), .A2(n9203), .A3(n9220), .A4(n8915), .ZN(n8916)
         );
  NOR4_X1 U10247 ( .A1(n9138), .A2(n9159), .A3(n9169), .A4(n8916), .ZN(n8917)
         );
  NAND4_X1 U10248 ( .A1(n9113), .A2(n9122), .A3(n8917), .A4(n9100), .ZN(n8918)
         );
  NOR4_X1 U10249 ( .A1(n9051), .A2(n9082), .A3(n9072), .A4(n8918), .ZN(n8920)
         );
  AND4_X1 U10250 ( .A1(n8921), .A2(n8920), .A3(n8924), .A4(n8919), .ZN(n8925)
         );
  INV_X1 U10251 ( .A(n8925), .ZN(n8922) );
  NOR2_X1 U10252 ( .A1(n8922), .A2(n8931), .ZN(n8929) );
  NAND2_X1 U10253 ( .A1(n8924), .A2(n8923), .ZN(n8926) );
  OAI22_X1 U10254 ( .A1(n8927), .A2(n8926), .B1(n8931), .B2(n8925), .ZN(n8928)
         );
  NAND4_X1 U10255 ( .A1(n8935), .A2(n9630), .A3(n8934), .A4(n8989), .ZN(n8936)
         );
  OAI211_X1 U10256 ( .C1(n5393), .C2(n8938), .A(n8936), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8937) );
  MUX2_X1 U10257 ( .A(n8939), .B(P1_DATAO_REG_30__SCAN_IN), .S(n8954), .Z(
        P1_U3585) );
  MUX2_X1 U10258 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8940), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10259 ( .A(n8941), .B(P1_DATAO_REG_28__SCAN_IN), .S(n8954), .Z(
        P1_U3583) );
  MUX2_X1 U10260 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9101), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10261 ( .A(n9114), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8954), .Z(
        P1_U3581) );
  MUX2_X1 U10262 ( .A(n9018), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8954), .Z(
        P1_U3580) );
  MUX2_X1 U10263 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9015), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10264 ( .A(n9160), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8954), .Z(
        P1_U3578) );
  MUX2_X1 U10265 ( .A(n9167), .B(P1_DATAO_REG_22__SCAN_IN), .S(n8954), .Z(
        P1_U3577) );
  MUX2_X1 U10266 ( .A(n9161), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8954), .Z(
        P1_U3576) );
  MUX2_X1 U10267 ( .A(n9204), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8954), .Z(
        P1_U3575) );
  MUX2_X1 U10268 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9222), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10269 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9205), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10270 ( .A(n9223), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8954), .Z(
        P1_U3572) );
  MUX2_X1 U10271 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8942), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10272 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8943), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10273 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8944), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10274 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8945), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10275 ( .A(n9356), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8954), .Z(
        P1_U3567) );
  MUX2_X1 U10276 ( .A(n8946), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8954), .Z(
        P1_U3566) );
  MUX2_X1 U10277 ( .A(n9358), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8954), .Z(
        P1_U3565) );
  MUX2_X1 U10278 ( .A(n8947), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8954), .Z(
        P1_U3564) );
  MUX2_X1 U10279 ( .A(n8948), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8954), .Z(
        P1_U3563) );
  MUX2_X1 U10280 ( .A(n8949), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8954), .Z(
        P1_U3562) );
  MUX2_X1 U10281 ( .A(n8950), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8954), .Z(
        P1_U3561) );
  MUX2_X1 U10282 ( .A(n8951), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8954), .Z(
        P1_U3560) );
  MUX2_X1 U10283 ( .A(n8952), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8954), .Z(
        P1_U3559) );
  MUX2_X1 U10284 ( .A(n8953), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8954), .Z(
        P1_U3558) );
  MUX2_X1 U10285 ( .A(n6029), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8954), .Z(
        P1_U3557) );
  MUX2_X1 U10286 ( .A(n5462), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8954), .Z(
        P1_U3556) );
  INV_X1 U10287 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8967) );
  XNOR2_X1 U10288 ( .A(n9571), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9574) );
  INV_X1 U10289 ( .A(n9555), .ZN(n8965) );
  INV_X1 U10290 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8964) );
  XOR2_X1 U10291 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9555), .Z(n9559) );
  INV_X1 U10292 ( .A(n9543), .ZN(n8963) );
  INV_X1 U10293 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9382) );
  NOR2_X1 U10294 ( .A1(n9543), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8955) );
  AOI21_X1 U10295 ( .B1(n9543), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8955), .ZN(
        n9546) );
  INV_X1 U10296 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9394) );
  INV_X1 U10297 ( .A(n9506), .ZN(n8960) );
  INV_X1 U10298 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9401) );
  INV_X1 U10299 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9407) );
  AOI21_X1 U10300 ( .B1(n8957), .B2(n9414), .A(n8956), .ZN(n9496) );
  NOR2_X1 U10301 ( .A1(n9493), .A2(n9407), .ZN(n8958) );
  AOI21_X1 U10302 ( .B1(n9493), .B2(n9407), .A(n8958), .ZN(n9495) );
  NOR2_X1 U10303 ( .A1(n9496), .A2(n9495), .ZN(n9494) );
  AOI21_X1 U10304 ( .B1(n4459), .B2(n9407), .A(n9494), .ZN(n9508) );
  NOR2_X1 U10305 ( .A1(n9506), .A2(n9401), .ZN(n8959) );
  AOI21_X1 U10306 ( .B1(n9506), .B2(n9401), .A(n8959), .ZN(n9509) );
  NOR2_X1 U10307 ( .A1(n9508), .A2(n9509), .ZN(n9507) );
  AOI21_X1 U10308 ( .B1(n8960), .B2(n9401), .A(n9507), .ZN(n9521) );
  NOR2_X1 U10309 ( .A1(n8973), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8961) );
  AOI21_X1 U10310 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n8973), .A(n8961), .ZN(
        n9522) );
  INV_X1 U10311 ( .A(n8962), .ZN(n9545) );
  NAND2_X1 U10312 ( .A1(n9546), .A2(n9545), .ZN(n9544) );
  OAI21_X1 U10313 ( .B1(n8963), .B2(n9382), .A(n9544), .ZN(n9558) );
  NAND2_X1 U10314 ( .A1(n9559), .A2(n9558), .ZN(n9556) );
  OAI21_X1 U10315 ( .B1(n8965), .B2(n8964), .A(n9556), .ZN(n9573) );
  INV_X1 U10316 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U10317 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9493), .ZN(n8968) );
  OAI21_X1 U10318 ( .B1(n9493), .B2(P1_REG2_REG_12__SCAN_IN), .A(n8968), .ZN(
        n9489) );
  NOR2_X1 U10319 ( .A1(n9489), .A2(n9490), .ZN(n9488) );
  NAND2_X1 U10320 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9506), .ZN(n8971) );
  OAI21_X1 U10321 ( .B1(n9506), .B2(P1_REG2_REG_13__SCAN_IN), .A(n8971), .ZN(
        n9502) );
  NOR2_X1 U10322 ( .A1(n8972), .A2(n8973), .ZN(n8974) );
  INV_X1 U10323 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9515) );
  NOR2_X1 U10324 ( .A1(n9515), .A2(n9516), .ZN(n9514) );
  INV_X1 U10325 ( .A(n8975), .ZN(n8976) );
  INV_X1 U10326 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U10327 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9543), .ZN(n8977) );
  OAI21_X1 U10328 ( .B1(n9543), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8977), .ZN(
        n9539) );
  NOR2_X1 U10329 ( .A1(n9540), .A2(n9539), .ZN(n9538) );
  AOI21_X1 U10330 ( .B1(n9543), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9538), .ZN(
        n9552) );
  NOR2_X1 U10331 ( .A1(n9555), .A2(n8979), .ZN(n8978) );
  AOI21_X1 U10332 ( .B1(n8979), .B2(n9555), .A(n8978), .ZN(n9551) );
  NOR2_X1 U10333 ( .A1(n9552), .A2(n9551), .ZN(n9550) );
  AOI21_X1 U10334 ( .B1(n9555), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9550), .ZN(
        n9567) );
  INV_X1 U10335 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8981) );
  NOR2_X1 U10336 ( .A1(n9571), .A2(n8981), .ZN(n8980) );
  AOI21_X1 U10337 ( .B1(n9571), .B2(n8981), .A(n8980), .ZN(n9566) );
  NOR2_X1 U10338 ( .A1(n9567), .A2(n9566), .ZN(n9565) );
  NAND2_X1 U10339 ( .A1(n8985), .A2(n9454), .ZN(n8982) );
  OAI211_X1 U10340 ( .C1(n8983), .C2(n9576), .A(n8982), .B(n9452), .ZN(n8986)
         );
  INV_X1 U10341 ( .A(n9292), .ZN(n9219) );
  OR2_X2 U10342 ( .A1(n9186), .A2(n9277), .ZN(n9172) );
  NOR2_X2 U10343 ( .A1(n9172), .A2(n9270), .ZN(n9153) );
  NAND2_X1 U10344 ( .A1(n9153), .A2(n9149), .ZN(n9142) );
  OR2_X2 U10345 ( .A1(n9142), .A2(n9261), .ZN(n9125) );
  NAND2_X1 U10346 ( .A1(n8996), .A2(n9056), .ZN(n8988) );
  XNOR2_X1 U10347 ( .A(n9229), .B(n8988), .ZN(n9231) );
  NAND2_X1 U10348 ( .A1(n8989), .A2(P1_B_REG_SCAN_IN), .ZN(n8990) );
  NAND2_X1 U10349 ( .A1(n9357), .A2(n8990), .ZN(n9055) );
  NOR2_X1 U10350 ( .A1(n9055), .A2(n8991), .ZN(n9372) );
  INV_X1 U10351 ( .A(n9372), .ZN(n8992) );
  NOR2_X1 U10352 ( .A1(n8992), .A2(n9598), .ZN(n8998) );
  NOR2_X1 U10353 ( .A1(n8993), .A2(n9619), .ZN(n8994) );
  AOI211_X1 U10354 ( .C1(n9598), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8998), .B(
        n8994), .ZN(n8995) );
  OAI21_X1 U10355 ( .B1(n9231), .B2(n9000), .A(n8995), .ZN(P1_U3261) );
  XNOR2_X1 U10356 ( .A(n8996), .B(n9056), .ZN(n9370) );
  NOR2_X1 U10357 ( .A1(n8996), .A2(n9619), .ZN(n8997) );
  AOI211_X1 U10358 ( .C1(n9598), .C2(P1_REG2_REG_30__SCAN_IN), .A(n8998), .B(
        n8997), .ZN(n8999) );
  OAI21_X1 U10359 ( .B1(n9000), .B2(n9370), .A(n8999), .ZN(P1_U3262) );
  NOR2_X1 U10360 ( .A1(n9299), .A2(n9223), .ZN(n9003) );
  NOR2_X1 U10361 ( .A1(n9288), .A2(n9222), .ZN(n9007) );
  INV_X1 U10362 ( .A(n9277), .ZN(n9176) );
  NAND2_X1 U10363 ( .A1(n9157), .A2(n9141), .ZN(n9011) );
  AOI21_X2 U10364 ( .B1(n9152), .B2(n9011), .A(n9010), .ZN(n9136) );
  NAND2_X1 U10365 ( .A1(n9267), .A2(n9160), .ZN(n9013) );
  INV_X1 U10366 ( .A(n9140), .ZN(n9015) );
  NAND2_X1 U10367 ( .A1(n9258), .A2(n9016), .ZN(n9107) );
  INV_X1 U10368 ( .A(n9017), .ZN(n9018) );
  NOR2_X1 U10369 ( .A1(n9023), .A2(n4808), .ZN(n9066) );
  NAND2_X1 U10370 ( .A1(n9066), .A2(n9072), .ZN(n9065) );
  NAND2_X1 U10371 ( .A1(n9065), .A2(n9024), .ZN(n9026) );
  XNOR2_X1 U10372 ( .A(n9026), .B(n9025), .ZN(n9232) );
  INV_X1 U10373 ( .A(n9232), .ZN(n9064) );
  NAND2_X1 U10374 ( .A1(n9221), .A2(n9220), .ZN(n9031) );
  NAND2_X1 U10375 ( .A1(n9036), .A2(n9035), .ZN(n9158) );
  NAND2_X1 U10376 ( .A1(n9158), .A2(n9037), .ZN(n9039) );
  NAND2_X1 U10377 ( .A1(n9039), .A2(n9038), .ZN(n9137) );
  INV_X1 U10378 ( .A(n9119), .ZN(n9040) );
  NOR2_X1 U10379 ( .A1(n9130), .A2(n9040), .ZN(n9041) );
  NAND2_X1 U10380 ( .A1(n9120), .A2(n9041), .ZN(n9121) );
  INV_X1 U10381 ( .A(n9048), .ZN(n9049) );
  XNOR2_X1 U10382 ( .A(n9052), .B(n9051), .ZN(n9053) );
  OAI222_X1 U10383 ( .A1(n9055), .A2(n9054), .B1(n9608), .B2(n9084), .C1(n9591), .C2(n9053), .ZN(n9233) );
  INV_X1 U10384 ( .A(n9235), .ZN(n9061) );
  AOI211_X1 U10385 ( .C1(n9235), .C2(n4300), .A(n9680), .B(n9056), .ZN(n9234)
         );
  NAND2_X1 U10386 ( .A1(n9234), .A2(n9209), .ZN(n9060) );
  INV_X1 U10387 ( .A(n9057), .ZN(n9058) );
  AOI22_X1 U10388 ( .A1(n9058), .A2(n9586), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9598), .ZN(n9059) );
  OAI211_X1 U10389 ( .C1(n9061), .C2(n9619), .A(n9060), .B(n9059), .ZN(n9062)
         );
  AOI21_X1 U10390 ( .B1(n9233), .B2(n9617), .A(n9062), .ZN(n9063) );
  OAI21_X1 U10391 ( .B1(n9064), .B2(n9228), .A(n9063), .ZN(P1_U3355) );
  NAND2_X1 U10392 ( .A1(n9086), .A2(n9238), .ZN(n9067) );
  NAND2_X1 U10393 ( .A1(n9238), .A2(n9132), .ZN(n9069) );
  NAND2_X1 U10394 ( .A1(n9598), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9068) );
  OAI211_X1 U10395 ( .C1(n9618), .C2(n9070), .A(n9069), .B(n9068), .ZN(n9071)
         );
  AOI21_X1 U10396 ( .B1(n9239), .B2(n9603), .A(n9071), .ZN(n9079) );
  XNOR2_X1 U10397 ( .A(n9073), .B(n9072), .ZN(n9077) );
  OAI22_X1 U10398 ( .A1(n9075), .A2(n9608), .B1(n9074), .B2(n9610), .ZN(n9076)
         );
  OR2_X1 U10399 ( .A1(n9241), .A2(n9598), .ZN(n9078) );
  OAI211_X1 U10400 ( .C1(n9242), .C2(n9228), .A(n9079), .B(n9078), .ZN(
        P1_U3263) );
  XNOR2_X1 U10401 ( .A(n9080), .B(n9082), .ZN(n9247) );
  XNOR2_X1 U10402 ( .A(n9081), .B(n9082), .ZN(n9083) );
  OAI222_X1 U10403 ( .A1(n9608), .A2(n9085), .B1(n9610), .B2(n9084), .C1(n9083), .C2(n9591), .ZN(n9243) );
  INV_X1 U10404 ( .A(n9094), .ZN(n9087) );
  AOI211_X1 U10405 ( .C1(n9245), .C2(n9087), .A(n9680), .B(n4481), .ZN(n9244)
         );
  NAND2_X1 U10406 ( .A1(n9244), .A2(n9209), .ZN(n9090) );
  AOI22_X1 U10407 ( .A1(n9088), .A2(n9586), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9598), .ZN(n9089) );
  OAI211_X1 U10408 ( .C1(n9091), .C2(n9619), .A(n9090), .B(n9089), .ZN(n9092)
         );
  AOI21_X1 U10409 ( .B1(n9243), .B2(n9617), .A(n9092), .ZN(n9093) );
  OAI21_X1 U10410 ( .B1(n9247), .B2(n9228), .A(n9093), .ZN(P1_U3264) );
  XOR2_X1 U10411 ( .A(n9100), .B(n4328), .Z(n9252) );
  INV_X1 U10412 ( .A(n9108), .ZN(n9095) );
  AOI21_X1 U10413 ( .B1(n9248), .B2(n9095), .A(n9094), .ZN(n9249) );
  AOI22_X1 U10414 ( .A1(n9096), .A2(n9586), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9598), .ZN(n9097) );
  OAI21_X1 U10415 ( .B1(n9098), .B2(n9619), .A(n9097), .ZN(n9104) );
  XOR2_X1 U10416 ( .A(n9100), .B(n9099), .Z(n9102) );
  AOI222_X1 U10417 ( .A1(n9612), .A2(n9102), .B1(n9101), .B2(n9357), .C1(n9018), .C2(n9359), .ZN(n9251) );
  NOR2_X1 U10418 ( .A1(n9251), .A2(n9598), .ZN(n9103) );
  AOI211_X1 U10419 ( .C1(n9603), .C2(n9249), .A(n9104), .B(n9103), .ZN(n9105)
         );
  OAI21_X1 U10420 ( .B1(n9252), .B2(n9228), .A(n9105), .ZN(P1_U3265) );
  AOI21_X1 U10421 ( .B1(n9113), .B2(n4273), .A(n9106), .ZN(n9257) );
  AOI21_X1 U10422 ( .B1(n9253), .B2(n9125), .A(n9108), .ZN(n9254) );
  INV_X1 U10423 ( .A(n9109), .ZN(n9110) );
  AOI22_X1 U10424 ( .A1(n9110), .A2(n9586), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9598), .ZN(n9111) );
  OAI21_X1 U10425 ( .B1(n4485), .B2(n9619), .A(n9111), .ZN(n9117) );
  XNOR2_X1 U10426 ( .A(n9112), .B(n9113), .ZN(n9115) );
  AOI222_X1 U10427 ( .A1(n9612), .A2(n9115), .B1(n9114), .B2(n9357), .C1(n9015), .C2(n9359), .ZN(n9256) );
  NOR2_X1 U10428 ( .A1(n9256), .A2(n9598), .ZN(n9116) );
  AOI211_X1 U10429 ( .C1(n9254), .C2(n9603), .A(n9117), .B(n9116), .ZN(n9118)
         );
  OAI21_X1 U10430 ( .B1(n9257), .B2(n9228), .A(n9118), .ZN(P1_U3266) );
  AND2_X1 U10431 ( .A1(n9120), .A2(n9119), .ZN(n9123) );
  OAI21_X1 U10432 ( .B1(n9123), .B2(n9122), .A(n9121), .ZN(n9124) );
  AOI222_X1 U10433 ( .A1(n9612), .A2(n9124), .B1(n9018), .B2(n9357), .C1(n9160), .C2(n9359), .ZN(n9263) );
  INV_X1 U10434 ( .A(n9125), .ZN(n9126) );
  AOI211_X1 U10435 ( .C1(n9261), .C2(n9142), .A(n9680), .B(n9126), .ZN(n9260)
         );
  AOI22_X1 U10436 ( .A1(n9260), .A2(n9128), .B1(n9586), .B2(n9127), .ZN(n9129)
         );
  AND2_X1 U10437 ( .A1(n9263), .A2(n9129), .ZN(n9135) );
  OR2_X1 U10438 ( .A1(n9131), .A2(n9130), .ZN(n9259) );
  NAND3_X1 U10439 ( .A1(n9259), .A2(n9258), .A3(n9171), .ZN(n9134) );
  AOI22_X1 U10440 ( .A1(n9261), .A2(n9132), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9598), .ZN(n9133) );
  OAI211_X1 U10441 ( .C1(n9598), .C2(n9135), .A(n9134), .B(n9133), .ZN(
        P1_U3267) );
  XOR2_X1 U10442 ( .A(n9136), .B(n9138), .Z(n9269) );
  XNOR2_X1 U10443 ( .A(n9137), .B(n9138), .ZN(n9139) );
  OAI222_X1 U10444 ( .A1(n9608), .A2(n9141), .B1(n9610), .B2(n9140), .C1(n9139), .C2(n9591), .ZN(n9265) );
  INV_X1 U10445 ( .A(n9153), .ZN(n9144) );
  INV_X1 U10446 ( .A(n9142), .ZN(n9143) );
  AOI211_X1 U10447 ( .C1(n9267), .C2(n9144), .A(n9680), .B(n9143), .ZN(n9266)
         );
  NAND2_X1 U10448 ( .A1(n9266), .A2(n9209), .ZN(n9148) );
  INV_X1 U10449 ( .A(n9145), .ZN(n9146) );
  AOI22_X1 U10450 ( .A1(n9146), .A2(n9586), .B1(n9598), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9147) );
  OAI211_X1 U10451 ( .C1(n9149), .C2(n9619), .A(n9148), .B(n9147), .ZN(n9150)
         );
  AOI21_X1 U10452 ( .B1(n9265), .B2(n9617), .A(n9150), .ZN(n9151) );
  OAI21_X1 U10453 ( .B1(n9269), .B2(n9228), .A(n9151), .ZN(P1_U3268) );
  XNOR2_X1 U10454 ( .A(n9152), .B(n9159), .ZN(n9274) );
  AOI21_X1 U10455 ( .B1(n9270), .B2(n9172), .A(n9153), .ZN(n9271) );
  INV_X1 U10456 ( .A(n9154), .ZN(n9155) );
  AOI22_X1 U10457 ( .A1(n9598), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9155), .B2(
        n9586), .ZN(n9156) );
  OAI21_X1 U10458 ( .B1(n9157), .B2(n9619), .A(n9156), .ZN(n9164) );
  XOR2_X1 U10459 ( .A(n9159), .B(n9158), .Z(n9162) );
  AOI222_X1 U10460 ( .A1(n9612), .A2(n9162), .B1(n9161), .B2(n9359), .C1(n9160), .C2(n9357), .ZN(n9273) );
  NOR2_X1 U10461 ( .A1(n9273), .A2(n9598), .ZN(n9163) );
  AOI211_X1 U10462 ( .C1(n9271), .C2(n9603), .A(n9164), .B(n9163), .ZN(n9165)
         );
  OAI21_X1 U10463 ( .B1(n9274), .B2(n9228), .A(n9165), .ZN(P1_U3269) );
  XNOR2_X1 U10464 ( .A(n9166), .B(n9169), .ZN(n9168) );
  AOI222_X1 U10465 ( .A1(n9612), .A2(n9168), .B1(n9167), .B2(n9357), .C1(n9204), .C2(n9359), .ZN(n9280) );
  OR2_X1 U10466 ( .A1(n9170), .A2(n9169), .ZN(n9276) );
  NAND3_X1 U10467 ( .A1(n9276), .A2(n9275), .A3(n9171), .ZN(n9179) );
  INV_X1 U10468 ( .A(n9172), .ZN(n9173) );
  AOI21_X1 U10469 ( .B1(n9277), .B2(n9186), .A(n9173), .ZN(n9278) );
  AOI22_X1 U10470 ( .A1(n9598), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9174), .B2(
        n9586), .ZN(n9175) );
  OAI21_X1 U10471 ( .B1(n9176), .B2(n9619), .A(n9175), .ZN(n9177) );
  AOI21_X1 U10472 ( .B1(n9278), .B2(n9603), .A(n9177), .ZN(n9178) );
  OAI211_X1 U10473 ( .C1(n9598), .C2(n9280), .A(n9179), .B(n9178), .ZN(
        P1_U3270) );
  XOR2_X1 U10474 ( .A(n9180), .B(n9182), .Z(n9286) );
  XOR2_X1 U10475 ( .A(n9182), .B(n9181), .Z(n9183) );
  OAI222_X1 U10476 ( .A1(n9608), .A2(n9185), .B1(n9610), .B2(n9184), .C1(n9183), .C2(n9591), .ZN(n9282) );
  AOI211_X1 U10477 ( .C1(n9284), .C2(n9195), .A(n9680), .B(n4476), .ZN(n9283)
         );
  NAND2_X1 U10478 ( .A1(n9283), .A2(n9209), .ZN(n9190) );
  INV_X1 U10479 ( .A(n9187), .ZN(n9188) );
  AOI22_X1 U10480 ( .A1(n9598), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9188), .B2(
        n9586), .ZN(n9189) );
  OAI211_X1 U10481 ( .C1(n9191), .C2(n9619), .A(n9190), .B(n9189), .ZN(n9192)
         );
  AOI21_X1 U10482 ( .B1(n9282), .B2(n9617), .A(n9192), .ZN(n9193) );
  OAI21_X1 U10483 ( .B1(n9286), .B2(n9228), .A(n9193), .ZN(P1_U3271) );
  XNOR2_X1 U10484 ( .A(n9194), .B(n9203), .ZN(n9291) );
  INV_X1 U10485 ( .A(n9214), .ZN(n9196) );
  AOI211_X1 U10486 ( .C1(n9288), .C2(n9196), .A(n9680), .B(n4477), .ZN(n9287)
         );
  INV_X1 U10487 ( .A(n9197), .ZN(n9198) );
  AOI22_X1 U10488 ( .A1(n9598), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9198), .B2(
        n9586), .ZN(n9199) );
  OAI21_X1 U10489 ( .B1(n9200), .B2(n9619), .A(n9199), .ZN(n9208) );
  OAI21_X1 U10490 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n9206) );
  AOI222_X1 U10491 ( .A1(n9612), .A2(n9206), .B1(n9205), .B2(n9359), .C1(n9204), .C2(n9357), .ZN(n9290) );
  NOR2_X1 U10492 ( .A1(n9290), .A2(n9598), .ZN(n9207) );
  AOI211_X1 U10493 ( .C1(n9287), .C2(n9209), .A(n9208), .B(n9207), .ZN(n9210)
         );
  OAI21_X1 U10494 ( .B1(n9291), .B2(n9228), .A(n9210), .ZN(P1_U3272) );
  XNOR2_X1 U10495 ( .A(n9212), .B(n9211), .ZN(n9296) );
  INV_X1 U10496 ( .A(n9213), .ZN(n9215) );
  AOI21_X1 U10497 ( .B1(n9292), .B2(n9215), .A(n9214), .ZN(n9293) );
  INV_X1 U10498 ( .A(n9216), .ZN(n9217) );
  AOI22_X1 U10499 ( .A1(n9598), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9217), .B2(
        n9586), .ZN(n9218) );
  OAI21_X1 U10500 ( .B1(n9219), .B2(n9619), .A(n9218), .ZN(n9226) );
  XNOR2_X1 U10501 ( .A(n9221), .B(n9220), .ZN(n9224) );
  AOI222_X1 U10502 ( .A1(n9612), .A2(n9224), .B1(n9223), .B2(n9359), .C1(n9222), .C2(n9357), .ZN(n9295) );
  NOR2_X1 U10503 ( .A1(n9295), .A2(n9598), .ZN(n9225) );
  AOI211_X1 U10504 ( .C1(n9293), .C2(n9603), .A(n9226), .B(n9225), .ZN(n9227)
         );
  OAI21_X1 U10505 ( .B1(n9296), .B2(n9228), .A(n9227), .ZN(P1_U3273) );
  AOI21_X1 U10506 ( .B1(n9229), .B2(n9632), .A(n9372), .ZN(n9230) );
  OAI21_X1 U10507 ( .B1(n9231), .B2(n9680), .A(n9230), .ZN(n9302) );
  MUX2_X1 U10508 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9302), .S(n4269), .Z(
        P1_U3554) );
  NAND2_X1 U10509 ( .A1(n9232), .A2(n9684), .ZN(n9237) );
  AOI211_X1 U10510 ( .C1(n9632), .C2(n9235), .A(n9234), .B(n9233), .ZN(n9236)
         );
  NAND2_X1 U10511 ( .A1(n9237), .A2(n9236), .ZN(n9303) );
  MUX2_X1 U10512 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9303), .S(n4269), .Z(
        P1_U3552) );
  AOI22_X1 U10513 ( .A1(n9239), .A2(n9633), .B1(n9632), .B2(n9238), .ZN(n9240)
         );
  OAI211_X1 U10514 ( .C1(n9242), .C2(n9375), .A(n9241), .B(n9240), .ZN(n9304)
         );
  MUX2_X1 U10515 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9304), .S(n4269), .Z(
        P1_U3551) );
  AOI211_X1 U10516 ( .C1(n9632), .C2(n9245), .A(n9244), .B(n9243), .ZN(n9246)
         );
  OAI21_X1 U10517 ( .B1(n9247), .B2(n9375), .A(n9246), .ZN(n9305) );
  MUX2_X1 U10518 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9305), .S(n4269), .Z(
        P1_U3550) );
  AOI22_X1 U10519 ( .A1(n9249), .A2(n9633), .B1(n9632), .B2(n9248), .ZN(n9250)
         );
  OAI211_X1 U10520 ( .C1(n9252), .C2(n9375), .A(n9251), .B(n9250), .ZN(n9306)
         );
  MUX2_X1 U10521 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9306), .S(n4269), .Z(
        P1_U3549) );
  AOI22_X1 U10522 ( .A1(n9254), .A2(n9633), .B1(n9632), .B2(n9253), .ZN(n9255)
         );
  OAI211_X1 U10523 ( .C1(n9257), .C2(n9375), .A(n9256), .B(n9255), .ZN(n9307)
         );
  MUX2_X1 U10524 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9307), .S(n4269), .Z(
        P1_U3548) );
  NAND3_X1 U10525 ( .A1(n9259), .A2(n9258), .A3(n9684), .ZN(n9264) );
  AOI21_X1 U10526 ( .B1(n9632), .B2(n9261), .A(n9260), .ZN(n9262) );
  NAND3_X1 U10527 ( .A1(n9264), .A2(n9263), .A3(n9262), .ZN(n9308) );
  MUX2_X1 U10528 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9308), .S(n4269), .Z(
        P1_U3547) );
  AOI211_X1 U10529 ( .C1(n9632), .C2(n9267), .A(n9266), .B(n9265), .ZN(n9268)
         );
  OAI21_X1 U10530 ( .B1(n9269), .B2(n9375), .A(n9268), .ZN(n9309) );
  MUX2_X1 U10531 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9309), .S(n4269), .Z(
        P1_U3546) );
  AOI22_X1 U10532 ( .A1(n9271), .A2(n9633), .B1(n9632), .B2(n9270), .ZN(n9272)
         );
  OAI211_X1 U10533 ( .C1(n9274), .C2(n9375), .A(n9273), .B(n9272), .ZN(n9310)
         );
  MUX2_X1 U10534 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9310), .S(n4269), .Z(
        P1_U3545) );
  NAND3_X1 U10535 ( .A1(n9276), .A2(n9275), .A3(n9684), .ZN(n9281) );
  AOI22_X1 U10536 ( .A1(n9278), .A2(n9633), .B1(n9632), .B2(n9277), .ZN(n9279)
         );
  NAND3_X1 U10537 ( .A1(n9281), .A2(n9280), .A3(n9279), .ZN(n9311) );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9311), .S(n4269), .Z(
        P1_U3544) );
  AOI211_X1 U10539 ( .C1(n9632), .C2(n9284), .A(n9283), .B(n9282), .ZN(n9285)
         );
  OAI21_X1 U10540 ( .B1(n9286), .B2(n9375), .A(n9285), .ZN(n9312) );
  MUX2_X1 U10541 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9312), .S(n4269), .Z(
        P1_U3543) );
  AOI21_X1 U10542 ( .B1(n9632), .B2(n9288), .A(n9287), .ZN(n9289) );
  OAI211_X1 U10543 ( .C1(n9291), .C2(n9375), .A(n9290), .B(n9289), .ZN(n9313)
         );
  MUX2_X1 U10544 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9313), .S(n4269), .Z(
        P1_U3542) );
  AOI22_X1 U10545 ( .A1(n9293), .A2(n9633), .B1(n9632), .B2(n9292), .ZN(n9294)
         );
  OAI211_X1 U10546 ( .C1(n9296), .C2(n9375), .A(n9295), .B(n9294), .ZN(n9314)
         );
  MUX2_X1 U10547 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9314), .S(n4269), .Z(
        P1_U3541) );
  AOI211_X1 U10548 ( .C1(n9632), .C2(n9299), .A(n9298), .B(n9297), .ZN(n9300)
         );
  OAI21_X1 U10549 ( .B1(n9301), .B2(n9375), .A(n9300), .ZN(n9315) );
  MUX2_X1 U10550 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9315), .S(n4269), .Z(
        P1_U3540) );
  MUX2_X1 U10551 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9302), .S(n10017), .Z(
        P1_U3522) );
  MUX2_X1 U10552 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9303), .S(n10017), .Z(
        P1_U3520) );
  MUX2_X1 U10553 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9304), .S(n10017), .Z(
        P1_U3519) );
  MUX2_X1 U10554 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9305), .S(n10017), .Z(
        P1_U3518) );
  MUX2_X1 U10555 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9306), .S(n10017), .Z(
        P1_U3517) );
  MUX2_X1 U10556 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9307), .S(n10017), .Z(
        P1_U3516) );
  MUX2_X1 U10557 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9308), .S(n10017), .Z(
        P1_U3515) );
  MUX2_X1 U10558 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9309), .S(n10017), .Z(
        P1_U3514) );
  MUX2_X1 U10559 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9310), .S(n10017), .Z(
        P1_U3513) );
  MUX2_X1 U10560 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9311), .S(n10017), .Z(
        P1_U3512) );
  MUX2_X1 U10561 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9312), .S(n10017), .Z(
        P1_U3511) );
  MUX2_X1 U10562 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9313), .S(n10017), .Z(
        P1_U3510) );
  MUX2_X1 U10563 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9314), .S(n10017), .Z(
        P1_U3508) );
  MUX2_X1 U10564 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9315), .S(n10017), .Z(
        P1_U3505) );
  NAND3_X1 U10565 ( .A1(n4487), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9316) );
  OAI22_X1 U10566 ( .A1(n5030), .A2(n9316), .B1(n4993), .B2(n9328), .ZN(n9317)
         );
  AOI21_X1 U10567 ( .B1(n8743), .B2(n9323), .A(n9317), .ZN(n9318) );
  INV_X1 U10568 ( .A(n9318), .ZN(P1_U3322) );
  OAI222_X1 U10569 ( .A1(n9328), .A2(n9322), .B1(n9319), .B2(P1_U3084), .C1(
        n8059), .C2(n9320), .ZN(P1_U3324) );
  NAND2_X1 U10570 ( .A1(n9324), .A2(n9323), .ZN(n9326) );
  OAI211_X1 U10571 ( .C1(n9328), .C2(n9327), .A(n9326), .B(n9325), .ZN(
        P1_U3325) );
  MUX2_X1 U10572 ( .A(n9329), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U10573 ( .A1(n9452), .A2(n9330), .ZN(n9331) );
  AOI211_X1 U10574 ( .C1(n9432), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9332), .B(
        n9331), .ZN(n9341) );
  OAI211_X1 U10575 ( .C1(n9335), .C2(n9334), .A(n9557), .B(n9333), .ZN(n9340)
         );
  OAI211_X1 U10576 ( .C1(n9338), .C2(n9337), .A(n9454), .B(n9336), .ZN(n9339)
         );
  NAND3_X1 U10577 ( .A1(n9341), .A2(n9340), .A3(n9339), .ZN(P1_U3244) );
  OAI21_X1 U10578 ( .B1(n9343), .B2(n9820), .A(n9342), .ZN(n9344) );
  AOI21_X1 U10579 ( .B1(n9345), .B2(n9810), .A(n9344), .ZN(n9347) );
  INV_X1 U10580 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U10581 ( .A1(n4268), .A2(n9347), .B1(n9994), .B2(n9833), .ZN(
        P2_U3550) );
  INV_X1 U10582 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9346) );
  AOI22_X1 U10583 ( .A1(n4267), .A2(n9347), .B1(n9346), .B2(n9825), .ZN(
        P2_U3518) );
  XNOR2_X1 U10584 ( .A(n9349), .B(n9348), .ZN(n9411) );
  OR2_X1 U10585 ( .A1(n9350), .A2(n9408), .ZN(n9351) );
  NAND2_X1 U10586 ( .A1(n9352), .A2(n9351), .ZN(n9409) );
  INV_X1 U10587 ( .A(n9409), .ZN(n9353) );
  AOI22_X1 U10588 ( .A1(n9411), .A2(n9604), .B1(n9603), .B2(n9353), .ZN(n9369)
         );
  XNOR2_X1 U10589 ( .A(n9354), .B(n9355), .ZN(n9361) );
  AOI22_X1 U10590 ( .A1(n9359), .A2(n9358), .B1(n9357), .B2(n9356), .ZN(n9360)
         );
  OAI21_X1 U10591 ( .B1(n9361), .B2(n9591), .A(n9360), .ZN(n9362) );
  AOI21_X1 U10592 ( .B1(n9411), .B2(n9363), .A(n9362), .ZN(n9413) );
  INV_X1 U10593 ( .A(n9413), .ZN(n9367) );
  AOI22_X1 U10594 ( .A1(n9598), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9364), .B2(
        n9586), .ZN(n9365) );
  OAI21_X1 U10595 ( .B1(n9408), .B2(n9619), .A(n9365), .ZN(n9366) );
  AOI21_X1 U10596 ( .B1(n9367), .B2(n9617), .A(n9366), .ZN(n9368) );
  NAND2_X1 U10597 ( .A1(n9369), .A2(n9368), .ZN(P1_U3280) );
  INV_X1 U10598 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9374) );
  AOI22_X1 U10599 ( .A1(n4269), .A2(n9416), .B1(n9374), .B2(n9697), .ZN(
        P1_U3553) );
  NOR3_X1 U10600 ( .A1(n4337), .A2(n9376), .A3(n9375), .ZN(n9381) );
  NOR2_X1 U10601 ( .A1(n9377), .A2(n9678), .ZN(n9379) );
  NOR4_X1 U10602 ( .A1(n9381), .A2(n9380), .A3(n9379), .A4(n9378), .ZN(n9418)
         );
  AOI22_X1 U10603 ( .A1(n4269), .A2(n9418), .B1(n9382), .B2(n9697), .ZN(
        P1_U3539) );
  OAI22_X1 U10604 ( .A1(n9384), .A2(n9680), .B1(n9383), .B2(n9678), .ZN(n9386)
         );
  AOI211_X1 U10605 ( .C1(n9684), .C2(n9387), .A(n9386), .B(n9385), .ZN(n9420)
         );
  INV_X1 U10606 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9388) );
  AOI22_X1 U10607 ( .A1(n4269), .A2(n9420), .B1(n9388), .B2(n9697), .ZN(
        P1_U3538) );
  OAI211_X1 U10608 ( .C1(n9391), .C2(n9678), .A(n9390), .B(n9389), .ZN(n9392)
         );
  AOI21_X1 U10609 ( .B1(n9393), .B2(n9684), .A(n9392), .ZN(n9422) );
  AOI22_X1 U10610 ( .A1(n4269), .A2(n9422), .B1(n9394), .B2(n9697), .ZN(
        P1_U3537) );
  INV_X1 U10611 ( .A(n9638), .ZN(n9677) );
  OAI21_X1 U10612 ( .B1(n9396), .B2(n9678), .A(n9395), .ZN(n9397) );
  AOI21_X1 U10613 ( .B1(n9398), .B2(n9677), .A(n9397), .ZN(n9399) );
  AND2_X1 U10614 ( .A1(n9400), .A2(n9399), .ZN(n9424) );
  AOI22_X1 U10615 ( .A1(n4269), .A2(n9424), .B1(n9401), .B2(n9697), .ZN(
        P1_U3536) );
  OAI21_X1 U10616 ( .B1(n4475), .B2(n9678), .A(n9402), .ZN(n9403) );
  AOI21_X1 U10617 ( .B1(n9404), .B2(n9677), .A(n9403), .ZN(n9405) );
  AND2_X1 U10618 ( .A1(n9406), .A2(n9405), .ZN(n9426) );
  AOI22_X1 U10619 ( .A1(n4269), .A2(n9426), .B1(n9407), .B2(n9697), .ZN(
        P1_U3535) );
  OAI22_X1 U10620 ( .A1(n9409), .A2(n9680), .B1(n9408), .B2(n9678), .ZN(n9410)
         );
  AOI21_X1 U10621 ( .B1(n9411), .B2(n9677), .A(n9410), .ZN(n9412) );
  AND2_X1 U10622 ( .A1(n9413), .A2(n9412), .ZN(n9428) );
  AOI22_X1 U10623 ( .A1(n4269), .A2(n9428), .B1(n9414), .B2(n9697), .ZN(
        P1_U3534) );
  INV_X1 U10624 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9415) );
  AOI22_X1 U10625 ( .A1(n10017), .A2(n9416), .B1(n9415), .B2(n9686), .ZN(
        P1_U3521) );
  INV_X1 U10626 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9417) );
  AOI22_X1 U10627 ( .A1(n10017), .A2(n9418), .B1(n9417), .B2(n9686), .ZN(
        P1_U3502) );
  INV_X1 U10628 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9419) );
  AOI22_X1 U10629 ( .A1(n10017), .A2(n9420), .B1(n9419), .B2(n9686), .ZN(
        P1_U3499) );
  INV_X1 U10630 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9421) );
  AOI22_X1 U10631 ( .A1(n10017), .A2(n9422), .B1(n9421), .B2(n9686), .ZN(
        P1_U3496) );
  INV_X1 U10632 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9423) );
  AOI22_X1 U10633 ( .A1(n10017), .A2(n9424), .B1(n9423), .B2(n9686), .ZN(
        P1_U3493) );
  INV_X1 U10634 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9425) );
  AOI22_X1 U10635 ( .A1(n10017), .A2(n9426), .B1(n9425), .B2(n9686), .ZN(
        P1_U3490) );
  INV_X1 U10636 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9427) );
  AOI22_X1 U10637 ( .A1(n10017), .A2(n9428), .B1(n9427), .B2(n9686), .ZN(
        P1_U3487) );
  XNOR2_X1 U10638 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10639 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI22_X1 U10640 ( .A1(n9452), .A2(n9430), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9429), .ZN(n9431) );
  AOI21_X1 U10641 ( .B1(n9432), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n9431), .ZN(
        n9446) );
  INV_X1 U10642 ( .A(n9433), .ZN(n9437) );
  OAI21_X1 U10643 ( .B1(n9435), .B2(n9440), .A(n9434), .ZN(n9436) );
  NAND3_X1 U10644 ( .A1(n9454), .A2(n9437), .A3(n9436), .ZN(n9445) );
  INV_X1 U10645 ( .A(n9438), .ZN(n9443) );
  OAI21_X1 U10646 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(n9442) );
  NAND3_X1 U10647 ( .A1(n9557), .A2(n9443), .A3(n9442), .ZN(n9444) );
  NAND3_X1 U10648 ( .A1(n9446), .A2(n9445), .A3(n9444), .ZN(P1_U3242) );
  INV_X1 U10649 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9461) );
  XNOR2_X1 U10650 ( .A(n9447), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n9448) );
  XNOR2_X1 U10651 ( .A(n9449), .B(n9448), .ZN(n9455) );
  OAI21_X1 U10652 ( .B1(n9452), .B2(n9451), .A(n9450), .ZN(n9453) );
  AOI21_X1 U10653 ( .B1(n9455), .B2(n9454), .A(n9453), .ZN(n9460) );
  OAI211_X1 U10654 ( .C1(n9458), .C2(n9457), .A(n9557), .B(n9456), .ZN(n9459)
         );
  OAI211_X1 U10655 ( .C1(n9461), .C2(n9579), .A(n9460), .B(n9459), .ZN(
        P1_U3249) );
  AOI211_X1 U10656 ( .C1(n9464), .C2(n9463), .A(n9564), .B(n9462), .ZN(n9465)
         );
  AOI211_X1 U10657 ( .C1(n9570), .C2(n9467), .A(n9466), .B(n9465), .ZN(n9473)
         );
  AOI21_X1 U10658 ( .B1(n9470), .B2(n9469), .A(n9468), .ZN(n9471) );
  OR2_X1 U10659 ( .A1(n9471), .A2(n9576), .ZN(n9472) );
  OAI211_X1 U10660 ( .C1(n10030), .C2(n9579), .A(n9473), .B(n9472), .ZN(
        P1_U3250) );
  INV_X1 U10661 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9487) );
  AOI211_X1 U10662 ( .C1(n9476), .C2(n9475), .A(n9564), .B(n9474), .ZN(n9477)
         );
  AOI211_X1 U10663 ( .C1(n9570), .C2(n9479), .A(n9478), .B(n9477), .ZN(n9486)
         );
  INV_X1 U10664 ( .A(n9480), .ZN(n9481) );
  AOI21_X1 U10665 ( .B1(n9483), .B2(n9482), .A(n9481), .ZN(n9484) );
  OR2_X1 U10666 ( .A1(n9484), .A2(n9576), .ZN(n9485) );
  OAI211_X1 U10667 ( .C1(n9487), .C2(n9579), .A(n9486), .B(n9485), .ZN(
        P1_U3251) );
  INV_X1 U10668 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9500) );
  AOI211_X1 U10669 ( .C1(n9490), .C2(n9489), .A(n9488), .B(n9564), .ZN(n9491)
         );
  AOI211_X1 U10670 ( .C1(n9570), .C2(n9493), .A(n9492), .B(n9491), .ZN(n9499)
         );
  AOI21_X1 U10671 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9497) );
  OR2_X1 U10672 ( .A1(n9576), .A2(n9497), .ZN(n9498) );
  OAI211_X1 U10673 ( .C1(n9500), .C2(n9579), .A(n9499), .B(n9498), .ZN(
        P1_U3253) );
  INV_X1 U10674 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9513) );
  AOI211_X1 U10675 ( .C1(n9503), .C2(n9502), .A(n9501), .B(n9564), .ZN(n9504)
         );
  AOI211_X1 U10676 ( .C1(n9570), .C2(n9506), .A(n9505), .B(n9504), .ZN(n9512)
         );
  AOI21_X1 U10677 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(n9510) );
  OR2_X1 U10678 ( .A1(n9576), .A2(n9510), .ZN(n9511) );
  OAI211_X1 U10679 ( .C1(n9513), .C2(n9579), .A(n9512), .B(n9511), .ZN(
        P1_U3254) );
  INV_X1 U10680 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9907) );
  AOI211_X1 U10681 ( .C1(n9516), .C2(n9515), .A(n9514), .B(n9564), .ZN(n9517)
         );
  AOI211_X1 U10682 ( .C1(n9570), .C2(n9519), .A(n9518), .B(n9517), .ZN(n9525)
         );
  AOI21_X1 U10683 ( .B1(n9522), .B2(n9521), .A(n9520), .ZN(n9523) );
  OR2_X1 U10684 ( .A1(n9576), .A2(n9523), .ZN(n9524) );
  OAI211_X1 U10685 ( .C1(n9907), .C2(n9579), .A(n9525), .B(n9524), .ZN(
        P1_U3255) );
  INV_X1 U10686 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9987) );
  INV_X1 U10687 ( .A(n9526), .ZN(n9531) );
  AOI211_X1 U10688 ( .C1(n9529), .C2(n9528), .A(n9564), .B(n9527), .ZN(n9530)
         );
  AOI211_X1 U10689 ( .C1(n9570), .C2(n9532), .A(n9531), .B(n9530), .ZN(n9536)
         );
  XOR2_X1 U10690 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9533), .Z(n9534) );
  NAND2_X1 U10691 ( .A1(n9557), .A2(n9534), .ZN(n9535) );
  OAI211_X1 U10692 ( .C1(n9987), .C2(n9579), .A(n9536), .B(n9535), .ZN(
        P1_U3256) );
  INV_X1 U10693 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9549) );
  INV_X1 U10694 ( .A(n9537), .ZN(n9542) );
  AOI211_X1 U10695 ( .C1(n9540), .C2(n9539), .A(n9538), .B(n9564), .ZN(n9541)
         );
  AOI211_X1 U10696 ( .C1(n9570), .C2(n9543), .A(n9542), .B(n9541), .ZN(n9548)
         );
  OAI211_X1 U10697 ( .C1(n9546), .C2(n9545), .A(n9557), .B(n9544), .ZN(n9547)
         );
  OAI211_X1 U10698 ( .C1(n9549), .C2(n9579), .A(n9548), .B(n9547), .ZN(
        P1_U3257) );
  INV_X1 U10699 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9562) );
  AOI211_X1 U10700 ( .C1(n9552), .C2(n9551), .A(n9550), .B(n9564), .ZN(n9553)
         );
  AOI211_X1 U10701 ( .C1(n9570), .C2(n9555), .A(n9554), .B(n9553), .ZN(n9561)
         );
  OAI211_X1 U10702 ( .C1(n9559), .C2(n9558), .A(n9557), .B(n9556), .ZN(n9560)
         );
  OAI211_X1 U10703 ( .C1(n9562), .C2(n9579), .A(n9561), .B(n9560), .ZN(
        P1_U3258) );
  INV_X1 U10704 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9979) );
  INV_X1 U10705 ( .A(n9563), .ZN(n9569) );
  AOI211_X1 U10706 ( .C1(n9567), .C2(n9566), .A(n9565), .B(n9564), .ZN(n9568)
         );
  AOI211_X1 U10707 ( .C1(n9571), .C2(n9570), .A(n9569), .B(n9568), .ZN(n9578)
         );
  AOI21_X1 U10708 ( .B1(n9574), .B2(n9573), .A(n9572), .ZN(n9575) );
  OR2_X1 U10709 ( .A1(n9576), .A2(n9575), .ZN(n9577) );
  OAI211_X1 U10710 ( .C1(n9979), .C2(n9579), .A(n9578), .B(n9577), .ZN(
        P1_U3259) );
  XNOR2_X1 U10711 ( .A(n9580), .B(n9590), .ZN(n9658) );
  AOI21_X1 U10712 ( .B1(n9581), .B2(n9584), .A(n9680), .ZN(n9583) );
  NAND2_X1 U10713 ( .A1(n9583), .A2(n9582), .ZN(n9654) );
  AOI22_X1 U10714 ( .A1(n9586), .A2(n9585), .B1(n4349), .B2(n9584), .ZN(n9587)
         );
  OAI21_X1 U10715 ( .B1(n9654), .B2(n9588), .A(n9587), .ZN(n9594) );
  XNOR2_X1 U10716 ( .A(n9589), .B(n9590), .ZN(n9592) );
  OAI222_X1 U10717 ( .A1(n9608), .A2(n9609), .B1(n9610), .B2(n9593), .C1(n9592), .C2(n9591), .ZN(n9656) );
  AOI211_X1 U10718 ( .C1(n9595), .C2(n9658), .A(n9594), .B(n9656), .ZN(n9596)
         );
  AOI22_X1 U10719 ( .A1(n9598), .A2(n9597), .B1(n9596), .B2(n9617), .ZN(
        P1_U3286) );
  XNOR2_X1 U10720 ( .A(n9599), .B(n9607), .ZN(n9616) );
  INV_X1 U10721 ( .A(n9616), .ZN(n9645) );
  OAI21_X1 U10722 ( .B1(n9601), .B2(n9641), .A(n9600), .ZN(n9642) );
  INV_X1 U10723 ( .A(n9642), .ZN(n9602) );
  AOI22_X1 U10724 ( .A1(n9645), .A2(n9604), .B1(n9603), .B2(n9602), .ZN(n9623)
         );
  OAI21_X1 U10725 ( .B1(n9607), .B2(n9606), .A(n9605), .ZN(n9613) );
  OAI22_X1 U10726 ( .A1(n9610), .A2(n9609), .B1(n6023), .B2(n9608), .ZN(n9611)
         );
  AOI21_X1 U10727 ( .B1(n9613), .B2(n9612), .A(n9611), .ZN(n9614) );
  OAI21_X1 U10728 ( .B1(n9616), .B2(n9615), .A(n9614), .ZN(n9643) );
  MUX2_X1 U10729 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9643), .S(n9617), .Z(n9621)
         );
  OAI22_X1 U10730 ( .A1(n9619), .A2(n9641), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9618), .ZN(n9620) );
  NOR2_X1 U10731 ( .A1(n9621), .A2(n9620), .ZN(n9622) );
  NAND2_X1 U10732 ( .A1(n9623), .A2(n9622), .ZN(P1_U3288) );
  INV_X1 U10733 ( .A(n9624), .ZN(n9625) );
  AND2_X1 U10734 ( .A1(n9630), .A2(n9625), .ZN(n9626) );
  AND2_X1 U10735 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9627), .ZN(P1_U3292) );
  AND2_X1 U10736 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9627), .ZN(P1_U3293) );
  INV_X1 U10737 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9892) );
  NOR2_X1 U10738 ( .A1(n9626), .A2(n9892), .ZN(P1_U3294) );
  AND2_X1 U10739 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9627), .ZN(P1_U3295) );
  AND2_X1 U10740 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9627), .ZN(P1_U3296) );
  AND2_X1 U10741 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9627), .ZN(P1_U3297) );
  AND2_X1 U10742 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9627), .ZN(P1_U3298) );
  AND2_X1 U10743 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9627), .ZN(P1_U3299) );
  AND2_X1 U10744 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9627), .ZN(P1_U3300) );
  AND2_X1 U10745 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9627), .ZN(P1_U3301) );
  INV_X1 U10746 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9966) );
  NOR2_X1 U10747 ( .A1(n9626), .A2(n9966), .ZN(P1_U3302) );
  AND2_X1 U10748 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9627), .ZN(P1_U3303) );
  AND2_X1 U10749 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9627), .ZN(P1_U3304) );
  AND2_X1 U10750 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9627), .ZN(P1_U3305) );
  AND2_X1 U10751 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9627), .ZN(P1_U3306) );
  INV_X1 U10752 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9986) );
  NOR2_X1 U10753 ( .A1(n9626), .A2(n9986), .ZN(P1_U3307) );
  AND2_X1 U10754 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9627), .ZN(P1_U3308) );
  AND2_X1 U10755 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9627), .ZN(P1_U3309) );
  AND2_X1 U10756 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9627), .ZN(P1_U3310) );
  AND2_X1 U10757 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9627), .ZN(P1_U3311) );
  AND2_X1 U10758 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9627), .ZN(P1_U3312) );
  AND2_X1 U10759 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9627), .ZN(P1_U3313) );
  AND2_X1 U10760 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9627), .ZN(P1_U3314) );
  INV_X1 U10761 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9891) );
  NOR2_X1 U10762 ( .A1(n9626), .A2(n9891), .ZN(P1_U3315) );
  AND2_X1 U10763 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9627), .ZN(P1_U3316) );
  INV_X1 U10764 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9954) );
  NOR2_X1 U10765 ( .A1(n9626), .A2(n9954), .ZN(P1_U3317) );
  AND2_X1 U10766 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9627), .ZN(P1_U3318) );
  AND2_X1 U10767 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9627), .ZN(P1_U3319) );
  AND2_X1 U10768 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9627), .ZN(P1_U3320) );
  AND2_X1 U10769 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9627), .ZN(P1_U3321) );
  NAND2_X1 U10770 ( .A1(n9628), .A2(n9630), .ZN(n9629) );
  OAI21_X1 U10771 ( .B1(n9631), .B2(n9630), .A(n9629), .ZN(P1_U3440) );
  AOI22_X1 U10772 ( .A1(n9634), .A2(n9633), .B1(n9632), .B2(n6022), .ZN(n9635)
         );
  OAI211_X1 U10773 ( .C1(n9638), .C2(n9637), .A(n9636), .B(n9635), .ZN(n9639)
         );
  INV_X1 U10774 ( .A(n9639), .ZN(n9689) );
  INV_X1 U10775 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9640) );
  AOI22_X1 U10776 ( .A1(n10017), .A2(n9689), .B1(n9640), .B2(n9686), .ZN(
        P1_U3460) );
  OAI22_X1 U10777 ( .A1(n9642), .A2(n9680), .B1(n9641), .B2(n9678), .ZN(n9644)
         );
  AOI211_X1 U10778 ( .C1(n9677), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9690)
         );
  INV_X1 U10779 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9646) );
  AOI22_X1 U10780 ( .A1(n10017), .A2(n9690), .B1(n9646), .B2(n9686), .ZN(
        P1_U3463) );
  INV_X1 U10781 ( .A(n9647), .ZN(n9652) );
  OAI22_X1 U10782 ( .A1(n9649), .A2(n9680), .B1(n9648), .B2(n9678), .ZN(n9651)
         );
  AOI211_X1 U10783 ( .C1(n9677), .C2(n9652), .A(n9651), .B(n9650), .ZN(n9691)
         );
  INV_X1 U10784 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9653) );
  AOI22_X1 U10785 ( .A1(n10017), .A2(n9691), .B1(n9653), .B2(n9686), .ZN(
        P1_U3466) );
  OAI21_X1 U10786 ( .B1(n9655), .B2(n9678), .A(n9654), .ZN(n9657) );
  AOI211_X1 U10787 ( .C1(n9684), .C2(n9658), .A(n9657), .B(n9656), .ZN(n9692)
         );
  INV_X1 U10788 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U10789 ( .A1(n10017), .A2(n9692), .B1(n9659), .B2(n9686), .ZN(
        P1_U3469) );
  OAI22_X1 U10790 ( .A1(n9661), .A2(n9680), .B1(n9660), .B2(n9678), .ZN(n9663)
         );
  AOI211_X1 U10791 ( .C1(n9677), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9693)
         );
  INV_X1 U10792 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9665) );
  AOI22_X1 U10793 ( .A1(n10017), .A2(n9693), .B1(n9665), .B2(n9686), .ZN(
        P1_U3472) );
  OAI211_X1 U10794 ( .C1(n9668), .C2(n9678), .A(n9667), .B(n9666), .ZN(n9669)
         );
  AOI21_X1 U10795 ( .B1(n9684), .B2(n9670), .A(n9669), .ZN(n9695) );
  INV_X1 U10796 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9671) );
  AOI22_X1 U10797 ( .A1(n10017), .A2(n9695), .B1(n9671), .B2(n9686), .ZN(
        P1_U3475) );
  OAI22_X1 U10798 ( .A1(n9673), .A2(n9680), .B1(n9672), .B2(n9678), .ZN(n9675)
         );
  AOI211_X1 U10799 ( .C1(n9677), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9696)
         );
  INV_X1 U10800 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9927) );
  AOI22_X1 U10801 ( .A1(n10017), .A2(n9696), .B1(n9927), .B2(n9686), .ZN(
        P1_U3478) );
  OAI22_X1 U10802 ( .A1(n9681), .A2(n9680), .B1(n9679), .B2(n9678), .ZN(n9683)
         );
  AOI211_X1 U10803 ( .C1(n9685), .C2(n9684), .A(n9683), .B(n9682), .ZN(n9698)
         );
  INV_X1 U10804 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9687) );
  AOI22_X1 U10805 ( .A1(n10017), .A2(n9698), .B1(n9687), .B2(n9686), .ZN(
        P1_U3481) );
  AOI22_X1 U10806 ( .A1(n4269), .A2(n9689), .B1(n9688), .B2(n9697), .ZN(
        P1_U3525) );
  AOI22_X1 U10807 ( .A1(n4269), .A2(n9690), .B1(n5182), .B2(n9697), .ZN(
        P1_U3526) );
  AOI22_X1 U10808 ( .A1(n4269), .A2(n9691), .B1(n5183), .B2(n9697), .ZN(
        P1_U3527) );
  AOI22_X1 U10809 ( .A1(n4269), .A2(n9692), .B1(n5180), .B2(n9697), .ZN(
        P1_U3528) );
  AOI22_X1 U10810 ( .A1(n4269), .A2(n9693), .B1(n5186), .B2(n9697), .ZN(
        P1_U3529) );
  AOI22_X1 U10811 ( .A1(n4269), .A2(n9695), .B1(n9694), .B2(n9697), .ZN(
        P1_U3530) );
  AOI22_X1 U10812 ( .A1(n4269), .A2(n9696), .B1(n5286), .B2(n9697), .ZN(
        P1_U3531) );
  AOI22_X1 U10813 ( .A1(n4269), .A2(n9698), .B1(n5287), .B2(n9697), .ZN(
        P1_U3532) );
  XOR2_X1 U10814 ( .A(n9700), .B(n9699), .Z(n9707) );
  OAI21_X1 U10815 ( .B1(n9714), .B2(n9702), .A(n9701), .ZN(n9703) );
  AOI21_X1 U10816 ( .B1(n9717), .B2(n9704), .A(n9703), .ZN(n9705) );
  OAI21_X1 U10817 ( .B1(n4540), .B2(n9731), .A(n9705), .ZN(n9706) );
  AOI21_X1 U10818 ( .B1(n9707), .B2(n9733), .A(n9706), .ZN(n9708) );
  OAI21_X1 U10819 ( .B1(n9737), .B2(n9709), .A(n9708), .ZN(P2_U3219) );
  XOR2_X1 U10820 ( .A(n9710), .B(n9711), .Z(n9721) );
  OAI21_X1 U10821 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9715) );
  AOI21_X1 U10822 ( .B1(n9717), .B2(n9716), .A(n9715), .ZN(n9718) );
  OAI21_X1 U10823 ( .B1(n9719), .B2(n9731), .A(n9718), .ZN(n9720) );
  AOI21_X1 U10824 ( .B1(n9721), .B2(n9733), .A(n9720), .ZN(n9722) );
  OAI21_X1 U10825 ( .B1(n9737), .B2(n9723), .A(n9722), .ZN(P2_U3223) );
  OAI21_X1 U10826 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(n9734) );
  AOI21_X1 U10827 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9730) );
  OAI21_X1 U10828 ( .B1(n9790), .B2(n9731), .A(n9730), .ZN(n9732) );
  AOI21_X1 U10829 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9735) );
  OAI21_X1 U10830 ( .B1(n9737), .B2(n9736), .A(n9735), .ZN(P2_U3229) );
  AOI21_X1 U10831 ( .B1(n9749), .B2(P2_REG2_REG_0__SCAN_IN), .A(n9738), .ZN(
        n9746) );
  OAI21_X1 U10832 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n9740), .A(n9739), .ZN(
        n9741) );
  AOI21_X1 U10833 ( .B1(n9749), .B2(n9742), .A(n9741), .ZN(n9744) );
  AOI22_X1 U10834 ( .A1(n9747), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9743) );
  OAI221_X1 U10835 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9746), .C1(n9745), .C2(
        n9744), .A(n9743), .ZN(P2_U3245) );
  AOI22_X1 U10836 ( .A1(n9747), .A2(P2_ADDR_REG_7__SCAN_IN), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(P2_U3152), .ZN(n9761) );
  OAI211_X1 U10837 ( .C1(n9751), .C2(n9750), .A(n9749), .B(n9748), .ZN(n9760)
         );
  OAI211_X1 U10838 ( .C1(n9755), .C2(n9754), .A(n9753), .B(n9752), .ZN(n9759)
         );
  NAND2_X1 U10839 ( .A1(n9757), .A2(n9756), .ZN(n9758) );
  NAND4_X1 U10840 ( .A1(n9761), .A2(n9760), .A3(n9759), .A4(n9758), .ZN(
        P2_U3252) );
  NOR2_X1 U10841 ( .A1(n9763), .A2(n9762), .ZN(n9764) );
  AND2_X1 U10842 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9767), .ZN(P2_U3297) );
  AND2_X1 U10843 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9767), .ZN(P2_U3298) );
  AND2_X1 U10844 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9767), .ZN(P2_U3299) );
  AND2_X1 U10845 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9767), .ZN(P2_U3300) );
  AND2_X1 U10846 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9767), .ZN(P2_U3301) );
  AND2_X1 U10847 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9767), .ZN(P2_U3302) );
  AND2_X1 U10848 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9767), .ZN(P2_U3303) );
  AND2_X1 U10849 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9767), .ZN(P2_U3304) );
  NOR2_X1 U10850 ( .A1(n9764), .A2(n9963), .ZN(P2_U3305) );
  AND2_X1 U10851 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9767), .ZN(P2_U3306) );
  AND2_X1 U10852 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9767), .ZN(P2_U3307) );
  AND2_X1 U10853 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9767), .ZN(P2_U3308) );
  AND2_X1 U10854 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9767), .ZN(P2_U3309) );
  AND2_X1 U10855 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9767), .ZN(P2_U3310) );
  AND2_X1 U10856 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9767), .ZN(P2_U3311) );
  AND2_X1 U10857 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9767), .ZN(P2_U3312) );
  AND2_X1 U10858 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9767), .ZN(P2_U3313) );
  AND2_X1 U10859 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9767), .ZN(P2_U3314) );
  AND2_X1 U10860 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9767), .ZN(P2_U3315) );
  AND2_X1 U10861 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9767), .ZN(P2_U3316) );
  AND2_X1 U10862 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9767), .ZN(P2_U3317) );
  NOR2_X1 U10863 ( .A1(n9764), .A2(n9983), .ZN(P2_U3318) );
  AND2_X1 U10864 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9767), .ZN(P2_U3319) );
  AND2_X1 U10865 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9767), .ZN(P2_U3320) );
  AND2_X1 U10866 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9767), .ZN(P2_U3321) );
  NOR2_X1 U10867 ( .A1(n9764), .A2(n9996), .ZN(P2_U3322) );
  NOR2_X1 U10868 ( .A1(n9764), .A2(n10003), .ZN(P2_U3323) );
  AND2_X1 U10869 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9767), .ZN(P2_U3324) );
  AND2_X1 U10870 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9767), .ZN(P2_U3325) );
  AND2_X1 U10871 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9767), .ZN(P2_U3326) );
  AOI22_X1 U10872 ( .A1(n9766), .A2(n9769), .B1(n9765), .B2(n9767), .ZN(
        P2_U3437) );
  AOI22_X1 U10873 ( .A1(n9770), .A2(n9769), .B1(n9768), .B2(n9767), .ZN(
        P2_U3438) );
  INV_X1 U10874 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9771) );
  AOI22_X1 U10875 ( .A1(n4267), .A2(n9772), .B1(n9771), .B2(n9825), .ZN(
        P2_U3451) );
  INV_X1 U10876 ( .A(n9773), .ZN(n9775) );
  OAI22_X1 U10877 ( .A1(n9775), .A2(n9781), .B1(n9774), .B2(n9820), .ZN(n9777)
         );
  AOI211_X1 U10878 ( .C1(n9823), .C2(n9778), .A(n9777), .B(n9776), .ZN(n9826)
         );
  INV_X1 U10879 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9779) );
  AOI22_X1 U10880 ( .A1(n4267), .A2(n9826), .B1(n9779), .B2(n9825), .ZN(
        P2_U3454) );
  OAI22_X1 U10881 ( .A1(n9782), .A2(n9781), .B1(n9780), .B2(n9820), .ZN(n9784)
         );
  AOI211_X1 U10882 ( .C1(n9786), .C2(n9785), .A(n9784), .B(n9783), .ZN(n9827)
         );
  INV_X1 U10883 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9787) );
  AOI22_X1 U10884 ( .A1(n4267), .A2(n9827), .B1(n9787), .B2(n9825), .ZN(
        P2_U3460) );
  OAI211_X1 U10885 ( .C1(n9790), .C2(n9820), .A(n9789), .B(n9788), .ZN(n9791)
         );
  AOI21_X1 U10886 ( .B1(n9823), .B2(n9792), .A(n9791), .ZN(n9829) );
  INV_X1 U10887 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9935) );
  AOI22_X1 U10888 ( .A1(n4267), .A2(n9829), .B1(n9935), .B2(n9825), .ZN(
        P2_U3466) );
  AOI22_X1 U10889 ( .A1(n9794), .A2(n9810), .B1(n9809), .B2(n9793), .ZN(n9795)
         );
  OAI211_X1 U10890 ( .C1(n9797), .C2(n9804), .A(n9796), .B(n9795), .ZN(n9798)
         );
  INV_X1 U10891 ( .A(n9798), .ZN(n9830) );
  INV_X1 U10892 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U10893 ( .A1(n4267), .A2(n9830), .B1(n9799), .B2(n9825), .ZN(
        P2_U3469) );
  AOI22_X1 U10894 ( .A1(n9801), .A2(n9810), .B1(n9809), .B2(n9800), .ZN(n9802)
         );
  OAI211_X1 U10895 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9806)
         );
  INV_X1 U10896 ( .A(n9806), .ZN(n9831) );
  INV_X1 U10897 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9807) );
  AOI22_X1 U10898 ( .A1(n4267), .A2(n9831), .B1(n9807), .B2(n9825), .ZN(
        P2_U3472) );
  AOI22_X1 U10899 ( .A1(n9811), .A2(n9810), .B1(n9809), .B2(n9808), .ZN(n9812)
         );
  OAI211_X1 U10900 ( .C1(n9815), .C2(n9814), .A(n9813), .B(n9812), .ZN(n9816)
         );
  INV_X1 U10901 ( .A(n9816), .ZN(n9832) );
  INV_X1 U10902 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9817) );
  AOI22_X1 U10903 ( .A1(n4267), .A2(n9832), .B1(n9817), .B2(n9825), .ZN(
        P2_U3478) );
  OAI211_X1 U10904 ( .C1(n9821), .C2(n9820), .A(n9819), .B(n9818), .ZN(n9822)
         );
  AOI21_X1 U10905 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9834) );
  INV_X1 U10906 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U10907 ( .A1(n4267), .A2(n9834), .B1(n9993), .B2(n9825), .ZN(
        P2_U3484) );
  AOI22_X1 U10908 ( .A1(n4268), .A2(n9826), .B1(n5205), .B2(n9833), .ZN(
        P2_U3521) );
  AOI22_X1 U10909 ( .A1(n4268), .A2(n9827), .B1(n5210), .B2(n9833), .ZN(
        P2_U3523) );
  AOI22_X1 U10910 ( .A1(n4268), .A2(n9829), .B1(n9828), .B2(n9833), .ZN(
        P2_U3525) );
  AOI22_X1 U10911 ( .A1(n4268), .A2(n9830), .B1(n5204), .B2(n9833), .ZN(
        P2_U3526) );
  AOI22_X1 U10912 ( .A1(n4268), .A2(n9831), .B1(n5203), .B2(n9833), .ZN(
        P2_U3527) );
  AOI22_X1 U10913 ( .A1(n4268), .A2(n9832), .B1(n5219), .B2(n9833), .ZN(
        P2_U3529) );
  AOI22_X1 U10914 ( .A1(n4268), .A2(n9834), .B1(n9952), .B2(n9833), .ZN(
        P2_U3531) );
  INV_X1 U10915 ( .A(n9835), .ZN(n9836) );
  NAND2_X1 U10916 ( .A1(n9837), .A2(n9836), .ZN(n9838) );
  XNOR2_X1 U10917 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9838), .ZN(ADD_1071_U5) );
  INV_X1 U10918 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U10919 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n9938), .B2(n5158), .ZN(ADD_1071_U46) );
  OAI21_X1 U10920 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(ADD_1071_U56) );
  OAI21_X1 U10921 ( .B1(n9844), .B2(n9843), .A(n9842), .ZN(ADD_1071_U57) );
  OAI21_X1 U10922 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(ADD_1071_U58) );
  OAI21_X1 U10923 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(ADD_1071_U59) );
  OAI21_X1 U10924 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(ADD_1071_U60) );
  OAI21_X1 U10925 ( .B1(n9856), .B2(n9855), .A(n9854), .ZN(ADD_1071_U61) );
  AOI21_X1 U10926 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(ADD_1071_U62) );
  AOI21_X1 U10927 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(ADD_1071_U63) );
  NAND4_X1 U10928 ( .A1(keyinput38), .A2(keyinput50), .A3(keyinput35), .A4(
        keyinput22), .ZN(n9867) );
  NAND3_X1 U10929 ( .A1(keyinput20), .A2(keyinput60), .A3(keyinput17), .ZN(
        n9866) );
  NOR2_X1 U10930 ( .A1(keyinput57), .A2(keyinput23), .ZN(n9864) );
  NOR4_X1 U10931 ( .A1(keyinput54), .A2(keyinput28), .A3(keyinput36), .A4(
        keyinput32), .ZN(n9863) );
  NAND4_X1 U10932 ( .A1(keyinput46), .A2(keyinput55), .A3(n9864), .A4(n9863), 
        .ZN(n9865) );
  NOR4_X1 U10933 ( .A1(keyinput51), .A2(n9867), .A3(n9866), .A4(n9865), .ZN(
        n10014) );
  NOR2_X1 U10934 ( .A1(keyinput4), .A2(keyinput24), .ZN(n9874) );
  NAND2_X1 U10935 ( .A1(keyinput11), .A2(keyinput47), .ZN(n9872) );
  NOR3_X1 U10936 ( .A1(keyinput14), .A2(keyinput48), .A3(keyinput56), .ZN(
        n9870) );
  INV_X1 U10937 ( .A(keyinput29), .ZN(n9868) );
  NOR3_X1 U10938 ( .A1(keyinput49), .A2(keyinput21), .A3(n9868), .ZN(n9869) );
  NAND4_X1 U10939 ( .A1(keyinput34), .A2(n9870), .A3(keyinput40), .A4(n9869), 
        .ZN(n9871) );
  NOR4_X1 U10940 ( .A1(keyinput8), .A2(keyinput58), .A3(n9872), .A4(n9871), 
        .ZN(n9873) );
  NAND4_X1 U10941 ( .A1(keyinput44), .A2(keyinput37), .A3(n9874), .A4(n9873), 
        .ZN(n9889) );
  NOR3_X1 U10942 ( .A1(keyinput41), .A2(keyinput31), .A3(keyinput26), .ZN(
        n9876) );
  NOR3_X1 U10943 ( .A1(keyinput7), .A2(keyinput5), .A3(keyinput33), .ZN(n9875)
         );
  NAND4_X1 U10944 ( .A1(keyinput18), .A2(n9876), .A3(keyinput19), .A4(n9875), 
        .ZN(n9888) );
  NOR3_X1 U10945 ( .A1(keyinput39), .A2(keyinput25), .A3(keyinput12), .ZN(
        n9878) );
  NOR4_X1 U10946 ( .A1(keyinput62), .A2(keyinput10), .A3(keyinput15), .A4(
        keyinput42), .ZN(n9877) );
  NAND3_X1 U10947 ( .A1(keyinput16), .A2(n9878), .A3(n9877), .ZN(n9887) );
  NAND2_X1 U10948 ( .A1(keyinput53), .A2(keyinput3), .ZN(n9879) );
  NOR3_X1 U10949 ( .A1(keyinput0), .A2(keyinput27), .A3(n9879), .ZN(n9885) );
  NOR3_X1 U10950 ( .A1(keyinput6), .A2(keyinput59), .A3(keyinput2), .ZN(n9884)
         );
  NAND3_X1 U10951 ( .A1(keyinput45), .A2(keyinput52), .A3(keyinput61), .ZN(
        n9882) );
  INV_X1 U10952 ( .A(keyinput30), .ZN(n9880) );
  NAND3_X1 U10953 ( .A1(keyinput1), .A2(keyinput9), .A3(n9880), .ZN(n9881) );
  NOR4_X1 U10954 ( .A1(keyinput63), .A2(keyinput43), .A3(n9882), .A4(n9881), 
        .ZN(n9883) );
  NAND4_X1 U10955 ( .A1(n9885), .A2(keyinput13), .A3(n9884), .A4(n9883), .ZN(
        n9886) );
  NOR4_X1 U10956 ( .A1(n9889), .A2(n9888), .A3(n9887), .A4(n9886), .ZN(n10013)
         );
  AOI22_X1 U10957 ( .A1(n9892), .A2(keyinput34), .B1(keyinput14), .B2(n9891), 
        .ZN(n9890) );
  OAI221_X1 U10958 ( .B1(n9892), .B2(keyinput34), .C1(n9891), .C2(keyinput14), 
        .A(n9890), .ZN(n9903) );
  INV_X1 U10959 ( .A(SI_29_), .ZN(n9894) );
  AOI22_X1 U10960 ( .A1(n9894), .A2(keyinput48), .B1(n4971), .B2(keyinput56), 
        .ZN(n9893) );
  OAI221_X1 U10961 ( .B1(n9894), .B2(keyinput48), .C1(n4971), .C2(keyinput56), 
        .A(n9893), .ZN(n9902) );
  AOI22_X1 U10962 ( .A1(n9897), .A2(keyinput44), .B1(keyinput4), .B2(n9896), 
        .ZN(n9895) );
  OAI221_X1 U10963 ( .B1(n9897), .B2(keyinput44), .C1(n9896), .C2(keyinput4), 
        .A(n9895), .ZN(n9901) );
  XNOR2_X1 U10964 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput24), .ZN(n9899) );
  XNOR2_X1 U10965 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput37), .ZN(n9898)
         );
  NAND2_X1 U10966 ( .A1(n9899), .A2(n9898), .ZN(n9900) );
  NOR4_X1 U10967 ( .A1(n9903), .A2(n9902), .A3(n9901), .A4(n9900), .ZN(n9949)
         );
  AOI22_X1 U10968 ( .A1(n9905), .A2(keyinput49), .B1(keyinput21), .B2(n5253), 
        .ZN(n9904) );
  OAI221_X1 U10969 ( .B1(n9905), .B2(keyinput49), .C1(n5253), .C2(keyinput21), 
        .A(n9904), .ZN(n9918) );
  AOI22_X1 U10970 ( .A1(n9908), .A2(keyinput8), .B1(keyinput58), .B2(n9907), 
        .ZN(n9906) );
  OAI221_X1 U10971 ( .B1(n9908), .B2(keyinput8), .C1(n9907), .C2(keyinput58), 
        .A(n9906), .ZN(n9917) );
  INV_X1 U10972 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U10973 ( .A1(n9911), .A2(keyinput40), .B1(n9910), .B2(keyinput29), 
        .ZN(n9909) );
  OAI221_X1 U10974 ( .B1(n9911), .B2(keyinput40), .C1(n9910), .C2(keyinput29), 
        .A(n9909), .ZN(n9916) );
  INV_X1 U10975 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9912) );
  XOR2_X1 U10976 ( .A(n9912), .B(keyinput47), .Z(n9914) );
  XNOR2_X1 U10977 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput11), .ZN(n9913) );
  NAND2_X1 U10978 ( .A1(n9914), .A2(n9913), .ZN(n9915) );
  NOR4_X1 U10979 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(n9948)
         );
  AOI22_X1 U10980 ( .A1(n9920), .A2(keyinput39), .B1(keyinput25), .B2(n7528), 
        .ZN(n9919) );
  OAI221_X1 U10981 ( .B1(n9920), .B2(keyinput39), .C1(n7528), .C2(keyinput25), 
        .A(n9919), .ZN(n9931) );
  INV_X1 U10982 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9922) );
  AOI22_X1 U10983 ( .A1(n9923), .A2(keyinput16), .B1(keyinput12), .B2(n9922), 
        .ZN(n9921) );
  OAI221_X1 U10984 ( .B1(n9923), .B2(keyinput16), .C1(n9922), .C2(keyinput12), 
        .A(n9921), .ZN(n9930) );
  AOI22_X1 U10985 ( .A1(n4984), .A2(keyinput62), .B1(n9925), .B2(keyinput10), 
        .ZN(n9924) );
  OAI221_X1 U10986 ( .B1(n4984), .B2(keyinput62), .C1(n9925), .C2(keyinput10), 
        .A(n9924), .ZN(n9929) );
  AOI22_X1 U10987 ( .A1(n9927), .A2(keyinput15), .B1(keyinput42), .B2(n8391), 
        .ZN(n9926) );
  OAI221_X1 U10988 ( .B1(n9927), .B2(keyinput15), .C1(n8391), .C2(keyinput42), 
        .A(n9926), .ZN(n9928) );
  NOR4_X1 U10989 ( .A1(n9931), .A2(n9930), .A3(n9929), .A4(n9928), .ZN(n9947)
         );
  INV_X1 U10990 ( .A(keyinput18), .ZN(n9933) );
  AOI22_X1 U10991 ( .A1(n5210), .A2(keyinput41), .B1(SI_31_), .B2(n9933), .ZN(
        n9932) );
  OAI221_X1 U10992 ( .B1(n5210), .B2(keyinput41), .C1(n9933), .C2(SI_31_), .A(
        n9932), .ZN(n9945) );
  AOI22_X1 U10993 ( .A1(n9935), .A2(keyinput31), .B1(n7833), .B2(keyinput26), 
        .ZN(n9934) );
  OAI221_X1 U10994 ( .B1(n9935), .B2(keyinput31), .C1(n7833), .C2(keyinput26), 
        .A(n9934), .ZN(n9944) );
  AOI22_X1 U10995 ( .A1(n9938), .A2(keyinput7), .B1(n9937), .B2(keyinput19), 
        .ZN(n9936) );
  OAI221_X1 U10996 ( .B1(n9938), .B2(keyinput7), .C1(n9937), .C2(keyinput19), 
        .A(n9936), .ZN(n9943) );
  AOI22_X1 U10997 ( .A1(n9941), .A2(keyinput5), .B1(keyinput33), .B2(n9940), 
        .ZN(n9939) );
  OAI221_X1 U10998 ( .B1(n9941), .B2(keyinput5), .C1(n9940), .C2(keyinput33), 
        .A(n9939), .ZN(n9942) );
  NOR4_X1 U10999 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(n9946)
         );
  NAND4_X1 U11000 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(n10012) );
  AOI22_X1 U11001 ( .A1(n9952), .A2(keyinput60), .B1(n9951), .B2(keyinput17), 
        .ZN(n9950) );
  OAI221_X1 U11002 ( .B1(n9952), .B2(keyinput60), .C1(n9951), .C2(keyinput17), 
        .A(n9950), .ZN(n9961) );
  AOI22_X1 U11003 ( .A1(n4907), .A2(keyinput20), .B1(keyinput51), .B2(n9954), 
        .ZN(n9953) );
  OAI221_X1 U11004 ( .B1(n4907), .B2(keyinput20), .C1(n9954), .C2(keyinput51), 
        .A(n9953), .ZN(n9960) );
  INV_X1 U11005 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U11006 ( .A1(n5287), .A2(keyinput36), .B1(keyinput32), .B2(n9956), 
        .ZN(n9955) );
  OAI221_X1 U11007 ( .B1(n5287), .B2(keyinput36), .C1(n9956), .C2(keyinput32), 
        .A(n9955), .ZN(n9959) );
  AOI22_X1 U11008 ( .A1(n5015), .A2(keyinput54), .B1(n5023), .B2(keyinput28), 
        .ZN(n9957) );
  OAI221_X1 U11009 ( .B1(n5015), .B2(keyinput54), .C1(n5023), .C2(keyinput28), 
        .A(n9957), .ZN(n9958) );
  NOR4_X1 U11010 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n10010)
         );
  AOI22_X1 U11011 ( .A1(n9964), .A2(keyinput55), .B1(n9963), .B2(keyinput23), 
        .ZN(n9962) );
  OAI221_X1 U11012 ( .B1(n9964), .B2(keyinput55), .C1(n9963), .C2(keyinput23), 
        .A(n9962), .ZN(n9976) );
  AOI22_X1 U11013 ( .A1(n9967), .A2(keyinput35), .B1(n9966), .B2(keyinput22), 
        .ZN(n9965) );
  OAI221_X1 U11014 ( .B1(n9967), .B2(keyinput35), .C1(n9966), .C2(keyinput22), 
        .A(n9965), .ZN(n9975) );
  AOI22_X1 U11015 ( .A1(n9970), .A2(keyinput38), .B1(keyinput50), .B2(n9969), 
        .ZN(n9968) );
  OAI221_X1 U11016 ( .B1(n9970), .B2(keyinput38), .C1(n9969), .C2(keyinput50), 
        .A(n9968), .ZN(n9974) );
  XNOR2_X1 U11017 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput57), .ZN(n9972) );
  XNOR2_X1 U11018 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput46), .ZN(n9971) );
  NAND2_X1 U11019 ( .A1(n9972), .A2(n9971), .ZN(n9973) );
  NOR4_X1 U11020 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), .ZN(n10009)
         );
  AOI22_X1 U11021 ( .A1(n9979), .A2(keyinput30), .B1(n9978), .B2(keyinput9), 
        .ZN(n9977) );
  OAI221_X1 U11022 ( .B1(n9979), .B2(keyinput30), .C1(n9978), .C2(keyinput9), 
        .A(n9977), .ZN(n9991) );
  AOI22_X1 U11023 ( .A1(n5186), .A2(keyinput43), .B1(keyinput1), .B2(n9981), 
        .ZN(n9980) );
  OAI221_X1 U11024 ( .B1(n5186), .B2(keyinput43), .C1(n9981), .C2(keyinput1), 
        .A(n9980), .ZN(n9990) );
  AOI22_X1 U11025 ( .A1(n9984), .A2(keyinput2), .B1(n9983), .B2(keyinput13), 
        .ZN(n9982) );
  OAI221_X1 U11026 ( .B1(n9984), .B2(keyinput2), .C1(n9983), .C2(keyinput13), 
        .A(n9982), .ZN(n9989) );
  AOI22_X1 U11027 ( .A1(n9987), .A2(keyinput6), .B1(n9986), .B2(keyinput59), 
        .ZN(n9985) );
  OAI221_X1 U11028 ( .B1(n9987), .B2(keyinput6), .C1(n9986), .C2(keyinput59), 
        .A(n9985), .ZN(n9988) );
  NOR4_X1 U11029 ( .A1(n9991), .A2(n9990), .A3(n9989), .A4(n9988), .ZN(n10008)
         );
  AOI22_X1 U11030 ( .A1(n9994), .A2(keyinput45), .B1(n9993), .B2(keyinput52), 
        .ZN(n9992) );
  OAI221_X1 U11031 ( .B1(n9994), .B2(keyinput45), .C1(n9993), .C2(keyinput52), 
        .A(n9992), .ZN(n9999) );
  XNOR2_X1 U11032 ( .A(n9995), .B(keyinput63), .ZN(n9998) );
  XNOR2_X1 U11033 ( .A(n9996), .B(keyinput61), .ZN(n9997) );
  OR3_X1 U11034 ( .A1(n9999), .A2(n9998), .A3(n9997), .ZN(n10006) );
  AOI22_X1 U11035 ( .A1(n10001), .A2(keyinput53), .B1(keyinput3), .B2(n5225), 
        .ZN(n10000) );
  OAI221_X1 U11036 ( .B1(n10001), .B2(keyinput53), .C1(n5225), .C2(keyinput3), 
        .A(n10000), .ZN(n10005) );
  AOI22_X1 U11037 ( .A1(n10003), .A2(keyinput0), .B1(keyinput27), .B2(n5515), 
        .ZN(n10002) );
  OAI221_X1 U11038 ( .B1(n10003), .B2(keyinput0), .C1(n5515), .C2(keyinput27), 
        .A(n10002), .ZN(n10004) );
  NOR3_X1 U11039 ( .A1(n10006), .A2(n10005), .A3(n10004), .ZN(n10007) );
  NAND4_X1 U11040 ( .A1(n10010), .A2(n10009), .A3(n10008), .A4(n10007), .ZN(
        n10011) );
  AOI211_X1 U11041 ( .C1(n10014), .C2(n10013), .A(n10012), .B(n10011), .ZN(
        n10019) );
  NAND2_X1 U11042 ( .A1(n10015), .A2(n10017), .ZN(n10016) );
  OAI21_X1 U11043 ( .B1(P1_REG0_REG_1__SCAN_IN), .B2(n10017), .A(n10016), .ZN(
        n10018) );
  XNOR2_X1 U11044 ( .A(n10019), .B(n10018), .ZN(P1_U3457) );
  XOR2_X1 U11045 ( .A(n10020), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11046 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  XOR2_X1 U11047 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10023), .Z(ADD_1071_U51) );
  OAI21_X1 U11048 ( .B1(n10026), .B2(n10025), .A(n10024), .ZN(n10027) );
  XNOR2_X1 U11049 ( .A(n10027), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11050 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(ADD_1071_U47) );
  AOI21_X1 U11051 ( .B1(n5253), .B2(n10032), .A(n10031), .ZN(ADD_1071_U48) );
  XOR2_X1 U11052 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10033), .Z(ADD_1071_U49) );
  XOR2_X1 U11053 ( .A(n10035), .B(n10034), .Z(ADD_1071_U54) );
  XOR2_X1 U11054 ( .A(n10037), .B(n10036), .Z(ADD_1071_U53) );
  XNOR2_X1 U11055 ( .A(n10039), .B(n10038), .ZN(ADD_1071_U52) );
  NAND2_X1 U9380 ( .A1(n7819), .A2(n7818), .ZN(n8640) );
  CLKBUF_X1 U4777 ( .A(n6561), .Z(n7995) );
  CLKBUF_X1 U4779 ( .A(n5750), .Z(n8043) );
  CLKBUF_X1 U4783 ( .A(n7320), .Z(n7525) );
  AND2_X1 U6077 ( .A1(n7422), .A2(n7421), .ZN(n10043) );
endmodule

